magic
tech sky130A
timestamp 1713605288
<< pwell >>
rect -200 -165 6570 12000
<< psubdiff >>
rect -152 11920 -140 11940
rect 6500 11920 6512 11940
rect -185 11870 -165 11885
rect -185 -50 -165 -35
rect -152 -105 -140 -85
rect 6500 -105 6512 -85
<< psubdiffcont >>
rect -140 11920 6500 11940
rect -185 -35 -165 11870
rect -140 -105 6500 -85
<< locali >>
rect -115 12065 -85 12085
rect -110 11940 -90 12065
rect 6485 12040 6515 12060
rect 6490 11940 6510 12040
rect -185 11870 -165 11940
rect -148 11920 -140 11940
rect 6500 11930 6510 11940
rect 6500 11920 6508 11930
rect -185 -70 -165 -35
rect -148 -105 -140 -85
rect 6500 -105 6508 -85
<< viali >>
rect -135 12065 -115 12085
rect -85 12065 -65 12085
rect 6465 12040 6485 12060
rect 6515 12040 6535 12060
rect -135 11920 6455 11940
rect -185 -25 -165 11870
rect -110 -105 6480 -85
<< metal1 >>
rect -145 12060 -140 12090
rect -195 11950 -190 11980
rect -160 11950 -155 11980
rect -195 11940 -155 11950
rect -110 11943 -90 12090
rect -60 12060 -55 12090
rect 6455 12035 6460 12065
rect 5 11950 10 11980
rect 40 11950 45 11980
rect 5 11943 45 11950
rect 205 11950 210 11980
rect 240 11950 245 11980
rect 205 11943 245 11950
rect 405 11950 410 11980
rect 440 11950 445 11980
rect 405 11943 445 11950
rect 605 11950 610 11980
rect 640 11950 645 11980
rect 605 11943 645 11950
rect 805 11950 810 11980
rect 840 11950 845 11980
rect 805 11943 845 11950
rect 1005 11950 1010 11980
rect 1040 11950 1045 11980
rect 1005 11943 1045 11950
rect 1205 11950 1210 11980
rect 1240 11950 1245 11980
rect 1205 11943 1245 11950
rect 1405 11950 1410 11980
rect 1440 11950 1445 11980
rect 1405 11943 1445 11950
rect 1605 11950 1610 11980
rect 1640 11950 1645 11980
rect 1605 11943 1645 11950
rect 1805 11950 1810 11980
rect 1840 11950 1845 11980
rect 1805 11943 1845 11950
rect 2005 11950 2010 11980
rect 2040 11950 2045 11980
rect 2005 11943 2045 11950
rect 2205 11950 2210 11980
rect 2240 11950 2245 11980
rect 2205 11943 2245 11950
rect 2405 11950 2410 11980
rect 2440 11950 2445 11980
rect 2405 11943 2445 11950
rect 2605 11950 2610 11980
rect 2640 11950 2645 11980
rect 2605 11943 2645 11950
rect 2805 11950 2810 11980
rect 2840 11950 2845 11980
rect 2805 11943 2845 11950
rect 3005 11950 3010 11980
rect 3040 11950 3045 11980
rect 3005 11943 3045 11950
rect 3205 11950 3210 11980
rect 3240 11950 3245 11980
rect 3205 11943 3245 11950
rect 3405 11950 3410 11980
rect 3440 11950 3445 11980
rect 3405 11943 3445 11950
rect 3605 11950 3610 11980
rect 3640 11950 3645 11980
rect 3605 11943 3645 11950
rect 3805 11950 3810 11980
rect 3840 11950 3845 11980
rect 3805 11943 3845 11950
rect 4005 11950 4010 11980
rect 4040 11950 4045 11980
rect 4005 11943 4045 11950
rect 4205 11950 4210 11980
rect 4240 11950 4245 11980
rect 4205 11943 4245 11950
rect 4405 11950 4410 11980
rect 4440 11950 4445 11980
rect 4405 11943 4445 11950
rect 4605 11950 4610 11980
rect 4640 11950 4645 11980
rect 4605 11943 4645 11950
rect 4805 11950 4810 11980
rect 4840 11950 4845 11980
rect 4805 11943 4845 11950
rect 5005 11950 5010 11980
rect 5040 11950 5045 11980
rect 5005 11943 5045 11950
rect 5205 11950 5210 11980
rect 5240 11950 5245 11980
rect 5205 11943 5245 11950
rect 5405 11950 5410 11980
rect 5440 11950 5445 11980
rect 5405 11943 5445 11950
rect 5605 11950 5610 11980
rect 5640 11950 5645 11980
rect 5605 11943 5645 11950
rect 5805 11950 5810 11980
rect 5840 11950 5845 11980
rect 5805 11943 5845 11950
rect 6005 11950 6010 11980
rect 6040 11950 6045 11980
rect 6005 11943 6045 11950
rect 6205 11950 6210 11980
rect 6240 11950 6245 11980
rect 6205 11943 6245 11950
rect 6405 11950 6410 11980
rect 6440 11950 6445 11980
rect 6405 11943 6445 11950
rect -141 11940 6461 11943
rect 6490 11940 6510 12065
rect 6540 12035 6545 12065
rect -195 11920 -135 11940
rect 6455 11920 6570 11940
rect -195 11910 -155 11920
rect -141 11917 6461 11920
rect -195 11880 -190 11910
rect -160 11880 -155 11910
rect 5 11910 45 11917
rect 5 11880 10 11910
rect 40 11880 45 11910
rect 205 11910 245 11917
rect 205 11880 210 11910
rect 240 11880 245 11910
rect 405 11910 445 11917
rect 405 11880 410 11910
rect 440 11880 445 11910
rect 605 11910 645 11917
rect 605 11880 610 11910
rect 640 11880 645 11910
rect 805 11910 845 11917
rect 805 11880 810 11910
rect 840 11880 845 11910
rect 1005 11910 1045 11917
rect 1005 11880 1010 11910
rect 1040 11880 1045 11910
rect 1205 11910 1245 11917
rect 1205 11880 1210 11910
rect 1240 11880 1245 11910
rect 1405 11910 1445 11917
rect 1405 11880 1410 11910
rect 1440 11880 1445 11910
rect 1605 11910 1645 11917
rect 1605 11880 1610 11910
rect 1640 11880 1645 11910
rect 1805 11910 1845 11917
rect 1805 11880 1810 11910
rect 1840 11880 1845 11910
rect 2005 11910 2045 11917
rect 2005 11880 2010 11910
rect 2040 11880 2045 11910
rect 2205 11910 2245 11917
rect 2205 11880 2210 11910
rect 2240 11880 2245 11910
rect 2405 11910 2445 11917
rect 2405 11880 2410 11910
rect 2440 11880 2445 11910
rect 2605 11910 2645 11917
rect 2605 11880 2610 11910
rect 2640 11880 2645 11910
rect 2805 11910 2845 11917
rect 2805 11880 2810 11910
rect 2840 11880 2845 11910
rect 3005 11910 3045 11917
rect 3005 11880 3010 11910
rect 3040 11880 3045 11910
rect 3205 11910 3245 11917
rect 3205 11880 3210 11910
rect 3240 11880 3245 11910
rect 3405 11910 3445 11917
rect 3405 11880 3410 11910
rect 3440 11880 3445 11910
rect 3605 11910 3645 11917
rect 3605 11880 3610 11910
rect 3640 11880 3645 11910
rect 3805 11910 3845 11917
rect 3805 11880 3810 11910
rect 3840 11880 3845 11910
rect 4005 11910 4045 11917
rect 4005 11880 4010 11910
rect 4040 11880 4045 11910
rect 4205 11910 4245 11917
rect 4205 11880 4210 11910
rect 4240 11880 4245 11910
rect 4405 11910 4445 11917
rect 4405 11880 4410 11910
rect 4440 11880 4445 11910
rect 4605 11910 4645 11917
rect 4605 11880 4610 11910
rect 4640 11880 4645 11910
rect 4805 11910 4845 11917
rect 4805 11880 4810 11910
rect 4840 11880 4845 11910
rect 5005 11910 5045 11917
rect 5005 11880 5010 11910
rect 5040 11880 5045 11910
rect 5205 11910 5245 11917
rect 5205 11880 5210 11910
rect 5240 11880 5245 11910
rect 5405 11910 5445 11917
rect 5405 11880 5410 11910
rect 5440 11880 5445 11910
rect 5605 11910 5645 11917
rect 5605 11880 5610 11910
rect 5640 11880 5645 11910
rect 5805 11910 5845 11917
rect 5805 11880 5810 11910
rect 5840 11880 5845 11910
rect 6005 11910 6045 11917
rect 6005 11880 6010 11910
rect 6040 11880 6045 11910
rect 6205 11910 6245 11917
rect 6205 11880 6210 11910
rect 6240 11880 6245 11910
rect 6405 11910 6445 11917
rect 6405 11880 6410 11910
rect 6440 11880 6445 11910
rect -188 11870 -162 11880
rect -188 11795 -185 11870
rect -165 11795 -162 11870
rect -195 11765 -190 11795
rect -160 11765 -155 11795
rect -195 11725 -185 11765
rect -165 11755 -155 11765
rect 5 11765 10 11795
rect 40 11765 45 11795
rect 5 11755 45 11765
rect 205 11765 210 11795
rect 240 11765 245 11795
rect 205 11755 245 11765
rect 405 11765 410 11795
rect 440 11765 445 11795
rect 405 11755 445 11765
rect 605 11765 610 11795
rect 640 11765 645 11795
rect 605 11755 645 11765
rect 805 11765 810 11795
rect 840 11765 845 11795
rect 805 11755 845 11765
rect 1005 11765 1010 11795
rect 1040 11765 1045 11795
rect 1005 11755 1045 11765
rect 1205 11765 1210 11795
rect 1240 11765 1245 11795
rect 1205 11755 1245 11765
rect 1405 11765 1410 11795
rect 1440 11765 1445 11795
rect 1405 11755 1445 11765
rect 1605 11765 1610 11795
rect 1640 11765 1645 11795
rect 1605 11755 1645 11765
rect 1805 11765 1810 11795
rect 1840 11765 1845 11795
rect 1805 11755 1845 11765
rect 2005 11765 2010 11795
rect 2040 11765 2045 11795
rect 2005 11755 2045 11765
rect 2205 11765 2210 11795
rect 2240 11765 2245 11795
rect 2205 11755 2245 11765
rect 2405 11765 2410 11795
rect 2440 11765 2445 11795
rect 2405 11755 2445 11765
rect 2605 11765 2610 11795
rect 2640 11765 2645 11795
rect 2605 11755 2645 11765
rect 2805 11765 2810 11795
rect 2840 11765 2845 11795
rect 2805 11755 2845 11765
rect 3005 11765 3010 11795
rect 3040 11765 3045 11795
rect 3005 11755 3045 11765
rect 3205 11765 3210 11795
rect 3240 11765 3245 11795
rect 3205 11755 3245 11765
rect 3405 11765 3410 11795
rect 3440 11765 3445 11795
rect 3405 11755 3445 11765
rect 3605 11765 3610 11795
rect 3640 11765 3645 11795
rect 3605 11755 3645 11765
rect 3805 11765 3810 11795
rect 3840 11765 3845 11795
rect 3805 11755 3845 11765
rect 4005 11765 4010 11795
rect 4040 11765 4045 11795
rect 4005 11755 4045 11765
rect 4205 11765 4210 11795
rect 4240 11765 4245 11795
rect 4205 11755 4245 11765
rect 4405 11765 4410 11795
rect 4440 11765 4445 11795
rect 4405 11755 4445 11765
rect 4605 11765 4610 11795
rect 4640 11765 4645 11795
rect 4605 11755 4645 11765
rect 4805 11765 4810 11795
rect 4840 11765 4845 11795
rect 4805 11755 4845 11765
rect 5005 11765 5010 11795
rect 5040 11765 5045 11795
rect 5005 11755 5045 11765
rect 5205 11765 5210 11795
rect 5240 11765 5245 11795
rect 5205 11755 5245 11765
rect 5405 11765 5410 11795
rect 5440 11765 5445 11795
rect 5405 11755 5445 11765
rect 5605 11765 5610 11795
rect 5640 11765 5645 11795
rect 5605 11755 5645 11765
rect 5805 11765 5810 11795
rect 5840 11765 5845 11795
rect 5805 11755 5845 11765
rect 6005 11765 6010 11795
rect 6040 11765 6045 11795
rect 6005 11755 6045 11765
rect 6205 11765 6210 11795
rect 6240 11765 6245 11795
rect 6205 11755 6245 11765
rect 6405 11765 6410 11795
rect 6440 11765 6445 11795
rect 6405 11755 6445 11765
rect -165 11735 -30 11755
rect 5 11735 6570 11755
rect -165 11725 -155 11735
rect -195 11695 -190 11725
rect -160 11695 -155 11725
rect 5 11725 45 11735
rect 5 11695 10 11725
rect 40 11695 45 11725
rect 205 11725 245 11735
rect 205 11695 210 11725
rect 240 11695 245 11725
rect 405 11725 445 11735
rect 405 11695 410 11725
rect 440 11695 445 11725
rect 605 11725 645 11735
rect 605 11695 610 11725
rect 640 11695 645 11725
rect 805 11725 845 11735
rect 805 11695 810 11725
rect 840 11695 845 11725
rect 1005 11725 1045 11735
rect 1005 11695 1010 11725
rect 1040 11695 1045 11725
rect 1205 11725 1245 11735
rect 1205 11695 1210 11725
rect 1240 11695 1245 11725
rect 1405 11725 1445 11735
rect 1405 11695 1410 11725
rect 1440 11695 1445 11725
rect 1605 11725 1645 11735
rect 1605 11695 1610 11725
rect 1640 11695 1645 11725
rect 1805 11725 1845 11735
rect 1805 11695 1810 11725
rect 1840 11695 1845 11725
rect 2005 11725 2045 11735
rect 2005 11695 2010 11725
rect 2040 11695 2045 11725
rect 2205 11725 2245 11735
rect 2205 11695 2210 11725
rect 2240 11695 2245 11725
rect 2405 11725 2445 11735
rect 2405 11695 2410 11725
rect 2440 11695 2445 11725
rect 2605 11725 2645 11735
rect 2605 11695 2610 11725
rect 2640 11695 2645 11725
rect 2805 11725 2845 11735
rect 2805 11695 2810 11725
rect 2840 11695 2845 11725
rect 3005 11725 3045 11735
rect 3005 11695 3010 11725
rect 3040 11695 3045 11725
rect 3205 11725 3245 11735
rect 3205 11695 3210 11725
rect 3240 11695 3245 11725
rect 3405 11725 3445 11735
rect 3405 11695 3410 11725
rect 3440 11695 3445 11725
rect 3605 11725 3645 11735
rect 3605 11695 3610 11725
rect 3640 11695 3645 11725
rect 3805 11725 3845 11735
rect 3805 11695 3810 11725
rect 3840 11695 3845 11725
rect 4005 11725 4045 11735
rect 4005 11695 4010 11725
rect 4040 11695 4045 11725
rect 4205 11725 4245 11735
rect 4205 11695 4210 11725
rect 4240 11695 4245 11725
rect 4405 11725 4445 11735
rect 4405 11695 4410 11725
rect 4440 11695 4445 11725
rect 4605 11725 4645 11735
rect 4605 11695 4610 11725
rect 4640 11695 4645 11725
rect 4805 11725 4845 11735
rect 4805 11695 4810 11725
rect 4840 11695 4845 11725
rect 5005 11725 5045 11735
rect 5005 11695 5010 11725
rect 5040 11695 5045 11725
rect 5205 11725 5245 11735
rect 5205 11695 5210 11725
rect 5240 11695 5245 11725
rect 5405 11725 5445 11735
rect 5405 11695 5410 11725
rect 5440 11695 5445 11725
rect 5605 11725 5645 11735
rect 5605 11695 5610 11725
rect 5640 11695 5645 11725
rect 5805 11725 5845 11735
rect 5805 11695 5810 11725
rect 5840 11695 5845 11725
rect 6005 11725 6045 11735
rect 6005 11695 6010 11725
rect 6040 11695 6045 11725
rect 6205 11725 6245 11735
rect 6205 11695 6210 11725
rect 6240 11695 6245 11725
rect 6405 11725 6445 11735
rect 6405 11695 6410 11725
rect 6440 11695 6445 11725
rect -188 11610 -185 11695
rect -165 11610 -162 11695
rect 15 11610 35 11695
rect 215 11610 235 11695
rect 415 11610 435 11695
rect 615 11610 635 11695
rect 815 11610 835 11695
rect 1015 11610 1035 11695
rect 1215 11610 1235 11695
rect 1415 11610 1435 11695
rect 1615 11610 1635 11695
rect 1815 11610 1835 11695
rect 2015 11610 2035 11695
rect 2215 11610 2235 11695
rect 2415 11610 2435 11695
rect 2615 11610 2635 11695
rect 2815 11610 2835 11695
rect 3015 11610 3035 11695
rect 3215 11610 3235 11695
rect 3415 11610 3435 11695
rect 3615 11610 3635 11695
rect 3815 11610 3835 11695
rect 4015 11610 4035 11695
rect 4215 11610 4235 11695
rect 4415 11610 4435 11695
rect 4615 11610 4635 11695
rect 4815 11610 4835 11695
rect 5015 11610 5035 11695
rect 5215 11610 5235 11695
rect 5415 11610 5435 11695
rect 5615 11610 5635 11695
rect 5815 11610 5835 11695
rect 6015 11610 6035 11695
rect 6215 11610 6235 11695
rect -195 11580 -190 11610
rect -160 11580 -155 11610
rect -195 11540 -185 11580
rect -165 11570 -155 11580
rect 5 11580 10 11610
rect 40 11580 45 11610
rect 5 11570 45 11580
rect 205 11580 210 11610
rect 240 11580 245 11610
rect 205 11570 245 11580
rect 405 11580 410 11610
rect 440 11580 445 11610
rect 405 11570 445 11580
rect 605 11580 610 11610
rect 640 11580 645 11610
rect 605 11570 645 11580
rect 805 11580 810 11610
rect 840 11580 845 11610
rect 805 11570 845 11580
rect 1005 11580 1010 11610
rect 1040 11580 1045 11610
rect 1005 11570 1045 11580
rect 1205 11580 1210 11610
rect 1240 11580 1245 11610
rect 1205 11570 1245 11580
rect 1405 11580 1410 11610
rect 1440 11580 1445 11610
rect 1405 11570 1445 11580
rect 1605 11580 1610 11610
rect 1640 11580 1645 11610
rect 1605 11570 1645 11580
rect 1805 11580 1810 11610
rect 1840 11580 1845 11610
rect 1805 11570 1845 11580
rect 2005 11580 2010 11610
rect 2040 11580 2045 11610
rect 2005 11570 2045 11580
rect 2205 11580 2210 11610
rect 2240 11580 2245 11610
rect 2205 11570 2245 11580
rect 2405 11580 2410 11610
rect 2440 11580 2445 11610
rect 2405 11570 2445 11580
rect 2605 11580 2610 11610
rect 2640 11580 2645 11610
rect 2605 11570 2645 11580
rect 2805 11580 2810 11610
rect 2840 11580 2845 11610
rect 2805 11570 2845 11580
rect 3005 11580 3010 11610
rect 3040 11580 3045 11610
rect 3005 11570 3045 11580
rect 3205 11580 3210 11610
rect 3240 11580 3245 11610
rect 3205 11570 3245 11580
rect 3405 11580 3410 11610
rect 3440 11580 3445 11610
rect 3405 11570 3445 11580
rect 3605 11580 3610 11610
rect 3640 11580 3645 11610
rect 3605 11570 3645 11580
rect 3805 11580 3810 11610
rect 3840 11580 3845 11610
rect 3805 11570 3845 11580
rect 4005 11580 4010 11610
rect 4040 11580 4045 11610
rect 4005 11570 4045 11580
rect 4205 11580 4210 11610
rect 4240 11580 4245 11610
rect 4205 11570 4245 11580
rect 4405 11580 4410 11610
rect 4440 11580 4445 11610
rect 4405 11570 4445 11580
rect 4605 11580 4610 11610
rect 4640 11580 4645 11610
rect 4605 11570 4645 11580
rect 4805 11580 4810 11610
rect 4840 11580 4845 11610
rect 4805 11570 4845 11580
rect 5005 11580 5010 11610
rect 5040 11580 5045 11610
rect 5005 11570 5045 11580
rect 5205 11580 5210 11610
rect 5240 11580 5245 11610
rect 5205 11570 5245 11580
rect 5405 11580 5410 11610
rect 5440 11580 5445 11610
rect 5405 11570 5445 11580
rect 5605 11580 5610 11610
rect 5640 11580 5645 11610
rect 5605 11570 5645 11580
rect 5805 11580 5810 11610
rect 5840 11580 5845 11610
rect 5805 11570 5845 11580
rect 6005 11580 6010 11610
rect 6040 11580 6045 11610
rect 6005 11570 6045 11580
rect 6205 11580 6210 11610
rect 6240 11580 6245 11610
rect 6205 11570 6245 11580
rect 6405 11580 6410 11610
rect 6440 11580 6445 11610
rect 6405 11570 6445 11580
rect -165 11550 -30 11570
rect 5 11550 6570 11570
rect -165 11540 -155 11550
rect -195 11510 -190 11540
rect -160 11510 -155 11540
rect 5 11540 45 11550
rect 5 11510 10 11540
rect 40 11510 45 11540
rect 205 11540 245 11550
rect 205 11510 210 11540
rect 240 11510 245 11540
rect 405 11540 445 11550
rect 405 11510 410 11540
rect 440 11510 445 11540
rect 605 11540 645 11550
rect 605 11510 610 11540
rect 640 11510 645 11540
rect 805 11540 845 11550
rect 805 11510 810 11540
rect 840 11510 845 11540
rect 1005 11540 1045 11550
rect 1005 11510 1010 11540
rect 1040 11510 1045 11540
rect 1205 11540 1245 11550
rect 1205 11510 1210 11540
rect 1240 11510 1245 11540
rect 1405 11540 1445 11550
rect 1405 11510 1410 11540
rect 1440 11510 1445 11540
rect 1605 11540 1645 11550
rect 1605 11510 1610 11540
rect 1640 11510 1645 11540
rect 1805 11540 1845 11550
rect 1805 11510 1810 11540
rect 1840 11510 1845 11540
rect 2005 11540 2045 11550
rect 2005 11510 2010 11540
rect 2040 11510 2045 11540
rect 2205 11540 2245 11550
rect 2205 11510 2210 11540
rect 2240 11510 2245 11540
rect 2405 11540 2445 11550
rect 2405 11510 2410 11540
rect 2440 11510 2445 11540
rect 2605 11540 2645 11550
rect 2605 11510 2610 11540
rect 2640 11510 2645 11540
rect 2805 11540 2845 11550
rect 2805 11510 2810 11540
rect 2840 11510 2845 11540
rect 3005 11540 3045 11550
rect 3005 11510 3010 11540
rect 3040 11510 3045 11540
rect 3205 11540 3245 11550
rect 3205 11510 3210 11540
rect 3240 11510 3245 11540
rect 3405 11540 3445 11550
rect 3405 11510 3410 11540
rect 3440 11510 3445 11540
rect 3605 11540 3645 11550
rect 3605 11510 3610 11540
rect 3640 11510 3645 11540
rect 3805 11540 3845 11550
rect 3805 11510 3810 11540
rect 3840 11510 3845 11540
rect 4005 11540 4045 11550
rect 4005 11510 4010 11540
rect 4040 11510 4045 11540
rect 4205 11540 4245 11550
rect 4205 11510 4210 11540
rect 4240 11510 4245 11540
rect 4405 11540 4445 11550
rect 4405 11510 4410 11540
rect 4440 11510 4445 11540
rect 4605 11540 4645 11550
rect 4605 11510 4610 11540
rect 4640 11510 4645 11540
rect 4805 11540 4845 11550
rect 4805 11510 4810 11540
rect 4840 11510 4845 11540
rect 5005 11540 5045 11550
rect 5005 11510 5010 11540
rect 5040 11510 5045 11540
rect 5205 11540 5245 11550
rect 5205 11510 5210 11540
rect 5240 11510 5245 11540
rect 5405 11540 5445 11550
rect 5405 11510 5410 11540
rect 5440 11510 5445 11540
rect 5605 11540 5645 11550
rect 5605 11510 5610 11540
rect 5640 11510 5645 11540
rect 5805 11540 5845 11550
rect 5805 11510 5810 11540
rect 5840 11510 5845 11540
rect 6005 11540 6045 11550
rect 6005 11510 6010 11540
rect 6040 11510 6045 11540
rect 6205 11540 6245 11550
rect 6205 11510 6210 11540
rect 6240 11510 6245 11540
rect 6405 11540 6445 11550
rect 6405 11510 6410 11540
rect 6440 11510 6445 11540
rect -188 11425 -185 11510
rect -165 11425 -162 11510
rect 15 11425 35 11510
rect 215 11425 235 11510
rect 415 11425 435 11510
rect 615 11425 635 11510
rect 815 11425 835 11510
rect 1015 11425 1035 11510
rect 1215 11425 1235 11510
rect 1415 11425 1435 11510
rect 1615 11425 1635 11510
rect 1815 11425 1835 11510
rect 2015 11425 2035 11510
rect 2215 11425 2235 11510
rect 2415 11425 2435 11510
rect 2615 11425 2635 11510
rect 2815 11425 2835 11510
rect 3015 11425 3035 11510
rect 3215 11425 3235 11510
rect 3415 11425 3435 11510
rect 3615 11425 3635 11510
rect 3815 11425 3835 11510
rect 4015 11425 4035 11510
rect 4215 11425 4235 11510
rect 4415 11425 4435 11510
rect 4615 11425 4635 11510
rect 4815 11425 4835 11510
rect 5015 11425 5035 11510
rect 5215 11425 5235 11510
rect 5415 11425 5435 11510
rect 5615 11425 5635 11510
rect 5815 11425 5835 11510
rect 6015 11425 6035 11510
rect 6215 11425 6235 11510
rect -195 11395 -190 11425
rect -160 11395 -155 11425
rect -195 11355 -185 11395
rect -165 11385 -155 11395
rect 5 11395 10 11425
rect 40 11395 45 11425
rect 5 11385 45 11395
rect 205 11395 210 11425
rect 240 11395 245 11425
rect 205 11385 245 11395
rect 405 11395 410 11425
rect 440 11395 445 11425
rect 405 11385 445 11395
rect 605 11395 610 11425
rect 640 11395 645 11425
rect 605 11385 645 11395
rect 805 11395 810 11425
rect 840 11395 845 11425
rect 805 11385 845 11395
rect 1005 11395 1010 11425
rect 1040 11395 1045 11425
rect 1005 11385 1045 11395
rect 1205 11395 1210 11425
rect 1240 11395 1245 11425
rect 1205 11385 1245 11395
rect 1405 11395 1410 11425
rect 1440 11395 1445 11425
rect 1405 11385 1445 11395
rect 1605 11395 1610 11425
rect 1640 11395 1645 11425
rect 1605 11385 1645 11395
rect 1805 11395 1810 11425
rect 1840 11395 1845 11425
rect 1805 11385 1845 11395
rect 2005 11395 2010 11425
rect 2040 11395 2045 11425
rect 2005 11385 2045 11395
rect 2205 11395 2210 11425
rect 2240 11395 2245 11425
rect 2205 11385 2245 11395
rect 2405 11395 2410 11425
rect 2440 11395 2445 11425
rect 2405 11385 2445 11395
rect 2605 11395 2610 11425
rect 2640 11395 2645 11425
rect 2605 11385 2645 11395
rect 2805 11395 2810 11425
rect 2840 11395 2845 11425
rect 2805 11385 2845 11395
rect 3005 11395 3010 11425
rect 3040 11395 3045 11425
rect 3005 11385 3045 11395
rect 3205 11395 3210 11425
rect 3240 11395 3245 11425
rect 3205 11385 3245 11395
rect 3405 11395 3410 11425
rect 3440 11395 3445 11425
rect 3405 11385 3445 11395
rect 3605 11395 3610 11425
rect 3640 11395 3645 11425
rect 3605 11385 3645 11395
rect 3805 11395 3810 11425
rect 3840 11395 3845 11425
rect 3805 11385 3845 11395
rect 4005 11395 4010 11425
rect 4040 11395 4045 11425
rect 4005 11385 4045 11395
rect 4205 11395 4210 11425
rect 4240 11395 4245 11425
rect 4205 11385 4245 11395
rect 4405 11395 4410 11425
rect 4440 11395 4445 11425
rect 4405 11385 4445 11395
rect 4605 11395 4610 11425
rect 4640 11395 4645 11425
rect 4605 11385 4645 11395
rect 4805 11395 4810 11425
rect 4840 11395 4845 11425
rect 4805 11385 4845 11395
rect 5005 11395 5010 11425
rect 5040 11395 5045 11425
rect 5005 11385 5045 11395
rect 5205 11395 5210 11425
rect 5240 11395 5245 11425
rect 5205 11385 5245 11395
rect 5405 11395 5410 11425
rect 5440 11395 5445 11425
rect 5405 11385 5445 11395
rect 5605 11395 5610 11425
rect 5640 11395 5645 11425
rect 5605 11385 5645 11395
rect 5805 11395 5810 11425
rect 5840 11395 5845 11425
rect 5805 11385 5845 11395
rect 6005 11395 6010 11425
rect 6040 11395 6045 11425
rect 6005 11385 6045 11395
rect 6205 11395 6210 11425
rect 6240 11395 6245 11425
rect 6205 11385 6245 11395
rect 6405 11395 6410 11425
rect 6440 11395 6445 11425
rect 6405 11385 6445 11395
rect -165 11365 -30 11385
rect 5 11365 6570 11385
rect -165 11355 -155 11365
rect -195 11325 -190 11355
rect -160 11325 -155 11355
rect 5 11355 45 11365
rect 5 11325 10 11355
rect 40 11325 45 11355
rect 205 11355 245 11365
rect 205 11325 210 11355
rect 240 11325 245 11355
rect 405 11355 445 11365
rect 405 11325 410 11355
rect 440 11325 445 11355
rect 605 11355 645 11365
rect 605 11325 610 11355
rect 640 11325 645 11355
rect 805 11355 845 11365
rect 805 11325 810 11355
rect 840 11325 845 11355
rect 1005 11355 1045 11365
rect 1005 11325 1010 11355
rect 1040 11325 1045 11355
rect 1205 11355 1245 11365
rect 1205 11325 1210 11355
rect 1240 11325 1245 11355
rect 1405 11355 1445 11365
rect 1405 11325 1410 11355
rect 1440 11325 1445 11355
rect 1605 11355 1645 11365
rect 1605 11325 1610 11355
rect 1640 11325 1645 11355
rect 1805 11355 1845 11365
rect 1805 11325 1810 11355
rect 1840 11325 1845 11355
rect 2005 11355 2045 11365
rect 2005 11325 2010 11355
rect 2040 11325 2045 11355
rect 2205 11355 2245 11365
rect 2205 11325 2210 11355
rect 2240 11325 2245 11355
rect 2405 11355 2445 11365
rect 2405 11325 2410 11355
rect 2440 11325 2445 11355
rect 2605 11355 2645 11365
rect 2605 11325 2610 11355
rect 2640 11325 2645 11355
rect 2805 11355 2845 11365
rect 2805 11325 2810 11355
rect 2840 11325 2845 11355
rect 3005 11355 3045 11365
rect 3005 11325 3010 11355
rect 3040 11325 3045 11355
rect 3205 11355 3245 11365
rect 3205 11325 3210 11355
rect 3240 11325 3245 11355
rect 3405 11355 3445 11365
rect 3405 11325 3410 11355
rect 3440 11325 3445 11355
rect 3605 11355 3645 11365
rect 3605 11325 3610 11355
rect 3640 11325 3645 11355
rect 3805 11355 3845 11365
rect 3805 11325 3810 11355
rect 3840 11325 3845 11355
rect 4005 11355 4045 11365
rect 4005 11325 4010 11355
rect 4040 11325 4045 11355
rect 4205 11355 4245 11365
rect 4205 11325 4210 11355
rect 4240 11325 4245 11355
rect 4405 11355 4445 11365
rect 4405 11325 4410 11355
rect 4440 11325 4445 11355
rect 4605 11355 4645 11365
rect 4605 11325 4610 11355
rect 4640 11325 4645 11355
rect 4805 11355 4845 11365
rect 4805 11325 4810 11355
rect 4840 11325 4845 11355
rect 5005 11355 5045 11365
rect 5005 11325 5010 11355
rect 5040 11325 5045 11355
rect 5205 11355 5245 11365
rect 5205 11325 5210 11355
rect 5240 11325 5245 11355
rect 5405 11355 5445 11365
rect 5405 11325 5410 11355
rect 5440 11325 5445 11355
rect 5605 11355 5645 11365
rect 5605 11325 5610 11355
rect 5640 11325 5645 11355
rect 5805 11355 5845 11365
rect 5805 11325 5810 11355
rect 5840 11325 5845 11355
rect 6005 11355 6045 11365
rect 6005 11325 6010 11355
rect 6040 11325 6045 11355
rect 6205 11355 6245 11365
rect 6205 11325 6210 11355
rect 6240 11325 6245 11355
rect 6405 11355 6445 11365
rect 6405 11325 6410 11355
rect 6440 11325 6445 11355
rect -188 11240 -185 11325
rect -165 11240 -162 11325
rect 15 11240 35 11325
rect 215 11240 235 11325
rect 415 11240 435 11325
rect 615 11240 635 11325
rect 815 11240 835 11325
rect 1015 11240 1035 11325
rect 1215 11240 1235 11325
rect 1415 11240 1435 11325
rect 1615 11240 1635 11325
rect 1815 11240 1835 11325
rect 2015 11240 2035 11325
rect 2215 11240 2235 11325
rect 2415 11240 2435 11325
rect 2615 11240 2635 11325
rect 2815 11240 2835 11325
rect 3015 11240 3035 11325
rect 3215 11240 3235 11325
rect 3415 11240 3435 11325
rect 3615 11240 3635 11325
rect 3815 11240 3835 11325
rect 4015 11240 4035 11325
rect 4215 11240 4235 11325
rect 4415 11240 4435 11325
rect 4615 11240 4635 11325
rect 4815 11240 4835 11325
rect 5015 11240 5035 11325
rect 5215 11240 5235 11325
rect 5415 11240 5435 11325
rect 5615 11240 5635 11325
rect 5815 11240 5835 11325
rect 6015 11240 6035 11325
rect 6215 11240 6235 11325
rect -195 11210 -190 11240
rect -160 11210 -155 11240
rect -195 11170 -185 11210
rect -165 11200 -155 11210
rect 5 11210 10 11240
rect 40 11210 45 11240
rect 5 11200 45 11210
rect 205 11210 210 11240
rect 240 11210 245 11240
rect 205 11200 245 11210
rect 405 11210 410 11240
rect 440 11210 445 11240
rect 405 11200 445 11210
rect 605 11210 610 11240
rect 640 11210 645 11240
rect 605 11200 645 11210
rect 805 11210 810 11240
rect 840 11210 845 11240
rect 805 11200 845 11210
rect 1005 11210 1010 11240
rect 1040 11210 1045 11240
rect 1005 11200 1045 11210
rect 1205 11210 1210 11240
rect 1240 11210 1245 11240
rect 1205 11200 1245 11210
rect 1405 11210 1410 11240
rect 1440 11210 1445 11240
rect 1405 11200 1445 11210
rect 1605 11210 1610 11240
rect 1640 11210 1645 11240
rect 1605 11200 1645 11210
rect 1805 11210 1810 11240
rect 1840 11210 1845 11240
rect 1805 11200 1845 11210
rect 2005 11210 2010 11240
rect 2040 11210 2045 11240
rect 2005 11200 2045 11210
rect 2205 11210 2210 11240
rect 2240 11210 2245 11240
rect 2205 11200 2245 11210
rect 2405 11210 2410 11240
rect 2440 11210 2445 11240
rect 2405 11200 2445 11210
rect 2605 11210 2610 11240
rect 2640 11210 2645 11240
rect 2605 11200 2645 11210
rect 2805 11210 2810 11240
rect 2840 11210 2845 11240
rect 2805 11200 2845 11210
rect 3005 11210 3010 11240
rect 3040 11210 3045 11240
rect 3005 11200 3045 11210
rect 3205 11210 3210 11240
rect 3240 11210 3245 11240
rect 3205 11200 3245 11210
rect 3405 11210 3410 11240
rect 3440 11210 3445 11240
rect 3405 11200 3445 11210
rect 3605 11210 3610 11240
rect 3640 11210 3645 11240
rect 3605 11200 3645 11210
rect 3805 11210 3810 11240
rect 3840 11210 3845 11240
rect 3805 11200 3845 11210
rect 4005 11210 4010 11240
rect 4040 11210 4045 11240
rect 4005 11200 4045 11210
rect 4205 11210 4210 11240
rect 4240 11210 4245 11240
rect 4205 11200 4245 11210
rect 4405 11210 4410 11240
rect 4440 11210 4445 11240
rect 4405 11200 4445 11210
rect 4605 11210 4610 11240
rect 4640 11210 4645 11240
rect 4605 11200 4645 11210
rect 4805 11210 4810 11240
rect 4840 11210 4845 11240
rect 4805 11200 4845 11210
rect 5005 11210 5010 11240
rect 5040 11210 5045 11240
rect 5005 11200 5045 11210
rect 5205 11210 5210 11240
rect 5240 11210 5245 11240
rect 5205 11200 5245 11210
rect 5405 11210 5410 11240
rect 5440 11210 5445 11240
rect 5405 11200 5445 11210
rect 5605 11210 5610 11240
rect 5640 11210 5645 11240
rect 5605 11200 5645 11210
rect 5805 11210 5810 11240
rect 5840 11210 5845 11240
rect 5805 11200 5845 11210
rect 6005 11210 6010 11240
rect 6040 11210 6045 11240
rect 6005 11200 6045 11210
rect 6205 11210 6210 11240
rect 6240 11210 6245 11240
rect 6205 11200 6245 11210
rect 6405 11210 6410 11240
rect 6440 11210 6445 11240
rect 6405 11200 6445 11210
rect -165 11180 -30 11200
rect 5 11180 6570 11200
rect -165 11170 -155 11180
rect -195 11140 -190 11170
rect -160 11140 -155 11170
rect 5 11170 45 11180
rect 5 11140 10 11170
rect 40 11140 45 11170
rect 205 11170 245 11180
rect 205 11140 210 11170
rect 240 11140 245 11170
rect 405 11170 445 11180
rect 405 11140 410 11170
rect 440 11140 445 11170
rect 605 11170 645 11180
rect 605 11140 610 11170
rect 640 11140 645 11170
rect 805 11170 845 11180
rect 805 11140 810 11170
rect 840 11140 845 11170
rect 1005 11170 1045 11180
rect 1005 11140 1010 11170
rect 1040 11140 1045 11170
rect 1205 11170 1245 11180
rect 1205 11140 1210 11170
rect 1240 11140 1245 11170
rect 1405 11170 1445 11180
rect 1405 11140 1410 11170
rect 1440 11140 1445 11170
rect 1605 11170 1645 11180
rect 1605 11140 1610 11170
rect 1640 11140 1645 11170
rect 1805 11170 1845 11180
rect 1805 11140 1810 11170
rect 1840 11140 1845 11170
rect 2005 11170 2045 11180
rect 2005 11140 2010 11170
rect 2040 11140 2045 11170
rect 2205 11170 2245 11180
rect 2205 11140 2210 11170
rect 2240 11140 2245 11170
rect 2405 11170 2445 11180
rect 2405 11140 2410 11170
rect 2440 11140 2445 11170
rect 2605 11170 2645 11180
rect 2605 11140 2610 11170
rect 2640 11140 2645 11170
rect 2805 11170 2845 11180
rect 2805 11140 2810 11170
rect 2840 11140 2845 11170
rect 3005 11170 3045 11180
rect 3005 11140 3010 11170
rect 3040 11140 3045 11170
rect 3205 11170 3245 11180
rect 3205 11140 3210 11170
rect 3240 11140 3245 11170
rect 3405 11170 3445 11180
rect 3405 11140 3410 11170
rect 3440 11140 3445 11170
rect 3605 11170 3645 11180
rect 3605 11140 3610 11170
rect 3640 11140 3645 11170
rect 3805 11170 3845 11180
rect 3805 11140 3810 11170
rect 3840 11140 3845 11170
rect 4005 11170 4045 11180
rect 4005 11140 4010 11170
rect 4040 11140 4045 11170
rect 4205 11170 4245 11180
rect 4205 11140 4210 11170
rect 4240 11140 4245 11170
rect 4405 11170 4445 11180
rect 4405 11140 4410 11170
rect 4440 11140 4445 11170
rect 4605 11170 4645 11180
rect 4605 11140 4610 11170
rect 4640 11140 4645 11170
rect 4805 11170 4845 11180
rect 4805 11140 4810 11170
rect 4840 11140 4845 11170
rect 5005 11170 5045 11180
rect 5005 11140 5010 11170
rect 5040 11140 5045 11170
rect 5205 11170 5245 11180
rect 5205 11140 5210 11170
rect 5240 11140 5245 11170
rect 5405 11170 5445 11180
rect 5405 11140 5410 11170
rect 5440 11140 5445 11170
rect 5605 11170 5645 11180
rect 5605 11140 5610 11170
rect 5640 11140 5645 11170
rect 5805 11170 5845 11180
rect 5805 11140 5810 11170
rect 5840 11140 5845 11170
rect 6005 11170 6045 11180
rect 6005 11140 6010 11170
rect 6040 11140 6045 11170
rect 6205 11170 6245 11180
rect 6205 11140 6210 11170
rect 6240 11140 6245 11170
rect 6405 11170 6445 11180
rect 6405 11140 6410 11170
rect 6440 11140 6445 11170
rect -188 11055 -185 11140
rect -165 11055 -162 11140
rect 15 11055 35 11140
rect 215 11055 235 11140
rect 415 11055 435 11140
rect 615 11055 635 11140
rect 815 11055 835 11140
rect 1015 11055 1035 11140
rect 1215 11055 1235 11140
rect 1415 11055 1435 11140
rect 1615 11055 1635 11140
rect 1815 11055 1835 11140
rect 2015 11055 2035 11140
rect 2215 11055 2235 11140
rect 2415 11055 2435 11140
rect 2615 11055 2635 11140
rect 2815 11055 2835 11140
rect 3015 11055 3035 11140
rect 3215 11055 3235 11140
rect 3415 11055 3435 11140
rect 3615 11055 3635 11140
rect 3815 11055 3835 11140
rect 4015 11055 4035 11140
rect 4215 11055 4235 11140
rect 4415 11055 4435 11140
rect 4615 11055 4635 11140
rect 4815 11055 4835 11140
rect 5015 11055 5035 11140
rect 5215 11055 5235 11140
rect 5415 11055 5435 11140
rect 5615 11055 5635 11140
rect 5815 11055 5835 11140
rect 6015 11055 6035 11140
rect 6215 11055 6235 11140
rect -195 11025 -190 11055
rect -160 11025 -155 11055
rect -195 10985 -185 11025
rect -165 11015 -155 11025
rect 5 11025 10 11055
rect 40 11025 45 11055
rect 5 11015 45 11025
rect 205 11025 210 11055
rect 240 11025 245 11055
rect 205 11015 245 11025
rect 405 11025 410 11055
rect 440 11025 445 11055
rect 405 11015 445 11025
rect 605 11025 610 11055
rect 640 11025 645 11055
rect 605 11015 645 11025
rect 805 11025 810 11055
rect 840 11025 845 11055
rect 805 11015 845 11025
rect 1005 11025 1010 11055
rect 1040 11025 1045 11055
rect 1005 11015 1045 11025
rect 1205 11025 1210 11055
rect 1240 11025 1245 11055
rect 1205 11015 1245 11025
rect 1405 11025 1410 11055
rect 1440 11025 1445 11055
rect 1405 11015 1445 11025
rect 1605 11025 1610 11055
rect 1640 11025 1645 11055
rect 1605 11015 1645 11025
rect 1805 11025 1810 11055
rect 1840 11025 1845 11055
rect 1805 11015 1845 11025
rect 2005 11025 2010 11055
rect 2040 11025 2045 11055
rect 2005 11015 2045 11025
rect 2205 11025 2210 11055
rect 2240 11025 2245 11055
rect 2205 11015 2245 11025
rect 2405 11025 2410 11055
rect 2440 11025 2445 11055
rect 2405 11015 2445 11025
rect 2605 11025 2610 11055
rect 2640 11025 2645 11055
rect 2605 11015 2645 11025
rect 2805 11025 2810 11055
rect 2840 11025 2845 11055
rect 2805 11015 2845 11025
rect 3005 11025 3010 11055
rect 3040 11025 3045 11055
rect 3005 11015 3045 11025
rect 3205 11025 3210 11055
rect 3240 11025 3245 11055
rect 3205 11015 3245 11025
rect 3405 11025 3410 11055
rect 3440 11025 3445 11055
rect 3405 11015 3445 11025
rect 3605 11025 3610 11055
rect 3640 11025 3645 11055
rect 3605 11015 3645 11025
rect 3805 11025 3810 11055
rect 3840 11025 3845 11055
rect 3805 11015 3845 11025
rect 4005 11025 4010 11055
rect 4040 11025 4045 11055
rect 4005 11015 4045 11025
rect 4205 11025 4210 11055
rect 4240 11025 4245 11055
rect 4205 11015 4245 11025
rect 4405 11025 4410 11055
rect 4440 11025 4445 11055
rect 4405 11015 4445 11025
rect 4605 11025 4610 11055
rect 4640 11025 4645 11055
rect 4605 11015 4645 11025
rect 4805 11025 4810 11055
rect 4840 11025 4845 11055
rect 4805 11015 4845 11025
rect 5005 11025 5010 11055
rect 5040 11025 5045 11055
rect 5005 11015 5045 11025
rect 5205 11025 5210 11055
rect 5240 11025 5245 11055
rect 5205 11015 5245 11025
rect 5405 11025 5410 11055
rect 5440 11025 5445 11055
rect 5405 11015 5445 11025
rect 5605 11025 5610 11055
rect 5640 11025 5645 11055
rect 5605 11015 5645 11025
rect 5805 11025 5810 11055
rect 5840 11025 5845 11055
rect 5805 11015 5845 11025
rect 6005 11025 6010 11055
rect 6040 11025 6045 11055
rect 6005 11015 6045 11025
rect 6205 11025 6210 11055
rect 6240 11025 6245 11055
rect 6205 11015 6245 11025
rect 6405 11025 6410 11055
rect 6440 11025 6445 11055
rect 6405 11015 6445 11025
rect -165 10995 -30 11015
rect 5 10995 6570 11015
rect -165 10985 -155 10995
rect -195 10955 -190 10985
rect -160 10955 -155 10985
rect 5 10985 45 10995
rect 5 10955 10 10985
rect 40 10955 45 10985
rect 205 10985 245 10995
rect 205 10955 210 10985
rect 240 10955 245 10985
rect 405 10985 445 10995
rect 405 10955 410 10985
rect 440 10955 445 10985
rect 605 10985 645 10995
rect 605 10955 610 10985
rect 640 10955 645 10985
rect 805 10985 845 10995
rect 805 10955 810 10985
rect 840 10955 845 10985
rect 1005 10985 1045 10995
rect 1005 10955 1010 10985
rect 1040 10955 1045 10985
rect 1205 10985 1245 10995
rect 1205 10955 1210 10985
rect 1240 10955 1245 10985
rect 1405 10985 1445 10995
rect 1405 10955 1410 10985
rect 1440 10955 1445 10985
rect 1605 10985 1645 10995
rect 1605 10955 1610 10985
rect 1640 10955 1645 10985
rect 1805 10985 1845 10995
rect 1805 10955 1810 10985
rect 1840 10955 1845 10985
rect 2005 10985 2045 10995
rect 2005 10955 2010 10985
rect 2040 10955 2045 10985
rect 2205 10985 2245 10995
rect 2205 10955 2210 10985
rect 2240 10955 2245 10985
rect 2405 10985 2445 10995
rect 2405 10955 2410 10985
rect 2440 10955 2445 10985
rect 2605 10985 2645 10995
rect 2605 10955 2610 10985
rect 2640 10955 2645 10985
rect 2805 10985 2845 10995
rect 2805 10955 2810 10985
rect 2840 10955 2845 10985
rect 3005 10985 3045 10995
rect 3005 10955 3010 10985
rect 3040 10955 3045 10985
rect 3205 10985 3245 10995
rect 3205 10955 3210 10985
rect 3240 10955 3245 10985
rect 3405 10985 3445 10995
rect 3405 10955 3410 10985
rect 3440 10955 3445 10985
rect 3605 10985 3645 10995
rect 3605 10955 3610 10985
rect 3640 10955 3645 10985
rect 3805 10985 3845 10995
rect 3805 10955 3810 10985
rect 3840 10955 3845 10985
rect 4005 10985 4045 10995
rect 4005 10955 4010 10985
rect 4040 10955 4045 10985
rect 4205 10985 4245 10995
rect 4205 10955 4210 10985
rect 4240 10955 4245 10985
rect 4405 10985 4445 10995
rect 4405 10955 4410 10985
rect 4440 10955 4445 10985
rect 4605 10985 4645 10995
rect 4605 10955 4610 10985
rect 4640 10955 4645 10985
rect 4805 10985 4845 10995
rect 4805 10955 4810 10985
rect 4840 10955 4845 10985
rect 5005 10985 5045 10995
rect 5005 10955 5010 10985
rect 5040 10955 5045 10985
rect 5205 10985 5245 10995
rect 5205 10955 5210 10985
rect 5240 10955 5245 10985
rect 5405 10985 5445 10995
rect 5405 10955 5410 10985
rect 5440 10955 5445 10985
rect 5605 10985 5645 10995
rect 5605 10955 5610 10985
rect 5640 10955 5645 10985
rect 5805 10985 5845 10995
rect 5805 10955 5810 10985
rect 5840 10955 5845 10985
rect 6005 10985 6045 10995
rect 6005 10955 6010 10985
rect 6040 10955 6045 10985
rect 6205 10985 6245 10995
rect 6205 10955 6210 10985
rect 6240 10955 6245 10985
rect 6405 10985 6445 10995
rect 6405 10955 6410 10985
rect 6440 10955 6445 10985
rect -188 10870 -185 10955
rect -165 10870 -162 10955
rect 15 10870 35 10955
rect 215 10870 235 10955
rect 415 10870 435 10955
rect 615 10870 635 10955
rect 815 10870 835 10955
rect 1015 10870 1035 10955
rect 1215 10870 1235 10955
rect 1415 10870 1435 10955
rect 1615 10870 1635 10955
rect 1815 10870 1835 10955
rect 2015 10870 2035 10955
rect 2215 10870 2235 10955
rect 2415 10870 2435 10955
rect 2615 10870 2635 10955
rect 2815 10870 2835 10955
rect 3015 10870 3035 10955
rect 3215 10870 3235 10955
rect 3415 10870 3435 10955
rect 3615 10870 3635 10955
rect 3815 10870 3835 10955
rect 4015 10870 4035 10955
rect 4215 10870 4235 10955
rect 4415 10870 4435 10955
rect 4615 10870 4635 10955
rect 4815 10870 4835 10955
rect 5015 10870 5035 10955
rect 5215 10870 5235 10955
rect 5415 10870 5435 10955
rect 5615 10870 5635 10955
rect 5815 10870 5835 10955
rect 6015 10870 6035 10955
rect 6215 10870 6235 10955
rect -195 10840 -190 10870
rect -160 10840 -155 10870
rect -195 10800 -185 10840
rect -165 10830 -155 10840
rect 5 10840 10 10870
rect 40 10840 45 10870
rect 5 10830 45 10840
rect 205 10840 210 10870
rect 240 10840 245 10870
rect 205 10830 245 10840
rect 405 10840 410 10870
rect 440 10840 445 10870
rect 405 10830 445 10840
rect 605 10840 610 10870
rect 640 10840 645 10870
rect 605 10830 645 10840
rect 805 10840 810 10870
rect 840 10840 845 10870
rect 805 10830 845 10840
rect 1005 10840 1010 10870
rect 1040 10840 1045 10870
rect 1005 10830 1045 10840
rect 1205 10840 1210 10870
rect 1240 10840 1245 10870
rect 1205 10830 1245 10840
rect 1405 10840 1410 10870
rect 1440 10840 1445 10870
rect 1405 10830 1445 10840
rect 1605 10840 1610 10870
rect 1640 10840 1645 10870
rect 1605 10830 1645 10840
rect 1805 10840 1810 10870
rect 1840 10840 1845 10870
rect 1805 10830 1845 10840
rect 2005 10840 2010 10870
rect 2040 10840 2045 10870
rect 2005 10830 2045 10840
rect 2205 10840 2210 10870
rect 2240 10840 2245 10870
rect 2205 10830 2245 10840
rect 2405 10840 2410 10870
rect 2440 10840 2445 10870
rect 2405 10830 2445 10840
rect 2605 10840 2610 10870
rect 2640 10840 2645 10870
rect 2605 10830 2645 10840
rect 2805 10840 2810 10870
rect 2840 10840 2845 10870
rect 2805 10830 2845 10840
rect 3005 10840 3010 10870
rect 3040 10840 3045 10870
rect 3005 10830 3045 10840
rect 3205 10840 3210 10870
rect 3240 10840 3245 10870
rect 3205 10830 3245 10840
rect 3405 10840 3410 10870
rect 3440 10840 3445 10870
rect 3405 10830 3445 10840
rect 3605 10840 3610 10870
rect 3640 10840 3645 10870
rect 3605 10830 3645 10840
rect 3805 10840 3810 10870
rect 3840 10840 3845 10870
rect 3805 10830 3845 10840
rect 4005 10840 4010 10870
rect 4040 10840 4045 10870
rect 4005 10830 4045 10840
rect 4205 10840 4210 10870
rect 4240 10840 4245 10870
rect 4205 10830 4245 10840
rect 4405 10840 4410 10870
rect 4440 10840 4445 10870
rect 4405 10830 4445 10840
rect 4605 10840 4610 10870
rect 4640 10840 4645 10870
rect 4605 10830 4645 10840
rect 4805 10840 4810 10870
rect 4840 10840 4845 10870
rect 4805 10830 4845 10840
rect 5005 10840 5010 10870
rect 5040 10840 5045 10870
rect 5005 10830 5045 10840
rect 5205 10840 5210 10870
rect 5240 10840 5245 10870
rect 5205 10830 5245 10840
rect 5405 10840 5410 10870
rect 5440 10840 5445 10870
rect 5405 10830 5445 10840
rect 5605 10840 5610 10870
rect 5640 10840 5645 10870
rect 5605 10830 5645 10840
rect 5805 10840 5810 10870
rect 5840 10840 5845 10870
rect 5805 10830 5845 10840
rect 6005 10840 6010 10870
rect 6040 10840 6045 10870
rect 6005 10830 6045 10840
rect 6205 10840 6210 10870
rect 6240 10840 6245 10870
rect 6205 10830 6245 10840
rect 6405 10840 6410 10870
rect 6440 10840 6445 10870
rect 6405 10830 6445 10840
rect -165 10810 -30 10830
rect 5 10810 6570 10830
rect -165 10800 -155 10810
rect -195 10770 -190 10800
rect -160 10770 -155 10800
rect 5 10800 45 10810
rect 5 10770 10 10800
rect 40 10770 45 10800
rect 205 10800 245 10810
rect 205 10770 210 10800
rect 240 10770 245 10800
rect 405 10800 445 10810
rect 405 10770 410 10800
rect 440 10770 445 10800
rect 605 10800 645 10810
rect 605 10770 610 10800
rect 640 10770 645 10800
rect 805 10800 845 10810
rect 805 10770 810 10800
rect 840 10770 845 10800
rect 1005 10800 1045 10810
rect 1005 10770 1010 10800
rect 1040 10770 1045 10800
rect 1205 10800 1245 10810
rect 1205 10770 1210 10800
rect 1240 10770 1245 10800
rect 1405 10800 1445 10810
rect 1405 10770 1410 10800
rect 1440 10770 1445 10800
rect 1605 10800 1645 10810
rect 1605 10770 1610 10800
rect 1640 10770 1645 10800
rect 1805 10800 1845 10810
rect 1805 10770 1810 10800
rect 1840 10770 1845 10800
rect 2005 10800 2045 10810
rect 2005 10770 2010 10800
rect 2040 10770 2045 10800
rect 2205 10800 2245 10810
rect 2205 10770 2210 10800
rect 2240 10770 2245 10800
rect 2405 10800 2445 10810
rect 2405 10770 2410 10800
rect 2440 10770 2445 10800
rect 2605 10800 2645 10810
rect 2605 10770 2610 10800
rect 2640 10770 2645 10800
rect 2805 10800 2845 10810
rect 2805 10770 2810 10800
rect 2840 10770 2845 10800
rect 3005 10800 3045 10810
rect 3005 10770 3010 10800
rect 3040 10770 3045 10800
rect 3205 10800 3245 10810
rect 3205 10770 3210 10800
rect 3240 10770 3245 10800
rect 3405 10800 3445 10810
rect 3405 10770 3410 10800
rect 3440 10770 3445 10800
rect 3605 10800 3645 10810
rect 3605 10770 3610 10800
rect 3640 10770 3645 10800
rect 3805 10800 3845 10810
rect 3805 10770 3810 10800
rect 3840 10770 3845 10800
rect 4005 10800 4045 10810
rect 4005 10770 4010 10800
rect 4040 10770 4045 10800
rect 4205 10800 4245 10810
rect 4205 10770 4210 10800
rect 4240 10770 4245 10800
rect 4405 10800 4445 10810
rect 4405 10770 4410 10800
rect 4440 10770 4445 10800
rect 4605 10800 4645 10810
rect 4605 10770 4610 10800
rect 4640 10770 4645 10800
rect 4805 10800 4845 10810
rect 4805 10770 4810 10800
rect 4840 10770 4845 10800
rect 5005 10800 5045 10810
rect 5005 10770 5010 10800
rect 5040 10770 5045 10800
rect 5205 10800 5245 10810
rect 5205 10770 5210 10800
rect 5240 10770 5245 10800
rect 5405 10800 5445 10810
rect 5405 10770 5410 10800
rect 5440 10770 5445 10800
rect 5605 10800 5645 10810
rect 5605 10770 5610 10800
rect 5640 10770 5645 10800
rect 5805 10800 5845 10810
rect 5805 10770 5810 10800
rect 5840 10770 5845 10800
rect 6005 10800 6045 10810
rect 6005 10770 6010 10800
rect 6040 10770 6045 10800
rect 6205 10800 6245 10810
rect 6205 10770 6210 10800
rect 6240 10770 6245 10800
rect 6405 10800 6445 10810
rect 6405 10770 6410 10800
rect 6440 10770 6445 10800
rect -188 10685 -185 10770
rect -165 10685 -162 10770
rect 15 10685 35 10770
rect 215 10685 235 10770
rect 415 10685 435 10770
rect 615 10685 635 10770
rect 815 10685 835 10770
rect 1015 10685 1035 10770
rect 1215 10685 1235 10770
rect 1415 10685 1435 10770
rect 1615 10685 1635 10770
rect 1815 10685 1835 10770
rect 2015 10685 2035 10770
rect 2215 10685 2235 10770
rect 2415 10685 2435 10770
rect 2615 10685 2635 10770
rect 2815 10685 2835 10770
rect 3015 10685 3035 10770
rect 3215 10685 3235 10770
rect 3415 10685 3435 10770
rect 3615 10685 3635 10770
rect 3815 10685 3835 10770
rect 4015 10685 4035 10770
rect 4215 10685 4235 10770
rect 4415 10685 4435 10770
rect 4615 10685 4635 10770
rect 4815 10685 4835 10770
rect 5015 10685 5035 10770
rect 5215 10685 5235 10770
rect 5415 10685 5435 10770
rect 5615 10685 5635 10770
rect 5815 10685 5835 10770
rect 6015 10685 6035 10770
rect 6215 10685 6235 10770
rect -195 10655 -190 10685
rect -160 10655 -155 10685
rect -195 10615 -185 10655
rect -165 10645 -155 10655
rect 5 10655 10 10685
rect 40 10655 45 10685
rect 5 10645 45 10655
rect 205 10655 210 10685
rect 240 10655 245 10685
rect 205 10645 245 10655
rect 405 10655 410 10685
rect 440 10655 445 10685
rect 405 10645 445 10655
rect 605 10655 610 10685
rect 640 10655 645 10685
rect 605 10645 645 10655
rect 805 10655 810 10685
rect 840 10655 845 10685
rect 805 10645 845 10655
rect 1005 10655 1010 10685
rect 1040 10655 1045 10685
rect 1005 10645 1045 10655
rect 1205 10655 1210 10685
rect 1240 10655 1245 10685
rect 1205 10645 1245 10655
rect 1405 10655 1410 10685
rect 1440 10655 1445 10685
rect 1405 10645 1445 10655
rect 1605 10655 1610 10685
rect 1640 10655 1645 10685
rect 1605 10645 1645 10655
rect 1805 10655 1810 10685
rect 1840 10655 1845 10685
rect 1805 10645 1845 10655
rect 2005 10655 2010 10685
rect 2040 10655 2045 10685
rect 2005 10645 2045 10655
rect 2205 10655 2210 10685
rect 2240 10655 2245 10685
rect 2205 10645 2245 10655
rect 2405 10655 2410 10685
rect 2440 10655 2445 10685
rect 2405 10645 2445 10655
rect 2605 10655 2610 10685
rect 2640 10655 2645 10685
rect 2605 10645 2645 10655
rect 2805 10655 2810 10685
rect 2840 10655 2845 10685
rect 2805 10645 2845 10655
rect 3005 10655 3010 10685
rect 3040 10655 3045 10685
rect 3005 10645 3045 10655
rect 3205 10655 3210 10685
rect 3240 10655 3245 10685
rect 3205 10645 3245 10655
rect 3405 10655 3410 10685
rect 3440 10655 3445 10685
rect 3405 10645 3445 10655
rect 3605 10655 3610 10685
rect 3640 10655 3645 10685
rect 3605 10645 3645 10655
rect 3805 10655 3810 10685
rect 3840 10655 3845 10685
rect 3805 10645 3845 10655
rect 4005 10655 4010 10685
rect 4040 10655 4045 10685
rect 4005 10645 4045 10655
rect 4205 10655 4210 10685
rect 4240 10655 4245 10685
rect 4205 10645 4245 10655
rect 4405 10655 4410 10685
rect 4440 10655 4445 10685
rect 4405 10645 4445 10655
rect 4605 10655 4610 10685
rect 4640 10655 4645 10685
rect 4605 10645 4645 10655
rect 4805 10655 4810 10685
rect 4840 10655 4845 10685
rect 4805 10645 4845 10655
rect 5005 10655 5010 10685
rect 5040 10655 5045 10685
rect 5005 10645 5045 10655
rect 5205 10655 5210 10685
rect 5240 10655 5245 10685
rect 5205 10645 5245 10655
rect 5405 10655 5410 10685
rect 5440 10655 5445 10685
rect 5405 10645 5445 10655
rect 5605 10655 5610 10685
rect 5640 10655 5645 10685
rect 5605 10645 5645 10655
rect 5805 10655 5810 10685
rect 5840 10655 5845 10685
rect 5805 10645 5845 10655
rect 6005 10655 6010 10685
rect 6040 10655 6045 10685
rect 6005 10645 6045 10655
rect 6205 10655 6210 10685
rect 6240 10655 6245 10685
rect 6205 10645 6245 10655
rect 6405 10655 6410 10685
rect 6440 10655 6445 10685
rect 6405 10645 6445 10655
rect -165 10625 -30 10645
rect 5 10625 6570 10645
rect -165 10615 -155 10625
rect -195 10585 -190 10615
rect -160 10585 -155 10615
rect 5 10615 45 10625
rect 5 10585 10 10615
rect 40 10585 45 10615
rect 205 10615 245 10625
rect 205 10585 210 10615
rect 240 10585 245 10615
rect 405 10615 445 10625
rect 405 10585 410 10615
rect 440 10585 445 10615
rect 605 10615 645 10625
rect 605 10585 610 10615
rect 640 10585 645 10615
rect 805 10615 845 10625
rect 805 10585 810 10615
rect 840 10585 845 10615
rect 1005 10615 1045 10625
rect 1005 10585 1010 10615
rect 1040 10585 1045 10615
rect 1205 10615 1245 10625
rect 1205 10585 1210 10615
rect 1240 10585 1245 10615
rect 1405 10615 1445 10625
rect 1405 10585 1410 10615
rect 1440 10585 1445 10615
rect 1605 10615 1645 10625
rect 1605 10585 1610 10615
rect 1640 10585 1645 10615
rect 1805 10615 1845 10625
rect 1805 10585 1810 10615
rect 1840 10585 1845 10615
rect 2005 10615 2045 10625
rect 2005 10585 2010 10615
rect 2040 10585 2045 10615
rect 2205 10615 2245 10625
rect 2205 10585 2210 10615
rect 2240 10585 2245 10615
rect 2405 10615 2445 10625
rect 2405 10585 2410 10615
rect 2440 10585 2445 10615
rect 2605 10615 2645 10625
rect 2605 10585 2610 10615
rect 2640 10585 2645 10615
rect 2805 10615 2845 10625
rect 2805 10585 2810 10615
rect 2840 10585 2845 10615
rect 3005 10615 3045 10625
rect 3005 10585 3010 10615
rect 3040 10585 3045 10615
rect 3205 10615 3245 10625
rect 3205 10585 3210 10615
rect 3240 10585 3245 10615
rect 3405 10615 3445 10625
rect 3405 10585 3410 10615
rect 3440 10585 3445 10615
rect 3605 10615 3645 10625
rect 3605 10585 3610 10615
rect 3640 10585 3645 10615
rect 3805 10615 3845 10625
rect 3805 10585 3810 10615
rect 3840 10585 3845 10615
rect 4005 10615 4045 10625
rect 4005 10585 4010 10615
rect 4040 10585 4045 10615
rect 4205 10615 4245 10625
rect 4205 10585 4210 10615
rect 4240 10585 4245 10615
rect 4405 10615 4445 10625
rect 4405 10585 4410 10615
rect 4440 10585 4445 10615
rect 4605 10615 4645 10625
rect 4605 10585 4610 10615
rect 4640 10585 4645 10615
rect 4805 10615 4845 10625
rect 4805 10585 4810 10615
rect 4840 10585 4845 10615
rect 5005 10615 5045 10625
rect 5005 10585 5010 10615
rect 5040 10585 5045 10615
rect 5205 10615 5245 10625
rect 5205 10585 5210 10615
rect 5240 10585 5245 10615
rect 5405 10615 5445 10625
rect 5405 10585 5410 10615
rect 5440 10585 5445 10615
rect 5605 10615 5645 10625
rect 5605 10585 5610 10615
rect 5640 10585 5645 10615
rect 5805 10615 5845 10625
rect 5805 10585 5810 10615
rect 5840 10585 5845 10615
rect 6005 10615 6045 10625
rect 6005 10585 6010 10615
rect 6040 10585 6045 10615
rect 6205 10615 6245 10625
rect 6205 10585 6210 10615
rect 6240 10585 6245 10615
rect 6405 10615 6445 10625
rect 6405 10585 6410 10615
rect 6440 10585 6445 10615
rect -188 10500 -185 10585
rect -165 10500 -162 10585
rect 15 10500 35 10585
rect 215 10500 235 10585
rect 415 10500 435 10585
rect 615 10500 635 10585
rect 815 10500 835 10585
rect 1015 10500 1035 10585
rect 1215 10500 1235 10585
rect 1415 10500 1435 10585
rect 1615 10500 1635 10585
rect 1815 10500 1835 10585
rect 2015 10500 2035 10585
rect 2215 10500 2235 10585
rect 2415 10500 2435 10585
rect 2615 10500 2635 10585
rect 2815 10500 2835 10585
rect 3015 10500 3035 10585
rect 3215 10500 3235 10585
rect 3415 10500 3435 10585
rect 3615 10500 3635 10585
rect 3815 10500 3835 10585
rect 4015 10500 4035 10585
rect 4215 10500 4235 10585
rect 4415 10500 4435 10585
rect 4615 10500 4635 10585
rect 4815 10500 4835 10585
rect 5015 10500 5035 10585
rect 5215 10500 5235 10585
rect 5415 10500 5435 10585
rect 5615 10500 5635 10585
rect 5815 10500 5835 10585
rect 6015 10500 6035 10585
rect 6215 10500 6235 10585
rect -195 10470 -190 10500
rect -160 10470 -155 10500
rect -195 10430 -185 10470
rect -165 10460 -155 10470
rect 5 10470 10 10500
rect 40 10470 45 10500
rect 5 10460 45 10470
rect 205 10470 210 10500
rect 240 10470 245 10500
rect 205 10460 245 10470
rect 405 10470 410 10500
rect 440 10470 445 10500
rect 405 10460 445 10470
rect 605 10470 610 10500
rect 640 10470 645 10500
rect 605 10460 645 10470
rect 805 10470 810 10500
rect 840 10470 845 10500
rect 805 10460 845 10470
rect 1005 10470 1010 10500
rect 1040 10470 1045 10500
rect 1005 10460 1045 10470
rect 1205 10470 1210 10500
rect 1240 10470 1245 10500
rect 1205 10460 1245 10470
rect 1405 10470 1410 10500
rect 1440 10470 1445 10500
rect 1405 10460 1445 10470
rect 1605 10470 1610 10500
rect 1640 10470 1645 10500
rect 1605 10460 1645 10470
rect 1805 10470 1810 10500
rect 1840 10470 1845 10500
rect 1805 10460 1845 10470
rect 2005 10470 2010 10500
rect 2040 10470 2045 10500
rect 2005 10460 2045 10470
rect 2205 10470 2210 10500
rect 2240 10470 2245 10500
rect 2205 10460 2245 10470
rect 2405 10470 2410 10500
rect 2440 10470 2445 10500
rect 2405 10460 2445 10470
rect 2605 10470 2610 10500
rect 2640 10470 2645 10500
rect 2605 10460 2645 10470
rect 2805 10470 2810 10500
rect 2840 10470 2845 10500
rect 2805 10460 2845 10470
rect 3005 10470 3010 10500
rect 3040 10470 3045 10500
rect 3005 10460 3045 10470
rect 3205 10470 3210 10500
rect 3240 10470 3245 10500
rect 3205 10460 3245 10470
rect 3405 10470 3410 10500
rect 3440 10470 3445 10500
rect 3405 10460 3445 10470
rect 3605 10470 3610 10500
rect 3640 10470 3645 10500
rect 3605 10460 3645 10470
rect 3805 10470 3810 10500
rect 3840 10470 3845 10500
rect 3805 10460 3845 10470
rect 4005 10470 4010 10500
rect 4040 10470 4045 10500
rect 4005 10460 4045 10470
rect 4205 10470 4210 10500
rect 4240 10470 4245 10500
rect 4205 10460 4245 10470
rect 4405 10470 4410 10500
rect 4440 10470 4445 10500
rect 4405 10460 4445 10470
rect 4605 10470 4610 10500
rect 4640 10470 4645 10500
rect 4605 10460 4645 10470
rect 4805 10470 4810 10500
rect 4840 10470 4845 10500
rect 4805 10460 4845 10470
rect 5005 10470 5010 10500
rect 5040 10470 5045 10500
rect 5005 10460 5045 10470
rect 5205 10470 5210 10500
rect 5240 10470 5245 10500
rect 5205 10460 5245 10470
rect 5405 10470 5410 10500
rect 5440 10470 5445 10500
rect 5405 10460 5445 10470
rect 5605 10470 5610 10500
rect 5640 10470 5645 10500
rect 5605 10460 5645 10470
rect 5805 10470 5810 10500
rect 5840 10470 5845 10500
rect 5805 10460 5845 10470
rect 6005 10470 6010 10500
rect 6040 10470 6045 10500
rect 6005 10460 6045 10470
rect 6205 10470 6210 10500
rect 6240 10470 6245 10500
rect 6205 10460 6245 10470
rect 6405 10470 6410 10500
rect 6440 10470 6445 10500
rect 6405 10460 6445 10470
rect -165 10440 -30 10460
rect 5 10440 6570 10460
rect -165 10430 -155 10440
rect -195 10400 -190 10430
rect -160 10400 -155 10430
rect 5 10430 45 10440
rect 5 10400 10 10430
rect 40 10400 45 10430
rect 205 10430 245 10440
rect 205 10400 210 10430
rect 240 10400 245 10430
rect 405 10430 445 10440
rect 405 10400 410 10430
rect 440 10400 445 10430
rect 605 10430 645 10440
rect 605 10400 610 10430
rect 640 10400 645 10430
rect 805 10430 845 10440
rect 805 10400 810 10430
rect 840 10400 845 10430
rect 1005 10430 1045 10440
rect 1005 10400 1010 10430
rect 1040 10400 1045 10430
rect 1205 10430 1245 10440
rect 1205 10400 1210 10430
rect 1240 10400 1245 10430
rect 1405 10430 1445 10440
rect 1405 10400 1410 10430
rect 1440 10400 1445 10430
rect 1605 10430 1645 10440
rect 1605 10400 1610 10430
rect 1640 10400 1645 10430
rect 1805 10430 1845 10440
rect 1805 10400 1810 10430
rect 1840 10400 1845 10430
rect 2005 10430 2045 10440
rect 2005 10400 2010 10430
rect 2040 10400 2045 10430
rect 2205 10430 2245 10440
rect 2205 10400 2210 10430
rect 2240 10400 2245 10430
rect 2405 10430 2445 10440
rect 2405 10400 2410 10430
rect 2440 10400 2445 10430
rect 2605 10430 2645 10440
rect 2605 10400 2610 10430
rect 2640 10400 2645 10430
rect 2805 10430 2845 10440
rect 2805 10400 2810 10430
rect 2840 10400 2845 10430
rect 3005 10430 3045 10440
rect 3005 10400 3010 10430
rect 3040 10400 3045 10430
rect 3205 10430 3245 10440
rect 3205 10400 3210 10430
rect 3240 10400 3245 10430
rect 3405 10430 3445 10440
rect 3405 10400 3410 10430
rect 3440 10400 3445 10430
rect 3605 10430 3645 10440
rect 3605 10400 3610 10430
rect 3640 10400 3645 10430
rect 3805 10430 3845 10440
rect 3805 10400 3810 10430
rect 3840 10400 3845 10430
rect 4005 10430 4045 10440
rect 4005 10400 4010 10430
rect 4040 10400 4045 10430
rect 4205 10430 4245 10440
rect 4205 10400 4210 10430
rect 4240 10400 4245 10430
rect 4405 10430 4445 10440
rect 4405 10400 4410 10430
rect 4440 10400 4445 10430
rect 4605 10430 4645 10440
rect 4605 10400 4610 10430
rect 4640 10400 4645 10430
rect 4805 10430 4845 10440
rect 4805 10400 4810 10430
rect 4840 10400 4845 10430
rect 5005 10430 5045 10440
rect 5005 10400 5010 10430
rect 5040 10400 5045 10430
rect 5205 10430 5245 10440
rect 5205 10400 5210 10430
rect 5240 10400 5245 10430
rect 5405 10430 5445 10440
rect 5405 10400 5410 10430
rect 5440 10400 5445 10430
rect 5605 10430 5645 10440
rect 5605 10400 5610 10430
rect 5640 10400 5645 10430
rect 5805 10430 5845 10440
rect 5805 10400 5810 10430
rect 5840 10400 5845 10430
rect 6005 10430 6045 10440
rect 6005 10400 6010 10430
rect 6040 10400 6045 10430
rect 6205 10430 6245 10440
rect 6205 10400 6210 10430
rect 6240 10400 6245 10430
rect 6405 10430 6445 10440
rect 6405 10400 6410 10430
rect 6440 10400 6445 10430
rect -188 10315 -185 10400
rect -165 10315 -162 10400
rect 15 10315 35 10400
rect 215 10315 235 10400
rect 415 10315 435 10400
rect 615 10315 635 10400
rect 815 10315 835 10400
rect 1015 10315 1035 10400
rect 1215 10315 1235 10400
rect 1415 10315 1435 10400
rect 1615 10315 1635 10400
rect 1815 10315 1835 10400
rect 2015 10315 2035 10400
rect 2215 10315 2235 10400
rect 2415 10315 2435 10400
rect 2615 10315 2635 10400
rect 2815 10315 2835 10400
rect 3015 10315 3035 10400
rect 3215 10315 3235 10400
rect 3415 10315 3435 10400
rect 3615 10315 3635 10400
rect 3815 10315 3835 10400
rect 4015 10315 4035 10400
rect 4215 10315 4235 10400
rect 4415 10315 4435 10400
rect 4615 10315 4635 10400
rect 4815 10315 4835 10400
rect 5015 10315 5035 10400
rect 5215 10315 5235 10400
rect 5415 10315 5435 10400
rect 5615 10315 5635 10400
rect 5815 10315 5835 10400
rect 6015 10315 6035 10400
rect 6215 10315 6235 10400
rect -195 10285 -190 10315
rect -160 10285 -155 10315
rect -195 10245 -185 10285
rect -165 10275 -155 10285
rect 5 10285 10 10315
rect 40 10285 45 10315
rect 5 10275 45 10285
rect 205 10285 210 10315
rect 240 10285 245 10315
rect 205 10275 245 10285
rect 405 10285 410 10315
rect 440 10285 445 10315
rect 405 10275 445 10285
rect 605 10285 610 10315
rect 640 10285 645 10315
rect 605 10275 645 10285
rect 805 10285 810 10315
rect 840 10285 845 10315
rect 805 10275 845 10285
rect 1005 10285 1010 10315
rect 1040 10285 1045 10315
rect 1005 10275 1045 10285
rect 1205 10285 1210 10315
rect 1240 10285 1245 10315
rect 1205 10275 1245 10285
rect 1405 10285 1410 10315
rect 1440 10285 1445 10315
rect 1405 10275 1445 10285
rect 1605 10285 1610 10315
rect 1640 10285 1645 10315
rect 1605 10275 1645 10285
rect 1805 10285 1810 10315
rect 1840 10285 1845 10315
rect 1805 10275 1845 10285
rect 2005 10285 2010 10315
rect 2040 10285 2045 10315
rect 2005 10275 2045 10285
rect 2205 10285 2210 10315
rect 2240 10285 2245 10315
rect 2205 10275 2245 10285
rect 2405 10285 2410 10315
rect 2440 10285 2445 10315
rect 2405 10275 2445 10285
rect 2605 10285 2610 10315
rect 2640 10285 2645 10315
rect 2605 10275 2645 10285
rect 2805 10285 2810 10315
rect 2840 10285 2845 10315
rect 2805 10275 2845 10285
rect 3005 10285 3010 10315
rect 3040 10285 3045 10315
rect 3005 10275 3045 10285
rect 3205 10285 3210 10315
rect 3240 10285 3245 10315
rect 3205 10275 3245 10285
rect 3405 10285 3410 10315
rect 3440 10285 3445 10315
rect 3405 10275 3445 10285
rect 3605 10285 3610 10315
rect 3640 10285 3645 10315
rect 3605 10275 3645 10285
rect 3805 10285 3810 10315
rect 3840 10285 3845 10315
rect 3805 10275 3845 10285
rect 4005 10285 4010 10315
rect 4040 10285 4045 10315
rect 4005 10275 4045 10285
rect 4205 10285 4210 10315
rect 4240 10285 4245 10315
rect 4205 10275 4245 10285
rect 4405 10285 4410 10315
rect 4440 10285 4445 10315
rect 4405 10275 4445 10285
rect 4605 10285 4610 10315
rect 4640 10285 4645 10315
rect 4605 10275 4645 10285
rect 4805 10285 4810 10315
rect 4840 10285 4845 10315
rect 4805 10275 4845 10285
rect 5005 10285 5010 10315
rect 5040 10285 5045 10315
rect 5005 10275 5045 10285
rect 5205 10285 5210 10315
rect 5240 10285 5245 10315
rect 5205 10275 5245 10285
rect 5405 10285 5410 10315
rect 5440 10285 5445 10315
rect 5405 10275 5445 10285
rect 5605 10285 5610 10315
rect 5640 10285 5645 10315
rect 5605 10275 5645 10285
rect 5805 10285 5810 10315
rect 5840 10285 5845 10315
rect 5805 10275 5845 10285
rect 6005 10285 6010 10315
rect 6040 10285 6045 10315
rect 6005 10275 6045 10285
rect 6205 10285 6210 10315
rect 6240 10285 6245 10315
rect 6205 10275 6245 10285
rect 6405 10285 6410 10315
rect 6440 10285 6445 10315
rect 6405 10275 6445 10285
rect -165 10255 -30 10275
rect 5 10255 6570 10275
rect -165 10245 -155 10255
rect -195 10215 -190 10245
rect -160 10215 -155 10245
rect 5 10245 45 10255
rect 5 10215 10 10245
rect 40 10215 45 10245
rect 205 10245 245 10255
rect 205 10215 210 10245
rect 240 10215 245 10245
rect 405 10245 445 10255
rect 405 10215 410 10245
rect 440 10215 445 10245
rect 605 10245 645 10255
rect 605 10215 610 10245
rect 640 10215 645 10245
rect 805 10245 845 10255
rect 805 10215 810 10245
rect 840 10215 845 10245
rect 1005 10245 1045 10255
rect 1005 10215 1010 10245
rect 1040 10215 1045 10245
rect 1205 10245 1245 10255
rect 1205 10215 1210 10245
rect 1240 10215 1245 10245
rect 1405 10245 1445 10255
rect 1405 10215 1410 10245
rect 1440 10215 1445 10245
rect 1605 10245 1645 10255
rect 1605 10215 1610 10245
rect 1640 10215 1645 10245
rect 1805 10245 1845 10255
rect 1805 10215 1810 10245
rect 1840 10215 1845 10245
rect 2005 10245 2045 10255
rect 2005 10215 2010 10245
rect 2040 10215 2045 10245
rect 2205 10245 2245 10255
rect 2205 10215 2210 10245
rect 2240 10215 2245 10245
rect 2405 10245 2445 10255
rect 2405 10215 2410 10245
rect 2440 10215 2445 10245
rect 2605 10245 2645 10255
rect 2605 10215 2610 10245
rect 2640 10215 2645 10245
rect 2805 10245 2845 10255
rect 2805 10215 2810 10245
rect 2840 10215 2845 10245
rect 3005 10245 3045 10255
rect 3005 10215 3010 10245
rect 3040 10215 3045 10245
rect 3205 10245 3245 10255
rect 3205 10215 3210 10245
rect 3240 10215 3245 10245
rect 3405 10245 3445 10255
rect 3405 10215 3410 10245
rect 3440 10215 3445 10245
rect 3605 10245 3645 10255
rect 3605 10215 3610 10245
rect 3640 10215 3645 10245
rect 3805 10245 3845 10255
rect 3805 10215 3810 10245
rect 3840 10215 3845 10245
rect 4005 10245 4045 10255
rect 4005 10215 4010 10245
rect 4040 10215 4045 10245
rect 4205 10245 4245 10255
rect 4205 10215 4210 10245
rect 4240 10215 4245 10245
rect 4405 10245 4445 10255
rect 4405 10215 4410 10245
rect 4440 10215 4445 10245
rect 4605 10245 4645 10255
rect 4605 10215 4610 10245
rect 4640 10215 4645 10245
rect 4805 10245 4845 10255
rect 4805 10215 4810 10245
rect 4840 10215 4845 10245
rect 5005 10245 5045 10255
rect 5005 10215 5010 10245
rect 5040 10215 5045 10245
rect 5205 10245 5245 10255
rect 5205 10215 5210 10245
rect 5240 10215 5245 10245
rect 5405 10245 5445 10255
rect 5405 10215 5410 10245
rect 5440 10215 5445 10245
rect 5605 10245 5645 10255
rect 5605 10215 5610 10245
rect 5640 10215 5645 10245
rect 5805 10245 5845 10255
rect 5805 10215 5810 10245
rect 5840 10215 5845 10245
rect 6005 10245 6045 10255
rect 6005 10215 6010 10245
rect 6040 10215 6045 10245
rect 6205 10245 6245 10255
rect 6205 10215 6210 10245
rect 6240 10215 6245 10245
rect 6405 10245 6445 10255
rect 6405 10215 6410 10245
rect 6440 10215 6445 10245
rect -188 10130 -185 10215
rect -165 10130 -162 10215
rect 15 10130 35 10215
rect 215 10130 235 10215
rect 415 10130 435 10215
rect 615 10130 635 10215
rect 815 10130 835 10215
rect 1015 10130 1035 10215
rect 1215 10130 1235 10215
rect 1415 10130 1435 10215
rect 1615 10130 1635 10215
rect 1815 10130 1835 10215
rect 2015 10130 2035 10215
rect 2215 10130 2235 10215
rect 2415 10130 2435 10215
rect 2615 10130 2635 10215
rect 2815 10130 2835 10215
rect 3015 10130 3035 10215
rect 3215 10130 3235 10215
rect 3415 10130 3435 10215
rect 3615 10130 3635 10215
rect 3815 10130 3835 10215
rect 4015 10130 4035 10215
rect 4215 10130 4235 10215
rect 4415 10130 4435 10215
rect 4615 10130 4635 10215
rect 4815 10130 4835 10215
rect 5015 10130 5035 10215
rect 5215 10130 5235 10215
rect 5415 10130 5435 10215
rect 5615 10130 5635 10215
rect 5815 10130 5835 10215
rect 6015 10130 6035 10215
rect 6215 10130 6235 10215
rect -195 10100 -190 10130
rect -160 10100 -155 10130
rect -195 10060 -185 10100
rect -165 10090 -155 10100
rect 5 10100 10 10130
rect 40 10100 45 10130
rect 5 10090 45 10100
rect 205 10100 210 10130
rect 240 10100 245 10130
rect 205 10090 245 10100
rect 405 10100 410 10130
rect 440 10100 445 10130
rect 405 10090 445 10100
rect 605 10100 610 10130
rect 640 10100 645 10130
rect 605 10090 645 10100
rect 805 10100 810 10130
rect 840 10100 845 10130
rect 805 10090 845 10100
rect 1005 10100 1010 10130
rect 1040 10100 1045 10130
rect 1005 10090 1045 10100
rect 1205 10100 1210 10130
rect 1240 10100 1245 10130
rect 1205 10090 1245 10100
rect 1405 10100 1410 10130
rect 1440 10100 1445 10130
rect 1405 10090 1445 10100
rect 1605 10100 1610 10130
rect 1640 10100 1645 10130
rect 1605 10090 1645 10100
rect 1805 10100 1810 10130
rect 1840 10100 1845 10130
rect 1805 10090 1845 10100
rect 2005 10100 2010 10130
rect 2040 10100 2045 10130
rect 2005 10090 2045 10100
rect 2205 10100 2210 10130
rect 2240 10100 2245 10130
rect 2205 10090 2245 10100
rect 2405 10100 2410 10130
rect 2440 10100 2445 10130
rect 2405 10090 2445 10100
rect 2605 10100 2610 10130
rect 2640 10100 2645 10130
rect 2605 10090 2645 10100
rect 2805 10100 2810 10130
rect 2840 10100 2845 10130
rect 2805 10090 2845 10100
rect 3005 10100 3010 10130
rect 3040 10100 3045 10130
rect 3005 10090 3045 10100
rect 3205 10100 3210 10130
rect 3240 10100 3245 10130
rect 3205 10090 3245 10100
rect 3405 10100 3410 10130
rect 3440 10100 3445 10130
rect 3405 10090 3445 10100
rect 3605 10100 3610 10130
rect 3640 10100 3645 10130
rect 3605 10090 3645 10100
rect 3805 10100 3810 10130
rect 3840 10100 3845 10130
rect 3805 10090 3845 10100
rect 4005 10100 4010 10130
rect 4040 10100 4045 10130
rect 4005 10090 4045 10100
rect 4205 10100 4210 10130
rect 4240 10100 4245 10130
rect 4205 10090 4245 10100
rect 4405 10100 4410 10130
rect 4440 10100 4445 10130
rect 4405 10090 4445 10100
rect 4605 10100 4610 10130
rect 4640 10100 4645 10130
rect 4605 10090 4645 10100
rect 4805 10100 4810 10130
rect 4840 10100 4845 10130
rect 4805 10090 4845 10100
rect 5005 10100 5010 10130
rect 5040 10100 5045 10130
rect 5005 10090 5045 10100
rect 5205 10100 5210 10130
rect 5240 10100 5245 10130
rect 5205 10090 5245 10100
rect 5405 10100 5410 10130
rect 5440 10100 5445 10130
rect 5405 10090 5445 10100
rect 5605 10100 5610 10130
rect 5640 10100 5645 10130
rect 5605 10090 5645 10100
rect 5805 10100 5810 10130
rect 5840 10100 5845 10130
rect 5805 10090 5845 10100
rect 6005 10100 6010 10130
rect 6040 10100 6045 10130
rect 6005 10090 6045 10100
rect 6205 10100 6210 10130
rect 6240 10100 6245 10130
rect 6205 10090 6245 10100
rect 6405 10100 6410 10130
rect 6440 10100 6445 10130
rect 6405 10090 6445 10100
rect -165 10070 -30 10090
rect 5 10070 6570 10090
rect -165 10060 -155 10070
rect -195 10030 -190 10060
rect -160 10030 -155 10060
rect 5 10060 45 10070
rect 5 10030 10 10060
rect 40 10030 45 10060
rect 205 10060 245 10070
rect 205 10030 210 10060
rect 240 10030 245 10060
rect 405 10060 445 10070
rect 405 10030 410 10060
rect 440 10030 445 10060
rect 605 10060 645 10070
rect 605 10030 610 10060
rect 640 10030 645 10060
rect 805 10060 845 10070
rect 805 10030 810 10060
rect 840 10030 845 10060
rect 1005 10060 1045 10070
rect 1005 10030 1010 10060
rect 1040 10030 1045 10060
rect 1205 10060 1245 10070
rect 1205 10030 1210 10060
rect 1240 10030 1245 10060
rect 1405 10060 1445 10070
rect 1405 10030 1410 10060
rect 1440 10030 1445 10060
rect 1605 10060 1645 10070
rect 1605 10030 1610 10060
rect 1640 10030 1645 10060
rect 1805 10060 1845 10070
rect 1805 10030 1810 10060
rect 1840 10030 1845 10060
rect 2005 10060 2045 10070
rect 2005 10030 2010 10060
rect 2040 10030 2045 10060
rect 2205 10060 2245 10070
rect 2205 10030 2210 10060
rect 2240 10030 2245 10060
rect 2405 10060 2445 10070
rect 2405 10030 2410 10060
rect 2440 10030 2445 10060
rect 2605 10060 2645 10070
rect 2605 10030 2610 10060
rect 2640 10030 2645 10060
rect 2805 10060 2845 10070
rect 2805 10030 2810 10060
rect 2840 10030 2845 10060
rect 3005 10060 3045 10070
rect 3005 10030 3010 10060
rect 3040 10030 3045 10060
rect 3205 10060 3245 10070
rect 3205 10030 3210 10060
rect 3240 10030 3245 10060
rect 3405 10060 3445 10070
rect 3405 10030 3410 10060
rect 3440 10030 3445 10060
rect 3605 10060 3645 10070
rect 3605 10030 3610 10060
rect 3640 10030 3645 10060
rect 3805 10060 3845 10070
rect 3805 10030 3810 10060
rect 3840 10030 3845 10060
rect 4005 10060 4045 10070
rect 4005 10030 4010 10060
rect 4040 10030 4045 10060
rect 4205 10060 4245 10070
rect 4205 10030 4210 10060
rect 4240 10030 4245 10060
rect 4405 10060 4445 10070
rect 4405 10030 4410 10060
rect 4440 10030 4445 10060
rect 4605 10060 4645 10070
rect 4605 10030 4610 10060
rect 4640 10030 4645 10060
rect 4805 10060 4845 10070
rect 4805 10030 4810 10060
rect 4840 10030 4845 10060
rect 5005 10060 5045 10070
rect 5005 10030 5010 10060
rect 5040 10030 5045 10060
rect 5205 10060 5245 10070
rect 5205 10030 5210 10060
rect 5240 10030 5245 10060
rect 5405 10060 5445 10070
rect 5405 10030 5410 10060
rect 5440 10030 5445 10060
rect 5605 10060 5645 10070
rect 5605 10030 5610 10060
rect 5640 10030 5645 10060
rect 5805 10060 5845 10070
rect 5805 10030 5810 10060
rect 5840 10030 5845 10060
rect 6005 10060 6045 10070
rect 6005 10030 6010 10060
rect 6040 10030 6045 10060
rect 6205 10060 6245 10070
rect 6205 10030 6210 10060
rect 6240 10030 6245 10060
rect 6405 10060 6445 10070
rect 6405 10030 6410 10060
rect 6440 10030 6445 10060
rect -188 9945 -185 10030
rect -165 9945 -162 10030
rect 15 9945 35 10030
rect 215 9945 235 10030
rect 415 9945 435 10030
rect 615 9945 635 10030
rect 815 9945 835 10030
rect 1015 9945 1035 10030
rect 1215 9945 1235 10030
rect 1415 9945 1435 10030
rect 1615 9945 1635 10030
rect 1815 9945 1835 10030
rect 2015 9945 2035 10030
rect 2215 9945 2235 10030
rect 2415 9945 2435 10030
rect 2615 9945 2635 10030
rect 2815 9945 2835 10030
rect 3015 9945 3035 10030
rect 3215 9945 3235 10030
rect 3415 9945 3435 10030
rect 3615 9945 3635 10030
rect 3815 9945 3835 10030
rect 4015 9945 4035 10030
rect 4215 9945 4235 10030
rect 4415 9945 4435 10030
rect 4615 9945 4635 10030
rect 4815 9945 4835 10030
rect 5015 9945 5035 10030
rect 5215 9945 5235 10030
rect 5415 9945 5435 10030
rect 5615 9945 5635 10030
rect 5815 9945 5835 10030
rect 6015 9945 6035 10030
rect 6215 9945 6235 10030
rect -195 9915 -190 9945
rect -160 9915 -155 9945
rect -195 9875 -185 9915
rect -165 9905 -155 9915
rect 5 9915 10 9945
rect 40 9915 45 9945
rect 5 9905 45 9915
rect 205 9915 210 9945
rect 240 9915 245 9945
rect 205 9905 245 9915
rect 405 9915 410 9945
rect 440 9915 445 9945
rect 405 9905 445 9915
rect 605 9915 610 9945
rect 640 9915 645 9945
rect 605 9905 645 9915
rect 805 9915 810 9945
rect 840 9915 845 9945
rect 805 9905 845 9915
rect 1005 9915 1010 9945
rect 1040 9915 1045 9945
rect 1005 9905 1045 9915
rect 1205 9915 1210 9945
rect 1240 9915 1245 9945
rect 1205 9905 1245 9915
rect 1405 9915 1410 9945
rect 1440 9915 1445 9945
rect 1405 9905 1445 9915
rect 1605 9915 1610 9945
rect 1640 9915 1645 9945
rect 1605 9905 1645 9915
rect 1805 9915 1810 9945
rect 1840 9915 1845 9945
rect 1805 9905 1845 9915
rect 2005 9915 2010 9945
rect 2040 9915 2045 9945
rect 2005 9905 2045 9915
rect 2205 9915 2210 9945
rect 2240 9915 2245 9945
rect 2205 9905 2245 9915
rect 2405 9915 2410 9945
rect 2440 9915 2445 9945
rect 2405 9905 2445 9915
rect 2605 9915 2610 9945
rect 2640 9915 2645 9945
rect 2605 9905 2645 9915
rect 2805 9915 2810 9945
rect 2840 9915 2845 9945
rect 2805 9905 2845 9915
rect 3005 9915 3010 9945
rect 3040 9915 3045 9945
rect 3005 9905 3045 9915
rect 3205 9915 3210 9945
rect 3240 9915 3245 9945
rect 3205 9905 3245 9915
rect 3405 9915 3410 9945
rect 3440 9915 3445 9945
rect 3405 9905 3445 9915
rect 3605 9915 3610 9945
rect 3640 9915 3645 9945
rect 3605 9905 3645 9915
rect 3805 9915 3810 9945
rect 3840 9915 3845 9945
rect 3805 9905 3845 9915
rect 4005 9915 4010 9945
rect 4040 9915 4045 9945
rect 4005 9905 4045 9915
rect 4205 9915 4210 9945
rect 4240 9915 4245 9945
rect 4205 9905 4245 9915
rect 4405 9915 4410 9945
rect 4440 9915 4445 9945
rect 4405 9905 4445 9915
rect 4605 9915 4610 9945
rect 4640 9915 4645 9945
rect 4605 9905 4645 9915
rect 4805 9915 4810 9945
rect 4840 9915 4845 9945
rect 4805 9905 4845 9915
rect 5005 9915 5010 9945
rect 5040 9915 5045 9945
rect 5005 9905 5045 9915
rect 5205 9915 5210 9945
rect 5240 9915 5245 9945
rect 5205 9905 5245 9915
rect 5405 9915 5410 9945
rect 5440 9915 5445 9945
rect 5405 9905 5445 9915
rect 5605 9915 5610 9945
rect 5640 9915 5645 9945
rect 5605 9905 5645 9915
rect 5805 9915 5810 9945
rect 5840 9915 5845 9945
rect 5805 9905 5845 9915
rect 6005 9915 6010 9945
rect 6040 9915 6045 9945
rect 6005 9905 6045 9915
rect 6205 9915 6210 9945
rect 6240 9915 6245 9945
rect 6205 9905 6245 9915
rect 6405 9915 6410 9945
rect 6440 9915 6445 9945
rect 6405 9905 6445 9915
rect -165 9885 -30 9905
rect 5 9885 6570 9905
rect -165 9875 -155 9885
rect -195 9845 -190 9875
rect -160 9845 -155 9875
rect 5 9875 45 9885
rect 5 9845 10 9875
rect 40 9845 45 9875
rect 205 9875 245 9885
rect 205 9845 210 9875
rect 240 9845 245 9875
rect 405 9875 445 9885
rect 405 9845 410 9875
rect 440 9845 445 9875
rect 605 9875 645 9885
rect 605 9845 610 9875
rect 640 9845 645 9875
rect 805 9875 845 9885
rect 805 9845 810 9875
rect 840 9845 845 9875
rect 1005 9875 1045 9885
rect 1005 9845 1010 9875
rect 1040 9845 1045 9875
rect 1205 9875 1245 9885
rect 1205 9845 1210 9875
rect 1240 9845 1245 9875
rect 1405 9875 1445 9885
rect 1405 9845 1410 9875
rect 1440 9845 1445 9875
rect 1605 9875 1645 9885
rect 1605 9845 1610 9875
rect 1640 9845 1645 9875
rect 1805 9875 1845 9885
rect 1805 9845 1810 9875
rect 1840 9845 1845 9875
rect 2005 9875 2045 9885
rect 2005 9845 2010 9875
rect 2040 9845 2045 9875
rect 2205 9875 2245 9885
rect 2205 9845 2210 9875
rect 2240 9845 2245 9875
rect 2405 9875 2445 9885
rect 2405 9845 2410 9875
rect 2440 9845 2445 9875
rect 2605 9875 2645 9885
rect 2605 9845 2610 9875
rect 2640 9845 2645 9875
rect 2805 9875 2845 9885
rect 2805 9845 2810 9875
rect 2840 9845 2845 9875
rect 3005 9875 3045 9885
rect 3005 9845 3010 9875
rect 3040 9845 3045 9875
rect 3205 9875 3245 9885
rect 3205 9845 3210 9875
rect 3240 9845 3245 9875
rect 3405 9875 3445 9885
rect 3405 9845 3410 9875
rect 3440 9845 3445 9875
rect 3605 9875 3645 9885
rect 3605 9845 3610 9875
rect 3640 9845 3645 9875
rect 3805 9875 3845 9885
rect 3805 9845 3810 9875
rect 3840 9845 3845 9875
rect 4005 9875 4045 9885
rect 4005 9845 4010 9875
rect 4040 9845 4045 9875
rect 4205 9875 4245 9885
rect 4205 9845 4210 9875
rect 4240 9845 4245 9875
rect 4405 9875 4445 9885
rect 4405 9845 4410 9875
rect 4440 9845 4445 9875
rect 4605 9875 4645 9885
rect 4605 9845 4610 9875
rect 4640 9845 4645 9875
rect 4805 9875 4845 9885
rect 4805 9845 4810 9875
rect 4840 9845 4845 9875
rect 5005 9875 5045 9885
rect 5005 9845 5010 9875
rect 5040 9845 5045 9875
rect 5205 9875 5245 9885
rect 5205 9845 5210 9875
rect 5240 9845 5245 9875
rect 5405 9875 5445 9885
rect 5405 9845 5410 9875
rect 5440 9845 5445 9875
rect 5605 9875 5645 9885
rect 5605 9845 5610 9875
rect 5640 9845 5645 9875
rect 5805 9875 5845 9885
rect 5805 9845 5810 9875
rect 5840 9845 5845 9875
rect 6005 9875 6045 9885
rect 6005 9845 6010 9875
rect 6040 9845 6045 9875
rect 6205 9875 6245 9885
rect 6205 9845 6210 9875
rect 6240 9845 6245 9875
rect 6405 9875 6445 9885
rect 6405 9845 6410 9875
rect 6440 9845 6445 9875
rect -188 9760 -185 9845
rect -165 9760 -162 9845
rect 15 9760 35 9845
rect 215 9760 235 9845
rect 415 9760 435 9845
rect 615 9760 635 9845
rect 815 9760 835 9845
rect 1015 9760 1035 9845
rect 1215 9760 1235 9845
rect 1415 9760 1435 9845
rect -195 9730 -190 9760
rect -160 9730 -155 9760
rect -195 9690 -185 9730
rect -165 9720 -155 9730
rect 5 9730 10 9760
rect 40 9730 45 9760
rect 5 9720 45 9730
rect 205 9730 210 9760
rect 240 9730 245 9760
rect 205 9720 245 9730
rect 405 9730 410 9760
rect 440 9730 445 9760
rect 405 9720 445 9730
rect 605 9730 610 9760
rect 640 9730 645 9760
rect 605 9720 645 9730
rect 805 9730 810 9760
rect 840 9730 845 9760
rect 805 9720 845 9730
rect 1005 9730 1010 9760
rect 1040 9730 1045 9760
rect 1005 9720 1045 9730
rect 1205 9730 1210 9760
rect 1240 9730 1245 9760
rect 1205 9720 1245 9730
rect 1405 9730 1410 9760
rect 1440 9730 1445 9760
rect 1405 9720 1445 9730
rect 1605 9730 1610 9760
rect 1640 9730 1645 9760
rect 1605 9720 1645 9730
rect 1805 9730 1810 9760
rect 1840 9730 1845 9760
rect 1805 9720 1845 9730
rect 2005 9730 2010 9760
rect 2040 9730 2045 9760
rect 2005 9720 2045 9730
rect 2205 9730 2210 9760
rect 2240 9730 2245 9760
rect 2205 9720 2245 9730
rect 2405 9730 2410 9760
rect 2440 9730 2445 9760
rect 2405 9720 2445 9730
rect 2605 9730 2610 9760
rect 2640 9730 2645 9760
rect 2605 9720 2645 9730
rect 2805 9730 2810 9760
rect 2840 9730 2845 9760
rect 2805 9720 2845 9730
rect 3005 9730 3010 9760
rect 3040 9730 3045 9760
rect 3005 9720 3045 9730
rect 3205 9730 3210 9760
rect 3240 9730 3245 9760
rect 3205 9720 3245 9730
rect 3405 9730 3410 9760
rect 3440 9730 3445 9760
rect 3405 9720 3445 9730
rect 3605 9730 3610 9760
rect 3640 9730 3645 9760
rect 3605 9720 3645 9730
rect 3805 9730 3810 9760
rect 3840 9730 3845 9760
rect 3805 9720 3845 9730
rect 4005 9730 4010 9760
rect 4040 9730 4045 9760
rect 4005 9720 4045 9730
rect 4205 9730 4210 9760
rect 4240 9730 4245 9760
rect 4205 9720 4245 9730
rect 4405 9730 4410 9760
rect 4440 9730 4445 9760
rect 4405 9720 4445 9730
rect 4605 9730 4610 9760
rect 4640 9730 4645 9760
rect 4605 9720 4645 9730
rect 4805 9730 4810 9760
rect 4840 9730 4845 9760
rect 4805 9720 4845 9730
rect 5005 9730 5010 9760
rect 5040 9730 5045 9760
rect 5005 9720 5045 9730
rect 5205 9730 5210 9760
rect 5240 9730 5245 9760
rect 5205 9720 5245 9730
rect 5405 9730 5410 9760
rect 5440 9730 5445 9760
rect 5405 9720 5445 9730
rect 5605 9730 5610 9760
rect 5640 9730 5645 9760
rect 5605 9720 5645 9730
rect 5805 9730 5810 9760
rect 5840 9730 5845 9760
rect 5805 9720 5845 9730
rect 6005 9730 6010 9760
rect 6040 9730 6045 9760
rect 6005 9720 6045 9730
rect 6205 9730 6210 9760
rect 6240 9730 6245 9760
rect 6205 9720 6245 9730
rect 6405 9730 6410 9760
rect 6440 9730 6445 9760
rect 6405 9720 6445 9730
rect -165 9700 -30 9720
rect 5 9700 1570 9720
rect 1605 9700 6570 9720
rect -165 9690 -155 9700
rect -195 9660 -190 9690
rect -160 9660 -155 9690
rect 5 9690 45 9700
rect 5 9660 10 9690
rect 40 9660 45 9690
rect 205 9690 245 9700
rect 205 9660 210 9690
rect 240 9660 245 9690
rect 405 9690 445 9700
rect 405 9660 410 9690
rect 440 9660 445 9690
rect 605 9690 645 9700
rect 605 9660 610 9690
rect 640 9660 645 9690
rect 805 9690 845 9700
rect 805 9660 810 9690
rect 840 9660 845 9690
rect 1005 9690 1045 9700
rect 1005 9660 1010 9690
rect 1040 9660 1045 9690
rect 1205 9690 1245 9700
rect 1205 9660 1210 9690
rect 1240 9660 1245 9690
rect 1405 9690 1445 9700
rect 1405 9660 1410 9690
rect 1440 9660 1445 9690
rect 1605 9690 1645 9700
rect 1605 9660 1610 9690
rect 1640 9660 1645 9690
rect 1805 9690 1845 9700
rect 1805 9660 1810 9690
rect 1840 9660 1845 9690
rect 2005 9690 2045 9700
rect 2005 9660 2010 9690
rect 2040 9660 2045 9690
rect 2205 9690 2245 9700
rect 2205 9660 2210 9690
rect 2240 9660 2245 9690
rect 2405 9690 2445 9700
rect 2405 9660 2410 9690
rect 2440 9660 2445 9690
rect 2605 9690 2645 9700
rect 2605 9660 2610 9690
rect 2640 9660 2645 9690
rect 2805 9690 2845 9700
rect 2805 9660 2810 9690
rect 2840 9660 2845 9690
rect 3005 9690 3045 9700
rect 3005 9660 3010 9690
rect 3040 9660 3045 9690
rect 3205 9690 3245 9700
rect 3205 9660 3210 9690
rect 3240 9660 3245 9690
rect 3405 9690 3445 9700
rect 3405 9660 3410 9690
rect 3440 9660 3445 9690
rect 3605 9690 3645 9700
rect 3605 9660 3610 9690
rect 3640 9660 3645 9690
rect 3805 9690 3845 9700
rect 3805 9660 3810 9690
rect 3840 9660 3845 9690
rect 4005 9690 4045 9700
rect 4005 9660 4010 9690
rect 4040 9660 4045 9690
rect 4205 9690 4245 9700
rect 4205 9660 4210 9690
rect 4240 9660 4245 9690
rect 4405 9690 4445 9700
rect 4405 9660 4410 9690
rect 4440 9660 4445 9690
rect 4605 9690 4645 9700
rect 4605 9660 4610 9690
rect 4640 9660 4645 9690
rect 4805 9690 4845 9700
rect 4805 9660 4810 9690
rect 4840 9660 4845 9690
rect 5005 9690 5045 9700
rect 5005 9660 5010 9690
rect 5040 9660 5045 9690
rect 5205 9690 5245 9700
rect 5205 9660 5210 9690
rect 5240 9660 5245 9690
rect 5405 9690 5445 9700
rect 5405 9660 5410 9690
rect 5440 9660 5445 9690
rect 5605 9690 5645 9700
rect 5605 9660 5610 9690
rect 5640 9660 5645 9690
rect 5805 9690 5845 9700
rect 5805 9660 5810 9690
rect 5840 9660 5845 9690
rect 6005 9690 6045 9700
rect 6005 9660 6010 9690
rect 6040 9660 6045 9690
rect 6205 9690 6245 9700
rect 6205 9660 6210 9690
rect 6240 9660 6245 9690
rect 6405 9690 6445 9700
rect 6405 9660 6410 9690
rect 6440 9660 6445 9690
rect -188 9575 -185 9660
rect -165 9575 -162 9660
rect 15 9575 35 9660
rect 215 9575 235 9660
rect 415 9575 435 9660
rect 615 9575 635 9660
rect 815 9575 835 9660
rect 1015 9575 1035 9660
rect 1215 9575 1235 9660
rect 1415 9575 1435 9660
rect 1615 9575 1635 9660
rect 1815 9575 1835 9660
rect 2015 9575 2035 9660
rect 2215 9575 2235 9660
rect 2415 9575 2435 9660
rect 2615 9575 2635 9660
rect 2815 9575 2835 9660
rect 3015 9575 3035 9660
rect 3215 9575 3235 9660
rect 3415 9575 3435 9660
rect 3615 9575 3635 9660
rect 3815 9575 3835 9660
rect 4015 9575 4035 9660
rect 4215 9575 4235 9660
rect 4415 9575 4435 9660
rect 4615 9575 4635 9660
rect 4815 9575 4835 9660
rect 5015 9575 5035 9660
rect 5215 9575 5235 9660
rect 5415 9575 5435 9660
rect 5615 9575 5635 9660
rect 5815 9575 5835 9660
rect 6015 9575 6035 9660
rect 6215 9575 6235 9660
rect -195 9545 -190 9575
rect -160 9545 -155 9575
rect -195 9505 -185 9545
rect -165 9535 -155 9545
rect 5 9545 10 9575
rect 40 9545 45 9575
rect 5 9535 45 9545
rect 205 9545 210 9575
rect 240 9545 245 9575
rect 205 9535 245 9545
rect 405 9545 410 9575
rect 440 9545 445 9575
rect 405 9535 445 9545
rect 605 9545 610 9575
rect 640 9545 645 9575
rect 605 9535 645 9545
rect 805 9545 810 9575
rect 840 9545 845 9575
rect 805 9535 845 9545
rect 1005 9545 1010 9575
rect 1040 9545 1045 9575
rect 1005 9535 1045 9545
rect 1205 9545 1210 9575
rect 1240 9545 1245 9575
rect 1205 9535 1245 9545
rect 1405 9545 1410 9575
rect 1440 9545 1445 9575
rect 1405 9535 1445 9545
rect 1605 9545 1610 9575
rect 1640 9545 1645 9575
rect 1605 9535 1645 9545
rect 1805 9545 1810 9575
rect 1840 9545 1845 9575
rect 1805 9535 1845 9545
rect 2005 9545 2010 9575
rect 2040 9545 2045 9575
rect 2005 9535 2045 9545
rect 2205 9545 2210 9575
rect 2240 9545 2245 9575
rect 2205 9535 2245 9545
rect 2405 9545 2410 9575
rect 2440 9545 2445 9575
rect 2405 9535 2445 9545
rect 2605 9545 2610 9575
rect 2640 9545 2645 9575
rect 2605 9535 2645 9545
rect 2805 9545 2810 9575
rect 2840 9545 2845 9575
rect 2805 9535 2845 9545
rect 3005 9545 3010 9575
rect 3040 9545 3045 9575
rect 3005 9535 3045 9545
rect 3205 9545 3210 9575
rect 3240 9545 3245 9575
rect 3205 9535 3245 9545
rect 3405 9545 3410 9575
rect 3440 9545 3445 9575
rect 3405 9535 3445 9545
rect 3605 9545 3610 9575
rect 3640 9545 3645 9575
rect 3605 9535 3645 9545
rect 3805 9545 3810 9575
rect 3840 9545 3845 9575
rect 3805 9535 3845 9545
rect 4005 9545 4010 9575
rect 4040 9545 4045 9575
rect 4005 9535 4045 9545
rect 4205 9545 4210 9575
rect 4240 9545 4245 9575
rect 4205 9535 4245 9545
rect 4405 9545 4410 9575
rect 4440 9545 4445 9575
rect 4405 9535 4445 9545
rect 4605 9545 4610 9575
rect 4640 9545 4645 9575
rect 4605 9535 4645 9545
rect 4805 9545 4810 9575
rect 4840 9545 4845 9575
rect 4805 9535 4845 9545
rect 5005 9545 5010 9575
rect 5040 9545 5045 9575
rect 5005 9535 5045 9545
rect 5205 9545 5210 9575
rect 5240 9545 5245 9575
rect 5205 9535 5245 9545
rect 5405 9545 5410 9575
rect 5440 9545 5445 9575
rect 5405 9535 5445 9545
rect 5605 9545 5610 9575
rect 5640 9545 5645 9575
rect 5605 9535 5645 9545
rect 5805 9545 5810 9575
rect 5840 9545 5845 9575
rect 5805 9535 5845 9545
rect 6005 9545 6010 9575
rect 6040 9545 6045 9575
rect 6005 9535 6045 9545
rect 6205 9545 6210 9575
rect 6240 9545 6245 9575
rect 6205 9535 6245 9545
rect 6405 9545 6410 9575
rect 6440 9545 6445 9575
rect 6405 9535 6445 9545
rect -165 9515 -30 9535
rect 5 9515 1570 9535
rect 1605 9515 6570 9535
rect -165 9505 -155 9515
rect -195 9475 -190 9505
rect -160 9475 -155 9505
rect 5 9505 45 9515
rect 5 9475 10 9505
rect 40 9475 45 9505
rect 205 9505 245 9515
rect 205 9475 210 9505
rect 240 9475 245 9505
rect 405 9505 445 9515
rect 405 9475 410 9505
rect 440 9475 445 9505
rect 605 9505 645 9515
rect 605 9475 610 9505
rect 640 9475 645 9505
rect 805 9505 845 9515
rect 805 9475 810 9505
rect 840 9475 845 9505
rect 1005 9505 1045 9515
rect 1005 9475 1010 9505
rect 1040 9475 1045 9505
rect 1205 9505 1245 9515
rect 1205 9475 1210 9505
rect 1240 9475 1245 9505
rect 1405 9505 1445 9515
rect 1405 9475 1410 9505
rect 1440 9475 1445 9505
rect 1605 9505 1645 9515
rect 1605 9475 1610 9505
rect 1640 9475 1645 9505
rect 1805 9505 1845 9515
rect 1805 9475 1810 9505
rect 1840 9475 1845 9505
rect 2005 9505 2045 9515
rect 2005 9475 2010 9505
rect 2040 9475 2045 9505
rect 2205 9505 2245 9515
rect 2205 9475 2210 9505
rect 2240 9475 2245 9505
rect 2405 9505 2445 9515
rect 2405 9475 2410 9505
rect 2440 9475 2445 9505
rect 2605 9505 2645 9515
rect 2605 9475 2610 9505
rect 2640 9475 2645 9505
rect 2805 9505 2845 9515
rect 2805 9475 2810 9505
rect 2840 9475 2845 9505
rect 3005 9505 3045 9515
rect 3005 9475 3010 9505
rect 3040 9475 3045 9505
rect 3205 9505 3245 9515
rect 3205 9475 3210 9505
rect 3240 9475 3245 9505
rect 3405 9505 3445 9515
rect 3405 9475 3410 9505
rect 3440 9475 3445 9505
rect 3605 9505 3645 9515
rect 3605 9475 3610 9505
rect 3640 9475 3645 9505
rect 3805 9505 3845 9515
rect 3805 9475 3810 9505
rect 3840 9475 3845 9505
rect 4005 9505 4045 9515
rect 4005 9475 4010 9505
rect 4040 9475 4045 9505
rect 4205 9505 4245 9515
rect 4205 9475 4210 9505
rect 4240 9475 4245 9505
rect 4405 9505 4445 9515
rect 4405 9475 4410 9505
rect 4440 9475 4445 9505
rect 4605 9505 4645 9515
rect 4605 9475 4610 9505
rect 4640 9475 4645 9505
rect 4805 9505 4845 9515
rect 4805 9475 4810 9505
rect 4840 9475 4845 9505
rect 5005 9505 5045 9515
rect 5005 9475 5010 9505
rect 5040 9475 5045 9505
rect 5205 9505 5245 9515
rect 5205 9475 5210 9505
rect 5240 9475 5245 9505
rect 5405 9505 5445 9515
rect 5405 9475 5410 9505
rect 5440 9475 5445 9505
rect 5605 9505 5645 9515
rect 5605 9475 5610 9505
rect 5640 9475 5645 9505
rect 5805 9505 5845 9515
rect 5805 9475 5810 9505
rect 5840 9475 5845 9505
rect 6005 9505 6045 9515
rect 6005 9475 6010 9505
rect 6040 9475 6045 9505
rect 6205 9505 6245 9515
rect 6205 9475 6210 9505
rect 6240 9475 6245 9505
rect 6405 9505 6445 9515
rect 6405 9475 6410 9505
rect 6440 9475 6445 9505
rect -188 9390 -185 9475
rect -165 9390 -162 9475
rect 15 9390 35 9475
rect 215 9390 235 9475
rect 415 9390 435 9475
rect 615 9390 635 9475
rect 815 9390 835 9475
rect 1015 9390 1035 9475
rect 1215 9390 1235 9475
rect 1415 9390 1435 9475
rect 1615 9390 1635 9475
rect 1815 9390 1835 9475
rect 2015 9390 2035 9475
rect 2215 9390 2235 9475
rect 2415 9390 2435 9475
rect 2615 9390 2635 9475
rect 2815 9390 2835 9475
rect 3015 9390 3035 9475
rect 3215 9390 3235 9475
rect 3415 9390 3435 9475
rect 3615 9390 3635 9475
rect 3815 9390 3835 9475
rect 4015 9390 4035 9475
rect 4215 9390 4235 9475
rect 4415 9390 4435 9475
rect 4615 9390 4635 9475
rect 4815 9390 4835 9475
rect 5015 9390 5035 9475
rect 5215 9390 5235 9475
rect 5415 9390 5435 9475
rect 5615 9390 5635 9475
rect 5815 9390 5835 9475
rect 6015 9390 6035 9475
rect 6215 9390 6235 9475
rect -195 9360 -190 9390
rect -160 9360 -155 9390
rect -195 9320 -185 9360
rect -165 9350 -155 9360
rect 5 9360 10 9390
rect 40 9360 45 9390
rect 5 9350 45 9360
rect 205 9360 210 9390
rect 240 9360 245 9390
rect 205 9350 245 9360
rect 405 9360 410 9390
rect 440 9360 445 9390
rect 405 9350 445 9360
rect 605 9360 610 9390
rect 640 9360 645 9390
rect 605 9350 645 9360
rect 805 9360 810 9390
rect 840 9360 845 9390
rect 805 9350 845 9360
rect 1005 9360 1010 9390
rect 1040 9360 1045 9390
rect 1005 9350 1045 9360
rect 1205 9360 1210 9390
rect 1240 9360 1245 9390
rect 1205 9350 1245 9360
rect 1405 9360 1410 9390
rect 1440 9360 1445 9390
rect 1405 9350 1445 9360
rect 1605 9360 1610 9390
rect 1640 9360 1645 9390
rect 1605 9350 1645 9360
rect 1805 9360 1810 9390
rect 1840 9360 1845 9390
rect 1805 9350 1845 9360
rect 2005 9360 2010 9390
rect 2040 9360 2045 9390
rect 2005 9350 2045 9360
rect 2205 9360 2210 9390
rect 2240 9360 2245 9390
rect 2205 9350 2245 9360
rect 2405 9360 2410 9390
rect 2440 9360 2445 9390
rect 2405 9350 2445 9360
rect 2605 9360 2610 9390
rect 2640 9360 2645 9390
rect 2605 9350 2645 9360
rect 2805 9360 2810 9390
rect 2840 9360 2845 9390
rect 2805 9350 2845 9360
rect 3005 9360 3010 9390
rect 3040 9360 3045 9390
rect 3005 9350 3045 9360
rect 3205 9360 3210 9390
rect 3240 9360 3245 9390
rect 3205 9350 3245 9360
rect 3405 9360 3410 9390
rect 3440 9360 3445 9390
rect 3405 9350 3445 9360
rect 3605 9360 3610 9390
rect 3640 9360 3645 9390
rect 3605 9350 3645 9360
rect 3805 9360 3810 9390
rect 3840 9360 3845 9390
rect 3805 9350 3845 9360
rect 4005 9360 4010 9390
rect 4040 9360 4045 9390
rect 4005 9350 4045 9360
rect 4205 9360 4210 9390
rect 4240 9360 4245 9390
rect 4205 9350 4245 9360
rect 4405 9360 4410 9390
rect 4440 9360 4445 9390
rect 4405 9350 4445 9360
rect 4605 9360 4610 9390
rect 4640 9360 4645 9390
rect 4605 9350 4645 9360
rect 4805 9360 4810 9390
rect 4840 9360 4845 9390
rect 4805 9350 4845 9360
rect 5005 9360 5010 9390
rect 5040 9360 5045 9390
rect 5005 9350 5045 9360
rect 5205 9360 5210 9390
rect 5240 9360 5245 9390
rect 5205 9350 5245 9360
rect 5405 9360 5410 9390
rect 5440 9360 5445 9390
rect 5405 9350 5445 9360
rect 5605 9360 5610 9390
rect 5640 9360 5645 9390
rect 5605 9350 5645 9360
rect 5805 9360 5810 9390
rect 5840 9360 5845 9390
rect 5805 9350 5845 9360
rect 6005 9360 6010 9390
rect 6040 9360 6045 9390
rect 6005 9350 6045 9360
rect 6205 9360 6210 9390
rect 6240 9360 6245 9390
rect 6205 9350 6245 9360
rect 6405 9360 6410 9390
rect 6440 9360 6445 9390
rect 6405 9350 6445 9360
rect -165 9330 -30 9350
rect 5 9330 1570 9350
rect 1605 9330 6570 9350
rect -165 9320 -155 9330
rect -195 9290 -190 9320
rect -160 9290 -155 9320
rect 5 9320 45 9330
rect 5 9290 10 9320
rect 40 9290 45 9320
rect 205 9320 245 9330
rect 205 9290 210 9320
rect 240 9290 245 9320
rect 405 9320 445 9330
rect 405 9290 410 9320
rect 440 9290 445 9320
rect 605 9320 645 9330
rect 605 9290 610 9320
rect 640 9290 645 9320
rect 805 9320 845 9330
rect 805 9290 810 9320
rect 840 9290 845 9320
rect 1005 9320 1045 9330
rect 1005 9290 1010 9320
rect 1040 9290 1045 9320
rect 1205 9320 1245 9330
rect 1205 9290 1210 9320
rect 1240 9290 1245 9320
rect 1405 9320 1445 9330
rect 1405 9290 1410 9320
rect 1440 9290 1445 9320
rect 1605 9320 1645 9330
rect 1605 9290 1610 9320
rect 1640 9290 1645 9320
rect 1805 9320 1845 9330
rect 1805 9290 1810 9320
rect 1840 9290 1845 9320
rect 2005 9320 2045 9330
rect 2005 9290 2010 9320
rect 2040 9290 2045 9320
rect 2205 9320 2245 9330
rect 2205 9290 2210 9320
rect 2240 9290 2245 9320
rect 2405 9320 2445 9330
rect 2405 9290 2410 9320
rect 2440 9290 2445 9320
rect 2605 9320 2645 9330
rect 2605 9290 2610 9320
rect 2640 9290 2645 9320
rect 2805 9320 2845 9330
rect 2805 9290 2810 9320
rect 2840 9290 2845 9320
rect 3005 9320 3045 9330
rect 3005 9290 3010 9320
rect 3040 9290 3045 9320
rect 3205 9320 3245 9330
rect 3205 9290 3210 9320
rect 3240 9290 3245 9320
rect 3405 9320 3445 9330
rect 3405 9290 3410 9320
rect 3440 9290 3445 9320
rect 3605 9320 3645 9330
rect 3605 9290 3610 9320
rect 3640 9290 3645 9320
rect 3805 9320 3845 9330
rect 3805 9290 3810 9320
rect 3840 9290 3845 9320
rect 4005 9320 4045 9330
rect 4005 9290 4010 9320
rect 4040 9290 4045 9320
rect 4205 9320 4245 9330
rect 4205 9290 4210 9320
rect 4240 9290 4245 9320
rect 4405 9320 4445 9330
rect 4405 9290 4410 9320
rect 4440 9290 4445 9320
rect 4605 9320 4645 9330
rect 4605 9290 4610 9320
rect 4640 9290 4645 9320
rect 4805 9320 4845 9330
rect 4805 9290 4810 9320
rect 4840 9290 4845 9320
rect 5005 9320 5045 9330
rect 5005 9290 5010 9320
rect 5040 9290 5045 9320
rect 5205 9320 5245 9330
rect 5205 9290 5210 9320
rect 5240 9290 5245 9320
rect 5405 9320 5445 9330
rect 5405 9290 5410 9320
rect 5440 9290 5445 9320
rect 5605 9320 5645 9330
rect 5605 9290 5610 9320
rect 5640 9290 5645 9320
rect 5805 9320 5845 9330
rect 5805 9290 5810 9320
rect 5840 9290 5845 9320
rect 6005 9320 6045 9330
rect 6005 9290 6010 9320
rect 6040 9290 6045 9320
rect 6205 9320 6245 9330
rect 6205 9290 6210 9320
rect 6240 9290 6245 9320
rect 6405 9320 6445 9330
rect 6405 9290 6410 9320
rect 6440 9290 6445 9320
rect -188 9205 -185 9290
rect -165 9205 -162 9290
rect 15 9205 35 9290
rect 215 9205 235 9290
rect 415 9205 435 9290
rect 615 9205 635 9290
rect 815 9205 835 9290
rect 1015 9205 1035 9290
rect 1215 9205 1235 9290
rect 1415 9205 1435 9290
rect 1615 9205 1635 9290
rect 1815 9205 1835 9290
rect 2015 9205 2035 9290
rect 2215 9205 2235 9290
rect 2415 9205 2435 9290
rect 2615 9205 2635 9290
rect 2815 9205 2835 9290
rect 3015 9205 3035 9290
rect 3215 9205 3235 9290
rect 3415 9205 3435 9290
rect 3615 9205 3635 9290
rect 3815 9205 3835 9290
rect 4015 9205 4035 9290
rect 4215 9205 4235 9290
rect 4415 9205 4435 9290
rect 4615 9205 4635 9290
rect 4815 9205 4835 9290
rect 5015 9205 5035 9290
rect 5215 9205 5235 9290
rect 5415 9205 5435 9290
rect 5615 9205 5635 9290
rect 5815 9205 5835 9290
rect 6015 9205 6035 9290
rect 6215 9205 6235 9290
rect -195 9175 -190 9205
rect -160 9175 -155 9205
rect -195 9135 -185 9175
rect -165 9165 -155 9175
rect 5 9175 10 9205
rect 40 9175 45 9205
rect 5 9165 45 9175
rect 205 9175 210 9205
rect 240 9175 245 9205
rect 205 9165 245 9175
rect 405 9175 410 9205
rect 440 9175 445 9205
rect 405 9165 445 9175
rect 605 9175 610 9205
rect 640 9175 645 9205
rect 605 9165 645 9175
rect 805 9175 810 9205
rect 840 9175 845 9205
rect 805 9165 845 9175
rect 1005 9175 1010 9205
rect 1040 9175 1045 9205
rect 1005 9165 1045 9175
rect 1205 9175 1210 9205
rect 1240 9175 1245 9205
rect 1205 9165 1245 9175
rect 1405 9175 1410 9205
rect 1440 9175 1445 9205
rect 1405 9165 1445 9175
rect 1605 9175 1610 9205
rect 1640 9175 1645 9205
rect 1605 9165 1645 9175
rect 1805 9175 1810 9205
rect 1840 9175 1845 9205
rect 1805 9165 1845 9175
rect 2005 9175 2010 9205
rect 2040 9175 2045 9205
rect 2005 9165 2045 9175
rect 2205 9175 2210 9205
rect 2240 9175 2245 9205
rect 2205 9165 2245 9175
rect 2405 9175 2410 9205
rect 2440 9175 2445 9205
rect 2405 9165 2445 9175
rect 2605 9175 2610 9205
rect 2640 9175 2645 9205
rect 2605 9165 2645 9175
rect 2805 9175 2810 9205
rect 2840 9175 2845 9205
rect 2805 9165 2845 9175
rect 3005 9175 3010 9205
rect 3040 9175 3045 9205
rect 3005 9165 3045 9175
rect 3205 9175 3210 9205
rect 3240 9175 3245 9205
rect 3205 9165 3245 9175
rect 3405 9175 3410 9205
rect 3440 9175 3445 9205
rect 3405 9165 3445 9175
rect 3605 9175 3610 9205
rect 3640 9175 3645 9205
rect 3605 9165 3645 9175
rect 3805 9175 3810 9205
rect 3840 9175 3845 9205
rect 3805 9165 3845 9175
rect 4005 9175 4010 9205
rect 4040 9175 4045 9205
rect 4005 9165 4045 9175
rect 4205 9175 4210 9205
rect 4240 9175 4245 9205
rect 4205 9165 4245 9175
rect 4405 9175 4410 9205
rect 4440 9175 4445 9205
rect 4405 9165 4445 9175
rect 4605 9175 4610 9205
rect 4640 9175 4645 9205
rect 4605 9165 4645 9175
rect 4805 9175 4810 9205
rect 4840 9175 4845 9205
rect 4805 9165 4845 9175
rect 5005 9175 5010 9205
rect 5040 9175 5045 9205
rect 5005 9165 5045 9175
rect 5205 9175 5210 9205
rect 5240 9175 5245 9205
rect 5205 9165 5245 9175
rect 5405 9175 5410 9205
rect 5440 9175 5445 9205
rect 5405 9165 5445 9175
rect 5605 9175 5610 9205
rect 5640 9175 5645 9205
rect 5605 9165 5645 9175
rect 5805 9175 5810 9205
rect 5840 9175 5845 9205
rect 5805 9165 5845 9175
rect 6005 9175 6010 9205
rect 6040 9175 6045 9205
rect 6005 9165 6045 9175
rect 6205 9175 6210 9205
rect 6240 9175 6245 9205
rect 6205 9165 6245 9175
rect 6405 9175 6410 9205
rect 6440 9175 6445 9205
rect 6405 9165 6445 9175
rect -165 9145 -30 9165
rect 5 9145 1570 9165
rect 1605 9145 6570 9165
rect -165 9135 -155 9145
rect -195 9105 -190 9135
rect -160 9105 -155 9135
rect 5 9135 45 9145
rect 5 9105 10 9135
rect 40 9105 45 9135
rect 205 9135 245 9145
rect 205 9105 210 9135
rect 240 9105 245 9135
rect 405 9135 445 9145
rect 405 9105 410 9135
rect 440 9105 445 9135
rect 605 9135 645 9145
rect 605 9105 610 9135
rect 640 9105 645 9135
rect 805 9135 845 9145
rect 805 9105 810 9135
rect 840 9105 845 9135
rect 1005 9135 1045 9145
rect 1005 9105 1010 9135
rect 1040 9105 1045 9135
rect 1205 9135 1245 9145
rect 1205 9105 1210 9135
rect 1240 9105 1245 9135
rect 1405 9135 1445 9145
rect 1405 9105 1410 9135
rect 1440 9105 1445 9135
rect 1605 9135 1645 9145
rect 1605 9105 1610 9135
rect 1640 9105 1645 9135
rect 1805 9135 1845 9145
rect 1805 9105 1810 9135
rect 1840 9105 1845 9135
rect 2005 9135 2045 9145
rect 2005 9105 2010 9135
rect 2040 9105 2045 9135
rect 2205 9135 2245 9145
rect 2205 9105 2210 9135
rect 2240 9105 2245 9135
rect 2405 9135 2445 9145
rect 2405 9105 2410 9135
rect 2440 9105 2445 9135
rect 2605 9135 2645 9145
rect 2605 9105 2610 9135
rect 2640 9105 2645 9135
rect 2805 9135 2845 9145
rect 2805 9105 2810 9135
rect 2840 9105 2845 9135
rect 3005 9135 3045 9145
rect 3005 9105 3010 9135
rect 3040 9105 3045 9135
rect 3205 9135 3245 9145
rect 3205 9105 3210 9135
rect 3240 9105 3245 9135
rect 3405 9135 3445 9145
rect 3405 9105 3410 9135
rect 3440 9105 3445 9135
rect 3605 9135 3645 9145
rect 3605 9105 3610 9135
rect 3640 9105 3645 9135
rect 3805 9135 3845 9145
rect 3805 9105 3810 9135
rect 3840 9105 3845 9135
rect 4005 9135 4045 9145
rect 4005 9105 4010 9135
rect 4040 9105 4045 9135
rect 4205 9135 4245 9145
rect 4205 9105 4210 9135
rect 4240 9105 4245 9135
rect 4405 9135 4445 9145
rect 4405 9105 4410 9135
rect 4440 9105 4445 9135
rect 4605 9135 4645 9145
rect 4605 9105 4610 9135
rect 4640 9105 4645 9135
rect 4805 9135 4845 9145
rect 4805 9105 4810 9135
rect 4840 9105 4845 9135
rect 5005 9135 5045 9145
rect 5005 9105 5010 9135
rect 5040 9105 5045 9135
rect 5205 9135 5245 9145
rect 5205 9105 5210 9135
rect 5240 9105 5245 9135
rect 5405 9135 5445 9145
rect 5405 9105 5410 9135
rect 5440 9105 5445 9135
rect 5605 9135 5645 9145
rect 5605 9105 5610 9135
rect 5640 9105 5645 9135
rect 5805 9135 5845 9145
rect 5805 9105 5810 9135
rect 5840 9105 5845 9135
rect 6005 9135 6045 9145
rect 6005 9105 6010 9135
rect 6040 9105 6045 9135
rect 6205 9135 6245 9145
rect 6205 9105 6210 9135
rect 6240 9105 6245 9135
rect 6405 9135 6445 9145
rect 6405 9105 6410 9135
rect 6440 9105 6445 9135
rect -188 9020 -185 9105
rect -165 9020 -162 9105
rect 15 9020 35 9105
rect 215 9020 235 9105
rect 415 9020 435 9105
rect 615 9020 635 9105
rect 815 9020 835 9105
rect 1015 9020 1035 9105
rect 1215 9020 1235 9105
rect 1415 9020 1435 9105
rect 1615 9020 1635 9105
rect 1815 9020 1835 9105
rect 2015 9020 2035 9105
rect 2215 9020 2235 9105
rect 2415 9020 2435 9105
rect 2615 9020 2635 9105
rect 2815 9020 2835 9105
rect 3015 9020 3035 9105
rect 3215 9020 3235 9105
rect 3415 9020 3435 9105
rect 3615 9020 3635 9105
rect 3815 9020 3835 9105
rect 4015 9020 4035 9105
rect 4215 9020 4235 9105
rect 4415 9020 4435 9105
rect 4615 9020 4635 9105
rect 4815 9020 4835 9105
rect 5015 9020 5035 9105
rect 5215 9020 5235 9105
rect 5415 9020 5435 9105
rect 5615 9020 5635 9105
rect 5815 9020 5835 9105
rect 6015 9020 6035 9105
rect 6215 9020 6235 9105
rect -195 8990 -190 9020
rect -160 8990 -155 9020
rect -195 8950 -185 8990
rect -165 8980 -155 8990
rect 5 8990 10 9020
rect 40 8990 45 9020
rect 5 8980 45 8990
rect 205 8990 210 9020
rect 240 8990 245 9020
rect 205 8980 245 8990
rect 405 8990 410 9020
rect 440 8990 445 9020
rect 405 8980 445 8990
rect 605 8990 610 9020
rect 640 8990 645 9020
rect 605 8980 645 8990
rect 805 8990 810 9020
rect 840 8990 845 9020
rect 805 8980 845 8990
rect 1005 8990 1010 9020
rect 1040 8990 1045 9020
rect 1005 8980 1045 8990
rect 1205 8990 1210 9020
rect 1240 8990 1245 9020
rect 1205 8980 1245 8990
rect 1405 8990 1410 9020
rect 1440 8990 1445 9020
rect 1405 8980 1445 8990
rect 1605 8990 1610 9020
rect 1640 8990 1645 9020
rect 1605 8980 1645 8990
rect 1805 8990 1810 9020
rect 1840 8990 1845 9020
rect 1805 8980 1845 8990
rect 2005 8990 2010 9020
rect 2040 8990 2045 9020
rect 2005 8980 2045 8990
rect 2205 8990 2210 9020
rect 2240 8990 2245 9020
rect 2205 8980 2245 8990
rect 2405 8990 2410 9020
rect 2440 8990 2445 9020
rect 2405 8980 2445 8990
rect 2605 8990 2610 9020
rect 2640 8990 2645 9020
rect 2605 8980 2645 8990
rect 2805 8990 2810 9020
rect 2840 8990 2845 9020
rect 2805 8980 2845 8990
rect 3005 8990 3010 9020
rect 3040 8990 3045 9020
rect 3005 8980 3045 8990
rect 3205 8990 3210 9020
rect 3240 8990 3245 9020
rect 3205 8980 3245 8990
rect 3405 8990 3410 9020
rect 3440 8990 3445 9020
rect 3405 8980 3445 8990
rect 3605 8990 3610 9020
rect 3640 8990 3645 9020
rect 3605 8980 3645 8990
rect 3805 8990 3810 9020
rect 3840 8990 3845 9020
rect 3805 8980 3845 8990
rect 4005 8990 4010 9020
rect 4040 8990 4045 9020
rect 4005 8980 4045 8990
rect 4205 8990 4210 9020
rect 4240 8990 4245 9020
rect 4205 8980 4245 8990
rect 4405 8990 4410 9020
rect 4440 8990 4445 9020
rect 4405 8980 4445 8990
rect 4605 8990 4610 9020
rect 4640 8990 4645 9020
rect 4605 8980 4645 8990
rect 4805 8990 4810 9020
rect 4840 8990 4845 9020
rect 4805 8980 4845 8990
rect 5005 8990 5010 9020
rect 5040 8990 5045 9020
rect 5005 8980 5045 8990
rect 5205 8990 5210 9020
rect 5240 8990 5245 9020
rect 5205 8980 5245 8990
rect 5405 8990 5410 9020
rect 5440 8990 5445 9020
rect 5405 8980 5445 8990
rect 5605 8990 5610 9020
rect 5640 8990 5645 9020
rect 5605 8980 5645 8990
rect 5805 8990 5810 9020
rect 5840 8990 5845 9020
rect 5805 8980 5845 8990
rect 6005 8990 6010 9020
rect 6040 8990 6045 9020
rect 6005 8980 6045 8990
rect 6205 8990 6210 9020
rect 6240 8990 6245 9020
rect 6205 8980 6245 8990
rect 6405 8990 6410 9020
rect 6440 8990 6445 9020
rect 6405 8980 6445 8990
rect -165 8960 -30 8980
rect 5 8960 1570 8980
rect 1605 8960 6570 8980
rect -165 8950 -155 8960
rect -195 8920 -190 8950
rect -160 8920 -155 8950
rect 5 8950 45 8960
rect 5 8920 10 8950
rect 40 8920 45 8950
rect 205 8950 245 8960
rect 205 8920 210 8950
rect 240 8920 245 8950
rect 405 8950 445 8960
rect 405 8920 410 8950
rect 440 8920 445 8950
rect 605 8950 645 8960
rect 605 8920 610 8950
rect 640 8920 645 8950
rect 805 8950 845 8960
rect 805 8920 810 8950
rect 840 8920 845 8950
rect 1005 8950 1045 8960
rect 1005 8920 1010 8950
rect 1040 8920 1045 8950
rect 1205 8950 1245 8960
rect 1205 8920 1210 8950
rect 1240 8920 1245 8950
rect 1405 8950 1445 8960
rect 1405 8920 1410 8950
rect 1440 8920 1445 8950
rect 1605 8950 1645 8960
rect 1605 8920 1610 8950
rect 1640 8920 1645 8950
rect 1805 8950 1845 8960
rect 1805 8920 1810 8950
rect 1840 8920 1845 8950
rect 2005 8950 2045 8960
rect 2005 8920 2010 8950
rect 2040 8920 2045 8950
rect 2205 8950 2245 8960
rect 2205 8920 2210 8950
rect 2240 8920 2245 8950
rect 2405 8950 2445 8960
rect 2405 8920 2410 8950
rect 2440 8920 2445 8950
rect 2605 8950 2645 8960
rect 2605 8920 2610 8950
rect 2640 8920 2645 8950
rect 2805 8950 2845 8960
rect 2805 8920 2810 8950
rect 2840 8920 2845 8950
rect 3005 8950 3045 8960
rect 3005 8920 3010 8950
rect 3040 8920 3045 8950
rect 3205 8950 3245 8960
rect 3205 8920 3210 8950
rect 3240 8920 3245 8950
rect 3405 8950 3445 8960
rect 3405 8920 3410 8950
rect 3440 8920 3445 8950
rect 3605 8950 3645 8960
rect 3605 8920 3610 8950
rect 3640 8920 3645 8950
rect 3805 8950 3845 8960
rect 3805 8920 3810 8950
rect 3840 8920 3845 8950
rect 4005 8950 4045 8960
rect 4005 8920 4010 8950
rect 4040 8920 4045 8950
rect 4205 8950 4245 8960
rect 4205 8920 4210 8950
rect 4240 8920 4245 8950
rect 4405 8950 4445 8960
rect 4405 8920 4410 8950
rect 4440 8920 4445 8950
rect 4605 8950 4645 8960
rect 4605 8920 4610 8950
rect 4640 8920 4645 8950
rect 4805 8950 4845 8960
rect 4805 8920 4810 8950
rect 4840 8920 4845 8950
rect 5005 8950 5045 8960
rect 5005 8920 5010 8950
rect 5040 8920 5045 8950
rect 5205 8950 5245 8960
rect 5205 8920 5210 8950
rect 5240 8920 5245 8950
rect 5405 8950 5445 8960
rect 5405 8920 5410 8950
rect 5440 8920 5445 8950
rect 5605 8950 5645 8960
rect 5605 8920 5610 8950
rect 5640 8920 5645 8950
rect 5805 8950 5845 8960
rect 5805 8920 5810 8950
rect 5840 8920 5845 8950
rect 6005 8950 6045 8960
rect 6005 8920 6010 8950
rect 6040 8920 6045 8950
rect 6205 8950 6245 8960
rect 6205 8920 6210 8950
rect 6240 8920 6245 8950
rect 6405 8950 6445 8960
rect 6405 8920 6410 8950
rect 6440 8920 6445 8950
rect -188 8835 -185 8920
rect -165 8835 -162 8920
rect 15 8835 35 8920
rect 215 8835 235 8920
rect 415 8835 435 8920
rect 615 8835 635 8920
rect 815 8835 835 8920
rect 1015 8835 1035 8920
rect 1215 8835 1235 8920
rect 1415 8835 1435 8920
rect 1615 8835 1635 8920
rect 1815 8835 1835 8920
rect 2015 8835 2035 8920
rect 2215 8835 2235 8920
rect 2415 8835 2435 8920
rect 2615 8835 2635 8920
rect 2815 8835 2835 8920
rect 3015 8835 3035 8920
rect 3215 8835 3235 8920
rect 3415 8835 3435 8920
rect 3615 8835 3635 8920
rect 3815 8835 3835 8920
rect 4015 8835 4035 8920
rect 4215 8835 4235 8920
rect 4415 8835 4435 8920
rect 4615 8835 4635 8920
rect 4815 8835 4835 8920
rect 5015 8835 5035 8920
rect 5215 8835 5235 8920
rect 5415 8835 5435 8920
rect 5615 8835 5635 8920
rect 5815 8835 5835 8920
rect 6015 8835 6035 8920
rect 6215 8835 6235 8920
rect -195 8805 -190 8835
rect -160 8805 -155 8835
rect -195 8765 -185 8805
rect -165 8795 -155 8805
rect 5 8805 10 8835
rect 40 8805 45 8835
rect 5 8795 45 8805
rect 205 8805 210 8835
rect 240 8805 245 8835
rect 205 8795 245 8805
rect 405 8805 410 8835
rect 440 8805 445 8835
rect 405 8795 445 8805
rect 605 8805 610 8835
rect 640 8805 645 8835
rect 605 8795 645 8805
rect 805 8805 810 8835
rect 840 8805 845 8835
rect 805 8795 845 8805
rect 1005 8805 1010 8835
rect 1040 8805 1045 8835
rect 1005 8795 1045 8805
rect 1205 8805 1210 8835
rect 1240 8805 1245 8835
rect 1205 8795 1245 8805
rect 1405 8805 1410 8835
rect 1440 8805 1445 8835
rect 1405 8795 1445 8805
rect 1605 8805 1610 8835
rect 1640 8805 1645 8835
rect 1605 8795 1645 8805
rect 1805 8805 1810 8835
rect 1840 8805 1845 8835
rect 1805 8795 1845 8805
rect 2005 8805 2010 8835
rect 2040 8805 2045 8835
rect 2005 8795 2045 8805
rect 2205 8805 2210 8835
rect 2240 8805 2245 8835
rect 2205 8795 2245 8805
rect 2405 8805 2410 8835
rect 2440 8805 2445 8835
rect 2405 8795 2445 8805
rect 2605 8805 2610 8835
rect 2640 8805 2645 8835
rect 2605 8795 2645 8805
rect 2805 8805 2810 8835
rect 2840 8805 2845 8835
rect 2805 8795 2845 8805
rect 3005 8805 3010 8835
rect 3040 8805 3045 8835
rect 3005 8795 3045 8805
rect 3205 8805 3210 8835
rect 3240 8805 3245 8835
rect 3205 8795 3245 8805
rect 3405 8805 3410 8835
rect 3440 8805 3445 8835
rect 3405 8795 3445 8805
rect 3605 8805 3610 8835
rect 3640 8805 3645 8835
rect 3605 8795 3645 8805
rect 3805 8805 3810 8835
rect 3840 8805 3845 8835
rect 3805 8795 3845 8805
rect 4005 8805 4010 8835
rect 4040 8805 4045 8835
rect 4005 8795 4045 8805
rect 4205 8805 4210 8835
rect 4240 8805 4245 8835
rect 4205 8795 4245 8805
rect 4405 8805 4410 8835
rect 4440 8805 4445 8835
rect 4405 8795 4445 8805
rect 4605 8805 4610 8835
rect 4640 8805 4645 8835
rect 4605 8795 4645 8805
rect 4805 8805 4810 8835
rect 4840 8805 4845 8835
rect 4805 8795 4845 8805
rect 5005 8805 5010 8835
rect 5040 8805 5045 8835
rect 5005 8795 5045 8805
rect 5205 8805 5210 8835
rect 5240 8805 5245 8835
rect 5205 8795 5245 8805
rect 5405 8805 5410 8835
rect 5440 8805 5445 8835
rect 5405 8795 5445 8805
rect 5605 8805 5610 8835
rect 5640 8805 5645 8835
rect 5605 8795 5645 8805
rect 5805 8805 5810 8835
rect 5840 8805 5845 8835
rect 5805 8795 5845 8805
rect 6005 8805 6010 8835
rect 6040 8805 6045 8835
rect 6005 8795 6045 8805
rect 6205 8805 6210 8835
rect 6240 8805 6245 8835
rect 6205 8795 6245 8805
rect 6405 8805 6410 8835
rect 6440 8805 6445 8835
rect 6405 8795 6445 8805
rect -165 8775 -30 8795
rect 5 8775 1570 8795
rect 1605 8775 6570 8795
rect -165 8765 -155 8775
rect -195 8735 -190 8765
rect -160 8735 -155 8765
rect 5 8765 45 8775
rect 5 8735 10 8765
rect 40 8735 45 8765
rect 205 8765 245 8775
rect 205 8735 210 8765
rect 240 8735 245 8765
rect 405 8765 445 8775
rect 405 8735 410 8765
rect 440 8735 445 8765
rect 605 8765 645 8775
rect 605 8735 610 8765
rect 640 8735 645 8765
rect 805 8765 845 8775
rect 805 8735 810 8765
rect 840 8735 845 8765
rect 1005 8765 1045 8775
rect 1005 8735 1010 8765
rect 1040 8735 1045 8765
rect 1205 8765 1245 8775
rect 1205 8735 1210 8765
rect 1240 8735 1245 8765
rect 1405 8765 1445 8775
rect 1405 8735 1410 8765
rect 1440 8735 1445 8765
rect 1605 8765 1645 8775
rect 1605 8735 1610 8765
rect 1640 8735 1645 8765
rect 1805 8765 1845 8775
rect 1805 8735 1810 8765
rect 1840 8735 1845 8765
rect 2005 8765 2045 8775
rect 2005 8735 2010 8765
rect 2040 8735 2045 8765
rect 2205 8765 2245 8775
rect 2205 8735 2210 8765
rect 2240 8735 2245 8765
rect 2405 8765 2445 8775
rect 2405 8735 2410 8765
rect 2440 8735 2445 8765
rect 2605 8765 2645 8775
rect 2605 8735 2610 8765
rect 2640 8735 2645 8765
rect 2805 8765 2845 8775
rect 2805 8735 2810 8765
rect 2840 8735 2845 8765
rect 3005 8765 3045 8775
rect 3005 8735 3010 8765
rect 3040 8735 3045 8765
rect 3205 8765 3245 8775
rect 3205 8735 3210 8765
rect 3240 8735 3245 8765
rect 3405 8765 3445 8775
rect 3405 8735 3410 8765
rect 3440 8735 3445 8765
rect 3605 8765 3645 8775
rect 3605 8735 3610 8765
rect 3640 8735 3645 8765
rect 3805 8765 3845 8775
rect 3805 8735 3810 8765
rect 3840 8735 3845 8765
rect 4005 8765 4045 8775
rect 4005 8735 4010 8765
rect 4040 8735 4045 8765
rect 4205 8765 4245 8775
rect 4205 8735 4210 8765
rect 4240 8735 4245 8765
rect 4405 8765 4445 8775
rect 4405 8735 4410 8765
rect 4440 8735 4445 8765
rect 4605 8765 4645 8775
rect 4605 8735 4610 8765
rect 4640 8735 4645 8765
rect 4805 8765 4845 8775
rect 4805 8735 4810 8765
rect 4840 8735 4845 8765
rect 5005 8765 5045 8775
rect 5005 8735 5010 8765
rect 5040 8735 5045 8765
rect 5205 8765 5245 8775
rect 5205 8735 5210 8765
rect 5240 8735 5245 8765
rect 5405 8765 5445 8775
rect 5405 8735 5410 8765
rect 5440 8735 5445 8765
rect 5605 8765 5645 8775
rect 5605 8735 5610 8765
rect 5640 8735 5645 8765
rect 5805 8765 5845 8775
rect 5805 8735 5810 8765
rect 5840 8735 5845 8765
rect 6005 8765 6045 8775
rect 6005 8735 6010 8765
rect 6040 8735 6045 8765
rect 6205 8765 6245 8775
rect 6205 8735 6210 8765
rect 6240 8735 6245 8765
rect 6405 8765 6445 8775
rect 6405 8735 6410 8765
rect 6440 8735 6445 8765
rect -188 8650 -185 8735
rect -165 8650 -162 8735
rect 15 8650 35 8735
rect 215 8650 235 8735
rect 415 8650 435 8735
rect 615 8650 635 8735
rect 815 8650 835 8735
rect 1015 8650 1035 8735
rect 1215 8650 1235 8735
rect 1415 8650 1435 8735
rect 1615 8650 1635 8735
rect 1815 8650 1835 8735
rect 2015 8650 2035 8735
rect 2215 8650 2235 8735
rect 2415 8650 2435 8735
rect 2615 8650 2635 8735
rect 2815 8650 2835 8735
rect -195 8620 -190 8650
rect -160 8620 -155 8650
rect -195 8580 -185 8620
rect -165 8610 -155 8620
rect 5 8620 10 8650
rect 40 8620 45 8650
rect 5 8610 45 8620
rect 205 8620 210 8650
rect 240 8620 245 8650
rect 205 8610 245 8620
rect 405 8620 410 8650
rect 440 8620 445 8650
rect 405 8610 445 8620
rect 605 8620 610 8650
rect 640 8620 645 8650
rect 605 8610 645 8620
rect 805 8620 810 8650
rect 840 8620 845 8650
rect 805 8610 845 8620
rect 1005 8620 1010 8650
rect 1040 8620 1045 8650
rect 1005 8610 1045 8620
rect 1205 8620 1210 8650
rect 1240 8620 1245 8650
rect 1205 8610 1245 8620
rect 1405 8620 1410 8650
rect 1440 8620 1445 8650
rect 1405 8610 1445 8620
rect 1605 8620 1610 8650
rect 1640 8620 1645 8650
rect 1605 8610 1645 8620
rect 1805 8620 1810 8650
rect 1840 8620 1845 8650
rect 1805 8610 1845 8620
rect 2005 8620 2010 8650
rect 2040 8620 2045 8650
rect 2005 8610 2045 8620
rect 2205 8620 2210 8650
rect 2240 8620 2245 8650
rect 2205 8610 2245 8620
rect 2405 8620 2410 8650
rect 2440 8620 2445 8650
rect 2405 8610 2445 8620
rect 2605 8620 2610 8650
rect 2640 8620 2645 8650
rect 2605 8610 2645 8620
rect 2805 8620 2810 8650
rect 2840 8620 2845 8650
rect 2805 8610 2845 8620
rect 3005 8620 3010 8650
rect 3040 8620 3045 8650
rect 3005 8610 3045 8620
rect 3205 8620 3210 8650
rect 3240 8620 3245 8650
rect 3205 8610 3245 8620
rect 3405 8620 3410 8650
rect 3440 8620 3445 8650
rect 3405 8610 3445 8620
rect 3605 8620 3610 8650
rect 3640 8620 3645 8650
rect 3605 8610 3645 8620
rect 3805 8620 3810 8650
rect 3840 8620 3845 8650
rect 3805 8610 3845 8620
rect 4005 8620 4010 8650
rect 4040 8620 4045 8650
rect 4005 8610 4045 8620
rect 4205 8620 4210 8650
rect 4240 8620 4245 8650
rect 4205 8610 4245 8620
rect 4405 8620 4410 8650
rect 4440 8620 4445 8650
rect 4405 8610 4445 8620
rect 4605 8620 4610 8650
rect 4640 8620 4645 8650
rect 4605 8610 4645 8620
rect 4805 8620 4810 8650
rect 4840 8620 4845 8650
rect 4805 8610 4845 8620
rect 5005 8620 5010 8650
rect 5040 8620 5045 8650
rect 5005 8610 5045 8620
rect 5205 8620 5210 8650
rect 5240 8620 5245 8650
rect 5205 8610 5245 8620
rect 5405 8620 5410 8650
rect 5440 8620 5445 8650
rect 5405 8610 5445 8620
rect 5605 8620 5610 8650
rect 5640 8620 5645 8650
rect 5605 8610 5645 8620
rect 5805 8620 5810 8650
rect 5840 8620 5845 8650
rect 5805 8610 5845 8620
rect 6005 8620 6010 8650
rect 6040 8620 6045 8650
rect 6005 8610 6045 8620
rect 6205 8620 6210 8650
rect 6240 8620 6245 8650
rect 6205 8610 6245 8620
rect 6405 8620 6410 8650
rect 6440 8620 6445 8650
rect 6405 8610 6445 8620
rect -165 8590 -30 8610
rect 5 8590 1570 8610
rect 1605 8590 2970 8610
rect 3005 8590 6570 8610
rect -165 8580 -155 8590
rect -195 8550 -190 8580
rect -160 8550 -155 8580
rect 5 8580 45 8590
rect 5 8550 10 8580
rect 40 8550 45 8580
rect 205 8580 245 8590
rect 205 8550 210 8580
rect 240 8550 245 8580
rect 405 8580 445 8590
rect 405 8550 410 8580
rect 440 8550 445 8580
rect 605 8580 645 8590
rect 605 8550 610 8580
rect 640 8550 645 8580
rect 805 8580 845 8590
rect 805 8550 810 8580
rect 840 8550 845 8580
rect 1005 8580 1045 8590
rect 1005 8550 1010 8580
rect 1040 8550 1045 8580
rect 1205 8580 1245 8590
rect 1205 8550 1210 8580
rect 1240 8550 1245 8580
rect 1405 8580 1445 8590
rect 1405 8550 1410 8580
rect 1440 8550 1445 8580
rect 1605 8580 1645 8590
rect 1605 8550 1610 8580
rect 1640 8550 1645 8580
rect 1805 8580 1845 8590
rect 1805 8550 1810 8580
rect 1840 8550 1845 8580
rect 2005 8580 2045 8590
rect 2005 8550 2010 8580
rect 2040 8550 2045 8580
rect 2205 8580 2245 8590
rect 2205 8550 2210 8580
rect 2240 8550 2245 8580
rect 2405 8580 2445 8590
rect 2405 8550 2410 8580
rect 2440 8550 2445 8580
rect 2605 8580 2645 8590
rect 2605 8550 2610 8580
rect 2640 8550 2645 8580
rect 2805 8580 2845 8590
rect 2805 8550 2810 8580
rect 2840 8550 2845 8580
rect 3005 8580 3045 8590
rect 3005 8550 3010 8580
rect 3040 8550 3045 8580
rect 3205 8580 3245 8590
rect 3205 8550 3210 8580
rect 3240 8550 3245 8580
rect 3405 8580 3445 8590
rect 3405 8550 3410 8580
rect 3440 8550 3445 8580
rect 3605 8580 3645 8590
rect 3605 8550 3610 8580
rect 3640 8550 3645 8580
rect 3805 8580 3845 8590
rect 3805 8550 3810 8580
rect 3840 8550 3845 8580
rect 4005 8580 4045 8590
rect 4005 8550 4010 8580
rect 4040 8550 4045 8580
rect 4205 8580 4245 8590
rect 4205 8550 4210 8580
rect 4240 8550 4245 8580
rect 4405 8580 4445 8590
rect 4405 8550 4410 8580
rect 4440 8550 4445 8580
rect 4605 8580 4645 8590
rect 4605 8550 4610 8580
rect 4640 8550 4645 8580
rect 4805 8580 4845 8590
rect 4805 8550 4810 8580
rect 4840 8550 4845 8580
rect 5005 8580 5045 8590
rect 5005 8550 5010 8580
rect 5040 8550 5045 8580
rect 5205 8580 5245 8590
rect 5205 8550 5210 8580
rect 5240 8550 5245 8580
rect 5405 8580 5445 8590
rect 5405 8550 5410 8580
rect 5440 8550 5445 8580
rect 5605 8580 5645 8590
rect 5605 8550 5610 8580
rect 5640 8550 5645 8580
rect 5805 8580 5845 8590
rect 5805 8550 5810 8580
rect 5840 8550 5845 8580
rect 6005 8580 6045 8590
rect 6005 8550 6010 8580
rect 6040 8550 6045 8580
rect 6205 8580 6245 8590
rect 6205 8550 6210 8580
rect 6240 8550 6245 8580
rect 6405 8580 6445 8590
rect 6405 8550 6410 8580
rect 6440 8550 6445 8580
rect -188 8465 -185 8550
rect -165 8465 -162 8550
rect 15 8465 35 8550
rect 215 8465 235 8550
rect 415 8465 435 8550
rect 615 8465 635 8550
rect 815 8465 835 8550
rect 1015 8465 1035 8550
rect 1215 8465 1235 8550
rect 1415 8465 1435 8550
rect 1615 8465 1635 8550
rect 1815 8465 1835 8550
rect 2015 8465 2035 8550
rect 2215 8465 2235 8550
rect 2415 8465 2435 8550
rect 2615 8465 2635 8550
rect 2815 8465 2835 8550
rect 3015 8465 3035 8550
rect 3215 8465 3235 8550
rect 3415 8465 3435 8550
rect 3615 8465 3635 8550
rect 3815 8465 3835 8550
rect 4015 8465 4035 8550
rect 4215 8465 4235 8550
rect 4415 8465 4435 8550
rect 4615 8465 4635 8550
rect 4815 8465 4835 8550
rect 5015 8465 5035 8550
rect 5215 8465 5235 8550
rect 5415 8465 5435 8550
rect 5615 8465 5635 8550
rect 5815 8465 5835 8550
rect 6015 8465 6035 8550
rect 6215 8465 6235 8550
rect -195 8435 -190 8465
rect -160 8435 -155 8465
rect -195 8395 -185 8435
rect -165 8425 -155 8435
rect 5 8435 10 8465
rect 40 8435 45 8465
rect 5 8425 45 8435
rect 205 8435 210 8465
rect 240 8435 245 8465
rect 205 8425 245 8435
rect 405 8435 410 8465
rect 440 8435 445 8465
rect 405 8425 445 8435
rect 605 8435 610 8465
rect 640 8435 645 8465
rect 605 8425 645 8435
rect 805 8435 810 8465
rect 840 8435 845 8465
rect 805 8425 845 8435
rect 1005 8435 1010 8465
rect 1040 8435 1045 8465
rect 1005 8425 1045 8435
rect 1205 8435 1210 8465
rect 1240 8435 1245 8465
rect 1205 8425 1245 8435
rect 1405 8435 1410 8465
rect 1440 8435 1445 8465
rect 1405 8425 1445 8435
rect 1605 8435 1610 8465
rect 1640 8435 1645 8465
rect 1605 8425 1645 8435
rect 1805 8435 1810 8465
rect 1840 8435 1845 8465
rect 1805 8425 1845 8435
rect 2005 8435 2010 8465
rect 2040 8435 2045 8465
rect 2005 8425 2045 8435
rect 2205 8435 2210 8465
rect 2240 8435 2245 8465
rect 2205 8425 2245 8435
rect 2405 8435 2410 8465
rect 2440 8435 2445 8465
rect 2405 8425 2445 8435
rect 2605 8435 2610 8465
rect 2640 8435 2645 8465
rect 2605 8425 2645 8435
rect 2805 8435 2810 8465
rect 2840 8435 2845 8465
rect 2805 8425 2845 8435
rect 3005 8435 3010 8465
rect 3040 8435 3045 8465
rect 3005 8425 3045 8435
rect 3205 8435 3210 8465
rect 3240 8435 3245 8465
rect 3205 8425 3245 8435
rect 3405 8435 3410 8465
rect 3440 8435 3445 8465
rect 3405 8425 3445 8435
rect 3605 8435 3610 8465
rect 3640 8435 3645 8465
rect 3605 8425 3645 8435
rect 3805 8435 3810 8465
rect 3840 8435 3845 8465
rect 3805 8425 3845 8435
rect 4005 8435 4010 8465
rect 4040 8435 4045 8465
rect 4005 8425 4045 8435
rect 4205 8435 4210 8465
rect 4240 8435 4245 8465
rect 4205 8425 4245 8435
rect 4405 8435 4410 8465
rect 4440 8435 4445 8465
rect 4405 8425 4445 8435
rect 4605 8435 4610 8465
rect 4640 8435 4645 8465
rect 4605 8425 4645 8435
rect 4805 8435 4810 8465
rect 4840 8435 4845 8465
rect 4805 8425 4845 8435
rect 5005 8435 5010 8465
rect 5040 8435 5045 8465
rect 5005 8425 5045 8435
rect 5205 8435 5210 8465
rect 5240 8435 5245 8465
rect 5205 8425 5245 8435
rect 5405 8435 5410 8465
rect 5440 8435 5445 8465
rect 5405 8425 5445 8435
rect 5605 8435 5610 8465
rect 5640 8435 5645 8465
rect 5605 8425 5645 8435
rect 5805 8435 5810 8465
rect 5840 8435 5845 8465
rect 5805 8425 5845 8435
rect 6005 8435 6010 8465
rect 6040 8435 6045 8465
rect 6005 8425 6045 8435
rect 6205 8435 6210 8465
rect 6240 8435 6245 8465
rect 6205 8425 6245 8435
rect 6405 8435 6410 8465
rect 6440 8435 6445 8465
rect 6405 8425 6445 8435
rect -165 8405 -30 8425
rect 5 8405 1570 8425
rect 1605 8405 2970 8425
rect 3005 8405 6570 8425
rect -165 8395 -155 8405
rect -195 8365 -190 8395
rect -160 8365 -155 8395
rect 5 8395 45 8405
rect 5 8365 10 8395
rect 40 8365 45 8395
rect 205 8395 245 8405
rect 205 8365 210 8395
rect 240 8365 245 8395
rect 405 8395 445 8405
rect 405 8365 410 8395
rect 440 8365 445 8395
rect 605 8395 645 8405
rect 605 8365 610 8395
rect 640 8365 645 8395
rect 805 8395 845 8405
rect 805 8365 810 8395
rect 840 8365 845 8395
rect 1005 8395 1045 8405
rect 1005 8365 1010 8395
rect 1040 8365 1045 8395
rect 1205 8395 1245 8405
rect 1205 8365 1210 8395
rect 1240 8365 1245 8395
rect 1405 8395 1445 8405
rect 1405 8365 1410 8395
rect 1440 8365 1445 8395
rect 1605 8395 1645 8405
rect 1605 8365 1610 8395
rect 1640 8365 1645 8395
rect 1805 8395 1845 8405
rect 1805 8365 1810 8395
rect 1840 8365 1845 8395
rect 2005 8395 2045 8405
rect 2005 8365 2010 8395
rect 2040 8365 2045 8395
rect 2205 8395 2245 8405
rect 2205 8365 2210 8395
rect 2240 8365 2245 8395
rect 2405 8395 2445 8405
rect 2405 8365 2410 8395
rect 2440 8365 2445 8395
rect 2605 8395 2645 8405
rect 2605 8365 2610 8395
rect 2640 8365 2645 8395
rect 2805 8395 2845 8405
rect 2805 8365 2810 8395
rect 2840 8365 2845 8395
rect 3005 8395 3045 8405
rect 3005 8365 3010 8395
rect 3040 8365 3045 8395
rect 3205 8395 3245 8405
rect 3205 8365 3210 8395
rect 3240 8365 3245 8395
rect 3405 8395 3445 8405
rect 3405 8365 3410 8395
rect 3440 8365 3445 8395
rect 3605 8395 3645 8405
rect 3605 8365 3610 8395
rect 3640 8365 3645 8395
rect 3805 8395 3845 8405
rect 3805 8365 3810 8395
rect 3840 8365 3845 8395
rect 4005 8395 4045 8405
rect 4005 8365 4010 8395
rect 4040 8365 4045 8395
rect 4205 8395 4245 8405
rect 4205 8365 4210 8395
rect 4240 8365 4245 8395
rect 4405 8395 4445 8405
rect 4405 8365 4410 8395
rect 4440 8365 4445 8395
rect 4605 8395 4645 8405
rect 4605 8365 4610 8395
rect 4640 8365 4645 8395
rect 4805 8395 4845 8405
rect 4805 8365 4810 8395
rect 4840 8365 4845 8395
rect 5005 8395 5045 8405
rect 5005 8365 5010 8395
rect 5040 8365 5045 8395
rect 5205 8395 5245 8405
rect 5205 8365 5210 8395
rect 5240 8365 5245 8395
rect 5405 8395 5445 8405
rect 5405 8365 5410 8395
rect 5440 8365 5445 8395
rect 5605 8395 5645 8405
rect 5605 8365 5610 8395
rect 5640 8365 5645 8395
rect 5805 8395 5845 8405
rect 5805 8365 5810 8395
rect 5840 8365 5845 8395
rect 6005 8395 6045 8405
rect 6005 8365 6010 8395
rect 6040 8365 6045 8395
rect 6205 8395 6245 8405
rect 6205 8365 6210 8395
rect 6240 8365 6245 8395
rect 6405 8395 6445 8405
rect 6405 8365 6410 8395
rect 6440 8365 6445 8395
rect -188 8280 -185 8365
rect -165 8280 -162 8365
rect 15 8280 35 8365
rect 215 8280 235 8365
rect 415 8280 435 8365
rect 615 8280 635 8365
rect 815 8280 835 8365
rect 1015 8280 1035 8365
rect 1215 8280 1235 8365
rect 1415 8280 1435 8365
rect 1615 8280 1635 8365
rect 1815 8280 1835 8365
rect 2015 8280 2035 8365
rect 2215 8280 2235 8365
rect 2415 8280 2435 8365
rect 2615 8280 2635 8365
rect 2815 8280 2835 8365
rect 3015 8280 3035 8365
rect 3215 8280 3235 8365
rect 3415 8280 3435 8365
rect 3615 8280 3635 8365
rect 3815 8280 3835 8365
rect 4015 8280 4035 8365
rect 4215 8280 4235 8365
rect 4415 8280 4435 8365
rect 4615 8280 4635 8365
rect 4815 8280 4835 8365
rect 5015 8280 5035 8365
rect 5215 8280 5235 8365
rect 5415 8280 5435 8365
rect 5615 8280 5635 8365
rect 5815 8280 5835 8365
rect 6015 8280 6035 8365
rect 6215 8280 6235 8365
rect -195 8250 -190 8280
rect -160 8250 -155 8280
rect -195 8210 -185 8250
rect -165 8240 -155 8250
rect 5 8250 10 8280
rect 40 8250 45 8280
rect 5 8240 45 8250
rect 205 8250 210 8280
rect 240 8250 245 8280
rect 205 8240 245 8250
rect 405 8250 410 8280
rect 440 8250 445 8280
rect 405 8240 445 8250
rect 605 8250 610 8280
rect 640 8250 645 8280
rect 605 8240 645 8250
rect 805 8250 810 8280
rect 840 8250 845 8280
rect 805 8240 845 8250
rect 1005 8250 1010 8280
rect 1040 8250 1045 8280
rect 1005 8240 1045 8250
rect 1205 8250 1210 8280
rect 1240 8250 1245 8280
rect 1205 8240 1245 8250
rect 1405 8250 1410 8280
rect 1440 8250 1445 8280
rect 1405 8240 1445 8250
rect 1605 8250 1610 8280
rect 1640 8250 1645 8280
rect 1605 8240 1645 8250
rect 1805 8250 1810 8280
rect 1840 8250 1845 8280
rect 1805 8240 1845 8250
rect 2005 8250 2010 8280
rect 2040 8250 2045 8280
rect 2005 8240 2045 8250
rect 2205 8250 2210 8280
rect 2240 8250 2245 8280
rect 2205 8240 2245 8250
rect 2405 8250 2410 8280
rect 2440 8250 2445 8280
rect 2405 8240 2445 8250
rect 2605 8250 2610 8280
rect 2640 8250 2645 8280
rect 2605 8240 2645 8250
rect 2805 8250 2810 8280
rect 2840 8250 2845 8280
rect 2805 8240 2845 8250
rect 3005 8250 3010 8280
rect 3040 8250 3045 8280
rect 3005 8240 3045 8250
rect 3205 8250 3210 8280
rect 3240 8250 3245 8280
rect 3205 8240 3245 8250
rect 3405 8250 3410 8280
rect 3440 8250 3445 8280
rect 3405 8240 3445 8250
rect 3605 8250 3610 8280
rect 3640 8250 3645 8280
rect 3605 8240 3645 8250
rect 3805 8250 3810 8280
rect 3840 8250 3845 8280
rect 3805 8240 3845 8250
rect 4005 8250 4010 8280
rect 4040 8250 4045 8280
rect 4005 8240 4045 8250
rect 4205 8250 4210 8280
rect 4240 8250 4245 8280
rect 4205 8240 4245 8250
rect 4405 8250 4410 8280
rect 4440 8250 4445 8280
rect 4405 8240 4445 8250
rect 4605 8250 4610 8280
rect 4640 8250 4645 8280
rect 4605 8240 4645 8250
rect 4805 8250 4810 8280
rect 4840 8250 4845 8280
rect 4805 8240 4845 8250
rect 5005 8250 5010 8280
rect 5040 8250 5045 8280
rect 5005 8240 5045 8250
rect 5205 8250 5210 8280
rect 5240 8250 5245 8280
rect 5205 8240 5245 8250
rect 5405 8250 5410 8280
rect 5440 8250 5445 8280
rect 5405 8240 5445 8250
rect 5605 8250 5610 8280
rect 5640 8250 5645 8280
rect 5605 8240 5645 8250
rect 5805 8250 5810 8280
rect 5840 8250 5845 8280
rect 5805 8240 5845 8250
rect 6005 8250 6010 8280
rect 6040 8250 6045 8280
rect 6005 8240 6045 8250
rect 6205 8250 6210 8280
rect 6240 8250 6245 8280
rect 6205 8240 6245 8250
rect 6405 8250 6410 8280
rect 6440 8250 6445 8280
rect 6405 8240 6445 8250
rect -165 8220 -30 8240
rect 5 8220 1570 8240
rect 1605 8220 2970 8240
rect 3005 8220 6570 8240
rect -165 8210 -155 8220
rect -195 8180 -190 8210
rect -160 8180 -155 8210
rect 5 8210 45 8220
rect 5 8180 10 8210
rect 40 8180 45 8210
rect 205 8210 245 8220
rect 205 8180 210 8210
rect 240 8180 245 8210
rect 405 8210 445 8220
rect 405 8180 410 8210
rect 440 8180 445 8210
rect 605 8210 645 8220
rect 605 8180 610 8210
rect 640 8180 645 8210
rect 805 8210 845 8220
rect 805 8180 810 8210
rect 840 8180 845 8210
rect 1005 8210 1045 8220
rect 1005 8180 1010 8210
rect 1040 8180 1045 8210
rect 1205 8210 1245 8220
rect 1205 8180 1210 8210
rect 1240 8180 1245 8210
rect 1405 8210 1445 8220
rect 1405 8180 1410 8210
rect 1440 8180 1445 8210
rect 1605 8210 1645 8220
rect 1605 8180 1610 8210
rect 1640 8180 1645 8210
rect 1805 8210 1845 8220
rect 1805 8180 1810 8210
rect 1840 8180 1845 8210
rect 2005 8210 2045 8220
rect 2005 8180 2010 8210
rect 2040 8180 2045 8210
rect 2205 8210 2245 8220
rect 2205 8180 2210 8210
rect 2240 8180 2245 8210
rect 2405 8210 2445 8220
rect 2405 8180 2410 8210
rect 2440 8180 2445 8210
rect 2605 8210 2645 8220
rect 2605 8180 2610 8210
rect 2640 8180 2645 8210
rect 2805 8210 2845 8220
rect 2805 8180 2810 8210
rect 2840 8180 2845 8210
rect 3005 8210 3045 8220
rect 3005 8180 3010 8210
rect 3040 8180 3045 8210
rect 3205 8210 3245 8220
rect 3205 8180 3210 8210
rect 3240 8180 3245 8210
rect 3405 8210 3445 8220
rect 3405 8180 3410 8210
rect 3440 8180 3445 8210
rect 3605 8210 3645 8220
rect 3605 8180 3610 8210
rect 3640 8180 3645 8210
rect 3805 8210 3845 8220
rect 3805 8180 3810 8210
rect 3840 8180 3845 8210
rect 4005 8210 4045 8220
rect 4005 8180 4010 8210
rect 4040 8180 4045 8210
rect 4205 8210 4245 8220
rect 4205 8180 4210 8210
rect 4240 8180 4245 8210
rect 4405 8210 4445 8220
rect 4405 8180 4410 8210
rect 4440 8180 4445 8210
rect 4605 8210 4645 8220
rect 4605 8180 4610 8210
rect 4640 8180 4645 8210
rect 4805 8210 4845 8220
rect 4805 8180 4810 8210
rect 4840 8180 4845 8210
rect 5005 8210 5045 8220
rect 5005 8180 5010 8210
rect 5040 8180 5045 8210
rect 5205 8210 5245 8220
rect 5205 8180 5210 8210
rect 5240 8180 5245 8210
rect 5405 8210 5445 8220
rect 5405 8180 5410 8210
rect 5440 8180 5445 8210
rect 5605 8210 5645 8220
rect 5605 8180 5610 8210
rect 5640 8180 5645 8210
rect 5805 8210 5845 8220
rect 5805 8180 5810 8210
rect 5840 8180 5845 8210
rect 6005 8210 6045 8220
rect 6005 8180 6010 8210
rect 6040 8180 6045 8210
rect 6205 8210 6245 8220
rect 6205 8180 6210 8210
rect 6240 8180 6245 8210
rect 6405 8210 6445 8220
rect 6405 8180 6410 8210
rect 6440 8180 6445 8210
rect -188 8095 -185 8180
rect -165 8095 -162 8180
rect 15 8095 35 8180
rect 215 8095 235 8180
rect 415 8095 435 8180
rect 615 8095 635 8180
rect 815 8095 835 8180
rect 1015 8095 1035 8180
rect 1215 8095 1235 8180
rect 1415 8095 1435 8180
rect 1615 8095 1635 8180
rect 1815 8095 1835 8180
rect 2015 8095 2035 8180
rect 2215 8095 2235 8180
rect 2415 8095 2435 8180
rect 2615 8095 2635 8180
rect 2815 8095 2835 8180
rect 3015 8095 3035 8180
rect 3215 8095 3235 8180
rect 3415 8095 3435 8180
rect 3615 8095 3635 8180
rect 3815 8095 3835 8180
rect 4015 8095 4035 8180
rect 4215 8095 4235 8180
rect 4415 8095 4435 8180
rect 4615 8095 4635 8180
rect 4815 8095 4835 8180
rect 5015 8095 5035 8180
rect 5215 8095 5235 8180
rect 5415 8095 5435 8180
rect 5615 8095 5635 8180
rect 5815 8095 5835 8180
rect 6015 8095 6035 8180
rect 6215 8095 6235 8180
rect -195 8065 -190 8095
rect -160 8065 -155 8095
rect -195 8025 -185 8065
rect -165 8055 -155 8065
rect 5 8065 10 8095
rect 40 8065 45 8095
rect 5 8055 45 8065
rect 205 8065 210 8095
rect 240 8065 245 8095
rect 205 8055 245 8065
rect 405 8065 410 8095
rect 440 8065 445 8095
rect 405 8055 445 8065
rect 605 8065 610 8095
rect 640 8065 645 8095
rect 605 8055 645 8065
rect 805 8065 810 8095
rect 840 8065 845 8095
rect 805 8055 845 8065
rect 1005 8065 1010 8095
rect 1040 8065 1045 8095
rect 1005 8055 1045 8065
rect 1205 8065 1210 8095
rect 1240 8065 1245 8095
rect 1205 8055 1245 8065
rect 1405 8065 1410 8095
rect 1440 8065 1445 8095
rect 1405 8055 1445 8065
rect 1605 8065 1610 8095
rect 1640 8065 1645 8095
rect 1605 8055 1645 8065
rect 1805 8065 1810 8095
rect 1840 8065 1845 8095
rect 1805 8055 1845 8065
rect 2005 8065 2010 8095
rect 2040 8065 2045 8095
rect 2005 8055 2045 8065
rect 2205 8065 2210 8095
rect 2240 8065 2245 8095
rect 2205 8055 2245 8065
rect 2405 8065 2410 8095
rect 2440 8065 2445 8095
rect 2405 8055 2445 8065
rect 2605 8065 2610 8095
rect 2640 8065 2645 8095
rect 2605 8055 2645 8065
rect 2805 8065 2810 8095
rect 2840 8065 2845 8095
rect 2805 8055 2845 8065
rect 3005 8065 3010 8095
rect 3040 8065 3045 8095
rect 3005 8055 3045 8065
rect 3205 8065 3210 8095
rect 3240 8065 3245 8095
rect 3205 8055 3245 8065
rect 3405 8065 3410 8095
rect 3440 8065 3445 8095
rect 3405 8055 3445 8065
rect 3605 8065 3610 8095
rect 3640 8065 3645 8095
rect 3605 8055 3645 8065
rect 3805 8065 3810 8095
rect 3840 8065 3845 8095
rect 3805 8055 3845 8065
rect 4005 8065 4010 8095
rect 4040 8065 4045 8095
rect 4005 8055 4045 8065
rect 4205 8065 4210 8095
rect 4240 8065 4245 8095
rect 4205 8055 4245 8065
rect 4405 8065 4410 8095
rect 4440 8065 4445 8095
rect 4405 8055 4445 8065
rect 4605 8065 4610 8095
rect 4640 8065 4645 8095
rect 4605 8055 4645 8065
rect 4805 8065 4810 8095
rect 4840 8065 4845 8095
rect 4805 8055 4845 8065
rect 5005 8065 5010 8095
rect 5040 8065 5045 8095
rect 5005 8055 5045 8065
rect 5205 8065 5210 8095
rect 5240 8065 5245 8095
rect 5205 8055 5245 8065
rect 5405 8065 5410 8095
rect 5440 8065 5445 8095
rect 5405 8055 5445 8065
rect 5605 8065 5610 8095
rect 5640 8065 5645 8095
rect 5605 8055 5645 8065
rect 5805 8065 5810 8095
rect 5840 8065 5845 8095
rect 5805 8055 5845 8065
rect 6005 8065 6010 8095
rect 6040 8065 6045 8095
rect 6005 8055 6045 8065
rect 6205 8065 6210 8095
rect 6240 8065 6245 8095
rect 6205 8055 6245 8065
rect 6405 8065 6410 8095
rect 6440 8065 6445 8095
rect 6405 8055 6445 8065
rect -165 8035 -30 8055
rect 5 8035 1570 8055
rect 1605 8035 2970 8055
rect 3005 8035 6570 8055
rect -165 8025 -155 8035
rect -195 7995 -190 8025
rect -160 7995 -155 8025
rect 5 8025 45 8035
rect 5 7995 10 8025
rect 40 7995 45 8025
rect 205 8025 245 8035
rect 205 7995 210 8025
rect 240 7995 245 8025
rect 405 8025 445 8035
rect 405 7995 410 8025
rect 440 7995 445 8025
rect 605 8025 645 8035
rect 605 7995 610 8025
rect 640 7995 645 8025
rect 805 8025 845 8035
rect 805 7995 810 8025
rect 840 7995 845 8025
rect 1005 8025 1045 8035
rect 1005 7995 1010 8025
rect 1040 7995 1045 8025
rect 1205 8025 1245 8035
rect 1205 7995 1210 8025
rect 1240 7995 1245 8025
rect 1405 8025 1445 8035
rect 1405 7995 1410 8025
rect 1440 7995 1445 8025
rect 1605 8025 1645 8035
rect 1605 7995 1610 8025
rect 1640 7995 1645 8025
rect 1805 8025 1845 8035
rect 1805 7995 1810 8025
rect 1840 7995 1845 8025
rect 2005 8025 2045 8035
rect 2005 7995 2010 8025
rect 2040 7995 2045 8025
rect 2205 8025 2245 8035
rect 2205 7995 2210 8025
rect 2240 7995 2245 8025
rect 2405 8025 2445 8035
rect 2405 7995 2410 8025
rect 2440 7995 2445 8025
rect 2605 8025 2645 8035
rect 2605 7995 2610 8025
rect 2640 7995 2645 8025
rect 2805 8025 2845 8035
rect 2805 7995 2810 8025
rect 2840 7995 2845 8025
rect 3005 8025 3045 8035
rect 3005 7995 3010 8025
rect 3040 7995 3045 8025
rect 3205 8025 3245 8035
rect 3205 7995 3210 8025
rect 3240 7995 3245 8025
rect 3405 8025 3445 8035
rect 3405 7995 3410 8025
rect 3440 7995 3445 8025
rect 3605 8025 3645 8035
rect 3605 7995 3610 8025
rect 3640 7995 3645 8025
rect 3805 8025 3845 8035
rect 3805 7995 3810 8025
rect 3840 7995 3845 8025
rect 4005 8025 4045 8035
rect 4005 7995 4010 8025
rect 4040 7995 4045 8025
rect 4205 8025 4245 8035
rect 4205 7995 4210 8025
rect 4240 7995 4245 8025
rect 4405 8025 4445 8035
rect 4405 7995 4410 8025
rect 4440 7995 4445 8025
rect 4605 8025 4645 8035
rect 4605 7995 4610 8025
rect 4640 7995 4645 8025
rect 4805 8025 4845 8035
rect 4805 7995 4810 8025
rect 4840 7995 4845 8025
rect 5005 8025 5045 8035
rect 5005 7995 5010 8025
rect 5040 7995 5045 8025
rect 5205 8025 5245 8035
rect 5205 7995 5210 8025
rect 5240 7995 5245 8025
rect 5405 8025 5445 8035
rect 5405 7995 5410 8025
rect 5440 7995 5445 8025
rect 5605 8025 5645 8035
rect 5605 7995 5610 8025
rect 5640 7995 5645 8025
rect 5805 8025 5845 8035
rect 5805 7995 5810 8025
rect 5840 7995 5845 8025
rect 6005 8025 6045 8035
rect 6005 7995 6010 8025
rect 6040 7995 6045 8025
rect 6205 8025 6245 8035
rect 6205 7995 6210 8025
rect 6240 7995 6245 8025
rect 6405 8025 6445 8035
rect 6405 7995 6410 8025
rect 6440 7995 6445 8025
rect -188 7910 -185 7995
rect -165 7910 -162 7995
rect 15 7910 35 7995
rect 215 7910 235 7995
rect 415 7910 435 7995
rect 615 7910 635 7995
rect 815 7910 835 7995
rect 1015 7910 1035 7995
rect 1215 7910 1235 7995
rect 1415 7910 1435 7995
rect 1615 7910 1635 7995
rect 1815 7910 1835 7995
rect 2015 7910 2035 7995
rect 2215 7910 2235 7995
rect 2415 7910 2435 7995
rect 2615 7910 2635 7995
rect 2815 7910 2835 7995
rect 3015 7910 3035 7995
rect 3215 7910 3235 7995
rect 3415 7910 3435 7995
rect 3615 7910 3635 7995
rect 3815 7910 3835 7995
rect 4015 7910 4035 7995
rect 4215 7910 4235 7995
rect 4415 7910 4435 7995
rect 4615 7910 4635 7995
rect 4815 7910 4835 7995
rect 5015 7910 5035 7995
rect 5215 7910 5235 7995
rect 5415 7910 5435 7995
rect 5615 7910 5635 7995
rect 5815 7910 5835 7995
rect 6015 7910 6035 7995
rect 6215 7910 6235 7995
rect -195 7880 -190 7910
rect -160 7880 -155 7910
rect -195 7840 -185 7880
rect -165 7870 -155 7880
rect 5 7880 10 7910
rect 40 7880 45 7910
rect 5 7870 45 7880
rect 205 7880 210 7910
rect 240 7880 245 7910
rect 205 7870 245 7880
rect 405 7880 410 7910
rect 440 7880 445 7910
rect 405 7870 445 7880
rect 605 7880 610 7910
rect 640 7880 645 7910
rect 605 7870 645 7880
rect 805 7880 810 7910
rect 840 7880 845 7910
rect 805 7870 845 7880
rect 1005 7880 1010 7910
rect 1040 7880 1045 7910
rect 1005 7870 1045 7880
rect 1205 7880 1210 7910
rect 1240 7880 1245 7910
rect 1205 7870 1245 7880
rect 1405 7880 1410 7910
rect 1440 7880 1445 7910
rect 1405 7870 1445 7880
rect 1605 7880 1610 7910
rect 1640 7880 1645 7910
rect 1605 7870 1645 7880
rect 1805 7880 1810 7910
rect 1840 7880 1845 7910
rect 1805 7870 1845 7880
rect 2005 7880 2010 7910
rect 2040 7880 2045 7910
rect 2005 7870 2045 7880
rect 2205 7880 2210 7910
rect 2240 7880 2245 7910
rect 2205 7870 2245 7880
rect 2405 7880 2410 7910
rect 2440 7880 2445 7910
rect 2405 7870 2445 7880
rect 2605 7880 2610 7910
rect 2640 7880 2645 7910
rect 2605 7870 2645 7880
rect 2805 7880 2810 7910
rect 2840 7880 2845 7910
rect 2805 7870 2845 7880
rect 3005 7880 3010 7910
rect 3040 7880 3045 7910
rect 3005 7870 3045 7880
rect 3205 7880 3210 7910
rect 3240 7880 3245 7910
rect 3205 7870 3245 7880
rect 3405 7880 3410 7910
rect 3440 7880 3445 7910
rect 3405 7870 3445 7880
rect 3605 7880 3610 7910
rect 3640 7880 3645 7910
rect 3605 7870 3645 7880
rect 3805 7880 3810 7910
rect 3840 7880 3845 7910
rect 3805 7870 3845 7880
rect 4005 7880 4010 7910
rect 4040 7880 4045 7910
rect 4005 7870 4045 7880
rect 4205 7880 4210 7910
rect 4240 7880 4245 7910
rect 4205 7870 4245 7880
rect 4405 7880 4410 7910
rect 4440 7880 4445 7910
rect 4405 7870 4445 7880
rect 4605 7880 4610 7910
rect 4640 7880 4645 7910
rect 4605 7870 4645 7880
rect 4805 7880 4810 7910
rect 4840 7880 4845 7910
rect 4805 7870 4845 7880
rect 5005 7880 5010 7910
rect 5040 7880 5045 7910
rect 5005 7870 5045 7880
rect 5205 7880 5210 7910
rect 5240 7880 5245 7910
rect 5205 7870 5245 7880
rect 5405 7880 5410 7910
rect 5440 7880 5445 7910
rect 5405 7870 5445 7880
rect 5605 7880 5610 7910
rect 5640 7880 5645 7910
rect 5605 7870 5645 7880
rect 5805 7880 5810 7910
rect 5840 7880 5845 7910
rect 5805 7870 5845 7880
rect 6005 7880 6010 7910
rect 6040 7880 6045 7910
rect 6005 7870 6045 7880
rect 6205 7880 6210 7910
rect 6240 7880 6245 7910
rect 6205 7870 6245 7880
rect 6405 7880 6410 7910
rect 6440 7880 6445 7910
rect 6405 7870 6445 7880
rect -165 7850 -30 7870
rect 5 7850 1570 7870
rect 1605 7850 2970 7870
rect 3005 7850 6570 7870
rect -165 7840 -155 7850
rect -195 7810 -190 7840
rect -160 7810 -155 7840
rect 5 7840 45 7850
rect 5 7810 10 7840
rect 40 7810 45 7840
rect 205 7840 245 7850
rect 205 7810 210 7840
rect 240 7810 245 7840
rect 405 7840 445 7850
rect 405 7810 410 7840
rect 440 7810 445 7840
rect 605 7840 645 7850
rect 605 7810 610 7840
rect 640 7810 645 7840
rect 805 7840 845 7850
rect 805 7810 810 7840
rect 840 7810 845 7840
rect 1005 7840 1045 7850
rect 1005 7810 1010 7840
rect 1040 7810 1045 7840
rect 1205 7840 1245 7850
rect 1205 7810 1210 7840
rect 1240 7810 1245 7840
rect 1405 7840 1445 7850
rect 1405 7810 1410 7840
rect 1440 7810 1445 7840
rect 1605 7840 1645 7850
rect 1605 7810 1610 7840
rect 1640 7810 1645 7840
rect 1805 7840 1845 7850
rect 1805 7810 1810 7840
rect 1840 7810 1845 7840
rect 2005 7840 2045 7850
rect 2005 7810 2010 7840
rect 2040 7810 2045 7840
rect 2205 7840 2245 7850
rect 2205 7810 2210 7840
rect 2240 7810 2245 7840
rect 2405 7840 2445 7850
rect 2405 7810 2410 7840
rect 2440 7810 2445 7840
rect 2605 7840 2645 7850
rect 2605 7810 2610 7840
rect 2640 7810 2645 7840
rect 2805 7840 2845 7850
rect 2805 7810 2810 7840
rect 2840 7810 2845 7840
rect 3005 7840 3045 7850
rect 3005 7810 3010 7840
rect 3040 7810 3045 7840
rect 3205 7840 3245 7850
rect 3205 7810 3210 7840
rect 3240 7810 3245 7840
rect 3405 7840 3445 7850
rect 3405 7810 3410 7840
rect 3440 7810 3445 7840
rect 3605 7840 3645 7850
rect 3605 7810 3610 7840
rect 3640 7810 3645 7840
rect 3805 7840 3845 7850
rect 3805 7810 3810 7840
rect 3840 7810 3845 7840
rect 4005 7840 4045 7850
rect 4005 7810 4010 7840
rect 4040 7810 4045 7840
rect 4205 7840 4245 7850
rect 4205 7810 4210 7840
rect 4240 7810 4245 7840
rect 4405 7840 4445 7850
rect 4405 7810 4410 7840
rect 4440 7810 4445 7840
rect 4605 7840 4645 7850
rect 4605 7810 4610 7840
rect 4640 7810 4645 7840
rect 4805 7840 4845 7850
rect 4805 7810 4810 7840
rect 4840 7810 4845 7840
rect 5005 7840 5045 7850
rect 5005 7810 5010 7840
rect 5040 7810 5045 7840
rect 5205 7840 5245 7850
rect 5205 7810 5210 7840
rect 5240 7810 5245 7840
rect 5405 7840 5445 7850
rect 5405 7810 5410 7840
rect 5440 7810 5445 7840
rect 5605 7840 5645 7850
rect 5605 7810 5610 7840
rect 5640 7810 5645 7840
rect 5805 7840 5845 7850
rect 5805 7810 5810 7840
rect 5840 7810 5845 7840
rect 6005 7840 6045 7850
rect 6005 7810 6010 7840
rect 6040 7810 6045 7840
rect 6205 7840 6245 7850
rect 6205 7810 6210 7840
rect 6240 7810 6245 7840
rect 6405 7840 6445 7850
rect 6405 7810 6410 7840
rect 6440 7810 6445 7840
rect -188 7725 -185 7810
rect -165 7725 -162 7810
rect 15 7725 35 7810
rect 215 7725 235 7810
rect 415 7725 435 7810
rect 615 7725 635 7810
rect 815 7725 835 7810
rect 1015 7725 1035 7810
rect 1215 7725 1235 7810
rect 1415 7725 1435 7810
rect 1615 7725 1635 7810
rect 1815 7725 1835 7810
rect 2015 7725 2035 7810
rect 2215 7725 2235 7810
rect 2415 7725 2435 7810
rect 2615 7725 2635 7810
rect 2815 7725 2835 7810
rect 3015 7725 3035 7810
rect 3215 7725 3235 7810
rect 3415 7725 3435 7810
rect 3615 7725 3635 7810
rect 3815 7725 3835 7810
rect -195 7695 -190 7725
rect -160 7695 -155 7725
rect -195 7655 -185 7695
rect -165 7685 -155 7695
rect 5 7695 10 7725
rect 40 7695 45 7725
rect 5 7685 45 7695
rect 205 7695 210 7725
rect 240 7695 245 7725
rect 205 7685 245 7695
rect 405 7695 410 7725
rect 440 7695 445 7725
rect 405 7685 445 7695
rect 605 7695 610 7725
rect 640 7695 645 7725
rect 605 7685 645 7695
rect 805 7695 810 7725
rect 840 7695 845 7725
rect 805 7685 845 7695
rect 1005 7695 1010 7725
rect 1040 7695 1045 7725
rect 1005 7685 1045 7695
rect 1205 7695 1210 7725
rect 1240 7695 1245 7725
rect 1205 7685 1245 7695
rect 1405 7695 1410 7725
rect 1440 7695 1445 7725
rect 1405 7685 1445 7695
rect 1605 7695 1610 7725
rect 1640 7695 1645 7725
rect 1605 7685 1645 7695
rect 1805 7695 1810 7725
rect 1840 7695 1845 7725
rect 1805 7685 1845 7695
rect 2005 7695 2010 7725
rect 2040 7695 2045 7725
rect 2005 7685 2045 7695
rect 2205 7695 2210 7725
rect 2240 7695 2245 7725
rect 2205 7685 2245 7695
rect 2405 7695 2410 7725
rect 2440 7695 2445 7725
rect 2405 7685 2445 7695
rect 2605 7695 2610 7725
rect 2640 7695 2645 7725
rect 2605 7685 2645 7695
rect 2805 7695 2810 7725
rect 2840 7695 2845 7725
rect 2805 7685 2845 7695
rect 3005 7695 3010 7725
rect 3040 7695 3045 7725
rect 3005 7685 3045 7695
rect 3205 7695 3210 7725
rect 3240 7695 3245 7725
rect 3205 7685 3245 7695
rect 3405 7695 3410 7725
rect 3440 7695 3445 7725
rect 3405 7685 3445 7695
rect 3605 7695 3610 7725
rect 3640 7695 3645 7725
rect 3605 7685 3645 7695
rect 3805 7695 3810 7725
rect 3840 7695 3845 7725
rect 3805 7685 3845 7695
rect 4005 7695 4010 7725
rect 4040 7695 4045 7725
rect 4005 7685 4045 7695
rect 4205 7695 4210 7725
rect 4240 7695 4245 7725
rect 4205 7685 4245 7695
rect 4405 7695 4410 7725
rect 4440 7695 4445 7725
rect 4405 7685 4445 7695
rect 4605 7695 4610 7725
rect 4640 7695 4645 7725
rect 4605 7685 4645 7695
rect 4805 7695 4810 7725
rect 4840 7695 4845 7725
rect 4805 7685 4845 7695
rect 5005 7695 5010 7725
rect 5040 7695 5045 7725
rect 5005 7685 5045 7695
rect 5205 7695 5210 7725
rect 5240 7695 5245 7725
rect 5205 7685 5245 7695
rect 5405 7695 5410 7725
rect 5440 7695 5445 7725
rect 5405 7685 5445 7695
rect 5605 7695 5610 7725
rect 5640 7695 5645 7725
rect 5605 7685 5645 7695
rect 5805 7695 5810 7725
rect 5840 7695 5845 7725
rect 5805 7685 5845 7695
rect 6005 7695 6010 7725
rect 6040 7695 6045 7725
rect 6005 7685 6045 7695
rect 6205 7695 6210 7725
rect 6240 7695 6245 7725
rect 6205 7685 6245 7695
rect 6405 7695 6410 7725
rect 6440 7695 6445 7725
rect 6405 7685 6445 7695
rect -165 7665 -30 7685
rect 5 7665 1570 7685
rect 1605 7665 2970 7685
rect 3005 7665 3970 7685
rect 4005 7665 6570 7685
rect -165 7655 -155 7665
rect -195 7625 -190 7655
rect -160 7625 -155 7655
rect 5 7655 45 7665
rect 5 7625 10 7655
rect 40 7625 45 7655
rect 205 7655 245 7665
rect 205 7625 210 7655
rect 240 7625 245 7655
rect 405 7655 445 7665
rect 405 7625 410 7655
rect 440 7625 445 7655
rect 605 7655 645 7665
rect 605 7625 610 7655
rect 640 7625 645 7655
rect 805 7655 845 7665
rect 805 7625 810 7655
rect 840 7625 845 7655
rect 1005 7655 1045 7665
rect 1005 7625 1010 7655
rect 1040 7625 1045 7655
rect 1205 7655 1245 7665
rect 1205 7625 1210 7655
rect 1240 7625 1245 7655
rect 1405 7655 1445 7665
rect 1405 7625 1410 7655
rect 1440 7625 1445 7655
rect 1605 7655 1645 7665
rect 1605 7625 1610 7655
rect 1640 7625 1645 7655
rect 1805 7655 1845 7665
rect 1805 7625 1810 7655
rect 1840 7625 1845 7655
rect 2005 7655 2045 7665
rect 2005 7625 2010 7655
rect 2040 7625 2045 7655
rect 2205 7655 2245 7665
rect 2205 7625 2210 7655
rect 2240 7625 2245 7655
rect 2405 7655 2445 7665
rect 2405 7625 2410 7655
rect 2440 7625 2445 7655
rect 2605 7655 2645 7665
rect 2605 7625 2610 7655
rect 2640 7625 2645 7655
rect 2805 7655 2845 7665
rect 2805 7625 2810 7655
rect 2840 7625 2845 7655
rect 3005 7655 3045 7665
rect 3005 7625 3010 7655
rect 3040 7625 3045 7655
rect 3205 7655 3245 7665
rect 3205 7625 3210 7655
rect 3240 7625 3245 7655
rect 3405 7655 3445 7665
rect 3405 7625 3410 7655
rect 3440 7625 3445 7655
rect 3605 7655 3645 7665
rect 3605 7625 3610 7655
rect 3640 7625 3645 7655
rect 3805 7655 3845 7665
rect 3805 7625 3810 7655
rect 3840 7625 3845 7655
rect 4005 7655 4045 7665
rect 4005 7625 4010 7655
rect 4040 7625 4045 7655
rect 4205 7655 4245 7665
rect 4205 7625 4210 7655
rect 4240 7625 4245 7655
rect 4405 7655 4445 7665
rect 4405 7625 4410 7655
rect 4440 7625 4445 7655
rect 4605 7655 4645 7665
rect 4605 7625 4610 7655
rect 4640 7625 4645 7655
rect 4805 7655 4845 7665
rect 4805 7625 4810 7655
rect 4840 7625 4845 7655
rect 5005 7655 5045 7665
rect 5005 7625 5010 7655
rect 5040 7625 5045 7655
rect 5205 7655 5245 7665
rect 5205 7625 5210 7655
rect 5240 7625 5245 7655
rect 5405 7655 5445 7665
rect 5405 7625 5410 7655
rect 5440 7625 5445 7655
rect 5605 7655 5645 7665
rect 5605 7625 5610 7655
rect 5640 7625 5645 7655
rect 5805 7655 5845 7665
rect 5805 7625 5810 7655
rect 5840 7625 5845 7655
rect 6005 7655 6045 7665
rect 6005 7625 6010 7655
rect 6040 7625 6045 7655
rect 6205 7655 6245 7665
rect 6205 7625 6210 7655
rect 6240 7625 6245 7655
rect 6405 7655 6445 7665
rect 6405 7625 6410 7655
rect 6440 7625 6445 7655
rect -188 7540 -185 7625
rect -165 7540 -162 7625
rect 15 7540 35 7625
rect 215 7540 235 7625
rect 415 7540 435 7625
rect 615 7540 635 7625
rect 815 7540 835 7625
rect 1015 7540 1035 7625
rect 1215 7540 1235 7625
rect 1415 7540 1435 7625
rect 1615 7540 1635 7625
rect 1815 7540 1835 7625
rect 2015 7540 2035 7625
rect 2215 7540 2235 7625
rect 2415 7540 2435 7625
rect 2615 7540 2635 7625
rect 2815 7540 2835 7625
rect 3015 7540 3035 7625
rect 3215 7540 3235 7625
rect 3415 7540 3435 7625
rect 3615 7540 3635 7625
rect 3815 7540 3835 7625
rect 4015 7540 4035 7625
rect 4215 7540 4235 7625
rect 4415 7540 4435 7625
rect 4615 7540 4635 7625
rect 4815 7540 4835 7625
rect 5015 7540 5035 7625
rect 5215 7540 5235 7625
rect 5415 7540 5435 7625
rect 5615 7540 5635 7625
rect 5815 7540 5835 7625
rect 6015 7540 6035 7625
rect 6215 7540 6235 7625
rect -195 7510 -190 7540
rect -160 7510 -155 7540
rect -195 7470 -185 7510
rect -165 7500 -155 7510
rect 5 7510 10 7540
rect 40 7510 45 7540
rect 5 7500 45 7510
rect 205 7510 210 7540
rect 240 7510 245 7540
rect 205 7500 245 7510
rect 405 7510 410 7540
rect 440 7510 445 7540
rect 405 7500 445 7510
rect 605 7510 610 7540
rect 640 7510 645 7540
rect 605 7500 645 7510
rect 805 7510 810 7540
rect 840 7510 845 7540
rect 805 7500 845 7510
rect 1005 7510 1010 7540
rect 1040 7510 1045 7540
rect 1005 7500 1045 7510
rect 1205 7510 1210 7540
rect 1240 7510 1245 7540
rect 1205 7500 1245 7510
rect 1405 7510 1410 7540
rect 1440 7510 1445 7540
rect 1405 7500 1445 7510
rect 1605 7510 1610 7540
rect 1640 7510 1645 7540
rect 1605 7500 1645 7510
rect 1805 7510 1810 7540
rect 1840 7510 1845 7540
rect 1805 7500 1845 7510
rect 2005 7510 2010 7540
rect 2040 7510 2045 7540
rect 2005 7500 2045 7510
rect 2205 7510 2210 7540
rect 2240 7510 2245 7540
rect 2205 7500 2245 7510
rect 2405 7510 2410 7540
rect 2440 7510 2445 7540
rect 2405 7500 2445 7510
rect 2605 7510 2610 7540
rect 2640 7510 2645 7540
rect 2605 7500 2645 7510
rect 2805 7510 2810 7540
rect 2840 7510 2845 7540
rect 2805 7500 2845 7510
rect 3005 7510 3010 7540
rect 3040 7510 3045 7540
rect 3005 7500 3045 7510
rect 3205 7510 3210 7540
rect 3240 7510 3245 7540
rect 3205 7500 3245 7510
rect 3405 7510 3410 7540
rect 3440 7510 3445 7540
rect 3405 7500 3445 7510
rect 3605 7510 3610 7540
rect 3640 7510 3645 7540
rect 3605 7500 3645 7510
rect 3805 7510 3810 7540
rect 3840 7510 3845 7540
rect 3805 7500 3845 7510
rect 4005 7510 4010 7540
rect 4040 7510 4045 7540
rect 4005 7500 4045 7510
rect 4205 7510 4210 7540
rect 4240 7510 4245 7540
rect 4205 7500 4245 7510
rect 4405 7510 4410 7540
rect 4440 7510 4445 7540
rect 4405 7500 4445 7510
rect 4605 7510 4610 7540
rect 4640 7510 4645 7540
rect 4605 7500 4645 7510
rect 4805 7510 4810 7540
rect 4840 7510 4845 7540
rect 4805 7500 4845 7510
rect 5005 7510 5010 7540
rect 5040 7510 5045 7540
rect 5005 7500 5045 7510
rect 5205 7510 5210 7540
rect 5240 7510 5245 7540
rect 5205 7500 5245 7510
rect 5405 7510 5410 7540
rect 5440 7510 5445 7540
rect 5405 7500 5445 7510
rect 5605 7510 5610 7540
rect 5640 7510 5645 7540
rect 5605 7500 5645 7510
rect 5805 7510 5810 7540
rect 5840 7510 5845 7540
rect 5805 7500 5845 7510
rect 6005 7510 6010 7540
rect 6040 7510 6045 7540
rect 6005 7500 6045 7510
rect 6205 7510 6210 7540
rect 6240 7510 6245 7540
rect 6205 7500 6245 7510
rect 6405 7510 6410 7540
rect 6440 7510 6445 7540
rect 6405 7500 6445 7510
rect -165 7480 -30 7500
rect 5 7480 1570 7500
rect 1605 7480 2970 7500
rect 3005 7480 3970 7500
rect 4005 7480 6570 7500
rect -165 7470 -155 7480
rect -195 7440 -190 7470
rect -160 7440 -155 7470
rect 5 7470 45 7480
rect 5 7440 10 7470
rect 40 7440 45 7470
rect 205 7470 245 7480
rect 205 7440 210 7470
rect 240 7440 245 7470
rect 405 7470 445 7480
rect 405 7440 410 7470
rect 440 7440 445 7470
rect 605 7470 645 7480
rect 605 7440 610 7470
rect 640 7440 645 7470
rect 805 7470 845 7480
rect 805 7440 810 7470
rect 840 7440 845 7470
rect 1005 7470 1045 7480
rect 1005 7440 1010 7470
rect 1040 7440 1045 7470
rect 1205 7470 1245 7480
rect 1205 7440 1210 7470
rect 1240 7440 1245 7470
rect 1405 7470 1445 7480
rect 1405 7440 1410 7470
rect 1440 7440 1445 7470
rect 1605 7470 1645 7480
rect 1605 7440 1610 7470
rect 1640 7440 1645 7470
rect 1805 7470 1845 7480
rect 1805 7440 1810 7470
rect 1840 7440 1845 7470
rect 2005 7470 2045 7480
rect 2005 7440 2010 7470
rect 2040 7440 2045 7470
rect 2205 7470 2245 7480
rect 2205 7440 2210 7470
rect 2240 7440 2245 7470
rect 2405 7470 2445 7480
rect 2405 7440 2410 7470
rect 2440 7440 2445 7470
rect 2605 7470 2645 7480
rect 2605 7440 2610 7470
rect 2640 7440 2645 7470
rect 2805 7470 2845 7480
rect 2805 7440 2810 7470
rect 2840 7440 2845 7470
rect 3005 7470 3045 7480
rect 3005 7440 3010 7470
rect 3040 7440 3045 7470
rect 3205 7470 3245 7480
rect 3205 7440 3210 7470
rect 3240 7440 3245 7470
rect 3405 7470 3445 7480
rect 3405 7440 3410 7470
rect 3440 7440 3445 7470
rect 3605 7470 3645 7480
rect 3605 7440 3610 7470
rect 3640 7440 3645 7470
rect 3805 7470 3845 7480
rect 3805 7440 3810 7470
rect 3840 7440 3845 7470
rect 4005 7470 4045 7480
rect 4005 7440 4010 7470
rect 4040 7440 4045 7470
rect 4205 7470 4245 7480
rect 4205 7440 4210 7470
rect 4240 7440 4245 7470
rect 4405 7470 4445 7480
rect 4405 7440 4410 7470
rect 4440 7440 4445 7470
rect 4605 7470 4645 7480
rect 4605 7440 4610 7470
rect 4640 7440 4645 7470
rect 4805 7470 4845 7480
rect 4805 7440 4810 7470
rect 4840 7440 4845 7470
rect 5005 7470 5045 7480
rect 5005 7440 5010 7470
rect 5040 7440 5045 7470
rect 5205 7470 5245 7480
rect 5205 7440 5210 7470
rect 5240 7440 5245 7470
rect 5405 7470 5445 7480
rect 5405 7440 5410 7470
rect 5440 7440 5445 7470
rect 5605 7470 5645 7480
rect 5605 7440 5610 7470
rect 5640 7440 5645 7470
rect 5805 7470 5845 7480
rect 5805 7440 5810 7470
rect 5840 7440 5845 7470
rect 6005 7470 6045 7480
rect 6005 7440 6010 7470
rect 6040 7440 6045 7470
rect 6205 7470 6245 7480
rect 6205 7440 6210 7470
rect 6240 7440 6245 7470
rect 6405 7470 6445 7480
rect 6405 7440 6410 7470
rect 6440 7440 6445 7470
rect -188 7355 -185 7440
rect -165 7355 -162 7440
rect 15 7355 35 7440
rect 215 7355 235 7440
rect 415 7355 435 7440
rect 615 7355 635 7440
rect 815 7355 835 7440
rect 1015 7355 1035 7440
rect 1215 7355 1235 7440
rect 1615 7355 1635 7440
rect 1815 7355 1835 7440
rect 2015 7355 2035 7440
rect 2215 7355 2235 7440
rect 2415 7355 2435 7440
rect 2615 7355 2635 7440
rect 2815 7355 2835 7440
rect 3015 7355 3035 7440
rect 3215 7355 3235 7440
rect 3415 7355 3435 7440
rect 3615 7355 3635 7440
rect 4015 7355 4035 7440
rect 4215 7355 4235 7440
rect 4415 7355 4435 7440
rect 4615 7355 4635 7440
rect 4815 7355 4835 7440
rect 5015 7355 5035 7440
rect 5215 7355 5235 7440
rect 5415 7355 5435 7440
rect 5615 7355 5635 7440
rect 5815 7355 5835 7440
rect 6015 7355 6035 7440
rect 6215 7355 6235 7440
rect -195 7325 -190 7355
rect -160 7325 -155 7355
rect -195 7285 -185 7325
rect -165 7315 -155 7325
rect 5 7325 10 7355
rect 40 7325 45 7355
rect 5 7315 45 7325
rect 205 7325 210 7355
rect 240 7325 245 7355
rect 205 7315 245 7325
rect 405 7325 410 7355
rect 440 7325 445 7355
rect 405 7315 445 7325
rect 605 7325 610 7355
rect 640 7325 645 7355
rect 605 7315 645 7325
rect 805 7325 810 7355
rect 840 7325 845 7355
rect 805 7315 845 7325
rect 1005 7325 1010 7355
rect 1040 7325 1045 7355
rect 1005 7315 1045 7325
rect 1205 7325 1210 7355
rect 1240 7325 1245 7355
rect 1205 7315 1245 7325
rect 1405 7325 1410 7355
rect 1440 7325 1445 7355
rect 1405 7315 1445 7325
rect 1605 7325 1610 7355
rect 1640 7325 1645 7355
rect 1605 7315 1645 7325
rect 1805 7325 1810 7355
rect 1840 7325 1845 7355
rect 1805 7315 1845 7325
rect 2005 7325 2010 7355
rect 2040 7325 2045 7355
rect 2005 7315 2045 7325
rect 2205 7325 2210 7355
rect 2240 7325 2245 7355
rect 2205 7315 2245 7325
rect 2405 7325 2410 7355
rect 2440 7325 2445 7355
rect 2405 7315 2445 7325
rect 2605 7325 2610 7355
rect 2640 7325 2645 7355
rect 2605 7315 2645 7325
rect 2805 7325 2810 7355
rect 2840 7325 2845 7355
rect 2805 7315 2845 7325
rect 3005 7325 3010 7355
rect 3040 7325 3045 7355
rect 3005 7315 3045 7325
rect 3205 7325 3210 7355
rect 3240 7325 3245 7355
rect 3205 7315 3245 7325
rect 3405 7325 3410 7355
rect 3440 7325 3445 7355
rect 3405 7315 3445 7325
rect 3605 7325 3610 7355
rect 3640 7325 3645 7355
rect 3605 7315 3645 7325
rect 3805 7325 3810 7355
rect 3840 7325 3845 7355
rect 3805 7315 3845 7325
rect 4005 7325 4010 7355
rect 4040 7325 4045 7355
rect 4005 7315 4045 7325
rect 4205 7325 4210 7355
rect 4240 7325 4245 7355
rect 4205 7315 4245 7325
rect 4405 7325 4410 7355
rect 4440 7325 4445 7355
rect 4405 7315 4445 7325
rect 4605 7325 4610 7355
rect 4640 7325 4645 7355
rect 4605 7315 4645 7325
rect 4805 7325 4810 7355
rect 4840 7325 4845 7355
rect 4805 7315 4845 7325
rect 5005 7325 5010 7355
rect 5040 7325 5045 7355
rect 5005 7315 5045 7325
rect 5205 7325 5210 7355
rect 5240 7325 5245 7355
rect 5205 7315 5245 7325
rect 5405 7325 5410 7355
rect 5440 7325 5445 7355
rect 5405 7315 5445 7325
rect 5605 7325 5610 7355
rect 5640 7325 5645 7355
rect 5605 7315 5645 7325
rect 5805 7325 5810 7355
rect 5840 7325 5845 7355
rect 5805 7315 5845 7325
rect 6005 7325 6010 7355
rect 6040 7325 6045 7355
rect 6005 7315 6045 7325
rect 6205 7325 6210 7355
rect 6240 7325 6245 7355
rect 6205 7315 6245 7325
rect 6405 7325 6410 7355
rect 6440 7325 6445 7355
rect 6405 7315 6445 7325
rect -165 7295 -30 7315
rect 5 7295 1370 7315
rect 1405 7295 2970 7315
rect 3005 7295 3770 7315
rect 3805 7295 6570 7315
rect -165 7285 -155 7295
rect -195 7255 -190 7285
rect -160 7255 -155 7285
rect 5 7285 45 7295
rect 5 7255 10 7285
rect 40 7255 45 7285
rect 205 7285 245 7295
rect 205 7255 210 7285
rect 240 7255 245 7285
rect 405 7285 445 7295
rect 405 7255 410 7285
rect 440 7255 445 7285
rect 605 7285 645 7295
rect 605 7255 610 7285
rect 640 7255 645 7285
rect 805 7285 845 7295
rect 805 7255 810 7285
rect 840 7255 845 7285
rect 1005 7285 1045 7295
rect 1005 7255 1010 7285
rect 1040 7255 1045 7285
rect 1205 7285 1245 7295
rect 1205 7255 1210 7285
rect 1240 7255 1245 7285
rect 1405 7285 1445 7295
rect 1405 7255 1410 7285
rect 1440 7255 1445 7285
rect 1605 7285 1645 7295
rect 1605 7255 1610 7285
rect 1640 7255 1645 7285
rect 1805 7285 1845 7295
rect 1805 7255 1810 7285
rect 1840 7255 1845 7285
rect 2005 7285 2045 7295
rect 2005 7255 2010 7285
rect 2040 7255 2045 7285
rect 2205 7285 2245 7295
rect 2205 7255 2210 7285
rect 2240 7255 2245 7285
rect 2405 7285 2445 7295
rect 2405 7255 2410 7285
rect 2440 7255 2445 7285
rect 2605 7285 2645 7295
rect 2605 7255 2610 7285
rect 2640 7255 2645 7285
rect 2805 7285 2845 7295
rect 2805 7255 2810 7285
rect 2840 7255 2845 7285
rect 3005 7285 3045 7295
rect 3005 7255 3010 7285
rect 3040 7255 3045 7285
rect 3205 7285 3245 7295
rect 3205 7255 3210 7285
rect 3240 7255 3245 7285
rect 3405 7285 3445 7295
rect 3405 7255 3410 7285
rect 3440 7255 3445 7285
rect 3605 7285 3645 7295
rect 3605 7255 3610 7285
rect 3640 7255 3645 7285
rect 3805 7285 3845 7295
rect 3805 7255 3810 7285
rect 3840 7255 3845 7285
rect 4005 7285 4045 7295
rect 4005 7255 4010 7285
rect 4040 7255 4045 7285
rect 4205 7285 4245 7295
rect 4205 7255 4210 7285
rect 4240 7255 4245 7285
rect 4405 7285 4445 7295
rect 4405 7255 4410 7285
rect 4440 7255 4445 7285
rect 4605 7285 4645 7295
rect 4605 7255 4610 7285
rect 4640 7255 4645 7285
rect 4805 7285 4845 7295
rect 4805 7255 4810 7285
rect 4840 7255 4845 7285
rect 5005 7285 5045 7295
rect 5005 7255 5010 7285
rect 5040 7255 5045 7285
rect 5205 7285 5245 7295
rect 5205 7255 5210 7285
rect 5240 7255 5245 7285
rect 5405 7285 5445 7295
rect 5405 7255 5410 7285
rect 5440 7255 5445 7285
rect 5605 7285 5645 7295
rect 5605 7255 5610 7285
rect 5640 7255 5645 7285
rect 5805 7285 5845 7295
rect 5805 7255 5810 7285
rect 5840 7255 5845 7285
rect 6005 7285 6045 7295
rect 6005 7255 6010 7285
rect 6040 7255 6045 7285
rect 6205 7285 6245 7295
rect 6205 7255 6210 7285
rect 6240 7255 6245 7285
rect 6405 7285 6445 7295
rect 6405 7255 6410 7285
rect 6440 7255 6445 7285
rect -188 7170 -185 7255
rect -165 7170 -162 7255
rect 15 7170 35 7255
rect 215 7170 235 7255
rect 415 7170 435 7255
rect 615 7170 635 7255
rect 815 7170 835 7255
rect 1015 7170 1035 7255
rect 1215 7170 1235 7255
rect 1415 7170 1435 7255
rect 1615 7170 1635 7255
rect 1815 7170 1835 7255
rect 2015 7170 2035 7255
rect 2215 7170 2235 7255
rect 2415 7170 2435 7255
rect 2615 7170 2635 7255
rect 2815 7170 2835 7255
rect 3015 7170 3035 7255
rect 3215 7170 3235 7255
rect 3415 7170 3435 7255
rect 3615 7170 3635 7255
rect 3815 7170 3835 7255
rect 4015 7170 4035 7255
rect 4215 7170 4235 7255
rect 4415 7170 4435 7255
rect -195 7140 -190 7170
rect -160 7140 -155 7170
rect -195 7100 -185 7140
rect -165 7130 -155 7140
rect 5 7140 10 7170
rect 40 7140 45 7170
rect 5 7130 45 7140
rect 205 7140 210 7170
rect 240 7140 245 7170
rect 205 7130 245 7140
rect 405 7140 410 7170
rect 440 7140 445 7170
rect 405 7130 445 7140
rect 605 7140 610 7170
rect 640 7140 645 7170
rect 605 7130 645 7140
rect 805 7140 810 7170
rect 840 7140 845 7170
rect 805 7130 845 7140
rect 1005 7140 1010 7170
rect 1040 7140 1045 7170
rect 1005 7130 1045 7140
rect 1205 7140 1210 7170
rect 1240 7140 1245 7170
rect 1205 7130 1245 7140
rect 1405 7140 1410 7170
rect 1440 7140 1445 7170
rect 1405 7130 1445 7140
rect 1605 7140 1610 7170
rect 1640 7140 1645 7170
rect 1605 7130 1645 7140
rect 1805 7140 1810 7170
rect 1840 7140 1845 7170
rect 1805 7130 1845 7140
rect 2005 7140 2010 7170
rect 2040 7140 2045 7170
rect 2005 7130 2045 7140
rect 2205 7140 2210 7170
rect 2240 7140 2245 7170
rect 2205 7130 2245 7140
rect 2405 7140 2410 7170
rect 2440 7140 2445 7170
rect 2405 7130 2445 7140
rect 2605 7140 2610 7170
rect 2640 7140 2645 7170
rect 2605 7130 2645 7140
rect 2805 7140 2810 7170
rect 2840 7140 2845 7170
rect 2805 7130 2845 7140
rect 3005 7140 3010 7170
rect 3040 7140 3045 7170
rect 3005 7130 3045 7140
rect 3205 7140 3210 7170
rect 3240 7140 3245 7170
rect 3205 7130 3245 7140
rect 3405 7140 3410 7170
rect 3440 7140 3445 7170
rect 3405 7130 3445 7140
rect 3605 7140 3610 7170
rect 3640 7140 3645 7170
rect 3605 7130 3645 7140
rect 3805 7140 3810 7170
rect 3840 7140 3845 7170
rect 3805 7130 3845 7140
rect 4005 7140 4010 7170
rect 4040 7140 4045 7170
rect 4005 7130 4045 7140
rect 4205 7140 4210 7170
rect 4240 7140 4245 7170
rect 4205 7130 4245 7140
rect 4405 7140 4410 7170
rect 4440 7140 4445 7170
rect 4405 7130 4445 7140
rect 4605 7140 4610 7170
rect 4640 7140 4645 7170
rect 4605 7130 4645 7140
rect 4805 7140 4810 7170
rect 4840 7140 4845 7170
rect 4805 7130 4845 7140
rect 5005 7140 5010 7170
rect 5040 7140 5045 7170
rect 5005 7130 5045 7140
rect 5205 7140 5210 7170
rect 5240 7140 5245 7170
rect 5205 7130 5245 7140
rect 5405 7140 5410 7170
rect 5440 7140 5445 7170
rect 5405 7130 5445 7140
rect 5605 7140 5610 7170
rect 5640 7140 5645 7170
rect 5605 7130 5645 7140
rect 5805 7140 5810 7170
rect 5840 7140 5845 7170
rect 5805 7130 5845 7140
rect 6005 7140 6010 7170
rect 6040 7140 6045 7170
rect 6005 7130 6045 7140
rect 6205 7140 6210 7170
rect 6240 7140 6245 7170
rect 6205 7130 6245 7140
rect 6405 7140 6410 7170
rect 6440 7140 6445 7170
rect 6405 7130 6445 7140
rect -165 7110 -30 7130
rect 5 7110 1370 7130
rect 1405 7110 2970 7130
rect 3005 7110 3770 7130
rect 3805 7110 4170 7130
rect 4205 7110 4370 7130
rect 4405 7110 4570 7130
rect 4605 7110 6570 7130
rect -165 7100 -155 7110
rect -195 7070 -190 7100
rect -160 7070 -155 7100
rect 5 7100 45 7110
rect 5 7070 10 7100
rect 40 7070 45 7100
rect 205 7100 245 7110
rect 205 7070 210 7100
rect 240 7070 245 7100
rect 405 7100 445 7110
rect 405 7070 410 7100
rect 440 7070 445 7100
rect 605 7100 645 7110
rect 605 7070 610 7100
rect 640 7070 645 7100
rect 805 7100 845 7110
rect 805 7070 810 7100
rect 840 7070 845 7100
rect 1005 7100 1045 7110
rect 1005 7070 1010 7100
rect 1040 7070 1045 7100
rect 1205 7100 1245 7110
rect 1205 7070 1210 7100
rect 1240 7070 1245 7100
rect 1405 7100 1445 7110
rect 1405 7070 1410 7100
rect 1440 7070 1445 7100
rect 1605 7100 1645 7110
rect 1605 7070 1610 7100
rect 1640 7070 1645 7100
rect 1805 7100 1845 7110
rect 1805 7070 1810 7100
rect 1840 7070 1845 7100
rect 2005 7100 2045 7110
rect 2005 7070 2010 7100
rect 2040 7070 2045 7100
rect 2205 7100 2245 7110
rect 2205 7070 2210 7100
rect 2240 7070 2245 7100
rect 2405 7100 2445 7110
rect 2405 7070 2410 7100
rect 2440 7070 2445 7100
rect 2605 7100 2645 7110
rect 2605 7070 2610 7100
rect 2640 7070 2645 7100
rect 2805 7100 2845 7110
rect 2805 7070 2810 7100
rect 2840 7070 2845 7100
rect 3005 7100 3045 7110
rect 3005 7070 3010 7100
rect 3040 7070 3045 7100
rect 3205 7100 3245 7110
rect 3205 7070 3210 7100
rect 3240 7070 3245 7100
rect 3405 7100 3445 7110
rect 3405 7070 3410 7100
rect 3440 7070 3445 7100
rect 3605 7100 3645 7110
rect 3605 7070 3610 7100
rect 3640 7070 3645 7100
rect 3805 7100 3845 7110
rect 3805 7070 3810 7100
rect 3840 7070 3845 7100
rect 4005 7100 4045 7110
rect 4005 7070 4010 7100
rect 4040 7070 4045 7100
rect 4205 7100 4245 7110
rect 4205 7070 4210 7100
rect 4240 7070 4245 7100
rect 4405 7100 4445 7110
rect 4405 7070 4410 7100
rect 4440 7070 4445 7100
rect 4605 7100 4645 7110
rect 4605 7070 4610 7100
rect 4640 7070 4645 7100
rect 4805 7100 4845 7110
rect 4805 7070 4810 7100
rect 4840 7070 4845 7100
rect 5005 7100 5045 7110
rect 5005 7070 5010 7100
rect 5040 7070 5045 7100
rect 5205 7100 5245 7110
rect 5205 7070 5210 7100
rect 5240 7070 5245 7100
rect 5405 7100 5445 7110
rect 5405 7070 5410 7100
rect 5440 7070 5445 7100
rect 5605 7100 5645 7110
rect 5605 7070 5610 7100
rect 5640 7070 5645 7100
rect 5805 7100 5845 7110
rect 5805 7070 5810 7100
rect 5840 7070 5845 7100
rect 6005 7100 6045 7110
rect 6005 7070 6010 7100
rect 6040 7070 6045 7100
rect 6205 7100 6245 7110
rect 6205 7070 6210 7100
rect 6240 7070 6245 7100
rect 6405 7100 6445 7110
rect 6405 7070 6410 7100
rect 6440 7070 6445 7100
rect -188 6985 -185 7070
rect -165 6985 -162 7070
rect 15 6985 35 7070
rect 215 6985 235 7070
rect 415 6985 435 7070
rect 615 6985 635 7070
rect 815 6985 835 7070
rect 1015 6985 1035 7070
rect 1215 6985 1235 7070
rect 1415 6985 1435 7070
rect 1615 6985 1635 7070
rect 1815 6985 1835 7070
rect 2015 6985 2035 7070
rect 2215 6985 2235 7070
rect 2415 6985 2435 7070
rect 2615 6985 2635 7070
rect 2815 6985 2835 7070
rect 3015 6985 3035 7070
rect 3215 6985 3235 7070
rect 3415 6985 3435 7070
rect 3615 6985 3635 7070
rect 3815 6985 3835 7070
rect 4015 6985 4035 7070
rect 4215 6985 4235 7070
rect 4415 6985 4435 7070
rect 4615 6985 4635 7070
rect 4815 6985 4835 7070
rect 5015 6985 5035 7070
rect 5215 6985 5235 7070
rect 5415 6985 5435 7070
rect 5615 6985 5635 7070
rect 5815 6985 5835 7070
rect 6015 6985 6035 7070
rect 6215 6985 6235 7070
rect -195 6955 -190 6985
rect -160 6955 -155 6985
rect -195 6915 -185 6955
rect -165 6945 -155 6955
rect 5 6955 10 6985
rect 40 6955 45 6985
rect 5 6945 45 6955
rect 205 6955 210 6985
rect 240 6955 245 6985
rect 205 6945 245 6955
rect 405 6955 410 6985
rect 440 6955 445 6985
rect 405 6945 445 6955
rect 605 6955 610 6985
rect 640 6955 645 6985
rect 605 6945 645 6955
rect 805 6955 810 6985
rect 840 6955 845 6985
rect 805 6945 845 6955
rect 1005 6955 1010 6985
rect 1040 6955 1045 6985
rect 1005 6945 1045 6955
rect 1205 6955 1210 6985
rect 1240 6955 1245 6985
rect 1205 6945 1245 6955
rect 1405 6955 1410 6985
rect 1440 6955 1445 6985
rect 1405 6945 1445 6955
rect 1605 6955 1610 6985
rect 1640 6955 1645 6985
rect 1605 6945 1645 6955
rect 1805 6955 1810 6985
rect 1840 6955 1845 6985
rect 1805 6945 1845 6955
rect 2005 6955 2010 6985
rect 2040 6955 2045 6985
rect 2005 6945 2045 6955
rect 2205 6955 2210 6985
rect 2240 6955 2245 6985
rect 2205 6945 2245 6955
rect 2405 6955 2410 6985
rect 2440 6955 2445 6985
rect 2405 6945 2445 6955
rect 2605 6955 2610 6985
rect 2640 6955 2645 6985
rect 2605 6945 2645 6955
rect 2805 6955 2810 6985
rect 2840 6955 2845 6985
rect 2805 6945 2845 6955
rect 3005 6955 3010 6985
rect 3040 6955 3045 6985
rect 3005 6945 3045 6955
rect 3205 6955 3210 6985
rect 3240 6955 3245 6985
rect 3205 6945 3245 6955
rect 3405 6955 3410 6985
rect 3440 6955 3445 6985
rect 3405 6945 3445 6955
rect 3605 6955 3610 6985
rect 3640 6955 3645 6985
rect 3605 6945 3645 6955
rect 3805 6955 3810 6985
rect 3840 6955 3845 6985
rect 3805 6945 3845 6955
rect 4005 6955 4010 6985
rect 4040 6955 4045 6985
rect 4005 6945 4045 6955
rect 4205 6955 4210 6985
rect 4240 6955 4245 6985
rect 4205 6945 4245 6955
rect 4405 6955 4410 6985
rect 4440 6955 4445 6985
rect 4405 6945 4445 6955
rect 4605 6955 4610 6985
rect 4640 6955 4645 6985
rect 4605 6945 4645 6955
rect 4805 6955 4810 6985
rect 4840 6955 4845 6985
rect 4805 6945 4845 6955
rect 5005 6955 5010 6985
rect 5040 6955 5045 6985
rect 5005 6945 5045 6955
rect 5205 6955 5210 6985
rect 5240 6955 5245 6985
rect 5205 6945 5245 6955
rect 5405 6955 5410 6985
rect 5440 6955 5445 6985
rect 5405 6945 5445 6955
rect 5605 6955 5610 6985
rect 5640 6955 5645 6985
rect 5605 6945 5645 6955
rect 5805 6955 5810 6985
rect 5840 6955 5845 6985
rect 5805 6945 5845 6955
rect 6005 6955 6010 6985
rect 6040 6955 6045 6985
rect 6005 6945 6045 6955
rect 6205 6955 6210 6985
rect 6240 6955 6245 6985
rect 6205 6945 6245 6955
rect 6405 6955 6410 6985
rect 6440 6955 6445 6985
rect 6405 6945 6445 6955
rect -165 6925 -30 6945
rect 5 6925 1370 6945
rect 1405 6925 2970 6945
rect 3005 6925 3770 6945
rect 3805 6925 4170 6945
rect 4205 6925 4370 6945
rect 4405 6925 4570 6945
rect 4605 6925 6570 6945
rect -165 6915 -155 6925
rect -195 6885 -190 6915
rect -160 6885 -155 6915
rect 5 6915 45 6925
rect 5 6885 10 6915
rect 40 6885 45 6915
rect 205 6915 245 6925
rect 205 6885 210 6915
rect 240 6885 245 6915
rect 405 6915 445 6925
rect 405 6885 410 6915
rect 440 6885 445 6915
rect 605 6915 645 6925
rect 605 6885 610 6915
rect 640 6885 645 6915
rect 805 6915 845 6925
rect 805 6885 810 6915
rect 840 6885 845 6915
rect 1005 6915 1045 6925
rect 1005 6885 1010 6915
rect 1040 6885 1045 6915
rect 1205 6915 1245 6925
rect 1205 6885 1210 6915
rect 1240 6885 1245 6915
rect 1405 6915 1445 6925
rect 1405 6885 1410 6915
rect 1440 6885 1445 6915
rect 1605 6915 1645 6925
rect 1605 6885 1610 6915
rect 1640 6885 1645 6915
rect 1805 6915 1845 6925
rect 1805 6885 1810 6915
rect 1840 6885 1845 6915
rect 2005 6915 2045 6925
rect 2005 6885 2010 6915
rect 2040 6885 2045 6915
rect 2205 6915 2245 6925
rect 2205 6885 2210 6915
rect 2240 6885 2245 6915
rect 2405 6915 2445 6925
rect 2405 6885 2410 6915
rect 2440 6885 2445 6915
rect 2605 6915 2645 6925
rect 2605 6885 2610 6915
rect 2640 6885 2645 6915
rect 2805 6915 2845 6925
rect 2805 6885 2810 6915
rect 2840 6885 2845 6915
rect 3005 6915 3045 6925
rect 3005 6885 3010 6915
rect 3040 6885 3045 6915
rect 3205 6915 3245 6925
rect 3205 6885 3210 6915
rect 3240 6885 3245 6915
rect 3405 6915 3445 6925
rect 3405 6885 3410 6915
rect 3440 6885 3445 6915
rect 3605 6915 3645 6925
rect 3605 6885 3610 6915
rect 3640 6885 3645 6915
rect 3805 6915 3845 6925
rect 3805 6885 3810 6915
rect 3840 6885 3845 6915
rect 4005 6915 4045 6925
rect 4005 6885 4010 6915
rect 4040 6885 4045 6915
rect 4205 6915 4245 6925
rect 4205 6885 4210 6915
rect 4240 6885 4245 6915
rect 4405 6915 4445 6925
rect 4405 6885 4410 6915
rect 4440 6885 4445 6915
rect 4605 6915 4645 6925
rect 4605 6885 4610 6915
rect 4640 6885 4645 6915
rect 4805 6915 4845 6925
rect 4805 6885 4810 6915
rect 4840 6885 4845 6915
rect 5005 6915 5045 6925
rect 5005 6885 5010 6915
rect 5040 6885 5045 6915
rect 5205 6915 5245 6925
rect 5205 6885 5210 6915
rect 5240 6885 5245 6915
rect 5405 6915 5445 6925
rect 5405 6885 5410 6915
rect 5440 6885 5445 6915
rect 5605 6915 5645 6925
rect 5605 6885 5610 6915
rect 5640 6885 5645 6915
rect 5805 6915 5845 6925
rect 5805 6885 5810 6915
rect 5840 6885 5845 6915
rect 6005 6915 6045 6925
rect 6005 6885 6010 6915
rect 6040 6885 6045 6915
rect 6205 6915 6245 6925
rect 6205 6885 6210 6915
rect 6240 6885 6245 6915
rect 6405 6915 6445 6925
rect 6405 6885 6410 6915
rect 6440 6885 6445 6915
rect -188 6800 -185 6885
rect -165 6800 -162 6885
rect 15 6800 35 6885
rect 215 6800 235 6885
rect 415 6800 435 6885
rect 615 6800 635 6885
rect 815 6800 835 6885
rect 1015 6800 1035 6885
rect 1215 6800 1235 6885
rect 1415 6800 1435 6885
rect 1615 6800 1635 6885
rect 1815 6800 1835 6885
rect 2015 6800 2035 6885
rect 2215 6800 2235 6885
rect 2415 6800 2435 6885
rect 2615 6800 2635 6885
rect 2815 6800 2835 6885
rect 3015 6800 3035 6885
rect 3215 6800 3235 6885
rect 3415 6800 3435 6885
rect 3615 6800 3635 6885
rect 3815 6800 3835 6885
rect 4015 6800 4035 6885
rect 4215 6800 4235 6885
rect 4415 6800 4435 6885
rect 4615 6800 4635 6885
rect 4815 6800 4835 6885
rect 5015 6800 5035 6885
rect -195 6770 -190 6800
rect -160 6770 -155 6800
rect -195 6730 -185 6770
rect -165 6760 -155 6770
rect 5 6770 10 6800
rect 40 6770 45 6800
rect 5 6760 45 6770
rect 205 6770 210 6800
rect 240 6770 245 6800
rect 205 6760 245 6770
rect 405 6770 410 6800
rect 440 6770 445 6800
rect 405 6760 445 6770
rect 605 6770 610 6800
rect 640 6770 645 6800
rect 605 6760 645 6770
rect 805 6770 810 6800
rect 840 6770 845 6800
rect 805 6760 845 6770
rect 1005 6770 1010 6800
rect 1040 6770 1045 6800
rect 1005 6760 1045 6770
rect 1205 6770 1210 6800
rect 1240 6770 1245 6800
rect 1205 6760 1245 6770
rect 1405 6770 1410 6800
rect 1440 6770 1445 6800
rect 1405 6760 1445 6770
rect 1605 6770 1610 6800
rect 1640 6770 1645 6800
rect 1605 6760 1645 6770
rect 1805 6770 1810 6800
rect 1840 6770 1845 6800
rect 1805 6760 1845 6770
rect 2005 6770 2010 6800
rect 2040 6770 2045 6800
rect 2005 6760 2045 6770
rect 2205 6770 2210 6800
rect 2240 6770 2245 6800
rect 2205 6760 2245 6770
rect 2405 6770 2410 6800
rect 2440 6770 2445 6800
rect 2405 6760 2445 6770
rect 2605 6770 2610 6800
rect 2640 6770 2645 6800
rect 2605 6760 2645 6770
rect 2805 6770 2810 6800
rect 2840 6770 2845 6800
rect 2805 6760 2845 6770
rect 3005 6770 3010 6800
rect 3040 6770 3045 6800
rect 3005 6760 3045 6770
rect 3205 6770 3210 6800
rect 3240 6770 3245 6800
rect 3205 6760 3245 6770
rect 3405 6770 3410 6800
rect 3440 6770 3445 6800
rect 3405 6760 3445 6770
rect 3605 6770 3610 6800
rect 3640 6770 3645 6800
rect 3605 6760 3645 6770
rect 3805 6770 3810 6800
rect 3840 6770 3845 6800
rect 3805 6760 3845 6770
rect 4005 6770 4010 6800
rect 4040 6770 4045 6800
rect 4005 6760 4045 6770
rect 4205 6770 4210 6800
rect 4240 6770 4245 6800
rect 4205 6760 4245 6770
rect 4405 6770 4410 6800
rect 4440 6770 4445 6800
rect 4405 6760 4445 6770
rect 4605 6770 4610 6800
rect 4640 6770 4645 6800
rect 4605 6760 4645 6770
rect 4805 6770 4810 6800
rect 4840 6770 4845 6800
rect 4805 6760 4845 6770
rect 5005 6770 5010 6800
rect 5040 6770 5045 6800
rect 5005 6760 5045 6770
rect 5205 6770 5210 6800
rect 5240 6770 5245 6800
rect 5205 6760 5245 6770
rect 5405 6770 5410 6800
rect 5440 6770 5445 6800
rect 5405 6760 5445 6770
rect 5605 6770 5610 6800
rect 5640 6770 5645 6800
rect 5605 6760 5645 6770
rect 5805 6770 5810 6800
rect 5840 6770 5845 6800
rect 5805 6760 5845 6770
rect 6005 6770 6010 6800
rect 6040 6770 6045 6800
rect 6005 6760 6045 6770
rect 6205 6770 6210 6800
rect 6240 6770 6245 6800
rect 6205 6760 6245 6770
rect 6405 6770 6410 6800
rect 6440 6770 6445 6800
rect 6405 6760 6445 6770
rect -165 6740 -30 6760
rect 5 6740 1370 6760
rect 1405 6740 2970 6760
rect 3005 6740 3770 6760
rect 3805 6740 4170 6760
rect 4205 6740 4370 6760
rect 4405 6740 4570 6760
rect 4605 6740 5170 6760
rect 5205 6740 6570 6760
rect -165 6730 -155 6740
rect -195 6700 -190 6730
rect -160 6700 -155 6730
rect 5 6730 45 6740
rect 5 6700 10 6730
rect 40 6700 45 6730
rect 205 6730 245 6740
rect 205 6700 210 6730
rect 240 6700 245 6730
rect 405 6730 445 6740
rect 405 6700 410 6730
rect 440 6700 445 6730
rect 605 6730 645 6740
rect 605 6700 610 6730
rect 640 6700 645 6730
rect 805 6730 845 6740
rect 805 6700 810 6730
rect 840 6700 845 6730
rect 1005 6730 1045 6740
rect 1005 6700 1010 6730
rect 1040 6700 1045 6730
rect 1205 6730 1245 6740
rect 1205 6700 1210 6730
rect 1240 6700 1245 6730
rect 1405 6730 1445 6740
rect 1405 6700 1410 6730
rect 1440 6700 1445 6730
rect 1605 6730 1645 6740
rect 1605 6700 1610 6730
rect 1640 6700 1645 6730
rect 1805 6730 1845 6740
rect 1805 6700 1810 6730
rect 1840 6700 1845 6730
rect 2005 6730 2045 6740
rect 2005 6700 2010 6730
rect 2040 6700 2045 6730
rect 2205 6730 2245 6740
rect 2205 6700 2210 6730
rect 2240 6700 2245 6730
rect 2405 6730 2445 6740
rect 2405 6700 2410 6730
rect 2440 6700 2445 6730
rect 2605 6730 2645 6740
rect 2605 6700 2610 6730
rect 2640 6700 2645 6730
rect 2805 6730 2845 6740
rect 2805 6700 2810 6730
rect 2840 6700 2845 6730
rect 3005 6730 3045 6740
rect 3005 6700 3010 6730
rect 3040 6700 3045 6730
rect 3205 6730 3245 6740
rect 3205 6700 3210 6730
rect 3240 6700 3245 6730
rect 3405 6730 3445 6740
rect 3405 6700 3410 6730
rect 3440 6700 3445 6730
rect 3605 6730 3645 6740
rect 3605 6700 3610 6730
rect 3640 6700 3645 6730
rect 3805 6730 3845 6740
rect 3805 6700 3810 6730
rect 3840 6700 3845 6730
rect 4005 6730 4045 6740
rect 4005 6700 4010 6730
rect 4040 6700 4045 6730
rect 4205 6730 4245 6740
rect 4205 6700 4210 6730
rect 4240 6700 4245 6730
rect 4405 6730 4445 6740
rect 4405 6700 4410 6730
rect 4440 6700 4445 6730
rect 4605 6730 4645 6740
rect 4605 6700 4610 6730
rect 4640 6700 4645 6730
rect 4805 6730 4845 6740
rect 4805 6700 4810 6730
rect 4840 6700 4845 6730
rect 5005 6730 5045 6740
rect 5005 6700 5010 6730
rect 5040 6700 5045 6730
rect 5205 6730 5245 6740
rect 5205 6700 5210 6730
rect 5240 6700 5245 6730
rect 5405 6730 5445 6740
rect 5405 6700 5410 6730
rect 5440 6700 5445 6730
rect 5605 6730 5645 6740
rect 5605 6700 5610 6730
rect 5640 6700 5645 6730
rect 5805 6730 5845 6740
rect 5805 6700 5810 6730
rect 5840 6700 5845 6730
rect 6005 6730 6045 6740
rect 6005 6700 6010 6730
rect 6040 6700 6045 6730
rect 6205 6730 6245 6740
rect 6205 6700 6210 6730
rect 6240 6700 6245 6730
rect 6405 6730 6445 6740
rect 6405 6700 6410 6730
rect 6440 6700 6445 6730
rect -188 6615 -185 6700
rect -165 6615 -162 6700
rect 15 6615 35 6700
rect 215 6615 235 6700
rect 415 6615 435 6700
rect 615 6615 635 6700
rect 815 6615 835 6700
rect 1015 6615 1035 6700
rect 1215 6615 1235 6700
rect 1415 6615 1435 6700
rect 1615 6615 1635 6700
rect 1815 6615 1835 6700
rect 2015 6615 2035 6700
rect 2215 6615 2235 6700
rect 2415 6615 2435 6700
rect 2615 6615 2635 6700
rect 2815 6615 2835 6700
rect 3015 6615 3035 6700
rect 3215 6615 3235 6700
rect 3415 6615 3435 6700
rect 3615 6615 3635 6700
rect 3815 6615 3835 6700
rect 4015 6615 4035 6700
rect 4215 6615 4235 6700
rect 4415 6615 4435 6700
rect 4615 6615 4635 6700
rect 4815 6615 4835 6700
rect 5015 6615 5035 6700
rect 5215 6615 5235 6700
rect 5415 6615 5435 6700
rect -195 6585 -190 6615
rect -160 6585 -155 6615
rect -195 6545 -185 6585
rect -165 6575 -155 6585
rect 5 6585 10 6615
rect 40 6585 45 6615
rect 5 6575 45 6585
rect 205 6585 210 6615
rect 240 6585 245 6615
rect 205 6575 245 6585
rect 405 6585 410 6615
rect 440 6585 445 6615
rect 405 6575 445 6585
rect 605 6585 610 6615
rect 640 6585 645 6615
rect 605 6575 645 6585
rect 805 6585 810 6615
rect 840 6585 845 6615
rect 805 6575 845 6585
rect 1005 6585 1010 6615
rect 1040 6585 1045 6615
rect 1005 6575 1045 6585
rect 1205 6585 1210 6615
rect 1240 6585 1245 6615
rect 1205 6575 1245 6585
rect 1405 6585 1410 6615
rect 1440 6585 1445 6615
rect 1405 6575 1445 6585
rect 1605 6585 1610 6615
rect 1640 6585 1645 6615
rect 1605 6575 1645 6585
rect 1805 6585 1810 6615
rect 1840 6585 1845 6615
rect 1805 6575 1845 6585
rect 2005 6585 2010 6615
rect 2040 6585 2045 6615
rect 2005 6575 2045 6585
rect 2205 6585 2210 6615
rect 2240 6585 2245 6615
rect 2205 6575 2245 6585
rect 2405 6585 2410 6615
rect 2440 6585 2445 6615
rect 2405 6575 2445 6585
rect 2605 6585 2610 6615
rect 2640 6585 2645 6615
rect 2605 6575 2645 6585
rect 2805 6585 2810 6615
rect 2840 6585 2845 6615
rect 2805 6575 2845 6585
rect 3005 6585 3010 6615
rect 3040 6585 3045 6615
rect 3005 6575 3045 6585
rect 3205 6585 3210 6615
rect 3240 6585 3245 6615
rect 3205 6575 3245 6585
rect 3405 6585 3410 6615
rect 3440 6585 3445 6615
rect 3405 6575 3445 6585
rect 3605 6585 3610 6615
rect 3640 6585 3645 6615
rect 3605 6575 3645 6585
rect 3805 6585 3810 6615
rect 3840 6585 3845 6615
rect 3805 6575 3845 6585
rect 4005 6585 4010 6615
rect 4040 6585 4045 6615
rect 4005 6575 4045 6585
rect 4205 6585 4210 6615
rect 4240 6585 4245 6615
rect 4205 6575 4245 6585
rect 4405 6585 4410 6615
rect 4440 6585 4445 6615
rect 4405 6575 4445 6585
rect 4605 6585 4610 6615
rect 4640 6585 4645 6615
rect 4605 6575 4645 6585
rect 4805 6585 4810 6615
rect 4840 6585 4845 6615
rect 4805 6575 4845 6585
rect 5005 6585 5010 6615
rect 5040 6585 5045 6615
rect 5005 6575 5045 6585
rect 5205 6585 5210 6615
rect 5240 6585 5245 6615
rect 5205 6575 5245 6585
rect 5405 6585 5410 6615
rect 5440 6585 5445 6615
rect 5405 6575 5445 6585
rect 5605 6585 5610 6615
rect 5640 6585 5645 6615
rect 5605 6575 5645 6585
rect 5805 6585 5810 6615
rect 5840 6585 5845 6615
rect 5805 6575 5845 6585
rect 6005 6585 6010 6615
rect 6040 6585 6045 6615
rect 6005 6575 6045 6585
rect 6205 6585 6210 6615
rect 6240 6585 6245 6615
rect 6205 6575 6245 6585
rect 6405 6585 6410 6615
rect 6440 6585 6445 6615
rect 6405 6575 6445 6585
rect -165 6555 -30 6575
rect 5 6555 1370 6575
rect 1405 6555 2970 6575
rect 3005 6555 3770 6575
rect 3805 6555 4170 6575
rect 4205 6555 4370 6575
rect 4405 6555 4570 6575
rect 4605 6555 5170 6575
rect 5205 6555 5570 6575
rect 5605 6555 6570 6575
rect -165 6545 -155 6555
rect -195 6515 -190 6545
rect -160 6515 -155 6545
rect 5 6545 45 6555
rect 5 6515 10 6545
rect 40 6515 45 6545
rect 205 6545 245 6555
rect 205 6515 210 6545
rect 240 6515 245 6545
rect 405 6545 445 6555
rect 405 6515 410 6545
rect 440 6515 445 6545
rect 605 6545 645 6555
rect 605 6515 610 6545
rect 640 6515 645 6545
rect 805 6545 845 6555
rect 805 6515 810 6545
rect 840 6515 845 6545
rect 1005 6545 1045 6555
rect 1005 6515 1010 6545
rect 1040 6515 1045 6545
rect 1205 6545 1245 6555
rect 1205 6515 1210 6545
rect 1240 6515 1245 6545
rect 1405 6545 1445 6555
rect 1405 6515 1410 6545
rect 1440 6515 1445 6545
rect 1605 6545 1645 6555
rect 1605 6515 1610 6545
rect 1640 6515 1645 6545
rect 1805 6545 1845 6555
rect 1805 6515 1810 6545
rect 1840 6515 1845 6545
rect 2005 6545 2045 6555
rect 2005 6515 2010 6545
rect 2040 6515 2045 6545
rect 2205 6545 2245 6555
rect 2205 6515 2210 6545
rect 2240 6515 2245 6545
rect 2405 6545 2445 6555
rect 2405 6515 2410 6545
rect 2440 6515 2445 6545
rect 2605 6545 2645 6555
rect 2605 6515 2610 6545
rect 2640 6515 2645 6545
rect 2805 6545 2845 6555
rect 2805 6515 2810 6545
rect 2840 6515 2845 6545
rect 3005 6545 3045 6555
rect 3005 6515 3010 6545
rect 3040 6515 3045 6545
rect 3205 6545 3245 6555
rect 3205 6515 3210 6545
rect 3240 6515 3245 6545
rect 3405 6545 3445 6555
rect 3405 6515 3410 6545
rect 3440 6515 3445 6545
rect 3605 6545 3645 6555
rect 3605 6515 3610 6545
rect 3640 6515 3645 6545
rect 3805 6545 3845 6555
rect 3805 6515 3810 6545
rect 3840 6515 3845 6545
rect 4005 6545 4045 6555
rect 4005 6515 4010 6545
rect 4040 6515 4045 6545
rect 4205 6545 4245 6555
rect 4205 6515 4210 6545
rect 4240 6515 4245 6545
rect 4405 6545 4445 6555
rect 4405 6515 4410 6545
rect 4440 6515 4445 6545
rect 4605 6545 4645 6555
rect 4605 6515 4610 6545
rect 4640 6515 4645 6545
rect 4805 6545 4845 6555
rect 4805 6515 4810 6545
rect 4840 6515 4845 6545
rect 5005 6545 5045 6555
rect 5005 6515 5010 6545
rect 5040 6515 5045 6545
rect 5205 6545 5245 6555
rect 5205 6515 5210 6545
rect 5240 6515 5245 6545
rect 5405 6545 5445 6555
rect 5405 6515 5410 6545
rect 5440 6515 5445 6545
rect 5605 6545 5645 6555
rect 5605 6515 5610 6545
rect 5640 6515 5645 6545
rect 5805 6545 5845 6555
rect 5805 6515 5810 6545
rect 5840 6515 5845 6545
rect 6005 6545 6045 6555
rect 6005 6515 6010 6545
rect 6040 6515 6045 6545
rect 6205 6545 6245 6555
rect 6205 6515 6210 6545
rect 6240 6515 6245 6545
rect 6405 6545 6445 6555
rect 6405 6515 6410 6545
rect 6440 6515 6445 6545
rect -188 6430 -185 6515
rect -165 6430 -162 6515
rect 15 6430 35 6515
rect 215 6430 235 6515
rect 415 6430 435 6515
rect 615 6430 635 6515
rect 815 6430 835 6515
rect 1015 6430 1035 6515
rect 1215 6430 1235 6515
rect 1415 6430 1435 6515
rect 1615 6430 1635 6515
rect 1815 6430 1835 6515
rect 2015 6430 2035 6515
rect 2215 6430 2235 6515
rect 2415 6430 2435 6515
rect 2615 6430 2635 6515
rect 2815 6430 2835 6515
rect 3015 6430 3035 6515
rect 3215 6430 3235 6515
rect 3415 6430 3435 6515
rect 3615 6430 3635 6515
rect 3815 6430 3835 6515
rect 4015 6430 4035 6515
rect 4215 6430 4235 6515
rect 4415 6430 4435 6515
rect 4615 6430 4635 6515
rect 4815 6430 4835 6515
rect 5015 6430 5035 6515
rect 5215 6430 5235 6515
rect 5415 6430 5435 6515
rect 5615 6430 5635 6515
rect -195 6400 -190 6430
rect -160 6400 -155 6430
rect -195 6360 -185 6400
rect -165 6390 -155 6400
rect 5 6400 10 6430
rect 40 6400 45 6430
rect 5 6390 45 6400
rect 205 6400 210 6430
rect 240 6400 245 6430
rect 205 6390 245 6400
rect 405 6400 410 6430
rect 440 6400 445 6430
rect 405 6390 445 6400
rect 605 6400 610 6430
rect 640 6400 645 6430
rect 605 6390 645 6400
rect 805 6400 810 6430
rect 840 6400 845 6430
rect 805 6390 845 6400
rect 1005 6400 1010 6430
rect 1040 6400 1045 6430
rect 1005 6390 1045 6400
rect 1205 6400 1210 6430
rect 1240 6400 1245 6430
rect 1205 6390 1245 6400
rect 1405 6400 1410 6430
rect 1440 6400 1445 6430
rect 1405 6390 1445 6400
rect 1605 6400 1610 6430
rect 1640 6400 1645 6430
rect 1605 6390 1645 6400
rect 1805 6400 1810 6430
rect 1840 6400 1845 6430
rect 1805 6390 1845 6400
rect 2005 6400 2010 6430
rect 2040 6400 2045 6430
rect 2005 6390 2045 6400
rect 2205 6400 2210 6430
rect 2240 6400 2245 6430
rect 2205 6390 2245 6400
rect 2405 6400 2410 6430
rect 2440 6400 2445 6430
rect 2405 6390 2445 6400
rect 2605 6400 2610 6430
rect 2640 6400 2645 6430
rect 2605 6390 2645 6400
rect 2805 6400 2810 6430
rect 2840 6400 2845 6430
rect 2805 6390 2845 6400
rect 3005 6400 3010 6430
rect 3040 6400 3045 6430
rect 3005 6390 3045 6400
rect 3205 6400 3210 6430
rect 3240 6400 3245 6430
rect 3205 6390 3245 6400
rect 3405 6400 3410 6430
rect 3440 6400 3445 6430
rect 3405 6390 3445 6400
rect 3605 6400 3610 6430
rect 3640 6400 3645 6430
rect 3605 6390 3645 6400
rect 3805 6400 3810 6430
rect 3840 6400 3845 6430
rect 3805 6390 3845 6400
rect 4005 6400 4010 6430
rect 4040 6400 4045 6430
rect 4005 6390 4045 6400
rect 4205 6400 4210 6430
rect 4240 6400 4245 6430
rect 4205 6390 4245 6400
rect 4405 6400 4410 6430
rect 4440 6400 4445 6430
rect 4405 6390 4445 6400
rect 4605 6400 4610 6430
rect 4640 6400 4645 6430
rect 4605 6390 4645 6400
rect 4805 6400 4810 6430
rect 4840 6400 4845 6430
rect 4805 6390 4845 6400
rect 5005 6400 5010 6430
rect 5040 6400 5045 6430
rect 5005 6390 5045 6400
rect 5205 6400 5210 6430
rect 5240 6400 5245 6430
rect 5205 6390 5245 6400
rect 5405 6400 5410 6430
rect 5440 6400 5445 6430
rect 5405 6390 5445 6400
rect 5605 6400 5610 6430
rect 5640 6400 5645 6430
rect 5605 6390 5645 6400
rect 5805 6400 5810 6430
rect 5840 6400 5845 6430
rect 5805 6390 5845 6400
rect 6005 6400 6010 6430
rect 6040 6400 6045 6430
rect 6005 6390 6045 6400
rect 6205 6400 6210 6430
rect 6240 6400 6245 6430
rect 6205 6390 6245 6400
rect 6405 6400 6410 6430
rect 6440 6400 6445 6430
rect 6405 6390 6445 6400
rect -165 6370 -30 6390
rect 5 6370 1370 6390
rect 1405 6370 2970 6390
rect 3005 6370 3770 6390
rect 3805 6370 4170 6390
rect 4205 6370 4370 6390
rect 4405 6370 4570 6390
rect 4605 6370 5170 6390
rect 5205 6370 5570 6390
rect 5605 6370 5770 6390
rect 5805 6370 6695 6390
rect -165 6360 -155 6370
rect -195 6330 -190 6360
rect -160 6330 -155 6360
rect 5 6360 45 6370
rect 5 6330 10 6360
rect 40 6330 45 6360
rect 205 6360 245 6370
rect 205 6330 210 6360
rect 240 6330 245 6360
rect 405 6360 445 6370
rect 405 6330 410 6360
rect 440 6330 445 6360
rect 605 6360 645 6370
rect 605 6330 610 6360
rect 640 6330 645 6360
rect 805 6360 845 6370
rect 805 6330 810 6360
rect 840 6330 845 6360
rect 1005 6360 1045 6370
rect 1005 6330 1010 6360
rect 1040 6330 1045 6360
rect 1205 6360 1245 6370
rect 1205 6330 1210 6360
rect 1240 6330 1245 6360
rect 1405 6360 1445 6370
rect 1405 6330 1410 6360
rect 1440 6330 1445 6360
rect 1605 6360 1645 6370
rect 1605 6330 1610 6360
rect 1640 6330 1645 6360
rect 1805 6360 1845 6370
rect 1805 6330 1810 6360
rect 1840 6330 1845 6360
rect 2005 6360 2045 6370
rect 2005 6330 2010 6360
rect 2040 6330 2045 6360
rect 2205 6360 2245 6370
rect 2205 6330 2210 6360
rect 2240 6330 2245 6360
rect 2405 6360 2445 6370
rect 2405 6330 2410 6360
rect 2440 6330 2445 6360
rect 2605 6360 2645 6370
rect 2605 6330 2610 6360
rect 2640 6330 2645 6360
rect 2805 6360 2845 6370
rect 2805 6330 2810 6360
rect 2840 6330 2845 6360
rect 3005 6360 3045 6370
rect 3005 6330 3010 6360
rect 3040 6330 3045 6360
rect 3205 6360 3245 6370
rect 3205 6330 3210 6360
rect 3240 6330 3245 6360
rect 3405 6360 3445 6370
rect 3405 6330 3410 6360
rect 3440 6330 3445 6360
rect 3605 6360 3645 6370
rect 3605 6330 3610 6360
rect 3640 6330 3645 6360
rect 3805 6360 3845 6370
rect 3805 6330 3810 6360
rect 3840 6330 3845 6360
rect 4005 6360 4045 6370
rect 4005 6330 4010 6360
rect 4040 6330 4045 6360
rect 4205 6360 4245 6370
rect 4205 6330 4210 6360
rect 4240 6330 4245 6360
rect 4405 6360 4445 6370
rect 4405 6330 4410 6360
rect 4440 6330 4445 6360
rect 4605 6360 4645 6370
rect 4605 6330 4610 6360
rect 4640 6330 4645 6360
rect 4805 6360 4845 6370
rect 4805 6330 4810 6360
rect 4840 6330 4845 6360
rect 5005 6360 5045 6370
rect 5005 6330 5010 6360
rect 5040 6330 5045 6360
rect 5205 6360 5245 6370
rect 5205 6330 5210 6360
rect 5240 6330 5245 6360
rect 5405 6360 5445 6370
rect 5405 6330 5410 6360
rect 5440 6330 5445 6360
rect 5605 6360 5645 6370
rect 5605 6330 5610 6360
rect 5640 6330 5645 6360
rect 5805 6360 5845 6370
rect 5805 6330 5810 6360
rect 5840 6330 5845 6360
rect 6005 6360 6045 6370
rect 6005 6330 6010 6360
rect 6040 6330 6045 6360
rect 6205 6360 6245 6370
rect 6205 6330 6210 6360
rect 6240 6330 6245 6360
rect 6405 6360 6445 6370
rect 6405 6330 6410 6360
rect 6440 6330 6445 6360
rect -188 6245 -185 6330
rect -165 6245 -162 6330
rect 15 6245 35 6330
rect 215 6245 235 6330
rect 415 6245 435 6330
rect 615 6245 635 6330
rect 815 6245 835 6330
rect 1015 6245 1035 6330
rect 1215 6245 1235 6330
rect 1415 6245 1435 6330
rect 1615 6245 1635 6330
rect 1815 6245 1835 6330
rect 2015 6245 2035 6330
rect 2215 6245 2235 6330
rect 2415 6245 2435 6330
rect 2615 6245 2635 6330
rect 2815 6245 2835 6330
rect 3015 6245 3035 6330
rect 3215 6245 3235 6330
rect 3415 6245 3435 6330
rect 3615 6245 3635 6330
rect 3815 6245 3835 6330
rect 4015 6245 4035 6330
rect 4215 6245 4235 6330
rect 4415 6245 4435 6330
rect 4615 6245 4635 6330
rect 4815 6245 4835 6330
rect 5215 6245 5235 6330
rect 5415 6245 5435 6330
rect 5615 6245 5635 6330
rect 5815 6245 5835 6330
rect -195 6215 -190 6245
rect -160 6215 -155 6245
rect -195 6175 -185 6215
rect -165 6205 -155 6215
rect 5 6215 10 6245
rect 40 6215 45 6245
rect 5 6205 45 6215
rect 205 6215 210 6245
rect 240 6215 245 6245
rect 205 6205 245 6215
rect 405 6215 410 6245
rect 440 6215 445 6245
rect 405 6205 445 6215
rect 605 6215 610 6245
rect 640 6215 645 6245
rect 605 6205 645 6215
rect 805 6215 810 6245
rect 840 6215 845 6245
rect 805 6205 845 6215
rect 1005 6215 1010 6245
rect 1040 6215 1045 6245
rect 1005 6205 1045 6215
rect 1205 6215 1210 6245
rect 1240 6215 1245 6245
rect 1205 6205 1245 6215
rect 1405 6215 1410 6245
rect 1440 6215 1445 6245
rect 1405 6205 1445 6215
rect 1605 6215 1610 6245
rect 1640 6215 1645 6245
rect 1605 6205 1645 6215
rect 1805 6215 1810 6245
rect 1840 6215 1845 6245
rect 1805 6205 1845 6215
rect 2005 6215 2010 6245
rect 2040 6215 2045 6245
rect 2005 6205 2045 6215
rect 2205 6215 2210 6245
rect 2240 6215 2245 6245
rect 2205 6205 2245 6215
rect 2405 6215 2410 6245
rect 2440 6215 2445 6245
rect 2405 6205 2445 6215
rect 2605 6215 2610 6245
rect 2640 6215 2645 6245
rect 2605 6205 2645 6215
rect 2805 6215 2810 6245
rect 2840 6215 2845 6245
rect 2805 6205 2845 6215
rect 3005 6215 3010 6245
rect 3040 6215 3045 6245
rect 3005 6205 3045 6215
rect 3205 6215 3210 6245
rect 3240 6215 3245 6245
rect 3205 6205 3245 6215
rect 3405 6215 3410 6245
rect 3440 6215 3445 6245
rect 3405 6205 3445 6215
rect 3605 6215 3610 6245
rect 3640 6215 3645 6245
rect 3605 6205 3645 6215
rect 3805 6215 3810 6245
rect 3840 6215 3845 6245
rect 3805 6205 3845 6215
rect 4005 6215 4010 6245
rect 4040 6215 4045 6245
rect 4005 6205 4045 6215
rect 4205 6215 4210 6245
rect 4240 6215 4245 6245
rect 4205 6205 4245 6215
rect 4405 6215 4410 6245
rect 4440 6215 4445 6245
rect 4405 6205 4445 6215
rect 4605 6215 4610 6245
rect 4640 6215 4645 6245
rect 4605 6205 4645 6215
rect 4805 6215 4810 6245
rect 4840 6215 4845 6245
rect 4805 6205 4845 6215
rect 5005 6215 5010 6245
rect 5040 6215 5045 6245
rect 5005 6205 5045 6215
rect 5205 6215 5210 6245
rect 5240 6215 5245 6245
rect 5205 6205 5245 6215
rect 5405 6215 5410 6245
rect 5440 6215 5445 6245
rect 5405 6205 5445 6215
rect 5605 6215 5610 6245
rect 5640 6215 5645 6245
rect 5605 6205 5645 6215
rect 5805 6215 5810 6245
rect 5840 6215 5845 6245
rect 5805 6205 5845 6215
rect 6005 6215 6010 6245
rect 6040 6215 6045 6245
rect 6005 6205 6045 6215
rect 6205 6215 6210 6245
rect 6240 6215 6245 6245
rect 6205 6205 6245 6215
rect 6405 6215 6410 6245
rect 6440 6215 6445 6245
rect 6405 6205 6445 6215
rect -165 6185 -30 6205
rect 5 6185 1370 6205
rect 1405 6185 2970 6205
rect 3005 6185 3770 6205
rect 3805 6185 4170 6205
rect 4205 6185 4370 6205
rect 4405 6185 4570 6205
rect 4605 6185 4970 6205
rect 5005 6185 5570 6205
rect 5605 6185 5770 6205
rect 5805 6185 5970 6205
rect 6005 6185 6695 6205
rect -165 6175 -155 6185
rect -195 6145 -190 6175
rect -160 6145 -155 6175
rect 5 6175 45 6185
rect 5 6145 10 6175
rect 40 6145 45 6175
rect 205 6175 245 6185
rect 205 6145 210 6175
rect 240 6145 245 6175
rect 405 6175 445 6185
rect 405 6145 410 6175
rect 440 6145 445 6175
rect 605 6175 645 6185
rect 605 6145 610 6175
rect 640 6145 645 6175
rect 805 6175 845 6185
rect 805 6145 810 6175
rect 840 6145 845 6175
rect 1005 6175 1045 6185
rect 1005 6145 1010 6175
rect 1040 6145 1045 6175
rect 1205 6175 1245 6185
rect 1205 6145 1210 6175
rect 1240 6145 1245 6175
rect 1405 6175 1445 6185
rect 1405 6145 1410 6175
rect 1440 6145 1445 6175
rect 1605 6175 1645 6185
rect 1605 6145 1610 6175
rect 1640 6145 1645 6175
rect 1805 6175 1845 6185
rect 1805 6145 1810 6175
rect 1840 6145 1845 6175
rect 2005 6175 2045 6185
rect 2005 6145 2010 6175
rect 2040 6145 2045 6175
rect 2205 6175 2245 6185
rect 2205 6145 2210 6175
rect 2240 6145 2245 6175
rect 2405 6175 2445 6185
rect 2405 6145 2410 6175
rect 2440 6145 2445 6175
rect 2605 6175 2645 6185
rect 2605 6145 2610 6175
rect 2640 6145 2645 6175
rect 2805 6175 2845 6185
rect 2805 6145 2810 6175
rect 2840 6145 2845 6175
rect 3005 6175 3045 6185
rect 3005 6145 3010 6175
rect 3040 6145 3045 6175
rect 3205 6175 3245 6185
rect 3205 6145 3210 6175
rect 3240 6145 3245 6175
rect 3405 6175 3445 6185
rect 3405 6145 3410 6175
rect 3440 6145 3445 6175
rect 3605 6175 3645 6185
rect 3605 6145 3610 6175
rect 3640 6145 3645 6175
rect 3805 6175 3845 6185
rect 3805 6145 3810 6175
rect 3840 6145 3845 6175
rect 4005 6175 4045 6185
rect 4005 6145 4010 6175
rect 4040 6145 4045 6175
rect 4205 6175 4245 6185
rect 4205 6145 4210 6175
rect 4240 6145 4245 6175
rect 4405 6175 4445 6185
rect 4405 6145 4410 6175
rect 4440 6145 4445 6175
rect 4605 6175 4645 6185
rect 4605 6145 4610 6175
rect 4640 6145 4645 6175
rect 4805 6175 4845 6185
rect 4805 6145 4810 6175
rect 4840 6145 4845 6175
rect 5005 6175 5045 6185
rect 5005 6145 5010 6175
rect 5040 6145 5045 6175
rect 5205 6175 5245 6185
rect 5205 6145 5210 6175
rect 5240 6145 5245 6175
rect 5405 6175 5445 6185
rect 5405 6145 5410 6175
rect 5440 6145 5445 6175
rect 5605 6175 5645 6185
rect 5605 6145 5610 6175
rect 5640 6145 5645 6175
rect 5805 6175 5845 6185
rect 5805 6145 5810 6175
rect 5840 6145 5845 6175
rect 6005 6175 6045 6185
rect 6005 6145 6010 6175
rect 6040 6145 6045 6175
rect 6205 6175 6245 6185
rect 6205 6145 6210 6175
rect 6240 6145 6245 6175
rect 6405 6175 6445 6185
rect 6405 6145 6410 6175
rect 6440 6145 6445 6175
rect -188 6060 -185 6145
rect -165 6060 -162 6145
rect 15 6060 35 6145
rect 215 6060 235 6145
rect 415 6060 435 6145
rect 615 6060 635 6145
rect 815 6060 835 6145
rect 1015 6060 1035 6145
rect 1215 6060 1235 6145
rect 1415 6060 1435 6145
rect 1615 6060 1635 6145
rect 1815 6060 1835 6145
rect 2015 6060 2035 6145
rect 2215 6060 2235 6145
rect 2415 6060 2435 6145
rect 2615 6060 2635 6145
rect 3015 6060 3035 6145
rect 3215 6060 3235 6145
rect 3415 6060 3435 6145
rect 3615 6060 3635 6145
rect 3815 6060 3835 6145
rect 4015 6060 4035 6145
rect 4215 6060 4235 6145
rect 4615 6060 4635 6145
rect 4815 6060 4835 6145
rect 5015 6060 5035 6145
rect 5215 6060 5235 6145
rect 5415 6060 5435 6145
rect 5615 6060 5635 6145
rect 5815 6060 5835 6145
rect -195 6030 -190 6060
rect -160 6030 -155 6060
rect -195 5990 -185 6030
rect -165 6020 -155 6030
rect 5 6030 10 6060
rect 40 6030 45 6060
rect 5 6020 45 6030
rect 205 6030 210 6060
rect 240 6030 245 6060
rect 205 6020 245 6030
rect 405 6030 410 6060
rect 440 6030 445 6060
rect 405 6020 445 6030
rect 605 6030 610 6060
rect 640 6030 645 6060
rect 605 6020 645 6030
rect 805 6030 810 6060
rect 840 6030 845 6060
rect 805 6020 845 6030
rect 1005 6030 1010 6060
rect 1040 6030 1045 6060
rect 1005 6020 1045 6030
rect 1205 6030 1210 6060
rect 1240 6030 1245 6060
rect 1205 6020 1245 6030
rect 1405 6030 1410 6060
rect 1440 6030 1445 6060
rect 1405 6020 1445 6030
rect 1605 6030 1610 6060
rect 1640 6030 1645 6060
rect 1605 6020 1645 6030
rect 1805 6030 1810 6060
rect 1840 6030 1845 6060
rect 1805 6020 1845 6030
rect 2005 6030 2010 6060
rect 2040 6030 2045 6060
rect 2005 6020 2045 6030
rect 2205 6030 2210 6060
rect 2240 6030 2245 6060
rect 2205 6020 2245 6030
rect 2405 6030 2410 6060
rect 2440 6030 2445 6060
rect 2405 6020 2445 6030
rect 2605 6030 2610 6060
rect 2640 6030 2645 6060
rect 2605 6020 2645 6030
rect 2805 6030 2810 6060
rect 2840 6030 2845 6060
rect 2805 6020 2845 6030
rect 3005 6030 3010 6060
rect 3040 6030 3045 6060
rect 3005 6020 3045 6030
rect 3205 6030 3210 6060
rect 3240 6030 3245 6060
rect 3205 6020 3245 6030
rect 3405 6030 3410 6060
rect 3440 6030 3445 6060
rect 3405 6020 3445 6030
rect 3605 6030 3610 6060
rect 3640 6030 3645 6060
rect 3605 6020 3645 6030
rect 3805 6030 3810 6060
rect 3840 6030 3845 6060
rect 3805 6020 3845 6030
rect 4005 6030 4010 6060
rect 4040 6030 4045 6060
rect 4005 6020 4045 6030
rect 4205 6030 4210 6060
rect 4240 6030 4245 6060
rect 4205 6020 4245 6030
rect 4405 6030 4410 6060
rect 4440 6030 4445 6060
rect 4405 6020 4445 6030
rect 4605 6030 4610 6060
rect 4640 6030 4645 6060
rect 4605 6020 4645 6030
rect 4805 6030 4810 6060
rect 4840 6030 4845 6060
rect 4805 6020 4845 6030
rect 5005 6030 5010 6060
rect 5040 6030 5045 6060
rect 5005 6020 5045 6030
rect 5205 6030 5210 6060
rect 5240 6030 5245 6060
rect 5205 6020 5245 6030
rect 5405 6030 5410 6060
rect 5440 6030 5445 6060
rect 5405 6020 5445 6030
rect 5605 6030 5610 6060
rect 5640 6030 5645 6060
rect 5605 6020 5645 6030
rect 5805 6030 5810 6060
rect 5840 6030 5845 6060
rect 5805 6020 5845 6030
rect 6005 6030 6010 6060
rect 6040 6030 6045 6060
rect 6005 6020 6045 6030
rect 6205 6030 6210 6060
rect 6240 6030 6245 6060
rect 6205 6020 6245 6030
rect 6405 6030 6410 6060
rect 6440 6030 6445 6060
rect 6405 6020 6445 6030
rect -165 6000 -30 6020
rect 5 6000 1370 6020
rect 1405 6000 2770 6020
rect 2805 6000 3770 6020
rect 3805 6000 4170 6020
rect 4205 6000 4370 6020
rect 4405 6000 4970 6020
rect 5005 6000 5570 6020
rect 5605 6000 5770 6020
rect 5805 6000 5970 6020
rect 6005 6000 6170 6020
rect 6205 6000 6695 6020
rect -165 5990 -155 6000
rect -195 5960 -190 5990
rect -160 5960 -155 5990
rect 5 5990 45 6000
rect 5 5960 10 5990
rect 40 5960 45 5990
rect 205 5990 245 6000
rect 205 5960 210 5990
rect 240 5960 245 5990
rect 405 5990 445 6000
rect 405 5960 410 5990
rect 440 5960 445 5990
rect 605 5990 645 6000
rect 605 5960 610 5990
rect 640 5960 645 5990
rect 805 5990 845 6000
rect 805 5960 810 5990
rect 840 5960 845 5990
rect 1005 5990 1045 6000
rect 1005 5960 1010 5990
rect 1040 5960 1045 5990
rect 1205 5990 1245 6000
rect 1205 5960 1210 5990
rect 1240 5960 1245 5990
rect 1405 5990 1445 6000
rect 1405 5960 1410 5990
rect 1440 5960 1445 5990
rect 1605 5990 1645 6000
rect 1605 5960 1610 5990
rect 1640 5960 1645 5990
rect 1805 5990 1845 6000
rect 1805 5960 1810 5990
rect 1840 5960 1845 5990
rect 2005 5990 2045 6000
rect 2005 5960 2010 5990
rect 2040 5960 2045 5990
rect 2205 5990 2245 6000
rect 2205 5960 2210 5990
rect 2240 5960 2245 5990
rect 2405 5990 2445 6000
rect 2405 5960 2410 5990
rect 2440 5960 2445 5990
rect 2605 5990 2645 6000
rect 2605 5960 2610 5990
rect 2640 5960 2645 5990
rect 2805 5990 2845 6000
rect 2805 5960 2810 5990
rect 2840 5960 2845 5990
rect 3005 5990 3045 6000
rect 3005 5960 3010 5990
rect 3040 5960 3045 5990
rect 3205 5990 3245 6000
rect 3205 5960 3210 5990
rect 3240 5960 3245 5990
rect 3405 5990 3445 6000
rect 3405 5960 3410 5990
rect 3440 5960 3445 5990
rect 3605 5990 3645 6000
rect 3605 5960 3610 5990
rect 3640 5960 3645 5990
rect 3805 5990 3845 6000
rect 3805 5960 3810 5990
rect 3840 5960 3845 5990
rect 4005 5990 4045 6000
rect 4005 5960 4010 5990
rect 4040 5960 4045 5990
rect 4205 5990 4245 6000
rect 4205 5960 4210 5990
rect 4240 5960 4245 5990
rect 4405 5990 4445 6000
rect 4405 5960 4410 5990
rect 4440 5960 4445 5990
rect 4605 5990 4645 6000
rect 4605 5960 4610 5990
rect 4640 5960 4645 5990
rect 4805 5990 4845 6000
rect 4805 5960 4810 5990
rect 4840 5960 4845 5990
rect 5005 5990 5045 6000
rect 5005 5960 5010 5990
rect 5040 5960 5045 5990
rect 5205 5990 5245 6000
rect 5205 5960 5210 5990
rect 5240 5960 5245 5990
rect 5405 5990 5445 6000
rect 5405 5960 5410 5990
rect 5440 5960 5445 5990
rect 5605 5990 5645 6000
rect 5605 5960 5610 5990
rect 5640 5960 5645 5990
rect 5805 5990 5845 6000
rect 5805 5960 5810 5990
rect 5840 5960 5845 5990
rect 6005 5990 6045 6000
rect 6005 5960 6010 5990
rect 6040 5960 6045 5990
rect 6205 5990 6245 6000
rect 6205 5960 6210 5990
rect 6240 5960 6245 5990
rect 6405 5990 6445 6000
rect 6405 5960 6410 5990
rect 6440 5960 6445 5990
rect -188 5875 -185 5960
rect -165 5875 -162 5960
rect 15 5875 35 5960
rect 215 5875 235 5960
rect 415 5875 435 5960
rect 615 5875 635 5960
rect 815 5875 835 5960
rect 1015 5875 1035 5960
rect 1215 5875 1235 5960
rect 1415 5875 1435 5960
rect 1615 5875 1635 5960
rect 1815 5875 1835 5960
rect 2015 5875 2035 5960
rect 2215 5875 2235 5960
rect 2415 5875 2435 5960
rect 2615 5875 2635 5960
rect 2815 5875 2835 5960
rect 3015 5875 3035 5960
rect 3215 5875 3235 5960
rect 3415 5875 3435 5960
rect 3615 5875 3635 5960
rect 3815 5875 3835 5960
rect 4015 5875 4035 5960
rect 4215 5875 4235 5960
rect 4415 5875 4435 5960
rect 4615 5875 4635 5960
rect 4815 5875 4835 5960
rect 5015 5875 5035 5960
rect 5215 5875 5235 5960
rect 5415 5875 5435 5960
rect 5615 5875 5635 5960
rect 5815 5875 5835 5960
rect 6015 5875 6035 5960
rect -195 5845 -190 5875
rect -160 5845 -155 5875
rect -195 5805 -185 5845
rect -165 5835 -155 5845
rect 5 5845 10 5875
rect 40 5845 45 5875
rect 5 5835 45 5845
rect 205 5845 210 5875
rect 240 5845 245 5875
rect 205 5835 245 5845
rect 405 5845 410 5875
rect 440 5845 445 5875
rect 405 5835 445 5845
rect 605 5845 610 5875
rect 640 5845 645 5875
rect 605 5835 645 5845
rect 805 5845 810 5875
rect 840 5845 845 5875
rect 805 5835 845 5845
rect 1005 5845 1010 5875
rect 1040 5845 1045 5875
rect 1005 5835 1045 5845
rect 1205 5845 1210 5875
rect 1240 5845 1245 5875
rect 1205 5835 1245 5845
rect 1405 5845 1410 5875
rect 1440 5845 1445 5875
rect 1405 5835 1445 5845
rect 1605 5845 1610 5875
rect 1640 5845 1645 5875
rect 1605 5835 1645 5845
rect 1805 5845 1810 5875
rect 1840 5845 1845 5875
rect 1805 5835 1845 5845
rect 2005 5845 2010 5875
rect 2040 5845 2045 5875
rect 2005 5835 2045 5845
rect 2205 5845 2210 5875
rect 2240 5845 2245 5875
rect 2205 5835 2245 5845
rect 2405 5845 2410 5875
rect 2440 5845 2445 5875
rect 2405 5835 2445 5845
rect 2605 5845 2610 5875
rect 2640 5845 2645 5875
rect 2605 5835 2645 5845
rect 2805 5845 2810 5875
rect 2840 5845 2845 5875
rect 2805 5835 2845 5845
rect 3005 5845 3010 5875
rect 3040 5845 3045 5875
rect 3005 5835 3045 5845
rect 3205 5845 3210 5875
rect 3240 5845 3245 5875
rect 3205 5835 3245 5845
rect 3405 5845 3410 5875
rect 3440 5845 3445 5875
rect 3405 5835 3445 5845
rect 3605 5845 3610 5875
rect 3640 5845 3645 5875
rect 3605 5835 3645 5845
rect 3805 5845 3810 5875
rect 3840 5845 3845 5875
rect 3805 5835 3845 5845
rect 4005 5845 4010 5875
rect 4040 5845 4045 5875
rect 4005 5835 4045 5845
rect 4205 5845 4210 5875
rect 4240 5845 4245 5875
rect 4205 5835 4245 5845
rect 4405 5845 4410 5875
rect 4440 5845 4445 5875
rect 4405 5835 4445 5845
rect 4605 5845 4610 5875
rect 4640 5845 4645 5875
rect 4605 5835 4645 5845
rect 4805 5845 4810 5875
rect 4840 5845 4845 5875
rect 4805 5835 4845 5845
rect 5005 5845 5010 5875
rect 5040 5845 5045 5875
rect 5005 5835 5045 5845
rect 5205 5845 5210 5875
rect 5240 5845 5245 5875
rect 5205 5835 5245 5845
rect 5405 5845 5410 5875
rect 5440 5845 5445 5875
rect 5405 5835 5445 5845
rect 5605 5845 5610 5875
rect 5640 5845 5645 5875
rect 5605 5835 5645 5845
rect 5805 5845 5810 5875
rect 5840 5845 5845 5875
rect 5805 5835 5845 5845
rect 6005 5845 6010 5875
rect 6040 5845 6045 5875
rect 6005 5835 6045 5845
rect 6205 5845 6210 5875
rect 6240 5845 6245 5875
rect 6205 5835 6245 5845
rect 6405 5845 6410 5875
rect 6440 5845 6445 5875
rect 6405 5835 6445 5845
rect -165 5815 -30 5835
rect 5 5815 1370 5835
rect 1405 5815 2770 5835
rect 2805 5815 3770 5835
rect 3805 5815 4170 5835
rect 4205 5815 4370 5835
rect 4405 5815 4970 5835
rect 5005 5815 5570 5835
rect 5605 5815 5770 5835
rect 5805 5815 5970 5835
rect 6005 5815 6170 5835
rect 6205 5815 6695 5835
rect -165 5805 -155 5815
rect -195 5775 -190 5805
rect -160 5775 -155 5805
rect 5 5805 45 5815
rect 5 5775 10 5805
rect 40 5775 45 5805
rect 205 5805 245 5815
rect 205 5775 210 5805
rect 240 5775 245 5805
rect 405 5805 445 5815
rect 405 5775 410 5805
rect 440 5775 445 5805
rect 605 5805 645 5815
rect 605 5775 610 5805
rect 640 5775 645 5805
rect 805 5805 845 5815
rect 805 5775 810 5805
rect 840 5775 845 5805
rect 1005 5805 1045 5815
rect 1005 5775 1010 5805
rect 1040 5775 1045 5805
rect 1205 5805 1245 5815
rect 1205 5775 1210 5805
rect 1240 5775 1245 5805
rect 1405 5805 1445 5815
rect 1405 5775 1410 5805
rect 1440 5775 1445 5805
rect 1605 5805 1645 5815
rect 1605 5775 1610 5805
rect 1640 5775 1645 5805
rect 1805 5805 1845 5815
rect 1805 5775 1810 5805
rect 1840 5775 1845 5805
rect 2005 5805 2045 5815
rect 2005 5775 2010 5805
rect 2040 5775 2045 5805
rect 2205 5805 2245 5815
rect 2205 5775 2210 5805
rect 2240 5775 2245 5805
rect 2405 5805 2445 5815
rect 2405 5775 2410 5805
rect 2440 5775 2445 5805
rect 2605 5805 2645 5815
rect 2605 5775 2610 5805
rect 2640 5775 2645 5805
rect 2805 5805 2845 5815
rect 2805 5775 2810 5805
rect 2840 5775 2845 5805
rect 3005 5805 3045 5815
rect 3005 5775 3010 5805
rect 3040 5775 3045 5805
rect 3205 5805 3245 5815
rect 3205 5775 3210 5805
rect 3240 5775 3245 5805
rect 3405 5805 3445 5815
rect 3405 5775 3410 5805
rect 3440 5775 3445 5805
rect 3605 5805 3645 5815
rect 3605 5775 3610 5805
rect 3640 5775 3645 5805
rect 3805 5805 3845 5815
rect 3805 5775 3810 5805
rect 3840 5775 3845 5805
rect 4005 5805 4045 5815
rect 4005 5775 4010 5805
rect 4040 5775 4045 5805
rect 4205 5805 4245 5815
rect 4205 5775 4210 5805
rect 4240 5775 4245 5805
rect 4405 5805 4445 5815
rect 4405 5775 4410 5805
rect 4440 5775 4445 5805
rect 4605 5805 4645 5815
rect 4605 5775 4610 5805
rect 4640 5775 4645 5805
rect 4805 5805 4845 5815
rect 4805 5775 4810 5805
rect 4840 5775 4845 5805
rect 5005 5805 5045 5815
rect 5005 5775 5010 5805
rect 5040 5775 5045 5805
rect 5205 5805 5245 5815
rect 5205 5775 5210 5805
rect 5240 5775 5245 5805
rect 5405 5805 5445 5815
rect 5405 5775 5410 5805
rect 5440 5775 5445 5805
rect 5605 5805 5645 5815
rect 5605 5775 5610 5805
rect 5640 5775 5645 5805
rect 5805 5805 5845 5815
rect 5805 5775 5810 5805
rect 5840 5775 5845 5805
rect 6005 5805 6045 5815
rect 6005 5775 6010 5805
rect 6040 5775 6045 5805
rect 6205 5805 6245 5815
rect 6205 5775 6210 5805
rect 6240 5775 6245 5805
rect 6405 5805 6445 5815
rect 6405 5775 6410 5805
rect 6440 5775 6445 5805
rect -188 5690 -185 5775
rect -165 5690 -162 5775
rect 15 5690 35 5775
rect 215 5690 235 5775
rect 415 5690 435 5775
rect 615 5690 635 5775
rect 815 5690 835 5775
rect 1015 5690 1035 5775
rect 1215 5690 1235 5775
rect 1415 5690 1435 5775
rect 1615 5690 1635 5775
rect 1815 5690 1835 5775
rect 2015 5690 2035 5775
rect 2215 5690 2235 5775
rect 2415 5690 2435 5775
rect 2615 5690 2635 5775
rect 3015 5690 3035 5775
rect 3215 5690 3235 5775
rect 3415 5690 3435 5775
rect 3615 5690 3635 5775
rect 3815 5690 3835 5775
rect 4015 5690 4035 5775
rect 4215 5690 4235 5775
rect 4615 5690 4635 5775
rect 4815 5690 4835 5775
rect 5015 5690 5035 5775
rect 5215 5690 5235 5775
rect 5415 5690 5435 5775
rect 5615 5690 5635 5775
rect 5815 5690 5835 5775
rect 6015 5690 6035 5775
rect -195 5660 -190 5690
rect -160 5660 -155 5690
rect -195 5620 -185 5660
rect -165 5650 -155 5660
rect 5 5660 10 5690
rect 40 5660 45 5690
rect 5 5650 45 5660
rect 205 5660 210 5690
rect 240 5660 245 5690
rect 205 5650 245 5660
rect 405 5660 410 5690
rect 440 5660 445 5690
rect 405 5650 445 5660
rect 605 5660 610 5690
rect 640 5660 645 5690
rect 605 5650 645 5660
rect 805 5660 810 5690
rect 840 5660 845 5690
rect 805 5650 845 5660
rect 1005 5660 1010 5690
rect 1040 5660 1045 5690
rect 1005 5650 1045 5660
rect 1205 5660 1210 5690
rect 1240 5660 1245 5690
rect 1205 5650 1245 5660
rect 1405 5660 1410 5690
rect 1440 5660 1445 5690
rect 1405 5650 1445 5660
rect 1605 5660 1610 5690
rect 1640 5660 1645 5690
rect 1605 5650 1645 5660
rect 1805 5660 1810 5690
rect 1840 5660 1845 5690
rect 1805 5650 1845 5660
rect 2005 5660 2010 5690
rect 2040 5660 2045 5690
rect 2005 5650 2045 5660
rect 2205 5660 2210 5690
rect 2240 5660 2245 5690
rect 2205 5650 2245 5660
rect 2405 5660 2410 5690
rect 2440 5660 2445 5690
rect 2405 5650 2445 5660
rect 2605 5660 2610 5690
rect 2640 5660 2645 5690
rect 2605 5650 2645 5660
rect 2805 5660 2810 5690
rect 2840 5660 2845 5690
rect 2805 5650 2845 5660
rect 3005 5660 3010 5690
rect 3040 5660 3045 5690
rect 3005 5650 3045 5660
rect 3205 5660 3210 5690
rect 3240 5660 3245 5690
rect 3205 5650 3245 5660
rect 3405 5660 3410 5690
rect 3440 5660 3445 5690
rect 3405 5650 3445 5660
rect 3605 5660 3610 5690
rect 3640 5660 3645 5690
rect 3605 5650 3645 5660
rect 3805 5660 3810 5690
rect 3840 5660 3845 5690
rect 3805 5650 3845 5660
rect 4005 5660 4010 5690
rect 4040 5660 4045 5690
rect 4005 5650 4045 5660
rect 4205 5660 4210 5690
rect 4240 5660 4245 5690
rect 4205 5650 4245 5660
rect 4405 5660 4410 5690
rect 4440 5660 4445 5690
rect 4405 5650 4445 5660
rect 4605 5660 4610 5690
rect 4640 5660 4645 5690
rect 4605 5650 4645 5660
rect 4805 5660 4810 5690
rect 4840 5660 4845 5690
rect 4805 5650 4845 5660
rect 5005 5660 5010 5690
rect 5040 5660 5045 5690
rect 5005 5650 5045 5660
rect 5205 5660 5210 5690
rect 5240 5660 5245 5690
rect 5205 5650 5245 5660
rect 5405 5660 5410 5690
rect 5440 5660 5445 5690
rect 5405 5650 5445 5660
rect 5605 5660 5610 5690
rect 5640 5660 5645 5690
rect 5605 5650 5645 5660
rect 5805 5660 5810 5690
rect 5840 5660 5845 5690
rect 5805 5650 5845 5660
rect 6005 5660 6010 5690
rect 6040 5660 6045 5690
rect 6005 5650 6045 5660
rect 6205 5660 6210 5690
rect 6240 5660 6245 5690
rect 6205 5650 6245 5660
rect 6405 5660 6410 5690
rect 6440 5660 6445 5690
rect 6405 5650 6445 5660
rect -165 5630 -30 5650
rect 5 5630 1370 5650
rect 1405 5630 2970 5650
rect 3005 5630 3770 5650
rect 3805 5630 4170 5650
rect 4205 5630 4370 5650
rect 4405 5630 4570 5650
rect 4605 5630 4970 5650
rect 5005 5630 5570 5650
rect 5605 5630 5770 5650
rect 5805 5630 5970 5650
rect 6005 5630 6695 5650
rect -165 5620 -155 5630
rect -195 5590 -190 5620
rect -160 5590 -155 5620
rect 5 5620 45 5630
rect 5 5590 10 5620
rect 40 5590 45 5620
rect 205 5620 245 5630
rect 205 5590 210 5620
rect 240 5590 245 5620
rect 405 5620 445 5630
rect 405 5590 410 5620
rect 440 5590 445 5620
rect 605 5620 645 5630
rect 605 5590 610 5620
rect 640 5590 645 5620
rect 805 5620 845 5630
rect 805 5590 810 5620
rect 840 5590 845 5620
rect 1005 5620 1045 5630
rect 1005 5590 1010 5620
rect 1040 5590 1045 5620
rect 1205 5620 1245 5630
rect 1205 5590 1210 5620
rect 1240 5590 1245 5620
rect 1405 5620 1445 5630
rect 1405 5590 1410 5620
rect 1440 5590 1445 5620
rect 1605 5620 1645 5630
rect 1605 5590 1610 5620
rect 1640 5590 1645 5620
rect 1805 5620 1845 5630
rect 1805 5590 1810 5620
rect 1840 5590 1845 5620
rect 2005 5620 2045 5630
rect 2005 5590 2010 5620
rect 2040 5590 2045 5620
rect 2205 5620 2245 5630
rect 2205 5590 2210 5620
rect 2240 5590 2245 5620
rect 2405 5620 2445 5630
rect 2405 5590 2410 5620
rect 2440 5590 2445 5620
rect 2605 5620 2645 5630
rect 2605 5590 2610 5620
rect 2640 5590 2645 5620
rect 2805 5620 2845 5630
rect 2805 5590 2810 5620
rect 2840 5590 2845 5620
rect 3005 5620 3045 5630
rect 3005 5590 3010 5620
rect 3040 5590 3045 5620
rect 3205 5620 3245 5630
rect 3205 5590 3210 5620
rect 3240 5590 3245 5620
rect 3405 5620 3445 5630
rect 3405 5590 3410 5620
rect 3440 5590 3445 5620
rect 3605 5620 3645 5630
rect 3605 5590 3610 5620
rect 3640 5590 3645 5620
rect 3805 5620 3845 5630
rect 3805 5590 3810 5620
rect 3840 5590 3845 5620
rect 4005 5620 4045 5630
rect 4005 5590 4010 5620
rect 4040 5590 4045 5620
rect 4205 5620 4245 5630
rect 4205 5590 4210 5620
rect 4240 5590 4245 5620
rect 4405 5620 4445 5630
rect 4405 5590 4410 5620
rect 4440 5590 4445 5620
rect 4605 5620 4645 5630
rect 4605 5590 4610 5620
rect 4640 5590 4645 5620
rect 4805 5620 4845 5630
rect 4805 5590 4810 5620
rect 4840 5590 4845 5620
rect 5005 5620 5045 5630
rect 5005 5590 5010 5620
rect 5040 5590 5045 5620
rect 5205 5620 5245 5630
rect 5205 5590 5210 5620
rect 5240 5590 5245 5620
rect 5405 5620 5445 5630
rect 5405 5590 5410 5620
rect 5440 5590 5445 5620
rect 5605 5620 5645 5630
rect 5605 5590 5610 5620
rect 5640 5590 5645 5620
rect 5805 5620 5845 5630
rect 5805 5590 5810 5620
rect 5840 5590 5845 5620
rect 6005 5620 6045 5630
rect 6005 5590 6010 5620
rect 6040 5590 6045 5620
rect 6205 5620 6245 5630
rect 6205 5590 6210 5620
rect 6240 5590 6245 5620
rect 6405 5620 6445 5630
rect 6405 5590 6410 5620
rect 6440 5590 6445 5620
rect -188 5505 -185 5590
rect -165 5505 -162 5590
rect 15 5505 35 5590
rect 215 5505 235 5590
rect 415 5505 435 5590
rect 615 5505 635 5590
rect 815 5505 835 5590
rect 1015 5505 1035 5590
rect 1215 5505 1235 5590
rect 1415 5505 1435 5590
rect 1615 5505 1635 5590
rect 1815 5505 1835 5590
rect 2015 5505 2035 5590
rect 2215 5505 2235 5590
rect 2415 5505 2435 5590
rect 2615 5505 2635 5590
rect 2815 5505 2835 5590
rect 3015 5505 3035 5590
rect 3215 5505 3235 5590
rect 3415 5505 3435 5590
rect 3615 5505 3635 5590
rect 3815 5505 3835 5590
rect 4015 5505 4035 5590
rect 4215 5505 4235 5590
rect 4415 5505 4435 5590
rect 4615 5505 4635 5590
rect 4815 5505 4835 5590
rect 5215 5505 5235 5590
rect 5415 5505 5435 5590
rect 5615 5505 5635 5590
rect 5815 5505 5835 5590
rect -195 5475 -190 5505
rect -160 5475 -155 5505
rect -195 5435 -185 5475
rect -165 5465 -155 5475
rect 5 5475 10 5505
rect 40 5475 45 5505
rect 5 5465 45 5475
rect 205 5475 210 5505
rect 240 5475 245 5505
rect 205 5465 245 5475
rect 405 5475 410 5505
rect 440 5475 445 5505
rect 405 5465 445 5475
rect 605 5475 610 5505
rect 640 5475 645 5505
rect 605 5465 645 5475
rect 805 5475 810 5505
rect 840 5475 845 5505
rect 805 5465 845 5475
rect 1005 5475 1010 5505
rect 1040 5475 1045 5505
rect 1005 5465 1045 5475
rect 1205 5475 1210 5505
rect 1240 5475 1245 5505
rect 1205 5465 1245 5475
rect 1405 5475 1410 5505
rect 1440 5475 1445 5505
rect 1405 5465 1445 5475
rect 1605 5475 1610 5505
rect 1640 5475 1645 5505
rect 1605 5465 1645 5475
rect 1805 5475 1810 5505
rect 1840 5475 1845 5505
rect 1805 5465 1845 5475
rect 2005 5475 2010 5505
rect 2040 5475 2045 5505
rect 2005 5465 2045 5475
rect 2205 5475 2210 5505
rect 2240 5475 2245 5505
rect 2205 5465 2245 5475
rect 2405 5475 2410 5505
rect 2440 5475 2445 5505
rect 2405 5465 2445 5475
rect 2605 5475 2610 5505
rect 2640 5475 2645 5505
rect 2605 5465 2645 5475
rect 2805 5475 2810 5505
rect 2840 5475 2845 5505
rect 2805 5465 2845 5475
rect 3005 5475 3010 5505
rect 3040 5475 3045 5505
rect 3005 5465 3045 5475
rect 3205 5475 3210 5505
rect 3240 5475 3245 5505
rect 3205 5465 3245 5475
rect 3405 5475 3410 5505
rect 3440 5475 3445 5505
rect 3405 5465 3445 5475
rect 3605 5475 3610 5505
rect 3640 5475 3645 5505
rect 3605 5465 3645 5475
rect 3805 5475 3810 5505
rect 3840 5475 3845 5505
rect 3805 5465 3845 5475
rect 4005 5475 4010 5505
rect 4040 5475 4045 5505
rect 4005 5465 4045 5475
rect 4205 5475 4210 5505
rect 4240 5475 4245 5505
rect 4205 5465 4245 5475
rect 4405 5475 4410 5505
rect 4440 5475 4445 5505
rect 4405 5465 4445 5475
rect 4605 5475 4610 5505
rect 4640 5475 4645 5505
rect 4605 5465 4645 5475
rect 4805 5475 4810 5505
rect 4840 5475 4845 5505
rect 4805 5465 4845 5475
rect 5005 5475 5010 5505
rect 5040 5475 5045 5505
rect 5005 5465 5045 5475
rect 5205 5475 5210 5505
rect 5240 5475 5245 5505
rect 5205 5465 5245 5475
rect 5405 5475 5410 5505
rect 5440 5475 5445 5505
rect 5405 5465 5445 5475
rect 5605 5475 5610 5505
rect 5640 5475 5645 5505
rect 5605 5465 5645 5475
rect 5805 5475 5810 5505
rect 5840 5475 5845 5505
rect 5805 5465 5845 5475
rect 6005 5475 6010 5505
rect 6040 5475 6045 5505
rect 6005 5465 6045 5475
rect 6205 5475 6210 5505
rect 6240 5475 6245 5505
rect 6205 5465 6245 5475
rect 6405 5475 6410 5505
rect 6440 5475 6445 5505
rect 6405 5465 6445 5475
rect -165 5445 -30 5465
rect 5 5445 1370 5465
rect 1405 5445 2970 5465
rect 3005 5445 3770 5465
rect 3805 5445 4170 5465
rect 4205 5445 4370 5465
rect 4405 5445 4570 5465
rect 4605 5445 5170 5465
rect 5205 5445 5570 5465
rect 5605 5445 5770 5465
rect 5805 5445 5970 5465
rect 6005 5445 6695 5465
rect -165 5435 -155 5445
rect -195 5405 -190 5435
rect -160 5405 -155 5435
rect 5 5435 45 5445
rect 5 5405 10 5435
rect 40 5405 45 5435
rect 205 5435 245 5445
rect 205 5405 210 5435
rect 240 5405 245 5435
rect 405 5435 445 5445
rect 405 5405 410 5435
rect 440 5405 445 5435
rect 605 5435 645 5445
rect 605 5405 610 5435
rect 640 5405 645 5435
rect 805 5435 845 5445
rect 805 5405 810 5435
rect 840 5405 845 5435
rect 1005 5435 1045 5445
rect 1005 5405 1010 5435
rect 1040 5405 1045 5435
rect 1205 5435 1245 5445
rect 1205 5405 1210 5435
rect 1240 5405 1245 5435
rect 1405 5435 1445 5445
rect 1405 5405 1410 5435
rect 1440 5405 1445 5435
rect 1605 5435 1645 5445
rect 1605 5405 1610 5435
rect 1640 5405 1645 5435
rect 1805 5435 1845 5445
rect 1805 5405 1810 5435
rect 1840 5405 1845 5435
rect 2005 5435 2045 5445
rect 2005 5405 2010 5435
rect 2040 5405 2045 5435
rect 2205 5435 2245 5445
rect 2205 5405 2210 5435
rect 2240 5405 2245 5435
rect 2405 5435 2445 5445
rect 2405 5405 2410 5435
rect 2440 5405 2445 5435
rect 2605 5435 2645 5445
rect 2605 5405 2610 5435
rect 2640 5405 2645 5435
rect 2805 5435 2845 5445
rect 2805 5405 2810 5435
rect 2840 5405 2845 5435
rect 3005 5435 3045 5445
rect 3005 5405 3010 5435
rect 3040 5405 3045 5435
rect 3205 5435 3245 5445
rect 3205 5405 3210 5435
rect 3240 5405 3245 5435
rect 3405 5435 3445 5445
rect 3405 5405 3410 5435
rect 3440 5405 3445 5435
rect 3605 5435 3645 5445
rect 3605 5405 3610 5435
rect 3640 5405 3645 5435
rect 3805 5435 3845 5445
rect 3805 5405 3810 5435
rect 3840 5405 3845 5435
rect 4005 5435 4045 5445
rect 4005 5405 4010 5435
rect 4040 5405 4045 5435
rect 4205 5435 4245 5445
rect 4205 5405 4210 5435
rect 4240 5405 4245 5435
rect 4405 5435 4445 5445
rect 4405 5405 4410 5435
rect 4440 5405 4445 5435
rect 4605 5435 4645 5445
rect 4605 5405 4610 5435
rect 4640 5405 4645 5435
rect 4805 5435 4845 5445
rect 4805 5405 4810 5435
rect 4840 5405 4845 5435
rect 5005 5435 5045 5445
rect 5005 5405 5010 5435
rect 5040 5405 5045 5435
rect 5205 5435 5245 5445
rect 5205 5405 5210 5435
rect 5240 5405 5245 5435
rect 5405 5435 5445 5445
rect 5405 5405 5410 5435
rect 5440 5405 5445 5435
rect 5605 5435 5645 5445
rect 5605 5405 5610 5435
rect 5640 5405 5645 5435
rect 5805 5435 5845 5445
rect 5805 5405 5810 5435
rect 5840 5405 5845 5435
rect 6005 5435 6045 5445
rect 6005 5405 6010 5435
rect 6040 5405 6045 5435
rect 6205 5435 6245 5445
rect 6205 5405 6210 5435
rect 6240 5405 6245 5435
rect 6405 5435 6445 5445
rect 6405 5405 6410 5435
rect 6440 5405 6445 5435
rect -188 5320 -185 5405
rect -165 5320 -162 5405
rect 15 5320 35 5405
rect 215 5320 235 5405
rect 415 5320 435 5405
rect 615 5320 635 5405
rect 815 5320 835 5405
rect 1015 5320 1035 5405
rect 1215 5320 1235 5405
rect 1415 5320 1435 5405
rect 1615 5320 1635 5405
rect 1815 5320 1835 5405
rect 2015 5320 2035 5405
rect 2215 5320 2235 5405
rect 2415 5320 2435 5405
rect 2615 5320 2635 5405
rect 2815 5320 2835 5405
rect 3015 5320 3035 5405
rect 3215 5320 3235 5405
rect 3415 5320 3435 5405
rect 3615 5320 3635 5405
rect 3815 5320 3835 5405
rect 4015 5320 4035 5405
rect 4215 5320 4235 5405
rect 4415 5320 4435 5405
rect 4615 5320 4635 5405
rect 4815 5320 4835 5405
rect 5015 5320 5035 5405
rect 5215 5320 5235 5405
rect 5415 5320 5435 5405
rect 5615 5320 5635 5405
rect 6015 5320 6035 5405
rect 6215 5320 6235 5405
rect -195 5290 -190 5320
rect -160 5290 -155 5320
rect -195 5250 -185 5290
rect -165 5280 -155 5290
rect 5 5290 10 5320
rect 40 5290 45 5320
rect 5 5280 45 5290
rect 205 5290 210 5320
rect 240 5290 245 5320
rect 205 5280 245 5290
rect 405 5290 410 5320
rect 440 5290 445 5320
rect 405 5280 445 5290
rect 605 5290 610 5320
rect 640 5290 645 5320
rect 605 5280 645 5290
rect 805 5290 810 5320
rect 840 5290 845 5320
rect 805 5280 845 5290
rect 1005 5290 1010 5320
rect 1040 5290 1045 5320
rect 1005 5280 1045 5290
rect 1205 5290 1210 5320
rect 1240 5290 1245 5320
rect 1205 5280 1245 5290
rect 1405 5290 1410 5320
rect 1440 5290 1445 5320
rect 1405 5280 1445 5290
rect 1605 5290 1610 5320
rect 1640 5290 1645 5320
rect 1605 5280 1645 5290
rect 1805 5290 1810 5320
rect 1840 5290 1845 5320
rect 1805 5280 1845 5290
rect 2005 5290 2010 5320
rect 2040 5290 2045 5320
rect 2005 5280 2045 5290
rect 2205 5290 2210 5320
rect 2240 5290 2245 5320
rect 2205 5280 2245 5290
rect 2405 5290 2410 5320
rect 2440 5290 2445 5320
rect 2405 5280 2445 5290
rect 2605 5290 2610 5320
rect 2640 5290 2645 5320
rect 2605 5280 2645 5290
rect 2805 5290 2810 5320
rect 2840 5290 2845 5320
rect 2805 5280 2845 5290
rect 3005 5290 3010 5320
rect 3040 5290 3045 5320
rect 3005 5280 3045 5290
rect 3205 5290 3210 5320
rect 3240 5290 3245 5320
rect 3205 5280 3245 5290
rect 3405 5290 3410 5320
rect 3440 5290 3445 5320
rect 3405 5280 3445 5290
rect 3605 5290 3610 5320
rect 3640 5290 3645 5320
rect 3605 5280 3645 5290
rect 3805 5290 3810 5320
rect 3840 5290 3845 5320
rect 3805 5280 3845 5290
rect 4005 5290 4010 5320
rect 4040 5290 4045 5320
rect 4005 5280 4045 5290
rect 4205 5290 4210 5320
rect 4240 5290 4245 5320
rect 4205 5280 4245 5290
rect 4405 5290 4410 5320
rect 4440 5290 4445 5320
rect 4405 5280 4445 5290
rect 4605 5290 4610 5320
rect 4640 5290 4645 5320
rect 4605 5280 4645 5290
rect 4805 5290 4810 5320
rect 4840 5290 4845 5320
rect 4805 5280 4845 5290
rect 5005 5290 5010 5320
rect 5040 5290 5045 5320
rect 5005 5280 5045 5290
rect 5205 5290 5210 5320
rect 5240 5290 5245 5320
rect 5205 5280 5245 5290
rect 5405 5290 5410 5320
rect 5440 5290 5445 5320
rect 5405 5280 5445 5290
rect 5605 5290 5610 5320
rect 5640 5290 5645 5320
rect 5605 5280 5645 5290
rect 5805 5290 5810 5320
rect 5840 5290 5845 5320
rect 5805 5280 5845 5290
rect 6005 5290 6010 5320
rect 6040 5290 6045 5320
rect 6005 5280 6045 5290
rect 6205 5290 6210 5320
rect 6240 5290 6245 5320
rect 6205 5280 6245 5290
rect 6405 5290 6410 5320
rect 6440 5290 6445 5320
rect 6405 5280 6445 5290
rect -165 5260 -30 5280
rect 5 5260 1370 5280
rect 1405 5260 2970 5280
rect 3005 5260 3770 5280
rect 3805 5260 4170 5280
rect 4205 5260 4370 5280
rect 4405 5260 4570 5280
rect 4605 5260 5170 5280
rect 5205 5260 5570 5280
rect 5605 5260 6570 5280
rect -165 5250 -155 5260
rect -195 5220 -190 5250
rect -160 5220 -155 5250
rect 5 5250 45 5260
rect 5 5220 10 5250
rect 40 5220 45 5250
rect 205 5250 245 5260
rect 205 5220 210 5250
rect 240 5220 245 5250
rect 405 5250 445 5260
rect 405 5220 410 5250
rect 440 5220 445 5250
rect 605 5250 645 5260
rect 605 5220 610 5250
rect 640 5220 645 5250
rect 805 5250 845 5260
rect 805 5220 810 5250
rect 840 5220 845 5250
rect 1005 5250 1045 5260
rect 1005 5220 1010 5250
rect 1040 5220 1045 5250
rect 1205 5250 1245 5260
rect 1205 5220 1210 5250
rect 1240 5220 1245 5250
rect 1405 5250 1445 5260
rect 1405 5220 1410 5250
rect 1440 5220 1445 5250
rect 1605 5250 1645 5260
rect 1605 5220 1610 5250
rect 1640 5220 1645 5250
rect 1805 5250 1845 5260
rect 1805 5220 1810 5250
rect 1840 5220 1845 5250
rect 2005 5250 2045 5260
rect 2005 5220 2010 5250
rect 2040 5220 2045 5250
rect 2205 5250 2245 5260
rect 2205 5220 2210 5250
rect 2240 5220 2245 5250
rect 2405 5250 2445 5260
rect 2405 5220 2410 5250
rect 2440 5220 2445 5250
rect 2605 5250 2645 5260
rect 2605 5220 2610 5250
rect 2640 5220 2645 5250
rect 2805 5250 2845 5260
rect 2805 5220 2810 5250
rect 2840 5220 2845 5250
rect 3005 5250 3045 5260
rect 3005 5220 3010 5250
rect 3040 5220 3045 5250
rect 3205 5250 3245 5260
rect 3205 5220 3210 5250
rect 3240 5220 3245 5250
rect 3405 5250 3445 5260
rect 3405 5220 3410 5250
rect 3440 5220 3445 5250
rect 3605 5250 3645 5260
rect 3605 5220 3610 5250
rect 3640 5220 3645 5250
rect 3805 5250 3845 5260
rect 3805 5220 3810 5250
rect 3840 5220 3845 5250
rect 4005 5250 4045 5260
rect 4005 5220 4010 5250
rect 4040 5220 4045 5250
rect 4205 5250 4245 5260
rect 4205 5220 4210 5250
rect 4240 5220 4245 5250
rect 4405 5250 4445 5260
rect 4405 5220 4410 5250
rect 4440 5220 4445 5250
rect 4605 5250 4645 5260
rect 4605 5220 4610 5250
rect 4640 5220 4645 5250
rect 4805 5250 4845 5260
rect 4805 5220 4810 5250
rect 4840 5220 4845 5250
rect 5005 5250 5045 5260
rect 5005 5220 5010 5250
rect 5040 5220 5045 5250
rect 5205 5250 5245 5260
rect 5205 5220 5210 5250
rect 5240 5220 5245 5250
rect 5405 5250 5445 5260
rect 5405 5220 5410 5250
rect 5440 5220 5445 5250
rect 5605 5250 5645 5260
rect 5605 5220 5610 5250
rect 5640 5220 5645 5250
rect 5805 5250 5845 5260
rect 5805 5220 5810 5250
rect 5840 5220 5845 5250
rect 6005 5250 6045 5260
rect 6005 5220 6010 5250
rect 6040 5220 6045 5250
rect 6205 5250 6245 5260
rect 6205 5220 6210 5250
rect 6240 5220 6245 5250
rect 6405 5250 6445 5260
rect 6405 5220 6410 5250
rect 6440 5220 6445 5250
rect -188 5135 -185 5220
rect -165 5135 -162 5220
rect 15 5135 35 5220
rect 215 5135 235 5220
rect 415 5135 435 5220
rect 615 5135 635 5220
rect 815 5135 835 5220
rect 1015 5135 1035 5220
rect 1215 5135 1235 5220
rect 1415 5135 1435 5220
rect 1615 5135 1635 5220
rect 1815 5135 1835 5220
rect 2015 5135 2035 5220
rect 2215 5135 2235 5220
rect 2415 5135 2435 5220
rect 2615 5135 2635 5220
rect 2815 5135 2835 5220
rect 3015 5135 3035 5220
rect 3215 5135 3235 5220
rect 3415 5135 3435 5220
rect 3615 5135 3635 5220
rect 3815 5135 3835 5220
rect 4015 5135 4035 5220
rect 4215 5135 4235 5220
rect 4415 5135 4435 5220
rect 4615 5135 4635 5220
rect 4815 5135 4835 5220
rect 5015 5135 5035 5220
rect 5215 5135 5235 5220
rect 5415 5135 5435 5220
rect -195 5105 -190 5135
rect -160 5105 -155 5135
rect -195 5065 -185 5105
rect -165 5095 -155 5105
rect 5 5105 10 5135
rect 40 5105 45 5135
rect 5 5095 45 5105
rect 205 5105 210 5135
rect 240 5105 245 5135
rect 205 5095 245 5105
rect 405 5105 410 5135
rect 440 5105 445 5135
rect 405 5095 445 5105
rect 605 5105 610 5135
rect 640 5105 645 5135
rect 605 5095 645 5105
rect 805 5105 810 5135
rect 840 5105 845 5135
rect 805 5095 845 5105
rect 1005 5105 1010 5135
rect 1040 5105 1045 5135
rect 1005 5095 1045 5105
rect 1205 5105 1210 5135
rect 1240 5105 1245 5135
rect 1205 5095 1245 5105
rect 1405 5105 1410 5135
rect 1440 5105 1445 5135
rect 1405 5095 1445 5105
rect 1605 5105 1610 5135
rect 1640 5105 1645 5135
rect 1605 5095 1645 5105
rect 1805 5105 1810 5135
rect 1840 5105 1845 5135
rect 1805 5095 1845 5105
rect 2005 5105 2010 5135
rect 2040 5105 2045 5135
rect 2005 5095 2045 5105
rect 2205 5105 2210 5135
rect 2240 5105 2245 5135
rect 2205 5095 2245 5105
rect 2405 5105 2410 5135
rect 2440 5105 2445 5135
rect 2405 5095 2445 5105
rect 2605 5105 2610 5135
rect 2640 5105 2645 5135
rect 2605 5095 2645 5105
rect 2805 5105 2810 5135
rect 2840 5105 2845 5135
rect 2805 5095 2845 5105
rect 3005 5105 3010 5135
rect 3040 5105 3045 5135
rect 3005 5095 3045 5105
rect 3205 5105 3210 5135
rect 3240 5105 3245 5135
rect 3205 5095 3245 5105
rect 3405 5105 3410 5135
rect 3440 5105 3445 5135
rect 3405 5095 3445 5105
rect 3605 5105 3610 5135
rect 3640 5105 3645 5135
rect 3605 5095 3645 5105
rect 3805 5105 3810 5135
rect 3840 5105 3845 5135
rect 3805 5095 3845 5105
rect 4005 5105 4010 5135
rect 4040 5105 4045 5135
rect 4005 5095 4045 5105
rect 4205 5105 4210 5135
rect 4240 5105 4245 5135
rect 4205 5095 4245 5105
rect 4405 5105 4410 5135
rect 4440 5105 4445 5135
rect 4405 5095 4445 5105
rect 4605 5105 4610 5135
rect 4640 5105 4645 5135
rect 4605 5095 4645 5105
rect 4805 5105 4810 5135
rect 4840 5105 4845 5135
rect 4805 5095 4845 5105
rect 5005 5105 5010 5135
rect 5040 5105 5045 5135
rect 5005 5095 5045 5105
rect 5205 5105 5210 5135
rect 5240 5105 5245 5135
rect 5205 5095 5245 5105
rect 5405 5105 5410 5135
rect 5440 5105 5445 5135
rect 5405 5095 5445 5105
rect 5605 5105 5610 5135
rect 5640 5105 5645 5135
rect 5605 5095 5645 5105
rect 5805 5105 5810 5135
rect 5840 5105 5845 5135
rect 5805 5095 5845 5105
rect 6005 5105 6010 5135
rect 6040 5105 6045 5135
rect 6005 5095 6045 5105
rect 6205 5105 6210 5135
rect 6240 5105 6245 5135
rect 6205 5095 6245 5105
rect 6405 5105 6410 5135
rect 6440 5105 6445 5135
rect 6405 5095 6445 5105
rect -165 5075 -30 5095
rect 5 5075 1370 5095
rect 1405 5075 2970 5095
rect 3005 5075 3770 5095
rect 3805 5075 4170 5095
rect 4205 5075 4370 5095
rect 4405 5075 4570 5095
rect 4605 5075 5170 5095
rect 5205 5075 6695 5095
rect -165 5065 -155 5075
rect -195 5035 -190 5065
rect -160 5035 -155 5065
rect 5 5065 45 5075
rect 5 5035 10 5065
rect 40 5035 45 5065
rect 205 5065 245 5075
rect 205 5035 210 5065
rect 240 5035 245 5065
rect 405 5065 445 5075
rect 405 5035 410 5065
rect 440 5035 445 5065
rect 605 5065 645 5075
rect 605 5035 610 5065
rect 640 5035 645 5065
rect 805 5065 845 5075
rect 805 5035 810 5065
rect 840 5035 845 5065
rect 1005 5065 1045 5075
rect 1005 5035 1010 5065
rect 1040 5035 1045 5065
rect 1205 5065 1245 5075
rect 1205 5035 1210 5065
rect 1240 5035 1245 5065
rect 1405 5065 1445 5075
rect 1405 5035 1410 5065
rect 1440 5035 1445 5065
rect 1605 5065 1645 5075
rect 1605 5035 1610 5065
rect 1640 5035 1645 5065
rect 1805 5065 1845 5075
rect 1805 5035 1810 5065
rect 1840 5035 1845 5065
rect 2005 5065 2045 5075
rect 2005 5035 2010 5065
rect 2040 5035 2045 5065
rect 2205 5065 2245 5075
rect 2205 5035 2210 5065
rect 2240 5035 2245 5065
rect 2405 5065 2445 5075
rect 2405 5035 2410 5065
rect 2440 5035 2445 5065
rect 2605 5065 2645 5075
rect 2605 5035 2610 5065
rect 2640 5035 2645 5065
rect 2805 5065 2845 5075
rect 2805 5035 2810 5065
rect 2840 5035 2845 5065
rect 3005 5065 3045 5075
rect 3005 5035 3010 5065
rect 3040 5035 3045 5065
rect 3205 5065 3245 5075
rect 3205 5035 3210 5065
rect 3240 5035 3245 5065
rect 3405 5065 3445 5075
rect 3405 5035 3410 5065
rect 3440 5035 3445 5065
rect 3605 5065 3645 5075
rect 3605 5035 3610 5065
rect 3640 5035 3645 5065
rect 3805 5065 3845 5075
rect 3805 5035 3810 5065
rect 3840 5035 3845 5065
rect 4005 5065 4045 5075
rect 4005 5035 4010 5065
rect 4040 5035 4045 5065
rect 4205 5065 4245 5075
rect 4205 5035 4210 5065
rect 4240 5035 4245 5065
rect 4405 5065 4445 5075
rect 4405 5035 4410 5065
rect 4440 5035 4445 5065
rect 4605 5065 4645 5075
rect 4605 5035 4610 5065
rect 4640 5035 4645 5065
rect 4805 5065 4845 5075
rect 4805 5035 4810 5065
rect 4840 5035 4845 5065
rect 5005 5065 5045 5075
rect 5005 5035 5010 5065
rect 5040 5035 5045 5065
rect 5205 5065 5245 5075
rect 5205 5035 5210 5065
rect 5240 5035 5245 5065
rect 5405 5065 5445 5075
rect 5405 5035 5410 5065
rect 5440 5035 5445 5065
rect 5605 5065 5645 5075
rect 5605 5035 5610 5065
rect 5640 5035 5645 5065
rect 5805 5065 5845 5075
rect 5805 5035 5810 5065
rect 5840 5035 5845 5065
rect 6005 5065 6045 5075
rect 6005 5035 6010 5065
rect 6040 5035 6045 5065
rect 6205 5065 6245 5075
rect 6205 5035 6210 5065
rect 6240 5035 6245 5065
rect 6405 5065 6445 5075
rect 6405 5035 6410 5065
rect 6440 5035 6445 5065
rect -188 4950 -185 5035
rect -165 4950 -162 5035
rect 15 4950 35 5035
rect 215 4950 235 5035
rect 415 4950 435 5035
rect 615 4950 635 5035
rect 815 4950 835 5035
rect 1015 4950 1035 5035
rect 1215 4950 1235 5035
rect 1415 4950 1435 5035
rect 1615 4950 1635 5035
rect 1815 4950 1835 5035
rect 2015 4950 2035 5035
rect 2215 4950 2235 5035
rect 2415 4950 2435 5035
rect 2615 4950 2635 5035
rect 2815 4950 2835 5035
rect 3015 4950 3035 5035
rect 3215 4950 3235 5035
rect 3415 4950 3435 5035
rect 3615 4950 3635 5035
rect 3815 4950 3835 5035
rect 4015 4950 4035 5035
rect 4215 4950 4235 5035
rect 4415 4950 4435 5035
rect 4615 4950 4635 5035
rect 4815 4950 4835 5035
rect 5015 4950 5035 5035
rect -195 4920 -190 4950
rect -160 4920 -155 4950
rect -195 4880 -185 4920
rect -165 4910 -155 4920
rect 5 4920 10 4950
rect 40 4920 45 4950
rect 5 4910 45 4920
rect 205 4920 210 4950
rect 240 4920 245 4950
rect 205 4910 245 4920
rect 405 4920 410 4950
rect 440 4920 445 4950
rect 405 4910 445 4920
rect 605 4920 610 4950
rect 640 4920 645 4950
rect 605 4910 645 4920
rect 805 4920 810 4950
rect 840 4920 845 4950
rect 805 4910 845 4920
rect 1005 4920 1010 4950
rect 1040 4920 1045 4950
rect 1005 4910 1045 4920
rect 1205 4920 1210 4950
rect 1240 4920 1245 4950
rect 1205 4910 1245 4920
rect 1405 4920 1410 4950
rect 1440 4920 1445 4950
rect 1405 4910 1445 4920
rect 1605 4920 1610 4950
rect 1640 4920 1645 4950
rect 1605 4910 1645 4920
rect 1805 4920 1810 4950
rect 1840 4920 1845 4950
rect 1805 4910 1845 4920
rect 2005 4920 2010 4950
rect 2040 4920 2045 4950
rect 2005 4910 2045 4920
rect 2205 4920 2210 4950
rect 2240 4920 2245 4950
rect 2205 4910 2245 4920
rect 2405 4920 2410 4950
rect 2440 4920 2445 4950
rect 2405 4910 2445 4920
rect 2605 4920 2610 4950
rect 2640 4920 2645 4950
rect 2605 4910 2645 4920
rect 2805 4920 2810 4950
rect 2840 4920 2845 4950
rect 2805 4910 2845 4920
rect 3005 4920 3010 4950
rect 3040 4920 3045 4950
rect 3005 4910 3045 4920
rect 3205 4920 3210 4950
rect 3240 4920 3245 4950
rect 3205 4910 3245 4920
rect 3405 4920 3410 4950
rect 3440 4920 3445 4950
rect 3405 4910 3445 4920
rect 3605 4920 3610 4950
rect 3640 4920 3645 4950
rect 3605 4910 3645 4920
rect 3805 4920 3810 4950
rect 3840 4920 3845 4950
rect 3805 4910 3845 4920
rect 4005 4920 4010 4950
rect 4040 4920 4045 4950
rect 4005 4910 4045 4920
rect 4205 4920 4210 4950
rect 4240 4920 4245 4950
rect 4205 4910 4245 4920
rect 4405 4920 4410 4950
rect 4440 4920 4445 4950
rect 4405 4910 4445 4920
rect 4605 4920 4610 4950
rect 4640 4920 4645 4950
rect 4605 4910 4645 4920
rect 4805 4920 4810 4950
rect 4840 4920 4845 4950
rect 4805 4910 4845 4920
rect 5005 4920 5010 4950
rect 5040 4920 5045 4950
rect 5005 4910 5045 4920
rect 5205 4920 5210 4950
rect 5240 4920 5245 4950
rect 5205 4910 5245 4920
rect 5405 4920 5410 4950
rect 5440 4920 5445 4950
rect 5405 4910 5445 4920
rect 5605 4920 5610 4950
rect 5640 4920 5645 4950
rect 5605 4910 5645 4920
rect 5805 4920 5810 4950
rect 5840 4920 5845 4950
rect 5805 4910 5845 4920
rect 6005 4920 6010 4950
rect 6040 4920 6045 4950
rect 6005 4910 6045 4920
rect 6205 4920 6210 4950
rect 6240 4920 6245 4950
rect 6205 4910 6245 4920
rect 6405 4920 6410 4950
rect 6440 4920 6445 4950
rect 6405 4910 6445 4920
rect -165 4890 -30 4910
rect 5 4890 1370 4910
rect 1405 4890 2970 4910
rect 3005 4890 3770 4910
rect 3805 4890 4170 4910
rect 4205 4890 4370 4910
rect 4405 4890 4570 4910
rect 4605 4890 6695 4910
rect -165 4880 -155 4890
rect -195 4850 -190 4880
rect -160 4850 -155 4880
rect 5 4880 45 4890
rect 5 4850 10 4880
rect 40 4850 45 4880
rect 205 4880 245 4890
rect 205 4850 210 4880
rect 240 4850 245 4880
rect 405 4880 445 4890
rect 405 4850 410 4880
rect 440 4850 445 4880
rect 605 4880 645 4890
rect 605 4850 610 4880
rect 640 4850 645 4880
rect 805 4880 845 4890
rect 805 4850 810 4880
rect 840 4850 845 4880
rect 1005 4880 1045 4890
rect 1005 4850 1010 4880
rect 1040 4850 1045 4880
rect 1205 4880 1245 4890
rect 1205 4850 1210 4880
rect 1240 4850 1245 4880
rect 1405 4880 1445 4890
rect 1405 4850 1410 4880
rect 1440 4850 1445 4880
rect 1605 4880 1645 4890
rect 1605 4850 1610 4880
rect 1640 4850 1645 4880
rect 1805 4880 1845 4890
rect 1805 4850 1810 4880
rect 1840 4850 1845 4880
rect 2005 4880 2045 4890
rect 2005 4850 2010 4880
rect 2040 4850 2045 4880
rect 2205 4880 2245 4890
rect 2205 4850 2210 4880
rect 2240 4850 2245 4880
rect 2405 4880 2445 4890
rect 2405 4850 2410 4880
rect 2440 4850 2445 4880
rect 2605 4880 2645 4890
rect 2605 4850 2610 4880
rect 2640 4850 2645 4880
rect 2805 4880 2845 4890
rect 2805 4850 2810 4880
rect 2840 4850 2845 4880
rect 3005 4880 3045 4890
rect 3005 4850 3010 4880
rect 3040 4850 3045 4880
rect 3205 4880 3245 4890
rect 3205 4850 3210 4880
rect 3240 4850 3245 4880
rect 3405 4880 3445 4890
rect 3405 4850 3410 4880
rect 3440 4850 3445 4880
rect 3605 4880 3645 4890
rect 3605 4850 3610 4880
rect 3640 4850 3645 4880
rect 3805 4880 3845 4890
rect 3805 4850 3810 4880
rect 3840 4850 3845 4880
rect 4005 4880 4045 4890
rect 4005 4850 4010 4880
rect 4040 4850 4045 4880
rect 4205 4880 4245 4890
rect 4205 4850 4210 4880
rect 4240 4850 4245 4880
rect 4405 4880 4445 4890
rect 4405 4850 4410 4880
rect 4440 4850 4445 4880
rect 4605 4880 4645 4890
rect 4605 4850 4610 4880
rect 4640 4850 4645 4880
rect 4805 4880 4845 4890
rect 4805 4850 4810 4880
rect 4840 4850 4845 4880
rect 5005 4880 5045 4890
rect 5005 4850 5010 4880
rect 5040 4850 5045 4880
rect 5205 4880 5245 4890
rect 5205 4850 5210 4880
rect 5240 4850 5245 4880
rect 5405 4880 5445 4890
rect 5405 4850 5410 4880
rect 5440 4850 5445 4880
rect 5605 4880 5645 4890
rect 5605 4850 5610 4880
rect 5640 4850 5645 4880
rect 5805 4880 5845 4890
rect 5805 4850 5810 4880
rect 5840 4850 5845 4880
rect 6005 4880 6045 4890
rect 6005 4850 6010 4880
rect 6040 4850 6045 4880
rect 6205 4880 6245 4890
rect 6205 4850 6210 4880
rect 6240 4850 6245 4880
rect 6405 4880 6445 4890
rect 6405 4850 6410 4880
rect 6440 4850 6445 4880
rect -188 4765 -185 4850
rect -165 4765 -162 4850
rect 15 4765 35 4850
rect 215 4765 235 4850
rect 415 4765 435 4850
rect 615 4765 635 4850
rect 815 4765 835 4850
rect 1015 4765 1035 4850
rect 1215 4765 1235 4850
rect 1415 4765 1435 4850
rect 1615 4765 1635 4850
rect 1815 4765 1835 4850
rect 2015 4765 2035 4850
rect 2215 4765 2235 4850
rect 2415 4765 2435 4850
rect 2615 4765 2635 4850
rect 2815 4765 2835 4850
rect 3015 4765 3035 4850
rect 3215 4765 3235 4850
rect 3415 4765 3435 4850
rect 3615 4765 3635 4850
rect 3815 4765 3835 4850
rect 4015 4765 4035 4850
rect 4215 4765 4235 4850
rect 4415 4765 4435 4850
rect 4615 4765 4635 4850
rect 4815 4765 4835 4850
rect 5015 4765 5035 4850
rect 5215 4765 5235 4850
rect 5415 4765 5435 4850
rect 5615 4765 5635 4850
rect 5815 4765 5835 4850
rect 6015 4765 6035 4850
rect 6215 4765 6235 4850
rect -195 4735 -190 4765
rect -160 4735 -155 4765
rect -195 4695 -185 4735
rect -165 4725 -155 4735
rect 5 4735 10 4765
rect 40 4735 45 4765
rect 5 4725 45 4735
rect 205 4735 210 4765
rect 240 4735 245 4765
rect 205 4725 245 4735
rect 405 4735 410 4765
rect 440 4735 445 4765
rect 405 4725 445 4735
rect 605 4735 610 4765
rect 640 4735 645 4765
rect 605 4725 645 4735
rect 805 4735 810 4765
rect 840 4735 845 4765
rect 805 4725 845 4735
rect 1005 4735 1010 4765
rect 1040 4735 1045 4765
rect 1005 4725 1045 4735
rect 1205 4735 1210 4765
rect 1240 4735 1245 4765
rect 1205 4725 1245 4735
rect 1405 4735 1410 4765
rect 1440 4735 1445 4765
rect 1405 4725 1445 4735
rect 1605 4735 1610 4765
rect 1640 4735 1645 4765
rect 1605 4725 1645 4735
rect 1805 4735 1810 4765
rect 1840 4735 1845 4765
rect 1805 4725 1845 4735
rect 2005 4735 2010 4765
rect 2040 4735 2045 4765
rect 2005 4725 2045 4735
rect 2205 4735 2210 4765
rect 2240 4735 2245 4765
rect 2205 4725 2245 4735
rect 2405 4735 2410 4765
rect 2440 4735 2445 4765
rect 2405 4725 2445 4735
rect 2605 4735 2610 4765
rect 2640 4735 2645 4765
rect 2605 4725 2645 4735
rect 2805 4735 2810 4765
rect 2840 4735 2845 4765
rect 2805 4725 2845 4735
rect 3005 4735 3010 4765
rect 3040 4735 3045 4765
rect 3005 4725 3045 4735
rect 3205 4735 3210 4765
rect 3240 4735 3245 4765
rect 3205 4725 3245 4735
rect 3405 4735 3410 4765
rect 3440 4735 3445 4765
rect 3405 4725 3445 4735
rect 3605 4735 3610 4765
rect 3640 4735 3645 4765
rect 3605 4725 3645 4735
rect 3805 4735 3810 4765
rect 3840 4735 3845 4765
rect 3805 4725 3845 4735
rect 4005 4735 4010 4765
rect 4040 4735 4045 4765
rect 4005 4725 4045 4735
rect 4205 4735 4210 4765
rect 4240 4735 4245 4765
rect 4205 4725 4245 4735
rect 4405 4735 4410 4765
rect 4440 4735 4445 4765
rect 4405 4725 4445 4735
rect 4605 4735 4610 4765
rect 4640 4735 4645 4765
rect 4605 4725 4645 4735
rect 4805 4735 4810 4765
rect 4840 4735 4845 4765
rect 4805 4725 4845 4735
rect 5005 4735 5010 4765
rect 5040 4735 5045 4765
rect 5005 4725 5045 4735
rect 5205 4735 5210 4765
rect 5240 4735 5245 4765
rect 5205 4725 5245 4735
rect 5405 4735 5410 4765
rect 5440 4735 5445 4765
rect 5405 4725 5445 4735
rect 5605 4735 5610 4765
rect 5640 4735 5645 4765
rect 5605 4725 5645 4735
rect 5805 4735 5810 4765
rect 5840 4735 5845 4765
rect 5805 4725 5845 4735
rect 6005 4735 6010 4765
rect 6040 4735 6045 4765
rect 6005 4725 6045 4735
rect 6205 4735 6210 4765
rect 6240 4735 6245 4765
rect 6205 4725 6245 4735
rect 6405 4735 6410 4765
rect 6440 4735 6445 4765
rect 6405 4725 6445 4735
rect -165 4705 -30 4725
rect 5 4705 1370 4725
rect 1405 4705 2970 4725
rect 3005 4705 3770 4725
rect 3805 4705 4170 4725
rect 4205 4705 4370 4725
rect 4405 4705 4570 4725
rect 4605 4705 6570 4725
rect -165 4695 -155 4705
rect -195 4665 -190 4695
rect -160 4665 -155 4695
rect 5 4695 45 4705
rect 5 4665 10 4695
rect 40 4665 45 4695
rect 205 4695 245 4705
rect 205 4665 210 4695
rect 240 4665 245 4695
rect 405 4695 445 4705
rect 405 4665 410 4695
rect 440 4665 445 4695
rect 605 4695 645 4705
rect 605 4665 610 4695
rect 640 4665 645 4695
rect 805 4695 845 4705
rect 805 4665 810 4695
rect 840 4665 845 4695
rect 1005 4695 1045 4705
rect 1005 4665 1010 4695
rect 1040 4665 1045 4695
rect 1205 4695 1245 4705
rect 1205 4665 1210 4695
rect 1240 4665 1245 4695
rect 1405 4695 1445 4705
rect 1405 4665 1410 4695
rect 1440 4665 1445 4695
rect 1605 4695 1645 4705
rect 1605 4665 1610 4695
rect 1640 4665 1645 4695
rect 1805 4695 1845 4705
rect 1805 4665 1810 4695
rect 1840 4665 1845 4695
rect 2005 4695 2045 4705
rect 2005 4665 2010 4695
rect 2040 4665 2045 4695
rect 2205 4695 2245 4705
rect 2205 4665 2210 4695
rect 2240 4665 2245 4695
rect 2405 4695 2445 4705
rect 2405 4665 2410 4695
rect 2440 4665 2445 4695
rect 2605 4695 2645 4705
rect 2605 4665 2610 4695
rect 2640 4665 2645 4695
rect 2805 4695 2845 4705
rect 2805 4665 2810 4695
rect 2840 4665 2845 4695
rect 3005 4695 3045 4705
rect 3005 4665 3010 4695
rect 3040 4665 3045 4695
rect 3205 4695 3245 4705
rect 3205 4665 3210 4695
rect 3240 4665 3245 4695
rect 3405 4695 3445 4705
rect 3405 4665 3410 4695
rect 3440 4665 3445 4695
rect 3605 4695 3645 4705
rect 3605 4665 3610 4695
rect 3640 4665 3645 4695
rect 3805 4695 3845 4705
rect 3805 4665 3810 4695
rect 3840 4665 3845 4695
rect 4005 4695 4045 4705
rect 4005 4665 4010 4695
rect 4040 4665 4045 4695
rect 4205 4695 4245 4705
rect 4205 4665 4210 4695
rect 4240 4665 4245 4695
rect 4405 4695 4445 4705
rect 4405 4665 4410 4695
rect 4440 4665 4445 4695
rect 4605 4695 4645 4705
rect 4605 4665 4610 4695
rect 4640 4665 4645 4695
rect 4805 4695 4845 4705
rect 4805 4665 4810 4695
rect 4840 4665 4845 4695
rect 5005 4695 5045 4705
rect 5005 4665 5010 4695
rect 5040 4665 5045 4695
rect 5205 4695 5245 4705
rect 5205 4665 5210 4695
rect 5240 4665 5245 4695
rect 5405 4695 5445 4705
rect 5405 4665 5410 4695
rect 5440 4665 5445 4695
rect 5605 4695 5645 4705
rect 5605 4665 5610 4695
rect 5640 4665 5645 4695
rect 5805 4695 5845 4705
rect 5805 4665 5810 4695
rect 5840 4665 5845 4695
rect 6005 4695 6045 4705
rect 6005 4665 6010 4695
rect 6040 4665 6045 4695
rect 6205 4695 6245 4705
rect 6205 4665 6210 4695
rect 6240 4665 6245 4695
rect 6405 4695 6445 4705
rect 6405 4665 6410 4695
rect 6440 4665 6445 4695
rect -188 4580 -185 4665
rect -165 4580 -162 4665
rect 15 4580 35 4665
rect 215 4580 235 4665
rect 415 4580 435 4665
rect 615 4580 635 4665
rect 815 4580 835 4665
rect 1015 4580 1035 4665
rect 1215 4580 1235 4665
rect 1415 4580 1435 4665
rect 1615 4580 1635 4665
rect 1815 4580 1835 4665
rect 2015 4580 2035 4665
rect 2215 4580 2235 4665
rect 2415 4580 2435 4665
rect 2615 4580 2635 4665
rect 2815 4580 2835 4665
rect 3015 4580 3035 4665
rect 3215 4580 3235 4665
rect 3415 4580 3435 4665
rect 3615 4580 3635 4665
rect 3815 4580 3835 4665
rect 4015 4580 4035 4665
rect 4215 4580 4235 4665
rect 4415 4580 4435 4665
rect -195 4550 -190 4580
rect -160 4550 -155 4580
rect -195 4510 -185 4550
rect -165 4540 -155 4550
rect 5 4550 10 4580
rect 40 4550 45 4580
rect 5 4540 45 4550
rect 205 4550 210 4580
rect 240 4550 245 4580
rect 205 4540 245 4550
rect 405 4550 410 4580
rect 440 4550 445 4580
rect 405 4540 445 4550
rect 605 4550 610 4580
rect 640 4550 645 4580
rect 605 4540 645 4550
rect 805 4550 810 4580
rect 840 4550 845 4580
rect 805 4540 845 4550
rect 1005 4550 1010 4580
rect 1040 4550 1045 4580
rect 1005 4540 1045 4550
rect 1205 4550 1210 4580
rect 1240 4550 1245 4580
rect 1205 4540 1245 4550
rect 1405 4550 1410 4580
rect 1440 4550 1445 4580
rect 1405 4540 1445 4550
rect 1605 4550 1610 4580
rect 1640 4550 1645 4580
rect 1605 4540 1645 4550
rect 1805 4550 1810 4580
rect 1840 4550 1845 4580
rect 1805 4540 1845 4550
rect 2005 4550 2010 4580
rect 2040 4550 2045 4580
rect 2005 4540 2045 4550
rect 2205 4550 2210 4580
rect 2240 4550 2245 4580
rect 2205 4540 2245 4550
rect 2405 4550 2410 4580
rect 2440 4550 2445 4580
rect 2405 4540 2445 4550
rect 2605 4550 2610 4580
rect 2640 4550 2645 4580
rect 2605 4540 2645 4550
rect 2805 4550 2810 4580
rect 2840 4550 2845 4580
rect 2805 4540 2845 4550
rect 3005 4550 3010 4580
rect 3040 4550 3045 4580
rect 3005 4540 3045 4550
rect 3205 4550 3210 4580
rect 3240 4550 3245 4580
rect 3205 4540 3245 4550
rect 3405 4550 3410 4580
rect 3440 4550 3445 4580
rect 3405 4540 3445 4550
rect 3605 4550 3610 4580
rect 3640 4550 3645 4580
rect 3605 4540 3645 4550
rect 3805 4550 3810 4580
rect 3840 4550 3845 4580
rect 3805 4540 3845 4550
rect 4005 4550 4010 4580
rect 4040 4550 4045 4580
rect 4005 4540 4045 4550
rect 4205 4550 4210 4580
rect 4240 4550 4245 4580
rect 4205 4540 4245 4550
rect 4405 4550 4410 4580
rect 4440 4550 4445 4580
rect 4405 4540 4445 4550
rect 4605 4550 4610 4580
rect 4640 4550 4645 4580
rect 4605 4540 4645 4550
rect 4805 4550 4810 4580
rect 4840 4550 4845 4580
rect 4805 4540 4845 4550
rect 5005 4550 5010 4580
rect 5040 4550 5045 4580
rect 5005 4540 5045 4550
rect 5205 4550 5210 4580
rect 5240 4550 5245 4580
rect 5205 4540 5245 4550
rect 5405 4550 5410 4580
rect 5440 4550 5445 4580
rect 5405 4540 5445 4550
rect 5605 4550 5610 4580
rect 5640 4550 5645 4580
rect 5605 4540 5645 4550
rect 5805 4550 5810 4580
rect 5840 4550 5845 4580
rect 5805 4540 5845 4550
rect 6005 4550 6010 4580
rect 6040 4550 6045 4580
rect 6005 4540 6045 4550
rect 6205 4550 6210 4580
rect 6240 4550 6245 4580
rect 6205 4540 6245 4550
rect 6405 4550 6410 4580
rect 6440 4550 6445 4580
rect 6405 4540 6445 4550
rect -165 4520 -30 4540
rect 5 4520 1370 4540
rect 1405 4520 2970 4540
rect 3005 4520 3770 4540
rect 3805 4520 6695 4540
rect -165 4510 -155 4520
rect -195 4480 -190 4510
rect -160 4480 -155 4510
rect 5 4510 45 4520
rect 5 4480 10 4510
rect 40 4480 45 4510
rect 205 4510 245 4520
rect 205 4480 210 4510
rect 240 4480 245 4510
rect 405 4510 445 4520
rect 405 4480 410 4510
rect 440 4480 445 4510
rect 605 4510 645 4520
rect 605 4480 610 4510
rect 640 4480 645 4510
rect 805 4510 845 4520
rect 805 4480 810 4510
rect 840 4480 845 4510
rect 1005 4510 1045 4520
rect 1005 4480 1010 4510
rect 1040 4480 1045 4510
rect 1205 4510 1245 4520
rect 1205 4480 1210 4510
rect 1240 4480 1245 4510
rect 1405 4510 1445 4520
rect 1405 4480 1410 4510
rect 1440 4480 1445 4510
rect 1605 4510 1645 4520
rect 1605 4480 1610 4510
rect 1640 4480 1645 4510
rect 1805 4510 1845 4520
rect 1805 4480 1810 4510
rect 1840 4480 1845 4510
rect 2005 4510 2045 4520
rect 2005 4480 2010 4510
rect 2040 4480 2045 4510
rect 2205 4510 2245 4520
rect 2205 4480 2210 4510
rect 2240 4480 2245 4510
rect 2405 4510 2445 4520
rect 2405 4480 2410 4510
rect 2440 4480 2445 4510
rect 2605 4510 2645 4520
rect 2605 4480 2610 4510
rect 2640 4480 2645 4510
rect 2805 4510 2845 4520
rect 2805 4480 2810 4510
rect 2840 4480 2845 4510
rect 3005 4510 3045 4520
rect 3005 4480 3010 4510
rect 3040 4480 3045 4510
rect 3205 4510 3245 4520
rect 3205 4480 3210 4510
rect 3240 4480 3245 4510
rect 3405 4510 3445 4520
rect 3405 4480 3410 4510
rect 3440 4480 3445 4510
rect 3605 4510 3645 4520
rect 3605 4480 3610 4510
rect 3640 4480 3645 4510
rect 3805 4510 3845 4520
rect 3805 4480 3810 4510
rect 3840 4480 3845 4510
rect 4005 4510 4045 4520
rect 4005 4480 4010 4510
rect 4040 4480 4045 4510
rect 4205 4510 4245 4520
rect 4205 4480 4210 4510
rect 4240 4480 4245 4510
rect 4405 4510 4445 4520
rect 4405 4480 4410 4510
rect 4440 4480 4445 4510
rect 4605 4510 4645 4520
rect 4605 4480 4610 4510
rect 4640 4480 4645 4510
rect 4805 4510 4845 4520
rect 4805 4480 4810 4510
rect 4840 4480 4845 4510
rect 5005 4510 5045 4520
rect 5005 4480 5010 4510
rect 5040 4480 5045 4510
rect 5205 4510 5245 4520
rect 5205 4480 5210 4510
rect 5240 4480 5245 4510
rect 5405 4510 5445 4520
rect 5405 4480 5410 4510
rect 5440 4480 5445 4510
rect 5605 4510 5645 4520
rect 5605 4480 5610 4510
rect 5640 4480 5645 4510
rect 5805 4510 5845 4520
rect 5805 4480 5810 4510
rect 5840 4480 5845 4510
rect 6005 4510 6045 4520
rect 6005 4480 6010 4510
rect 6040 4480 6045 4510
rect 6205 4510 6245 4520
rect 6205 4480 6210 4510
rect 6240 4480 6245 4510
rect 6405 4510 6445 4520
rect 6405 4480 6410 4510
rect 6440 4480 6445 4510
rect -188 4395 -185 4480
rect -165 4395 -162 4480
rect 15 4395 35 4480
rect 215 4395 235 4480
rect 415 4395 435 4480
rect 615 4395 635 4480
rect 815 4395 835 4480
rect 1015 4395 1035 4480
rect 1215 4395 1235 4480
rect 1615 4395 1635 4480
rect 1815 4395 1835 4480
rect 2015 4395 2035 4480
rect 2215 4395 2235 4480
rect 2415 4395 2435 4480
rect 2615 4395 2635 4480
rect 2815 4395 2835 4480
rect 3015 4395 3035 4480
rect 3215 4395 3235 4480
rect 3415 4395 3435 4480
rect 3615 4395 3635 4480
rect 4015 4395 4035 4480
rect 4215 4395 4235 4480
rect 4415 4395 4435 4480
rect 4615 4395 4635 4480
rect 4815 4395 4835 4480
rect 5015 4395 5035 4480
rect 5215 4395 5235 4480
rect 5415 4395 5435 4480
rect 5615 4395 5635 4480
rect 5815 4395 5835 4480
rect 6015 4395 6035 4480
rect 6215 4395 6235 4480
rect -195 4365 -190 4395
rect -160 4365 -155 4395
rect -195 4325 -185 4365
rect -165 4355 -155 4365
rect 5 4365 10 4395
rect 40 4365 45 4395
rect 5 4355 45 4365
rect 205 4365 210 4395
rect 240 4365 245 4395
rect 205 4355 245 4365
rect 405 4365 410 4395
rect 440 4365 445 4395
rect 405 4355 445 4365
rect 605 4365 610 4395
rect 640 4365 645 4395
rect 605 4355 645 4365
rect 805 4365 810 4395
rect 840 4365 845 4395
rect 805 4355 845 4365
rect 1005 4365 1010 4395
rect 1040 4365 1045 4395
rect 1005 4355 1045 4365
rect 1205 4365 1210 4395
rect 1240 4365 1245 4395
rect 1205 4355 1245 4365
rect 1405 4365 1410 4395
rect 1440 4365 1445 4395
rect 1405 4355 1445 4365
rect 1605 4365 1610 4395
rect 1640 4365 1645 4395
rect 1605 4355 1645 4365
rect 1805 4365 1810 4395
rect 1840 4365 1845 4395
rect 1805 4355 1845 4365
rect 2005 4365 2010 4395
rect 2040 4365 2045 4395
rect 2005 4355 2045 4365
rect 2205 4365 2210 4395
rect 2240 4365 2245 4395
rect 2205 4355 2245 4365
rect 2405 4365 2410 4395
rect 2440 4365 2445 4395
rect 2405 4355 2445 4365
rect 2605 4365 2610 4395
rect 2640 4365 2645 4395
rect 2605 4355 2645 4365
rect 2805 4365 2810 4395
rect 2840 4365 2845 4395
rect 2805 4355 2845 4365
rect 3005 4365 3010 4395
rect 3040 4365 3045 4395
rect 3005 4355 3045 4365
rect 3205 4365 3210 4395
rect 3240 4365 3245 4395
rect 3205 4355 3245 4365
rect 3405 4365 3410 4395
rect 3440 4365 3445 4395
rect 3405 4355 3445 4365
rect 3605 4365 3610 4395
rect 3640 4365 3645 4395
rect 3605 4355 3645 4365
rect 3805 4365 3810 4395
rect 3840 4365 3845 4395
rect 3805 4355 3845 4365
rect 4005 4365 4010 4395
rect 4040 4365 4045 4395
rect 4005 4355 4045 4365
rect 4205 4365 4210 4395
rect 4240 4365 4245 4395
rect 4205 4355 4245 4365
rect 4405 4365 4410 4395
rect 4440 4365 4445 4395
rect 4405 4355 4445 4365
rect 4605 4365 4610 4395
rect 4640 4365 4645 4395
rect 4605 4355 4645 4365
rect 4805 4365 4810 4395
rect 4840 4365 4845 4395
rect 4805 4355 4845 4365
rect 5005 4365 5010 4395
rect 5040 4365 5045 4395
rect 5005 4355 5045 4365
rect 5205 4365 5210 4395
rect 5240 4365 5245 4395
rect 5205 4355 5245 4365
rect 5405 4365 5410 4395
rect 5440 4365 5445 4395
rect 5405 4355 5445 4365
rect 5605 4365 5610 4395
rect 5640 4365 5645 4395
rect 5605 4355 5645 4365
rect 5805 4365 5810 4395
rect 5840 4365 5845 4395
rect 5805 4355 5845 4365
rect 6005 4365 6010 4395
rect 6040 4365 6045 4395
rect 6005 4355 6045 4365
rect 6205 4365 6210 4395
rect 6240 4365 6245 4395
rect 6205 4355 6245 4365
rect 6405 4365 6410 4395
rect 6440 4365 6445 4395
rect 6405 4355 6445 4365
rect -165 4335 -30 4355
rect 5 4335 1570 4355
rect 1605 4335 2970 4355
rect 3005 4335 3970 4355
rect 4005 4335 6570 4355
rect -165 4325 -155 4335
rect -195 4295 -190 4325
rect -160 4295 -155 4325
rect 5 4325 45 4335
rect 5 4295 10 4325
rect 40 4295 45 4325
rect 205 4325 245 4335
rect 205 4295 210 4325
rect 240 4295 245 4325
rect 405 4325 445 4335
rect 405 4295 410 4325
rect 440 4295 445 4325
rect 605 4325 645 4335
rect 605 4295 610 4325
rect 640 4295 645 4325
rect 805 4325 845 4335
rect 805 4295 810 4325
rect 840 4295 845 4325
rect 1005 4325 1045 4335
rect 1005 4295 1010 4325
rect 1040 4295 1045 4325
rect 1205 4325 1245 4335
rect 1205 4295 1210 4325
rect 1240 4295 1245 4325
rect 1405 4325 1445 4335
rect 1405 4295 1410 4325
rect 1440 4295 1445 4325
rect 1605 4325 1645 4335
rect 1605 4295 1610 4325
rect 1640 4295 1645 4325
rect 1805 4325 1845 4335
rect 1805 4295 1810 4325
rect 1840 4295 1845 4325
rect 2005 4325 2045 4335
rect 2005 4295 2010 4325
rect 2040 4295 2045 4325
rect 2205 4325 2245 4335
rect 2205 4295 2210 4325
rect 2240 4295 2245 4325
rect 2405 4325 2445 4335
rect 2405 4295 2410 4325
rect 2440 4295 2445 4325
rect 2605 4325 2645 4335
rect 2605 4295 2610 4325
rect 2640 4295 2645 4325
rect 2805 4325 2845 4335
rect 2805 4295 2810 4325
rect 2840 4295 2845 4325
rect 3005 4325 3045 4335
rect 3005 4295 3010 4325
rect 3040 4295 3045 4325
rect 3205 4325 3245 4335
rect 3205 4295 3210 4325
rect 3240 4295 3245 4325
rect 3405 4325 3445 4335
rect 3405 4295 3410 4325
rect 3440 4295 3445 4325
rect 3605 4325 3645 4335
rect 3605 4295 3610 4325
rect 3640 4295 3645 4325
rect 3805 4325 3845 4335
rect 3805 4295 3810 4325
rect 3840 4295 3845 4325
rect 4005 4325 4045 4335
rect 4005 4295 4010 4325
rect 4040 4295 4045 4325
rect 4205 4325 4245 4335
rect 4205 4295 4210 4325
rect 4240 4295 4245 4325
rect 4405 4325 4445 4335
rect 4405 4295 4410 4325
rect 4440 4295 4445 4325
rect 4605 4325 4645 4335
rect 4605 4295 4610 4325
rect 4640 4295 4645 4325
rect 4805 4325 4845 4335
rect 4805 4295 4810 4325
rect 4840 4295 4845 4325
rect 5005 4325 5045 4335
rect 5005 4295 5010 4325
rect 5040 4295 5045 4325
rect 5205 4325 5245 4335
rect 5205 4295 5210 4325
rect 5240 4295 5245 4325
rect 5405 4325 5445 4335
rect 5405 4295 5410 4325
rect 5440 4295 5445 4325
rect 5605 4325 5645 4335
rect 5605 4295 5610 4325
rect 5640 4295 5645 4325
rect 5805 4325 5845 4335
rect 5805 4295 5810 4325
rect 5840 4295 5845 4325
rect 6005 4325 6045 4335
rect 6005 4295 6010 4325
rect 6040 4295 6045 4325
rect 6205 4325 6245 4335
rect 6205 4295 6210 4325
rect 6240 4295 6245 4325
rect 6405 4325 6445 4335
rect 6405 4295 6410 4325
rect 6440 4295 6445 4325
rect -188 4210 -185 4295
rect -165 4210 -162 4295
rect 15 4210 35 4295
rect 215 4210 235 4295
rect 415 4210 435 4295
rect 615 4210 635 4295
rect 815 4210 835 4295
rect 1015 4210 1035 4295
rect 1215 4210 1235 4295
rect 1415 4210 1435 4295
rect 1615 4210 1635 4295
rect 1815 4210 1835 4295
rect 2015 4210 2035 4295
rect 2215 4210 2235 4295
rect 2415 4210 2435 4295
rect 2615 4210 2635 4295
rect 2815 4210 2835 4295
rect 3015 4210 3035 4295
rect 3215 4210 3235 4295
rect 3415 4210 3435 4295
rect 3615 4210 3635 4295
rect 3815 4210 3835 4295
rect 4015 4210 4035 4295
rect 4215 4210 4235 4295
rect 4415 4210 4435 4295
rect 4615 4210 4635 4295
rect 4815 4210 4835 4295
rect 5015 4210 5035 4295
rect 5215 4210 5235 4295
rect 5415 4210 5435 4295
rect 5615 4210 5635 4295
rect 5815 4210 5835 4295
rect 6015 4210 6035 4295
rect 6215 4210 6235 4295
rect -195 4180 -190 4210
rect -160 4180 -155 4210
rect -195 4140 -185 4180
rect -165 4170 -155 4180
rect 5 4180 10 4210
rect 40 4180 45 4210
rect 5 4170 45 4180
rect 205 4180 210 4210
rect 240 4180 245 4210
rect 205 4170 245 4180
rect 405 4180 410 4210
rect 440 4180 445 4210
rect 405 4170 445 4180
rect 605 4180 610 4210
rect 640 4180 645 4210
rect 605 4170 645 4180
rect 805 4180 810 4210
rect 840 4180 845 4210
rect 805 4170 845 4180
rect 1005 4180 1010 4210
rect 1040 4180 1045 4210
rect 1005 4170 1045 4180
rect 1205 4180 1210 4210
rect 1240 4180 1245 4210
rect 1205 4170 1245 4180
rect 1405 4180 1410 4210
rect 1440 4180 1445 4210
rect 1405 4170 1445 4180
rect 1605 4180 1610 4210
rect 1640 4180 1645 4210
rect 1605 4170 1645 4180
rect 1805 4180 1810 4210
rect 1840 4180 1845 4210
rect 1805 4170 1845 4180
rect 2005 4180 2010 4210
rect 2040 4180 2045 4210
rect 2005 4170 2045 4180
rect 2205 4180 2210 4210
rect 2240 4180 2245 4210
rect 2205 4170 2245 4180
rect 2405 4180 2410 4210
rect 2440 4180 2445 4210
rect 2405 4170 2445 4180
rect 2605 4180 2610 4210
rect 2640 4180 2645 4210
rect 2605 4170 2645 4180
rect 2805 4180 2810 4210
rect 2840 4180 2845 4210
rect 2805 4170 2845 4180
rect 3005 4180 3010 4210
rect 3040 4180 3045 4210
rect 3005 4170 3045 4180
rect 3205 4180 3210 4210
rect 3240 4180 3245 4210
rect 3205 4170 3245 4180
rect 3405 4180 3410 4210
rect 3440 4180 3445 4210
rect 3405 4170 3445 4180
rect 3605 4180 3610 4210
rect 3640 4180 3645 4210
rect 3605 4170 3645 4180
rect 3805 4180 3810 4210
rect 3840 4180 3845 4210
rect 3805 4170 3845 4180
rect 4005 4180 4010 4210
rect 4040 4180 4045 4210
rect 4005 4170 4045 4180
rect 4205 4180 4210 4210
rect 4240 4180 4245 4210
rect 4205 4170 4245 4180
rect 4405 4180 4410 4210
rect 4440 4180 4445 4210
rect 4405 4170 4445 4180
rect 4605 4180 4610 4210
rect 4640 4180 4645 4210
rect 4605 4170 4645 4180
rect 4805 4180 4810 4210
rect 4840 4180 4845 4210
rect 4805 4170 4845 4180
rect 5005 4180 5010 4210
rect 5040 4180 5045 4210
rect 5005 4170 5045 4180
rect 5205 4180 5210 4210
rect 5240 4180 5245 4210
rect 5205 4170 5245 4180
rect 5405 4180 5410 4210
rect 5440 4180 5445 4210
rect 5405 4170 5445 4180
rect 5605 4180 5610 4210
rect 5640 4180 5645 4210
rect 5605 4170 5645 4180
rect 5805 4180 5810 4210
rect 5840 4180 5845 4210
rect 5805 4170 5845 4180
rect 6005 4180 6010 4210
rect 6040 4180 6045 4210
rect 6005 4170 6045 4180
rect 6205 4180 6210 4210
rect 6240 4180 6245 4210
rect 6205 4170 6245 4180
rect 6405 4180 6410 4210
rect 6440 4180 6445 4210
rect 6405 4170 6445 4180
rect -165 4150 -30 4170
rect 5 4150 1570 4170
rect 1605 4150 2970 4170
rect 3005 4150 3970 4170
rect 4005 4150 6570 4170
rect -165 4140 -155 4150
rect -195 4110 -190 4140
rect -160 4110 -155 4140
rect 5 4140 45 4150
rect 5 4110 10 4140
rect 40 4110 45 4140
rect 205 4140 245 4150
rect 205 4110 210 4140
rect 240 4110 245 4140
rect 405 4140 445 4150
rect 405 4110 410 4140
rect 440 4110 445 4140
rect 605 4140 645 4150
rect 605 4110 610 4140
rect 640 4110 645 4140
rect 805 4140 845 4150
rect 805 4110 810 4140
rect 840 4110 845 4140
rect 1005 4140 1045 4150
rect 1005 4110 1010 4140
rect 1040 4110 1045 4140
rect 1205 4140 1245 4150
rect 1205 4110 1210 4140
rect 1240 4110 1245 4140
rect 1405 4140 1445 4150
rect 1405 4110 1410 4140
rect 1440 4110 1445 4140
rect 1605 4140 1645 4150
rect 1605 4110 1610 4140
rect 1640 4110 1645 4140
rect 1805 4140 1845 4150
rect 1805 4110 1810 4140
rect 1840 4110 1845 4140
rect 2005 4140 2045 4150
rect 2005 4110 2010 4140
rect 2040 4110 2045 4140
rect 2205 4140 2245 4150
rect 2205 4110 2210 4140
rect 2240 4110 2245 4140
rect 2405 4140 2445 4150
rect 2405 4110 2410 4140
rect 2440 4110 2445 4140
rect 2605 4140 2645 4150
rect 2605 4110 2610 4140
rect 2640 4110 2645 4140
rect 2805 4140 2845 4150
rect 2805 4110 2810 4140
rect 2840 4110 2845 4140
rect 3005 4140 3045 4150
rect 3005 4110 3010 4140
rect 3040 4110 3045 4140
rect 3205 4140 3245 4150
rect 3205 4110 3210 4140
rect 3240 4110 3245 4140
rect 3405 4140 3445 4150
rect 3405 4110 3410 4140
rect 3440 4110 3445 4140
rect 3605 4140 3645 4150
rect 3605 4110 3610 4140
rect 3640 4110 3645 4140
rect 3805 4140 3845 4150
rect 3805 4110 3810 4140
rect 3840 4110 3845 4140
rect 4005 4140 4045 4150
rect 4005 4110 4010 4140
rect 4040 4110 4045 4140
rect 4205 4140 4245 4150
rect 4205 4110 4210 4140
rect 4240 4110 4245 4140
rect 4405 4140 4445 4150
rect 4405 4110 4410 4140
rect 4440 4110 4445 4140
rect 4605 4140 4645 4150
rect 4605 4110 4610 4140
rect 4640 4110 4645 4140
rect 4805 4140 4845 4150
rect 4805 4110 4810 4140
rect 4840 4110 4845 4140
rect 5005 4140 5045 4150
rect 5005 4110 5010 4140
rect 5040 4110 5045 4140
rect 5205 4140 5245 4150
rect 5205 4110 5210 4140
rect 5240 4110 5245 4140
rect 5405 4140 5445 4150
rect 5405 4110 5410 4140
rect 5440 4110 5445 4140
rect 5605 4140 5645 4150
rect 5605 4110 5610 4140
rect 5640 4110 5645 4140
rect 5805 4140 5845 4150
rect 5805 4110 5810 4140
rect 5840 4110 5845 4140
rect 6005 4140 6045 4150
rect 6005 4110 6010 4140
rect 6040 4110 6045 4140
rect 6205 4140 6245 4150
rect 6205 4110 6210 4140
rect 6240 4110 6245 4140
rect 6405 4140 6445 4150
rect 6405 4110 6410 4140
rect 6440 4110 6445 4140
rect -188 4025 -185 4110
rect -165 4025 -162 4110
rect 15 4025 35 4110
rect 215 4025 235 4110
rect 415 4025 435 4110
rect 615 4025 635 4110
rect 815 4025 835 4110
rect 1015 4025 1035 4110
rect 1215 4025 1235 4110
rect 1415 4025 1435 4110
rect 1615 4025 1635 4110
rect 1815 4025 1835 4110
rect 2015 4025 2035 4110
rect 2215 4025 2235 4110
rect 2415 4025 2435 4110
rect 2615 4025 2635 4110
rect 2815 4025 2835 4110
rect 3015 4025 3035 4110
rect 3215 4025 3235 4110
rect 3415 4025 3435 4110
rect 3615 4025 3635 4110
rect 3815 4025 3835 4110
rect -195 3995 -190 4025
rect -160 3995 -155 4025
rect -195 3955 -185 3995
rect -165 3985 -155 3995
rect 5 3995 10 4025
rect 40 3995 45 4025
rect 5 3985 45 3995
rect 205 3995 210 4025
rect 240 3995 245 4025
rect 205 3985 245 3995
rect 405 3995 410 4025
rect 440 3995 445 4025
rect 405 3985 445 3995
rect 605 3995 610 4025
rect 640 3995 645 4025
rect 605 3985 645 3995
rect 805 3995 810 4025
rect 840 3995 845 4025
rect 805 3985 845 3995
rect 1005 3995 1010 4025
rect 1040 3995 1045 4025
rect 1005 3985 1045 3995
rect 1205 3995 1210 4025
rect 1240 3995 1245 4025
rect 1205 3985 1245 3995
rect 1405 3995 1410 4025
rect 1440 3995 1445 4025
rect 1405 3985 1445 3995
rect 1605 3995 1610 4025
rect 1640 3995 1645 4025
rect 1605 3985 1645 3995
rect 1805 3995 1810 4025
rect 1840 3995 1845 4025
rect 1805 3985 1845 3995
rect 2005 3995 2010 4025
rect 2040 3995 2045 4025
rect 2005 3985 2045 3995
rect 2205 3995 2210 4025
rect 2240 3995 2245 4025
rect 2205 3985 2245 3995
rect 2405 3995 2410 4025
rect 2440 3995 2445 4025
rect 2405 3985 2445 3995
rect 2605 3995 2610 4025
rect 2640 3995 2645 4025
rect 2605 3985 2645 3995
rect 2805 3995 2810 4025
rect 2840 3995 2845 4025
rect 2805 3985 2845 3995
rect 3005 3995 3010 4025
rect 3040 3995 3045 4025
rect 3005 3985 3045 3995
rect 3205 3995 3210 4025
rect 3240 3995 3245 4025
rect 3205 3985 3245 3995
rect 3405 3995 3410 4025
rect 3440 3995 3445 4025
rect 3405 3985 3445 3995
rect 3605 3995 3610 4025
rect 3640 3995 3645 4025
rect 3605 3985 3645 3995
rect 3805 3995 3810 4025
rect 3840 3995 3845 4025
rect 3805 3985 3845 3995
rect 4005 3995 4010 4025
rect 4040 3995 4045 4025
rect 4005 3985 4045 3995
rect 4205 3995 4210 4025
rect 4240 3995 4245 4025
rect 4205 3985 4245 3995
rect 4405 3995 4410 4025
rect 4440 3995 4445 4025
rect 4405 3985 4445 3995
rect 4605 3995 4610 4025
rect 4640 3995 4645 4025
rect 4605 3985 4645 3995
rect 4805 3995 4810 4025
rect 4840 3995 4845 4025
rect 4805 3985 4845 3995
rect 5005 3995 5010 4025
rect 5040 3995 5045 4025
rect 5005 3985 5045 3995
rect 5205 3995 5210 4025
rect 5240 3995 5245 4025
rect 5205 3985 5245 3995
rect 5405 3995 5410 4025
rect 5440 3995 5445 4025
rect 5405 3985 5445 3995
rect 5605 3995 5610 4025
rect 5640 3995 5645 4025
rect 5605 3985 5645 3995
rect 5805 3995 5810 4025
rect 5840 3995 5845 4025
rect 5805 3985 5845 3995
rect 6005 3995 6010 4025
rect 6040 3995 6045 4025
rect 6005 3985 6045 3995
rect 6205 3995 6210 4025
rect 6240 3995 6245 4025
rect 6205 3985 6245 3995
rect 6405 3995 6410 4025
rect 6440 3995 6445 4025
rect 6405 3985 6445 3995
rect -165 3965 -30 3985
rect 5 3965 1570 3985
rect 1605 3965 2970 3985
rect 3005 3965 6695 3985
rect -165 3955 -155 3965
rect -195 3925 -190 3955
rect -160 3925 -155 3955
rect 5 3955 45 3965
rect 5 3925 10 3955
rect 40 3925 45 3955
rect 205 3955 245 3965
rect 205 3925 210 3955
rect 240 3925 245 3955
rect 405 3955 445 3965
rect 405 3925 410 3955
rect 440 3925 445 3955
rect 605 3955 645 3965
rect 605 3925 610 3955
rect 640 3925 645 3955
rect 805 3955 845 3965
rect 805 3925 810 3955
rect 840 3925 845 3955
rect 1005 3955 1045 3965
rect 1005 3925 1010 3955
rect 1040 3925 1045 3955
rect 1205 3955 1245 3965
rect 1205 3925 1210 3955
rect 1240 3925 1245 3955
rect 1405 3955 1445 3965
rect 1405 3925 1410 3955
rect 1440 3925 1445 3955
rect 1605 3955 1645 3965
rect 1605 3925 1610 3955
rect 1640 3925 1645 3955
rect 1805 3955 1845 3965
rect 1805 3925 1810 3955
rect 1840 3925 1845 3955
rect 2005 3955 2045 3965
rect 2005 3925 2010 3955
rect 2040 3925 2045 3955
rect 2205 3955 2245 3965
rect 2205 3925 2210 3955
rect 2240 3925 2245 3955
rect 2405 3955 2445 3965
rect 2405 3925 2410 3955
rect 2440 3925 2445 3955
rect 2605 3955 2645 3965
rect 2605 3925 2610 3955
rect 2640 3925 2645 3955
rect 2805 3955 2845 3965
rect 2805 3925 2810 3955
rect 2840 3925 2845 3955
rect 3005 3955 3045 3965
rect 3005 3925 3010 3955
rect 3040 3925 3045 3955
rect 3205 3955 3245 3965
rect 3205 3925 3210 3955
rect 3240 3925 3245 3955
rect 3405 3955 3445 3965
rect 3405 3925 3410 3955
rect 3440 3925 3445 3955
rect 3605 3955 3645 3965
rect 3605 3925 3610 3955
rect 3640 3925 3645 3955
rect 3805 3955 3845 3965
rect 3805 3925 3810 3955
rect 3840 3925 3845 3955
rect 4005 3955 4045 3965
rect 4005 3925 4010 3955
rect 4040 3925 4045 3955
rect 4205 3955 4245 3965
rect 4205 3925 4210 3955
rect 4240 3925 4245 3955
rect 4405 3955 4445 3965
rect 4405 3925 4410 3955
rect 4440 3925 4445 3955
rect 4605 3955 4645 3965
rect 4605 3925 4610 3955
rect 4640 3925 4645 3955
rect 4805 3955 4845 3965
rect 4805 3925 4810 3955
rect 4840 3925 4845 3955
rect 5005 3955 5045 3965
rect 5005 3925 5010 3955
rect 5040 3925 5045 3955
rect 5205 3955 5245 3965
rect 5205 3925 5210 3955
rect 5240 3925 5245 3955
rect 5405 3955 5445 3965
rect 5405 3925 5410 3955
rect 5440 3925 5445 3955
rect 5605 3955 5645 3965
rect 5605 3925 5610 3955
rect 5640 3925 5645 3955
rect 5805 3955 5845 3965
rect 5805 3925 5810 3955
rect 5840 3925 5845 3955
rect 6005 3955 6045 3965
rect 6005 3925 6010 3955
rect 6040 3925 6045 3955
rect 6205 3955 6245 3965
rect 6205 3925 6210 3955
rect 6240 3925 6245 3955
rect 6405 3955 6445 3965
rect 6405 3925 6410 3955
rect 6440 3925 6445 3955
rect -188 3840 -185 3925
rect -165 3840 -162 3925
rect 15 3840 35 3925
rect 215 3840 235 3925
rect 415 3840 435 3925
rect 615 3840 635 3925
rect 815 3840 835 3925
rect 1015 3840 1035 3925
rect 1215 3840 1235 3925
rect 1415 3840 1435 3925
rect 1615 3840 1635 3925
rect 1815 3840 1835 3925
rect 2015 3840 2035 3925
rect 2215 3840 2235 3925
rect 2415 3840 2435 3925
rect 2615 3840 2635 3925
rect 2815 3840 2835 3925
rect 3015 3840 3035 3925
rect 3215 3840 3235 3925
rect 3415 3840 3435 3925
rect 3615 3840 3635 3925
rect 3815 3840 3835 3925
rect 4015 3840 4035 3925
rect 4215 3840 4235 3925
rect 4415 3840 4435 3925
rect 4615 3840 4635 3925
rect 4815 3840 4835 3925
rect 5015 3840 5035 3925
rect 5215 3840 5235 3925
rect 5415 3840 5435 3925
rect 5615 3840 5635 3925
rect 5815 3840 5835 3925
rect 6015 3840 6035 3925
rect 6215 3840 6235 3925
rect -195 3810 -190 3840
rect -160 3810 -155 3840
rect -195 3770 -185 3810
rect -165 3800 -155 3810
rect 5 3810 10 3840
rect 40 3810 45 3840
rect 5 3800 45 3810
rect 205 3810 210 3840
rect 240 3810 245 3840
rect 205 3800 245 3810
rect 405 3810 410 3840
rect 440 3810 445 3840
rect 405 3800 445 3810
rect 605 3810 610 3840
rect 640 3810 645 3840
rect 605 3800 645 3810
rect 805 3810 810 3840
rect 840 3810 845 3840
rect 805 3800 845 3810
rect 1005 3810 1010 3840
rect 1040 3810 1045 3840
rect 1005 3800 1045 3810
rect 1205 3810 1210 3840
rect 1240 3810 1245 3840
rect 1205 3800 1245 3810
rect 1405 3810 1410 3840
rect 1440 3810 1445 3840
rect 1405 3800 1445 3810
rect 1605 3810 1610 3840
rect 1640 3810 1645 3840
rect 1605 3800 1645 3810
rect 1805 3810 1810 3840
rect 1840 3810 1845 3840
rect 1805 3800 1845 3810
rect 2005 3810 2010 3840
rect 2040 3810 2045 3840
rect 2005 3800 2045 3810
rect 2205 3810 2210 3840
rect 2240 3810 2245 3840
rect 2205 3800 2245 3810
rect 2405 3810 2410 3840
rect 2440 3810 2445 3840
rect 2405 3800 2445 3810
rect 2605 3810 2610 3840
rect 2640 3810 2645 3840
rect 2605 3800 2645 3810
rect 2805 3810 2810 3840
rect 2840 3810 2845 3840
rect 2805 3800 2845 3810
rect 3005 3810 3010 3840
rect 3040 3810 3045 3840
rect 3005 3800 3045 3810
rect 3205 3810 3210 3840
rect 3240 3810 3245 3840
rect 3205 3800 3245 3810
rect 3405 3810 3410 3840
rect 3440 3810 3445 3840
rect 3405 3800 3445 3810
rect 3605 3810 3610 3840
rect 3640 3810 3645 3840
rect 3605 3800 3645 3810
rect 3805 3810 3810 3840
rect 3840 3810 3845 3840
rect 3805 3800 3845 3810
rect 4005 3810 4010 3840
rect 4040 3810 4045 3840
rect 4005 3800 4045 3810
rect 4205 3810 4210 3840
rect 4240 3810 4245 3840
rect 4205 3800 4245 3810
rect 4405 3810 4410 3840
rect 4440 3810 4445 3840
rect 4405 3800 4445 3810
rect 4605 3810 4610 3840
rect 4640 3810 4645 3840
rect 4605 3800 4645 3810
rect 4805 3810 4810 3840
rect 4840 3810 4845 3840
rect 4805 3800 4845 3810
rect 5005 3810 5010 3840
rect 5040 3810 5045 3840
rect 5005 3800 5045 3810
rect 5205 3810 5210 3840
rect 5240 3810 5245 3840
rect 5205 3800 5245 3810
rect 5405 3810 5410 3840
rect 5440 3810 5445 3840
rect 5405 3800 5445 3810
rect 5605 3810 5610 3840
rect 5640 3810 5645 3840
rect 5605 3800 5645 3810
rect 5805 3810 5810 3840
rect 5840 3810 5845 3840
rect 5805 3800 5845 3810
rect 6005 3810 6010 3840
rect 6040 3810 6045 3840
rect 6005 3800 6045 3810
rect 6205 3810 6210 3840
rect 6240 3810 6245 3840
rect 6205 3800 6245 3810
rect 6405 3810 6410 3840
rect 6440 3810 6445 3840
rect 6405 3800 6445 3810
rect -165 3780 -30 3800
rect 5 3780 1570 3800
rect 1605 3780 2970 3800
rect 3005 3780 6570 3800
rect -165 3770 -155 3780
rect -195 3740 -190 3770
rect -160 3740 -155 3770
rect 5 3770 45 3780
rect 5 3740 10 3770
rect 40 3740 45 3770
rect 205 3770 245 3780
rect 205 3740 210 3770
rect 240 3740 245 3770
rect 405 3770 445 3780
rect 405 3740 410 3770
rect 440 3740 445 3770
rect 605 3770 645 3780
rect 605 3740 610 3770
rect 640 3740 645 3770
rect 805 3770 845 3780
rect 805 3740 810 3770
rect 840 3740 845 3770
rect 1005 3770 1045 3780
rect 1005 3740 1010 3770
rect 1040 3740 1045 3770
rect 1205 3770 1245 3780
rect 1205 3740 1210 3770
rect 1240 3740 1245 3770
rect 1405 3770 1445 3780
rect 1405 3740 1410 3770
rect 1440 3740 1445 3770
rect 1605 3770 1645 3780
rect 1605 3740 1610 3770
rect 1640 3740 1645 3770
rect 1805 3770 1845 3780
rect 1805 3740 1810 3770
rect 1840 3740 1845 3770
rect 2005 3770 2045 3780
rect 2005 3740 2010 3770
rect 2040 3740 2045 3770
rect 2205 3770 2245 3780
rect 2205 3740 2210 3770
rect 2240 3740 2245 3770
rect 2405 3770 2445 3780
rect 2405 3740 2410 3770
rect 2440 3740 2445 3770
rect 2605 3770 2645 3780
rect 2605 3740 2610 3770
rect 2640 3740 2645 3770
rect 2805 3770 2845 3780
rect 2805 3740 2810 3770
rect 2840 3740 2845 3770
rect 3005 3770 3045 3780
rect 3005 3740 3010 3770
rect 3040 3740 3045 3770
rect 3205 3770 3245 3780
rect 3205 3740 3210 3770
rect 3240 3740 3245 3770
rect 3405 3770 3445 3780
rect 3405 3740 3410 3770
rect 3440 3740 3445 3770
rect 3605 3770 3645 3780
rect 3605 3740 3610 3770
rect 3640 3740 3645 3770
rect 3805 3770 3845 3780
rect 3805 3740 3810 3770
rect 3840 3740 3845 3770
rect 4005 3770 4045 3780
rect 4005 3740 4010 3770
rect 4040 3740 4045 3770
rect 4205 3770 4245 3780
rect 4205 3740 4210 3770
rect 4240 3740 4245 3770
rect 4405 3770 4445 3780
rect 4405 3740 4410 3770
rect 4440 3740 4445 3770
rect 4605 3770 4645 3780
rect 4605 3740 4610 3770
rect 4640 3740 4645 3770
rect 4805 3770 4845 3780
rect 4805 3740 4810 3770
rect 4840 3740 4845 3770
rect 5005 3770 5045 3780
rect 5005 3740 5010 3770
rect 5040 3740 5045 3770
rect 5205 3770 5245 3780
rect 5205 3740 5210 3770
rect 5240 3740 5245 3770
rect 5405 3770 5445 3780
rect 5405 3740 5410 3770
rect 5440 3740 5445 3770
rect 5605 3770 5645 3780
rect 5605 3740 5610 3770
rect 5640 3740 5645 3770
rect 5805 3770 5845 3780
rect 5805 3740 5810 3770
rect 5840 3740 5845 3770
rect 6005 3770 6045 3780
rect 6005 3740 6010 3770
rect 6040 3740 6045 3770
rect 6205 3770 6245 3780
rect 6205 3740 6210 3770
rect 6240 3740 6245 3770
rect 6405 3770 6445 3780
rect 6405 3740 6410 3770
rect 6440 3740 6445 3770
rect -188 3655 -185 3740
rect -165 3655 -162 3740
rect 15 3655 35 3740
rect 215 3655 235 3740
rect 415 3655 435 3740
rect 615 3655 635 3740
rect 815 3655 835 3740
rect 1015 3655 1035 3740
rect 1215 3655 1235 3740
rect 1415 3655 1435 3740
rect 1615 3655 1635 3740
rect 1815 3655 1835 3740
rect 2015 3655 2035 3740
rect 2215 3655 2235 3740
rect 2415 3655 2435 3740
rect 2615 3655 2635 3740
rect 2815 3655 2835 3740
rect 3015 3655 3035 3740
rect 3215 3655 3235 3740
rect 3415 3655 3435 3740
rect 3615 3655 3635 3740
rect 3815 3655 3835 3740
rect 4015 3655 4035 3740
rect 4215 3655 4235 3740
rect 4415 3655 4435 3740
rect 4615 3655 4635 3740
rect 4815 3655 4835 3740
rect 5015 3655 5035 3740
rect 5215 3655 5235 3740
rect 5415 3655 5435 3740
rect 5615 3655 5635 3740
rect 5815 3655 5835 3740
rect 6015 3655 6035 3740
rect 6215 3655 6235 3740
rect -195 3625 -190 3655
rect -160 3625 -155 3655
rect -195 3585 -185 3625
rect -165 3615 -155 3625
rect 5 3625 10 3655
rect 40 3625 45 3655
rect 5 3615 45 3625
rect 205 3625 210 3655
rect 240 3625 245 3655
rect 205 3615 245 3625
rect 405 3625 410 3655
rect 440 3625 445 3655
rect 405 3615 445 3625
rect 605 3625 610 3655
rect 640 3625 645 3655
rect 605 3615 645 3625
rect 805 3625 810 3655
rect 840 3625 845 3655
rect 805 3615 845 3625
rect 1005 3625 1010 3655
rect 1040 3625 1045 3655
rect 1005 3615 1045 3625
rect 1205 3625 1210 3655
rect 1240 3625 1245 3655
rect 1205 3615 1245 3625
rect 1405 3625 1410 3655
rect 1440 3625 1445 3655
rect 1405 3615 1445 3625
rect 1605 3625 1610 3655
rect 1640 3625 1645 3655
rect 1605 3615 1645 3625
rect 1805 3625 1810 3655
rect 1840 3625 1845 3655
rect 1805 3615 1845 3625
rect 2005 3625 2010 3655
rect 2040 3625 2045 3655
rect 2005 3615 2045 3625
rect 2205 3625 2210 3655
rect 2240 3625 2245 3655
rect 2205 3615 2245 3625
rect 2405 3625 2410 3655
rect 2440 3625 2445 3655
rect 2405 3615 2445 3625
rect 2605 3625 2610 3655
rect 2640 3625 2645 3655
rect 2605 3615 2645 3625
rect 2805 3625 2810 3655
rect 2840 3625 2845 3655
rect 2805 3615 2845 3625
rect 3005 3625 3010 3655
rect 3040 3625 3045 3655
rect 3005 3615 3045 3625
rect 3205 3625 3210 3655
rect 3240 3625 3245 3655
rect 3205 3615 3245 3625
rect 3405 3625 3410 3655
rect 3440 3625 3445 3655
rect 3405 3615 3445 3625
rect 3605 3625 3610 3655
rect 3640 3625 3645 3655
rect 3605 3615 3645 3625
rect 3805 3625 3810 3655
rect 3840 3625 3845 3655
rect 3805 3615 3845 3625
rect 4005 3625 4010 3655
rect 4040 3625 4045 3655
rect 4005 3615 4045 3625
rect 4205 3625 4210 3655
rect 4240 3625 4245 3655
rect 4205 3615 4245 3625
rect 4405 3625 4410 3655
rect 4440 3625 4445 3655
rect 4405 3615 4445 3625
rect 4605 3625 4610 3655
rect 4640 3625 4645 3655
rect 4605 3615 4645 3625
rect 4805 3625 4810 3655
rect 4840 3625 4845 3655
rect 4805 3615 4845 3625
rect 5005 3625 5010 3655
rect 5040 3625 5045 3655
rect 5005 3615 5045 3625
rect 5205 3625 5210 3655
rect 5240 3625 5245 3655
rect 5205 3615 5245 3625
rect 5405 3625 5410 3655
rect 5440 3625 5445 3655
rect 5405 3615 5445 3625
rect 5605 3625 5610 3655
rect 5640 3625 5645 3655
rect 5605 3615 5645 3625
rect 5805 3625 5810 3655
rect 5840 3625 5845 3655
rect 5805 3615 5845 3625
rect 6005 3625 6010 3655
rect 6040 3625 6045 3655
rect 6005 3615 6045 3625
rect 6205 3625 6210 3655
rect 6240 3625 6245 3655
rect 6205 3615 6245 3625
rect 6405 3625 6410 3655
rect 6440 3625 6445 3655
rect 6405 3615 6445 3625
rect -165 3595 -30 3615
rect 5 3595 1570 3615
rect 1605 3595 2970 3615
rect 3005 3595 6570 3615
rect -165 3585 -155 3595
rect -195 3555 -190 3585
rect -160 3555 -155 3585
rect 5 3585 45 3595
rect 5 3555 10 3585
rect 40 3555 45 3585
rect 205 3585 245 3595
rect 205 3555 210 3585
rect 240 3555 245 3585
rect 405 3585 445 3595
rect 405 3555 410 3585
rect 440 3555 445 3585
rect 605 3585 645 3595
rect 605 3555 610 3585
rect 640 3555 645 3585
rect 805 3585 845 3595
rect 805 3555 810 3585
rect 840 3555 845 3585
rect 1005 3585 1045 3595
rect 1005 3555 1010 3585
rect 1040 3555 1045 3585
rect 1205 3585 1245 3595
rect 1205 3555 1210 3585
rect 1240 3555 1245 3585
rect 1405 3585 1445 3595
rect 1405 3555 1410 3585
rect 1440 3555 1445 3585
rect 1605 3585 1645 3595
rect 1605 3555 1610 3585
rect 1640 3555 1645 3585
rect 1805 3585 1845 3595
rect 1805 3555 1810 3585
rect 1840 3555 1845 3585
rect 2005 3585 2045 3595
rect 2005 3555 2010 3585
rect 2040 3555 2045 3585
rect 2205 3585 2245 3595
rect 2205 3555 2210 3585
rect 2240 3555 2245 3585
rect 2405 3585 2445 3595
rect 2405 3555 2410 3585
rect 2440 3555 2445 3585
rect 2605 3585 2645 3595
rect 2605 3555 2610 3585
rect 2640 3555 2645 3585
rect 2805 3585 2845 3595
rect 2805 3555 2810 3585
rect 2840 3555 2845 3585
rect 3005 3585 3045 3595
rect 3005 3555 3010 3585
rect 3040 3555 3045 3585
rect 3205 3585 3245 3595
rect 3205 3555 3210 3585
rect 3240 3555 3245 3585
rect 3405 3585 3445 3595
rect 3405 3555 3410 3585
rect 3440 3555 3445 3585
rect 3605 3585 3645 3595
rect 3605 3555 3610 3585
rect 3640 3555 3645 3585
rect 3805 3585 3845 3595
rect 3805 3555 3810 3585
rect 3840 3555 3845 3585
rect 4005 3585 4045 3595
rect 4005 3555 4010 3585
rect 4040 3555 4045 3585
rect 4205 3585 4245 3595
rect 4205 3555 4210 3585
rect 4240 3555 4245 3585
rect 4405 3585 4445 3595
rect 4405 3555 4410 3585
rect 4440 3555 4445 3585
rect 4605 3585 4645 3595
rect 4605 3555 4610 3585
rect 4640 3555 4645 3585
rect 4805 3585 4845 3595
rect 4805 3555 4810 3585
rect 4840 3555 4845 3585
rect 5005 3585 5045 3595
rect 5005 3555 5010 3585
rect 5040 3555 5045 3585
rect 5205 3585 5245 3595
rect 5205 3555 5210 3585
rect 5240 3555 5245 3585
rect 5405 3585 5445 3595
rect 5405 3555 5410 3585
rect 5440 3555 5445 3585
rect 5605 3585 5645 3595
rect 5605 3555 5610 3585
rect 5640 3555 5645 3585
rect 5805 3585 5845 3595
rect 5805 3555 5810 3585
rect 5840 3555 5845 3585
rect 6005 3585 6045 3595
rect 6005 3555 6010 3585
rect 6040 3555 6045 3585
rect 6205 3585 6245 3595
rect 6205 3555 6210 3585
rect 6240 3555 6245 3585
rect 6405 3585 6445 3595
rect 6405 3555 6410 3585
rect 6440 3555 6445 3585
rect -188 3470 -185 3555
rect -165 3470 -162 3555
rect 15 3470 35 3555
rect 215 3470 235 3555
rect 415 3470 435 3555
rect 615 3470 635 3555
rect 815 3470 835 3555
rect 1015 3470 1035 3555
rect 1215 3470 1235 3555
rect 1415 3470 1435 3555
rect 1615 3470 1635 3555
rect 1815 3470 1835 3555
rect 2015 3470 2035 3555
rect 2215 3470 2235 3555
rect 2415 3470 2435 3555
rect 2615 3470 2635 3555
rect 2815 3470 2835 3555
rect 3015 3470 3035 3555
rect 3215 3470 3235 3555
rect 3415 3470 3435 3555
rect 3615 3470 3635 3555
rect 3815 3470 3835 3555
rect 4015 3470 4035 3555
rect 4215 3470 4235 3555
rect 4415 3470 4435 3555
rect 4615 3470 4635 3555
rect 4815 3470 4835 3555
rect 5015 3470 5035 3555
rect 5215 3470 5235 3555
rect 5415 3470 5435 3555
rect 5615 3470 5635 3555
rect 5815 3470 5835 3555
rect 6015 3470 6035 3555
rect 6215 3470 6235 3555
rect -195 3440 -190 3470
rect -160 3440 -155 3470
rect -195 3400 -185 3440
rect -165 3430 -155 3440
rect 5 3440 10 3470
rect 40 3440 45 3470
rect 5 3430 45 3440
rect 205 3440 210 3470
rect 240 3440 245 3470
rect 205 3430 245 3440
rect 405 3440 410 3470
rect 440 3440 445 3470
rect 405 3430 445 3440
rect 605 3440 610 3470
rect 640 3440 645 3470
rect 605 3430 645 3440
rect 805 3440 810 3470
rect 840 3440 845 3470
rect 805 3430 845 3440
rect 1005 3440 1010 3470
rect 1040 3440 1045 3470
rect 1005 3430 1045 3440
rect 1205 3440 1210 3470
rect 1240 3440 1245 3470
rect 1205 3430 1245 3440
rect 1405 3440 1410 3470
rect 1440 3440 1445 3470
rect 1405 3430 1445 3440
rect 1605 3440 1610 3470
rect 1640 3440 1645 3470
rect 1605 3430 1645 3440
rect 1805 3440 1810 3470
rect 1840 3440 1845 3470
rect 1805 3430 1845 3440
rect 2005 3440 2010 3470
rect 2040 3440 2045 3470
rect 2005 3430 2045 3440
rect 2205 3440 2210 3470
rect 2240 3440 2245 3470
rect 2205 3430 2245 3440
rect 2405 3440 2410 3470
rect 2440 3440 2445 3470
rect 2405 3430 2445 3440
rect 2605 3440 2610 3470
rect 2640 3440 2645 3470
rect 2605 3430 2645 3440
rect 2805 3440 2810 3470
rect 2840 3440 2845 3470
rect 2805 3430 2845 3440
rect 3005 3440 3010 3470
rect 3040 3440 3045 3470
rect 3005 3430 3045 3440
rect 3205 3440 3210 3470
rect 3240 3440 3245 3470
rect 3205 3430 3245 3440
rect 3405 3440 3410 3470
rect 3440 3440 3445 3470
rect 3405 3430 3445 3440
rect 3605 3440 3610 3470
rect 3640 3440 3645 3470
rect 3605 3430 3645 3440
rect 3805 3440 3810 3470
rect 3840 3440 3845 3470
rect 3805 3430 3845 3440
rect 4005 3440 4010 3470
rect 4040 3440 4045 3470
rect 4005 3430 4045 3440
rect 4205 3440 4210 3470
rect 4240 3440 4245 3470
rect 4205 3430 4245 3440
rect 4405 3440 4410 3470
rect 4440 3440 4445 3470
rect 4405 3430 4445 3440
rect 4605 3440 4610 3470
rect 4640 3440 4645 3470
rect 4605 3430 4645 3440
rect 4805 3440 4810 3470
rect 4840 3440 4845 3470
rect 4805 3430 4845 3440
rect 5005 3440 5010 3470
rect 5040 3440 5045 3470
rect 5005 3430 5045 3440
rect 5205 3440 5210 3470
rect 5240 3440 5245 3470
rect 5205 3430 5245 3440
rect 5405 3440 5410 3470
rect 5440 3440 5445 3470
rect 5405 3430 5445 3440
rect 5605 3440 5610 3470
rect 5640 3440 5645 3470
rect 5605 3430 5645 3440
rect 5805 3440 5810 3470
rect 5840 3440 5845 3470
rect 5805 3430 5845 3440
rect 6005 3440 6010 3470
rect 6040 3440 6045 3470
rect 6005 3430 6045 3440
rect 6205 3440 6210 3470
rect 6240 3440 6245 3470
rect 6205 3430 6245 3440
rect 6405 3440 6410 3470
rect 6440 3440 6445 3470
rect 6405 3430 6445 3440
rect -165 3410 -30 3430
rect 5 3410 1570 3430
rect 1605 3410 2970 3430
rect 3005 3410 6570 3430
rect -165 3400 -155 3410
rect -195 3370 -190 3400
rect -160 3370 -155 3400
rect 5 3400 45 3410
rect 5 3370 10 3400
rect 40 3370 45 3400
rect 205 3400 245 3410
rect 205 3370 210 3400
rect 240 3370 245 3400
rect 405 3400 445 3410
rect 405 3370 410 3400
rect 440 3370 445 3400
rect 605 3400 645 3410
rect 605 3370 610 3400
rect 640 3370 645 3400
rect 805 3400 845 3410
rect 805 3370 810 3400
rect 840 3370 845 3400
rect 1005 3400 1045 3410
rect 1005 3370 1010 3400
rect 1040 3370 1045 3400
rect 1205 3400 1245 3410
rect 1205 3370 1210 3400
rect 1240 3370 1245 3400
rect 1405 3400 1445 3410
rect 1405 3370 1410 3400
rect 1440 3370 1445 3400
rect 1605 3400 1645 3410
rect 1605 3370 1610 3400
rect 1640 3370 1645 3400
rect 1805 3400 1845 3410
rect 1805 3370 1810 3400
rect 1840 3370 1845 3400
rect 2005 3400 2045 3410
rect 2005 3370 2010 3400
rect 2040 3370 2045 3400
rect 2205 3400 2245 3410
rect 2205 3370 2210 3400
rect 2240 3370 2245 3400
rect 2405 3400 2445 3410
rect 2405 3370 2410 3400
rect 2440 3370 2445 3400
rect 2605 3400 2645 3410
rect 2605 3370 2610 3400
rect 2640 3370 2645 3400
rect 2805 3400 2845 3410
rect 2805 3370 2810 3400
rect 2840 3370 2845 3400
rect 3005 3400 3045 3410
rect 3005 3370 3010 3400
rect 3040 3370 3045 3400
rect 3205 3400 3245 3410
rect 3205 3370 3210 3400
rect 3240 3370 3245 3400
rect 3405 3400 3445 3410
rect 3405 3370 3410 3400
rect 3440 3370 3445 3400
rect 3605 3400 3645 3410
rect 3605 3370 3610 3400
rect 3640 3370 3645 3400
rect 3805 3400 3845 3410
rect 3805 3370 3810 3400
rect 3840 3370 3845 3400
rect 4005 3400 4045 3410
rect 4005 3370 4010 3400
rect 4040 3370 4045 3400
rect 4205 3400 4245 3410
rect 4205 3370 4210 3400
rect 4240 3370 4245 3400
rect 4405 3400 4445 3410
rect 4405 3370 4410 3400
rect 4440 3370 4445 3400
rect 4605 3400 4645 3410
rect 4605 3370 4610 3400
rect 4640 3370 4645 3400
rect 4805 3400 4845 3410
rect 4805 3370 4810 3400
rect 4840 3370 4845 3400
rect 5005 3400 5045 3410
rect 5005 3370 5010 3400
rect 5040 3370 5045 3400
rect 5205 3400 5245 3410
rect 5205 3370 5210 3400
rect 5240 3370 5245 3400
rect 5405 3400 5445 3410
rect 5405 3370 5410 3400
rect 5440 3370 5445 3400
rect 5605 3400 5645 3410
rect 5605 3370 5610 3400
rect 5640 3370 5645 3400
rect 5805 3400 5845 3410
rect 5805 3370 5810 3400
rect 5840 3370 5845 3400
rect 6005 3400 6045 3410
rect 6005 3370 6010 3400
rect 6040 3370 6045 3400
rect 6205 3400 6245 3410
rect 6205 3370 6210 3400
rect 6240 3370 6245 3400
rect 6405 3400 6445 3410
rect 6405 3370 6410 3400
rect 6440 3370 6445 3400
rect -188 3285 -185 3370
rect -165 3285 -162 3370
rect 15 3285 35 3370
rect 215 3285 235 3370
rect 415 3285 435 3370
rect 615 3285 635 3370
rect 815 3285 835 3370
rect 1015 3285 1035 3370
rect 1215 3285 1235 3370
rect 1415 3285 1435 3370
rect 1615 3285 1635 3370
rect 1815 3285 1835 3370
rect 2015 3285 2035 3370
rect 2215 3285 2235 3370
rect 2415 3285 2435 3370
rect 2615 3285 2635 3370
rect 2815 3285 2835 3370
rect 3015 3285 3035 3370
rect 3215 3285 3235 3370
rect 3415 3285 3435 3370
rect 3615 3285 3635 3370
rect 3815 3285 3835 3370
rect 4015 3285 4035 3370
rect 4215 3285 4235 3370
rect 4415 3285 4435 3370
rect 4615 3285 4635 3370
rect 4815 3285 4835 3370
rect 5015 3285 5035 3370
rect 5215 3285 5235 3370
rect 5415 3285 5435 3370
rect 5615 3285 5635 3370
rect 5815 3285 5835 3370
rect 6015 3285 6035 3370
rect 6215 3285 6235 3370
rect -195 3255 -190 3285
rect -160 3255 -155 3285
rect -195 3215 -185 3255
rect -165 3245 -155 3255
rect 5 3255 10 3285
rect 40 3255 45 3285
rect 5 3245 45 3255
rect 205 3255 210 3285
rect 240 3255 245 3285
rect 205 3245 245 3255
rect 405 3255 410 3285
rect 440 3255 445 3285
rect 405 3245 445 3255
rect 605 3255 610 3285
rect 640 3255 645 3285
rect 605 3245 645 3255
rect 805 3255 810 3285
rect 840 3255 845 3285
rect 805 3245 845 3255
rect 1005 3255 1010 3285
rect 1040 3255 1045 3285
rect 1005 3245 1045 3255
rect 1205 3255 1210 3285
rect 1240 3255 1245 3285
rect 1205 3245 1245 3255
rect 1405 3255 1410 3285
rect 1440 3255 1445 3285
rect 1405 3245 1445 3255
rect 1605 3255 1610 3285
rect 1640 3255 1645 3285
rect 1605 3245 1645 3255
rect 1805 3255 1810 3285
rect 1840 3255 1845 3285
rect 1805 3245 1845 3255
rect 2005 3255 2010 3285
rect 2040 3255 2045 3285
rect 2005 3245 2045 3255
rect 2205 3255 2210 3285
rect 2240 3255 2245 3285
rect 2205 3245 2245 3255
rect 2405 3255 2410 3285
rect 2440 3255 2445 3285
rect 2405 3245 2445 3255
rect 2605 3255 2610 3285
rect 2640 3255 2645 3285
rect 2605 3245 2645 3255
rect 2805 3255 2810 3285
rect 2840 3255 2845 3285
rect 2805 3245 2845 3255
rect 3005 3255 3010 3285
rect 3040 3255 3045 3285
rect 3005 3245 3045 3255
rect 3205 3255 3210 3285
rect 3240 3255 3245 3285
rect 3205 3245 3245 3255
rect 3405 3255 3410 3285
rect 3440 3255 3445 3285
rect 3405 3245 3445 3255
rect 3605 3255 3610 3285
rect 3640 3255 3645 3285
rect 3605 3245 3645 3255
rect 3805 3255 3810 3285
rect 3840 3255 3845 3285
rect 3805 3245 3845 3255
rect 4005 3255 4010 3285
rect 4040 3255 4045 3285
rect 4005 3245 4045 3255
rect 4205 3255 4210 3285
rect 4240 3255 4245 3285
rect 4205 3245 4245 3255
rect 4405 3255 4410 3285
rect 4440 3255 4445 3285
rect 4405 3245 4445 3255
rect 4605 3255 4610 3285
rect 4640 3255 4645 3285
rect 4605 3245 4645 3255
rect 4805 3255 4810 3285
rect 4840 3255 4845 3285
rect 4805 3245 4845 3255
rect 5005 3255 5010 3285
rect 5040 3255 5045 3285
rect 5005 3245 5045 3255
rect 5205 3255 5210 3285
rect 5240 3255 5245 3285
rect 5205 3245 5245 3255
rect 5405 3255 5410 3285
rect 5440 3255 5445 3285
rect 5405 3245 5445 3255
rect 5605 3255 5610 3285
rect 5640 3255 5645 3285
rect 5605 3245 5645 3255
rect 5805 3255 5810 3285
rect 5840 3255 5845 3285
rect 5805 3245 5845 3255
rect 6005 3255 6010 3285
rect 6040 3255 6045 3285
rect 6005 3245 6045 3255
rect 6205 3255 6210 3285
rect 6240 3255 6245 3285
rect 6205 3245 6245 3255
rect 6405 3255 6410 3285
rect 6440 3255 6445 3285
rect 6405 3245 6445 3255
rect -165 3225 -30 3245
rect 5 3225 1570 3245
rect 1605 3225 2970 3245
rect 3005 3225 6570 3245
rect -165 3215 -155 3225
rect -195 3185 -190 3215
rect -160 3185 -155 3215
rect 5 3215 45 3225
rect 5 3185 10 3215
rect 40 3185 45 3215
rect 205 3215 245 3225
rect 205 3185 210 3215
rect 240 3185 245 3215
rect 405 3215 445 3225
rect 405 3185 410 3215
rect 440 3185 445 3215
rect 605 3215 645 3225
rect 605 3185 610 3215
rect 640 3185 645 3215
rect 805 3215 845 3225
rect 805 3185 810 3215
rect 840 3185 845 3215
rect 1005 3215 1045 3225
rect 1005 3185 1010 3215
rect 1040 3185 1045 3215
rect 1205 3215 1245 3225
rect 1205 3185 1210 3215
rect 1240 3185 1245 3215
rect 1405 3215 1445 3225
rect 1405 3185 1410 3215
rect 1440 3185 1445 3215
rect 1605 3215 1645 3225
rect 1605 3185 1610 3215
rect 1640 3185 1645 3215
rect 1805 3215 1845 3225
rect 1805 3185 1810 3215
rect 1840 3185 1845 3215
rect 2005 3215 2045 3225
rect 2005 3185 2010 3215
rect 2040 3185 2045 3215
rect 2205 3215 2245 3225
rect 2205 3185 2210 3215
rect 2240 3185 2245 3215
rect 2405 3215 2445 3225
rect 2405 3185 2410 3215
rect 2440 3185 2445 3215
rect 2605 3215 2645 3225
rect 2605 3185 2610 3215
rect 2640 3185 2645 3215
rect 2805 3215 2845 3225
rect 2805 3185 2810 3215
rect 2840 3185 2845 3215
rect 3005 3215 3045 3225
rect 3005 3185 3010 3215
rect 3040 3185 3045 3215
rect 3205 3215 3245 3225
rect 3205 3185 3210 3215
rect 3240 3185 3245 3215
rect 3405 3215 3445 3225
rect 3405 3185 3410 3215
rect 3440 3185 3445 3215
rect 3605 3215 3645 3225
rect 3605 3185 3610 3215
rect 3640 3185 3645 3215
rect 3805 3215 3845 3225
rect 3805 3185 3810 3215
rect 3840 3185 3845 3215
rect 4005 3215 4045 3225
rect 4005 3185 4010 3215
rect 4040 3185 4045 3215
rect 4205 3215 4245 3225
rect 4205 3185 4210 3215
rect 4240 3185 4245 3215
rect 4405 3215 4445 3225
rect 4405 3185 4410 3215
rect 4440 3185 4445 3215
rect 4605 3215 4645 3225
rect 4605 3185 4610 3215
rect 4640 3185 4645 3215
rect 4805 3215 4845 3225
rect 4805 3185 4810 3215
rect 4840 3185 4845 3215
rect 5005 3215 5045 3225
rect 5005 3185 5010 3215
rect 5040 3185 5045 3215
rect 5205 3215 5245 3225
rect 5205 3185 5210 3215
rect 5240 3185 5245 3215
rect 5405 3215 5445 3225
rect 5405 3185 5410 3215
rect 5440 3185 5445 3215
rect 5605 3215 5645 3225
rect 5605 3185 5610 3215
rect 5640 3185 5645 3215
rect 5805 3215 5845 3225
rect 5805 3185 5810 3215
rect 5840 3185 5845 3215
rect 6005 3215 6045 3225
rect 6005 3185 6010 3215
rect 6040 3185 6045 3215
rect 6205 3215 6245 3225
rect 6205 3185 6210 3215
rect 6240 3185 6245 3215
rect 6405 3215 6445 3225
rect 6405 3185 6410 3215
rect 6440 3185 6445 3215
rect -188 3100 -185 3185
rect -165 3100 -162 3185
rect 15 3100 35 3185
rect 215 3100 235 3185
rect 415 3100 435 3185
rect 615 3100 635 3185
rect 815 3100 835 3185
rect 1015 3100 1035 3185
rect 1215 3100 1235 3185
rect 1415 3100 1435 3185
rect 1615 3100 1635 3185
rect 1815 3100 1835 3185
rect 2015 3100 2035 3185
rect 2215 3100 2235 3185
rect 2415 3100 2435 3185
rect 2615 3100 2635 3185
rect 2815 3100 2835 3185
rect -195 3070 -190 3100
rect -160 3070 -155 3100
rect -195 3030 -185 3070
rect -165 3060 -155 3070
rect 5 3070 10 3100
rect 40 3070 45 3100
rect 5 3060 45 3070
rect 205 3070 210 3100
rect 240 3070 245 3100
rect 205 3060 245 3070
rect 405 3070 410 3100
rect 440 3070 445 3100
rect 405 3060 445 3070
rect 605 3070 610 3100
rect 640 3070 645 3100
rect 605 3060 645 3070
rect 805 3070 810 3100
rect 840 3070 845 3100
rect 805 3060 845 3070
rect 1005 3070 1010 3100
rect 1040 3070 1045 3100
rect 1005 3060 1045 3070
rect 1205 3070 1210 3100
rect 1240 3070 1245 3100
rect 1205 3060 1245 3070
rect 1405 3070 1410 3100
rect 1440 3070 1445 3100
rect 1405 3060 1445 3070
rect 1605 3070 1610 3100
rect 1640 3070 1645 3100
rect 1605 3060 1645 3070
rect 1805 3070 1810 3100
rect 1840 3070 1845 3100
rect 1805 3060 1845 3070
rect 2005 3070 2010 3100
rect 2040 3070 2045 3100
rect 2005 3060 2045 3070
rect 2205 3070 2210 3100
rect 2240 3070 2245 3100
rect 2205 3060 2245 3070
rect 2405 3070 2410 3100
rect 2440 3070 2445 3100
rect 2405 3060 2445 3070
rect 2605 3070 2610 3100
rect 2640 3070 2645 3100
rect 2605 3060 2645 3070
rect 2805 3070 2810 3100
rect 2840 3070 2845 3100
rect 2805 3060 2845 3070
rect 3005 3070 3010 3100
rect 3040 3070 3045 3100
rect 3005 3060 3045 3070
rect 3205 3070 3210 3100
rect 3240 3070 3245 3100
rect 3205 3060 3245 3070
rect 3405 3070 3410 3100
rect 3440 3070 3445 3100
rect 3405 3060 3445 3070
rect 3605 3070 3610 3100
rect 3640 3070 3645 3100
rect 3605 3060 3645 3070
rect 3805 3070 3810 3100
rect 3840 3070 3845 3100
rect 3805 3060 3845 3070
rect 4005 3070 4010 3100
rect 4040 3070 4045 3100
rect 4005 3060 4045 3070
rect 4205 3070 4210 3100
rect 4240 3070 4245 3100
rect 4205 3060 4245 3070
rect 4405 3070 4410 3100
rect 4440 3070 4445 3100
rect 4405 3060 4445 3070
rect 4605 3070 4610 3100
rect 4640 3070 4645 3100
rect 4605 3060 4645 3070
rect 4805 3070 4810 3100
rect 4840 3070 4845 3100
rect 4805 3060 4845 3070
rect 5005 3070 5010 3100
rect 5040 3070 5045 3100
rect 5005 3060 5045 3070
rect 5205 3070 5210 3100
rect 5240 3070 5245 3100
rect 5205 3060 5245 3070
rect 5405 3070 5410 3100
rect 5440 3070 5445 3100
rect 5405 3060 5445 3070
rect 5605 3070 5610 3100
rect 5640 3070 5645 3100
rect 5605 3060 5645 3070
rect 5805 3070 5810 3100
rect 5840 3070 5845 3100
rect 5805 3060 5845 3070
rect 6005 3070 6010 3100
rect 6040 3070 6045 3100
rect 6005 3060 6045 3070
rect 6205 3070 6210 3100
rect 6240 3070 6245 3100
rect 6205 3060 6245 3070
rect 6405 3070 6410 3100
rect 6440 3070 6445 3100
rect 6405 3060 6445 3070
rect -165 3040 -30 3060
rect 5 3040 1570 3060
rect 1605 3040 6695 3060
rect -165 3030 -155 3040
rect -195 3000 -190 3030
rect -160 3000 -155 3030
rect 5 3030 45 3040
rect 5 3000 10 3030
rect 40 3000 45 3030
rect 205 3030 245 3040
rect 205 3000 210 3030
rect 240 3000 245 3030
rect 405 3030 445 3040
rect 405 3000 410 3030
rect 440 3000 445 3030
rect 605 3030 645 3040
rect 605 3000 610 3030
rect 640 3000 645 3030
rect 805 3030 845 3040
rect 805 3000 810 3030
rect 840 3000 845 3030
rect 1005 3030 1045 3040
rect 1005 3000 1010 3030
rect 1040 3000 1045 3030
rect 1205 3030 1245 3040
rect 1205 3000 1210 3030
rect 1240 3000 1245 3030
rect 1405 3030 1445 3040
rect 1405 3000 1410 3030
rect 1440 3000 1445 3030
rect 1605 3030 1645 3040
rect 1605 3000 1610 3030
rect 1640 3000 1645 3030
rect 1805 3030 1845 3040
rect 1805 3000 1810 3030
rect 1840 3000 1845 3030
rect 2005 3030 2045 3040
rect 2005 3000 2010 3030
rect 2040 3000 2045 3030
rect 2205 3030 2245 3040
rect 2205 3000 2210 3030
rect 2240 3000 2245 3030
rect 2405 3030 2445 3040
rect 2405 3000 2410 3030
rect 2440 3000 2445 3030
rect 2605 3030 2645 3040
rect 2605 3000 2610 3030
rect 2640 3000 2645 3030
rect 2805 3030 2845 3040
rect 2805 3000 2810 3030
rect 2840 3000 2845 3030
rect 3005 3030 3045 3040
rect 3005 3000 3010 3030
rect 3040 3000 3045 3030
rect 3205 3030 3245 3040
rect 3205 3000 3210 3030
rect 3240 3000 3245 3030
rect 3405 3030 3445 3040
rect 3405 3000 3410 3030
rect 3440 3000 3445 3030
rect 3605 3030 3645 3040
rect 3605 3000 3610 3030
rect 3640 3000 3645 3030
rect 3805 3030 3845 3040
rect 3805 3000 3810 3030
rect 3840 3000 3845 3030
rect 4005 3030 4045 3040
rect 4005 3000 4010 3030
rect 4040 3000 4045 3030
rect 4205 3030 4245 3040
rect 4205 3000 4210 3030
rect 4240 3000 4245 3030
rect 4405 3030 4445 3040
rect 4405 3000 4410 3030
rect 4440 3000 4445 3030
rect 4605 3030 4645 3040
rect 4605 3000 4610 3030
rect 4640 3000 4645 3030
rect 4805 3030 4845 3040
rect 4805 3000 4810 3030
rect 4840 3000 4845 3030
rect 5005 3030 5045 3040
rect 5005 3000 5010 3030
rect 5040 3000 5045 3030
rect 5205 3030 5245 3040
rect 5205 3000 5210 3030
rect 5240 3000 5245 3030
rect 5405 3030 5445 3040
rect 5405 3000 5410 3030
rect 5440 3000 5445 3030
rect 5605 3030 5645 3040
rect 5605 3000 5610 3030
rect 5640 3000 5645 3030
rect 5805 3030 5845 3040
rect 5805 3000 5810 3030
rect 5840 3000 5845 3030
rect 6005 3030 6045 3040
rect 6005 3000 6010 3030
rect 6040 3000 6045 3030
rect 6205 3030 6245 3040
rect 6205 3000 6210 3030
rect 6240 3000 6245 3030
rect 6405 3030 6445 3040
rect 6405 3000 6410 3030
rect 6440 3000 6445 3030
rect -188 2915 -185 3000
rect -165 2915 -162 3000
rect 15 2915 35 3000
rect 215 2915 235 3000
rect 415 2915 435 3000
rect 615 2915 635 3000
rect 815 2915 835 3000
rect 1015 2915 1035 3000
rect 1215 2915 1235 3000
rect 1415 2915 1435 3000
rect 1615 2915 1635 3000
rect 1815 2915 1835 3000
rect 2015 2915 2035 3000
rect 2215 2915 2235 3000
rect 2415 2915 2435 3000
rect 2615 2915 2635 3000
rect 2815 2915 2835 3000
rect 3015 2915 3035 3000
rect 3215 2915 3235 3000
rect 3415 2915 3435 3000
rect 3615 2915 3635 3000
rect 3815 2915 3835 3000
rect 4015 2915 4035 3000
rect 4215 2915 4235 3000
rect 4415 2915 4435 3000
rect 4615 2915 4635 3000
rect 4815 2915 4835 3000
rect 5015 2915 5035 3000
rect 5215 2915 5235 3000
rect 5415 2915 5435 3000
rect 5615 2915 5635 3000
rect 5815 2915 5835 3000
rect 6015 2915 6035 3000
rect 6215 2915 6235 3000
rect -195 2885 -190 2915
rect -160 2885 -155 2915
rect -195 2845 -185 2885
rect -165 2875 -155 2885
rect 5 2885 10 2915
rect 40 2885 45 2915
rect 5 2875 45 2885
rect 205 2885 210 2915
rect 240 2885 245 2915
rect 205 2875 245 2885
rect 405 2885 410 2915
rect 440 2885 445 2915
rect 405 2875 445 2885
rect 605 2885 610 2915
rect 640 2885 645 2915
rect 605 2875 645 2885
rect 805 2885 810 2915
rect 840 2885 845 2915
rect 805 2875 845 2885
rect 1005 2885 1010 2915
rect 1040 2885 1045 2915
rect 1005 2875 1045 2885
rect 1205 2885 1210 2915
rect 1240 2885 1245 2915
rect 1205 2875 1245 2885
rect 1405 2885 1410 2915
rect 1440 2885 1445 2915
rect 1405 2875 1445 2885
rect 1605 2885 1610 2915
rect 1640 2885 1645 2915
rect 1605 2875 1645 2885
rect 1805 2885 1810 2915
rect 1840 2885 1845 2915
rect 1805 2875 1845 2885
rect 2005 2885 2010 2915
rect 2040 2885 2045 2915
rect 2005 2875 2045 2885
rect 2205 2885 2210 2915
rect 2240 2885 2245 2915
rect 2205 2875 2245 2885
rect 2405 2885 2410 2915
rect 2440 2885 2445 2915
rect 2405 2875 2445 2885
rect 2605 2885 2610 2915
rect 2640 2885 2645 2915
rect 2605 2875 2645 2885
rect 2805 2885 2810 2915
rect 2840 2885 2845 2915
rect 2805 2875 2845 2885
rect 3005 2885 3010 2915
rect 3040 2885 3045 2915
rect 3005 2875 3045 2885
rect 3205 2885 3210 2915
rect 3240 2885 3245 2915
rect 3205 2875 3245 2885
rect 3405 2885 3410 2915
rect 3440 2885 3445 2915
rect 3405 2875 3445 2885
rect 3605 2885 3610 2915
rect 3640 2885 3645 2915
rect 3605 2875 3645 2885
rect 3805 2885 3810 2915
rect 3840 2885 3845 2915
rect 3805 2875 3845 2885
rect 4005 2885 4010 2915
rect 4040 2885 4045 2915
rect 4005 2875 4045 2885
rect 4205 2885 4210 2915
rect 4240 2885 4245 2915
rect 4205 2875 4245 2885
rect 4405 2885 4410 2915
rect 4440 2885 4445 2915
rect 4405 2875 4445 2885
rect 4605 2885 4610 2915
rect 4640 2885 4645 2915
rect 4605 2875 4645 2885
rect 4805 2885 4810 2915
rect 4840 2885 4845 2915
rect 4805 2875 4845 2885
rect 5005 2885 5010 2915
rect 5040 2885 5045 2915
rect 5005 2875 5045 2885
rect 5205 2885 5210 2915
rect 5240 2885 5245 2915
rect 5205 2875 5245 2885
rect 5405 2885 5410 2915
rect 5440 2885 5445 2915
rect 5405 2875 5445 2885
rect 5605 2885 5610 2915
rect 5640 2885 5645 2915
rect 5605 2875 5645 2885
rect 5805 2885 5810 2915
rect 5840 2885 5845 2915
rect 5805 2875 5845 2885
rect 6005 2885 6010 2915
rect 6040 2885 6045 2915
rect 6005 2875 6045 2885
rect 6205 2885 6210 2915
rect 6240 2885 6245 2915
rect 6205 2875 6245 2885
rect 6405 2885 6410 2915
rect 6440 2885 6445 2915
rect 6405 2875 6445 2885
rect -165 2855 -30 2875
rect 5 2855 1570 2875
rect 1605 2855 6570 2875
rect -165 2845 -155 2855
rect -195 2815 -190 2845
rect -160 2815 -155 2845
rect 5 2845 45 2855
rect 5 2815 10 2845
rect 40 2815 45 2845
rect 205 2845 245 2855
rect 205 2815 210 2845
rect 240 2815 245 2845
rect 405 2845 445 2855
rect 405 2815 410 2845
rect 440 2815 445 2845
rect 605 2845 645 2855
rect 605 2815 610 2845
rect 640 2815 645 2845
rect 805 2845 845 2855
rect 805 2815 810 2845
rect 840 2815 845 2845
rect 1005 2845 1045 2855
rect 1005 2815 1010 2845
rect 1040 2815 1045 2845
rect 1205 2845 1245 2855
rect 1205 2815 1210 2845
rect 1240 2815 1245 2845
rect 1405 2845 1445 2855
rect 1405 2815 1410 2845
rect 1440 2815 1445 2845
rect 1605 2845 1645 2855
rect 1605 2815 1610 2845
rect 1640 2815 1645 2845
rect 1805 2845 1845 2855
rect 1805 2815 1810 2845
rect 1840 2815 1845 2845
rect 2005 2845 2045 2855
rect 2005 2815 2010 2845
rect 2040 2815 2045 2845
rect 2205 2845 2245 2855
rect 2205 2815 2210 2845
rect 2240 2815 2245 2845
rect 2405 2845 2445 2855
rect 2405 2815 2410 2845
rect 2440 2815 2445 2845
rect 2605 2845 2645 2855
rect 2605 2815 2610 2845
rect 2640 2815 2645 2845
rect 2805 2845 2845 2855
rect 2805 2815 2810 2845
rect 2840 2815 2845 2845
rect 3005 2845 3045 2855
rect 3005 2815 3010 2845
rect 3040 2815 3045 2845
rect 3205 2845 3245 2855
rect 3205 2815 3210 2845
rect 3240 2815 3245 2845
rect 3405 2845 3445 2855
rect 3405 2815 3410 2845
rect 3440 2815 3445 2845
rect 3605 2845 3645 2855
rect 3605 2815 3610 2845
rect 3640 2815 3645 2845
rect 3805 2845 3845 2855
rect 3805 2815 3810 2845
rect 3840 2815 3845 2845
rect 4005 2845 4045 2855
rect 4005 2815 4010 2845
rect 4040 2815 4045 2845
rect 4205 2845 4245 2855
rect 4205 2815 4210 2845
rect 4240 2815 4245 2845
rect 4405 2845 4445 2855
rect 4405 2815 4410 2845
rect 4440 2815 4445 2845
rect 4605 2845 4645 2855
rect 4605 2815 4610 2845
rect 4640 2815 4645 2845
rect 4805 2845 4845 2855
rect 4805 2815 4810 2845
rect 4840 2815 4845 2845
rect 5005 2845 5045 2855
rect 5005 2815 5010 2845
rect 5040 2815 5045 2845
rect 5205 2845 5245 2855
rect 5205 2815 5210 2845
rect 5240 2815 5245 2845
rect 5405 2845 5445 2855
rect 5405 2815 5410 2845
rect 5440 2815 5445 2845
rect 5605 2845 5645 2855
rect 5605 2815 5610 2845
rect 5640 2815 5645 2845
rect 5805 2845 5845 2855
rect 5805 2815 5810 2845
rect 5840 2815 5845 2845
rect 6005 2845 6045 2855
rect 6005 2815 6010 2845
rect 6040 2815 6045 2845
rect 6205 2845 6245 2855
rect 6205 2815 6210 2845
rect 6240 2815 6245 2845
rect 6405 2845 6445 2855
rect 6405 2815 6410 2845
rect 6440 2815 6445 2845
rect -188 2730 -185 2815
rect -165 2730 -162 2815
rect 15 2730 35 2815
rect 215 2730 235 2815
rect 415 2730 435 2815
rect 615 2730 635 2815
rect 815 2730 835 2815
rect 1015 2730 1035 2815
rect 1215 2730 1235 2815
rect 1415 2730 1435 2815
rect 1615 2730 1635 2815
rect 1815 2730 1835 2815
rect 2015 2730 2035 2815
rect 2215 2730 2235 2815
rect 2415 2730 2435 2815
rect 2615 2730 2635 2815
rect 2815 2730 2835 2815
rect 3015 2730 3035 2815
rect 3215 2730 3235 2815
rect 3415 2730 3435 2815
rect 3615 2730 3635 2815
rect 3815 2730 3835 2815
rect 4015 2730 4035 2815
rect 4215 2730 4235 2815
rect 4415 2730 4435 2815
rect 4615 2730 4635 2815
rect 4815 2730 4835 2815
rect 5015 2730 5035 2815
rect 5215 2730 5235 2815
rect 5415 2730 5435 2815
rect 5615 2730 5635 2815
rect 5815 2730 5835 2815
rect 6015 2730 6035 2815
rect 6215 2730 6235 2815
rect -195 2700 -190 2730
rect -160 2700 -155 2730
rect -195 2660 -185 2700
rect -165 2690 -155 2700
rect 5 2700 10 2730
rect 40 2700 45 2730
rect 5 2690 45 2700
rect 205 2700 210 2730
rect 240 2700 245 2730
rect 205 2690 245 2700
rect 405 2700 410 2730
rect 440 2700 445 2730
rect 405 2690 445 2700
rect 605 2700 610 2730
rect 640 2700 645 2730
rect 605 2690 645 2700
rect 805 2700 810 2730
rect 840 2700 845 2730
rect 805 2690 845 2700
rect 1005 2700 1010 2730
rect 1040 2700 1045 2730
rect 1005 2690 1045 2700
rect 1205 2700 1210 2730
rect 1240 2700 1245 2730
rect 1205 2690 1245 2700
rect 1405 2700 1410 2730
rect 1440 2700 1445 2730
rect 1405 2690 1445 2700
rect 1605 2700 1610 2730
rect 1640 2700 1645 2730
rect 1605 2690 1645 2700
rect 1805 2700 1810 2730
rect 1840 2700 1845 2730
rect 1805 2690 1845 2700
rect 2005 2700 2010 2730
rect 2040 2700 2045 2730
rect 2005 2690 2045 2700
rect 2205 2700 2210 2730
rect 2240 2700 2245 2730
rect 2205 2690 2245 2700
rect 2405 2700 2410 2730
rect 2440 2700 2445 2730
rect 2405 2690 2445 2700
rect 2605 2700 2610 2730
rect 2640 2700 2645 2730
rect 2605 2690 2645 2700
rect 2805 2700 2810 2730
rect 2840 2700 2845 2730
rect 2805 2690 2845 2700
rect 3005 2700 3010 2730
rect 3040 2700 3045 2730
rect 3005 2690 3045 2700
rect 3205 2700 3210 2730
rect 3240 2700 3245 2730
rect 3205 2690 3245 2700
rect 3405 2700 3410 2730
rect 3440 2700 3445 2730
rect 3405 2690 3445 2700
rect 3605 2700 3610 2730
rect 3640 2700 3645 2730
rect 3605 2690 3645 2700
rect 3805 2700 3810 2730
rect 3840 2700 3845 2730
rect 3805 2690 3845 2700
rect 4005 2700 4010 2730
rect 4040 2700 4045 2730
rect 4005 2690 4045 2700
rect 4205 2700 4210 2730
rect 4240 2700 4245 2730
rect 4205 2690 4245 2700
rect 4405 2700 4410 2730
rect 4440 2700 4445 2730
rect 4405 2690 4445 2700
rect 4605 2700 4610 2730
rect 4640 2700 4645 2730
rect 4605 2690 4645 2700
rect 4805 2700 4810 2730
rect 4840 2700 4845 2730
rect 4805 2690 4845 2700
rect 5005 2700 5010 2730
rect 5040 2700 5045 2730
rect 5005 2690 5045 2700
rect 5205 2700 5210 2730
rect 5240 2700 5245 2730
rect 5205 2690 5245 2700
rect 5405 2700 5410 2730
rect 5440 2700 5445 2730
rect 5405 2690 5445 2700
rect 5605 2700 5610 2730
rect 5640 2700 5645 2730
rect 5605 2690 5645 2700
rect 5805 2700 5810 2730
rect 5840 2700 5845 2730
rect 5805 2690 5845 2700
rect 6005 2700 6010 2730
rect 6040 2700 6045 2730
rect 6005 2690 6045 2700
rect 6205 2700 6210 2730
rect 6240 2700 6245 2730
rect 6205 2690 6245 2700
rect 6405 2700 6410 2730
rect 6440 2700 6445 2730
rect 6405 2690 6445 2700
rect -165 2670 -30 2690
rect 5 2670 1570 2690
rect 1605 2670 6570 2690
rect -165 2660 -155 2670
rect -195 2630 -190 2660
rect -160 2630 -155 2660
rect 5 2660 45 2670
rect 5 2630 10 2660
rect 40 2630 45 2660
rect 205 2660 245 2670
rect 205 2630 210 2660
rect 240 2630 245 2660
rect 405 2660 445 2670
rect 405 2630 410 2660
rect 440 2630 445 2660
rect 605 2660 645 2670
rect 605 2630 610 2660
rect 640 2630 645 2660
rect 805 2660 845 2670
rect 805 2630 810 2660
rect 840 2630 845 2660
rect 1005 2660 1045 2670
rect 1005 2630 1010 2660
rect 1040 2630 1045 2660
rect 1205 2660 1245 2670
rect 1205 2630 1210 2660
rect 1240 2630 1245 2660
rect 1405 2660 1445 2670
rect 1405 2630 1410 2660
rect 1440 2630 1445 2660
rect 1605 2660 1645 2670
rect 1605 2630 1610 2660
rect 1640 2630 1645 2660
rect 1805 2660 1845 2670
rect 1805 2630 1810 2660
rect 1840 2630 1845 2660
rect 2005 2660 2045 2670
rect 2005 2630 2010 2660
rect 2040 2630 2045 2660
rect 2205 2660 2245 2670
rect 2205 2630 2210 2660
rect 2240 2630 2245 2660
rect 2405 2660 2445 2670
rect 2405 2630 2410 2660
rect 2440 2630 2445 2660
rect 2605 2660 2645 2670
rect 2605 2630 2610 2660
rect 2640 2630 2645 2660
rect 2805 2660 2845 2670
rect 2805 2630 2810 2660
rect 2840 2630 2845 2660
rect 3005 2660 3045 2670
rect 3005 2630 3010 2660
rect 3040 2630 3045 2660
rect 3205 2660 3245 2670
rect 3205 2630 3210 2660
rect 3240 2630 3245 2660
rect 3405 2660 3445 2670
rect 3405 2630 3410 2660
rect 3440 2630 3445 2660
rect 3605 2660 3645 2670
rect 3605 2630 3610 2660
rect 3640 2630 3645 2660
rect 3805 2660 3845 2670
rect 3805 2630 3810 2660
rect 3840 2630 3845 2660
rect 4005 2660 4045 2670
rect 4005 2630 4010 2660
rect 4040 2630 4045 2660
rect 4205 2660 4245 2670
rect 4205 2630 4210 2660
rect 4240 2630 4245 2660
rect 4405 2660 4445 2670
rect 4405 2630 4410 2660
rect 4440 2630 4445 2660
rect 4605 2660 4645 2670
rect 4605 2630 4610 2660
rect 4640 2630 4645 2660
rect 4805 2660 4845 2670
rect 4805 2630 4810 2660
rect 4840 2630 4845 2660
rect 5005 2660 5045 2670
rect 5005 2630 5010 2660
rect 5040 2630 5045 2660
rect 5205 2660 5245 2670
rect 5205 2630 5210 2660
rect 5240 2630 5245 2660
rect 5405 2660 5445 2670
rect 5405 2630 5410 2660
rect 5440 2630 5445 2660
rect 5605 2660 5645 2670
rect 5605 2630 5610 2660
rect 5640 2630 5645 2660
rect 5805 2660 5845 2670
rect 5805 2630 5810 2660
rect 5840 2630 5845 2660
rect 6005 2660 6045 2670
rect 6005 2630 6010 2660
rect 6040 2630 6045 2660
rect 6205 2660 6245 2670
rect 6205 2630 6210 2660
rect 6240 2630 6245 2660
rect 6405 2660 6445 2670
rect 6405 2630 6410 2660
rect 6440 2630 6445 2660
rect -188 2545 -185 2630
rect -165 2545 -162 2630
rect 15 2545 35 2630
rect 215 2545 235 2630
rect 415 2545 435 2630
rect 615 2545 635 2630
rect 815 2545 835 2630
rect 1015 2545 1035 2630
rect 1215 2545 1235 2630
rect 1415 2545 1435 2630
rect 1615 2545 1635 2630
rect 1815 2545 1835 2630
rect 2015 2545 2035 2630
rect 2215 2545 2235 2630
rect 2415 2545 2435 2630
rect 2615 2545 2635 2630
rect 2815 2545 2835 2630
rect 3015 2545 3035 2630
rect 3215 2545 3235 2630
rect 3415 2545 3435 2630
rect 3615 2545 3635 2630
rect 3815 2545 3835 2630
rect 4015 2545 4035 2630
rect 4215 2545 4235 2630
rect 4415 2545 4435 2630
rect 4615 2545 4635 2630
rect 4815 2545 4835 2630
rect 5015 2545 5035 2630
rect 5215 2545 5235 2630
rect 5415 2545 5435 2630
rect 5615 2545 5635 2630
rect 5815 2545 5835 2630
rect 6015 2545 6035 2630
rect 6215 2545 6235 2630
rect -195 2515 -190 2545
rect -160 2515 -155 2545
rect -195 2475 -185 2515
rect -165 2505 -155 2515
rect 5 2515 10 2545
rect 40 2515 45 2545
rect 5 2505 45 2515
rect 205 2515 210 2545
rect 240 2515 245 2545
rect 205 2505 245 2515
rect 405 2515 410 2545
rect 440 2515 445 2545
rect 405 2505 445 2515
rect 605 2515 610 2545
rect 640 2515 645 2545
rect 605 2505 645 2515
rect 805 2515 810 2545
rect 840 2515 845 2545
rect 805 2505 845 2515
rect 1005 2515 1010 2545
rect 1040 2515 1045 2545
rect 1005 2505 1045 2515
rect 1205 2515 1210 2545
rect 1240 2515 1245 2545
rect 1205 2505 1245 2515
rect 1405 2515 1410 2545
rect 1440 2515 1445 2545
rect 1405 2505 1445 2515
rect 1605 2515 1610 2545
rect 1640 2515 1645 2545
rect 1605 2505 1645 2515
rect 1805 2515 1810 2545
rect 1840 2515 1845 2545
rect 1805 2505 1845 2515
rect 2005 2515 2010 2545
rect 2040 2515 2045 2545
rect 2005 2505 2045 2515
rect 2205 2515 2210 2545
rect 2240 2515 2245 2545
rect 2205 2505 2245 2515
rect 2405 2515 2410 2545
rect 2440 2515 2445 2545
rect 2405 2505 2445 2515
rect 2605 2515 2610 2545
rect 2640 2515 2645 2545
rect 2605 2505 2645 2515
rect 2805 2515 2810 2545
rect 2840 2515 2845 2545
rect 2805 2505 2845 2515
rect 3005 2515 3010 2545
rect 3040 2515 3045 2545
rect 3005 2505 3045 2515
rect 3205 2515 3210 2545
rect 3240 2515 3245 2545
rect 3205 2505 3245 2515
rect 3405 2515 3410 2545
rect 3440 2515 3445 2545
rect 3405 2505 3445 2515
rect 3605 2515 3610 2545
rect 3640 2515 3645 2545
rect 3605 2505 3645 2515
rect 3805 2515 3810 2545
rect 3840 2515 3845 2545
rect 3805 2505 3845 2515
rect 4005 2515 4010 2545
rect 4040 2515 4045 2545
rect 4005 2505 4045 2515
rect 4205 2515 4210 2545
rect 4240 2515 4245 2545
rect 4205 2505 4245 2515
rect 4405 2515 4410 2545
rect 4440 2515 4445 2545
rect 4405 2505 4445 2515
rect 4605 2515 4610 2545
rect 4640 2515 4645 2545
rect 4605 2505 4645 2515
rect 4805 2515 4810 2545
rect 4840 2515 4845 2545
rect 4805 2505 4845 2515
rect 5005 2515 5010 2545
rect 5040 2515 5045 2545
rect 5005 2505 5045 2515
rect 5205 2515 5210 2545
rect 5240 2515 5245 2545
rect 5205 2505 5245 2515
rect 5405 2515 5410 2545
rect 5440 2515 5445 2545
rect 5405 2505 5445 2515
rect 5605 2515 5610 2545
rect 5640 2515 5645 2545
rect 5605 2505 5645 2515
rect 5805 2515 5810 2545
rect 5840 2515 5845 2545
rect 5805 2505 5845 2515
rect 6005 2515 6010 2545
rect 6040 2515 6045 2545
rect 6005 2505 6045 2515
rect 6205 2515 6210 2545
rect 6240 2515 6245 2545
rect 6205 2505 6245 2515
rect 6405 2515 6410 2545
rect 6440 2515 6445 2545
rect 6405 2505 6445 2515
rect -165 2485 -30 2505
rect 5 2485 1570 2505
rect 1605 2485 6570 2505
rect -165 2475 -155 2485
rect -195 2445 -190 2475
rect -160 2445 -155 2475
rect 5 2475 45 2485
rect 5 2445 10 2475
rect 40 2445 45 2475
rect 205 2475 245 2485
rect 205 2445 210 2475
rect 240 2445 245 2475
rect 405 2475 445 2485
rect 405 2445 410 2475
rect 440 2445 445 2475
rect 605 2475 645 2485
rect 605 2445 610 2475
rect 640 2445 645 2475
rect 805 2475 845 2485
rect 805 2445 810 2475
rect 840 2445 845 2475
rect 1005 2475 1045 2485
rect 1005 2445 1010 2475
rect 1040 2445 1045 2475
rect 1205 2475 1245 2485
rect 1205 2445 1210 2475
rect 1240 2445 1245 2475
rect 1405 2475 1445 2485
rect 1405 2445 1410 2475
rect 1440 2445 1445 2475
rect 1605 2475 1645 2485
rect 1605 2445 1610 2475
rect 1640 2445 1645 2475
rect 1805 2475 1845 2485
rect 1805 2445 1810 2475
rect 1840 2445 1845 2475
rect 2005 2475 2045 2485
rect 2005 2445 2010 2475
rect 2040 2445 2045 2475
rect 2205 2475 2245 2485
rect 2205 2445 2210 2475
rect 2240 2445 2245 2475
rect 2405 2475 2445 2485
rect 2405 2445 2410 2475
rect 2440 2445 2445 2475
rect 2605 2475 2645 2485
rect 2605 2445 2610 2475
rect 2640 2445 2645 2475
rect 2805 2475 2845 2485
rect 2805 2445 2810 2475
rect 2840 2445 2845 2475
rect 3005 2475 3045 2485
rect 3005 2445 3010 2475
rect 3040 2445 3045 2475
rect 3205 2475 3245 2485
rect 3205 2445 3210 2475
rect 3240 2445 3245 2475
rect 3405 2475 3445 2485
rect 3405 2445 3410 2475
rect 3440 2445 3445 2475
rect 3605 2475 3645 2485
rect 3605 2445 3610 2475
rect 3640 2445 3645 2475
rect 3805 2475 3845 2485
rect 3805 2445 3810 2475
rect 3840 2445 3845 2475
rect 4005 2475 4045 2485
rect 4005 2445 4010 2475
rect 4040 2445 4045 2475
rect 4205 2475 4245 2485
rect 4205 2445 4210 2475
rect 4240 2445 4245 2475
rect 4405 2475 4445 2485
rect 4405 2445 4410 2475
rect 4440 2445 4445 2475
rect 4605 2475 4645 2485
rect 4605 2445 4610 2475
rect 4640 2445 4645 2475
rect 4805 2475 4845 2485
rect 4805 2445 4810 2475
rect 4840 2445 4845 2475
rect 5005 2475 5045 2485
rect 5005 2445 5010 2475
rect 5040 2445 5045 2475
rect 5205 2475 5245 2485
rect 5205 2445 5210 2475
rect 5240 2445 5245 2475
rect 5405 2475 5445 2485
rect 5405 2445 5410 2475
rect 5440 2445 5445 2475
rect 5605 2475 5645 2485
rect 5605 2445 5610 2475
rect 5640 2445 5645 2475
rect 5805 2475 5845 2485
rect 5805 2445 5810 2475
rect 5840 2445 5845 2475
rect 6005 2475 6045 2485
rect 6005 2445 6010 2475
rect 6040 2445 6045 2475
rect 6205 2475 6245 2485
rect 6205 2445 6210 2475
rect 6240 2445 6245 2475
rect 6405 2475 6445 2485
rect 6405 2445 6410 2475
rect 6440 2445 6445 2475
rect -188 2360 -185 2445
rect -165 2360 -162 2445
rect 15 2360 35 2445
rect 215 2360 235 2445
rect 415 2360 435 2445
rect 615 2360 635 2445
rect 815 2360 835 2445
rect 1015 2360 1035 2445
rect 1215 2360 1235 2445
rect 1415 2360 1435 2445
rect 1615 2360 1635 2445
rect 1815 2360 1835 2445
rect 2015 2360 2035 2445
rect 2215 2360 2235 2445
rect 2415 2360 2435 2445
rect 2615 2360 2635 2445
rect 2815 2360 2835 2445
rect 3015 2360 3035 2445
rect 3215 2360 3235 2445
rect 3415 2360 3435 2445
rect 3615 2360 3635 2445
rect 3815 2360 3835 2445
rect 4015 2360 4035 2445
rect 4215 2360 4235 2445
rect 4415 2360 4435 2445
rect 4615 2360 4635 2445
rect 4815 2360 4835 2445
rect 5015 2360 5035 2445
rect 5215 2360 5235 2445
rect 5415 2360 5435 2445
rect 5615 2360 5635 2445
rect 5815 2360 5835 2445
rect 6015 2360 6035 2445
rect 6215 2360 6235 2445
rect -195 2330 -190 2360
rect -160 2330 -155 2360
rect -195 2290 -185 2330
rect -165 2320 -155 2330
rect 5 2330 10 2360
rect 40 2330 45 2360
rect 5 2320 45 2330
rect 205 2330 210 2360
rect 240 2330 245 2360
rect 205 2320 245 2330
rect 405 2330 410 2360
rect 440 2330 445 2360
rect 405 2320 445 2330
rect 605 2330 610 2360
rect 640 2330 645 2360
rect 605 2320 645 2330
rect 805 2330 810 2360
rect 840 2330 845 2360
rect 805 2320 845 2330
rect 1005 2330 1010 2360
rect 1040 2330 1045 2360
rect 1005 2320 1045 2330
rect 1205 2330 1210 2360
rect 1240 2330 1245 2360
rect 1205 2320 1245 2330
rect 1405 2330 1410 2360
rect 1440 2330 1445 2360
rect 1405 2320 1445 2330
rect 1605 2330 1610 2360
rect 1640 2330 1645 2360
rect 1605 2320 1645 2330
rect 1805 2330 1810 2360
rect 1840 2330 1845 2360
rect 1805 2320 1845 2330
rect 2005 2330 2010 2360
rect 2040 2330 2045 2360
rect 2005 2320 2045 2330
rect 2205 2330 2210 2360
rect 2240 2330 2245 2360
rect 2205 2320 2245 2330
rect 2405 2330 2410 2360
rect 2440 2330 2445 2360
rect 2405 2320 2445 2330
rect 2605 2330 2610 2360
rect 2640 2330 2645 2360
rect 2605 2320 2645 2330
rect 2805 2330 2810 2360
rect 2840 2330 2845 2360
rect 2805 2320 2845 2330
rect 3005 2330 3010 2360
rect 3040 2330 3045 2360
rect 3005 2320 3045 2330
rect 3205 2330 3210 2360
rect 3240 2330 3245 2360
rect 3205 2320 3245 2330
rect 3405 2330 3410 2360
rect 3440 2330 3445 2360
rect 3405 2320 3445 2330
rect 3605 2330 3610 2360
rect 3640 2330 3645 2360
rect 3605 2320 3645 2330
rect 3805 2330 3810 2360
rect 3840 2330 3845 2360
rect 3805 2320 3845 2330
rect 4005 2330 4010 2360
rect 4040 2330 4045 2360
rect 4005 2320 4045 2330
rect 4205 2330 4210 2360
rect 4240 2330 4245 2360
rect 4205 2320 4245 2330
rect 4405 2330 4410 2360
rect 4440 2330 4445 2360
rect 4405 2320 4445 2330
rect 4605 2330 4610 2360
rect 4640 2330 4645 2360
rect 4605 2320 4645 2330
rect 4805 2330 4810 2360
rect 4840 2330 4845 2360
rect 4805 2320 4845 2330
rect 5005 2330 5010 2360
rect 5040 2330 5045 2360
rect 5005 2320 5045 2330
rect 5205 2330 5210 2360
rect 5240 2330 5245 2360
rect 5205 2320 5245 2330
rect 5405 2330 5410 2360
rect 5440 2330 5445 2360
rect 5405 2320 5445 2330
rect 5605 2330 5610 2360
rect 5640 2330 5645 2360
rect 5605 2320 5645 2330
rect 5805 2330 5810 2360
rect 5840 2330 5845 2360
rect 5805 2320 5845 2330
rect 6005 2330 6010 2360
rect 6040 2330 6045 2360
rect 6005 2320 6045 2330
rect 6205 2330 6210 2360
rect 6240 2330 6245 2360
rect 6205 2320 6245 2330
rect 6405 2330 6410 2360
rect 6440 2330 6445 2360
rect 6405 2320 6445 2330
rect -165 2300 -30 2320
rect 5 2300 1570 2320
rect 1605 2300 6570 2320
rect -165 2290 -155 2300
rect -195 2260 -190 2290
rect -160 2260 -155 2290
rect 5 2290 45 2300
rect 5 2260 10 2290
rect 40 2260 45 2290
rect 205 2290 245 2300
rect 205 2260 210 2290
rect 240 2260 245 2290
rect 405 2290 445 2300
rect 405 2260 410 2290
rect 440 2260 445 2290
rect 605 2290 645 2300
rect 605 2260 610 2290
rect 640 2260 645 2290
rect 805 2290 845 2300
rect 805 2260 810 2290
rect 840 2260 845 2290
rect 1005 2290 1045 2300
rect 1005 2260 1010 2290
rect 1040 2260 1045 2290
rect 1205 2290 1245 2300
rect 1205 2260 1210 2290
rect 1240 2260 1245 2290
rect 1405 2290 1445 2300
rect 1405 2260 1410 2290
rect 1440 2260 1445 2290
rect 1605 2290 1645 2300
rect 1605 2260 1610 2290
rect 1640 2260 1645 2290
rect 1805 2290 1845 2300
rect 1805 2260 1810 2290
rect 1840 2260 1845 2290
rect 2005 2290 2045 2300
rect 2005 2260 2010 2290
rect 2040 2260 2045 2290
rect 2205 2290 2245 2300
rect 2205 2260 2210 2290
rect 2240 2260 2245 2290
rect 2405 2290 2445 2300
rect 2405 2260 2410 2290
rect 2440 2260 2445 2290
rect 2605 2290 2645 2300
rect 2605 2260 2610 2290
rect 2640 2260 2645 2290
rect 2805 2290 2845 2300
rect 2805 2260 2810 2290
rect 2840 2260 2845 2290
rect 3005 2290 3045 2300
rect 3005 2260 3010 2290
rect 3040 2260 3045 2290
rect 3205 2290 3245 2300
rect 3205 2260 3210 2290
rect 3240 2260 3245 2290
rect 3405 2290 3445 2300
rect 3405 2260 3410 2290
rect 3440 2260 3445 2290
rect 3605 2290 3645 2300
rect 3605 2260 3610 2290
rect 3640 2260 3645 2290
rect 3805 2290 3845 2300
rect 3805 2260 3810 2290
rect 3840 2260 3845 2290
rect 4005 2290 4045 2300
rect 4005 2260 4010 2290
rect 4040 2260 4045 2290
rect 4205 2290 4245 2300
rect 4205 2260 4210 2290
rect 4240 2260 4245 2290
rect 4405 2290 4445 2300
rect 4405 2260 4410 2290
rect 4440 2260 4445 2290
rect 4605 2290 4645 2300
rect 4605 2260 4610 2290
rect 4640 2260 4645 2290
rect 4805 2290 4845 2300
rect 4805 2260 4810 2290
rect 4840 2260 4845 2290
rect 5005 2290 5045 2300
rect 5005 2260 5010 2290
rect 5040 2260 5045 2290
rect 5205 2290 5245 2300
rect 5205 2260 5210 2290
rect 5240 2260 5245 2290
rect 5405 2290 5445 2300
rect 5405 2260 5410 2290
rect 5440 2260 5445 2290
rect 5605 2290 5645 2300
rect 5605 2260 5610 2290
rect 5640 2260 5645 2290
rect 5805 2290 5845 2300
rect 5805 2260 5810 2290
rect 5840 2260 5845 2290
rect 6005 2290 6045 2300
rect 6005 2260 6010 2290
rect 6040 2260 6045 2290
rect 6205 2290 6245 2300
rect 6205 2260 6210 2290
rect 6240 2260 6245 2290
rect 6405 2290 6445 2300
rect 6405 2260 6410 2290
rect 6440 2260 6445 2290
rect -188 2175 -185 2260
rect -165 2175 -162 2260
rect 15 2175 35 2260
rect 215 2175 235 2260
rect 415 2175 435 2260
rect 615 2175 635 2260
rect 815 2175 835 2260
rect 1015 2175 1035 2260
rect 1215 2175 1235 2260
rect 1415 2175 1435 2260
rect 1615 2175 1635 2260
rect 1815 2175 1835 2260
rect 2015 2175 2035 2260
rect 2215 2175 2235 2260
rect 2415 2175 2435 2260
rect 2615 2175 2635 2260
rect 2815 2175 2835 2260
rect 3015 2175 3035 2260
rect 3215 2175 3235 2260
rect 3415 2175 3435 2260
rect 3615 2175 3635 2260
rect 3815 2175 3835 2260
rect 4015 2175 4035 2260
rect 4215 2175 4235 2260
rect 4415 2175 4435 2260
rect 4615 2175 4635 2260
rect 4815 2175 4835 2260
rect 5015 2175 5035 2260
rect 5215 2175 5235 2260
rect 5415 2175 5435 2260
rect 5615 2175 5635 2260
rect 5815 2175 5835 2260
rect 6015 2175 6035 2260
rect 6215 2175 6235 2260
rect -195 2145 -190 2175
rect -160 2145 -155 2175
rect -195 2105 -185 2145
rect -165 2135 -155 2145
rect 5 2145 10 2175
rect 40 2145 45 2175
rect 5 2135 45 2145
rect 205 2145 210 2175
rect 240 2145 245 2175
rect 205 2135 245 2145
rect 405 2145 410 2175
rect 440 2145 445 2175
rect 405 2135 445 2145
rect 605 2145 610 2175
rect 640 2145 645 2175
rect 605 2135 645 2145
rect 805 2145 810 2175
rect 840 2145 845 2175
rect 805 2135 845 2145
rect 1005 2145 1010 2175
rect 1040 2145 1045 2175
rect 1005 2135 1045 2145
rect 1205 2145 1210 2175
rect 1240 2145 1245 2175
rect 1205 2135 1245 2145
rect 1405 2145 1410 2175
rect 1440 2145 1445 2175
rect 1405 2135 1445 2145
rect 1605 2145 1610 2175
rect 1640 2145 1645 2175
rect 1605 2135 1645 2145
rect 1805 2145 1810 2175
rect 1840 2145 1845 2175
rect 1805 2135 1845 2145
rect 2005 2145 2010 2175
rect 2040 2145 2045 2175
rect 2005 2135 2045 2145
rect 2205 2145 2210 2175
rect 2240 2145 2245 2175
rect 2205 2135 2245 2145
rect 2405 2145 2410 2175
rect 2440 2145 2445 2175
rect 2405 2135 2445 2145
rect 2605 2145 2610 2175
rect 2640 2145 2645 2175
rect 2605 2135 2645 2145
rect 2805 2145 2810 2175
rect 2840 2145 2845 2175
rect 2805 2135 2845 2145
rect 3005 2145 3010 2175
rect 3040 2145 3045 2175
rect 3005 2135 3045 2145
rect 3205 2145 3210 2175
rect 3240 2145 3245 2175
rect 3205 2135 3245 2145
rect 3405 2145 3410 2175
rect 3440 2145 3445 2175
rect 3405 2135 3445 2145
rect 3605 2145 3610 2175
rect 3640 2145 3645 2175
rect 3605 2135 3645 2145
rect 3805 2145 3810 2175
rect 3840 2145 3845 2175
rect 3805 2135 3845 2145
rect 4005 2145 4010 2175
rect 4040 2145 4045 2175
rect 4005 2135 4045 2145
rect 4205 2145 4210 2175
rect 4240 2145 4245 2175
rect 4205 2135 4245 2145
rect 4405 2145 4410 2175
rect 4440 2145 4445 2175
rect 4405 2135 4445 2145
rect 4605 2145 4610 2175
rect 4640 2145 4645 2175
rect 4605 2135 4645 2145
rect 4805 2145 4810 2175
rect 4840 2145 4845 2175
rect 4805 2135 4845 2145
rect 5005 2145 5010 2175
rect 5040 2145 5045 2175
rect 5005 2135 5045 2145
rect 5205 2145 5210 2175
rect 5240 2145 5245 2175
rect 5205 2135 5245 2145
rect 5405 2145 5410 2175
rect 5440 2145 5445 2175
rect 5405 2135 5445 2145
rect 5605 2145 5610 2175
rect 5640 2145 5645 2175
rect 5605 2135 5645 2145
rect 5805 2145 5810 2175
rect 5840 2145 5845 2175
rect 5805 2135 5845 2145
rect 6005 2145 6010 2175
rect 6040 2145 6045 2175
rect 6005 2135 6045 2145
rect 6205 2145 6210 2175
rect 6240 2145 6245 2175
rect 6205 2135 6245 2145
rect 6405 2145 6410 2175
rect 6440 2145 6445 2175
rect 6405 2135 6445 2145
rect -165 2115 -30 2135
rect 5 2115 1570 2135
rect 1605 2115 6570 2135
rect -165 2105 -155 2115
rect -195 2075 -190 2105
rect -160 2075 -155 2105
rect 5 2105 45 2115
rect 5 2075 10 2105
rect 40 2075 45 2105
rect 205 2105 245 2115
rect 205 2075 210 2105
rect 240 2075 245 2105
rect 405 2105 445 2115
rect 405 2075 410 2105
rect 440 2075 445 2105
rect 605 2105 645 2115
rect 605 2075 610 2105
rect 640 2075 645 2105
rect 805 2105 845 2115
rect 805 2075 810 2105
rect 840 2075 845 2105
rect 1005 2105 1045 2115
rect 1005 2075 1010 2105
rect 1040 2075 1045 2105
rect 1205 2105 1245 2115
rect 1205 2075 1210 2105
rect 1240 2075 1245 2105
rect 1405 2105 1445 2115
rect 1405 2075 1410 2105
rect 1440 2075 1445 2105
rect 1605 2105 1645 2115
rect 1605 2075 1610 2105
rect 1640 2075 1645 2105
rect 1805 2105 1845 2115
rect 1805 2075 1810 2105
rect 1840 2075 1845 2105
rect 2005 2105 2045 2115
rect 2005 2075 2010 2105
rect 2040 2075 2045 2105
rect 2205 2105 2245 2115
rect 2205 2075 2210 2105
rect 2240 2075 2245 2105
rect 2405 2105 2445 2115
rect 2405 2075 2410 2105
rect 2440 2075 2445 2105
rect 2605 2105 2645 2115
rect 2605 2075 2610 2105
rect 2640 2075 2645 2105
rect 2805 2105 2845 2115
rect 2805 2075 2810 2105
rect 2840 2075 2845 2105
rect 3005 2105 3045 2115
rect 3005 2075 3010 2105
rect 3040 2075 3045 2105
rect 3205 2105 3245 2115
rect 3205 2075 3210 2105
rect 3240 2075 3245 2105
rect 3405 2105 3445 2115
rect 3405 2075 3410 2105
rect 3440 2075 3445 2105
rect 3605 2105 3645 2115
rect 3605 2075 3610 2105
rect 3640 2075 3645 2105
rect 3805 2105 3845 2115
rect 3805 2075 3810 2105
rect 3840 2075 3845 2105
rect 4005 2105 4045 2115
rect 4005 2075 4010 2105
rect 4040 2075 4045 2105
rect 4205 2105 4245 2115
rect 4205 2075 4210 2105
rect 4240 2075 4245 2105
rect 4405 2105 4445 2115
rect 4405 2075 4410 2105
rect 4440 2075 4445 2105
rect 4605 2105 4645 2115
rect 4605 2075 4610 2105
rect 4640 2075 4645 2105
rect 4805 2105 4845 2115
rect 4805 2075 4810 2105
rect 4840 2075 4845 2105
rect 5005 2105 5045 2115
rect 5005 2075 5010 2105
rect 5040 2075 5045 2105
rect 5205 2105 5245 2115
rect 5205 2075 5210 2105
rect 5240 2075 5245 2105
rect 5405 2105 5445 2115
rect 5405 2075 5410 2105
rect 5440 2075 5445 2105
rect 5605 2105 5645 2115
rect 5605 2075 5610 2105
rect 5640 2075 5645 2105
rect 5805 2105 5845 2115
rect 5805 2075 5810 2105
rect 5840 2075 5845 2105
rect 6005 2105 6045 2115
rect 6005 2075 6010 2105
rect 6040 2075 6045 2105
rect 6205 2105 6245 2115
rect 6205 2075 6210 2105
rect 6240 2075 6245 2105
rect 6405 2105 6445 2115
rect 6405 2075 6410 2105
rect 6440 2075 6445 2105
rect -188 1990 -185 2075
rect -165 1990 -162 2075
rect 15 1990 35 2075
rect 215 1990 235 2075
rect 415 1990 435 2075
rect 615 1990 635 2075
rect 815 1990 835 2075
rect 1015 1990 1035 2075
rect 1215 1990 1235 2075
rect 1415 1990 1435 2075
rect -195 1960 -190 1990
rect -160 1960 -155 1990
rect -195 1920 -185 1960
rect -165 1950 -155 1960
rect 5 1960 10 1990
rect 40 1960 45 1990
rect 5 1950 45 1960
rect 205 1960 210 1990
rect 240 1960 245 1990
rect 205 1950 245 1960
rect 405 1960 410 1990
rect 440 1960 445 1990
rect 405 1950 445 1960
rect 605 1960 610 1990
rect 640 1960 645 1990
rect 605 1950 645 1960
rect 805 1960 810 1990
rect 840 1960 845 1990
rect 805 1950 845 1960
rect 1005 1960 1010 1990
rect 1040 1960 1045 1990
rect 1005 1950 1045 1960
rect 1205 1960 1210 1990
rect 1240 1960 1245 1990
rect 1205 1950 1245 1960
rect 1405 1960 1410 1990
rect 1440 1960 1445 1990
rect 1405 1950 1445 1960
rect 1605 1960 1610 1990
rect 1640 1960 1645 1990
rect 1605 1950 1645 1960
rect 1805 1960 1810 1990
rect 1840 1960 1845 1990
rect 1805 1950 1845 1960
rect 2005 1960 2010 1990
rect 2040 1960 2045 1990
rect 2005 1950 2045 1960
rect 2205 1960 2210 1990
rect 2240 1960 2245 1990
rect 2205 1950 2245 1960
rect 2405 1960 2410 1990
rect 2440 1960 2445 1990
rect 2405 1950 2445 1960
rect 2605 1960 2610 1990
rect 2640 1960 2645 1990
rect 2605 1950 2645 1960
rect 2805 1960 2810 1990
rect 2840 1960 2845 1990
rect 2805 1950 2845 1960
rect 3005 1960 3010 1990
rect 3040 1960 3045 1990
rect 3005 1950 3045 1960
rect 3205 1960 3210 1990
rect 3240 1960 3245 1990
rect 3205 1950 3245 1960
rect 3405 1960 3410 1990
rect 3440 1960 3445 1990
rect 3405 1950 3445 1960
rect 3605 1960 3610 1990
rect 3640 1960 3645 1990
rect 3605 1950 3645 1960
rect 3805 1960 3810 1990
rect 3840 1960 3845 1990
rect 3805 1950 3845 1960
rect 4005 1960 4010 1990
rect 4040 1960 4045 1990
rect 4005 1950 4045 1960
rect 4205 1960 4210 1990
rect 4240 1960 4245 1990
rect 4205 1950 4245 1960
rect 4405 1960 4410 1990
rect 4440 1960 4445 1990
rect 4405 1950 4445 1960
rect 4605 1960 4610 1990
rect 4640 1960 4645 1990
rect 4605 1950 4645 1960
rect 4805 1960 4810 1990
rect 4840 1960 4845 1990
rect 4805 1950 4845 1960
rect 5005 1960 5010 1990
rect 5040 1960 5045 1990
rect 5005 1950 5045 1960
rect 5205 1960 5210 1990
rect 5240 1960 5245 1990
rect 5205 1950 5245 1960
rect 5405 1960 5410 1990
rect 5440 1960 5445 1990
rect 5405 1950 5445 1960
rect 5605 1960 5610 1990
rect 5640 1960 5645 1990
rect 5605 1950 5645 1960
rect 5805 1960 5810 1990
rect 5840 1960 5845 1990
rect 5805 1950 5845 1960
rect 6005 1960 6010 1990
rect 6040 1960 6045 1990
rect 6005 1950 6045 1960
rect 6205 1960 6210 1990
rect 6240 1960 6245 1990
rect 6205 1950 6245 1960
rect 6405 1960 6410 1990
rect 6440 1960 6445 1990
rect 6405 1950 6445 1960
rect -165 1930 -30 1950
rect 5 1930 6695 1950
rect -165 1920 -155 1930
rect -195 1890 -190 1920
rect -160 1890 -155 1920
rect 5 1920 45 1930
rect 5 1890 10 1920
rect 40 1890 45 1920
rect 205 1920 245 1930
rect 205 1890 210 1920
rect 240 1890 245 1920
rect 405 1920 445 1930
rect 405 1890 410 1920
rect 440 1890 445 1920
rect 605 1920 645 1930
rect 605 1890 610 1920
rect 640 1890 645 1920
rect 805 1920 845 1930
rect 805 1890 810 1920
rect 840 1890 845 1920
rect 1005 1920 1045 1930
rect 1005 1890 1010 1920
rect 1040 1890 1045 1920
rect 1205 1920 1245 1930
rect 1205 1890 1210 1920
rect 1240 1890 1245 1920
rect 1405 1920 1445 1930
rect 1405 1890 1410 1920
rect 1440 1890 1445 1920
rect 1605 1920 1645 1930
rect 1605 1890 1610 1920
rect 1640 1890 1645 1920
rect 1805 1920 1845 1930
rect 1805 1890 1810 1920
rect 1840 1890 1845 1920
rect 2005 1920 2045 1930
rect 2005 1890 2010 1920
rect 2040 1890 2045 1920
rect 2205 1920 2245 1930
rect 2205 1890 2210 1920
rect 2240 1890 2245 1920
rect 2405 1920 2445 1930
rect 2405 1890 2410 1920
rect 2440 1890 2445 1920
rect 2605 1920 2645 1930
rect 2605 1890 2610 1920
rect 2640 1890 2645 1920
rect 2805 1920 2845 1930
rect 2805 1890 2810 1920
rect 2840 1890 2845 1920
rect 3005 1920 3045 1930
rect 3005 1890 3010 1920
rect 3040 1890 3045 1920
rect 3205 1920 3245 1930
rect 3205 1890 3210 1920
rect 3240 1890 3245 1920
rect 3405 1920 3445 1930
rect 3405 1890 3410 1920
rect 3440 1890 3445 1920
rect 3605 1920 3645 1930
rect 3605 1890 3610 1920
rect 3640 1890 3645 1920
rect 3805 1920 3845 1930
rect 3805 1890 3810 1920
rect 3840 1890 3845 1920
rect 4005 1920 4045 1930
rect 4005 1890 4010 1920
rect 4040 1890 4045 1920
rect 4205 1920 4245 1930
rect 4205 1890 4210 1920
rect 4240 1890 4245 1920
rect 4405 1920 4445 1930
rect 4405 1890 4410 1920
rect 4440 1890 4445 1920
rect 4605 1920 4645 1930
rect 4605 1890 4610 1920
rect 4640 1890 4645 1920
rect 4805 1920 4845 1930
rect 4805 1890 4810 1920
rect 4840 1890 4845 1920
rect 5005 1920 5045 1930
rect 5005 1890 5010 1920
rect 5040 1890 5045 1920
rect 5205 1920 5245 1930
rect 5205 1890 5210 1920
rect 5240 1890 5245 1920
rect 5405 1920 5445 1930
rect 5405 1890 5410 1920
rect 5440 1890 5445 1920
rect 5605 1920 5645 1930
rect 5605 1890 5610 1920
rect 5640 1890 5645 1920
rect 5805 1920 5845 1930
rect 5805 1890 5810 1920
rect 5840 1890 5845 1920
rect 6005 1920 6045 1930
rect 6005 1890 6010 1920
rect 6040 1890 6045 1920
rect 6205 1920 6245 1930
rect 6205 1890 6210 1920
rect 6240 1890 6245 1920
rect 6405 1920 6445 1930
rect 6405 1890 6410 1920
rect 6440 1890 6445 1920
rect -188 1805 -185 1890
rect -165 1805 -162 1890
rect 15 1805 35 1890
rect 215 1805 235 1890
rect 415 1805 435 1890
rect 615 1805 635 1890
rect 815 1805 835 1890
rect 1015 1805 1035 1890
rect 1215 1805 1235 1890
rect 1415 1805 1435 1890
rect 1615 1805 1635 1890
rect 1815 1805 1835 1890
rect 2015 1805 2035 1890
rect 2215 1805 2235 1890
rect 2415 1805 2435 1890
rect 2615 1805 2635 1890
rect 2815 1805 2835 1890
rect 3015 1805 3035 1890
rect 3215 1805 3235 1890
rect 3415 1805 3435 1890
rect 3615 1805 3635 1890
rect 3815 1805 3835 1890
rect 4015 1805 4035 1890
rect 4215 1805 4235 1890
rect 4415 1805 4435 1890
rect 4615 1805 4635 1890
rect 4815 1805 4835 1890
rect 5015 1805 5035 1890
rect 5215 1805 5235 1890
rect 5415 1805 5435 1890
rect 5615 1805 5635 1890
rect 5815 1805 5835 1890
rect 6015 1805 6035 1890
rect 6215 1805 6235 1890
rect -195 1775 -190 1805
rect -160 1775 -155 1805
rect -195 1735 -185 1775
rect -165 1765 -155 1775
rect 5 1775 10 1805
rect 40 1775 45 1805
rect 5 1765 45 1775
rect 205 1775 210 1805
rect 240 1775 245 1805
rect 205 1765 245 1775
rect 405 1775 410 1805
rect 440 1775 445 1805
rect 405 1765 445 1775
rect 605 1775 610 1805
rect 640 1775 645 1805
rect 605 1765 645 1775
rect 805 1775 810 1805
rect 840 1775 845 1805
rect 805 1765 845 1775
rect 1005 1775 1010 1805
rect 1040 1775 1045 1805
rect 1005 1765 1045 1775
rect 1205 1775 1210 1805
rect 1240 1775 1245 1805
rect 1205 1765 1245 1775
rect 1405 1775 1410 1805
rect 1440 1775 1445 1805
rect 1405 1765 1445 1775
rect 1605 1775 1610 1805
rect 1640 1775 1645 1805
rect 1605 1765 1645 1775
rect 1805 1775 1810 1805
rect 1840 1775 1845 1805
rect 1805 1765 1845 1775
rect 2005 1775 2010 1805
rect 2040 1775 2045 1805
rect 2005 1765 2045 1775
rect 2205 1775 2210 1805
rect 2240 1775 2245 1805
rect 2205 1765 2245 1775
rect 2405 1775 2410 1805
rect 2440 1775 2445 1805
rect 2405 1765 2445 1775
rect 2605 1775 2610 1805
rect 2640 1775 2645 1805
rect 2605 1765 2645 1775
rect 2805 1775 2810 1805
rect 2840 1775 2845 1805
rect 2805 1765 2845 1775
rect 3005 1775 3010 1805
rect 3040 1775 3045 1805
rect 3005 1765 3045 1775
rect 3205 1775 3210 1805
rect 3240 1775 3245 1805
rect 3205 1765 3245 1775
rect 3405 1775 3410 1805
rect 3440 1775 3445 1805
rect 3405 1765 3445 1775
rect 3605 1775 3610 1805
rect 3640 1775 3645 1805
rect 3605 1765 3645 1775
rect 3805 1775 3810 1805
rect 3840 1775 3845 1805
rect 3805 1765 3845 1775
rect 4005 1775 4010 1805
rect 4040 1775 4045 1805
rect 4005 1765 4045 1775
rect 4205 1775 4210 1805
rect 4240 1775 4245 1805
rect 4205 1765 4245 1775
rect 4405 1775 4410 1805
rect 4440 1775 4445 1805
rect 4405 1765 4445 1775
rect 4605 1775 4610 1805
rect 4640 1775 4645 1805
rect 4605 1765 4645 1775
rect 4805 1775 4810 1805
rect 4840 1775 4845 1805
rect 4805 1765 4845 1775
rect 5005 1775 5010 1805
rect 5040 1775 5045 1805
rect 5005 1765 5045 1775
rect 5205 1775 5210 1805
rect 5240 1775 5245 1805
rect 5205 1765 5245 1775
rect 5405 1775 5410 1805
rect 5440 1775 5445 1805
rect 5405 1765 5445 1775
rect 5605 1775 5610 1805
rect 5640 1775 5645 1805
rect 5605 1765 5645 1775
rect 5805 1775 5810 1805
rect 5840 1775 5845 1805
rect 5805 1765 5845 1775
rect 6005 1775 6010 1805
rect 6040 1775 6045 1805
rect 6005 1765 6045 1775
rect 6205 1775 6210 1805
rect 6240 1775 6245 1805
rect 6205 1765 6245 1775
rect 6405 1775 6410 1805
rect 6440 1775 6445 1805
rect 6405 1765 6445 1775
rect -165 1745 -30 1765
rect 5 1745 6570 1765
rect -165 1735 -155 1745
rect -195 1705 -190 1735
rect -160 1705 -155 1735
rect 5 1735 45 1745
rect 5 1705 10 1735
rect 40 1705 45 1735
rect 205 1735 245 1745
rect 205 1705 210 1735
rect 240 1705 245 1735
rect 405 1735 445 1745
rect 405 1705 410 1735
rect 440 1705 445 1735
rect 605 1735 645 1745
rect 605 1705 610 1735
rect 640 1705 645 1735
rect 805 1735 845 1745
rect 805 1705 810 1735
rect 840 1705 845 1735
rect 1005 1735 1045 1745
rect 1005 1705 1010 1735
rect 1040 1705 1045 1735
rect 1205 1735 1245 1745
rect 1205 1705 1210 1735
rect 1240 1705 1245 1735
rect 1405 1735 1445 1745
rect 1405 1705 1410 1735
rect 1440 1705 1445 1735
rect 1605 1735 1645 1745
rect 1605 1705 1610 1735
rect 1640 1705 1645 1735
rect 1805 1735 1845 1745
rect 1805 1705 1810 1735
rect 1840 1705 1845 1735
rect 2005 1735 2045 1745
rect 2005 1705 2010 1735
rect 2040 1705 2045 1735
rect 2205 1735 2245 1745
rect 2205 1705 2210 1735
rect 2240 1705 2245 1735
rect 2405 1735 2445 1745
rect 2405 1705 2410 1735
rect 2440 1705 2445 1735
rect 2605 1735 2645 1745
rect 2605 1705 2610 1735
rect 2640 1705 2645 1735
rect 2805 1735 2845 1745
rect 2805 1705 2810 1735
rect 2840 1705 2845 1735
rect 3005 1735 3045 1745
rect 3005 1705 3010 1735
rect 3040 1705 3045 1735
rect 3205 1735 3245 1745
rect 3205 1705 3210 1735
rect 3240 1705 3245 1735
rect 3405 1735 3445 1745
rect 3405 1705 3410 1735
rect 3440 1705 3445 1735
rect 3605 1735 3645 1745
rect 3605 1705 3610 1735
rect 3640 1705 3645 1735
rect 3805 1735 3845 1745
rect 3805 1705 3810 1735
rect 3840 1705 3845 1735
rect 4005 1735 4045 1745
rect 4005 1705 4010 1735
rect 4040 1705 4045 1735
rect 4205 1735 4245 1745
rect 4205 1705 4210 1735
rect 4240 1705 4245 1735
rect 4405 1735 4445 1745
rect 4405 1705 4410 1735
rect 4440 1705 4445 1735
rect 4605 1735 4645 1745
rect 4605 1705 4610 1735
rect 4640 1705 4645 1735
rect 4805 1735 4845 1745
rect 4805 1705 4810 1735
rect 4840 1705 4845 1735
rect 5005 1735 5045 1745
rect 5005 1705 5010 1735
rect 5040 1705 5045 1735
rect 5205 1735 5245 1745
rect 5205 1705 5210 1735
rect 5240 1705 5245 1735
rect 5405 1735 5445 1745
rect 5405 1705 5410 1735
rect 5440 1705 5445 1735
rect 5605 1735 5645 1745
rect 5605 1705 5610 1735
rect 5640 1705 5645 1735
rect 5805 1735 5845 1745
rect 5805 1705 5810 1735
rect 5840 1705 5845 1735
rect 6005 1735 6045 1745
rect 6005 1705 6010 1735
rect 6040 1705 6045 1735
rect 6205 1735 6245 1745
rect 6205 1705 6210 1735
rect 6240 1705 6245 1735
rect 6405 1735 6445 1745
rect 6405 1705 6410 1735
rect 6440 1705 6445 1735
rect -188 1620 -185 1705
rect -165 1620 -162 1705
rect 15 1620 35 1705
rect 215 1620 235 1705
rect 415 1620 435 1705
rect 615 1620 635 1705
rect 815 1620 835 1705
rect 1015 1620 1035 1705
rect 1215 1620 1235 1705
rect 1415 1620 1435 1705
rect 1615 1620 1635 1705
rect 1815 1620 1835 1705
rect 2015 1620 2035 1705
rect 2215 1620 2235 1705
rect 2415 1620 2435 1705
rect 2615 1620 2635 1705
rect 2815 1620 2835 1705
rect 3015 1620 3035 1705
rect 3215 1620 3235 1705
rect 3415 1620 3435 1705
rect 3615 1620 3635 1705
rect 3815 1620 3835 1705
rect 4015 1620 4035 1705
rect 4215 1620 4235 1705
rect 4415 1620 4435 1705
rect 4615 1620 4635 1705
rect 4815 1620 4835 1705
rect 5015 1620 5035 1705
rect 5215 1620 5235 1705
rect 5415 1620 5435 1705
rect 5615 1620 5635 1705
rect 5815 1620 5835 1705
rect 6015 1620 6035 1705
rect 6215 1620 6235 1705
rect -195 1590 -190 1620
rect -160 1590 -155 1620
rect -195 1550 -185 1590
rect -165 1580 -155 1590
rect 5 1590 10 1620
rect 40 1590 45 1620
rect 5 1580 45 1590
rect 205 1590 210 1620
rect 240 1590 245 1620
rect 205 1580 245 1590
rect 405 1590 410 1620
rect 440 1590 445 1620
rect 405 1580 445 1590
rect 605 1590 610 1620
rect 640 1590 645 1620
rect 605 1580 645 1590
rect 805 1590 810 1620
rect 840 1590 845 1620
rect 805 1580 845 1590
rect 1005 1590 1010 1620
rect 1040 1590 1045 1620
rect 1005 1580 1045 1590
rect 1205 1590 1210 1620
rect 1240 1590 1245 1620
rect 1205 1580 1245 1590
rect 1405 1590 1410 1620
rect 1440 1590 1445 1620
rect 1405 1580 1445 1590
rect 1605 1590 1610 1620
rect 1640 1590 1645 1620
rect 1605 1580 1645 1590
rect 1805 1590 1810 1620
rect 1840 1590 1845 1620
rect 1805 1580 1845 1590
rect 2005 1590 2010 1620
rect 2040 1590 2045 1620
rect 2005 1580 2045 1590
rect 2205 1590 2210 1620
rect 2240 1590 2245 1620
rect 2205 1580 2245 1590
rect 2405 1590 2410 1620
rect 2440 1590 2445 1620
rect 2405 1580 2445 1590
rect 2605 1590 2610 1620
rect 2640 1590 2645 1620
rect 2605 1580 2645 1590
rect 2805 1590 2810 1620
rect 2840 1590 2845 1620
rect 2805 1580 2845 1590
rect 3005 1590 3010 1620
rect 3040 1590 3045 1620
rect 3005 1580 3045 1590
rect 3205 1590 3210 1620
rect 3240 1590 3245 1620
rect 3205 1580 3245 1590
rect 3405 1590 3410 1620
rect 3440 1590 3445 1620
rect 3405 1580 3445 1590
rect 3605 1590 3610 1620
rect 3640 1590 3645 1620
rect 3605 1580 3645 1590
rect 3805 1590 3810 1620
rect 3840 1590 3845 1620
rect 3805 1580 3845 1590
rect 4005 1590 4010 1620
rect 4040 1590 4045 1620
rect 4005 1580 4045 1590
rect 4205 1590 4210 1620
rect 4240 1590 4245 1620
rect 4205 1580 4245 1590
rect 4405 1590 4410 1620
rect 4440 1590 4445 1620
rect 4405 1580 4445 1590
rect 4605 1590 4610 1620
rect 4640 1590 4645 1620
rect 4605 1580 4645 1590
rect 4805 1590 4810 1620
rect 4840 1590 4845 1620
rect 4805 1580 4845 1590
rect 5005 1590 5010 1620
rect 5040 1590 5045 1620
rect 5005 1580 5045 1590
rect 5205 1590 5210 1620
rect 5240 1590 5245 1620
rect 5205 1580 5245 1590
rect 5405 1590 5410 1620
rect 5440 1590 5445 1620
rect 5405 1580 5445 1590
rect 5605 1590 5610 1620
rect 5640 1590 5645 1620
rect 5605 1580 5645 1590
rect 5805 1590 5810 1620
rect 5840 1590 5845 1620
rect 5805 1580 5845 1590
rect 6005 1590 6010 1620
rect 6040 1590 6045 1620
rect 6005 1580 6045 1590
rect 6205 1590 6210 1620
rect 6240 1590 6245 1620
rect 6205 1580 6245 1590
rect 6405 1590 6410 1620
rect 6440 1590 6445 1620
rect 6405 1580 6445 1590
rect -165 1560 -30 1580
rect 5 1560 6570 1580
rect -165 1550 -155 1560
rect -195 1520 -190 1550
rect -160 1520 -155 1550
rect 5 1550 45 1560
rect 5 1520 10 1550
rect 40 1520 45 1550
rect 205 1550 245 1560
rect 205 1520 210 1550
rect 240 1520 245 1550
rect 405 1550 445 1560
rect 405 1520 410 1550
rect 440 1520 445 1550
rect 605 1550 645 1560
rect 605 1520 610 1550
rect 640 1520 645 1550
rect 805 1550 845 1560
rect 805 1520 810 1550
rect 840 1520 845 1550
rect 1005 1550 1045 1560
rect 1005 1520 1010 1550
rect 1040 1520 1045 1550
rect 1205 1550 1245 1560
rect 1205 1520 1210 1550
rect 1240 1520 1245 1550
rect 1405 1550 1445 1560
rect 1405 1520 1410 1550
rect 1440 1520 1445 1550
rect 1605 1550 1645 1560
rect 1605 1520 1610 1550
rect 1640 1520 1645 1550
rect 1805 1550 1845 1560
rect 1805 1520 1810 1550
rect 1840 1520 1845 1550
rect 2005 1550 2045 1560
rect 2005 1520 2010 1550
rect 2040 1520 2045 1550
rect 2205 1550 2245 1560
rect 2205 1520 2210 1550
rect 2240 1520 2245 1550
rect 2405 1550 2445 1560
rect 2405 1520 2410 1550
rect 2440 1520 2445 1550
rect 2605 1550 2645 1560
rect 2605 1520 2610 1550
rect 2640 1520 2645 1550
rect 2805 1550 2845 1560
rect 2805 1520 2810 1550
rect 2840 1520 2845 1550
rect 3005 1550 3045 1560
rect 3005 1520 3010 1550
rect 3040 1520 3045 1550
rect 3205 1550 3245 1560
rect 3205 1520 3210 1550
rect 3240 1520 3245 1550
rect 3405 1550 3445 1560
rect 3405 1520 3410 1550
rect 3440 1520 3445 1550
rect 3605 1550 3645 1560
rect 3605 1520 3610 1550
rect 3640 1520 3645 1550
rect 3805 1550 3845 1560
rect 3805 1520 3810 1550
rect 3840 1520 3845 1550
rect 4005 1550 4045 1560
rect 4005 1520 4010 1550
rect 4040 1520 4045 1550
rect 4205 1550 4245 1560
rect 4205 1520 4210 1550
rect 4240 1520 4245 1550
rect 4405 1550 4445 1560
rect 4405 1520 4410 1550
rect 4440 1520 4445 1550
rect 4605 1550 4645 1560
rect 4605 1520 4610 1550
rect 4640 1520 4645 1550
rect 4805 1550 4845 1560
rect 4805 1520 4810 1550
rect 4840 1520 4845 1550
rect 5005 1550 5045 1560
rect 5005 1520 5010 1550
rect 5040 1520 5045 1550
rect 5205 1550 5245 1560
rect 5205 1520 5210 1550
rect 5240 1520 5245 1550
rect 5405 1550 5445 1560
rect 5405 1520 5410 1550
rect 5440 1520 5445 1550
rect 5605 1550 5645 1560
rect 5605 1520 5610 1550
rect 5640 1520 5645 1550
rect 5805 1550 5845 1560
rect 5805 1520 5810 1550
rect 5840 1520 5845 1550
rect 6005 1550 6045 1560
rect 6005 1520 6010 1550
rect 6040 1520 6045 1550
rect 6205 1550 6245 1560
rect 6205 1520 6210 1550
rect 6240 1520 6245 1550
rect 6405 1550 6445 1560
rect 6405 1520 6410 1550
rect 6440 1520 6445 1550
rect -188 1435 -185 1520
rect -165 1435 -162 1520
rect 15 1435 35 1520
rect 215 1435 235 1520
rect 415 1435 435 1520
rect 615 1435 635 1520
rect 815 1435 835 1520
rect 1015 1435 1035 1520
rect 1215 1435 1235 1520
rect 1415 1435 1435 1520
rect 1615 1435 1635 1520
rect 1815 1435 1835 1520
rect 2015 1435 2035 1520
rect 2215 1435 2235 1520
rect 2415 1435 2435 1520
rect 2615 1435 2635 1520
rect 2815 1435 2835 1520
rect 3015 1435 3035 1520
rect 3215 1435 3235 1520
rect 3415 1435 3435 1520
rect 3615 1435 3635 1520
rect 3815 1435 3835 1520
rect 4015 1435 4035 1520
rect 4215 1435 4235 1520
rect 4415 1435 4435 1520
rect 4615 1435 4635 1520
rect 4815 1435 4835 1520
rect 5015 1435 5035 1520
rect 5215 1435 5235 1520
rect 5415 1435 5435 1520
rect 5615 1435 5635 1520
rect 5815 1435 5835 1520
rect 6015 1435 6035 1520
rect 6215 1435 6235 1520
rect -195 1405 -190 1435
rect -160 1405 -155 1435
rect -195 1365 -185 1405
rect -165 1395 -155 1405
rect 5 1405 10 1435
rect 40 1405 45 1435
rect 5 1395 45 1405
rect 205 1405 210 1435
rect 240 1405 245 1435
rect 205 1395 245 1405
rect 405 1405 410 1435
rect 440 1405 445 1435
rect 405 1395 445 1405
rect 605 1405 610 1435
rect 640 1405 645 1435
rect 605 1395 645 1405
rect 805 1405 810 1435
rect 840 1405 845 1435
rect 805 1395 845 1405
rect 1005 1405 1010 1435
rect 1040 1405 1045 1435
rect 1005 1395 1045 1405
rect 1205 1405 1210 1435
rect 1240 1405 1245 1435
rect 1205 1395 1245 1405
rect 1405 1405 1410 1435
rect 1440 1405 1445 1435
rect 1405 1395 1445 1405
rect 1605 1405 1610 1435
rect 1640 1405 1645 1435
rect 1605 1395 1645 1405
rect 1805 1405 1810 1435
rect 1840 1405 1845 1435
rect 1805 1395 1845 1405
rect 2005 1405 2010 1435
rect 2040 1405 2045 1435
rect 2005 1395 2045 1405
rect 2205 1405 2210 1435
rect 2240 1405 2245 1435
rect 2205 1395 2245 1405
rect 2405 1405 2410 1435
rect 2440 1405 2445 1435
rect 2405 1395 2445 1405
rect 2605 1405 2610 1435
rect 2640 1405 2645 1435
rect 2605 1395 2645 1405
rect 2805 1405 2810 1435
rect 2840 1405 2845 1435
rect 2805 1395 2845 1405
rect 3005 1405 3010 1435
rect 3040 1405 3045 1435
rect 3005 1395 3045 1405
rect 3205 1405 3210 1435
rect 3240 1405 3245 1435
rect 3205 1395 3245 1405
rect 3405 1405 3410 1435
rect 3440 1405 3445 1435
rect 3405 1395 3445 1405
rect 3605 1405 3610 1435
rect 3640 1405 3645 1435
rect 3605 1395 3645 1405
rect 3805 1405 3810 1435
rect 3840 1405 3845 1435
rect 3805 1395 3845 1405
rect 4005 1405 4010 1435
rect 4040 1405 4045 1435
rect 4005 1395 4045 1405
rect 4205 1405 4210 1435
rect 4240 1405 4245 1435
rect 4205 1395 4245 1405
rect 4405 1405 4410 1435
rect 4440 1405 4445 1435
rect 4405 1395 4445 1405
rect 4605 1405 4610 1435
rect 4640 1405 4645 1435
rect 4605 1395 4645 1405
rect 4805 1405 4810 1435
rect 4840 1405 4845 1435
rect 4805 1395 4845 1405
rect 5005 1405 5010 1435
rect 5040 1405 5045 1435
rect 5005 1395 5045 1405
rect 5205 1405 5210 1435
rect 5240 1405 5245 1435
rect 5205 1395 5245 1405
rect 5405 1405 5410 1435
rect 5440 1405 5445 1435
rect 5405 1395 5445 1405
rect 5605 1405 5610 1435
rect 5640 1405 5645 1435
rect 5605 1395 5645 1405
rect 5805 1405 5810 1435
rect 5840 1405 5845 1435
rect 5805 1395 5845 1405
rect 6005 1405 6010 1435
rect 6040 1405 6045 1435
rect 6005 1395 6045 1405
rect 6205 1405 6210 1435
rect 6240 1405 6245 1435
rect 6205 1395 6245 1405
rect 6405 1405 6410 1435
rect 6440 1405 6445 1435
rect 6405 1395 6445 1405
rect -165 1375 -30 1395
rect 5 1375 6570 1395
rect -165 1365 -155 1375
rect -195 1335 -190 1365
rect -160 1335 -155 1365
rect 5 1365 45 1375
rect 5 1335 10 1365
rect 40 1335 45 1365
rect 205 1365 245 1375
rect 205 1335 210 1365
rect 240 1335 245 1365
rect 405 1365 445 1375
rect 405 1335 410 1365
rect 440 1335 445 1365
rect 605 1365 645 1375
rect 605 1335 610 1365
rect 640 1335 645 1365
rect 805 1365 845 1375
rect 805 1335 810 1365
rect 840 1335 845 1365
rect 1005 1365 1045 1375
rect 1005 1335 1010 1365
rect 1040 1335 1045 1365
rect 1205 1365 1245 1375
rect 1205 1335 1210 1365
rect 1240 1335 1245 1365
rect 1405 1365 1445 1375
rect 1405 1335 1410 1365
rect 1440 1335 1445 1365
rect 1605 1365 1645 1375
rect 1605 1335 1610 1365
rect 1640 1335 1645 1365
rect 1805 1365 1845 1375
rect 1805 1335 1810 1365
rect 1840 1335 1845 1365
rect 2005 1365 2045 1375
rect 2005 1335 2010 1365
rect 2040 1335 2045 1365
rect 2205 1365 2245 1375
rect 2205 1335 2210 1365
rect 2240 1335 2245 1365
rect 2405 1365 2445 1375
rect 2405 1335 2410 1365
rect 2440 1335 2445 1365
rect 2605 1365 2645 1375
rect 2605 1335 2610 1365
rect 2640 1335 2645 1365
rect 2805 1365 2845 1375
rect 2805 1335 2810 1365
rect 2840 1335 2845 1365
rect 3005 1365 3045 1375
rect 3005 1335 3010 1365
rect 3040 1335 3045 1365
rect 3205 1365 3245 1375
rect 3205 1335 3210 1365
rect 3240 1335 3245 1365
rect 3405 1365 3445 1375
rect 3405 1335 3410 1365
rect 3440 1335 3445 1365
rect 3605 1365 3645 1375
rect 3605 1335 3610 1365
rect 3640 1335 3645 1365
rect 3805 1365 3845 1375
rect 3805 1335 3810 1365
rect 3840 1335 3845 1365
rect 4005 1365 4045 1375
rect 4005 1335 4010 1365
rect 4040 1335 4045 1365
rect 4205 1365 4245 1375
rect 4205 1335 4210 1365
rect 4240 1335 4245 1365
rect 4405 1365 4445 1375
rect 4405 1335 4410 1365
rect 4440 1335 4445 1365
rect 4605 1365 4645 1375
rect 4605 1335 4610 1365
rect 4640 1335 4645 1365
rect 4805 1365 4845 1375
rect 4805 1335 4810 1365
rect 4840 1335 4845 1365
rect 5005 1365 5045 1375
rect 5005 1335 5010 1365
rect 5040 1335 5045 1365
rect 5205 1365 5245 1375
rect 5205 1335 5210 1365
rect 5240 1335 5245 1365
rect 5405 1365 5445 1375
rect 5405 1335 5410 1365
rect 5440 1335 5445 1365
rect 5605 1365 5645 1375
rect 5605 1335 5610 1365
rect 5640 1335 5645 1365
rect 5805 1365 5845 1375
rect 5805 1335 5810 1365
rect 5840 1335 5845 1365
rect 6005 1365 6045 1375
rect 6005 1335 6010 1365
rect 6040 1335 6045 1365
rect 6205 1365 6245 1375
rect 6205 1335 6210 1365
rect 6240 1335 6245 1365
rect 6405 1365 6445 1375
rect 6405 1335 6410 1365
rect 6440 1335 6445 1365
rect -188 1250 -185 1335
rect -165 1250 -162 1335
rect 15 1250 35 1335
rect 215 1250 235 1335
rect 415 1250 435 1335
rect 615 1250 635 1335
rect 815 1250 835 1335
rect 1015 1250 1035 1335
rect 1215 1250 1235 1335
rect 1415 1250 1435 1335
rect 1615 1250 1635 1335
rect 1815 1250 1835 1335
rect 2015 1250 2035 1335
rect 2215 1250 2235 1335
rect 2415 1250 2435 1335
rect 2615 1250 2635 1335
rect 2815 1250 2835 1335
rect 3015 1250 3035 1335
rect 3215 1250 3235 1335
rect 3415 1250 3435 1335
rect 3615 1250 3635 1335
rect 3815 1250 3835 1335
rect 4015 1250 4035 1335
rect 4215 1250 4235 1335
rect 4415 1250 4435 1335
rect 4615 1250 4635 1335
rect 4815 1250 4835 1335
rect 5015 1250 5035 1335
rect 5215 1250 5235 1335
rect 5415 1250 5435 1335
rect 5615 1250 5635 1335
rect 5815 1250 5835 1335
rect 6015 1250 6035 1335
rect 6215 1250 6235 1335
rect -195 1220 -190 1250
rect -160 1220 -155 1250
rect -195 1180 -185 1220
rect -165 1210 -155 1220
rect 5 1220 10 1250
rect 40 1220 45 1250
rect 5 1210 45 1220
rect 205 1220 210 1250
rect 240 1220 245 1250
rect 205 1210 245 1220
rect 405 1220 410 1250
rect 440 1220 445 1250
rect 405 1210 445 1220
rect 605 1220 610 1250
rect 640 1220 645 1250
rect 605 1210 645 1220
rect 805 1220 810 1250
rect 840 1220 845 1250
rect 805 1210 845 1220
rect 1005 1220 1010 1250
rect 1040 1220 1045 1250
rect 1005 1210 1045 1220
rect 1205 1220 1210 1250
rect 1240 1220 1245 1250
rect 1205 1210 1245 1220
rect 1405 1220 1410 1250
rect 1440 1220 1445 1250
rect 1405 1210 1445 1220
rect 1605 1220 1610 1250
rect 1640 1220 1645 1250
rect 1605 1210 1645 1220
rect 1805 1220 1810 1250
rect 1840 1220 1845 1250
rect 1805 1210 1845 1220
rect 2005 1220 2010 1250
rect 2040 1220 2045 1250
rect 2005 1210 2045 1220
rect 2205 1220 2210 1250
rect 2240 1220 2245 1250
rect 2205 1210 2245 1220
rect 2405 1220 2410 1250
rect 2440 1220 2445 1250
rect 2405 1210 2445 1220
rect 2605 1220 2610 1250
rect 2640 1220 2645 1250
rect 2605 1210 2645 1220
rect 2805 1220 2810 1250
rect 2840 1220 2845 1250
rect 2805 1210 2845 1220
rect 3005 1220 3010 1250
rect 3040 1220 3045 1250
rect 3005 1210 3045 1220
rect 3205 1220 3210 1250
rect 3240 1220 3245 1250
rect 3205 1210 3245 1220
rect 3405 1220 3410 1250
rect 3440 1220 3445 1250
rect 3405 1210 3445 1220
rect 3605 1220 3610 1250
rect 3640 1220 3645 1250
rect 3605 1210 3645 1220
rect 3805 1220 3810 1250
rect 3840 1220 3845 1250
rect 3805 1210 3845 1220
rect 4005 1220 4010 1250
rect 4040 1220 4045 1250
rect 4005 1210 4045 1220
rect 4205 1220 4210 1250
rect 4240 1220 4245 1250
rect 4205 1210 4245 1220
rect 4405 1220 4410 1250
rect 4440 1220 4445 1250
rect 4405 1210 4445 1220
rect 4605 1220 4610 1250
rect 4640 1220 4645 1250
rect 4605 1210 4645 1220
rect 4805 1220 4810 1250
rect 4840 1220 4845 1250
rect 4805 1210 4845 1220
rect 5005 1220 5010 1250
rect 5040 1220 5045 1250
rect 5005 1210 5045 1220
rect 5205 1220 5210 1250
rect 5240 1220 5245 1250
rect 5205 1210 5245 1220
rect 5405 1220 5410 1250
rect 5440 1220 5445 1250
rect 5405 1210 5445 1220
rect 5605 1220 5610 1250
rect 5640 1220 5645 1250
rect 5605 1210 5645 1220
rect 5805 1220 5810 1250
rect 5840 1220 5845 1250
rect 5805 1210 5845 1220
rect 6005 1220 6010 1250
rect 6040 1220 6045 1250
rect 6005 1210 6045 1220
rect 6205 1220 6210 1250
rect 6240 1220 6245 1250
rect 6205 1210 6245 1220
rect 6405 1220 6410 1250
rect 6440 1220 6445 1250
rect 6405 1210 6445 1220
rect -165 1190 -30 1210
rect 5 1190 6570 1210
rect -165 1180 -155 1190
rect -195 1150 -190 1180
rect -160 1150 -155 1180
rect 5 1180 45 1190
rect 5 1150 10 1180
rect 40 1150 45 1180
rect 205 1180 245 1190
rect 205 1150 210 1180
rect 240 1150 245 1180
rect 405 1180 445 1190
rect 405 1150 410 1180
rect 440 1150 445 1180
rect 605 1180 645 1190
rect 605 1150 610 1180
rect 640 1150 645 1180
rect 805 1180 845 1190
rect 805 1150 810 1180
rect 840 1150 845 1180
rect 1005 1180 1045 1190
rect 1005 1150 1010 1180
rect 1040 1150 1045 1180
rect 1205 1180 1245 1190
rect 1205 1150 1210 1180
rect 1240 1150 1245 1180
rect 1405 1180 1445 1190
rect 1405 1150 1410 1180
rect 1440 1150 1445 1180
rect 1605 1180 1645 1190
rect 1605 1150 1610 1180
rect 1640 1150 1645 1180
rect 1805 1180 1845 1190
rect 1805 1150 1810 1180
rect 1840 1150 1845 1180
rect 2005 1180 2045 1190
rect 2005 1150 2010 1180
rect 2040 1150 2045 1180
rect 2205 1180 2245 1190
rect 2205 1150 2210 1180
rect 2240 1150 2245 1180
rect 2405 1180 2445 1190
rect 2405 1150 2410 1180
rect 2440 1150 2445 1180
rect 2605 1180 2645 1190
rect 2605 1150 2610 1180
rect 2640 1150 2645 1180
rect 2805 1180 2845 1190
rect 2805 1150 2810 1180
rect 2840 1150 2845 1180
rect 3005 1180 3045 1190
rect 3005 1150 3010 1180
rect 3040 1150 3045 1180
rect 3205 1180 3245 1190
rect 3205 1150 3210 1180
rect 3240 1150 3245 1180
rect 3405 1180 3445 1190
rect 3405 1150 3410 1180
rect 3440 1150 3445 1180
rect 3605 1180 3645 1190
rect 3605 1150 3610 1180
rect 3640 1150 3645 1180
rect 3805 1180 3845 1190
rect 3805 1150 3810 1180
rect 3840 1150 3845 1180
rect 4005 1180 4045 1190
rect 4005 1150 4010 1180
rect 4040 1150 4045 1180
rect 4205 1180 4245 1190
rect 4205 1150 4210 1180
rect 4240 1150 4245 1180
rect 4405 1180 4445 1190
rect 4405 1150 4410 1180
rect 4440 1150 4445 1180
rect 4605 1180 4645 1190
rect 4605 1150 4610 1180
rect 4640 1150 4645 1180
rect 4805 1180 4845 1190
rect 4805 1150 4810 1180
rect 4840 1150 4845 1180
rect 5005 1180 5045 1190
rect 5005 1150 5010 1180
rect 5040 1150 5045 1180
rect 5205 1180 5245 1190
rect 5205 1150 5210 1180
rect 5240 1150 5245 1180
rect 5405 1180 5445 1190
rect 5405 1150 5410 1180
rect 5440 1150 5445 1180
rect 5605 1180 5645 1190
rect 5605 1150 5610 1180
rect 5640 1150 5645 1180
rect 5805 1180 5845 1190
rect 5805 1150 5810 1180
rect 5840 1150 5845 1180
rect 6005 1180 6045 1190
rect 6005 1150 6010 1180
rect 6040 1150 6045 1180
rect 6205 1180 6245 1190
rect 6205 1150 6210 1180
rect 6240 1150 6245 1180
rect 6405 1180 6445 1190
rect 6405 1150 6410 1180
rect 6440 1150 6445 1180
rect -188 1065 -185 1150
rect -165 1065 -162 1150
rect 15 1065 35 1150
rect 215 1065 235 1150
rect 415 1065 435 1150
rect 615 1065 635 1150
rect 815 1065 835 1150
rect 1015 1065 1035 1150
rect 1215 1065 1235 1150
rect 1415 1065 1435 1150
rect 1615 1065 1635 1150
rect 1815 1065 1835 1150
rect 2015 1065 2035 1150
rect 2215 1065 2235 1150
rect 2415 1065 2435 1150
rect 2615 1065 2635 1150
rect 2815 1065 2835 1150
rect 3015 1065 3035 1150
rect 3215 1065 3235 1150
rect 3415 1065 3435 1150
rect 3615 1065 3635 1150
rect 3815 1065 3835 1150
rect 4015 1065 4035 1150
rect 4215 1065 4235 1150
rect 4415 1065 4435 1150
rect 4615 1065 4635 1150
rect 4815 1065 4835 1150
rect 5015 1065 5035 1150
rect 5215 1065 5235 1150
rect 5415 1065 5435 1150
rect 5615 1065 5635 1150
rect 5815 1065 5835 1150
rect 6015 1065 6035 1150
rect 6215 1065 6235 1150
rect -195 1035 -190 1065
rect -160 1035 -155 1065
rect -195 995 -185 1035
rect -165 1025 -155 1035
rect 5 1035 10 1065
rect 40 1035 45 1065
rect 5 1025 45 1035
rect 205 1035 210 1065
rect 240 1035 245 1065
rect 205 1025 245 1035
rect 405 1035 410 1065
rect 440 1035 445 1065
rect 405 1025 445 1035
rect 605 1035 610 1065
rect 640 1035 645 1065
rect 605 1025 645 1035
rect 805 1035 810 1065
rect 840 1035 845 1065
rect 805 1025 845 1035
rect 1005 1035 1010 1065
rect 1040 1035 1045 1065
rect 1005 1025 1045 1035
rect 1205 1035 1210 1065
rect 1240 1035 1245 1065
rect 1205 1025 1245 1035
rect 1405 1035 1410 1065
rect 1440 1035 1445 1065
rect 1405 1025 1445 1035
rect 1605 1035 1610 1065
rect 1640 1035 1645 1065
rect 1605 1025 1645 1035
rect 1805 1035 1810 1065
rect 1840 1035 1845 1065
rect 1805 1025 1845 1035
rect 2005 1035 2010 1065
rect 2040 1035 2045 1065
rect 2005 1025 2045 1035
rect 2205 1035 2210 1065
rect 2240 1035 2245 1065
rect 2205 1025 2245 1035
rect 2405 1035 2410 1065
rect 2440 1035 2445 1065
rect 2405 1025 2445 1035
rect 2605 1035 2610 1065
rect 2640 1035 2645 1065
rect 2605 1025 2645 1035
rect 2805 1035 2810 1065
rect 2840 1035 2845 1065
rect 2805 1025 2845 1035
rect 3005 1035 3010 1065
rect 3040 1035 3045 1065
rect 3005 1025 3045 1035
rect 3205 1035 3210 1065
rect 3240 1035 3245 1065
rect 3205 1025 3245 1035
rect 3405 1035 3410 1065
rect 3440 1035 3445 1065
rect 3405 1025 3445 1035
rect 3605 1035 3610 1065
rect 3640 1035 3645 1065
rect 3605 1025 3645 1035
rect 3805 1035 3810 1065
rect 3840 1035 3845 1065
rect 3805 1025 3845 1035
rect 4005 1035 4010 1065
rect 4040 1035 4045 1065
rect 4005 1025 4045 1035
rect 4205 1035 4210 1065
rect 4240 1035 4245 1065
rect 4205 1025 4245 1035
rect 4405 1035 4410 1065
rect 4440 1035 4445 1065
rect 4405 1025 4445 1035
rect 4605 1035 4610 1065
rect 4640 1035 4645 1065
rect 4605 1025 4645 1035
rect 4805 1035 4810 1065
rect 4840 1035 4845 1065
rect 4805 1025 4845 1035
rect 5005 1035 5010 1065
rect 5040 1035 5045 1065
rect 5005 1025 5045 1035
rect 5205 1035 5210 1065
rect 5240 1035 5245 1065
rect 5205 1025 5245 1035
rect 5405 1035 5410 1065
rect 5440 1035 5445 1065
rect 5405 1025 5445 1035
rect 5605 1035 5610 1065
rect 5640 1035 5645 1065
rect 5605 1025 5645 1035
rect 5805 1035 5810 1065
rect 5840 1035 5845 1065
rect 5805 1025 5845 1035
rect 6005 1035 6010 1065
rect 6040 1035 6045 1065
rect 6005 1025 6045 1035
rect 6205 1035 6210 1065
rect 6240 1035 6245 1065
rect 6205 1025 6245 1035
rect 6405 1035 6410 1065
rect 6440 1035 6445 1065
rect 6405 1025 6445 1035
rect -165 1005 -30 1025
rect 5 1005 6570 1025
rect -165 995 -155 1005
rect -195 965 -190 995
rect -160 965 -155 995
rect 5 995 45 1005
rect 5 965 10 995
rect 40 965 45 995
rect 205 995 245 1005
rect 205 965 210 995
rect 240 965 245 995
rect 405 995 445 1005
rect 405 965 410 995
rect 440 965 445 995
rect 605 995 645 1005
rect 605 965 610 995
rect 640 965 645 995
rect 805 995 845 1005
rect 805 965 810 995
rect 840 965 845 995
rect 1005 995 1045 1005
rect 1005 965 1010 995
rect 1040 965 1045 995
rect 1205 995 1245 1005
rect 1205 965 1210 995
rect 1240 965 1245 995
rect 1405 995 1445 1005
rect 1405 965 1410 995
rect 1440 965 1445 995
rect 1605 995 1645 1005
rect 1605 965 1610 995
rect 1640 965 1645 995
rect 1805 995 1845 1005
rect 1805 965 1810 995
rect 1840 965 1845 995
rect 2005 995 2045 1005
rect 2005 965 2010 995
rect 2040 965 2045 995
rect 2205 995 2245 1005
rect 2205 965 2210 995
rect 2240 965 2245 995
rect 2405 995 2445 1005
rect 2405 965 2410 995
rect 2440 965 2445 995
rect 2605 995 2645 1005
rect 2605 965 2610 995
rect 2640 965 2645 995
rect 2805 995 2845 1005
rect 2805 965 2810 995
rect 2840 965 2845 995
rect 3005 995 3045 1005
rect 3005 965 3010 995
rect 3040 965 3045 995
rect 3205 995 3245 1005
rect 3205 965 3210 995
rect 3240 965 3245 995
rect 3405 995 3445 1005
rect 3405 965 3410 995
rect 3440 965 3445 995
rect 3605 995 3645 1005
rect 3605 965 3610 995
rect 3640 965 3645 995
rect 3805 995 3845 1005
rect 3805 965 3810 995
rect 3840 965 3845 995
rect 4005 995 4045 1005
rect 4005 965 4010 995
rect 4040 965 4045 995
rect 4205 995 4245 1005
rect 4205 965 4210 995
rect 4240 965 4245 995
rect 4405 995 4445 1005
rect 4405 965 4410 995
rect 4440 965 4445 995
rect 4605 995 4645 1005
rect 4605 965 4610 995
rect 4640 965 4645 995
rect 4805 995 4845 1005
rect 4805 965 4810 995
rect 4840 965 4845 995
rect 5005 995 5045 1005
rect 5005 965 5010 995
rect 5040 965 5045 995
rect 5205 995 5245 1005
rect 5205 965 5210 995
rect 5240 965 5245 995
rect 5405 995 5445 1005
rect 5405 965 5410 995
rect 5440 965 5445 995
rect 5605 995 5645 1005
rect 5605 965 5610 995
rect 5640 965 5645 995
rect 5805 995 5845 1005
rect 5805 965 5810 995
rect 5840 965 5845 995
rect 6005 995 6045 1005
rect 6005 965 6010 995
rect 6040 965 6045 995
rect 6205 995 6245 1005
rect 6205 965 6210 995
rect 6240 965 6245 995
rect 6405 995 6445 1005
rect 6405 965 6410 995
rect 6440 965 6445 995
rect -188 880 -185 965
rect -165 880 -162 965
rect 15 880 35 965
rect 215 880 235 965
rect 415 880 435 965
rect 615 880 635 965
rect 815 880 835 965
rect 1015 880 1035 965
rect 1215 880 1235 965
rect 1415 880 1435 965
rect 1615 880 1635 965
rect 1815 880 1835 965
rect 2015 880 2035 965
rect 2215 880 2235 965
rect 2415 880 2435 965
rect 2615 880 2635 965
rect 2815 880 2835 965
rect 3015 880 3035 965
rect 3215 880 3235 965
rect 3415 880 3435 965
rect 3615 880 3635 965
rect 3815 880 3835 965
rect 4015 880 4035 965
rect 4215 880 4235 965
rect 4415 880 4435 965
rect 4615 880 4635 965
rect 4815 880 4835 965
rect 5015 880 5035 965
rect 5215 880 5235 965
rect 5415 880 5435 965
rect 5615 880 5635 965
rect 5815 880 5835 965
rect 6015 880 6035 965
rect 6215 880 6235 965
rect -195 850 -190 880
rect -160 850 -155 880
rect -195 810 -185 850
rect -165 840 -155 850
rect 5 850 10 880
rect 40 850 45 880
rect 5 840 45 850
rect 205 850 210 880
rect 240 850 245 880
rect 205 840 245 850
rect 405 850 410 880
rect 440 850 445 880
rect 405 840 445 850
rect 605 850 610 880
rect 640 850 645 880
rect 605 840 645 850
rect 805 850 810 880
rect 840 850 845 880
rect 805 840 845 850
rect 1005 850 1010 880
rect 1040 850 1045 880
rect 1005 840 1045 850
rect 1205 850 1210 880
rect 1240 850 1245 880
rect 1205 840 1245 850
rect 1405 850 1410 880
rect 1440 850 1445 880
rect 1405 840 1445 850
rect 1605 850 1610 880
rect 1640 850 1645 880
rect 1605 840 1645 850
rect 1805 850 1810 880
rect 1840 850 1845 880
rect 1805 840 1845 850
rect 2005 850 2010 880
rect 2040 850 2045 880
rect 2005 840 2045 850
rect 2205 850 2210 880
rect 2240 850 2245 880
rect 2205 840 2245 850
rect 2405 850 2410 880
rect 2440 850 2445 880
rect 2405 840 2445 850
rect 2605 850 2610 880
rect 2640 850 2645 880
rect 2605 840 2645 850
rect 2805 850 2810 880
rect 2840 850 2845 880
rect 2805 840 2845 850
rect 3005 850 3010 880
rect 3040 850 3045 880
rect 3005 840 3045 850
rect 3205 850 3210 880
rect 3240 850 3245 880
rect 3205 840 3245 850
rect 3405 850 3410 880
rect 3440 850 3445 880
rect 3405 840 3445 850
rect 3605 850 3610 880
rect 3640 850 3645 880
rect 3605 840 3645 850
rect 3805 850 3810 880
rect 3840 850 3845 880
rect 3805 840 3845 850
rect 4005 850 4010 880
rect 4040 850 4045 880
rect 4005 840 4045 850
rect 4205 850 4210 880
rect 4240 850 4245 880
rect 4205 840 4245 850
rect 4405 850 4410 880
rect 4440 850 4445 880
rect 4405 840 4445 850
rect 4605 850 4610 880
rect 4640 850 4645 880
rect 4605 840 4645 850
rect 4805 850 4810 880
rect 4840 850 4845 880
rect 4805 840 4845 850
rect 5005 850 5010 880
rect 5040 850 5045 880
rect 5005 840 5045 850
rect 5205 850 5210 880
rect 5240 850 5245 880
rect 5205 840 5245 850
rect 5405 850 5410 880
rect 5440 850 5445 880
rect 5405 840 5445 850
rect 5605 850 5610 880
rect 5640 850 5645 880
rect 5605 840 5645 850
rect 5805 850 5810 880
rect 5840 850 5845 880
rect 5805 840 5845 850
rect 6005 850 6010 880
rect 6040 850 6045 880
rect 6005 840 6045 850
rect 6205 850 6210 880
rect 6240 850 6245 880
rect 6205 840 6245 850
rect 6405 850 6410 880
rect 6440 850 6445 880
rect 6405 840 6445 850
rect -165 820 -30 840
rect 5 820 6570 840
rect -165 810 -155 820
rect -195 780 -190 810
rect -160 780 -155 810
rect 5 810 45 820
rect 5 780 10 810
rect 40 780 45 810
rect 205 810 245 820
rect 205 780 210 810
rect 240 780 245 810
rect 405 810 445 820
rect 405 780 410 810
rect 440 780 445 810
rect 605 810 645 820
rect 605 780 610 810
rect 640 780 645 810
rect 805 810 845 820
rect 805 780 810 810
rect 840 780 845 810
rect 1005 810 1045 820
rect 1005 780 1010 810
rect 1040 780 1045 810
rect 1205 810 1245 820
rect 1205 780 1210 810
rect 1240 780 1245 810
rect 1405 810 1445 820
rect 1405 780 1410 810
rect 1440 780 1445 810
rect 1605 810 1645 820
rect 1605 780 1610 810
rect 1640 780 1645 810
rect 1805 810 1845 820
rect 1805 780 1810 810
rect 1840 780 1845 810
rect 2005 810 2045 820
rect 2005 780 2010 810
rect 2040 780 2045 810
rect 2205 810 2245 820
rect 2205 780 2210 810
rect 2240 780 2245 810
rect 2405 810 2445 820
rect 2405 780 2410 810
rect 2440 780 2445 810
rect 2605 810 2645 820
rect 2605 780 2610 810
rect 2640 780 2645 810
rect 2805 810 2845 820
rect 2805 780 2810 810
rect 2840 780 2845 810
rect 3005 810 3045 820
rect 3005 780 3010 810
rect 3040 780 3045 810
rect 3205 810 3245 820
rect 3205 780 3210 810
rect 3240 780 3245 810
rect 3405 810 3445 820
rect 3405 780 3410 810
rect 3440 780 3445 810
rect 3605 810 3645 820
rect 3605 780 3610 810
rect 3640 780 3645 810
rect 3805 810 3845 820
rect 3805 780 3810 810
rect 3840 780 3845 810
rect 4005 810 4045 820
rect 4005 780 4010 810
rect 4040 780 4045 810
rect 4205 810 4245 820
rect 4205 780 4210 810
rect 4240 780 4245 810
rect 4405 810 4445 820
rect 4405 780 4410 810
rect 4440 780 4445 810
rect 4605 810 4645 820
rect 4605 780 4610 810
rect 4640 780 4645 810
rect 4805 810 4845 820
rect 4805 780 4810 810
rect 4840 780 4845 810
rect 5005 810 5045 820
rect 5005 780 5010 810
rect 5040 780 5045 810
rect 5205 810 5245 820
rect 5205 780 5210 810
rect 5240 780 5245 810
rect 5405 810 5445 820
rect 5405 780 5410 810
rect 5440 780 5445 810
rect 5605 810 5645 820
rect 5605 780 5610 810
rect 5640 780 5645 810
rect 5805 810 5845 820
rect 5805 780 5810 810
rect 5840 780 5845 810
rect 6005 810 6045 820
rect 6005 780 6010 810
rect 6040 780 6045 810
rect 6205 810 6245 820
rect 6205 780 6210 810
rect 6240 780 6245 810
rect 6405 810 6445 820
rect 6405 780 6410 810
rect 6440 780 6445 810
rect -188 695 -185 780
rect -165 695 -162 780
rect 15 695 35 780
rect 215 695 235 780
rect 415 695 435 780
rect 615 695 635 780
rect 815 695 835 780
rect 1015 695 1035 780
rect 1215 695 1235 780
rect 1415 695 1435 780
rect 1615 695 1635 780
rect 1815 695 1835 780
rect 2015 695 2035 780
rect 2215 695 2235 780
rect 2415 695 2435 780
rect 2615 695 2635 780
rect 2815 695 2835 780
rect 3015 695 3035 780
rect 3215 695 3235 780
rect 3415 695 3435 780
rect 3615 695 3635 780
rect 3815 695 3835 780
rect 4015 695 4035 780
rect 4215 695 4235 780
rect 4415 695 4435 780
rect 4615 695 4635 780
rect 4815 695 4835 780
rect 5015 695 5035 780
rect 5215 695 5235 780
rect 5415 695 5435 780
rect 5615 695 5635 780
rect 5815 695 5835 780
rect 6015 695 6035 780
rect 6215 695 6235 780
rect -195 665 -190 695
rect -160 665 -155 695
rect -195 625 -185 665
rect -165 655 -155 665
rect 5 665 10 695
rect 40 665 45 695
rect 5 655 45 665
rect 205 665 210 695
rect 240 665 245 695
rect 205 655 245 665
rect 405 665 410 695
rect 440 665 445 695
rect 405 655 445 665
rect 605 665 610 695
rect 640 665 645 695
rect 605 655 645 665
rect 805 665 810 695
rect 840 665 845 695
rect 805 655 845 665
rect 1005 665 1010 695
rect 1040 665 1045 695
rect 1005 655 1045 665
rect 1205 665 1210 695
rect 1240 665 1245 695
rect 1205 655 1245 665
rect 1405 665 1410 695
rect 1440 665 1445 695
rect 1405 655 1445 665
rect 1605 665 1610 695
rect 1640 665 1645 695
rect 1605 655 1645 665
rect 1805 665 1810 695
rect 1840 665 1845 695
rect 1805 655 1845 665
rect 2005 665 2010 695
rect 2040 665 2045 695
rect 2005 655 2045 665
rect 2205 665 2210 695
rect 2240 665 2245 695
rect 2205 655 2245 665
rect 2405 665 2410 695
rect 2440 665 2445 695
rect 2405 655 2445 665
rect 2605 665 2610 695
rect 2640 665 2645 695
rect 2605 655 2645 665
rect 2805 665 2810 695
rect 2840 665 2845 695
rect 2805 655 2845 665
rect 3005 665 3010 695
rect 3040 665 3045 695
rect 3005 655 3045 665
rect 3205 665 3210 695
rect 3240 665 3245 695
rect 3205 655 3245 665
rect 3405 665 3410 695
rect 3440 665 3445 695
rect 3405 655 3445 665
rect 3605 665 3610 695
rect 3640 665 3645 695
rect 3605 655 3645 665
rect 3805 665 3810 695
rect 3840 665 3845 695
rect 3805 655 3845 665
rect 4005 665 4010 695
rect 4040 665 4045 695
rect 4005 655 4045 665
rect 4205 665 4210 695
rect 4240 665 4245 695
rect 4205 655 4245 665
rect 4405 665 4410 695
rect 4440 665 4445 695
rect 4405 655 4445 665
rect 4605 665 4610 695
rect 4640 665 4645 695
rect 4605 655 4645 665
rect 4805 665 4810 695
rect 4840 665 4845 695
rect 4805 655 4845 665
rect 5005 665 5010 695
rect 5040 665 5045 695
rect 5005 655 5045 665
rect 5205 665 5210 695
rect 5240 665 5245 695
rect 5205 655 5245 665
rect 5405 665 5410 695
rect 5440 665 5445 695
rect 5405 655 5445 665
rect 5605 665 5610 695
rect 5640 665 5645 695
rect 5605 655 5645 665
rect 5805 665 5810 695
rect 5840 665 5845 695
rect 5805 655 5845 665
rect 6005 665 6010 695
rect 6040 665 6045 695
rect 6005 655 6045 665
rect 6205 665 6210 695
rect 6240 665 6245 695
rect 6205 655 6245 665
rect 6405 665 6410 695
rect 6440 665 6445 695
rect 6405 655 6445 665
rect -165 635 -30 655
rect 5 635 6570 655
rect -165 625 -155 635
rect -195 595 -190 625
rect -160 595 -155 625
rect 5 625 45 635
rect 5 595 10 625
rect 40 595 45 625
rect 205 625 245 635
rect 205 595 210 625
rect 240 595 245 625
rect 405 625 445 635
rect 405 595 410 625
rect 440 595 445 625
rect 605 625 645 635
rect 605 595 610 625
rect 640 595 645 625
rect 805 625 845 635
rect 805 595 810 625
rect 840 595 845 625
rect 1005 625 1045 635
rect 1005 595 1010 625
rect 1040 595 1045 625
rect 1205 625 1245 635
rect 1205 595 1210 625
rect 1240 595 1245 625
rect 1405 625 1445 635
rect 1405 595 1410 625
rect 1440 595 1445 625
rect 1605 625 1645 635
rect 1605 595 1610 625
rect 1640 595 1645 625
rect 1805 625 1845 635
rect 1805 595 1810 625
rect 1840 595 1845 625
rect 2005 625 2045 635
rect 2005 595 2010 625
rect 2040 595 2045 625
rect 2205 625 2245 635
rect 2205 595 2210 625
rect 2240 595 2245 625
rect 2405 625 2445 635
rect 2405 595 2410 625
rect 2440 595 2445 625
rect 2605 625 2645 635
rect 2605 595 2610 625
rect 2640 595 2645 625
rect 2805 625 2845 635
rect 2805 595 2810 625
rect 2840 595 2845 625
rect 3005 625 3045 635
rect 3005 595 3010 625
rect 3040 595 3045 625
rect 3205 625 3245 635
rect 3205 595 3210 625
rect 3240 595 3245 625
rect 3405 625 3445 635
rect 3405 595 3410 625
rect 3440 595 3445 625
rect 3605 625 3645 635
rect 3605 595 3610 625
rect 3640 595 3645 625
rect 3805 625 3845 635
rect 3805 595 3810 625
rect 3840 595 3845 625
rect 4005 625 4045 635
rect 4005 595 4010 625
rect 4040 595 4045 625
rect 4205 625 4245 635
rect 4205 595 4210 625
rect 4240 595 4245 625
rect 4405 625 4445 635
rect 4405 595 4410 625
rect 4440 595 4445 625
rect 4605 625 4645 635
rect 4605 595 4610 625
rect 4640 595 4645 625
rect 4805 625 4845 635
rect 4805 595 4810 625
rect 4840 595 4845 625
rect 5005 625 5045 635
rect 5005 595 5010 625
rect 5040 595 5045 625
rect 5205 625 5245 635
rect 5205 595 5210 625
rect 5240 595 5245 625
rect 5405 625 5445 635
rect 5405 595 5410 625
rect 5440 595 5445 625
rect 5605 625 5645 635
rect 5605 595 5610 625
rect 5640 595 5645 625
rect 5805 625 5845 635
rect 5805 595 5810 625
rect 5840 595 5845 625
rect 6005 625 6045 635
rect 6005 595 6010 625
rect 6040 595 6045 625
rect 6205 625 6245 635
rect 6205 595 6210 625
rect 6240 595 6245 625
rect 6405 625 6445 635
rect 6405 595 6410 625
rect 6440 595 6445 625
rect -188 510 -185 595
rect -165 510 -162 595
rect 15 510 35 595
rect 215 510 235 595
rect 415 510 435 595
rect 615 510 635 595
rect 815 510 835 595
rect 1015 510 1035 595
rect 1215 510 1235 595
rect 1415 510 1435 595
rect 1615 510 1635 595
rect 1815 510 1835 595
rect 2015 510 2035 595
rect 2215 510 2235 595
rect 2415 510 2435 595
rect 2615 510 2635 595
rect 2815 510 2835 595
rect 3015 510 3035 595
rect 3215 510 3235 595
rect 3415 510 3435 595
rect 3615 510 3635 595
rect 3815 510 3835 595
rect 4015 510 4035 595
rect 4215 510 4235 595
rect 4415 510 4435 595
rect 4615 510 4635 595
rect 4815 510 4835 595
rect 5015 510 5035 595
rect 5215 510 5235 595
rect 5415 510 5435 595
rect 5615 510 5635 595
rect 5815 510 5835 595
rect 6015 510 6035 595
rect 6215 510 6235 595
rect -195 480 -190 510
rect -160 480 -155 510
rect -195 440 -185 480
rect -165 470 -155 480
rect 5 480 10 510
rect 40 480 45 510
rect 5 470 45 480
rect 205 480 210 510
rect 240 480 245 510
rect 205 470 245 480
rect 405 480 410 510
rect 440 480 445 510
rect 405 470 445 480
rect 605 480 610 510
rect 640 480 645 510
rect 605 470 645 480
rect 805 480 810 510
rect 840 480 845 510
rect 805 470 845 480
rect 1005 480 1010 510
rect 1040 480 1045 510
rect 1005 470 1045 480
rect 1205 480 1210 510
rect 1240 480 1245 510
rect 1205 470 1245 480
rect 1405 480 1410 510
rect 1440 480 1445 510
rect 1405 470 1445 480
rect 1605 480 1610 510
rect 1640 480 1645 510
rect 1605 470 1645 480
rect 1805 480 1810 510
rect 1840 480 1845 510
rect 1805 470 1845 480
rect 2005 480 2010 510
rect 2040 480 2045 510
rect 2005 470 2045 480
rect 2205 480 2210 510
rect 2240 480 2245 510
rect 2205 470 2245 480
rect 2405 480 2410 510
rect 2440 480 2445 510
rect 2405 470 2445 480
rect 2605 480 2610 510
rect 2640 480 2645 510
rect 2605 470 2645 480
rect 2805 480 2810 510
rect 2840 480 2845 510
rect 2805 470 2845 480
rect 3005 480 3010 510
rect 3040 480 3045 510
rect 3005 470 3045 480
rect 3205 480 3210 510
rect 3240 480 3245 510
rect 3205 470 3245 480
rect 3405 480 3410 510
rect 3440 480 3445 510
rect 3405 470 3445 480
rect 3605 480 3610 510
rect 3640 480 3645 510
rect 3605 470 3645 480
rect 3805 480 3810 510
rect 3840 480 3845 510
rect 3805 470 3845 480
rect 4005 480 4010 510
rect 4040 480 4045 510
rect 4005 470 4045 480
rect 4205 480 4210 510
rect 4240 480 4245 510
rect 4205 470 4245 480
rect 4405 480 4410 510
rect 4440 480 4445 510
rect 4405 470 4445 480
rect 4605 480 4610 510
rect 4640 480 4645 510
rect 4605 470 4645 480
rect 4805 480 4810 510
rect 4840 480 4845 510
rect 4805 470 4845 480
rect 5005 480 5010 510
rect 5040 480 5045 510
rect 5005 470 5045 480
rect 5205 480 5210 510
rect 5240 480 5245 510
rect 5205 470 5245 480
rect 5405 480 5410 510
rect 5440 480 5445 510
rect 5405 470 5445 480
rect 5605 480 5610 510
rect 5640 480 5645 510
rect 5605 470 5645 480
rect 5805 480 5810 510
rect 5840 480 5845 510
rect 5805 470 5845 480
rect 6005 480 6010 510
rect 6040 480 6045 510
rect 6005 470 6045 480
rect 6205 480 6210 510
rect 6240 480 6245 510
rect 6205 470 6245 480
rect 6405 480 6410 510
rect 6440 480 6445 510
rect 6405 470 6445 480
rect -165 450 -30 470
rect 5 450 6570 470
rect -165 440 -155 450
rect -195 410 -190 440
rect -160 410 -155 440
rect 5 440 45 450
rect 5 410 10 440
rect 40 410 45 440
rect 205 440 245 450
rect 205 410 210 440
rect 240 410 245 440
rect 405 440 445 450
rect 405 410 410 440
rect 440 410 445 440
rect 605 440 645 450
rect 605 410 610 440
rect 640 410 645 440
rect 805 440 845 450
rect 805 410 810 440
rect 840 410 845 440
rect 1005 440 1045 450
rect 1005 410 1010 440
rect 1040 410 1045 440
rect 1205 440 1245 450
rect 1205 410 1210 440
rect 1240 410 1245 440
rect 1405 440 1445 450
rect 1405 410 1410 440
rect 1440 410 1445 440
rect 1605 440 1645 450
rect 1605 410 1610 440
rect 1640 410 1645 440
rect 1805 440 1845 450
rect 1805 410 1810 440
rect 1840 410 1845 440
rect 2005 440 2045 450
rect 2005 410 2010 440
rect 2040 410 2045 440
rect 2205 440 2245 450
rect 2205 410 2210 440
rect 2240 410 2245 440
rect 2405 440 2445 450
rect 2405 410 2410 440
rect 2440 410 2445 440
rect 2605 440 2645 450
rect 2605 410 2610 440
rect 2640 410 2645 440
rect 2805 440 2845 450
rect 2805 410 2810 440
rect 2840 410 2845 440
rect 3005 440 3045 450
rect 3005 410 3010 440
rect 3040 410 3045 440
rect 3205 440 3245 450
rect 3205 410 3210 440
rect 3240 410 3245 440
rect 3405 440 3445 450
rect 3405 410 3410 440
rect 3440 410 3445 440
rect 3605 440 3645 450
rect 3605 410 3610 440
rect 3640 410 3645 440
rect 3805 440 3845 450
rect 3805 410 3810 440
rect 3840 410 3845 440
rect 4005 440 4045 450
rect 4005 410 4010 440
rect 4040 410 4045 440
rect 4205 440 4245 450
rect 4205 410 4210 440
rect 4240 410 4245 440
rect 4405 440 4445 450
rect 4405 410 4410 440
rect 4440 410 4445 440
rect 4605 440 4645 450
rect 4605 410 4610 440
rect 4640 410 4645 440
rect 4805 440 4845 450
rect 4805 410 4810 440
rect 4840 410 4845 440
rect 5005 440 5045 450
rect 5005 410 5010 440
rect 5040 410 5045 440
rect 5205 440 5245 450
rect 5205 410 5210 440
rect 5240 410 5245 440
rect 5405 440 5445 450
rect 5405 410 5410 440
rect 5440 410 5445 440
rect 5605 440 5645 450
rect 5605 410 5610 440
rect 5640 410 5645 440
rect 5805 440 5845 450
rect 5805 410 5810 440
rect 5840 410 5845 440
rect 6005 440 6045 450
rect 6005 410 6010 440
rect 6040 410 6045 440
rect 6205 440 6245 450
rect 6205 410 6210 440
rect 6240 410 6245 440
rect 6405 440 6445 450
rect 6405 410 6410 440
rect 6440 410 6445 440
rect -188 325 -185 410
rect -165 325 -162 410
rect 15 325 35 410
rect 215 325 235 410
rect 415 325 435 410
rect 615 325 635 410
rect 815 325 835 410
rect 1015 325 1035 410
rect 1215 325 1235 410
rect 1415 325 1435 410
rect 1615 325 1635 410
rect 1815 325 1835 410
rect 2015 325 2035 410
rect 2215 325 2235 410
rect 2415 325 2435 410
rect 2615 325 2635 410
rect 2815 325 2835 410
rect 3015 325 3035 410
rect 3215 325 3235 410
rect 3415 325 3435 410
rect 3615 325 3635 410
rect 3815 325 3835 410
rect 4015 325 4035 410
rect 4215 325 4235 410
rect 4415 325 4435 410
rect 4615 325 4635 410
rect 4815 325 4835 410
rect 5015 325 5035 410
rect 5215 325 5235 410
rect 5415 325 5435 410
rect 5615 325 5635 410
rect 5815 325 5835 410
rect 6015 325 6035 410
rect 6215 325 6235 410
rect -195 295 -190 325
rect -160 295 -155 325
rect -195 255 -185 295
rect -165 285 -155 295
rect 5 295 10 325
rect 40 295 45 325
rect 5 285 45 295
rect 205 295 210 325
rect 240 295 245 325
rect 205 285 245 295
rect 405 295 410 325
rect 440 295 445 325
rect 405 285 445 295
rect 605 295 610 325
rect 640 295 645 325
rect 605 285 645 295
rect 805 295 810 325
rect 840 295 845 325
rect 805 285 845 295
rect 1005 295 1010 325
rect 1040 295 1045 325
rect 1005 285 1045 295
rect 1205 295 1210 325
rect 1240 295 1245 325
rect 1205 285 1245 295
rect 1405 295 1410 325
rect 1440 295 1445 325
rect 1405 285 1445 295
rect 1605 295 1610 325
rect 1640 295 1645 325
rect 1605 285 1645 295
rect 1805 295 1810 325
rect 1840 295 1845 325
rect 1805 285 1845 295
rect 2005 295 2010 325
rect 2040 295 2045 325
rect 2005 285 2045 295
rect 2205 295 2210 325
rect 2240 295 2245 325
rect 2205 285 2245 295
rect 2405 295 2410 325
rect 2440 295 2445 325
rect 2405 285 2445 295
rect 2605 295 2610 325
rect 2640 295 2645 325
rect 2605 285 2645 295
rect 2805 295 2810 325
rect 2840 295 2845 325
rect 2805 285 2845 295
rect 3005 295 3010 325
rect 3040 295 3045 325
rect 3005 285 3045 295
rect 3205 295 3210 325
rect 3240 295 3245 325
rect 3205 285 3245 295
rect 3405 295 3410 325
rect 3440 295 3445 325
rect 3405 285 3445 295
rect 3605 295 3610 325
rect 3640 295 3645 325
rect 3605 285 3645 295
rect 3805 295 3810 325
rect 3840 295 3845 325
rect 3805 285 3845 295
rect 4005 295 4010 325
rect 4040 295 4045 325
rect 4005 285 4045 295
rect 4205 295 4210 325
rect 4240 295 4245 325
rect 4205 285 4245 295
rect 4405 295 4410 325
rect 4440 295 4445 325
rect 4405 285 4445 295
rect 4605 295 4610 325
rect 4640 295 4645 325
rect 4605 285 4645 295
rect 4805 295 4810 325
rect 4840 295 4845 325
rect 4805 285 4845 295
rect 5005 295 5010 325
rect 5040 295 5045 325
rect 5005 285 5045 295
rect 5205 295 5210 325
rect 5240 295 5245 325
rect 5205 285 5245 295
rect 5405 295 5410 325
rect 5440 295 5445 325
rect 5405 285 5445 295
rect 5605 295 5610 325
rect 5640 295 5645 325
rect 5605 285 5645 295
rect 5805 295 5810 325
rect 5840 295 5845 325
rect 5805 285 5845 295
rect 6005 295 6010 325
rect 6040 295 6045 325
rect 6005 285 6045 295
rect 6205 295 6210 325
rect 6240 295 6245 325
rect 6205 285 6245 295
rect 6405 295 6410 325
rect 6440 295 6445 325
rect 6405 285 6445 295
rect -165 265 -30 285
rect 5 265 6570 285
rect -165 255 -155 265
rect -195 225 -190 255
rect -160 225 -155 255
rect 5 255 45 265
rect 5 225 10 255
rect 40 225 45 255
rect 205 255 245 265
rect 205 225 210 255
rect 240 225 245 255
rect 405 255 445 265
rect 405 225 410 255
rect 440 225 445 255
rect 605 255 645 265
rect 605 225 610 255
rect 640 225 645 255
rect 805 255 845 265
rect 805 225 810 255
rect 840 225 845 255
rect 1005 255 1045 265
rect 1005 225 1010 255
rect 1040 225 1045 255
rect 1205 255 1245 265
rect 1205 225 1210 255
rect 1240 225 1245 255
rect 1405 255 1445 265
rect 1405 225 1410 255
rect 1440 225 1445 255
rect 1605 255 1645 265
rect 1605 225 1610 255
rect 1640 225 1645 255
rect 1805 255 1845 265
rect 1805 225 1810 255
rect 1840 225 1845 255
rect 2005 255 2045 265
rect 2005 225 2010 255
rect 2040 225 2045 255
rect 2205 255 2245 265
rect 2205 225 2210 255
rect 2240 225 2245 255
rect 2405 255 2445 265
rect 2405 225 2410 255
rect 2440 225 2445 255
rect 2605 255 2645 265
rect 2605 225 2610 255
rect 2640 225 2645 255
rect 2805 255 2845 265
rect 2805 225 2810 255
rect 2840 225 2845 255
rect 3005 255 3045 265
rect 3005 225 3010 255
rect 3040 225 3045 255
rect 3205 255 3245 265
rect 3205 225 3210 255
rect 3240 225 3245 255
rect 3405 255 3445 265
rect 3405 225 3410 255
rect 3440 225 3445 255
rect 3605 255 3645 265
rect 3605 225 3610 255
rect 3640 225 3645 255
rect 3805 255 3845 265
rect 3805 225 3810 255
rect 3840 225 3845 255
rect 4005 255 4045 265
rect 4005 225 4010 255
rect 4040 225 4045 255
rect 4205 255 4245 265
rect 4205 225 4210 255
rect 4240 225 4245 255
rect 4405 255 4445 265
rect 4405 225 4410 255
rect 4440 225 4445 255
rect 4605 255 4645 265
rect 4605 225 4610 255
rect 4640 225 4645 255
rect 4805 255 4845 265
rect 4805 225 4810 255
rect 4840 225 4845 255
rect 5005 255 5045 265
rect 5005 225 5010 255
rect 5040 225 5045 255
rect 5205 255 5245 265
rect 5205 225 5210 255
rect 5240 225 5245 255
rect 5405 255 5445 265
rect 5405 225 5410 255
rect 5440 225 5445 255
rect 5605 255 5645 265
rect 5605 225 5610 255
rect 5640 225 5645 255
rect 5805 255 5845 265
rect 5805 225 5810 255
rect 5840 225 5845 255
rect 6005 255 6045 265
rect 6005 225 6010 255
rect 6040 225 6045 255
rect 6205 255 6245 265
rect 6205 225 6210 255
rect 6240 225 6245 255
rect 6405 255 6445 265
rect 6405 225 6410 255
rect 6440 225 6445 255
rect -188 140 -185 225
rect -165 140 -162 225
rect 15 140 35 225
rect 215 140 235 225
rect 415 140 435 225
rect 615 140 635 225
rect 815 140 835 225
rect 1015 140 1035 225
rect 1215 140 1235 225
rect 1415 140 1435 225
rect 1615 140 1635 225
rect 1815 140 1835 225
rect 2015 140 2035 225
rect 2215 140 2235 225
rect 2415 140 2435 225
rect 2615 140 2635 225
rect 2815 140 2835 225
rect 3015 140 3035 225
rect 3215 140 3235 225
rect 3415 140 3435 225
rect 3615 140 3635 225
rect 3815 140 3835 225
rect 4015 140 4035 225
rect 4215 140 4235 225
rect 4415 140 4435 225
rect 4615 140 4635 225
rect 4815 140 4835 225
rect 5015 140 5035 225
rect 5215 140 5235 225
rect 5415 140 5435 225
rect 5615 140 5635 225
rect 5815 140 5835 225
rect 6015 140 6035 225
rect 6215 140 6235 225
rect -195 110 -190 140
rect -160 110 -155 140
rect -195 70 -185 110
rect -165 100 -155 110
rect 5 110 10 140
rect 40 110 45 140
rect 5 100 45 110
rect 205 110 210 140
rect 240 110 245 140
rect 205 100 245 110
rect 405 110 410 140
rect 440 110 445 140
rect 405 100 445 110
rect 605 110 610 140
rect 640 110 645 140
rect 605 100 645 110
rect 805 110 810 140
rect 840 110 845 140
rect 805 100 845 110
rect 1005 110 1010 140
rect 1040 110 1045 140
rect 1005 100 1045 110
rect 1205 110 1210 140
rect 1240 110 1245 140
rect 1205 100 1245 110
rect 1405 110 1410 140
rect 1440 110 1445 140
rect 1405 100 1445 110
rect 1605 110 1610 140
rect 1640 110 1645 140
rect 1605 100 1645 110
rect 1805 110 1810 140
rect 1840 110 1845 140
rect 1805 100 1845 110
rect 2005 110 2010 140
rect 2040 110 2045 140
rect 2005 100 2045 110
rect 2205 110 2210 140
rect 2240 110 2245 140
rect 2205 100 2245 110
rect 2405 110 2410 140
rect 2440 110 2445 140
rect 2405 100 2445 110
rect 2605 110 2610 140
rect 2640 110 2645 140
rect 2605 100 2645 110
rect 2805 110 2810 140
rect 2840 110 2845 140
rect 2805 100 2845 110
rect 3005 110 3010 140
rect 3040 110 3045 140
rect 3005 100 3045 110
rect 3205 110 3210 140
rect 3240 110 3245 140
rect 3205 100 3245 110
rect 3405 110 3410 140
rect 3440 110 3445 140
rect 3405 100 3445 110
rect 3605 110 3610 140
rect 3640 110 3645 140
rect 3605 100 3645 110
rect 3805 110 3810 140
rect 3840 110 3845 140
rect 3805 100 3845 110
rect 4005 110 4010 140
rect 4040 110 4045 140
rect 4005 100 4045 110
rect 4205 110 4210 140
rect 4240 110 4245 140
rect 4205 100 4245 110
rect 4405 110 4410 140
rect 4440 110 4445 140
rect 4405 100 4445 110
rect 4605 110 4610 140
rect 4640 110 4645 140
rect 4605 100 4645 110
rect 4805 110 4810 140
rect 4840 110 4845 140
rect 4805 100 4845 110
rect 5005 110 5010 140
rect 5040 110 5045 140
rect 5005 100 5045 110
rect 5205 110 5210 140
rect 5240 110 5245 140
rect 5205 100 5245 110
rect 5405 110 5410 140
rect 5440 110 5445 140
rect 5405 100 5445 110
rect 5605 110 5610 140
rect 5640 110 5645 140
rect 5605 100 5645 110
rect 5805 110 5810 140
rect 5840 110 5845 140
rect 5805 100 5845 110
rect 6005 110 6010 140
rect 6040 110 6045 140
rect 6005 100 6045 110
rect 6205 110 6210 140
rect 6240 110 6245 140
rect 6205 100 6245 110
rect 6405 110 6410 140
rect 6440 110 6445 140
rect 6405 100 6445 110
rect -165 80 -30 100
rect 5 80 6570 100
rect -165 70 -155 80
rect -195 40 -190 70
rect -160 40 -155 70
rect 5 70 45 80
rect 5 40 10 70
rect 40 40 45 70
rect 205 70 245 80
rect 205 40 210 70
rect 240 40 245 70
rect 405 70 445 80
rect 405 40 410 70
rect 440 40 445 70
rect 605 70 645 80
rect 605 40 610 70
rect 640 40 645 70
rect 805 70 845 80
rect 805 40 810 70
rect 840 40 845 70
rect 1005 70 1045 80
rect 1005 40 1010 70
rect 1040 40 1045 70
rect 1205 70 1245 80
rect 1205 40 1210 70
rect 1240 40 1245 70
rect 1405 70 1445 80
rect 1405 40 1410 70
rect 1440 40 1445 70
rect 1605 70 1645 80
rect 1605 40 1610 70
rect 1640 40 1645 70
rect 1805 70 1845 80
rect 1805 40 1810 70
rect 1840 40 1845 70
rect 2005 70 2045 80
rect 2005 40 2010 70
rect 2040 40 2045 70
rect 2205 70 2245 80
rect 2205 40 2210 70
rect 2240 40 2245 70
rect 2405 70 2445 80
rect 2405 40 2410 70
rect 2440 40 2445 70
rect 2605 70 2645 80
rect 2605 40 2610 70
rect 2640 40 2645 70
rect 2805 70 2845 80
rect 2805 40 2810 70
rect 2840 40 2845 70
rect 3005 70 3045 80
rect 3005 40 3010 70
rect 3040 40 3045 70
rect 3205 70 3245 80
rect 3205 40 3210 70
rect 3240 40 3245 70
rect 3405 70 3445 80
rect 3405 40 3410 70
rect 3440 40 3445 70
rect 3605 70 3645 80
rect 3605 40 3610 70
rect 3640 40 3645 70
rect 3805 70 3845 80
rect 3805 40 3810 70
rect 3840 40 3845 70
rect 4005 70 4045 80
rect 4005 40 4010 70
rect 4040 40 4045 70
rect 4205 70 4245 80
rect 4205 40 4210 70
rect 4240 40 4245 70
rect 4405 70 4445 80
rect 4405 40 4410 70
rect 4440 40 4445 70
rect 4605 70 4645 80
rect 4605 40 4610 70
rect 4640 40 4645 70
rect 4805 70 4845 80
rect 4805 40 4810 70
rect 4840 40 4845 70
rect 5005 70 5045 80
rect 5005 40 5010 70
rect 5040 40 5045 70
rect 5205 70 5245 80
rect 5205 40 5210 70
rect 5240 40 5245 70
rect 5405 70 5445 80
rect 5405 40 5410 70
rect 5440 40 5445 70
rect 5605 70 5645 80
rect 5605 40 5610 70
rect 5640 40 5645 70
rect 5805 70 5845 80
rect 5805 40 5810 70
rect 5840 40 5845 70
rect 6005 70 6045 80
rect 6005 40 6010 70
rect 6040 40 6045 70
rect 6205 70 6245 80
rect 6205 40 6210 70
rect 6240 40 6245 70
rect 6405 70 6445 80
rect 6405 40 6410 70
rect 6440 40 6445 70
rect -188 -25 -185 40
rect -165 -25 -162 40
rect -188 -45 -162 -25
rect -195 -75 -190 -45
rect -160 -75 -155 -45
rect -195 -85 -155 -75
rect 5 -75 10 -45
rect 40 -75 45 -45
rect 5 -82 45 -75
rect 205 -75 210 -45
rect 240 -75 245 -45
rect 205 -82 245 -75
rect 405 -75 410 -45
rect 440 -75 445 -45
rect 405 -82 445 -75
rect 605 -75 610 -45
rect 640 -75 645 -45
rect 605 -82 645 -75
rect 805 -75 810 -45
rect 840 -75 845 -45
rect 805 -82 845 -75
rect 1005 -75 1010 -45
rect 1040 -75 1045 -45
rect 1005 -82 1045 -75
rect 1205 -75 1210 -45
rect 1240 -75 1245 -45
rect 1205 -82 1245 -75
rect 1405 -75 1410 -45
rect 1440 -75 1445 -45
rect 1405 -82 1445 -75
rect 1605 -75 1610 -45
rect 1640 -75 1645 -45
rect 1605 -82 1645 -75
rect 1805 -75 1810 -45
rect 1840 -75 1845 -45
rect 1805 -82 1845 -75
rect 2005 -75 2010 -45
rect 2040 -75 2045 -45
rect 2005 -82 2045 -75
rect 2205 -75 2210 -45
rect 2240 -75 2245 -45
rect 2205 -82 2245 -75
rect 2405 -75 2410 -45
rect 2440 -75 2445 -45
rect 2405 -82 2445 -75
rect 2605 -75 2610 -45
rect 2640 -75 2645 -45
rect 2605 -82 2645 -75
rect 2805 -75 2810 -45
rect 2840 -75 2845 -45
rect 2805 -82 2845 -75
rect 3005 -75 3010 -45
rect 3040 -75 3045 -45
rect 3005 -82 3045 -75
rect 3205 -75 3210 -45
rect 3240 -75 3245 -45
rect 3205 -82 3245 -75
rect 3405 -75 3410 -45
rect 3440 -75 3445 -45
rect 3405 -82 3445 -75
rect 3605 -75 3610 -45
rect 3640 -75 3645 -45
rect 3605 -82 3645 -75
rect 3805 -75 3810 -45
rect 3840 -75 3845 -45
rect 3805 -82 3845 -75
rect 4005 -75 4010 -45
rect 4040 -75 4045 -45
rect 4005 -82 4045 -75
rect 4205 -75 4210 -45
rect 4240 -75 4245 -45
rect 4205 -82 4245 -75
rect 4405 -75 4410 -45
rect 4440 -75 4445 -45
rect 4405 -82 4445 -75
rect 4605 -75 4610 -45
rect 4640 -75 4645 -45
rect 4605 -82 4645 -75
rect 4805 -75 4810 -45
rect 4840 -75 4845 -45
rect 4805 -82 4845 -75
rect 5005 -75 5010 -45
rect 5040 -75 5045 -45
rect 5005 -82 5045 -75
rect 5205 -75 5210 -45
rect 5240 -75 5245 -45
rect 5205 -82 5245 -75
rect 5405 -75 5410 -45
rect 5440 -75 5445 -45
rect 5405 -82 5445 -75
rect 5605 -75 5610 -45
rect 5640 -75 5645 -45
rect 5605 -82 5645 -75
rect 5805 -75 5810 -45
rect 5840 -75 5845 -45
rect 5805 -82 5845 -75
rect 6005 -75 6010 -45
rect 6040 -75 6045 -45
rect 6005 -82 6045 -75
rect 6205 -75 6210 -45
rect 6240 -75 6245 -45
rect 6205 -82 6245 -75
rect 6405 -75 6410 -45
rect 6440 -75 6445 -45
rect 6405 -82 6445 -75
rect -116 -85 6486 -82
rect -195 -105 -110 -85
rect 6480 -105 6570 -85
rect -195 -115 -155 -105
rect -116 -108 6486 -105
rect -195 -145 -190 -115
rect -160 -145 -155 -115
rect 5 -115 45 -108
rect 5 -145 10 -115
rect 40 -145 45 -115
rect 205 -115 245 -108
rect 205 -145 210 -115
rect 240 -145 245 -115
rect 405 -115 445 -108
rect 405 -145 410 -115
rect 440 -145 445 -115
rect 605 -115 645 -108
rect 605 -145 610 -115
rect 640 -145 645 -115
rect 805 -115 845 -108
rect 805 -145 810 -115
rect 840 -145 845 -115
rect 1005 -115 1045 -108
rect 1005 -145 1010 -115
rect 1040 -145 1045 -115
rect 1205 -115 1245 -108
rect 1205 -145 1210 -115
rect 1240 -145 1245 -115
rect 1405 -115 1445 -108
rect 1405 -145 1410 -115
rect 1440 -145 1445 -115
rect 1605 -115 1645 -108
rect 1605 -145 1610 -115
rect 1640 -145 1645 -115
rect 1805 -115 1845 -108
rect 1805 -145 1810 -115
rect 1840 -145 1845 -115
rect 2005 -115 2045 -108
rect 2005 -145 2010 -115
rect 2040 -145 2045 -115
rect 2205 -115 2245 -108
rect 2205 -145 2210 -115
rect 2240 -145 2245 -115
rect 2405 -115 2445 -108
rect 2405 -145 2410 -115
rect 2440 -145 2445 -115
rect 2605 -115 2645 -108
rect 2605 -145 2610 -115
rect 2640 -145 2645 -115
rect 2805 -115 2845 -108
rect 2805 -145 2810 -115
rect 2840 -145 2845 -115
rect 3005 -115 3045 -108
rect 3005 -145 3010 -115
rect 3040 -145 3045 -115
rect 3205 -115 3245 -108
rect 3205 -145 3210 -115
rect 3240 -145 3245 -115
rect 3405 -115 3445 -108
rect 3405 -145 3410 -115
rect 3440 -145 3445 -115
rect 3605 -115 3645 -108
rect 3605 -145 3610 -115
rect 3640 -145 3645 -115
rect 3805 -115 3845 -108
rect 3805 -145 3810 -115
rect 3840 -145 3845 -115
rect 4005 -115 4045 -108
rect 4005 -145 4010 -115
rect 4040 -145 4045 -115
rect 4205 -115 4245 -108
rect 4205 -145 4210 -115
rect 4240 -145 4245 -115
rect 4405 -115 4445 -108
rect 4405 -145 4410 -115
rect 4440 -145 4445 -115
rect 4605 -115 4645 -108
rect 4605 -145 4610 -115
rect 4640 -145 4645 -115
rect 4805 -115 4845 -108
rect 4805 -145 4810 -115
rect 4840 -145 4845 -115
rect 5005 -115 5045 -108
rect 5005 -145 5010 -115
rect 5040 -145 5045 -115
rect 5205 -115 5245 -108
rect 5205 -145 5210 -115
rect 5240 -145 5245 -115
rect 5405 -115 5445 -108
rect 5405 -145 5410 -115
rect 5440 -145 5445 -115
rect 5605 -115 5645 -108
rect 5605 -145 5610 -115
rect 5640 -145 5645 -115
rect 5805 -115 5845 -108
rect 5805 -145 5810 -115
rect 5840 -145 5845 -115
rect 6005 -115 6045 -108
rect 6005 -145 6010 -115
rect 6040 -145 6045 -115
rect 6205 -115 6245 -108
rect 6205 -145 6210 -115
rect 6240 -145 6245 -115
rect 6405 -115 6445 -108
rect 6405 -145 6410 -115
rect 6440 -145 6445 -115
<< via1 >>
rect -140 12085 -110 12090
rect -140 12065 -135 12085
rect -135 12065 -115 12085
rect -115 12065 -110 12085
rect -140 12060 -110 12065
rect -190 11950 -160 11980
rect -90 12085 -60 12090
rect -90 12065 -85 12085
rect -85 12065 -65 12085
rect -65 12065 -60 12085
rect -90 12060 -60 12065
rect 6460 12060 6490 12065
rect 6460 12040 6465 12060
rect 6465 12040 6485 12060
rect 6485 12040 6490 12060
rect 6460 12035 6490 12040
rect 10 11950 40 11980
rect 210 11950 240 11980
rect 410 11950 440 11980
rect 610 11950 640 11980
rect 810 11950 840 11980
rect 1010 11950 1040 11980
rect 1210 11950 1240 11980
rect 1410 11950 1440 11980
rect 1610 11950 1640 11980
rect 1810 11950 1840 11980
rect 2010 11950 2040 11980
rect 2210 11950 2240 11980
rect 2410 11950 2440 11980
rect 2610 11950 2640 11980
rect 2810 11950 2840 11980
rect 3010 11950 3040 11980
rect 3210 11950 3240 11980
rect 3410 11950 3440 11980
rect 3610 11950 3640 11980
rect 3810 11950 3840 11980
rect 4010 11950 4040 11980
rect 4210 11950 4240 11980
rect 4410 11950 4440 11980
rect 4610 11950 4640 11980
rect 4810 11950 4840 11980
rect 5010 11950 5040 11980
rect 5210 11950 5240 11980
rect 5410 11950 5440 11980
rect 5610 11950 5640 11980
rect 5810 11950 5840 11980
rect 6010 11950 6040 11980
rect 6210 11950 6240 11980
rect 6410 11950 6440 11980
rect 6510 12060 6540 12065
rect 6510 12040 6515 12060
rect 6515 12040 6535 12060
rect 6535 12040 6540 12060
rect 6510 12035 6540 12040
rect -190 11880 -160 11910
rect 10 11880 40 11910
rect 210 11880 240 11910
rect 410 11880 440 11910
rect 610 11880 640 11910
rect 810 11880 840 11910
rect 1010 11880 1040 11910
rect 1210 11880 1240 11910
rect 1410 11880 1440 11910
rect 1610 11880 1640 11910
rect 1810 11880 1840 11910
rect 2010 11880 2040 11910
rect 2210 11880 2240 11910
rect 2410 11880 2440 11910
rect 2610 11880 2640 11910
rect 2810 11880 2840 11910
rect 3010 11880 3040 11910
rect 3210 11880 3240 11910
rect 3410 11880 3440 11910
rect 3610 11880 3640 11910
rect 3810 11880 3840 11910
rect 4010 11880 4040 11910
rect 4210 11880 4240 11910
rect 4410 11880 4440 11910
rect 4610 11880 4640 11910
rect 4810 11880 4840 11910
rect 5010 11880 5040 11910
rect 5210 11880 5240 11910
rect 5410 11880 5440 11910
rect 5610 11880 5640 11910
rect 5810 11880 5840 11910
rect 6010 11880 6040 11910
rect 6210 11880 6240 11910
rect 6410 11880 6440 11910
rect -190 11765 -185 11795
rect -185 11765 -165 11795
rect -165 11765 -160 11795
rect 10 11765 40 11795
rect 210 11765 240 11795
rect 410 11765 440 11795
rect 610 11765 640 11795
rect 810 11765 840 11795
rect 1010 11765 1040 11795
rect 1210 11765 1240 11795
rect 1410 11765 1440 11795
rect 1610 11765 1640 11795
rect 1810 11765 1840 11795
rect 2010 11765 2040 11795
rect 2210 11765 2240 11795
rect 2410 11765 2440 11795
rect 2610 11765 2640 11795
rect 2810 11765 2840 11795
rect 3010 11765 3040 11795
rect 3210 11765 3240 11795
rect 3410 11765 3440 11795
rect 3610 11765 3640 11795
rect 3810 11765 3840 11795
rect 4010 11765 4040 11795
rect 4210 11765 4240 11795
rect 4410 11765 4440 11795
rect 4610 11765 4640 11795
rect 4810 11765 4840 11795
rect 5010 11765 5040 11795
rect 5210 11765 5240 11795
rect 5410 11765 5440 11795
rect 5610 11765 5640 11795
rect 5810 11765 5840 11795
rect 6010 11765 6040 11795
rect 6210 11765 6240 11795
rect 6410 11765 6440 11795
rect -190 11695 -185 11725
rect -185 11695 -165 11725
rect -165 11695 -160 11725
rect 10 11695 40 11725
rect 210 11695 240 11725
rect 410 11695 440 11725
rect 610 11695 640 11725
rect 810 11695 840 11725
rect 1010 11695 1040 11725
rect 1210 11695 1240 11725
rect 1410 11695 1440 11725
rect 1610 11695 1640 11725
rect 1810 11695 1840 11725
rect 2010 11695 2040 11725
rect 2210 11695 2240 11725
rect 2410 11695 2440 11725
rect 2610 11695 2640 11725
rect 2810 11695 2840 11725
rect 3010 11695 3040 11725
rect 3210 11695 3240 11725
rect 3410 11695 3440 11725
rect 3610 11695 3640 11725
rect 3810 11695 3840 11725
rect 4010 11695 4040 11725
rect 4210 11695 4240 11725
rect 4410 11695 4440 11725
rect 4610 11695 4640 11725
rect 4810 11695 4840 11725
rect 5010 11695 5040 11725
rect 5210 11695 5240 11725
rect 5410 11695 5440 11725
rect 5610 11695 5640 11725
rect 5810 11695 5840 11725
rect 6010 11695 6040 11725
rect 6210 11695 6240 11725
rect 6410 11695 6440 11725
rect -190 11580 -185 11610
rect -185 11580 -165 11610
rect -165 11580 -160 11610
rect 10 11580 40 11610
rect 210 11580 240 11610
rect 410 11580 440 11610
rect 610 11580 640 11610
rect 810 11580 840 11610
rect 1010 11580 1040 11610
rect 1210 11580 1240 11610
rect 1410 11580 1440 11610
rect 1610 11580 1640 11610
rect 1810 11580 1840 11610
rect 2010 11580 2040 11610
rect 2210 11580 2240 11610
rect 2410 11580 2440 11610
rect 2610 11580 2640 11610
rect 2810 11580 2840 11610
rect 3010 11580 3040 11610
rect 3210 11580 3240 11610
rect 3410 11580 3440 11610
rect 3610 11580 3640 11610
rect 3810 11580 3840 11610
rect 4010 11580 4040 11610
rect 4210 11580 4240 11610
rect 4410 11580 4440 11610
rect 4610 11580 4640 11610
rect 4810 11580 4840 11610
rect 5010 11580 5040 11610
rect 5210 11580 5240 11610
rect 5410 11580 5440 11610
rect 5610 11580 5640 11610
rect 5810 11580 5840 11610
rect 6010 11580 6040 11610
rect 6210 11580 6240 11610
rect 6410 11580 6440 11610
rect -190 11510 -185 11540
rect -185 11510 -165 11540
rect -165 11510 -160 11540
rect 10 11510 40 11540
rect 210 11510 240 11540
rect 410 11510 440 11540
rect 610 11510 640 11540
rect 810 11510 840 11540
rect 1010 11510 1040 11540
rect 1210 11510 1240 11540
rect 1410 11510 1440 11540
rect 1610 11510 1640 11540
rect 1810 11510 1840 11540
rect 2010 11510 2040 11540
rect 2210 11510 2240 11540
rect 2410 11510 2440 11540
rect 2610 11510 2640 11540
rect 2810 11510 2840 11540
rect 3010 11510 3040 11540
rect 3210 11510 3240 11540
rect 3410 11510 3440 11540
rect 3610 11510 3640 11540
rect 3810 11510 3840 11540
rect 4010 11510 4040 11540
rect 4210 11510 4240 11540
rect 4410 11510 4440 11540
rect 4610 11510 4640 11540
rect 4810 11510 4840 11540
rect 5010 11510 5040 11540
rect 5210 11510 5240 11540
rect 5410 11510 5440 11540
rect 5610 11510 5640 11540
rect 5810 11510 5840 11540
rect 6010 11510 6040 11540
rect 6210 11510 6240 11540
rect 6410 11510 6440 11540
rect -190 11395 -185 11425
rect -185 11395 -165 11425
rect -165 11395 -160 11425
rect 10 11395 40 11425
rect 210 11395 240 11425
rect 410 11395 440 11425
rect 610 11395 640 11425
rect 810 11395 840 11425
rect 1010 11395 1040 11425
rect 1210 11395 1240 11425
rect 1410 11395 1440 11425
rect 1610 11395 1640 11425
rect 1810 11395 1840 11425
rect 2010 11395 2040 11425
rect 2210 11395 2240 11425
rect 2410 11395 2440 11425
rect 2610 11395 2640 11425
rect 2810 11395 2840 11425
rect 3010 11395 3040 11425
rect 3210 11395 3240 11425
rect 3410 11395 3440 11425
rect 3610 11395 3640 11425
rect 3810 11395 3840 11425
rect 4010 11395 4040 11425
rect 4210 11395 4240 11425
rect 4410 11395 4440 11425
rect 4610 11395 4640 11425
rect 4810 11395 4840 11425
rect 5010 11395 5040 11425
rect 5210 11395 5240 11425
rect 5410 11395 5440 11425
rect 5610 11395 5640 11425
rect 5810 11395 5840 11425
rect 6010 11395 6040 11425
rect 6210 11395 6240 11425
rect 6410 11395 6440 11425
rect -190 11325 -185 11355
rect -185 11325 -165 11355
rect -165 11325 -160 11355
rect 10 11325 40 11355
rect 210 11325 240 11355
rect 410 11325 440 11355
rect 610 11325 640 11355
rect 810 11325 840 11355
rect 1010 11325 1040 11355
rect 1210 11325 1240 11355
rect 1410 11325 1440 11355
rect 1610 11325 1640 11355
rect 1810 11325 1840 11355
rect 2010 11325 2040 11355
rect 2210 11325 2240 11355
rect 2410 11325 2440 11355
rect 2610 11325 2640 11355
rect 2810 11325 2840 11355
rect 3010 11325 3040 11355
rect 3210 11325 3240 11355
rect 3410 11325 3440 11355
rect 3610 11325 3640 11355
rect 3810 11325 3840 11355
rect 4010 11325 4040 11355
rect 4210 11325 4240 11355
rect 4410 11325 4440 11355
rect 4610 11325 4640 11355
rect 4810 11325 4840 11355
rect 5010 11325 5040 11355
rect 5210 11325 5240 11355
rect 5410 11325 5440 11355
rect 5610 11325 5640 11355
rect 5810 11325 5840 11355
rect 6010 11325 6040 11355
rect 6210 11325 6240 11355
rect 6410 11325 6440 11355
rect -190 11210 -185 11240
rect -185 11210 -165 11240
rect -165 11210 -160 11240
rect 10 11210 40 11240
rect 210 11210 240 11240
rect 410 11210 440 11240
rect 610 11210 640 11240
rect 810 11210 840 11240
rect 1010 11210 1040 11240
rect 1210 11210 1240 11240
rect 1410 11210 1440 11240
rect 1610 11210 1640 11240
rect 1810 11210 1840 11240
rect 2010 11210 2040 11240
rect 2210 11210 2240 11240
rect 2410 11210 2440 11240
rect 2610 11210 2640 11240
rect 2810 11210 2840 11240
rect 3010 11210 3040 11240
rect 3210 11210 3240 11240
rect 3410 11210 3440 11240
rect 3610 11210 3640 11240
rect 3810 11210 3840 11240
rect 4010 11210 4040 11240
rect 4210 11210 4240 11240
rect 4410 11210 4440 11240
rect 4610 11210 4640 11240
rect 4810 11210 4840 11240
rect 5010 11210 5040 11240
rect 5210 11210 5240 11240
rect 5410 11210 5440 11240
rect 5610 11210 5640 11240
rect 5810 11210 5840 11240
rect 6010 11210 6040 11240
rect 6210 11210 6240 11240
rect 6410 11210 6440 11240
rect -190 11140 -185 11170
rect -185 11140 -165 11170
rect -165 11140 -160 11170
rect 10 11140 40 11170
rect 210 11140 240 11170
rect 410 11140 440 11170
rect 610 11140 640 11170
rect 810 11140 840 11170
rect 1010 11140 1040 11170
rect 1210 11140 1240 11170
rect 1410 11140 1440 11170
rect 1610 11140 1640 11170
rect 1810 11140 1840 11170
rect 2010 11140 2040 11170
rect 2210 11140 2240 11170
rect 2410 11140 2440 11170
rect 2610 11140 2640 11170
rect 2810 11140 2840 11170
rect 3010 11140 3040 11170
rect 3210 11140 3240 11170
rect 3410 11140 3440 11170
rect 3610 11140 3640 11170
rect 3810 11140 3840 11170
rect 4010 11140 4040 11170
rect 4210 11140 4240 11170
rect 4410 11140 4440 11170
rect 4610 11140 4640 11170
rect 4810 11140 4840 11170
rect 5010 11140 5040 11170
rect 5210 11140 5240 11170
rect 5410 11140 5440 11170
rect 5610 11140 5640 11170
rect 5810 11140 5840 11170
rect 6010 11140 6040 11170
rect 6210 11140 6240 11170
rect 6410 11140 6440 11170
rect -190 11025 -185 11055
rect -185 11025 -165 11055
rect -165 11025 -160 11055
rect 10 11025 40 11055
rect 210 11025 240 11055
rect 410 11025 440 11055
rect 610 11025 640 11055
rect 810 11025 840 11055
rect 1010 11025 1040 11055
rect 1210 11025 1240 11055
rect 1410 11025 1440 11055
rect 1610 11025 1640 11055
rect 1810 11025 1840 11055
rect 2010 11025 2040 11055
rect 2210 11025 2240 11055
rect 2410 11025 2440 11055
rect 2610 11025 2640 11055
rect 2810 11025 2840 11055
rect 3010 11025 3040 11055
rect 3210 11025 3240 11055
rect 3410 11025 3440 11055
rect 3610 11025 3640 11055
rect 3810 11025 3840 11055
rect 4010 11025 4040 11055
rect 4210 11025 4240 11055
rect 4410 11025 4440 11055
rect 4610 11025 4640 11055
rect 4810 11025 4840 11055
rect 5010 11025 5040 11055
rect 5210 11025 5240 11055
rect 5410 11025 5440 11055
rect 5610 11025 5640 11055
rect 5810 11025 5840 11055
rect 6010 11025 6040 11055
rect 6210 11025 6240 11055
rect 6410 11025 6440 11055
rect -190 10955 -185 10985
rect -185 10955 -165 10985
rect -165 10955 -160 10985
rect 10 10955 40 10985
rect 210 10955 240 10985
rect 410 10955 440 10985
rect 610 10955 640 10985
rect 810 10955 840 10985
rect 1010 10955 1040 10985
rect 1210 10955 1240 10985
rect 1410 10955 1440 10985
rect 1610 10955 1640 10985
rect 1810 10955 1840 10985
rect 2010 10955 2040 10985
rect 2210 10955 2240 10985
rect 2410 10955 2440 10985
rect 2610 10955 2640 10985
rect 2810 10955 2840 10985
rect 3010 10955 3040 10985
rect 3210 10955 3240 10985
rect 3410 10955 3440 10985
rect 3610 10955 3640 10985
rect 3810 10955 3840 10985
rect 4010 10955 4040 10985
rect 4210 10955 4240 10985
rect 4410 10955 4440 10985
rect 4610 10955 4640 10985
rect 4810 10955 4840 10985
rect 5010 10955 5040 10985
rect 5210 10955 5240 10985
rect 5410 10955 5440 10985
rect 5610 10955 5640 10985
rect 5810 10955 5840 10985
rect 6010 10955 6040 10985
rect 6210 10955 6240 10985
rect 6410 10955 6440 10985
rect -190 10840 -185 10870
rect -185 10840 -165 10870
rect -165 10840 -160 10870
rect 10 10840 40 10870
rect 210 10840 240 10870
rect 410 10840 440 10870
rect 610 10840 640 10870
rect 810 10840 840 10870
rect 1010 10840 1040 10870
rect 1210 10840 1240 10870
rect 1410 10840 1440 10870
rect 1610 10840 1640 10870
rect 1810 10840 1840 10870
rect 2010 10840 2040 10870
rect 2210 10840 2240 10870
rect 2410 10840 2440 10870
rect 2610 10840 2640 10870
rect 2810 10840 2840 10870
rect 3010 10840 3040 10870
rect 3210 10840 3240 10870
rect 3410 10840 3440 10870
rect 3610 10840 3640 10870
rect 3810 10840 3840 10870
rect 4010 10840 4040 10870
rect 4210 10840 4240 10870
rect 4410 10840 4440 10870
rect 4610 10840 4640 10870
rect 4810 10840 4840 10870
rect 5010 10840 5040 10870
rect 5210 10840 5240 10870
rect 5410 10840 5440 10870
rect 5610 10840 5640 10870
rect 5810 10840 5840 10870
rect 6010 10840 6040 10870
rect 6210 10840 6240 10870
rect 6410 10840 6440 10870
rect -190 10770 -185 10800
rect -185 10770 -165 10800
rect -165 10770 -160 10800
rect 10 10770 40 10800
rect 210 10770 240 10800
rect 410 10770 440 10800
rect 610 10770 640 10800
rect 810 10770 840 10800
rect 1010 10770 1040 10800
rect 1210 10770 1240 10800
rect 1410 10770 1440 10800
rect 1610 10770 1640 10800
rect 1810 10770 1840 10800
rect 2010 10770 2040 10800
rect 2210 10770 2240 10800
rect 2410 10770 2440 10800
rect 2610 10770 2640 10800
rect 2810 10770 2840 10800
rect 3010 10770 3040 10800
rect 3210 10770 3240 10800
rect 3410 10770 3440 10800
rect 3610 10770 3640 10800
rect 3810 10770 3840 10800
rect 4010 10770 4040 10800
rect 4210 10770 4240 10800
rect 4410 10770 4440 10800
rect 4610 10770 4640 10800
rect 4810 10770 4840 10800
rect 5010 10770 5040 10800
rect 5210 10770 5240 10800
rect 5410 10770 5440 10800
rect 5610 10770 5640 10800
rect 5810 10770 5840 10800
rect 6010 10770 6040 10800
rect 6210 10770 6240 10800
rect 6410 10770 6440 10800
rect -190 10655 -185 10685
rect -185 10655 -165 10685
rect -165 10655 -160 10685
rect 10 10655 40 10685
rect 210 10655 240 10685
rect 410 10655 440 10685
rect 610 10655 640 10685
rect 810 10655 840 10685
rect 1010 10655 1040 10685
rect 1210 10655 1240 10685
rect 1410 10655 1440 10685
rect 1610 10655 1640 10685
rect 1810 10655 1840 10685
rect 2010 10655 2040 10685
rect 2210 10655 2240 10685
rect 2410 10655 2440 10685
rect 2610 10655 2640 10685
rect 2810 10655 2840 10685
rect 3010 10655 3040 10685
rect 3210 10655 3240 10685
rect 3410 10655 3440 10685
rect 3610 10655 3640 10685
rect 3810 10655 3840 10685
rect 4010 10655 4040 10685
rect 4210 10655 4240 10685
rect 4410 10655 4440 10685
rect 4610 10655 4640 10685
rect 4810 10655 4840 10685
rect 5010 10655 5040 10685
rect 5210 10655 5240 10685
rect 5410 10655 5440 10685
rect 5610 10655 5640 10685
rect 5810 10655 5840 10685
rect 6010 10655 6040 10685
rect 6210 10655 6240 10685
rect 6410 10655 6440 10685
rect -190 10585 -185 10615
rect -185 10585 -165 10615
rect -165 10585 -160 10615
rect 10 10585 40 10615
rect 210 10585 240 10615
rect 410 10585 440 10615
rect 610 10585 640 10615
rect 810 10585 840 10615
rect 1010 10585 1040 10615
rect 1210 10585 1240 10615
rect 1410 10585 1440 10615
rect 1610 10585 1640 10615
rect 1810 10585 1840 10615
rect 2010 10585 2040 10615
rect 2210 10585 2240 10615
rect 2410 10585 2440 10615
rect 2610 10585 2640 10615
rect 2810 10585 2840 10615
rect 3010 10585 3040 10615
rect 3210 10585 3240 10615
rect 3410 10585 3440 10615
rect 3610 10585 3640 10615
rect 3810 10585 3840 10615
rect 4010 10585 4040 10615
rect 4210 10585 4240 10615
rect 4410 10585 4440 10615
rect 4610 10585 4640 10615
rect 4810 10585 4840 10615
rect 5010 10585 5040 10615
rect 5210 10585 5240 10615
rect 5410 10585 5440 10615
rect 5610 10585 5640 10615
rect 5810 10585 5840 10615
rect 6010 10585 6040 10615
rect 6210 10585 6240 10615
rect 6410 10585 6440 10615
rect -190 10470 -185 10500
rect -185 10470 -165 10500
rect -165 10470 -160 10500
rect 10 10470 40 10500
rect 210 10470 240 10500
rect 410 10470 440 10500
rect 610 10470 640 10500
rect 810 10470 840 10500
rect 1010 10470 1040 10500
rect 1210 10470 1240 10500
rect 1410 10470 1440 10500
rect 1610 10470 1640 10500
rect 1810 10470 1840 10500
rect 2010 10470 2040 10500
rect 2210 10470 2240 10500
rect 2410 10470 2440 10500
rect 2610 10470 2640 10500
rect 2810 10470 2840 10500
rect 3010 10470 3040 10500
rect 3210 10470 3240 10500
rect 3410 10470 3440 10500
rect 3610 10470 3640 10500
rect 3810 10470 3840 10500
rect 4010 10470 4040 10500
rect 4210 10470 4240 10500
rect 4410 10470 4440 10500
rect 4610 10470 4640 10500
rect 4810 10470 4840 10500
rect 5010 10470 5040 10500
rect 5210 10470 5240 10500
rect 5410 10470 5440 10500
rect 5610 10470 5640 10500
rect 5810 10470 5840 10500
rect 6010 10470 6040 10500
rect 6210 10470 6240 10500
rect 6410 10470 6440 10500
rect -190 10400 -185 10430
rect -185 10400 -165 10430
rect -165 10400 -160 10430
rect 10 10400 40 10430
rect 210 10400 240 10430
rect 410 10400 440 10430
rect 610 10400 640 10430
rect 810 10400 840 10430
rect 1010 10400 1040 10430
rect 1210 10400 1240 10430
rect 1410 10400 1440 10430
rect 1610 10400 1640 10430
rect 1810 10400 1840 10430
rect 2010 10400 2040 10430
rect 2210 10400 2240 10430
rect 2410 10400 2440 10430
rect 2610 10400 2640 10430
rect 2810 10400 2840 10430
rect 3010 10400 3040 10430
rect 3210 10400 3240 10430
rect 3410 10400 3440 10430
rect 3610 10400 3640 10430
rect 3810 10400 3840 10430
rect 4010 10400 4040 10430
rect 4210 10400 4240 10430
rect 4410 10400 4440 10430
rect 4610 10400 4640 10430
rect 4810 10400 4840 10430
rect 5010 10400 5040 10430
rect 5210 10400 5240 10430
rect 5410 10400 5440 10430
rect 5610 10400 5640 10430
rect 5810 10400 5840 10430
rect 6010 10400 6040 10430
rect 6210 10400 6240 10430
rect 6410 10400 6440 10430
rect -190 10285 -185 10315
rect -185 10285 -165 10315
rect -165 10285 -160 10315
rect 10 10285 40 10315
rect 210 10285 240 10315
rect 410 10285 440 10315
rect 610 10285 640 10315
rect 810 10285 840 10315
rect 1010 10285 1040 10315
rect 1210 10285 1240 10315
rect 1410 10285 1440 10315
rect 1610 10285 1640 10315
rect 1810 10285 1840 10315
rect 2010 10285 2040 10315
rect 2210 10285 2240 10315
rect 2410 10285 2440 10315
rect 2610 10285 2640 10315
rect 2810 10285 2840 10315
rect 3010 10285 3040 10315
rect 3210 10285 3240 10315
rect 3410 10285 3440 10315
rect 3610 10285 3640 10315
rect 3810 10285 3840 10315
rect 4010 10285 4040 10315
rect 4210 10285 4240 10315
rect 4410 10285 4440 10315
rect 4610 10285 4640 10315
rect 4810 10285 4840 10315
rect 5010 10285 5040 10315
rect 5210 10285 5240 10315
rect 5410 10285 5440 10315
rect 5610 10285 5640 10315
rect 5810 10285 5840 10315
rect 6010 10285 6040 10315
rect 6210 10285 6240 10315
rect 6410 10285 6440 10315
rect -190 10215 -185 10245
rect -185 10215 -165 10245
rect -165 10215 -160 10245
rect 10 10215 40 10245
rect 210 10215 240 10245
rect 410 10215 440 10245
rect 610 10215 640 10245
rect 810 10215 840 10245
rect 1010 10215 1040 10245
rect 1210 10215 1240 10245
rect 1410 10215 1440 10245
rect 1610 10215 1640 10245
rect 1810 10215 1840 10245
rect 2010 10215 2040 10245
rect 2210 10215 2240 10245
rect 2410 10215 2440 10245
rect 2610 10215 2640 10245
rect 2810 10215 2840 10245
rect 3010 10215 3040 10245
rect 3210 10215 3240 10245
rect 3410 10215 3440 10245
rect 3610 10215 3640 10245
rect 3810 10215 3840 10245
rect 4010 10215 4040 10245
rect 4210 10215 4240 10245
rect 4410 10215 4440 10245
rect 4610 10215 4640 10245
rect 4810 10215 4840 10245
rect 5010 10215 5040 10245
rect 5210 10215 5240 10245
rect 5410 10215 5440 10245
rect 5610 10215 5640 10245
rect 5810 10215 5840 10245
rect 6010 10215 6040 10245
rect 6210 10215 6240 10245
rect 6410 10215 6440 10245
rect -190 10100 -185 10130
rect -185 10100 -165 10130
rect -165 10100 -160 10130
rect 10 10100 40 10130
rect 210 10100 240 10130
rect 410 10100 440 10130
rect 610 10100 640 10130
rect 810 10100 840 10130
rect 1010 10100 1040 10130
rect 1210 10100 1240 10130
rect 1410 10100 1440 10130
rect 1610 10100 1640 10130
rect 1810 10100 1840 10130
rect 2010 10100 2040 10130
rect 2210 10100 2240 10130
rect 2410 10100 2440 10130
rect 2610 10100 2640 10130
rect 2810 10100 2840 10130
rect 3010 10100 3040 10130
rect 3210 10100 3240 10130
rect 3410 10100 3440 10130
rect 3610 10100 3640 10130
rect 3810 10100 3840 10130
rect 4010 10100 4040 10130
rect 4210 10100 4240 10130
rect 4410 10100 4440 10130
rect 4610 10100 4640 10130
rect 4810 10100 4840 10130
rect 5010 10100 5040 10130
rect 5210 10100 5240 10130
rect 5410 10100 5440 10130
rect 5610 10100 5640 10130
rect 5810 10100 5840 10130
rect 6010 10100 6040 10130
rect 6210 10100 6240 10130
rect 6410 10100 6440 10130
rect -190 10030 -185 10060
rect -185 10030 -165 10060
rect -165 10030 -160 10060
rect 10 10030 40 10060
rect 210 10030 240 10060
rect 410 10030 440 10060
rect 610 10030 640 10060
rect 810 10030 840 10060
rect 1010 10030 1040 10060
rect 1210 10030 1240 10060
rect 1410 10030 1440 10060
rect 1610 10030 1640 10060
rect 1810 10030 1840 10060
rect 2010 10030 2040 10060
rect 2210 10030 2240 10060
rect 2410 10030 2440 10060
rect 2610 10030 2640 10060
rect 2810 10030 2840 10060
rect 3010 10030 3040 10060
rect 3210 10030 3240 10060
rect 3410 10030 3440 10060
rect 3610 10030 3640 10060
rect 3810 10030 3840 10060
rect 4010 10030 4040 10060
rect 4210 10030 4240 10060
rect 4410 10030 4440 10060
rect 4610 10030 4640 10060
rect 4810 10030 4840 10060
rect 5010 10030 5040 10060
rect 5210 10030 5240 10060
rect 5410 10030 5440 10060
rect 5610 10030 5640 10060
rect 5810 10030 5840 10060
rect 6010 10030 6040 10060
rect 6210 10030 6240 10060
rect 6410 10030 6440 10060
rect -190 9915 -185 9945
rect -185 9915 -165 9945
rect -165 9915 -160 9945
rect 10 9915 40 9945
rect 210 9915 240 9945
rect 410 9915 440 9945
rect 610 9915 640 9945
rect 810 9915 840 9945
rect 1010 9915 1040 9945
rect 1210 9915 1240 9945
rect 1410 9915 1440 9945
rect 1610 9915 1640 9945
rect 1810 9915 1840 9945
rect 2010 9915 2040 9945
rect 2210 9915 2240 9945
rect 2410 9915 2440 9945
rect 2610 9915 2640 9945
rect 2810 9915 2840 9945
rect 3010 9915 3040 9945
rect 3210 9915 3240 9945
rect 3410 9915 3440 9945
rect 3610 9915 3640 9945
rect 3810 9915 3840 9945
rect 4010 9915 4040 9945
rect 4210 9915 4240 9945
rect 4410 9915 4440 9945
rect 4610 9915 4640 9945
rect 4810 9915 4840 9945
rect 5010 9915 5040 9945
rect 5210 9915 5240 9945
rect 5410 9915 5440 9945
rect 5610 9915 5640 9945
rect 5810 9915 5840 9945
rect 6010 9915 6040 9945
rect 6210 9915 6240 9945
rect 6410 9915 6440 9945
rect -190 9845 -185 9875
rect -185 9845 -165 9875
rect -165 9845 -160 9875
rect 10 9845 40 9875
rect 210 9845 240 9875
rect 410 9845 440 9875
rect 610 9845 640 9875
rect 810 9845 840 9875
rect 1010 9845 1040 9875
rect 1210 9845 1240 9875
rect 1410 9845 1440 9875
rect 1610 9845 1640 9875
rect 1810 9845 1840 9875
rect 2010 9845 2040 9875
rect 2210 9845 2240 9875
rect 2410 9845 2440 9875
rect 2610 9845 2640 9875
rect 2810 9845 2840 9875
rect 3010 9845 3040 9875
rect 3210 9845 3240 9875
rect 3410 9845 3440 9875
rect 3610 9845 3640 9875
rect 3810 9845 3840 9875
rect 4010 9845 4040 9875
rect 4210 9845 4240 9875
rect 4410 9845 4440 9875
rect 4610 9845 4640 9875
rect 4810 9845 4840 9875
rect 5010 9845 5040 9875
rect 5210 9845 5240 9875
rect 5410 9845 5440 9875
rect 5610 9845 5640 9875
rect 5810 9845 5840 9875
rect 6010 9845 6040 9875
rect 6210 9845 6240 9875
rect 6410 9845 6440 9875
rect -190 9730 -185 9760
rect -185 9730 -165 9760
rect -165 9730 -160 9760
rect 10 9730 40 9760
rect 210 9730 240 9760
rect 410 9730 440 9760
rect 610 9730 640 9760
rect 810 9730 840 9760
rect 1010 9730 1040 9760
rect 1210 9730 1240 9760
rect 1410 9730 1440 9760
rect 1610 9730 1640 9760
rect 1810 9730 1840 9760
rect 2010 9730 2040 9760
rect 2210 9730 2240 9760
rect 2410 9730 2440 9760
rect 2610 9730 2640 9760
rect 2810 9730 2840 9760
rect 3010 9730 3040 9760
rect 3210 9730 3240 9760
rect 3410 9730 3440 9760
rect 3610 9730 3640 9760
rect 3810 9730 3840 9760
rect 4010 9730 4040 9760
rect 4210 9730 4240 9760
rect 4410 9730 4440 9760
rect 4610 9730 4640 9760
rect 4810 9730 4840 9760
rect 5010 9730 5040 9760
rect 5210 9730 5240 9760
rect 5410 9730 5440 9760
rect 5610 9730 5640 9760
rect 5810 9730 5840 9760
rect 6010 9730 6040 9760
rect 6210 9730 6240 9760
rect 6410 9730 6440 9760
rect -190 9660 -185 9690
rect -185 9660 -165 9690
rect -165 9660 -160 9690
rect 10 9660 40 9690
rect 210 9660 240 9690
rect 410 9660 440 9690
rect 610 9660 640 9690
rect 810 9660 840 9690
rect 1010 9660 1040 9690
rect 1210 9660 1240 9690
rect 1410 9660 1440 9690
rect 1610 9660 1640 9690
rect 1810 9660 1840 9690
rect 2010 9660 2040 9690
rect 2210 9660 2240 9690
rect 2410 9660 2440 9690
rect 2610 9660 2640 9690
rect 2810 9660 2840 9690
rect 3010 9660 3040 9690
rect 3210 9660 3240 9690
rect 3410 9660 3440 9690
rect 3610 9660 3640 9690
rect 3810 9660 3840 9690
rect 4010 9660 4040 9690
rect 4210 9660 4240 9690
rect 4410 9660 4440 9690
rect 4610 9660 4640 9690
rect 4810 9660 4840 9690
rect 5010 9660 5040 9690
rect 5210 9660 5240 9690
rect 5410 9660 5440 9690
rect 5610 9660 5640 9690
rect 5810 9660 5840 9690
rect 6010 9660 6040 9690
rect 6210 9660 6240 9690
rect 6410 9660 6440 9690
rect -190 9545 -185 9575
rect -185 9545 -165 9575
rect -165 9545 -160 9575
rect 10 9545 40 9575
rect 210 9545 240 9575
rect 410 9545 440 9575
rect 610 9545 640 9575
rect 810 9545 840 9575
rect 1010 9545 1040 9575
rect 1210 9545 1240 9575
rect 1410 9545 1440 9575
rect 1610 9545 1640 9575
rect 1810 9545 1840 9575
rect 2010 9545 2040 9575
rect 2210 9545 2240 9575
rect 2410 9545 2440 9575
rect 2610 9545 2640 9575
rect 2810 9545 2840 9575
rect 3010 9545 3040 9575
rect 3210 9545 3240 9575
rect 3410 9545 3440 9575
rect 3610 9545 3640 9575
rect 3810 9545 3840 9575
rect 4010 9545 4040 9575
rect 4210 9545 4240 9575
rect 4410 9545 4440 9575
rect 4610 9545 4640 9575
rect 4810 9545 4840 9575
rect 5010 9545 5040 9575
rect 5210 9545 5240 9575
rect 5410 9545 5440 9575
rect 5610 9545 5640 9575
rect 5810 9545 5840 9575
rect 6010 9545 6040 9575
rect 6210 9545 6240 9575
rect 6410 9545 6440 9575
rect -190 9475 -185 9505
rect -185 9475 -165 9505
rect -165 9475 -160 9505
rect 10 9475 40 9505
rect 210 9475 240 9505
rect 410 9475 440 9505
rect 610 9475 640 9505
rect 810 9475 840 9505
rect 1010 9475 1040 9505
rect 1210 9475 1240 9505
rect 1410 9475 1440 9505
rect 1610 9475 1640 9505
rect 1810 9475 1840 9505
rect 2010 9475 2040 9505
rect 2210 9475 2240 9505
rect 2410 9475 2440 9505
rect 2610 9475 2640 9505
rect 2810 9475 2840 9505
rect 3010 9475 3040 9505
rect 3210 9475 3240 9505
rect 3410 9475 3440 9505
rect 3610 9475 3640 9505
rect 3810 9475 3840 9505
rect 4010 9475 4040 9505
rect 4210 9475 4240 9505
rect 4410 9475 4440 9505
rect 4610 9475 4640 9505
rect 4810 9475 4840 9505
rect 5010 9475 5040 9505
rect 5210 9475 5240 9505
rect 5410 9475 5440 9505
rect 5610 9475 5640 9505
rect 5810 9475 5840 9505
rect 6010 9475 6040 9505
rect 6210 9475 6240 9505
rect 6410 9475 6440 9505
rect -190 9360 -185 9390
rect -185 9360 -165 9390
rect -165 9360 -160 9390
rect 10 9360 40 9390
rect 210 9360 240 9390
rect 410 9360 440 9390
rect 610 9360 640 9390
rect 810 9360 840 9390
rect 1010 9360 1040 9390
rect 1210 9360 1240 9390
rect 1410 9360 1440 9390
rect 1610 9360 1640 9390
rect 1810 9360 1840 9390
rect 2010 9360 2040 9390
rect 2210 9360 2240 9390
rect 2410 9360 2440 9390
rect 2610 9360 2640 9390
rect 2810 9360 2840 9390
rect 3010 9360 3040 9390
rect 3210 9360 3240 9390
rect 3410 9360 3440 9390
rect 3610 9360 3640 9390
rect 3810 9360 3840 9390
rect 4010 9360 4040 9390
rect 4210 9360 4240 9390
rect 4410 9360 4440 9390
rect 4610 9360 4640 9390
rect 4810 9360 4840 9390
rect 5010 9360 5040 9390
rect 5210 9360 5240 9390
rect 5410 9360 5440 9390
rect 5610 9360 5640 9390
rect 5810 9360 5840 9390
rect 6010 9360 6040 9390
rect 6210 9360 6240 9390
rect 6410 9360 6440 9390
rect -190 9290 -185 9320
rect -185 9290 -165 9320
rect -165 9290 -160 9320
rect 10 9290 40 9320
rect 210 9290 240 9320
rect 410 9290 440 9320
rect 610 9290 640 9320
rect 810 9290 840 9320
rect 1010 9290 1040 9320
rect 1210 9290 1240 9320
rect 1410 9290 1440 9320
rect 1610 9290 1640 9320
rect 1810 9290 1840 9320
rect 2010 9290 2040 9320
rect 2210 9290 2240 9320
rect 2410 9290 2440 9320
rect 2610 9290 2640 9320
rect 2810 9290 2840 9320
rect 3010 9290 3040 9320
rect 3210 9290 3240 9320
rect 3410 9290 3440 9320
rect 3610 9290 3640 9320
rect 3810 9290 3840 9320
rect 4010 9290 4040 9320
rect 4210 9290 4240 9320
rect 4410 9290 4440 9320
rect 4610 9290 4640 9320
rect 4810 9290 4840 9320
rect 5010 9290 5040 9320
rect 5210 9290 5240 9320
rect 5410 9290 5440 9320
rect 5610 9290 5640 9320
rect 5810 9290 5840 9320
rect 6010 9290 6040 9320
rect 6210 9290 6240 9320
rect 6410 9290 6440 9320
rect -190 9175 -185 9205
rect -185 9175 -165 9205
rect -165 9175 -160 9205
rect 10 9175 40 9205
rect 210 9175 240 9205
rect 410 9175 440 9205
rect 610 9175 640 9205
rect 810 9175 840 9205
rect 1010 9175 1040 9205
rect 1210 9175 1240 9205
rect 1410 9175 1440 9205
rect 1610 9175 1640 9205
rect 1810 9175 1840 9205
rect 2010 9175 2040 9205
rect 2210 9175 2240 9205
rect 2410 9175 2440 9205
rect 2610 9175 2640 9205
rect 2810 9175 2840 9205
rect 3010 9175 3040 9205
rect 3210 9175 3240 9205
rect 3410 9175 3440 9205
rect 3610 9175 3640 9205
rect 3810 9175 3840 9205
rect 4010 9175 4040 9205
rect 4210 9175 4240 9205
rect 4410 9175 4440 9205
rect 4610 9175 4640 9205
rect 4810 9175 4840 9205
rect 5010 9175 5040 9205
rect 5210 9175 5240 9205
rect 5410 9175 5440 9205
rect 5610 9175 5640 9205
rect 5810 9175 5840 9205
rect 6010 9175 6040 9205
rect 6210 9175 6240 9205
rect 6410 9175 6440 9205
rect -190 9105 -185 9135
rect -185 9105 -165 9135
rect -165 9105 -160 9135
rect 10 9105 40 9135
rect 210 9105 240 9135
rect 410 9105 440 9135
rect 610 9105 640 9135
rect 810 9105 840 9135
rect 1010 9105 1040 9135
rect 1210 9105 1240 9135
rect 1410 9105 1440 9135
rect 1610 9105 1640 9135
rect 1810 9105 1840 9135
rect 2010 9105 2040 9135
rect 2210 9105 2240 9135
rect 2410 9105 2440 9135
rect 2610 9105 2640 9135
rect 2810 9105 2840 9135
rect 3010 9105 3040 9135
rect 3210 9105 3240 9135
rect 3410 9105 3440 9135
rect 3610 9105 3640 9135
rect 3810 9105 3840 9135
rect 4010 9105 4040 9135
rect 4210 9105 4240 9135
rect 4410 9105 4440 9135
rect 4610 9105 4640 9135
rect 4810 9105 4840 9135
rect 5010 9105 5040 9135
rect 5210 9105 5240 9135
rect 5410 9105 5440 9135
rect 5610 9105 5640 9135
rect 5810 9105 5840 9135
rect 6010 9105 6040 9135
rect 6210 9105 6240 9135
rect 6410 9105 6440 9135
rect -190 8990 -185 9020
rect -185 8990 -165 9020
rect -165 8990 -160 9020
rect 10 8990 40 9020
rect 210 8990 240 9020
rect 410 8990 440 9020
rect 610 8990 640 9020
rect 810 8990 840 9020
rect 1010 8990 1040 9020
rect 1210 8990 1240 9020
rect 1410 8990 1440 9020
rect 1610 8990 1640 9020
rect 1810 8990 1840 9020
rect 2010 8990 2040 9020
rect 2210 8990 2240 9020
rect 2410 8990 2440 9020
rect 2610 8990 2640 9020
rect 2810 8990 2840 9020
rect 3010 8990 3040 9020
rect 3210 8990 3240 9020
rect 3410 8990 3440 9020
rect 3610 8990 3640 9020
rect 3810 8990 3840 9020
rect 4010 8990 4040 9020
rect 4210 8990 4240 9020
rect 4410 8990 4440 9020
rect 4610 8990 4640 9020
rect 4810 8990 4840 9020
rect 5010 8990 5040 9020
rect 5210 8990 5240 9020
rect 5410 8990 5440 9020
rect 5610 8990 5640 9020
rect 5810 8990 5840 9020
rect 6010 8990 6040 9020
rect 6210 8990 6240 9020
rect 6410 8990 6440 9020
rect -190 8920 -185 8950
rect -185 8920 -165 8950
rect -165 8920 -160 8950
rect 10 8920 40 8950
rect 210 8920 240 8950
rect 410 8920 440 8950
rect 610 8920 640 8950
rect 810 8920 840 8950
rect 1010 8920 1040 8950
rect 1210 8920 1240 8950
rect 1410 8920 1440 8950
rect 1610 8920 1640 8950
rect 1810 8920 1840 8950
rect 2010 8920 2040 8950
rect 2210 8920 2240 8950
rect 2410 8920 2440 8950
rect 2610 8920 2640 8950
rect 2810 8920 2840 8950
rect 3010 8920 3040 8950
rect 3210 8920 3240 8950
rect 3410 8920 3440 8950
rect 3610 8920 3640 8950
rect 3810 8920 3840 8950
rect 4010 8920 4040 8950
rect 4210 8920 4240 8950
rect 4410 8920 4440 8950
rect 4610 8920 4640 8950
rect 4810 8920 4840 8950
rect 5010 8920 5040 8950
rect 5210 8920 5240 8950
rect 5410 8920 5440 8950
rect 5610 8920 5640 8950
rect 5810 8920 5840 8950
rect 6010 8920 6040 8950
rect 6210 8920 6240 8950
rect 6410 8920 6440 8950
rect -190 8805 -185 8835
rect -185 8805 -165 8835
rect -165 8805 -160 8835
rect 10 8805 40 8835
rect 210 8805 240 8835
rect 410 8805 440 8835
rect 610 8805 640 8835
rect 810 8805 840 8835
rect 1010 8805 1040 8835
rect 1210 8805 1240 8835
rect 1410 8805 1440 8835
rect 1610 8805 1640 8835
rect 1810 8805 1840 8835
rect 2010 8805 2040 8835
rect 2210 8805 2240 8835
rect 2410 8805 2440 8835
rect 2610 8805 2640 8835
rect 2810 8805 2840 8835
rect 3010 8805 3040 8835
rect 3210 8805 3240 8835
rect 3410 8805 3440 8835
rect 3610 8805 3640 8835
rect 3810 8805 3840 8835
rect 4010 8805 4040 8835
rect 4210 8805 4240 8835
rect 4410 8805 4440 8835
rect 4610 8805 4640 8835
rect 4810 8805 4840 8835
rect 5010 8805 5040 8835
rect 5210 8805 5240 8835
rect 5410 8805 5440 8835
rect 5610 8805 5640 8835
rect 5810 8805 5840 8835
rect 6010 8805 6040 8835
rect 6210 8805 6240 8835
rect 6410 8805 6440 8835
rect -190 8735 -185 8765
rect -185 8735 -165 8765
rect -165 8735 -160 8765
rect 10 8735 40 8765
rect 210 8735 240 8765
rect 410 8735 440 8765
rect 610 8735 640 8765
rect 810 8735 840 8765
rect 1010 8735 1040 8765
rect 1210 8735 1240 8765
rect 1410 8735 1440 8765
rect 1610 8735 1640 8765
rect 1810 8735 1840 8765
rect 2010 8735 2040 8765
rect 2210 8735 2240 8765
rect 2410 8735 2440 8765
rect 2610 8735 2640 8765
rect 2810 8735 2840 8765
rect 3010 8735 3040 8765
rect 3210 8735 3240 8765
rect 3410 8735 3440 8765
rect 3610 8735 3640 8765
rect 3810 8735 3840 8765
rect 4010 8735 4040 8765
rect 4210 8735 4240 8765
rect 4410 8735 4440 8765
rect 4610 8735 4640 8765
rect 4810 8735 4840 8765
rect 5010 8735 5040 8765
rect 5210 8735 5240 8765
rect 5410 8735 5440 8765
rect 5610 8735 5640 8765
rect 5810 8735 5840 8765
rect 6010 8735 6040 8765
rect 6210 8735 6240 8765
rect 6410 8735 6440 8765
rect -190 8620 -185 8650
rect -185 8620 -165 8650
rect -165 8620 -160 8650
rect 10 8620 40 8650
rect 210 8620 240 8650
rect 410 8620 440 8650
rect 610 8620 640 8650
rect 810 8620 840 8650
rect 1010 8620 1040 8650
rect 1210 8620 1240 8650
rect 1410 8620 1440 8650
rect 1610 8620 1640 8650
rect 1810 8620 1840 8650
rect 2010 8620 2040 8650
rect 2210 8620 2240 8650
rect 2410 8620 2440 8650
rect 2610 8620 2640 8650
rect 2810 8620 2840 8650
rect 3010 8620 3040 8650
rect 3210 8620 3240 8650
rect 3410 8620 3440 8650
rect 3610 8620 3640 8650
rect 3810 8620 3840 8650
rect 4010 8620 4040 8650
rect 4210 8620 4240 8650
rect 4410 8620 4440 8650
rect 4610 8620 4640 8650
rect 4810 8620 4840 8650
rect 5010 8620 5040 8650
rect 5210 8620 5240 8650
rect 5410 8620 5440 8650
rect 5610 8620 5640 8650
rect 5810 8620 5840 8650
rect 6010 8620 6040 8650
rect 6210 8620 6240 8650
rect 6410 8620 6440 8650
rect -190 8550 -185 8580
rect -185 8550 -165 8580
rect -165 8550 -160 8580
rect 10 8550 40 8580
rect 210 8550 240 8580
rect 410 8550 440 8580
rect 610 8550 640 8580
rect 810 8550 840 8580
rect 1010 8550 1040 8580
rect 1210 8550 1240 8580
rect 1410 8550 1440 8580
rect 1610 8550 1640 8580
rect 1810 8550 1840 8580
rect 2010 8550 2040 8580
rect 2210 8550 2240 8580
rect 2410 8550 2440 8580
rect 2610 8550 2640 8580
rect 2810 8550 2840 8580
rect 3010 8550 3040 8580
rect 3210 8550 3240 8580
rect 3410 8550 3440 8580
rect 3610 8550 3640 8580
rect 3810 8550 3840 8580
rect 4010 8550 4040 8580
rect 4210 8550 4240 8580
rect 4410 8550 4440 8580
rect 4610 8550 4640 8580
rect 4810 8550 4840 8580
rect 5010 8550 5040 8580
rect 5210 8550 5240 8580
rect 5410 8550 5440 8580
rect 5610 8550 5640 8580
rect 5810 8550 5840 8580
rect 6010 8550 6040 8580
rect 6210 8550 6240 8580
rect 6410 8550 6440 8580
rect -190 8435 -185 8465
rect -185 8435 -165 8465
rect -165 8435 -160 8465
rect 10 8435 40 8465
rect 210 8435 240 8465
rect 410 8435 440 8465
rect 610 8435 640 8465
rect 810 8435 840 8465
rect 1010 8435 1040 8465
rect 1210 8435 1240 8465
rect 1410 8435 1440 8465
rect 1610 8435 1640 8465
rect 1810 8435 1840 8465
rect 2010 8435 2040 8465
rect 2210 8435 2240 8465
rect 2410 8435 2440 8465
rect 2610 8435 2640 8465
rect 2810 8435 2840 8465
rect 3010 8435 3040 8465
rect 3210 8435 3240 8465
rect 3410 8435 3440 8465
rect 3610 8435 3640 8465
rect 3810 8435 3840 8465
rect 4010 8435 4040 8465
rect 4210 8435 4240 8465
rect 4410 8435 4440 8465
rect 4610 8435 4640 8465
rect 4810 8435 4840 8465
rect 5010 8435 5040 8465
rect 5210 8435 5240 8465
rect 5410 8435 5440 8465
rect 5610 8435 5640 8465
rect 5810 8435 5840 8465
rect 6010 8435 6040 8465
rect 6210 8435 6240 8465
rect 6410 8435 6440 8465
rect -190 8365 -185 8395
rect -185 8365 -165 8395
rect -165 8365 -160 8395
rect 10 8365 40 8395
rect 210 8365 240 8395
rect 410 8365 440 8395
rect 610 8365 640 8395
rect 810 8365 840 8395
rect 1010 8365 1040 8395
rect 1210 8365 1240 8395
rect 1410 8365 1440 8395
rect 1610 8365 1640 8395
rect 1810 8365 1840 8395
rect 2010 8365 2040 8395
rect 2210 8365 2240 8395
rect 2410 8365 2440 8395
rect 2610 8365 2640 8395
rect 2810 8365 2840 8395
rect 3010 8365 3040 8395
rect 3210 8365 3240 8395
rect 3410 8365 3440 8395
rect 3610 8365 3640 8395
rect 3810 8365 3840 8395
rect 4010 8365 4040 8395
rect 4210 8365 4240 8395
rect 4410 8365 4440 8395
rect 4610 8365 4640 8395
rect 4810 8365 4840 8395
rect 5010 8365 5040 8395
rect 5210 8365 5240 8395
rect 5410 8365 5440 8395
rect 5610 8365 5640 8395
rect 5810 8365 5840 8395
rect 6010 8365 6040 8395
rect 6210 8365 6240 8395
rect 6410 8365 6440 8395
rect -190 8250 -185 8280
rect -185 8250 -165 8280
rect -165 8250 -160 8280
rect 10 8250 40 8280
rect 210 8250 240 8280
rect 410 8250 440 8280
rect 610 8250 640 8280
rect 810 8250 840 8280
rect 1010 8250 1040 8280
rect 1210 8250 1240 8280
rect 1410 8250 1440 8280
rect 1610 8250 1640 8280
rect 1810 8250 1840 8280
rect 2010 8250 2040 8280
rect 2210 8250 2240 8280
rect 2410 8250 2440 8280
rect 2610 8250 2640 8280
rect 2810 8250 2840 8280
rect 3010 8250 3040 8280
rect 3210 8250 3240 8280
rect 3410 8250 3440 8280
rect 3610 8250 3640 8280
rect 3810 8250 3840 8280
rect 4010 8250 4040 8280
rect 4210 8250 4240 8280
rect 4410 8250 4440 8280
rect 4610 8250 4640 8280
rect 4810 8250 4840 8280
rect 5010 8250 5040 8280
rect 5210 8250 5240 8280
rect 5410 8250 5440 8280
rect 5610 8250 5640 8280
rect 5810 8250 5840 8280
rect 6010 8250 6040 8280
rect 6210 8250 6240 8280
rect 6410 8250 6440 8280
rect -190 8180 -185 8210
rect -185 8180 -165 8210
rect -165 8180 -160 8210
rect 10 8180 40 8210
rect 210 8180 240 8210
rect 410 8180 440 8210
rect 610 8180 640 8210
rect 810 8180 840 8210
rect 1010 8180 1040 8210
rect 1210 8180 1240 8210
rect 1410 8180 1440 8210
rect 1610 8180 1640 8210
rect 1810 8180 1840 8210
rect 2010 8180 2040 8210
rect 2210 8180 2240 8210
rect 2410 8180 2440 8210
rect 2610 8180 2640 8210
rect 2810 8180 2840 8210
rect 3010 8180 3040 8210
rect 3210 8180 3240 8210
rect 3410 8180 3440 8210
rect 3610 8180 3640 8210
rect 3810 8180 3840 8210
rect 4010 8180 4040 8210
rect 4210 8180 4240 8210
rect 4410 8180 4440 8210
rect 4610 8180 4640 8210
rect 4810 8180 4840 8210
rect 5010 8180 5040 8210
rect 5210 8180 5240 8210
rect 5410 8180 5440 8210
rect 5610 8180 5640 8210
rect 5810 8180 5840 8210
rect 6010 8180 6040 8210
rect 6210 8180 6240 8210
rect 6410 8180 6440 8210
rect -190 8065 -185 8095
rect -185 8065 -165 8095
rect -165 8065 -160 8095
rect 10 8065 40 8095
rect 210 8065 240 8095
rect 410 8065 440 8095
rect 610 8065 640 8095
rect 810 8065 840 8095
rect 1010 8065 1040 8095
rect 1210 8065 1240 8095
rect 1410 8065 1440 8095
rect 1610 8065 1640 8095
rect 1810 8065 1840 8095
rect 2010 8065 2040 8095
rect 2210 8065 2240 8095
rect 2410 8065 2440 8095
rect 2610 8065 2640 8095
rect 2810 8065 2840 8095
rect 3010 8065 3040 8095
rect 3210 8065 3240 8095
rect 3410 8065 3440 8095
rect 3610 8065 3640 8095
rect 3810 8065 3840 8095
rect 4010 8065 4040 8095
rect 4210 8065 4240 8095
rect 4410 8065 4440 8095
rect 4610 8065 4640 8095
rect 4810 8065 4840 8095
rect 5010 8065 5040 8095
rect 5210 8065 5240 8095
rect 5410 8065 5440 8095
rect 5610 8065 5640 8095
rect 5810 8065 5840 8095
rect 6010 8065 6040 8095
rect 6210 8065 6240 8095
rect 6410 8065 6440 8095
rect -190 7995 -185 8025
rect -185 7995 -165 8025
rect -165 7995 -160 8025
rect 10 7995 40 8025
rect 210 7995 240 8025
rect 410 7995 440 8025
rect 610 7995 640 8025
rect 810 7995 840 8025
rect 1010 7995 1040 8025
rect 1210 7995 1240 8025
rect 1410 7995 1440 8025
rect 1610 7995 1640 8025
rect 1810 7995 1840 8025
rect 2010 7995 2040 8025
rect 2210 7995 2240 8025
rect 2410 7995 2440 8025
rect 2610 7995 2640 8025
rect 2810 7995 2840 8025
rect 3010 7995 3040 8025
rect 3210 7995 3240 8025
rect 3410 7995 3440 8025
rect 3610 7995 3640 8025
rect 3810 7995 3840 8025
rect 4010 7995 4040 8025
rect 4210 7995 4240 8025
rect 4410 7995 4440 8025
rect 4610 7995 4640 8025
rect 4810 7995 4840 8025
rect 5010 7995 5040 8025
rect 5210 7995 5240 8025
rect 5410 7995 5440 8025
rect 5610 7995 5640 8025
rect 5810 7995 5840 8025
rect 6010 7995 6040 8025
rect 6210 7995 6240 8025
rect 6410 7995 6440 8025
rect -190 7880 -185 7910
rect -185 7880 -165 7910
rect -165 7880 -160 7910
rect 10 7880 40 7910
rect 210 7880 240 7910
rect 410 7880 440 7910
rect 610 7880 640 7910
rect 810 7880 840 7910
rect 1010 7880 1040 7910
rect 1210 7880 1240 7910
rect 1410 7880 1440 7910
rect 1610 7880 1640 7910
rect 1810 7880 1840 7910
rect 2010 7880 2040 7910
rect 2210 7880 2240 7910
rect 2410 7880 2440 7910
rect 2610 7880 2640 7910
rect 2810 7880 2840 7910
rect 3010 7880 3040 7910
rect 3210 7880 3240 7910
rect 3410 7880 3440 7910
rect 3610 7880 3640 7910
rect 3810 7880 3840 7910
rect 4010 7880 4040 7910
rect 4210 7880 4240 7910
rect 4410 7880 4440 7910
rect 4610 7880 4640 7910
rect 4810 7880 4840 7910
rect 5010 7880 5040 7910
rect 5210 7880 5240 7910
rect 5410 7880 5440 7910
rect 5610 7880 5640 7910
rect 5810 7880 5840 7910
rect 6010 7880 6040 7910
rect 6210 7880 6240 7910
rect 6410 7880 6440 7910
rect -190 7810 -185 7840
rect -185 7810 -165 7840
rect -165 7810 -160 7840
rect 10 7810 40 7840
rect 210 7810 240 7840
rect 410 7810 440 7840
rect 610 7810 640 7840
rect 810 7810 840 7840
rect 1010 7810 1040 7840
rect 1210 7810 1240 7840
rect 1410 7810 1440 7840
rect 1610 7810 1640 7840
rect 1810 7810 1840 7840
rect 2010 7810 2040 7840
rect 2210 7810 2240 7840
rect 2410 7810 2440 7840
rect 2610 7810 2640 7840
rect 2810 7810 2840 7840
rect 3010 7810 3040 7840
rect 3210 7810 3240 7840
rect 3410 7810 3440 7840
rect 3610 7810 3640 7840
rect 3810 7810 3840 7840
rect 4010 7810 4040 7840
rect 4210 7810 4240 7840
rect 4410 7810 4440 7840
rect 4610 7810 4640 7840
rect 4810 7810 4840 7840
rect 5010 7810 5040 7840
rect 5210 7810 5240 7840
rect 5410 7810 5440 7840
rect 5610 7810 5640 7840
rect 5810 7810 5840 7840
rect 6010 7810 6040 7840
rect 6210 7810 6240 7840
rect 6410 7810 6440 7840
rect -190 7695 -185 7725
rect -185 7695 -165 7725
rect -165 7695 -160 7725
rect 10 7695 40 7725
rect 210 7695 240 7725
rect 410 7695 440 7725
rect 610 7695 640 7725
rect 810 7695 840 7725
rect 1010 7695 1040 7725
rect 1210 7695 1240 7725
rect 1410 7695 1440 7725
rect 1610 7695 1640 7725
rect 1810 7695 1840 7725
rect 2010 7695 2040 7725
rect 2210 7695 2240 7725
rect 2410 7695 2440 7725
rect 2610 7695 2640 7725
rect 2810 7695 2840 7725
rect 3010 7695 3040 7725
rect 3210 7695 3240 7725
rect 3410 7695 3440 7725
rect 3610 7695 3640 7725
rect 3810 7695 3840 7725
rect 4010 7695 4040 7725
rect 4210 7695 4240 7725
rect 4410 7695 4440 7725
rect 4610 7695 4640 7725
rect 4810 7695 4840 7725
rect 5010 7695 5040 7725
rect 5210 7695 5240 7725
rect 5410 7695 5440 7725
rect 5610 7695 5640 7725
rect 5810 7695 5840 7725
rect 6010 7695 6040 7725
rect 6210 7695 6240 7725
rect 6410 7695 6440 7725
rect -190 7625 -185 7655
rect -185 7625 -165 7655
rect -165 7625 -160 7655
rect 10 7625 40 7655
rect 210 7625 240 7655
rect 410 7625 440 7655
rect 610 7625 640 7655
rect 810 7625 840 7655
rect 1010 7625 1040 7655
rect 1210 7625 1240 7655
rect 1410 7625 1440 7655
rect 1610 7625 1640 7655
rect 1810 7625 1840 7655
rect 2010 7625 2040 7655
rect 2210 7625 2240 7655
rect 2410 7625 2440 7655
rect 2610 7625 2640 7655
rect 2810 7625 2840 7655
rect 3010 7625 3040 7655
rect 3210 7625 3240 7655
rect 3410 7625 3440 7655
rect 3610 7625 3640 7655
rect 3810 7625 3840 7655
rect 4010 7625 4040 7655
rect 4210 7625 4240 7655
rect 4410 7625 4440 7655
rect 4610 7625 4640 7655
rect 4810 7625 4840 7655
rect 5010 7625 5040 7655
rect 5210 7625 5240 7655
rect 5410 7625 5440 7655
rect 5610 7625 5640 7655
rect 5810 7625 5840 7655
rect 6010 7625 6040 7655
rect 6210 7625 6240 7655
rect 6410 7625 6440 7655
rect -190 7510 -185 7540
rect -185 7510 -165 7540
rect -165 7510 -160 7540
rect 10 7510 40 7540
rect 210 7510 240 7540
rect 410 7510 440 7540
rect 610 7510 640 7540
rect 810 7510 840 7540
rect 1010 7510 1040 7540
rect 1210 7510 1240 7540
rect 1410 7510 1440 7540
rect 1610 7510 1640 7540
rect 1810 7510 1840 7540
rect 2010 7510 2040 7540
rect 2210 7510 2240 7540
rect 2410 7510 2440 7540
rect 2610 7510 2640 7540
rect 2810 7510 2840 7540
rect 3010 7510 3040 7540
rect 3210 7510 3240 7540
rect 3410 7510 3440 7540
rect 3610 7510 3640 7540
rect 3810 7510 3840 7540
rect 4010 7510 4040 7540
rect 4210 7510 4240 7540
rect 4410 7510 4440 7540
rect 4610 7510 4640 7540
rect 4810 7510 4840 7540
rect 5010 7510 5040 7540
rect 5210 7510 5240 7540
rect 5410 7510 5440 7540
rect 5610 7510 5640 7540
rect 5810 7510 5840 7540
rect 6010 7510 6040 7540
rect 6210 7510 6240 7540
rect 6410 7510 6440 7540
rect -190 7440 -185 7470
rect -185 7440 -165 7470
rect -165 7440 -160 7470
rect 10 7440 40 7470
rect 210 7440 240 7470
rect 410 7440 440 7470
rect 610 7440 640 7470
rect 810 7440 840 7470
rect 1010 7440 1040 7470
rect 1210 7440 1240 7470
rect 1410 7440 1440 7470
rect 1610 7440 1640 7470
rect 1810 7440 1840 7470
rect 2010 7440 2040 7470
rect 2210 7440 2240 7470
rect 2410 7440 2440 7470
rect 2610 7440 2640 7470
rect 2810 7440 2840 7470
rect 3010 7440 3040 7470
rect 3210 7440 3240 7470
rect 3410 7440 3440 7470
rect 3610 7440 3640 7470
rect 3810 7440 3840 7470
rect 4010 7440 4040 7470
rect 4210 7440 4240 7470
rect 4410 7440 4440 7470
rect 4610 7440 4640 7470
rect 4810 7440 4840 7470
rect 5010 7440 5040 7470
rect 5210 7440 5240 7470
rect 5410 7440 5440 7470
rect 5610 7440 5640 7470
rect 5810 7440 5840 7470
rect 6010 7440 6040 7470
rect 6210 7440 6240 7470
rect 6410 7440 6440 7470
rect -190 7325 -185 7355
rect -185 7325 -165 7355
rect -165 7325 -160 7355
rect 10 7325 40 7355
rect 210 7325 240 7355
rect 410 7325 440 7355
rect 610 7325 640 7355
rect 810 7325 840 7355
rect 1010 7325 1040 7355
rect 1210 7325 1240 7355
rect 1410 7325 1440 7355
rect 1610 7325 1640 7355
rect 1810 7325 1840 7355
rect 2010 7325 2040 7355
rect 2210 7325 2240 7355
rect 2410 7325 2440 7355
rect 2610 7325 2640 7355
rect 2810 7325 2840 7355
rect 3010 7325 3040 7355
rect 3210 7325 3240 7355
rect 3410 7325 3440 7355
rect 3610 7325 3640 7355
rect 3810 7325 3840 7355
rect 4010 7325 4040 7355
rect 4210 7325 4240 7355
rect 4410 7325 4440 7355
rect 4610 7325 4640 7355
rect 4810 7325 4840 7355
rect 5010 7325 5040 7355
rect 5210 7325 5240 7355
rect 5410 7325 5440 7355
rect 5610 7325 5640 7355
rect 5810 7325 5840 7355
rect 6010 7325 6040 7355
rect 6210 7325 6240 7355
rect 6410 7325 6440 7355
rect -190 7255 -185 7285
rect -185 7255 -165 7285
rect -165 7255 -160 7285
rect 10 7255 40 7285
rect 210 7255 240 7285
rect 410 7255 440 7285
rect 610 7255 640 7285
rect 810 7255 840 7285
rect 1010 7255 1040 7285
rect 1210 7255 1240 7285
rect 1410 7255 1440 7285
rect 1610 7255 1640 7285
rect 1810 7255 1840 7285
rect 2010 7255 2040 7285
rect 2210 7255 2240 7285
rect 2410 7255 2440 7285
rect 2610 7255 2640 7285
rect 2810 7255 2840 7285
rect 3010 7255 3040 7285
rect 3210 7255 3240 7285
rect 3410 7255 3440 7285
rect 3610 7255 3640 7285
rect 3810 7255 3840 7285
rect 4010 7255 4040 7285
rect 4210 7255 4240 7285
rect 4410 7255 4440 7285
rect 4610 7255 4640 7285
rect 4810 7255 4840 7285
rect 5010 7255 5040 7285
rect 5210 7255 5240 7285
rect 5410 7255 5440 7285
rect 5610 7255 5640 7285
rect 5810 7255 5840 7285
rect 6010 7255 6040 7285
rect 6210 7255 6240 7285
rect 6410 7255 6440 7285
rect -190 7140 -185 7170
rect -185 7140 -165 7170
rect -165 7140 -160 7170
rect 10 7140 40 7170
rect 210 7140 240 7170
rect 410 7140 440 7170
rect 610 7140 640 7170
rect 810 7140 840 7170
rect 1010 7140 1040 7170
rect 1210 7140 1240 7170
rect 1410 7140 1440 7170
rect 1610 7140 1640 7170
rect 1810 7140 1840 7170
rect 2010 7140 2040 7170
rect 2210 7140 2240 7170
rect 2410 7140 2440 7170
rect 2610 7140 2640 7170
rect 2810 7140 2840 7170
rect 3010 7140 3040 7170
rect 3210 7140 3240 7170
rect 3410 7140 3440 7170
rect 3610 7140 3640 7170
rect 3810 7140 3840 7170
rect 4010 7140 4040 7170
rect 4210 7140 4240 7170
rect 4410 7140 4440 7170
rect 4610 7140 4640 7170
rect 4810 7140 4840 7170
rect 5010 7140 5040 7170
rect 5210 7140 5240 7170
rect 5410 7140 5440 7170
rect 5610 7140 5640 7170
rect 5810 7140 5840 7170
rect 6010 7140 6040 7170
rect 6210 7140 6240 7170
rect 6410 7140 6440 7170
rect -190 7070 -185 7100
rect -185 7070 -165 7100
rect -165 7070 -160 7100
rect 10 7070 40 7100
rect 210 7070 240 7100
rect 410 7070 440 7100
rect 610 7070 640 7100
rect 810 7070 840 7100
rect 1010 7070 1040 7100
rect 1210 7070 1240 7100
rect 1410 7070 1440 7100
rect 1610 7070 1640 7100
rect 1810 7070 1840 7100
rect 2010 7070 2040 7100
rect 2210 7070 2240 7100
rect 2410 7070 2440 7100
rect 2610 7070 2640 7100
rect 2810 7070 2840 7100
rect 3010 7070 3040 7100
rect 3210 7070 3240 7100
rect 3410 7070 3440 7100
rect 3610 7070 3640 7100
rect 3810 7070 3840 7100
rect 4010 7070 4040 7100
rect 4210 7070 4240 7100
rect 4410 7070 4440 7100
rect 4610 7070 4640 7100
rect 4810 7070 4840 7100
rect 5010 7070 5040 7100
rect 5210 7070 5240 7100
rect 5410 7070 5440 7100
rect 5610 7070 5640 7100
rect 5810 7070 5840 7100
rect 6010 7070 6040 7100
rect 6210 7070 6240 7100
rect 6410 7070 6440 7100
rect -190 6955 -185 6985
rect -185 6955 -165 6985
rect -165 6955 -160 6985
rect 10 6955 40 6985
rect 210 6955 240 6985
rect 410 6955 440 6985
rect 610 6955 640 6985
rect 810 6955 840 6985
rect 1010 6955 1040 6985
rect 1210 6955 1240 6985
rect 1410 6955 1440 6985
rect 1610 6955 1640 6985
rect 1810 6955 1840 6985
rect 2010 6955 2040 6985
rect 2210 6955 2240 6985
rect 2410 6955 2440 6985
rect 2610 6955 2640 6985
rect 2810 6955 2840 6985
rect 3010 6955 3040 6985
rect 3210 6955 3240 6985
rect 3410 6955 3440 6985
rect 3610 6955 3640 6985
rect 3810 6955 3840 6985
rect 4010 6955 4040 6985
rect 4210 6955 4240 6985
rect 4410 6955 4440 6985
rect 4610 6955 4640 6985
rect 4810 6955 4840 6985
rect 5010 6955 5040 6985
rect 5210 6955 5240 6985
rect 5410 6955 5440 6985
rect 5610 6955 5640 6985
rect 5810 6955 5840 6985
rect 6010 6955 6040 6985
rect 6210 6955 6240 6985
rect 6410 6955 6440 6985
rect -190 6885 -185 6915
rect -185 6885 -165 6915
rect -165 6885 -160 6915
rect 10 6885 40 6915
rect 210 6885 240 6915
rect 410 6885 440 6915
rect 610 6885 640 6915
rect 810 6885 840 6915
rect 1010 6885 1040 6915
rect 1210 6885 1240 6915
rect 1410 6885 1440 6915
rect 1610 6885 1640 6915
rect 1810 6885 1840 6915
rect 2010 6885 2040 6915
rect 2210 6885 2240 6915
rect 2410 6885 2440 6915
rect 2610 6885 2640 6915
rect 2810 6885 2840 6915
rect 3010 6885 3040 6915
rect 3210 6885 3240 6915
rect 3410 6885 3440 6915
rect 3610 6885 3640 6915
rect 3810 6885 3840 6915
rect 4010 6885 4040 6915
rect 4210 6885 4240 6915
rect 4410 6885 4440 6915
rect 4610 6885 4640 6915
rect 4810 6885 4840 6915
rect 5010 6885 5040 6915
rect 5210 6885 5240 6915
rect 5410 6885 5440 6915
rect 5610 6885 5640 6915
rect 5810 6885 5840 6915
rect 6010 6885 6040 6915
rect 6210 6885 6240 6915
rect 6410 6885 6440 6915
rect -190 6770 -185 6800
rect -185 6770 -165 6800
rect -165 6770 -160 6800
rect 10 6770 40 6800
rect 210 6770 240 6800
rect 410 6770 440 6800
rect 610 6770 640 6800
rect 810 6770 840 6800
rect 1010 6770 1040 6800
rect 1210 6770 1240 6800
rect 1410 6770 1440 6800
rect 1610 6770 1640 6800
rect 1810 6770 1840 6800
rect 2010 6770 2040 6800
rect 2210 6770 2240 6800
rect 2410 6770 2440 6800
rect 2610 6770 2640 6800
rect 2810 6770 2840 6800
rect 3010 6770 3040 6800
rect 3210 6770 3240 6800
rect 3410 6770 3440 6800
rect 3610 6770 3640 6800
rect 3810 6770 3840 6800
rect 4010 6770 4040 6800
rect 4210 6770 4240 6800
rect 4410 6770 4440 6800
rect 4610 6770 4640 6800
rect 4810 6770 4840 6800
rect 5010 6770 5040 6800
rect 5210 6770 5240 6800
rect 5410 6770 5440 6800
rect 5610 6770 5640 6800
rect 5810 6770 5840 6800
rect 6010 6770 6040 6800
rect 6210 6770 6240 6800
rect 6410 6770 6440 6800
rect -190 6700 -185 6730
rect -185 6700 -165 6730
rect -165 6700 -160 6730
rect 10 6700 40 6730
rect 210 6700 240 6730
rect 410 6700 440 6730
rect 610 6700 640 6730
rect 810 6700 840 6730
rect 1010 6700 1040 6730
rect 1210 6700 1240 6730
rect 1410 6700 1440 6730
rect 1610 6700 1640 6730
rect 1810 6700 1840 6730
rect 2010 6700 2040 6730
rect 2210 6700 2240 6730
rect 2410 6700 2440 6730
rect 2610 6700 2640 6730
rect 2810 6700 2840 6730
rect 3010 6700 3040 6730
rect 3210 6700 3240 6730
rect 3410 6700 3440 6730
rect 3610 6700 3640 6730
rect 3810 6700 3840 6730
rect 4010 6700 4040 6730
rect 4210 6700 4240 6730
rect 4410 6700 4440 6730
rect 4610 6700 4640 6730
rect 4810 6700 4840 6730
rect 5010 6700 5040 6730
rect 5210 6700 5240 6730
rect 5410 6700 5440 6730
rect 5610 6700 5640 6730
rect 5810 6700 5840 6730
rect 6010 6700 6040 6730
rect 6210 6700 6240 6730
rect 6410 6700 6440 6730
rect -190 6585 -185 6615
rect -185 6585 -165 6615
rect -165 6585 -160 6615
rect 10 6585 40 6615
rect 210 6585 240 6615
rect 410 6585 440 6615
rect 610 6585 640 6615
rect 810 6585 840 6615
rect 1010 6585 1040 6615
rect 1210 6585 1240 6615
rect 1410 6585 1440 6615
rect 1610 6585 1640 6615
rect 1810 6585 1840 6615
rect 2010 6585 2040 6615
rect 2210 6585 2240 6615
rect 2410 6585 2440 6615
rect 2610 6585 2640 6615
rect 2810 6585 2840 6615
rect 3010 6585 3040 6615
rect 3210 6585 3240 6615
rect 3410 6585 3440 6615
rect 3610 6585 3640 6615
rect 3810 6585 3840 6615
rect 4010 6585 4040 6615
rect 4210 6585 4240 6615
rect 4410 6585 4440 6615
rect 4610 6585 4640 6615
rect 4810 6585 4840 6615
rect 5010 6585 5040 6615
rect 5210 6585 5240 6615
rect 5410 6585 5440 6615
rect 5610 6585 5640 6615
rect 5810 6585 5840 6615
rect 6010 6585 6040 6615
rect 6210 6585 6240 6615
rect 6410 6585 6440 6615
rect -190 6515 -185 6545
rect -185 6515 -165 6545
rect -165 6515 -160 6545
rect 10 6515 40 6545
rect 210 6515 240 6545
rect 410 6515 440 6545
rect 610 6515 640 6545
rect 810 6515 840 6545
rect 1010 6515 1040 6545
rect 1210 6515 1240 6545
rect 1410 6515 1440 6545
rect 1610 6515 1640 6545
rect 1810 6515 1840 6545
rect 2010 6515 2040 6545
rect 2210 6515 2240 6545
rect 2410 6515 2440 6545
rect 2610 6515 2640 6545
rect 2810 6515 2840 6545
rect 3010 6515 3040 6545
rect 3210 6515 3240 6545
rect 3410 6515 3440 6545
rect 3610 6515 3640 6545
rect 3810 6515 3840 6545
rect 4010 6515 4040 6545
rect 4210 6515 4240 6545
rect 4410 6515 4440 6545
rect 4610 6515 4640 6545
rect 4810 6515 4840 6545
rect 5010 6515 5040 6545
rect 5210 6515 5240 6545
rect 5410 6515 5440 6545
rect 5610 6515 5640 6545
rect 5810 6515 5840 6545
rect 6010 6515 6040 6545
rect 6210 6515 6240 6545
rect 6410 6515 6440 6545
rect -190 6400 -185 6430
rect -185 6400 -165 6430
rect -165 6400 -160 6430
rect 10 6400 40 6430
rect 210 6400 240 6430
rect 410 6400 440 6430
rect 610 6400 640 6430
rect 810 6400 840 6430
rect 1010 6400 1040 6430
rect 1210 6400 1240 6430
rect 1410 6400 1440 6430
rect 1610 6400 1640 6430
rect 1810 6400 1840 6430
rect 2010 6400 2040 6430
rect 2210 6400 2240 6430
rect 2410 6400 2440 6430
rect 2610 6400 2640 6430
rect 2810 6400 2840 6430
rect 3010 6400 3040 6430
rect 3210 6400 3240 6430
rect 3410 6400 3440 6430
rect 3610 6400 3640 6430
rect 3810 6400 3840 6430
rect 4010 6400 4040 6430
rect 4210 6400 4240 6430
rect 4410 6400 4440 6430
rect 4610 6400 4640 6430
rect 4810 6400 4840 6430
rect 5010 6400 5040 6430
rect 5210 6400 5240 6430
rect 5410 6400 5440 6430
rect 5610 6400 5640 6430
rect 5810 6400 5840 6430
rect 6010 6400 6040 6430
rect 6210 6400 6240 6430
rect 6410 6400 6440 6430
rect -190 6330 -185 6360
rect -185 6330 -165 6360
rect -165 6330 -160 6360
rect 10 6330 40 6360
rect 210 6330 240 6360
rect 410 6330 440 6360
rect 610 6330 640 6360
rect 810 6330 840 6360
rect 1010 6330 1040 6360
rect 1210 6330 1240 6360
rect 1410 6330 1440 6360
rect 1610 6330 1640 6360
rect 1810 6330 1840 6360
rect 2010 6330 2040 6360
rect 2210 6330 2240 6360
rect 2410 6330 2440 6360
rect 2610 6330 2640 6360
rect 2810 6330 2840 6360
rect 3010 6330 3040 6360
rect 3210 6330 3240 6360
rect 3410 6330 3440 6360
rect 3610 6330 3640 6360
rect 3810 6330 3840 6360
rect 4010 6330 4040 6360
rect 4210 6330 4240 6360
rect 4410 6330 4440 6360
rect 4610 6330 4640 6360
rect 4810 6330 4840 6360
rect 5010 6330 5040 6360
rect 5210 6330 5240 6360
rect 5410 6330 5440 6360
rect 5610 6330 5640 6360
rect 5810 6330 5840 6360
rect 6010 6330 6040 6360
rect 6210 6330 6240 6360
rect 6410 6330 6440 6360
rect -190 6215 -185 6245
rect -185 6215 -165 6245
rect -165 6215 -160 6245
rect 10 6215 40 6245
rect 210 6215 240 6245
rect 410 6215 440 6245
rect 610 6215 640 6245
rect 810 6215 840 6245
rect 1010 6215 1040 6245
rect 1210 6215 1240 6245
rect 1410 6215 1440 6245
rect 1610 6215 1640 6245
rect 1810 6215 1840 6245
rect 2010 6215 2040 6245
rect 2210 6215 2240 6245
rect 2410 6215 2440 6245
rect 2610 6215 2640 6245
rect 2810 6215 2840 6245
rect 3010 6215 3040 6245
rect 3210 6215 3240 6245
rect 3410 6215 3440 6245
rect 3610 6215 3640 6245
rect 3810 6215 3840 6245
rect 4010 6215 4040 6245
rect 4210 6215 4240 6245
rect 4410 6215 4440 6245
rect 4610 6215 4640 6245
rect 4810 6215 4840 6245
rect 5010 6215 5040 6245
rect 5210 6215 5240 6245
rect 5410 6215 5440 6245
rect 5610 6215 5640 6245
rect 5810 6215 5840 6245
rect 6010 6215 6040 6245
rect 6210 6215 6240 6245
rect 6410 6215 6440 6245
rect -190 6145 -185 6175
rect -185 6145 -165 6175
rect -165 6145 -160 6175
rect 10 6145 40 6175
rect 210 6145 240 6175
rect 410 6145 440 6175
rect 610 6145 640 6175
rect 810 6145 840 6175
rect 1010 6145 1040 6175
rect 1210 6145 1240 6175
rect 1410 6145 1440 6175
rect 1610 6145 1640 6175
rect 1810 6145 1840 6175
rect 2010 6145 2040 6175
rect 2210 6145 2240 6175
rect 2410 6145 2440 6175
rect 2610 6145 2640 6175
rect 2810 6145 2840 6175
rect 3010 6145 3040 6175
rect 3210 6145 3240 6175
rect 3410 6145 3440 6175
rect 3610 6145 3640 6175
rect 3810 6145 3840 6175
rect 4010 6145 4040 6175
rect 4210 6145 4240 6175
rect 4410 6145 4440 6175
rect 4610 6145 4640 6175
rect 4810 6145 4840 6175
rect 5010 6145 5040 6175
rect 5210 6145 5240 6175
rect 5410 6145 5440 6175
rect 5610 6145 5640 6175
rect 5810 6145 5840 6175
rect 6010 6145 6040 6175
rect 6210 6145 6240 6175
rect 6410 6145 6440 6175
rect -190 6030 -185 6060
rect -185 6030 -165 6060
rect -165 6030 -160 6060
rect 10 6030 40 6060
rect 210 6030 240 6060
rect 410 6030 440 6060
rect 610 6030 640 6060
rect 810 6030 840 6060
rect 1010 6030 1040 6060
rect 1210 6030 1240 6060
rect 1410 6030 1440 6060
rect 1610 6030 1640 6060
rect 1810 6030 1840 6060
rect 2010 6030 2040 6060
rect 2210 6030 2240 6060
rect 2410 6030 2440 6060
rect 2610 6030 2640 6060
rect 2810 6030 2840 6060
rect 3010 6030 3040 6060
rect 3210 6030 3240 6060
rect 3410 6030 3440 6060
rect 3610 6030 3640 6060
rect 3810 6030 3840 6060
rect 4010 6030 4040 6060
rect 4210 6030 4240 6060
rect 4410 6030 4440 6060
rect 4610 6030 4640 6060
rect 4810 6030 4840 6060
rect 5010 6030 5040 6060
rect 5210 6030 5240 6060
rect 5410 6030 5440 6060
rect 5610 6030 5640 6060
rect 5810 6030 5840 6060
rect 6010 6030 6040 6060
rect 6210 6030 6240 6060
rect 6410 6030 6440 6060
rect -190 5960 -185 5990
rect -185 5960 -165 5990
rect -165 5960 -160 5990
rect 10 5960 40 5990
rect 210 5960 240 5990
rect 410 5960 440 5990
rect 610 5960 640 5990
rect 810 5960 840 5990
rect 1010 5960 1040 5990
rect 1210 5960 1240 5990
rect 1410 5960 1440 5990
rect 1610 5960 1640 5990
rect 1810 5960 1840 5990
rect 2010 5960 2040 5990
rect 2210 5960 2240 5990
rect 2410 5960 2440 5990
rect 2610 5960 2640 5990
rect 2810 5960 2840 5990
rect 3010 5960 3040 5990
rect 3210 5960 3240 5990
rect 3410 5960 3440 5990
rect 3610 5960 3640 5990
rect 3810 5960 3840 5990
rect 4010 5960 4040 5990
rect 4210 5960 4240 5990
rect 4410 5960 4440 5990
rect 4610 5960 4640 5990
rect 4810 5960 4840 5990
rect 5010 5960 5040 5990
rect 5210 5960 5240 5990
rect 5410 5960 5440 5990
rect 5610 5960 5640 5990
rect 5810 5960 5840 5990
rect 6010 5960 6040 5990
rect 6210 5960 6240 5990
rect 6410 5960 6440 5990
rect -190 5845 -185 5875
rect -185 5845 -165 5875
rect -165 5845 -160 5875
rect 10 5845 40 5875
rect 210 5845 240 5875
rect 410 5845 440 5875
rect 610 5845 640 5875
rect 810 5845 840 5875
rect 1010 5845 1040 5875
rect 1210 5845 1240 5875
rect 1410 5845 1440 5875
rect 1610 5845 1640 5875
rect 1810 5845 1840 5875
rect 2010 5845 2040 5875
rect 2210 5845 2240 5875
rect 2410 5845 2440 5875
rect 2610 5845 2640 5875
rect 2810 5845 2840 5875
rect 3010 5845 3040 5875
rect 3210 5845 3240 5875
rect 3410 5845 3440 5875
rect 3610 5845 3640 5875
rect 3810 5845 3840 5875
rect 4010 5845 4040 5875
rect 4210 5845 4240 5875
rect 4410 5845 4440 5875
rect 4610 5845 4640 5875
rect 4810 5845 4840 5875
rect 5010 5845 5040 5875
rect 5210 5845 5240 5875
rect 5410 5845 5440 5875
rect 5610 5845 5640 5875
rect 5810 5845 5840 5875
rect 6010 5845 6040 5875
rect 6210 5845 6240 5875
rect 6410 5845 6440 5875
rect -190 5775 -185 5805
rect -185 5775 -165 5805
rect -165 5775 -160 5805
rect 10 5775 40 5805
rect 210 5775 240 5805
rect 410 5775 440 5805
rect 610 5775 640 5805
rect 810 5775 840 5805
rect 1010 5775 1040 5805
rect 1210 5775 1240 5805
rect 1410 5775 1440 5805
rect 1610 5775 1640 5805
rect 1810 5775 1840 5805
rect 2010 5775 2040 5805
rect 2210 5775 2240 5805
rect 2410 5775 2440 5805
rect 2610 5775 2640 5805
rect 2810 5775 2840 5805
rect 3010 5775 3040 5805
rect 3210 5775 3240 5805
rect 3410 5775 3440 5805
rect 3610 5775 3640 5805
rect 3810 5775 3840 5805
rect 4010 5775 4040 5805
rect 4210 5775 4240 5805
rect 4410 5775 4440 5805
rect 4610 5775 4640 5805
rect 4810 5775 4840 5805
rect 5010 5775 5040 5805
rect 5210 5775 5240 5805
rect 5410 5775 5440 5805
rect 5610 5775 5640 5805
rect 5810 5775 5840 5805
rect 6010 5775 6040 5805
rect 6210 5775 6240 5805
rect 6410 5775 6440 5805
rect -190 5660 -185 5690
rect -185 5660 -165 5690
rect -165 5660 -160 5690
rect 10 5660 40 5690
rect 210 5660 240 5690
rect 410 5660 440 5690
rect 610 5660 640 5690
rect 810 5660 840 5690
rect 1010 5660 1040 5690
rect 1210 5660 1240 5690
rect 1410 5660 1440 5690
rect 1610 5660 1640 5690
rect 1810 5660 1840 5690
rect 2010 5660 2040 5690
rect 2210 5660 2240 5690
rect 2410 5660 2440 5690
rect 2610 5660 2640 5690
rect 2810 5660 2840 5690
rect 3010 5660 3040 5690
rect 3210 5660 3240 5690
rect 3410 5660 3440 5690
rect 3610 5660 3640 5690
rect 3810 5660 3840 5690
rect 4010 5660 4040 5690
rect 4210 5660 4240 5690
rect 4410 5660 4440 5690
rect 4610 5660 4640 5690
rect 4810 5660 4840 5690
rect 5010 5660 5040 5690
rect 5210 5660 5240 5690
rect 5410 5660 5440 5690
rect 5610 5660 5640 5690
rect 5810 5660 5840 5690
rect 6010 5660 6040 5690
rect 6210 5660 6240 5690
rect 6410 5660 6440 5690
rect -190 5590 -185 5620
rect -185 5590 -165 5620
rect -165 5590 -160 5620
rect 10 5590 40 5620
rect 210 5590 240 5620
rect 410 5590 440 5620
rect 610 5590 640 5620
rect 810 5590 840 5620
rect 1010 5590 1040 5620
rect 1210 5590 1240 5620
rect 1410 5590 1440 5620
rect 1610 5590 1640 5620
rect 1810 5590 1840 5620
rect 2010 5590 2040 5620
rect 2210 5590 2240 5620
rect 2410 5590 2440 5620
rect 2610 5590 2640 5620
rect 2810 5590 2840 5620
rect 3010 5590 3040 5620
rect 3210 5590 3240 5620
rect 3410 5590 3440 5620
rect 3610 5590 3640 5620
rect 3810 5590 3840 5620
rect 4010 5590 4040 5620
rect 4210 5590 4240 5620
rect 4410 5590 4440 5620
rect 4610 5590 4640 5620
rect 4810 5590 4840 5620
rect 5010 5590 5040 5620
rect 5210 5590 5240 5620
rect 5410 5590 5440 5620
rect 5610 5590 5640 5620
rect 5810 5590 5840 5620
rect 6010 5590 6040 5620
rect 6210 5590 6240 5620
rect 6410 5590 6440 5620
rect -190 5475 -185 5505
rect -185 5475 -165 5505
rect -165 5475 -160 5505
rect 10 5475 40 5505
rect 210 5475 240 5505
rect 410 5475 440 5505
rect 610 5475 640 5505
rect 810 5475 840 5505
rect 1010 5475 1040 5505
rect 1210 5475 1240 5505
rect 1410 5475 1440 5505
rect 1610 5475 1640 5505
rect 1810 5475 1840 5505
rect 2010 5475 2040 5505
rect 2210 5475 2240 5505
rect 2410 5475 2440 5505
rect 2610 5475 2640 5505
rect 2810 5475 2840 5505
rect 3010 5475 3040 5505
rect 3210 5475 3240 5505
rect 3410 5475 3440 5505
rect 3610 5475 3640 5505
rect 3810 5475 3840 5505
rect 4010 5475 4040 5505
rect 4210 5475 4240 5505
rect 4410 5475 4440 5505
rect 4610 5475 4640 5505
rect 4810 5475 4840 5505
rect 5010 5475 5040 5505
rect 5210 5475 5240 5505
rect 5410 5475 5440 5505
rect 5610 5475 5640 5505
rect 5810 5475 5840 5505
rect 6010 5475 6040 5505
rect 6210 5475 6240 5505
rect 6410 5475 6440 5505
rect -190 5405 -185 5435
rect -185 5405 -165 5435
rect -165 5405 -160 5435
rect 10 5405 40 5435
rect 210 5405 240 5435
rect 410 5405 440 5435
rect 610 5405 640 5435
rect 810 5405 840 5435
rect 1010 5405 1040 5435
rect 1210 5405 1240 5435
rect 1410 5405 1440 5435
rect 1610 5405 1640 5435
rect 1810 5405 1840 5435
rect 2010 5405 2040 5435
rect 2210 5405 2240 5435
rect 2410 5405 2440 5435
rect 2610 5405 2640 5435
rect 2810 5405 2840 5435
rect 3010 5405 3040 5435
rect 3210 5405 3240 5435
rect 3410 5405 3440 5435
rect 3610 5405 3640 5435
rect 3810 5405 3840 5435
rect 4010 5405 4040 5435
rect 4210 5405 4240 5435
rect 4410 5405 4440 5435
rect 4610 5405 4640 5435
rect 4810 5405 4840 5435
rect 5010 5405 5040 5435
rect 5210 5405 5240 5435
rect 5410 5405 5440 5435
rect 5610 5405 5640 5435
rect 5810 5405 5840 5435
rect 6010 5405 6040 5435
rect 6210 5405 6240 5435
rect 6410 5405 6440 5435
rect -190 5290 -185 5320
rect -185 5290 -165 5320
rect -165 5290 -160 5320
rect 10 5290 40 5320
rect 210 5290 240 5320
rect 410 5290 440 5320
rect 610 5290 640 5320
rect 810 5290 840 5320
rect 1010 5290 1040 5320
rect 1210 5290 1240 5320
rect 1410 5290 1440 5320
rect 1610 5290 1640 5320
rect 1810 5290 1840 5320
rect 2010 5290 2040 5320
rect 2210 5290 2240 5320
rect 2410 5290 2440 5320
rect 2610 5290 2640 5320
rect 2810 5290 2840 5320
rect 3010 5290 3040 5320
rect 3210 5290 3240 5320
rect 3410 5290 3440 5320
rect 3610 5290 3640 5320
rect 3810 5290 3840 5320
rect 4010 5290 4040 5320
rect 4210 5290 4240 5320
rect 4410 5290 4440 5320
rect 4610 5290 4640 5320
rect 4810 5290 4840 5320
rect 5010 5290 5040 5320
rect 5210 5290 5240 5320
rect 5410 5290 5440 5320
rect 5610 5290 5640 5320
rect 5810 5290 5840 5320
rect 6010 5290 6040 5320
rect 6210 5290 6240 5320
rect 6410 5290 6440 5320
rect -190 5220 -185 5250
rect -185 5220 -165 5250
rect -165 5220 -160 5250
rect 10 5220 40 5250
rect 210 5220 240 5250
rect 410 5220 440 5250
rect 610 5220 640 5250
rect 810 5220 840 5250
rect 1010 5220 1040 5250
rect 1210 5220 1240 5250
rect 1410 5220 1440 5250
rect 1610 5220 1640 5250
rect 1810 5220 1840 5250
rect 2010 5220 2040 5250
rect 2210 5220 2240 5250
rect 2410 5220 2440 5250
rect 2610 5220 2640 5250
rect 2810 5220 2840 5250
rect 3010 5220 3040 5250
rect 3210 5220 3240 5250
rect 3410 5220 3440 5250
rect 3610 5220 3640 5250
rect 3810 5220 3840 5250
rect 4010 5220 4040 5250
rect 4210 5220 4240 5250
rect 4410 5220 4440 5250
rect 4610 5220 4640 5250
rect 4810 5220 4840 5250
rect 5010 5220 5040 5250
rect 5210 5220 5240 5250
rect 5410 5220 5440 5250
rect 5610 5220 5640 5250
rect 5810 5220 5840 5250
rect 6010 5220 6040 5250
rect 6210 5220 6240 5250
rect 6410 5220 6440 5250
rect -190 5105 -185 5135
rect -185 5105 -165 5135
rect -165 5105 -160 5135
rect 10 5105 40 5135
rect 210 5105 240 5135
rect 410 5105 440 5135
rect 610 5105 640 5135
rect 810 5105 840 5135
rect 1010 5105 1040 5135
rect 1210 5105 1240 5135
rect 1410 5105 1440 5135
rect 1610 5105 1640 5135
rect 1810 5105 1840 5135
rect 2010 5105 2040 5135
rect 2210 5105 2240 5135
rect 2410 5105 2440 5135
rect 2610 5105 2640 5135
rect 2810 5105 2840 5135
rect 3010 5105 3040 5135
rect 3210 5105 3240 5135
rect 3410 5105 3440 5135
rect 3610 5105 3640 5135
rect 3810 5105 3840 5135
rect 4010 5105 4040 5135
rect 4210 5105 4240 5135
rect 4410 5105 4440 5135
rect 4610 5105 4640 5135
rect 4810 5105 4840 5135
rect 5010 5105 5040 5135
rect 5210 5105 5240 5135
rect 5410 5105 5440 5135
rect 5610 5105 5640 5135
rect 5810 5105 5840 5135
rect 6010 5105 6040 5135
rect 6210 5105 6240 5135
rect 6410 5105 6440 5135
rect -190 5035 -185 5065
rect -185 5035 -165 5065
rect -165 5035 -160 5065
rect 10 5035 40 5065
rect 210 5035 240 5065
rect 410 5035 440 5065
rect 610 5035 640 5065
rect 810 5035 840 5065
rect 1010 5035 1040 5065
rect 1210 5035 1240 5065
rect 1410 5035 1440 5065
rect 1610 5035 1640 5065
rect 1810 5035 1840 5065
rect 2010 5035 2040 5065
rect 2210 5035 2240 5065
rect 2410 5035 2440 5065
rect 2610 5035 2640 5065
rect 2810 5035 2840 5065
rect 3010 5035 3040 5065
rect 3210 5035 3240 5065
rect 3410 5035 3440 5065
rect 3610 5035 3640 5065
rect 3810 5035 3840 5065
rect 4010 5035 4040 5065
rect 4210 5035 4240 5065
rect 4410 5035 4440 5065
rect 4610 5035 4640 5065
rect 4810 5035 4840 5065
rect 5010 5035 5040 5065
rect 5210 5035 5240 5065
rect 5410 5035 5440 5065
rect 5610 5035 5640 5065
rect 5810 5035 5840 5065
rect 6010 5035 6040 5065
rect 6210 5035 6240 5065
rect 6410 5035 6440 5065
rect -190 4920 -185 4950
rect -185 4920 -165 4950
rect -165 4920 -160 4950
rect 10 4920 40 4950
rect 210 4920 240 4950
rect 410 4920 440 4950
rect 610 4920 640 4950
rect 810 4920 840 4950
rect 1010 4920 1040 4950
rect 1210 4920 1240 4950
rect 1410 4920 1440 4950
rect 1610 4920 1640 4950
rect 1810 4920 1840 4950
rect 2010 4920 2040 4950
rect 2210 4920 2240 4950
rect 2410 4920 2440 4950
rect 2610 4920 2640 4950
rect 2810 4920 2840 4950
rect 3010 4920 3040 4950
rect 3210 4920 3240 4950
rect 3410 4920 3440 4950
rect 3610 4920 3640 4950
rect 3810 4920 3840 4950
rect 4010 4920 4040 4950
rect 4210 4920 4240 4950
rect 4410 4920 4440 4950
rect 4610 4920 4640 4950
rect 4810 4920 4840 4950
rect 5010 4920 5040 4950
rect 5210 4920 5240 4950
rect 5410 4920 5440 4950
rect 5610 4920 5640 4950
rect 5810 4920 5840 4950
rect 6010 4920 6040 4950
rect 6210 4920 6240 4950
rect 6410 4920 6440 4950
rect -190 4850 -185 4880
rect -185 4850 -165 4880
rect -165 4850 -160 4880
rect 10 4850 40 4880
rect 210 4850 240 4880
rect 410 4850 440 4880
rect 610 4850 640 4880
rect 810 4850 840 4880
rect 1010 4850 1040 4880
rect 1210 4850 1240 4880
rect 1410 4850 1440 4880
rect 1610 4850 1640 4880
rect 1810 4850 1840 4880
rect 2010 4850 2040 4880
rect 2210 4850 2240 4880
rect 2410 4850 2440 4880
rect 2610 4850 2640 4880
rect 2810 4850 2840 4880
rect 3010 4850 3040 4880
rect 3210 4850 3240 4880
rect 3410 4850 3440 4880
rect 3610 4850 3640 4880
rect 3810 4850 3840 4880
rect 4010 4850 4040 4880
rect 4210 4850 4240 4880
rect 4410 4850 4440 4880
rect 4610 4850 4640 4880
rect 4810 4850 4840 4880
rect 5010 4850 5040 4880
rect 5210 4850 5240 4880
rect 5410 4850 5440 4880
rect 5610 4850 5640 4880
rect 5810 4850 5840 4880
rect 6010 4850 6040 4880
rect 6210 4850 6240 4880
rect 6410 4850 6440 4880
rect -190 4735 -185 4765
rect -185 4735 -165 4765
rect -165 4735 -160 4765
rect 10 4735 40 4765
rect 210 4735 240 4765
rect 410 4735 440 4765
rect 610 4735 640 4765
rect 810 4735 840 4765
rect 1010 4735 1040 4765
rect 1210 4735 1240 4765
rect 1410 4735 1440 4765
rect 1610 4735 1640 4765
rect 1810 4735 1840 4765
rect 2010 4735 2040 4765
rect 2210 4735 2240 4765
rect 2410 4735 2440 4765
rect 2610 4735 2640 4765
rect 2810 4735 2840 4765
rect 3010 4735 3040 4765
rect 3210 4735 3240 4765
rect 3410 4735 3440 4765
rect 3610 4735 3640 4765
rect 3810 4735 3840 4765
rect 4010 4735 4040 4765
rect 4210 4735 4240 4765
rect 4410 4735 4440 4765
rect 4610 4735 4640 4765
rect 4810 4735 4840 4765
rect 5010 4735 5040 4765
rect 5210 4735 5240 4765
rect 5410 4735 5440 4765
rect 5610 4735 5640 4765
rect 5810 4735 5840 4765
rect 6010 4735 6040 4765
rect 6210 4735 6240 4765
rect 6410 4735 6440 4765
rect -190 4665 -185 4695
rect -185 4665 -165 4695
rect -165 4665 -160 4695
rect 10 4665 40 4695
rect 210 4665 240 4695
rect 410 4665 440 4695
rect 610 4665 640 4695
rect 810 4665 840 4695
rect 1010 4665 1040 4695
rect 1210 4665 1240 4695
rect 1410 4665 1440 4695
rect 1610 4665 1640 4695
rect 1810 4665 1840 4695
rect 2010 4665 2040 4695
rect 2210 4665 2240 4695
rect 2410 4665 2440 4695
rect 2610 4665 2640 4695
rect 2810 4665 2840 4695
rect 3010 4665 3040 4695
rect 3210 4665 3240 4695
rect 3410 4665 3440 4695
rect 3610 4665 3640 4695
rect 3810 4665 3840 4695
rect 4010 4665 4040 4695
rect 4210 4665 4240 4695
rect 4410 4665 4440 4695
rect 4610 4665 4640 4695
rect 4810 4665 4840 4695
rect 5010 4665 5040 4695
rect 5210 4665 5240 4695
rect 5410 4665 5440 4695
rect 5610 4665 5640 4695
rect 5810 4665 5840 4695
rect 6010 4665 6040 4695
rect 6210 4665 6240 4695
rect 6410 4665 6440 4695
rect -190 4550 -185 4580
rect -185 4550 -165 4580
rect -165 4550 -160 4580
rect 10 4550 40 4580
rect 210 4550 240 4580
rect 410 4550 440 4580
rect 610 4550 640 4580
rect 810 4550 840 4580
rect 1010 4550 1040 4580
rect 1210 4550 1240 4580
rect 1410 4550 1440 4580
rect 1610 4550 1640 4580
rect 1810 4550 1840 4580
rect 2010 4550 2040 4580
rect 2210 4550 2240 4580
rect 2410 4550 2440 4580
rect 2610 4550 2640 4580
rect 2810 4550 2840 4580
rect 3010 4550 3040 4580
rect 3210 4550 3240 4580
rect 3410 4550 3440 4580
rect 3610 4550 3640 4580
rect 3810 4550 3840 4580
rect 4010 4550 4040 4580
rect 4210 4550 4240 4580
rect 4410 4550 4440 4580
rect 4610 4550 4640 4580
rect 4810 4550 4840 4580
rect 5010 4550 5040 4580
rect 5210 4550 5240 4580
rect 5410 4550 5440 4580
rect 5610 4550 5640 4580
rect 5810 4550 5840 4580
rect 6010 4550 6040 4580
rect 6210 4550 6240 4580
rect 6410 4550 6440 4580
rect -190 4480 -185 4510
rect -185 4480 -165 4510
rect -165 4480 -160 4510
rect 10 4480 40 4510
rect 210 4480 240 4510
rect 410 4480 440 4510
rect 610 4480 640 4510
rect 810 4480 840 4510
rect 1010 4480 1040 4510
rect 1210 4480 1240 4510
rect 1410 4480 1440 4510
rect 1610 4480 1640 4510
rect 1810 4480 1840 4510
rect 2010 4480 2040 4510
rect 2210 4480 2240 4510
rect 2410 4480 2440 4510
rect 2610 4480 2640 4510
rect 2810 4480 2840 4510
rect 3010 4480 3040 4510
rect 3210 4480 3240 4510
rect 3410 4480 3440 4510
rect 3610 4480 3640 4510
rect 3810 4480 3840 4510
rect 4010 4480 4040 4510
rect 4210 4480 4240 4510
rect 4410 4480 4440 4510
rect 4610 4480 4640 4510
rect 4810 4480 4840 4510
rect 5010 4480 5040 4510
rect 5210 4480 5240 4510
rect 5410 4480 5440 4510
rect 5610 4480 5640 4510
rect 5810 4480 5840 4510
rect 6010 4480 6040 4510
rect 6210 4480 6240 4510
rect 6410 4480 6440 4510
rect -190 4365 -185 4395
rect -185 4365 -165 4395
rect -165 4365 -160 4395
rect 10 4365 40 4395
rect 210 4365 240 4395
rect 410 4365 440 4395
rect 610 4365 640 4395
rect 810 4365 840 4395
rect 1010 4365 1040 4395
rect 1210 4365 1240 4395
rect 1410 4365 1440 4395
rect 1610 4365 1640 4395
rect 1810 4365 1840 4395
rect 2010 4365 2040 4395
rect 2210 4365 2240 4395
rect 2410 4365 2440 4395
rect 2610 4365 2640 4395
rect 2810 4365 2840 4395
rect 3010 4365 3040 4395
rect 3210 4365 3240 4395
rect 3410 4365 3440 4395
rect 3610 4365 3640 4395
rect 3810 4365 3840 4395
rect 4010 4365 4040 4395
rect 4210 4365 4240 4395
rect 4410 4365 4440 4395
rect 4610 4365 4640 4395
rect 4810 4365 4840 4395
rect 5010 4365 5040 4395
rect 5210 4365 5240 4395
rect 5410 4365 5440 4395
rect 5610 4365 5640 4395
rect 5810 4365 5840 4395
rect 6010 4365 6040 4395
rect 6210 4365 6240 4395
rect 6410 4365 6440 4395
rect -190 4295 -185 4325
rect -185 4295 -165 4325
rect -165 4295 -160 4325
rect 10 4295 40 4325
rect 210 4295 240 4325
rect 410 4295 440 4325
rect 610 4295 640 4325
rect 810 4295 840 4325
rect 1010 4295 1040 4325
rect 1210 4295 1240 4325
rect 1410 4295 1440 4325
rect 1610 4295 1640 4325
rect 1810 4295 1840 4325
rect 2010 4295 2040 4325
rect 2210 4295 2240 4325
rect 2410 4295 2440 4325
rect 2610 4295 2640 4325
rect 2810 4295 2840 4325
rect 3010 4295 3040 4325
rect 3210 4295 3240 4325
rect 3410 4295 3440 4325
rect 3610 4295 3640 4325
rect 3810 4295 3840 4325
rect 4010 4295 4040 4325
rect 4210 4295 4240 4325
rect 4410 4295 4440 4325
rect 4610 4295 4640 4325
rect 4810 4295 4840 4325
rect 5010 4295 5040 4325
rect 5210 4295 5240 4325
rect 5410 4295 5440 4325
rect 5610 4295 5640 4325
rect 5810 4295 5840 4325
rect 6010 4295 6040 4325
rect 6210 4295 6240 4325
rect 6410 4295 6440 4325
rect -190 4180 -185 4210
rect -185 4180 -165 4210
rect -165 4180 -160 4210
rect 10 4180 40 4210
rect 210 4180 240 4210
rect 410 4180 440 4210
rect 610 4180 640 4210
rect 810 4180 840 4210
rect 1010 4180 1040 4210
rect 1210 4180 1240 4210
rect 1410 4180 1440 4210
rect 1610 4180 1640 4210
rect 1810 4180 1840 4210
rect 2010 4180 2040 4210
rect 2210 4180 2240 4210
rect 2410 4180 2440 4210
rect 2610 4180 2640 4210
rect 2810 4180 2840 4210
rect 3010 4180 3040 4210
rect 3210 4180 3240 4210
rect 3410 4180 3440 4210
rect 3610 4180 3640 4210
rect 3810 4180 3840 4210
rect 4010 4180 4040 4210
rect 4210 4180 4240 4210
rect 4410 4180 4440 4210
rect 4610 4180 4640 4210
rect 4810 4180 4840 4210
rect 5010 4180 5040 4210
rect 5210 4180 5240 4210
rect 5410 4180 5440 4210
rect 5610 4180 5640 4210
rect 5810 4180 5840 4210
rect 6010 4180 6040 4210
rect 6210 4180 6240 4210
rect 6410 4180 6440 4210
rect -190 4110 -185 4140
rect -185 4110 -165 4140
rect -165 4110 -160 4140
rect 10 4110 40 4140
rect 210 4110 240 4140
rect 410 4110 440 4140
rect 610 4110 640 4140
rect 810 4110 840 4140
rect 1010 4110 1040 4140
rect 1210 4110 1240 4140
rect 1410 4110 1440 4140
rect 1610 4110 1640 4140
rect 1810 4110 1840 4140
rect 2010 4110 2040 4140
rect 2210 4110 2240 4140
rect 2410 4110 2440 4140
rect 2610 4110 2640 4140
rect 2810 4110 2840 4140
rect 3010 4110 3040 4140
rect 3210 4110 3240 4140
rect 3410 4110 3440 4140
rect 3610 4110 3640 4140
rect 3810 4110 3840 4140
rect 4010 4110 4040 4140
rect 4210 4110 4240 4140
rect 4410 4110 4440 4140
rect 4610 4110 4640 4140
rect 4810 4110 4840 4140
rect 5010 4110 5040 4140
rect 5210 4110 5240 4140
rect 5410 4110 5440 4140
rect 5610 4110 5640 4140
rect 5810 4110 5840 4140
rect 6010 4110 6040 4140
rect 6210 4110 6240 4140
rect 6410 4110 6440 4140
rect -190 3995 -185 4025
rect -185 3995 -165 4025
rect -165 3995 -160 4025
rect 10 3995 40 4025
rect 210 3995 240 4025
rect 410 3995 440 4025
rect 610 3995 640 4025
rect 810 3995 840 4025
rect 1010 3995 1040 4025
rect 1210 3995 1240 4025
rect 1410 3995 1440 4025
rect 1610 3995 1640 4025
rect 1810 3995 1840 4025
rect 2010 3995 2040 4025
rect 2210 3995 2240 4025
rect 2410 3995 2440 4025
rect 2610 3995 2640 4025
rect 2810 3995 2840 4025
rect 3010 3995 3040 4025
rect 3210 3995 3240 4025
rect 3410 3995 3440 4025
rect 3610 3995 3640 4025
rect 3810 3995 3840 4025
rect 4010 3995 4040 4025
rect 4210 3995 4240 4025
rect 4410 3995 4440 4025
rect 4610 3995 4640 4025
rect 4810 3995 4840 4025
rect 5010 3995 5040 4025
rect 5210 3995 5240 4025
rect 5410 3995 5440 4025
rect 5610 3995 5640 4025
rect 5810 3995 5840 4025
rect 6010 3995 6040 4025
rect 6210 3995 6240 4025
rect 6410 3995 6440 4025
rect -190 3925 -185 3955
rect -185 3925 -165 3955
rect -165 3925 -160 3955
rect 10 3925 40 3955
rect 210 3925 240 3955
rect 410 3925 440 3955
rect 610 3925 640 3955
rect 810 3925 840 3955
rect 1010 3925 1040 3955
rect 1210 3925 1240 3955
rect 1410 3925 1440 3955
rect 1610 3925 1640 3955
rect 1810 3925 1840 3955
rect 2010 3925 2040 3955
rect 2210 3925 2240 3955
rect 2410 3925 2440 3955
rect 2610 3925 2640 3955
rect 2810 3925 2840 3955
rect 3010 3925 3040 3955
rect 3210 3925 3240 3955
rect 3410 3925 3440 3955
rect 3610 3925 3640 3955
rect 3810 3925 3840 3955
rect 4010 3925 4040 3955
rect 4210 3925 4240 3955
rect 4410 3925 4440 3955
rect 4610 3925 4640 3955
rect 4810 3925 4840 3955
rect 5010 3925 5040 3955
rect 5210 3925 5240 3955
rect 5410 3925 5440 3955
rect 5610 3925 5640 3955
rect 5810 3925 5840 3955
rect 6010 3925 6040 3955
rect 6210 3925 6240 3955
rect 6410 3925 6440 3955
rect -190 3810 -185 3840
rect -185 3810 -165 3840
rect -165 3810 -160 3840
rect 10 3810 40 3840
rect 210 3810 240 3840
rect 410 3810 440 3840
rect 610 3810 640 3840
rect 810 3810 840 3840
rect 1010 3810 1040 3840
rect 1210 3810 1240 3840
rect 1410 3810 1440 3840
rect 1610 3810 1640 3840
rect 1810 3810 1840 3840
rect 2010 3810 2040 3840
rect 2210 3810 2240 3840
rect 2410 3810 2440 3840
rect 2610 3810 2640 3840
rect 2810 3810 2840 3840
rect 3010 3810 3040 3840
rect 3210 3810 3240 3840
rect 3410 3810 3440 3840
rect 3610 3810 3640 3840
rect 3810 3810 3840 3840
rect 4010 3810 4040 3840
rect 4210 3810 4240 3840
rect 4410 3810 4440 3840
rect 4610 3810 4640 3840
rect 4810 3810 4840 3840
rect 5010 3810 5040 3840
rect 5210 3810 5240 3840
rect 5410 3810 5440 3840
rect 5610 3810 5640 3840
rect 5810 3810 5840 3840
rect 6010 3810 6040 3840
rect 6210 3810 6240 3840
rect 6410 3810 6440 3840
rect -190 3740 -185 3770
rect -185 3740 -165 3770
rect -165 3740 -160 3770
rect 10 3740 40 3770
rect 210 3740 240 3770
rect 410 3740 440 3770
rect 610 3740 640 3770
rect 810 3740 840 3770
rect 1010 3740 1040 3770
rect 1210 3740 1240 3770
rect 1410 3740 1440 3770
rect 1610 3740 1640 3770
rect 1810 3740 1840 3770
rect 2010 3740 2040 3770
rect 2210 3740 2240 3770
rect 2410 3740 2440 3770
rect 2610 3740 2640 3770
rect 2810 3740 2840 3770
rect 3010 3740 3040 3770
rect 3210 3740 3240 3770
rect 3410 3740 3440 3770
rect 3610 3740 3640 3770
rect 3810 3740 3840 3770
rect 4010 3740 4040 3770
rect 4210 3740 4240 3770
rect 4410 3740 4440 3770
rect 4610 3740 4640 3770
rect 4810 3740 4840 3770
rect 5010 3740 5040 3770
rect 5210 3740 5240 3770
rect 5410 3740 5440 3770
rect 5610 3740 5640 3770
rect 5810 3740 5840 3770
rect 6010 3740 6040 3770
rect 6210 3740 6240 3770
rect 6410 3740 6440 3770
rect -190 3625 -185 3655
rect -185 3625 -165 3655
rect -165 3625 -160 3655
rect 10 3625 40 3655
rect 210 3625 240 3655
rect 410 3625 440 3655
rect 610 3625 640 3655
rect 810 3625 840 3655
rect 1010 3625 1040 3655
rect 1210 3625 1240 3655
rect 1410 3625 1440 3655
rect 1610 3625 1640 3655
rect 1810 3625 1840 3655
rect 2010 3625 2040 3655
rect 2210 3625 2240 3655
rect 2410 3625 2440 3655
rect 2610 3625 2640 3655
rect 2810 3625 2840 3655
rect 3010 3625 3040 3655
rect 3210 3625 3240 3655
rect 3410 3625 3440 3655
rect 3610 3625 3640 3655
rect 3810 3625 3840 3655
rect 4010 3625 4040 3655
rect 4210 3625 4240 3655
rect 4410 3625 4440 3655
rect 4610 3625 4640 3655
rect 4810 3625 4840 3655
rect 5010 3625 5040 3655
rect 5210 3625 5240 3655
rect 5410 3625 5440 3655
rect 5610 3625 5640 3655
rect 5810 3625 5840 3655
rect 6010 3625 6040 3655
rect 6210 3625 6240 3655
rect 6410 3625 6440 3655
rect -190 3555 -185 3585
rect -185 3555 -165 3585
rect -165 3555 -160 3585
rect 10 3555 40 3585
rect 210 3555 240 3585
rect 410 3555 440 3585
rect 610 3555 640 3585
rect 810 3555 840 3585
rect 1010 3555 1040 3585
rect 1210 3555 1240 3585
rect 1410 3555 1440 3585
rect 1610 3555 1640 3585
rect 1810 3555 1840 3585
rect 2010 3555 2040 3585
rect 2210 3555 2240 3585
rect 2410 3555 2440 3585
rect 2610 3555 2640 3585
rect 2810 3555 2840 3585
rect 3010 3555 3040 3585
rect 3210 3555 3240 3585
rect 3410 3555 3440 3585
rect 3610 3555 3640 3585
rect 3810 3555 3840 3585
rect 4010 3555 4040 3585
rect 4210 3555 4240 3585
rect 4410 3555 4440 3585
rect 4610 3555 4640 3585
rect 4810 3555 4840 3585
rect 5010 3555 5040 3585
rect 5210 3555 5240 3585
rect 5410 3555 5440 3585
rect 5610 3555 5640 3585
rect 5810 3555 5840 3585
rect 6010 3555 6040 3585
rect 6210 3555 6240 3585
rect 6410 3555 6440 3585
rect -190 3440 -185 3470
rect -185 3440 -165 3470
rect -165 3440 -160 3470
rect 10 3440 40 3470
rect 210 3440 240 3470
rect 410 3440 440 3470
rect 610 3440 640 3470
rect 810 3440 840 3470
rect 1010 3440 1040 3470
rect 1210 3440 1240 3470
rect 1410 3440 1440 3470
rect 1610 3440 1640 3470
rect 1810 3440 1840 3470
rect 2010 3440 2040 3470
rect 2210 3440 2240 3470
rect 2410 3440 2440 3470
rect 2610 3440 2640 3470
rect 2810 3440 2840 3470
rect 3010 3440 3040 3470
rect 3210 3440 3240 3470
rect 3410 3440 3440 3470
rect 3610 3440 3640 3470
rect 3810 3440 3840 3470
rect 4010 3440 4040 3470
rect 4210 3440 4240 3470
rect 4410 3440 4440 3470
rect 4610 3440 4640 3470
rect 4810 3440 4840 3470
rect 5010 3440 5040 3470
rect 5210 3440 5240 3470
rect 5410 3440 5440 3470
rect 5610 3440 5640 3470
rect 5810 3440 5840 3470
rect 6010 3440 6040 3470
rect 6210 3440 6240 3470
rect 6410 3440 6440 3470
rect -190 3370 -185 3400
rect -185 3370 -165 3400
rect -165 3370 -160 3400
rect 10 3370 40 3400
rect 210 3370 240 3400
rect 410 3370 440 3400
rect 610 3370 640 3400
rect 810 3370 840 3400
rect 1010 3370 1040 3400
rect 1210 3370 1240 3400
rect 1410 3370 1440 3400
rect 1610 3370 1640 3400
rect 1810 3370 1840 3400
rect 2010 3370 2040 3400
rect 2210 3370 2240 3400
rect 2410 3370 2440 3400
rect 2610 3370 2640 3400
rect 2810 3370 2840 3400
rect 3010 3370 3040 3400
rect 3210 3370 3240 3400
rect 3410 3370 3440 3400
rect 3610 3370 3640 3400
rect 3810 3370 3840 3400
rect 4010 3370 4040 3400
rect 4210 3370 4240 3400
rect 4410 3370 4440 3400
rect 4610 3370 4640 3400
rect 4810 3370 4840 3400
rect 5010 3370 5040 3400
rect 5210 3370 5240 3400
rect 5410 3370 5440 3400
rect 5610 3370 5640 3400
rect 5810 3370 5840 3400
rect 6010 3370 6040 3400
rect 6210 3370 6240 3400
rect 6410 3370 6440 3400
rect -190 3255 -185 3285
rect -185 3255 -165 3285
rect -165 3255 -160 3285
rect 10 3255 40 3285
rect 210 3255 240 3285
rect 410 3255 440 3285
rect 610 3255 640 3285
rect 810 3255 840 3285
rect 1010 3255 1040 3285
rect 1210 3255 1240 3285
rect 1410 3255 1440 3285
rect 1610 3255 1640 3285
rect 1810 3255 1840 3285
rect 2010 3255 2040 3285
rect 2210 3255 2240 3285
rect 2410 3255 2440 3285
rect 2610 3255 2640 3285
rect 2810 3255 2840 3285
rect 3010 3255 3040 3285
rect 3210 3255 3240 3285
rect 3410 3255 3440 3285
rect 3610 3255 3640 3285
rect 3810 3255 3840 3285
rect 4010 3255 4040 3285
rect 4210 3255 4240 3285
rect 4410 3255 4440 3285
rect 4610 3255 4640 3285
rect 4810 3255 4840 3285
rect 5010 3255 5040 3285
rect 5210 3255 5240 3285
rect 5410 3255 5440 3285
rect 5610 3255 5640 3285
rect 5810 3255 5840 3285
rect 6010 3255 6040 3285
rect 6210 3255 6240 3285
rect 6410 3255 6440 3285
rect -190 3185 -185 3215
rect -185 3185 -165 3215
rect -165 3185 -160 3215
rect 10 3185 40 3215
rect 210 3185 240 3215
rect 410 3185 440 3215
rect 610 3185 640 3215
rect 810 3185 840 3215
rect 1010 3185 1040 3215
rect 1210 3185 1240 3215
rect 1410 3185 1440 3215
rect 1610 3185 1640 3215
rect 1810 3185 1840 3215
rect 2010 3185 2040 3215
rect 2210 3185 2240 3215
rect 2410 3185 2440 3215
rect 2610 3185 2640 3215
rect 2810 3185 2840 3215
rect 3010 3185 3040 3215
rect 3210 3185 3240 3215
rect 3410 3185 3440 3215
rect 3610 3185 3640 3215
rect 3810 3185 3840 3215
rect 4010 3185 4040 3215
rect 4210 3185 4240 3215
rect 4410 3185 4440 3215
rect 4610 3185 4640 3215
rect 4810 3185 4840 3215
rect 5010 3185 5040 3215
rect 5210 3185 5240 3215
rect 5410 3185 5440 3215
rect 5610 3185 5640 3215
rect 5810 3185 5840 3215
rect 6010 3185 6040 3215
rect 6210 3185 6240 3215
rect 6410 3185 6440 3215
rect -190 3070 -185 3100
rect -185 3070 -165 3100
rect -165 3070 -160 3100
rect 10 3070 40 3100
rect 210 3070 240 3100
rect 410 3070 440 3100
rect 610 3070 640 3100
rect 810 3070 840 3100
rect 1010 3070 1040 3100
rect 1210 3070 1240 3100
rect 1410 3070 1440 3100
rect 1610 3070 1640 3100
rect 1810 3070 1840 3100
rect 2010 3070 2040 3100
rect 2210 3070 2240 3100
rect 2410 3070 2440 3100
rect 2610 3070 2640 3100
rect 2810 3070 2840 3100
rect 3010 3070 3040 3100
rect 3210 3070 3240 3100
rect 3410 3070 3440 3100
rect 3610 3070 3640 3100
rect 3810 3070 3840 3100
rect 4010 3070 4040 3100
rect 4210 3070 4240 3100
rect 4410 3070 4440 3100
rect 4610 3070 4640 3100
rect 4810 3070 4840 3100
rect 5010 3070 5040 3100
rect 5210 3070 5240 3100
rect 5410 3070 5440 3100
rect 5610 3070 5640 3100
rect 5810 3070 5840 3100
rect 6010 3070 6040 3100
rect 6210 3070 6240 3100
rect 6410 3070 6440 3100
rect -190 3000 -185 3030
rect -185 3000 -165 3030
rect -165 3000 -160 3030
rect 10 3000 40 3030
rect 210 3000 240 3030
rect 410 3000 440 3030
rect 610 3000 640 3030
rect 810 3000 840 3030
rect 1010 3000 1040 3030
rect 1210 3000 1240 3030
rect 1410 3000 1440 3030
rect 1610 3000 1640 3030
rect 1810 3000 1840 3030
rect 2010 3000 2040 3030
rect 2210 3000 2240 3030
rect 2410 3000 2440 3030
rect 2610 3000 2640 3030
rect 2810 3000 2840 3030
rect 3010 3000 3040 3030
rect 3210 3000 3240 3030
rect 3410 3000 3440 3030
rect 3610 3000 3640 3030
rect 3810 3000 3840 3030
rect 4010 3000 4040 3030
rect 4210 3000 4240 3030
rect 4410 3000 4440 3030
rect 4610 3000 4640 3030
rect 4810 3000 4840 3030
rect 5010 3000 5040 3030
rect 5210 3000 5240 3030
rect 5410 3000 5440 3030
rect 5610 3000 5640 3030
rect 5810 3000 5840 3030
rect 6010 3000 6040 3030
rect 6210 3000 6240 3030
rect 6410 3000 6440 3030
rect -190 2885 -185 2915
rect -185 2885 -165 2915
rect -165 2885 -160 2915
rect 10 2885 40 2915
rect 210 2885 240 2915
rect 410 2885 440 2915
rect 610 2885 640 2915
rect 810 2885 840 2915
rect 1010 2885 1040 2915
rect 1210 2885 1240 2915
rect 1410 2885 1440 2915
rect 1610 2885 1640 2915
rect 1810 2885 1840 2915
rect 2010 2885 2040 2915
rect 2210 2885 2240 2915
rect 2410 2885 2440 2915
rect 2610 2885 2640 2915
rect 2810 2885 2840 2915
rect 3010 2885 3040 2915
rect 3210 2885 3240 2915
rect 3410 2885 3440 2915
rect 3610 2885 3640 2915
rect 3810 2885 3840 2915
rect 4010 2885 4040 2915
rect 4210 2885 4240 2915
rect 4410 2885 4440 2915
rect 4610 2885 4640 2915
rect 4810 2885 4840 2915
rect 5010 2885 5040 2915
rect 5210 2885 5240 2915
rect 5410 2885 5440 2915
rect 5610 2885 5640 2915
rect 5810 2885 5840 2915
rect 6010 2885 6040 2915
rect 6210 2885 6240 2915
rect 6410 2885 6440 2915
rect -190 2815 -185 2845
rect -185 2815 -165 2845
rect -165 2815 -160 2845
rect 10 2815 40 2845
rect 210 2815 240 2845
rect 410 2815 440 2845
rect 610 2815 640 2845
rect 810 2815 840 2845
rect 1010 2815 1040 2845
rect 1210 2815 1240 2845
rect 1410 2815 1440 2845
rect 1610 2815 1640 2845
rect 1810 2815 1840 2845
rect 2010 2815 2040 2845
rect 2210 2815 2240 2845
rect 2410 2815 2440 2845
rect 2610 2815 2640 2845
rect 2810 2815 2840 2845
rect 3010 2815 3040 2845
rect 3210 2815 3240 2845
rect 3410 2815 3440 2845
rect 3610 2815 3640 2845
rect 3810 2815 3840 2845
rect 4010 2815 4040 2845
rect 4210 2815 4240 2845
rect 4410 2815 4440 2845
rect 4610 2815 4640 2845
rect 4810 2815 4840 2845
rect 5010 2815 5040 2845
rect 5210 2815 5240 2845
rect 5410 2815 5440 2845
rect 5610 2815 5640 2845
rect 5810 2815 5840 2845
rect 6010 2815 6040 2845
rect 6210 2815 6240 2845
rect 6410 2815 6440 2845
rect -190 2700 -185 2730
rect -185 2700 -165 2730
rect -165 2700 -160 2730
rect 10 2700 40 2730
rect 210 2700 240 2730
rect 410 2700 440 2730
rect 610 2700 640 2730
rect 810 2700 840 2730
rect 1010 2700 1040 2730
rect 1210 2700 1240 2730
rect 1410 2700 1440 2730
rect 1610 2700 1640 2730
rect 1810 2700 1840 2730
rect 2010 2700 2040 2730
rect 2210 2700 2240 2730
rect 2410 2700 2440 2730
rect 2610 2700 2640 2730
rect 2810 2700 2840 2730
rect 3010 2700 3040 2730
rect 3210 2700 3240 2730
rect 3410 2700 3440 2730
rect 3610 2700 3640 2730
rect 3810 2700 3840 2730
rect 4010 2700 4040 2730
rect 4210 2700 4240 2730
rect 4410 2700 4440 2730
rect 4610 2700 4640 2730
rect 4810 2700 4840 2730
rect 5010 2700 5040 2730
rect 5210 2700 5240 2730
rect 5410 2700 5440 2730
rect 5610 2700 5640 2730
rect 5810 2700 5840 2730
rect 6010 2700 6040 2730
rect 6210 2700 6240 2730
rect 6410 2700 6440 2730
rect -190 2630 -185 2660
rect -185 2630 -165 2660
rect -165 2630 -160 2660
rect 10 2630 40 2660
rect 210 2630 240 2660
rect 410 2630 440 2660
rect 610 2630 640 2660
rect 810 2630 840 2660
rect 1010 2630 1040 2660
rect 1210 2630 1240 2660
rect 1410 2630 1440 2660
rect 1610 2630 1640 2660
rect 1810 2630 1840 2660
rect 2010 2630 2040 2660
rect 2210 2630 2240 2660
rect 2410 2630 2440 2660
rect 2610 2630 2640 2660
rect 2810 2630 2840 2660
rect 3010 2630 3040 2660
rect 3210 2630 3240 2660
rect 3410 2630 3440 2660
rect 3610 2630 3640 2660
rect 3810 2630 3840 2660
rect 4010 2630 4040 2660
rect 4210 2630 4240 2660
rect 4410 2630 4440 2660
rect 4610 2630 4640 2660
rect 4810 2630 4840 2660
rect 5010 2630 5040 2660
rect 5210 2630 5240 2660
rect 5410 2630 5440 2660
rect 5610 2630 5640 2660
rect 5810 2630 5840 2660
rect 6010 2630 6040 2660
rect 6210 2630 6240 2660
rect 6410 2630 6440 2660
rect -190 2515 -185 2545
rect -185 2515 -165 2545
rect -165 2515 -160 2545
rect 10 2515 40 2545
rect 210 2515 240 2545
rect 410 2515 440 2545
rect 610 2515 640 2545
rect 810 2515 840 2545
rect 1010 2515 1040 2545
rect 1210 2515 1240 2545
rect 1410 2515 1440 2545
rect 1610 2515 1640 2545
rect 1810 2515 1840 2545
rect 2010 2515 2040 2545
rect 2210 2515 2240 2545
rect 2410 2515 2440 2545
rect 2610 2515 2640 2545
rect 2810 2515 2840 2545
rect 3010 2515 3040 2545
rect 3210 2515 3240 2545
rect 3410 2515 3440 2545
rect 3610 2515 3640 2545
rect 3810 2515 3840 2545
rect 4010 2515 4040 2545
rect 4210 2515 4240 2545
rect 4410 2515 4440 2545
rect 4610 2515 4640 2545
rect 4810 2515 4840 2545
rect 5010 2515 5040 2545
rect 5210 2515 5240 2545
rect 5410 2515 5440 2545
rect 5610 2515 5640 2545
rect 5810 2515 5840 2545
rect 6010 2515 6040 2545
rect 6210 2515 6240 2545
rect 6410 2515 6440 2545
rect -190 2445 -185 2475
rect -185 2445 -165 2475
rect -165 2445 -160 2475
rect 10 2445 40 2475
rect 210 2445 240 2475
rect 410 2445 440 2475
rect 610 2445 640 2475
rect 810 2445 840 2475
rect 1010 2445 1040 2475
rect 1210 2445 1240 2475
rect 1410 2445 1440 2475
rect 1610 2445 1640 2475
rect 1810 2445 1840 2475
rect 2010 2445 2040 2475
rect 2210 2445 2240 2475
rect 2410 2445 2440 2475
rect 2610 2445 2640 2475
rect 2810 2445 2840 2475
rect 3010 2445 3040 2475
rect 3210 2445 3240 2475
rect 3410 2445 3440 2475
rect 3610 2445 3640 2475
rect 3810 2445 3840 2475
rect 4010 2445 4040 2475
rect 4210 2445 4240 2475
rect 4410 2445 4440 2475
rect 4610 2445 4640 2475
rect 4810 2445 4840 2475
rect 5010 2445 5040 2475
rect 5210 2445 5240 2475
rect 5410 2445 5440 2475
rect 5610 2445 5640 2475
rect 5810 2445 5840 2475
rect 6010 2445 6040 2475
rect 6210 2445 6240 2475
rect 6410 2445 6440 2475
rect -190 2330 -185 2360
rect -185 2330 -165 2360
rect -165 2330 -160 2360
rect 10 2330 40 2360
rect 210 2330 240 2360
rect 410 2330 440 2360
rect 610 2330 640 2360
rect 810 2330 840 2360
rect 1010 2330 1040 2360
rect 1210 2330 1240 2360
rect 1410 2330 1440 2360
rect 1610 2330 1640 2360
rect 1810 2330 1840 2360
rect 2010 2330 2040 2360
rect 2210 2330 2240 2360
rect 2410 2330 2440 2360
rect 2610 2330 2640 2360
rect 2810 2330 2840 2360
rect 3010 2330 3040 2360
rect 3210 2330 3240 2360
rect 3410 2330 3440 2360
rect 3610 2330 3640 2360
rect 3810 2330 3840 2360
rect 4010 2330 4040 2360
rect 4210 2330 4240 2360
rect 4410 2330 4440 2360
rect 4610 2330 4640 2360
rect 4810 2330 4840 2360
rect 5010 2330 5040 2360
rect 5210 2330 5240 2360
rect 5410 2330 5440 2360
rect 5610 2330 5640 2360
rect 5810 2330 5840 2360
rect 6010 2330 6040 2360
rect 6210 2330 6240 2360
rect 6410 2330 6440 2360
rect -190 2260 -185 2290
rect -185 2260 -165 2290
rect -165 2260 -160 2290
rect 10 2260 40 2290
rect 210 2260 240 2290
rect 410 2260 440 2290
rect 610 2260 640 2290
rect 810 2260 840 2290
rect 1010 2260 1040 2290
rect 1210 2260 1240 2290
rect 1410 2260 1440 2290
rect 1610 2260 1640 2290
rect 1810 2260 1840 2290
rect 2010 2260 2040 2290
rect 2210 2260 2240 2290
rect 2410 2260 2440 2290
rect 2610 2260 2640 2290
rect 2810 2260 2840 2290
rect 3010 2260 3040 2290
rect 3210 2260 3240 2290
rect 3410 2260 3440 2290
rect 3610 2260 3640 2290
rect 3810 2260 3840 2290
rect 4010 2260 4040 2290
rect 4210 2260 4240 2290
rect 4410 2260 4440 2290
rect 4610 2260 4640 2290
rect 4810 2260 4840 2290
rect 5010 2260 5040 2290
rect 5210 2260 5240 2290
rect 5410 2260 5440 2290
rect 5610 2260 5640 2290
rect 5810 2260 5840 2290
rect 6010 2260 6040 2290
rect 6210 2260 6240 2290
rect 6410 2260 6440 2290
rect -190 2145 -185 2175
rect -185 2145 -165 2175
rect -165 2145 -160 2175
rect 10 2145 40 2175
rect 210 2145 240 2175
rect 410 2145 440 2175
rect 610 2145 640 2175
rect 810 2145 840 2175
rect 1010 2145 1040 2175
rect 1210 2145 1240 2175
rect 1410 2145 1440 2175
rect 1610 2145 1640 2175
rect 1810 2145 1840 2175
rect 2010 2145 2040 2175
rect 2210 2145 2240 2175
rect 2410 2145 2440 2175
rect 2610 2145 2640 2175
rect 2810 2145 2840 2175
rect 3010 2145 3040 2175
rect 3210 2145 3240 2175
rect 3410 2145 3440 2175
rect 3610 2145 3640 2175
rect 3810 2145 3840 2175
rect 4010 2145 4040 2175
rect 4210 2145 4240 2175
rect 4410 2145 4440 2175
rect 4610 2145 4640 2175
rect 4810 2145 4840 2175
rect 5010 2145 5040 2175
rect 5210 2145 5240 2175
rect 5410 2145 5440 2175
rect 5610 2145 5640 2175
rect 5810 2145 5840 2175
rect 6010 2145 6040 2175
rect 6210 2145 6240 2175
rect 6410 2145 6440 2175
rect -190 2075 -185 2105
rect -185 2075 -165 2105
rect -165 2075 -160 2105
rect 10 2075 40 2105
rect 210 2075 240 2105
rect 410 2075 440 2105
rect 610 2075 640 2105
rect 810 2075 840 2105
rect 1010 2075 1040 2105
rect 1210 2075 1240 2105
rect 1410 2075 1440 2105
rect 1610 2075 1640 2105
rect 1810 2075 1840 2105
rect 2010 2075 2040 2105
rect 2210 2075 2240 2105
rect 2410 2075 2440 2105
rect 2610 2075 2640 2105
rect 2810 2075 2840 2105
rect 3010 2075 3040 2105
rect 3210 2075 3240 2105
rect 3410 2075 3440 2105
rect 3610 2075 3640 2105
rect 3810 2075 3840 2105
rect 4010 2075 4040 2105
rect 4210 2075 4240 2105
rect 4410 2075 4440 2105
rect 4610 2075 4640 2105
rect 4810 2075 4840 2105
rect 5010 2075 5040 2105
rect 5210 2075 5240 2105
rect 5410 2075 5440 2105
rect 5610 2075 5640 2105
rect 5810 2075 5840 2105
rect 6010 2075 6040 2105
rect 6210 2075 6240 2105
rect 6410 2075 6440 2105
rect -190 1960 -185 1990
rect -185 1960 -165 1990
rect -165 1960 -160 1990
rect 10 1960 40 1990
rect 210 1960 240 1990
rect 410 1960 440 1990
rect 610 1960 640 1990
rect 810 1960 840 1990
rect 1010 1960 1040 1990
rect 1210 1960 1240 1990
rect 1410 1960 1440 1990
rect 1610 1960 1640 1990
rect 1810 1960 1840 1990
rect 2010 1960 2040 1990
rect 2210 1960 2240 1990
rect 2410 1960 2440 1990
rect 2610 1960 2640 1990
rect 2810 1960 2840 1990
rect 3010 1960 3040 1990
rect 3210 1960 3240 1990
rect 3410 1960 3440 1990
rect 3610 1960 3640 1990
rect 3810 1960 3840 1990
rect 4010 1960 4040 1990
rect 4210 1960 4240 1990
rect 4410 1960 4440 1990
rect 4610 1960 4640 1990
rect 4810 1960 4840 1990
rect 5010 1960 5040 1990
rect 5210 1960 5240 1990
rect 5410 1960 5440 1990
rect 5610 1960 5640 1990
rect 5810 1960 5840 1990
rect 6010 1960 6040 1990
rect 6210 1960 6240 1990
rect 6410 1960 6440 1990
rect -190 1890 -185 1920
rect -185 1890 -165 1920
rect -165 1890 -160 1920
rect 10 1890 40 1920
rect 210 1890 240 1920
rect 410 1890 440 1920
rect 610 1890 640 1920
rect 810 1890 840 1920
rect 1010 1890 1040 1920
rect 1210 1890 1240 1920
rect 1410 1890 1440 1920
rect 1610 1890 1640 1920
rect 1810 1890 1840 1920
rect 2010 1890 2040 1920
rect 2210 1890 2240 1920
rect 2410 1890 2440 1920
rect 2610 1890 2640 1920
rect 2810 1890 2840 1920
rect 3010 1890 3040 1920
rect 3210 1890 3240 1920
rect 3410 1890 3440 1920
rect 3610 1890 3640 1920
rect 3810 1890 3840 1920
rect 4010 1890 4040 1920
rect 4210 1890 4240 1920
rect 4410 1890 4440 1920
rect 4610 1890 4640 1920
rect 4810 1890 4840 1920
rect 5010 1890 5040 1920
rect 5210 1890 5240 1920
rect 5410 1890 5440 1920
rect 5610 1890 5640 1920
rect 5810 1890 5840 1920
rect 6010 1890 6040 1920
rect 6210 1890 6240 1920
rect 6410 1890 6440 1920
rect -190 1775 -185 1805
rect -185 1775 -165 1805
rect -165 1775 -160 1805
rect 10 1775 40 1805
rect 210 1775 240 1805
rect 410 1775 440 1805
rect 610 1775 640 1805
rect 810 1775 840 1805
rect 1010 1775 1040 1805
rect 1210 1775 1240 1805
rect 1410 1775 1440 1805
rect 1610 1775 1640 1805
rect 1810 1775 1840 1805
rect 2010 1775 2040 1805
rect 2210 1775 2240 1805
rect 2410 1775 2440 1805
rect 2610 1775 2640 1805
rect 2810 1775 2840 1805
rect 3010 1775 3040 1805
rect 3210 1775 3240 1805
rect 3410 1775 3440 1805
rect 3610 1775 3640 1805
rect 3810 1775 3840 1805
rect 4010 1775 4040 1805
rect 4210 1775 4240 1805
rect 4410 1775 4440 1805
rect 4610 1775 4640 1805
rect 4810 1775 4840 1805
rect 5010 1775 5040 1805
rect 5210 1775 5240 1805
rect 5410 1775 5440 1805
rect 5610 1775 5640 1805
rect 5810 1775 5840 1805
rect 6010 1775 6040 1805
rect 6210 1775 6240 1805
rect 6410 1775 6440 1805
rect -190 1705 -185 1735
rect -185 1705 -165 1735
rect -165 1705 -160 1735
rect 10 1705 40 1735
rect 210 1705 240 1735
rect 410 1705 440 1735
rect 610 1705 640 1735
rect 810 1705 840 1735
rect 1010 1705 1040 1735
rect 1210 1705 1240 1735
rect 1410 1705 1440 1735
rect 1610 1705 1640 1735
rect 1810 1705 1840 1735
rect 2010 1705 2040 1735
rect 2210 1705 2240 1735
rect 2410 1705 2440 1735
rect 2610 1705 2640 1735
rect 2810 1705 2840 1735
rect 3010 1705 3040 1735
rect 3210 1705 3240 1735
rect 3410 1705 3440 1735
rect 3610 1705 3640 1735
rect 3810 1705 3840 1735
rect 4010 1705 4040 1735
rect 4210 1705 4240 1735
rect 4410 1705 4440 1735
rect 4610 1705 4640 1735
rect 4810 1705 4840 1735
rect 5010 1705 5040 1735
rect 5210 1705 5240 1735
rect 5410 1705 5440 1735
rect 5610 1705 5640 1735
rect 5810 1705 5840 1735
rect 6010 1705 6040 1735
rect 6210 1705 6240 1735
rect 6410 1705 6440 1735
rect -190 1590 -185 1620
rect -185 1590 -165 1620
rect -165 1590 -160 1620
rect 10 1590 40 1620
rect 210 1590 240 1620
rect 410 1590 440 1620
rect 610 1590 640 1620
rect 810 1590 840 1620
rect 1010 1590 1040 1620
rect 1210 1590 1240 1620
rect 1410 1590 1440 1620
rect 1610 1590 1640 1620
rect 1810 1590 1840 1620
rect 2010 1590 2040 1620
rect 2210 1590 2240 1620
rect 2410 1590 2440 1620
rect 2610 1590 2640 1620
rect 2810 1590 2840 1620
rect 3010 1590 3040 1620
rect 3210 1590 3240 1620
rect 3410 1590 3440 1620
rect 3610 1590 3640 1620
rect 3810 1590 3840 1620
rect 4010 1590 4040 1620
rect 4210 1590 4240 1620
rect 4410 1590 4440 1620
rect 4610 1590 4640 1620
rect 4810 1590 4840 1620
rect 5010 1590 5040 1620
rect 5210 1590 5240 1620
rect 5410 1590 5440 1620
rect 5610 1590 5640 1620
rect 5810 1590 5840 1620
rect 6010 1590 6040 1620
rect 6210 1590 6240 1620
rect 6410 1590 6440 1620
rect -190 1520 -185 1550
rect -185 1520 -165 1550
rect -165 1520 -160 1550
rect 10 1520 40 1550
rect 210 1520 240 1550
rect 410 1520 440 1550
rect 610 1520 640 1550
rect 810 1520 840 1550
rect 1010 1520 1040 1550
rect 1210 1520 1240 1550
rect 1410 1520 1440 1550
rect 1610 1520 1640 1550
rect 1810 1520 1840 1550
rect 2010 1520 2040 1550
rect 2210 1520 2240 1550
rect 2410 1520 2440 1550
rect 2610 1520 2640 1550
rect 2810 1520 2840 1550
rect 3010 1520 3040 1550
rect 3210 1520 3240 1550
rect 3410 1520 3440 1550
rect 3610 1520 3640 1550
rect 3810 1520 3840 1550
rect 4010 1520 4040 1550
rect 4210 1520 4240 1550
rect 4410 1520 4440 1550
rect 4610 1520 4640 1550
rect 4810 1520 4840 1550
rect 5010 1520 5040 1550
rect 5210 1520 5240 1550
rect 5410 1520 5440 1550
rect 5610 1520 5640 1550
rect 5810 1520 5840 1550
rect 6010 1520 6040 1550
rect 6210 1520 6240 1550
rect 6410 1520 6440 1550
rect -190 1405 -185 1435
rect -185 1405 -165 1435
rect -165 1405 -160 1435
rect 10 1405 40 1435
rect 210 1405 240 1435
rect 410 1405 440 1435
rect 610 1405 640 1435
rect 810 1405 840 1435
rect 1010 1405 1040 1435
rect 1210 1405 1240 1435
rect 1410 1405 1440 1435
rect 1610 1405 1640 1435
rect 1810 1405 1840 1435
rect 2010 1405 2040 1435
rect 2210 1405 2240 1435
rect 2410 1405 2440 1435
rect 2610 1405 2640 1435
rect 2810 1405 2840 1435
rect 3010 1405 3040 1435
rect 3210 1405 3240 1435
rect 3410 1405 3440 1435
rect 3610 1405 3640 1435
rect 3810 1405 3840 1435
rect 4010 1405 4040 1435
rect 4210 1405 4240 1435
rect 4410 1405 4440 1435
rect 4610 1405 4640 1435
rect 4810 1405 4840 1435
rect 5010 1405 5040 1435
rect 5210 1405 5240 1435
rect 5410 1405 5440 1435
rect 5610 1405 5640 1435
rect 5810 1405 5840 1435
rect 6010 1405 6040 1435
rect 6210 1405 6240 1435
rect 6410 1405 6440 1435
rect -190 1335 -185 1365
rect -185 1335 -165 1365
rect -165 1335 -160 1365
rect 10 1335 40 1365
rect 210 1335 240 1365
rect 410 1335 440 1365
rect 610 1335 640 1365
rect 810 1335 840 1365
rect 1010 1335 1040 1365
rect 1210 1335 1240 1365
rect 1410 1335 1440 1365
rect 1610 1335 1640 1365
rect 1810 1335 1840 1365
rect 2010 1335 2040 1365
rect 2210 1335 2240 1365
rect 2410 1335 2440 1365
rect 2610 1335 2640 1365
rect 2810 1335 2840 1365
rect 3010 1335 3040 1365
rect 3210 1335 3240 1365
rect 3410 1335 3440 1365
rect 3610 1335 3640 1365
rect 3810 1335 3840 1365
rect 4010 1335 4040 1365
rect 4210 1335 4240 1365
rect 4410 1335 4440 1365
rect 4610 1335 4640 1365
rect 4810 1335 4840 1365
rect 5010 1335 5040 1365
rect 5210 1335 5240 1365
rect 5410 1335 5440 1365
rect 5610 1335 5640 1365
rect 5810 1335 5840 1365
rect 6010 1335 6040 1365
rect 6210 1335 6240 1365
rect 6410 1335 6440 1365
rect -190 1220 -185 1250
rect -185 1220 -165 1250
rect -165 1220 -160 1250
rect 10 1220 40 1250
rect 210 1220 240 1250
rect 410 1220 440 1250
rect 610 1220 640 1250
rect 810 1220 840 1250
rect 1010 1220 1040 1250
rect 1210 1220 1240 1250
rect 1410 1220 1440 1250
rect 1610 1220 1640 1250
rect 1810 1220 1840 1250
rect 2010 1220 2040 1250
rect 2210 1220 2240 1250
rect 2410 1220 2440 1250
rect 2610 1220 2640 1250
rect 2810 1220 2840 1250
rect 3010 1220 3040 1250
rect 3210 1220 3240 1250
rect 3410 1220 3440 1250
rect 3610 1220 3640 1250
rect 3810 1220 3840 1250
rect 4010 1220 4040 1250
rect 4210 1220 4240 1250
rect 4410 1220 4440 1250
rect 4610 1220 4640 1250
rect 4810 1220 4840 1250
rect 5010 1220 5040 1250
rect 5210 1220 5240 1250
rect 5410 1220 5440 1250
rect 5610 1220 5640 1250
rect 5810 1220 5840 1250
rect 6010 1220 6040 1250
rect 6210 1220 6240 1250
rect 6410 1220 6440 1250
rect -190 1150 -185 1180
rect -185 1150 -165 1180
rect -165 1150 -160 1180
rect 10 1150 40 1180
rect 210 1150 240 1180
rect 410 1150 440 1180
rect 610 1150 640 1180
rect 810 1150 840 1180
rect 1010 1150 1040 1180
rect 1210 1150 1240 1180
rect 1410 1150 1440 1180
rect 1610 1150 1640 1180
rect 1810 1150 1840 1180
rect 2010 1150 2040 1180
rect 2210 1150 2240 1180
rect 2410 1150 2440 1180
rect 2610 1150 2640 1180
rect 2810 1150 2840 1180
rect 3010 1150 3040 1180
rect 3210 1150 3240 1180
rect 3410 1150 3440 1180
rect 3610 1150 3640 1180
rect 3810 1150 3840 1180
rect 4010 1150 4040 1180
rect 4210 1150 4240 1180
rect 4410 1150 4440 1180
rect 4610 1150 4640 1180
rect 4810 1150 4840 1180
rect 5010 1150 5040 1180
rect 5210 1150 5240 1180
rect 5410 1150 5440 1180
rect 5610 1150 5640 1180
rect 5810 1150 5840 1180
rect 6010 1150 6040 1180
rect 6210 1150 6240 1180
rect 6410 1150 6440 1180
rect -190 1035 -185 1065
rect -185 1035 -165 1065
rect -165 1035 -160 1065
rect 10 1035 40 1065
rect 210 1035 240 1065
rect 410 1035 440 1065
rect 610 1035 640 1065
rect 810 1035 840 1065
rect 1010 1035 1040 1065
rect 1210 1035 1240 1065
rect 1410 1035 1440 1065
rect 1610 1035 1640 1065
rect 1810 1035 1840 1065
rect 2010 1035 2040 1065
rect 2210 1035 2240 1065
rect 2410 1035 2440 1065
rect 2610 1035 2640 1065
rect 2810 1035 2840 1065
rect 3010 1035 3040 1065
rect 3210 1035 3240 1065
rect 3410 1035 3440 1065
rect 3610 1035 3640 1065
rect 3810 1035 3840 1065
rect 4010 1035 4040 1065
rect 4210 1035 4240 1065
rect 4410 1035 4440 1065
rect 4610 1035 4640 1065
rect 4810 1035 4840 1065
rect 5010 1035 5040 1065
rect 5210 1035 5240 1065
rect 5410 1035 5440 1065
rect 5610 1035 5640 1065
rect 5810 1035 5840 1065
rect 6010 1035 6040 1065
rect 6210 1035 6240 1065
rect 6410 1035 6440 1065
rect -190 965 -185 995
rect -185 965 -165 995
rect -165 965 -160 995
rect 10 965 40 995
rect 210 965 240 995
rect 410 965 440 995
rect 610 965 640 995
rect 810 965 840 995
rect 1010 965 1040 995
rect 1210 965 1240 995
rect 1410 965 1440 995
rect 1610 965 1640 995
rect 1810 965 1840 995
rect 2010 965 2040 995
rect 2210 965 2240 995
rect 2410 965 2440 995
rect 2610 965 2640 995
rect 2810 965 2840 995
rect 3010 965 3040 995
rect 3210 965 3240 995
rect 3410 965 3440 995
rect 3610 965 3640 995
rect 3810 965 3840 995
rect 4010 965 4040 995
rect 4210 965 4240 995
rect 4410 965 4440 995
rect 4610 965 4640 995
rect 4810 965 4840 995
rect 5010 965 5040 995
rect 5210 965 5240 995
rect 5410 965 5440 995
rect 5610 965 5640 995
rect 5810 965 5840 995
rect 6010 965 6040 995
rect 6210 965 6240 995
rect 6410 965 6440 995
rect -190 850 -185 880
rect -185 850 -165 880
rect -165 850 -160 880
rect 10 850 40 880
rect 210 850 240 880
rect 410 850 440 880
rect 610 850 640 880
rect 810 850 840 880
rect 1010 850 1040 880
rect 1210 850 1240 880
rect 1410 850 1440 880
rect 1610 850 1640 880
rect 1810 850 1840 880
rect 2010 850 2040 880
rect 2210 850 2240 880
rect 2410 850 2440 880
rect 2610 850 2640 880
rect 2810 850 2840 880
rect 3010 850 3040 880
rect 3210 850 3240 880
rect 3410 850 3440 880
rect 3610 850 3640 880
rect 3810 850 3840 880
rect 4010 850 4040 880
rect 4210 850 4240 880
rect 4410 850 4440 880
rect 4610 850 4640 880
rect 4810 850 4840 880
rect 5010 850 5040 880
rect 5210 850 5240 880
rect 5410 850 5440 880
rect 5610 850 5640 880
rect 5810 850 5840 880
rect 6010 850 6040 880
rect 6210 850 6240 880
rect 6410 850 6440 880
rect -190 780 -185 810
rect -185 780 -165 810
rect -165 780 -160 810
rect 10 780 40 810
rect 210 780 240 810
rect 410 780 440 810
rect 610 780 640 810
rect 810 780 840 810
rect 1010 780 1040 810
rect 1210 780 1240 810
rect 1410 780 1440 810
rect 1610 780 1640 810
rect 1810 780 1840 810
rect 2010 780 2040 810
rect 2210 780 2240 810
rect 2410 780 2440 810
rect 2610 780 2640 810
rect 2810 780 2840 810
rect 3010 780 3040 810
rect 3210 780 3240 810
rect 3410 780 3440 810
rect 3610 780 3640 810
rect 3810 780 3840 810
rect 4010 780 4040 810
rect 4210 780 4240 810
rect 4410 780 4440 810
rect 4610 780 4640 810
rect 4810 780 4840 810
rect 5010 780 5040 810
rect 5210 780 5240 810
rect 5410 780 5440 810
rect 5610 780 5640 810
rect 5810 780 5840 810
rect 6010 780 6040 810
rect 6210 780 6240 810
rect 6410 780 6440 810
rect -190 665 -185 695
rect -185 665 -165 695
rect -165 665 -160 695
rect 10 665 40 695
rect 210 665 240 695
rect 410 665 440 695
rect 610 665 640 695
rect 810 665 840 695
rect 1010 665 1040 695
rect 1210 665 1240 695
rect 1410 665 1440 695
rect 1610 665 1640 695
rect 1810 665 1840 695
rect 2010 665 2040 695
rect 2210 665 2240 695
rect 2410 665 2440 695
rect 2610 665 2640 695
rect 2810 665 2840 695
rect 3010 665 3040 695
rect 3210 665 3240 695
rect 3410 665 3440 695
rect 3610 665 3640 695
rect 3810 665 3840 695
rect 4010 665 4040 695
rect 4210 665 4240 695
rect 4410 665 4440 695
rect 4610 665 4640 695
rect 4810 665 4840 695
rect 5010 665 5040 695
rect 5210 665 5240 695
rect 5410 665 5440 695
rect 5610 665 5640 695
rect 5810 665 5840 695
rect 6010 665 6040 695
rect 6210 665 6240 695
rect 6410 665 6440 695
rect -190 595 -185 625
rect -185 595 -165 625
rect -165 595 -160 625
rect 10 595 40 625
rect 210 595 240 625
rect 410 595 440 625
rect 610 595 640 625
rect 810 595 840 625
rect 1010 595 1040 625
rect 1210 595 1240 625
rect 1410 595 1440 625
rect 1610 595 1640 625
rect 1810 595 1840 625
rect 2010 595 2040 625
rect 2210 595 2240 625
rect 2410 595 2440 625
rect 2610 595 2640 625
rect 2810 595 2840 625
rect 3010 595 3040 625
rect 3210 595 3240 625
rect 3410 595 3440 625
rect 3610 595 3640 625
rect 3810 595 3840 625
rect 4010 595 4040 625
rect 4210 595 4240 625
rect 4410 595 4440 625
rect 4610 595 4640 625
rect 4810 595 4840 625
rect 5010 595 5040 625
rect 5210 595 5240 625
rect 5410 595 5440 625
rect 5610 595 5640 625
rect 5810 595 5840 625
rect 6010 595 6040 625
rect 6210 595 6240 625
rect 6410 595 6440 625
rect -190 480 -185 510
rect -185 480 -165 510
rect -165 480 -160 510
rect 10 480 40 510
rect 210 480 240 510
rect 410 480 440 510
rect 610 480 640 510
rect 810 480 840 510
rect 1010 480 1040 510
rect 1210 480 1240 510
rect 1410 480 1440 510
rect 1610 480 1640 510
rect 1810 480 1840 510
rect 2010 480 2040 510
rect 2210 480 2240 510
rect 2410 480 2440 510
rect 2610 480 2640 510
rect 2810 480 2840 510
rect 3010 480 3040 510
rect 3210 480 3240 510
rect 3410 480 3440 510
rect 3610 480 3640 510
rect 3810 480 3840 510
rect 4010 480 4040 510
rect 4210 480 4240 510
rect 4410 480 4440 510
rect 4610 480 4640 510
rect 4810 480 4840 510
rect 5010 480 5040 510
rect 5210 480 5240 510
rect 5410 480 5440 510
rect 5610 480 5640 510
rect 5810 480 5840 510
rect 6010 480 6040 510
rect 6210 480 6240 510
rect 6410 480 6440 510
rect -190 410 -185 440
rect -185 410 -165 440
rect -165 410 -160 440
rect 10 410 40 440
rect 210 410 240 440
rect 410 410 440 440
rect 610 410 640 440
rect 810 410 840 440
rect 1010 410 1040 440
rect 1210 410 1240 440
rect 1410 410 1440 440
rect 1610 410 1640 440
rect 1810 410 1840 440
rect 2010 410 2040 440
rect 2210 410 2240 440
rect 2410 410 2440 440
rect 2610 410 2640 440
rect 2810 410 2840 440
rect 3010 410 3040 440
rect 3210 410 3240 440
rect 3410 410 3440 440
rect 3610 410 3640 440
rect 3810 410 3840 440
rect 4010 410 4040 440
rect 4210 410 4240 440
rect 4410 410 4440 440
rect 4610 410 4640 440
rect 4810 410 4840 440
rect 5010 410 5040 440
rect 5210 410 5240 440
rect 5410 410 5440 440
rect 5610 410 5640 440
rect 5810 410 5840 440
rect 6010 410 6040 440
rect 6210 410 6240 440
rect 6410 410 6440 440
rect -190 295 -185 325
rect -185 295 -165 325
rect -165 295 -160 325
rect 10 295 40 325
rect 210 295 240 325
rect 410 295 440 325
rect 610 295 640 325
rect 810 295 840 325
rect 1010 295 1040 325
rect 1210 295 1240 325
rect 1410 295 1440 325
rect 1610 295 1640 325
rect 1810 295 1840 325
rect 2010 295 2040 325
rect 2210 295 2240 325
rect 2410 295 2440 325
rect 2610 295 2640 325
rect 2810 295 2840 325
rect 3010 295 3040 325
rect 3210 295 3240 325
rect 3410 295 3440 325
rect 3610 295 3640 325
rect 3810 295 3840 325
rect 4010 295 4040 325
rect 4210 295 4240 325
rect 4410 295 4440 325
rect 4610 295 4640 325
rect 4810 295 4840 325
rect 5010 295 5040 325
rect 5210 295 5240 325
rect 5410 295 5440 325
rect 5610 295 5640 325
rect 5810 295 5840 325
rect 6010 295 6040 325
rect 6210 295 6240 325
rect 6410 295 6440 325
rect -190 225 -185 255
rect -185 225 -165 255
rect -165 225 -160 255
rect 10 225 40 255
rect 210 225 240 255
rect 410 225 440 255
rect 610 225 640 255
rect 810 225 840 255
rect 1010 225 1040 255
rect 1210 225 1240 255
rect 1410 225 1440 255
rect 1610 225 1640 255
rect 1810 225 1840 255
rect 2010 225 2040 255
rect 2210 225 2240 255
rect 2410 225 2440 255
rect 2610 225 2640 255
rect 2810 225 2840 255
rect 3010 225 3040 255
rect 3210 225 3240 255
rect 3410 225 3440 255
rect 3610 225 3640 255
rect 3810 225 3840 255
rect 4010 225 4040 255
rect 4210 225 4240 255
rect 4410 225 4440 255
rect 4610 225 4640 255
rect 4810 225 4840 255
rect 5010 225 5040 255
rect 5210 225 5240 255
rect 5410 225 5440 255
rect 5610 225 5640 255
rect 5810 225 5840 255
rect 6010 225 6040 255
rect 6210 225 6240 255
rect 6410 225 6440 255
rect -190 110 -185 140
rect -185 110 -165 140
rect -165 110 -160 140
rect 10 110 40 140
rect 210 110 240 140
rect 410 110 440 140
rect 610 110 640 140
rect 810 110 840 140
rect 1010 110 1040 140
rect 1210 110 1240 140
rect 1410 110 1440 140
rect 1610 110 1640 140
rect 1810 110 1840 140
rect 2010 110 2040 140
rect 2210 110 2240 140
rect 2410 110 2440 140
rect 2610 110 2640 140
rect 2810 110 2840 140
rect 3010 110 3040 140
rect 3210 110 3240 140
rect 3410 110 3440 140
rect 3610 110 3640 140
rect 3810 110 3840 140
rect 4010 110 4040 140
rect 4210 110 4240 140
rect 4410 110 4440 140
rect 4610 110 4640 140
rect 4810 110 4840 140
rect 5010 110 5040 140
rect 5210 110 5240 140
rect 5410 110 5440 140
rect 5610 110 5640 140
rect 5810 110 5840 140
rect 6010 110 6040 140
rect 6210 110 6240 140
rect 6410 110 6440 140
rect -190 40 -185 70
rect -185 40 -165 70
rect -165 40 -160 70
rect 10 40 40 70
rect 210 40 240 70
rect 410 40 440 70
rect 610 40 640 70
rect 810 40 840 70
rect 1010 40 1040 70
rect 1210 40 1240 70
rect 1410 40 1440 70
rect 1610 40 1640 70
rect 1810 40 1840 70
rect 2010 40 2040 70
rect 2210 40 2240 70
rect 2410 40 2440 70
rect 2610 40 2640 70
rect 2810 40 2840 70
rect 3010 40 3040 70
rect 3210 40 3240 70
rect 3410 40 3440 70
rect 3610 40 3640 70
rect 3810 40 3840 70
rect 4010 40 4040 70
rect 4210 40 4240 70
rect 4410 40 4440 70
rect 4610 40 4640 70
rect 4810 40 4840 70
rect 5010 40 5040 70
rect 5210 40 5240 70
rect 5410 40 5440 70
rect 5610 40 5640 70
rect 5810 40 5840 70
rect 6010 40 6040 70
rect 6210 40 6240 70
rect 6410 40 6440 70
rect -190 -75 -160 -45
rect 10 -75 40 -45
rect 210 -75 240 -45
rect 410 -75 440 -45
rect 610 -75 640 -45
rect 810 -75 840 -45
rect 1010 -75 1040 -45
rect 1210 -75 1240 -45
rect 1410 -75 1440 -45
rect 1610 -75 1640 -45
rect 1810 -75 1840 -45
rect 2010 -75 2040 -45
rect 2210 -75 2240 -45
rect 2410 -75 2440 -45
rect 2610 -75 2640 -45
rect 2810 -75 2840 -45
rect 3010 -75 3040 -45
rect 3210 -75 3240 -45
rect 3410 -75 3440 -45
rect 3610 -75 3640 -45
rect 3810 -75 3840 -45
rect 4010 -75 4040 -45
rect 4210 -75 4240 -45
rect 4410 -75 4440 -45
rect 4610 -75 4640 -45
rect 4810 -75 4840 -45
rect 5010 -75 5040 -45
rect 5210 -75 5240 -45
rect 5410 -75 5440 -45
rect 5610 -75 5640 -45
rect 5810 -75 5840 -45
rect 6010 -75 6040 -45
rect 6210 -75 6240 -45
rect 6410 -75 6440 -45
rect -190 -145 -160 -115
rect 10 -145 40 -115
rect 210 -145 240 -115
rect 410 -145 440 -115
rect 610 -145 640 -115
rect 810 -145 840 -115
rect 1010 -145 1040 -115
rect 1210 -145 1240 -115
rect 1410 -145 1440 -115
rect 1610 -145 1640 -115
rect 1810 -145 1840 -115
rect 2010 -145 2040 -115
rect 2210 -145 2240 -115
rect 2410 -145 2440 -115
rect 2610 -145 2640 -115
rect 2810 -145 2840 -115
rect 3010 -145 3040 -115
rect 3210 -145 3240 -115
rect 3410 -145 3440 -115
rect 3610 -145 3640 -115
rect 3810 -145 3840 -115
rect 4010 -145 4040 -115
rect 4210 -145 4240 -115
rect 4410 -145 4440 -115
rect 4610 -145 4640 -115
rect 4810 -145 4840 -115
rect 5010 -145 5040 -115
rect 5210 -145 5240 -115
rect 5410 -145 5440 -115
rect 5610 -145 5640 -115
rect 5810 -145 5840 -115
rect 6010 -145 6040 -115
rect 6210 -145 6240 -115
rect 6410 -145 6440 -115
<< metal2 >>
rect -145 12090 -55 12095
rect -145 12060 -140 12090
rect -110 12060 -90 12090
rect -60 12060 -55 12090
rect -145 12055 -55 12060
rect 6455 12065 6545 12070
rect 6455 12035 6460 12065
rect 6490 12035 6510 12065
rect 6540 12035 6545 12065
rect 6455 12030 6545 12035
rect -195 11980 -155 11985
rect -195 11950 -190 11980
rect -160 11950 -155 11980
rect -195 11910 -155 11950
rect -195 11880 -190 11910
rect -160 11880 -155 11910
rect -195 11875 -155 11880
rect 5 11980 45 11985
rect 5 11950 10 11980
rect 40 11950 45 11980
rect 5 11910 45 11950
rect 5 11880 10 11910
rect 40 11880 45 11910
rect 5 11875 45 11880
rect 205 11980 245 11985
rect 205 11950 210 11980
rect 240 11950 245 11980
rect 205 11910 245 11950
rect 205 11880 210 11910
rect 240 11880 245 11910
rect 205 11875 245 11880
rect 405 11980 445 11985
rect 405 11950 410 11980
rect 440 11950 445 11980
rect 405 11910 445 11950
rect 405 11880 410 11910
rect 440 11880 445 11910
rect 405 11875 445 11880
rect 605 11980 645 11985
rect 605 11950 610 11980
rect 640 11950 645 11980
rect 605 11910 645 11950
rect 605 11880 610 11910
rect 640 11880 645 11910
rect 605 11875 645 11880
rect 805 11980 845 11985
rect 805 11950 810 11980
rect 840 11950 845 11980
rect 805 11910 845 11950
rect 805 11880 810 11910
rect 840 11880 845 11910
rect 805 11875 845 11880
rect 1005 11980 1045 11985
rect 1005 11950 1010 11980
rect 1040 11950 1045 11980
rect 1005 11910 1045 11950
rect 1005 11880 1010 11910
rect 1040 11880 1045 11910
rect 1005 11875 1045 11880
rect 1205 11980 1245 11985
rect 1205 11950 1210 11980
rect 1240 11950 1245 11980
rect 1205 11910 1245 11950
rect 1205 11880 1210 11910
rect 1240 11880 1245 11910
rect 1205 11875 1245 11880
rect 1405 11980 1445 11985
rect 1405 11950 1410 11980
rect 1440 11950 1445 11980
rect 1405 11910 1445 11950
rect 1405 11880 1410 11910
rect 1440 11880 1445 11910
rect 1405 11875 1445 11880
rect 1605 11980 1645 11985
rect 1605 11950 1610 11980
rect 1640 11950 1645 11980
rect 1605 11910 1645 11950
rect 1605 11880 1610 11910
rect 1640 11880 1645 11910
rect 1605 11875 1645 11880
rect 1805 11980 1845 11985
rect 1805 11950 1810 11980
rect 1840 11950 1845 11980
rect 1805 11910 1845 11950
rect 1805 11880 1810 11910
rect 1840 11880 1845 11910
rect 1805 11875 1845 11880
rect 2005 11980 2045 11985
rect 2005 11950 2010 11980
rect 2040 11950 2045 11980
rect 2005 11910 2045 11950
rect 2005 11880 2010 11910
rect 2040 11880 2045 11910
rect 2005 11875 2045 11880
rect 2205 11980 2245 11985
rect 2205 11950 2210 11980
rect 2240 11950 2245 11980
rect 2205 11910 2245 11950
rect 2205 11880 2210 11910
rect 2240 11880 2245 11910
rect 2205 11875 2245 11880
rect 2405 11980 2445 11985
rect 2405 11950 2410 11980
rect 2440 11950 2445 11980
rect 2405 11910 2445 11950
rect 2405 11880 2410 11910
rect 2440 11880 2445 11910
rect 2405 11875 2445 11880
rect 2605 11980 2645 11985
rect 2605 11950 2610 11980
rect 2640 11950 2645 11980
rect 2605 11910 2645 11950
rect 2605 11880 2610 11910
rect 2640 11880 2645 11910
rect 2605 11875 2645 11880
rect 2805 11980 2845 11985
rect 2805 11950 2810 11980
rect 2840 11950 2845 11980
rect 2805 11910 2845 11950
rect 2805 11880 2810 11910
rect 2840 11880 2845 11910
rect 2805 11875 2845 11880
rect 3005 11980 3045 11985
rect 3005 11950 3010 11980
rect 3040 11950 3045 11980
rect 3005 11910 3045 11950
rect 3005 11880 3010 11910
rect 3040 11880 3045 11910
rect 3005 11875 3045 11880
rect 3205 11980 3245 11985
rect 3205 11950 3210 11980
rect 3240 11950 3245 11980
rect 3205 11910 3245 11950
rect 3205 11880 3210 11910
rect 3240 11880 3245 11910
rect 3205 11875 3245 11880
rect 3405 11980 3445 11985
rect 3405 11950 3410 11980
rect 3440 11950 3445 11980
rect 3405 11910 3445 11950
rect 3405 11880 3410 11910
rect 3440 11880 3445 11910
rect 3405 11875 3445 11880
rect 3605 11980 3645 11985
rect 3605 11950 3610 11980
rect 3640 11950 3645 11980
rect 3605 11910 3645 11950
rect 3605 11880 3610 11910
rect 3640 11880 3645 11910
rect 3605 11875 3645 11880
rect 3805 11980 3845 11985
rect 3805 11950 3810 11980
rect 3840 11950 3845 11980
rect 3805 11910 3845 11950
rect 3805 11880 3810 11910
rect 3840 11880 3845 11910
rect 3805 11875 3845 11880
rect 4005 11980 4045 11985
rect 4005 11950 4010 11980
rect 4040 11950 4045 11980
rect 4005 11910 4045 11950
rect 4005 11880 4010 11910
rect 4040 11880 4045 11910
rect 4005 11875 4045 11880
rect 4205 11980 4245 11985
rect 4205 11950 4210 11980
rect 4240 11950 4245 11980
rect 4205 11910 4245 11950
rect 4205 11880 4210 11910
rect 4240 11880 4245 11910
rect 4205 11875 4245 11880
rect 4405 11980 4445 11985
rect 4405 11950 4410 11980
rect 4440 11950 4445 11980
rect 4405 11910 4445 11950
rect 4405 11880 4410 11910
rect 4440 11880 4445 11910
rect 4405 11875 4445 11880
rect 4605 11980 4645 11985
rect 4605 11950 4610 11980
rect 4640 11950 4645 11980
rect 4605 11910 4645 11950
rect 4605 11880 4610 11910
rect 4640 11880 4645 11910
rect 4605 11875 4645 11880
rect 4805 11980 4845 11985
rect 4805 11950 4810 11980
rect 4840 11950 4845 11980
rect 4805 11910 4845 11950
rect 4805 11880 4810 11910
rect 4840 11880 4845 11910
rect 4805 11875 4845 11880
rect 5005 11980 5045 11985
rect 5005 11950 5010 11980
rect 5040 11950 5045 11980
rect 5005 11910 5045 11950
rect 5005 11880 5010 11910
rect 5040 11880 5045 11910
rect 5005 11875 5045 11880
rect 5205 11980 5245 11985
rect 5205 11950 5210 11980
rect 5240 11950 5245 11980
rect 5205 11910 5245 11950
rect 5205 11880 5210 11910
rect 5240 11880 5245 11910
rect 5205 11875 5245 11880
rect 5405 11980 5445 11985
rect 5405 11950 5410 11980
rect 5440 11950 5445 11980
rect 5405 11910 5445 11950
rect 5405 11880 5410 11910
rect 5440 11880 5445 11910
rect 5405 11875 5445 11880
rect 5605 11980 5645 11985
rect 5605 11950 5610 11980
rect 5640 11950 5645 11980
rect 5605 11910 5645 11950
rect 5605 11880 5610 11910
rect 5640 11880 5645 11910
rect 5605 11875 5645 11880
rect 5805 11980 5845 11985
rect 5805 11950 5810 11980
rect 5840 11950 5845 11980
rect 5805 11910 5845 11950
rect 5805 11880 5810 11910
rect 5840 11880 5845 11910
rect 5805 11875 5845 11880
rect 6005 11980 6045 11985
rect 6005 11950 6010 11980
rect 6040 11950 6045 11980
rect 6005 11910 6045 11950
rect 6005 11880 6010 11910
rect 6040 11880 6045 11910
rect 6005 11875 6045 11880
rect 6205 11980 6245 11985
rect 6205 11950 6210 11980
rect 6240 11950 6245 11980
rect 6205 11910 6245 11950
rect 6205 11880 6210 11910
rect 6240 11880 6245 11910
rect 6205 11875 6245 11880
rect 6405 11980 6445 11985
rect 6405 11950 6410 11980
rect 6440 11950 6445 11980
rect 6405 11910 6445 11950
rect 6405 11880 6410 11910
rect 6440 11880 6445 11910
rect 6405 11875 6445 11880
rect -195 11795 -155 11800
rect -195 11765 -190 11795
rect -160 11765 -155 11795
rect -195 11725 -155 11765
rect -195 11695 -190 11725
rect -160 11695 -155 11725
rect -195 11690 -155 11695
rect 5 11795 45 11800
rect 5 11765 10 11795
rect 40 11765 45 11795
rect 5 11725 45 11765
rect 5 11695 10 11725
rect 40 11695 45 11725
rect 5 11690 45 11695
rect 205 11795 245 11800
rect 205 11765 210 11795
rect 240 11765 245 11795
rect 205 11725 245 11765
rect 205 11695 210 11725
rect 240 11695 245 11725
rect 205 11690 245 11695
rect 405 11795 445 11800
rect 405 11765 410 11795
rect 440 11765 445 11795
rect 405 11725 445 11765
rect 405 11695 410 11725
rect 440 11695 445 11725
rect 405 11690 445 11695
rect 605 11795 645 11800
rect 605 11765 610 11795
rect 640 11765 645 11795
rect 605 11725 645 11765
rect 605 11695 610 11725
rect 640 11695 645 11725
rect 605 11690 645 11695
rect 805 11795 845 11800
rect 805 11765 810 11795
rect 840 11765 845 11795
rect 805 11725 845 11765
rect 805 11695 810 11725
rect 840 11695 845 11725
rect 805 11690 845 11695
rect 1005 11795 1045 11800
rect 1005 11765 1010 11795
rect 1040 11765 1045 11795
rect 1005 11725 1045 11765
rect 1005 11695 1010 11725
rect 1040 11695 1045 11725
rect 1005 11690 1045 11695
rect 1205 11795 1245 11800
rect 1205 11765 1210 11795
rect 1240 11765 1245 11795
rect 1205 11725 1245 11765
rect 1205 11695 1210 11725
rect 1240 11695 1245 11725
rect 1205 11690 1245 11695
rect 1405 11795 1445 11800
rect 1405 11765 1410 11795
rect 1440 11765 1445 11795
rect 1405 11725 1445 11765
rect 1405 11695 1410 11725
rect 1440 11695 1445 11725
rect 1405 11690 1445 11695
rect 1605 11795 1645 11800
rect 1605 11765 1610 11795
rect 1640 11765 1645 11795
rect 1605 11725 1645 11765
rect 1605 11695 1610 11725
rect 1640 11695 1645 11725
rect 1605 11690 1645 11695
rect 1805 11795 1845 11800
rect 1805 11765 1810 11795
rect 1840 11765 1845 11795
rect 1805 11725 1845 11765
rect 1805 11695 1810 11725
rect 1840 11695 1845 11725
rect 1805 11690 1845 11695
rect 2005 11795 2045 11800
rect 2005 11765 2010 11795
rect 2040 11765 2045 11795
rect 2005 11725 2045 11765
rect 2005 11695 2010 11725
rect 2040 11695 2045 11725
rect 2005 11690 2045 11695
rect 2205 11795 2245 11800
rect 2205 11765 2210 11795
rect 2240 11765 2245 11795
rect 2205 11725 2245 11765
rect 2205 11695 2210 11725
rect 2240 11695 2245 11725
rect 2205 11690 2245 11695
rect 2405 11795 2445 11800
rect 2405 11765 2410 11795
rect 2440 11765 2445 11795
rect 2405 11725 2445 11765
rect 2405 11695 2410 11725
rect 2440 11695 2445 11725
rect 2405 11690 2445 11695
rect 2605 11795 2645 11800
rect 2605 11765 2610 11795
rect 2640 11765 2645 11795
rect 2605 11725 2645 11765
rect 2605 11695 2610 11725
rect 2640 11695 2645 11725
rect 2605 11690 2645 11695
rect 2805 11795 2845 11800
rect 2805 11765 2810 11795
rect 2840 11765 2845 11795
rect 2805 11725 2845 11765
rect 2805 11695 2810 11725
rect 2840 11695 2845 11725
rect 2805 11690 2845 11695
rect 3005 11795 3045 11800
rect 3005 11765 3010 11795
rect 3040 11765 3045 11795
rect 3005 11725 3045 11765
rect 3005 11695 3010 11725
rect 3040 11695 3045 11725
rect 3005 11690 3045 11695
rect 3205 11795 3245 11800
rect 3205 11765 3210 11795
rect 3240 11765 3245 11795
rect 3205 11725 3245 11765
rect 3205 11695 3210 11725
rect 3240 11695 3245 11725
rect 3205 11690 3245 11695
rect 3405 11795 3445 11800
rect 3405 11765 3410 11795
rect 3440 11765 3445 11795
rect 3405 11725 3445 11765
rect 3405 11695 3410 11725
rect 3440 11695 3445 11725
rect 3405 11690 3445 11695
rect 3605 11795 3645 11800
rect 3605 11765 3610 11795
rect 3640 11765 3645 11795
rect 3605 11725 3645 11765
rect 3605 11695 3610 11725
rect 3640 11695 3645 11725
rect 3605 11690 3645 11695
rect 3805 11795 3845 11800
rect 3805 11765 3810 11795
rect 3840 11765 3845 11795
rect 3805 11725 3845 11765
rect 3805 11695 3810 11725
rect 3840 11695 3845 11725
rect 3805 11690 3845 11695
rect 4005 11795 4045 11800
rect 4005 11765 4010 11795
rect 4040 11765 4045 11795
rect 4005 11725 4045 11765
rect 4005 11695 4010 11725
rect 4040 11695 4045 11725
rect 4005 11690 4045 11695
rect 4205 11795 4245 11800
rect 4205 11765 4210 11795
rect 4240 11765 4245 11795
rect 4205 11725 4245 11765
rect 4205 11695 4210 11725
rect 4240 11695 4245 11725
rect 4205 11690 4245 11695
rect 4405 11795 4445 11800
rect 4405 11765 4410 11795
rect 4440 11765 4445 11795
rect 4405 11725 4445 11765
rect 4405 11695 4410 11725
rect 4440 11695 4445 11725
rect 4405 11690 4445 11695
rect 4605 11795 4645 11800
rect 4605 11765 4610 11795
rect 4640 11765 4645 11795
rect 4605 11725 4645 11765
rect 4605 11695 4610 11725
rect 4640 11695 4645 11725
rect 4605 11690 4645 11695
rect 4805 11795 4845 11800
rect 4805 11765 4810 11795
rect 4840 11765 4845 11795
rect 4805 11725 4845 11765
rect 4805 11695 4810 11725
rect 4840 11695 4845 11725
rect 4805 11690 4845 11695
rect 5005 11795 5045 11800
rect 5005 11765 5010 11795
rect 5040 11765 5045 11795
rect 5005 11725 5045 11765
rect 5005 11695 5010 11725
rect 5040 11695 5045 11725
rect 5005 11690 5045 11695
rect 5205 11795 5245 11800
rect 5205 11765 5210 11795
rect 5240 11765 5245 11795
rect 5205 11725 5245 11765
rect 5205 11695 5210 11725
rect 5240 11695 5245 11725
rect 5205 11690 5245 11695
rect 5405 11795 5445 11800
rect 5405 11765 5410 11795
rect 5440 11765 5445 11795
rect 5405 11725 5445 11765
rect 5405 11695 5410 11725
rect 5440 11695 5445 11725
rect 5405 11690 5445 11695
rect 5605 11795 5645 11800
rect 5605 11765 5610 11795
rect 5640 11765 5645 11795
rect 5605 11725 5645 11765
rect 5605 11695 5610 11725
rect 5640 11695 5645 11725
rect 5605 11690 5645 11695
rect 5805 11795 5845 11800
rect 5805 11765 5810 11795
rect 5840 11765 5845 11795
rect 5805 11725 5845 11765
rect 5805 11695 5810 11725
rect 5840 11695 5845 11725
rect 5805 11690 5845 11695
rect 6005 11795 6045 11800
rect 6005 11765 6010 11795
rect 6040 11765 6045 11795
rect 6005 11725 6045 11765
rect 6005 11695 6010 11725
rect 6040 11695 6045 11725
rect 6005 11690 6045 11695
rect 6205 11795 6245 11800
rect 6205 11765 6210 11795
rect 6240 11765 6245 11795
rect 6205 11725 6245 11765
rect 6205 11695 6210 11725
rect 6240 11695 6245 11725
rect 6205 11690 6245 11695
rect 6405 11795 6445 11800
rect 6405 11765 6410 11795
rect 6440 11765 6445 11795
rect 6405 11725 6445 11765
rect 6405 11695 6410 11725
rect 6440 11695 6445 11725
rect 6405 11690 6445 11695
rect -195 11610 -155 11615
rect -195 11580 -190 11610
rect -160 11580 -155 11610
rect -195 11540 -155 11580
rect -195 11510 -190 11540
rect -160 11510 -155 11540
rect -195 11505 -155 11510
rect 5 11610 45 11615
rect 5 11580 10 11610
rect 40 11580 45 11610
rect 5 11540 45 11580
rect 5 11510 10 11540
rect 40 11510 45 11540
rect 5 11505 45 11510
rect 205 11610 245 11615
rect 205 11580 210 11610
rect 240 11580 245 11610
rect 205 11540 245 11580
rect 205 11510 210 11540
rect 240 11510 245 11540
rect 205 11505 245 11510
rect 405 11610 445 11615
rect 405 11580 410 11610
rect 440 11580 445 11610
rect 405 11540 445 11580
rect 405 11510 410 11540
rect 440 11510 445 11540
rect 405 11505 445 11510
rect 605 11610 645 11615
rect 605 11580 610 11610
rect 640 11580 645 11610
rect 605 11540 645 11580
rect 605 11510 610 11540
rect 640 11510 645 11540
rect 605 11505 645 11510
rect 805 11610 845 11615
rect 805 11580 810 11610
rect 840 11580 845 11610
rect 805 11540 845 11580
rect 805 11510 810 11540
rect 840 11510 845 11540
rect 805 11505 845 11510
rect 1005 11610 1045 11615
rect 1005 11580 1010 11610
rect 1040 11580 1045 11610
rect 1005 11540 1045 11580
rect 1005 11510 1010 11540
rect 1040 11510 1045 11540
rect 1005 11505 1045 11510
rect 1205 11610 1245 11615
rect 1205 11580 1210 11610
rect 1240 11580 1245 11610
rect 1205 11540 1245 11580
rect 1205 11510 1210 11540
rect 1240 11510 1245 11540
rect 1205 11505 1245 11510
rect 1405 11610 1445 11615
rect 1405 11580 1410 11610
rect 1440 11580 1445 11610
rect 1405 11540 1445 11580
rect 1405 11510 1410 11540
rect 1440 11510 1445 11540
rect 1405 11505 1445 11510
rect 1605 11610 1645 11615
rect 1605 11580 1610 11610
rect 1640 11580 1645 11610
rect 1605 11540 1645 11580
rect 1605 11510 1610 11540
rect 1640 11510 1645 11540
rect 1605 11505 1645 11510
rect 1805 11610 1845 11615
rect 1805 11580 1810 11610
rect 1840 11580 1845 11610
rect 1805 11540 1845 11580
rect 1805 11510 1810 11540
rect 1840 11510 1845 11540
rect 1805 11505 1845 11510
rect 2005 11610 2045 11615
rect 2005 11580 2010 11610
rect 2040 11580 2045 11610
rect 2005 11540 2045 11580
rect 2005 11510 2010 11540
rect 2040 11510 2045 11540
rect 2005 11505 2045 11510
rect 2205 11610 2245 11615
rect 2205 11580 2210 11610
rect 2240 11580 2245 11610
rect 2205 11540 2245 11580
rect 2205 11510 2210 11540
rect 2240 11510 2245 11540
rect 2205 11505 2245 11510
rect 2405 11610 2445 11615
rect 2405 11580 2410 11610
rect 2440 11580 2445 11610
rect 2405 11540 2445 11580
rect 2405 11510 2410 11540
rect 2440 11510 2445 11540
rect 2405 11505 2445 11510
rect 2605 11610 2645 11615
rect 2605 11580 2610 11610
rect 2640 11580 2645 11610
rect 2605 11540 2645 11580
rect 2605 11510 2610 11540
rect 2640 11510 2645 11540
rect 2605 11505 2645 11510
rect 2805 11610 2845 11615
rect 2805 11580 2810 11610
rect 2840 11580 2845 11610
rect 2805 11540 2845 11580
rect 2805 11510 2810 11540
rect 2840 11510 2845 11540
rect 2805 11505 2845 11510
rect 3005 11610 3045 11615
rect 3005 11580 3010 11610
rect 3040 11580 3045 11610
rect 3005 11540 3045 11580
rect 3005 11510 3010 11540
rect 3040 11510 3045 11540
rect 3005 11505 3045 11510
rect 3205 11610 3245 11615
rect 3205 11580 3210 11610
rect 3240 11580 3245 11610
rect 3205 11540 3245 11580
rect 3205 11510 3210 11540
rect 3240 11510 3245 11540
rect 3205 11505 3245 11510
rect 3405 11610 3445 11615
rect 3405 11580 3410 11610
rect 3440 11580 3445 11610
rect 3405 11540 3445 11580
rect 3405 11510 3410 11540
rect 3440 11510 3445 11540
rect 3405 11505 3445 11510
rect 3605 11610 3645 11615
rect 3605 11580 3610 11610
rect 3640 11580 3645 11610
rect 3605 11540 3645 11580
rect 3605 11510 3610 11540
rect 3640 11510 3645 11540
rect 3605 11505 3645 11510
rect 3805 11610 3845 11615
rect 3805 11580 3810 11610
rect 3840 11580 3845 11610
rect 3805 11540 3845 11580
rect 3805 11510 3810 11540
rect 3840 11510 3845 11540
rect 3805 11505 3845 11510
rect 4005 11610 4045 11615
rect 4005 11580 4010 11610
rect 4040 11580 4045 11610
rect 4005 11540 4045 11580
rect 4005 11510 4010 11540
rect 4040 11510 4045 11540
rect 4005 11505 4045 11510
rect 4205 11610 4245 11615
rect 4205 11580 4210 11610
rect 4240 11580 4245 11610
rect 4205 11540 4245 11580
rect 4205 11510 4210 11540
rect 4240 11510 4245 11540
rect 4205 11505 4245 11510
rect 4405 11610 4445 11615
rect 4405 11580 4410 11610
rect 4440 11580 4445 11610
rect 4405 11540 4445 11580
rect 4405 11510 4410 11540
rect 4440 11510 4445 11540
rect 4405 11505 4445 11510
rect 4605 11610 4645 11615
rect 4605 11580 4610 11610
rect 4640 11580 4645 11610
rect 4605 11540 4645 11580
rect 4605 11510 4610 11540
rect 4640 11510 4645 11540
rect 4605 11505 4645 11510
rect 4805 11610 4845 11615
rect 4805 11580 4810 11610
rect 4840 11580 4845 11610
rect 4805 11540 4845 11580
rect 4805 11510 4810 11540
rect 4840 11510 4845 11540
rect 4805 11505 4845 11510
rect 5005 11610 5045 11615
rect 5005 11580 5010 11610
rect 5040 11580 5045 11610
rect 5005 11540 5045 11580
rect 5005 11510 5010 11540
rect 5040 11510 5045 11540
rect 5005 11505 5045 11510
rect 5205 11610 5245 11615
rect 5205 11580 5210 11610
rect 5240 11580 5245 11610
rect 5205 11540 5245 11580
rect 5205 11510 5210 11540
rect 5240 11510 5245 11540
rect 5205 11505 5245 11510
rect 5405 11610 5445 11615
rect 5405 11580 5410 11610
rect 5440 11580 5445 11610
rect 5405 11540 5445 11580
rect 5405 11510 5410 11540
rect 5440 11510 5445 11540
rect 5405 11505 5445 11510
rect 5605 11610 5645 11615
rect 5605 11580 5610 11610
rect 5640 11580 5645 11610
rect 5605 11540 5645 11580
rect 5605 11510 5610 11540
rect 5640 11510 5645 11540
rect 5605 11505 5645 11510
rect 5805 11610 5845 11615
rect 5805 11580 5810 11610
rect 5840 11580 5845 11610
rect 5805 11540 5845 11580
rect 5805 11510 5810 11540
rect 5840 11510 5845 11540
rect 5805 11505 5845 11510
rect 6005 11610 6045 11615
rect 6005 11580 6010 11610
rect 6040 11580 6045 11610
rect 6005 11540 6045 11580
rect 6005 11510 6010 11540
rect 6040 11510 6045 11540
rect 6005 11505 6045 11510
rect 6205 11610 6245 11615
rect 6205 11580 6210 11610
rect 6240 11580 6245 11610
rect 6205 11540 6245 11580
rect 6205 11510 6210 11540
rect 6240 11510 6245 11540
rect 6205 11505 6245 11510
rect 6405 11610 6445 11615
rect 6405 11580 6410 11610
rect 6440 11580 6445 11610
rect 6405 11540 6445 11580
rect 6405 11510 6410 11540
rect 6440 11510 6445 11540
rect 6405 11505 6445 11510
rect -195 11425 -155 11430
rect -195 11395 -190 11425
rect -160 11395 -155 11425
rect -195 11355 -155 11395
rect -195 11325 -190 11355
rect -160 11325 -155 11355
rect -195 11320 -155 11325
rect 5 11425 45 11430
rect 5 11395 10 11425
rect 40 11395 45 11425
rect 5 11355 45 11395
rect 5 11325 10 11355
rect 40 11325 45 11355
rect 5 11320 45 11325
rect 205 11425 245 11430
rect 205 11395 210 11425
rect 240 11395 245 11425
rect 205 11355 245 11395
rect 205 11325 210 11355
rect 240 11325 245 11355
rect 205 11320 245 11325
rect 405 11425 445 11430
rect 405 11395 410 11425
rect 440 11395 445 11425
rect 405 11355 445 11395
rect 405 11325 410 11355
rect 440 11325 445 11355
rect 405 11320 445 11325
rect 605 11425 645 11430
rect 605 11395 610 11425
rect 640 11395 645 11425
rect 605 11355 645 11395
rect 605 11325 610 11355
rect 640 11325 645 11355
rect 605 11320 645 11325
rect 805 11425 845 11430
rect 805 11395 810 11425
rect 840 11395 845 11425
rect 805 11355 845 11395
rect 805 11325 810 11355
rect 840 11325 845 11355
rect 805 11320 845 11325
rect 1005 11425 1045 11430
rect 1005 11395 1010 11425
rect 1040 11395 1045 11425
rect 1005 11355 1045 11395
rect 1005 11325 1010 11355
rect 1040 11325 1045 11355
rect 1005 11320 1045 11325
rect 1205 11425 1245 11430
rect 1205 11395 1210 11425
rect 1240 11395 1245 11425
rect 1205 11355 1245 11395
rect 1205 11325 1210 11355
rect 1240 11325 1245 11355
rect 1205 11320 1245 11325
rect 1405 11425 1445 11430
rect 1405 11395 1410 11425
rect 1440 11395 1445 11425
rect 1405 11355 1445 11395
rect 1405 11325 1410 11355
rect 1440 11325 1445 11355
rect 1405 11320 1445 11325
rect 1605 11425 1645 11430
rect 1605 11395 1610 11425
rect 1640 11395 1645 11425
rect 1605 11355 1645 11395
rect 1605 11325 1610 11355
rect 1640 11325 1645 11355
rect 1605 11320 1645 11325
rect 1805 11425 1845 11430
rect 1805 11395 1810 11425
rect 1840 11395 1845 11425
rect 1805 11355 1845 11395
rect 1805 11325 1810 11355
rect 1840 11325 1845 11355
rect 1805 11320 1845 11325
rect 2005 11425 2045 11430
rect 2005 11395 2010 11425
rect 2040 11395 2045 11425
rect 2005 11355 2045 11395
rect 2005 11325 2010 11355
rect 2040 11325 2045 11355
rect 2005 11320 2045 11325
rect 2205 11425 2245 11430
rect 2205 11395 2210 11425
rect 2240 11395 2245 11425
rect 2205 11355 2245 11395
rect 2205 11325 2210 11355
rect 2240 11325 2245 11355
rect 2205 11320 2245 11325
rect 2405 11425 2445 11430
rect 2405 11395 2410 11425
rect 2440 11395 2445 11425
rect 2405 11355 2445 11395
rect 2405 11325 2410 11355
rect 2440 11325 2445 11355
rect 2405 11320 2445 11325
rect 2605 11425 2645 11430
rect 2605 11395 2610 11425
rect 2640 11395 2645 11425
rect 2605 11355 2645 11395
rect 2605 11325 2610 11355
rect 2640 11325 2645 11355
rect 2605 11320 2645 11325
rect 2805 11425 2845 11430
rect 2805 11395 2810 11425
rect 2840 11395 2845 11425
rect 2805 11355 2845 11395
rect 2805 11325 2810 11355
rect 2840 11325 2845 11355
rect 2805 11320 2845 11325
rect 3005 11425 3045 11430
rect 3005 11395 3010 11425
rect 3040 11395 3045 11425
rect 3005 11355 3045 11395
rect 3005 11325 3010 11355
rect 3040 11325 3045 11355
rect 3005 11320 3045 11325
rect 3205 11425 3245 11430
rect 3205 11395 3210 11425
rect 3240 11395 3245 11425
rect 3205 11355 3245 11395
rect 3205 11325 3210 11355
rect 3240 11325 3245 11355
rect 3205 11320 3245 11325
rect 3405 11425 3445 11430
rect 3405 11395 3410 11425
rect 3440 11395 3445 11425
rect 3405 11355 3445 11395
rect 3405 11325 3410 11355
rect 3440 11325 3445 11355
rect 3405 11320 3445 11325
rect 3605 11425 3645 11430
rect 3605 11395 3610 11425
rect 3640 11395 3645 11425
rect 3605 11355 3645 11395
rect 3605 11325 3610 11355
rect 3640 11325 3645 11355
rect 3605 11320 3645 11325
rect 3805 11425 3845 11430
rect 3805 11395 3810 11425
rect 3840 11395 3845 11425
rect 3805 11355 3845 11395
rect 3805 11325 3810 11355
rect 3840 11325 3845 11355
rect 3805 11320 3845 11325
rect 4005 11425 4045 11430
rect 4005 11395 4010 11425
rect 4040 11395 4045 11425
rect 4005 11355 4045 11395
rect 4005 11325 4010 11355
rect 4040 11325 4045 11355
rect 4005 11320 4045 11325
rect 4205 11425 4245 11430
rect 4205 11395 4210 11425
rect 4240 11395 4245 11425
rect 4205 11355 4245 11395
rect 4205 11325 4210 11355
rect 4240 11325 4245 11355
rect 4205 11320 4245 11325
rect 4405 11425 4445 11430
rect 4405 11395 4410 11425
rect 4440 11395 4445 11425
rect 4405 11355 4445 11395
rect 4405 11325 4410 11355
rect 4440 11325 4445 11355
rect 4405 11320 4445 11325
rect 4605 11425 4645 11430
rect 4605 11395 4610 11425
rect 4640 11395 4645 11425
rect 4605 11355 4645 11395
rect 4605 11325 4610 11355
rect 4640 11325 4645 11355
rect 4605 11320 4645 11325
rect 4805 11425 4845 11430
rect 4805 11395 4810 11425
rect 4840 11395 4845 11425
rect 4805 11355 4845 11395
rect 4805 11325 4810 11355
rect 4840 11325 4845 11355
rect 4805 11320 4845 11325
rect 5005 11425 5045 11430
rect 5005 11395 5010 11425
rect 5040 11395 5045 11425
rect 5005 11355 5045 11395
rect 5005 11325 5010 11355
rect 5040 11325 5045 11355
rect 5005 11320 5045 11325
rect 5205 11425 5245 11430
rect 5205 11395 5210 11425
rect 5240 11395 5245 11425
rect 5205 11355 5245 11395
rect 5205 11325 5210 11355
rect 5240 11325 5245 11355
rect 5205 11320 5245 11325
rect 5405 11425 5445 11430
rect 5405 11395 5410 11425
rect 5440 11395 5445 11425
rect 5405 11355 5445 11395
rect 5405 11325 5410 11355
rect 5440 11325 5445 11355
rect 5405 11320 5445 11325
rect 5605 11425 5645 11430
rect 5605 11395 5610 11425
rect 5640 11395 5645 11425
rect 5605 11355 5645 11395
rect 5605 11325 5610 11355
rect 5640 11325 5645 11355
rect 5605 11320 5645 11325
rect 5805 11425 5845 11430
rect 5805 11395 5810 11425
rect 5840 11395 5845 11425
rect 5805 11355 5845 11395
rect 5805 11325 5810 11355
rect 5840 11325 5845 11355
rect 5805 11320 5845 11325
rect 6005 11425 6045 11430
rect 6005 11395 6010 11425
rect 6040 11395 6045 11425
rect 6005 11355 6045 11395
rect 6005 11325 6010 11355
rect 6040 11325 6045 11355
rect 6005 11320 6045 11325
rect 6205 11425 6245 11430
rect 6205 11395 6210 11425
rect 6240 11395 6245 11425
rect 6205 11355 6245 11395
rect 6205 11325 6210 11355
rect 6240 11325 6245 11355
rect 6205 11320 6245 11325
rect 6405 11425 6445 11430
rect 6405 11395 6410 11425
rect 6440 11395 6445 11425
rect 6405 11355 6445 11395
rect 6405 11325 6410 11355
rect 6440 11325 6445 11355
rect 6405 11320 6445 11325
rect -195 11240 -155 11245
rect -195 11210 -190 11240
rect -160 11210 -155 11240
rect -195 11170 -155 11210
rect -195 11140 -190 11170
rect -160 11140 -155 11170
rect -195 11135 -155 11140
rect 5 11240 45 11245
rect 5 11210 10 11240
rect 40 11210 45 11240
rect 5 11170 45 11210
rect 5 11140 10 11170
rect 40 11140 45 11170
rect 5 11135 45 11140
rect 205 11240 245 11245
rect 205 11210 210 11240
rect 240 11210 245 11240
rect 205 11170 245 11210
rect 205 11140 210 11170
rect 240 11140 245 11170
rect 205 11135 245 11140
rect 405 11240 445 11245
rect 405 11210 410 11240
rect 440 11210 445 11240
rect 405 11170 445 11210
rect 405 11140 410 11170
rect 440 11140 445 11170
rect 405 11135 445 11140
rect 605 11240 645 11245
rect 605 11210 610 11240
rect 640 11210 645 11240
rect 605 11170 645 11210
rect 605 11140 610 11170
rect 640 11140 645 11170
rect 605 11135 645 11140
rect 805 11240 845 11245
rect 805 11210 810 11240
rect 840 11210 845 11240
rect 805 11170 845 11210
rect 805 11140 810 11170
rect 840 11140 845 11170
rect 805 11135 845 11140
rect 1005 11240 1045 11245
rect 1005 11210 1010 11240
rect 1040 11210 1045 11240
rect 1005 11170 1045 11210
rect 1005 11140 1010 11170
rect 1040 11140 1045 11170
rect 1005 11135 1045 11140
rect 1205 11240 1245 11245
rect 1205 11210 1210 11240
rect 1240 11210 1245 11240
rect 1205 11170 1245 11210
rect 1205 11140 1210 11170
rect 1240 11140 1245 11170
rect 1205 11135 1245 11140
rect 1405 11240 1445 11245
rect 1405 11210 1410 11240
rect 1440 11210 1445 11240
rect 1405 11170 1445 11210
rect 1405 11140 1410 11170
rect 1440 11140 1445 11170
rect 1405 11135 1445 11140
rect 1605 11240 1645 11245
rect 1605 11210 1610 11240
rect 1640 11210 1645 11240
rect 1605 11170 1645 11210
rect 1605 11140 1610 11170
rect 1640 11140 1645 11170
rect 1605 11135 1645 11140
rect 1805 11240 1845 11245
rect 1805 11210 1810 11240
rect 1840 11210 1845 11240
rect 1805 11170 1845 11210
rect 1805 11140 1810 11170
rect 1840 11140 1845 11170
rect 1805 11135 1845 11140
rect 2005 11240 2045 11245
rect 2005 11210 2010 11240
rect 2040 11210 2045 11240
rect 2005 11170 2045 11210
rect 2005 11140 2010 11170
rect 2040 11140 2045 11170
rect 2005 11135 2045 11140
rect 2205 11240 2245 11245
rect 2205 11210 2210 11240
rect 2240 11210 2245 11240
rect 2205 11170 2245 11210
rect 2205 11140 2210 11170
rect 2240 11140 2245 11170
rect 2205 11135 2245 11140
rect 2405 11240 2445 11245
rect 2405 11210 2410 11240
rect 2440 11210 2445 11240
rect 2405 11170 2445 11210
rect 2405 11140 2410 11170
rect 2440 11140 2445 11170
rect 2405 11135 2445 11140
rect 2605 11240 2645 11245
rect 2605 11210 2610 11240
rect 2640 11210 2645 11240
rect 2605 11170 2645 11210
rect 2605 11140 2610 11170
rect 2640 11140 2645 11170
rect 2605 11135 2645 11140
rect 2805 11240 2845 11245
rect 2805 11210 2810 11240
rect 2840 11210 2845 11240
rect 2805 11170 2845 11210
rect 2805 11140 2810 11170
rect 2840 11140 2845 11170
rect 2805 11135 2845 11140
rect 3005 11240 3045 11245
rect 3005 11210 3010 11240
rect 3040 11210 3045 11240
rect 3005 11170 3045 11210
rect 3005 11140 3010 11170
rect 3040 11140 3045 11170
rect 3005 11135 3045 11140
rect 3205 11240 3245 11245
rect 3205 11210 3210 11240
rect 3240 11210 3245 11240
rect 3205 11170 3245 11210
rect 3205 11140 3210 11170
rect 3240 11140 3245 11170
rect 3205 11135 3245 11140
rect 3405 11240 3445 11245
rect 3405 11210 3410 11240
rect 3440 11210 3445 11240
rect 3405 11170 3445 11210
rect 3405 11140 3410 11170
rect 3440 11140 3445 11170
rect 3405 11135 3445 11140
rect 3605 11240 3645 11245
rect 3605 11210 3610 11240
rect 3640 11210 3645 11240
rect 3605 11170 3645 11210
rect 3605 11140 3610 11170
rect 3640 11140 3645 11170
rect 3605 11135 3645 11140
rect 3805 11240 3845 11245
rect 3805 11210 3810 11240
rect 3840 11210 3845 11240
rect 3805 11170 3845 11210
rect 3805 11140 3810 11170
rect 3840 11140 3845 11170
rect 3805 11135 3845 11140
rect 4005 11240 4045 11245
rect 4005 11210 4010 11240
rect 4040 11210 4045 11240
rect 4005 11170 4045 11210
rect 4005 11140 4010 11170
rect 4040 11140 4045 11170
rect 4005 11135 4045 11140
rect 4205 11240 4245 11245
rect 4205 11210 4210 11240
rect 4240 11210 4245 11240
rect 4205 11170 4245 11210
rect 4205 11140 4210 11170
rect 4240 11140 4245 11170
rect 4205 11135 4245 11140
rect 4405 11240 4445 11245
rect 4405 11210 4410 11240
rect 4440 11210 4445 11240
rect 4405 11170 4445 11210
rect 4405 11140 4410 11170
rect 4440 11140 4445 11170
rect 4405 11135 4445 11140
rect 4605 11240 4645 11245
rect 4605 11210 4610 11240
rect 4640 11210 4645 11240
rect 4605 11170 4645 11210
rect 4605 11140 4610 11170
rect 4640 11140 4645 11170
rect 4605 11135 4645 11140
rect 4805 11240 4845 11245
rect 4805 11210 4810 11240
rect 4840 11210 4845 11240
rect 4805 11170 4845 11210
rect 4805 11140 4810 11170
rect 4840 11140 4845 11170
rect 4805 11135 4845 11140
rect 5005 11240 5045 11245
rect 5005 11210 5010 11240
rect 5040 11210 5045 11240
rect 5005 11170 5045 11210
rect 5005 11140 5010 11170
rect 5040 11140 5045 11170
rect 5005 11135 5045 11140
rect 5205 11240 5245 11245
rect 5205 11210 5210 11240
rect 5240 11210 5245 11240
rect 5205 11170 5245 11210
rect 5205 11140 5210 11170
rect 5240 11140 5245 11170
rect 5205 11135 5245 11140
rect 5405 11240 5445 11245
rect 5405 11210 5410 11240
rect 5440 11210 5445 11240
rect 5405 11170 5445 11210
rect 5405 11140 5410 11170
rect 5440 11140 5445 11170
rect 5405 11135 5445 11140
rect 5605 11240 5645 11245
rect 5605 11210 5610 11240
rect 5640 11210 5645 11240
rect 5605 11170 5645 11210
rect 5605 11140 5610 11170
rect 5640 11140 5645 11170
rect 5605 11135 5645 11140
rect 5805 11240 5845 11245
rect 5805 11210 5810 11240
rect 5840 11210 5845 11240
rect 5805 11170 5845 11210
rect 5805 11140 5810 11170
rect 5840 11140 5845 11170
rect 5805 11135 5845 11140
rect 6005 11240 6045 11245
rect 6005 11210 6010 11240
rect 6040 11210 6045 11240
rect 6005 11170 6045 11210
rect 6005 11140 6010 11170
rect 6040 11140 6045 11170
rect 6005 11135 6045 11140
rect 6205 11240 6245 11245
rect 6205 11210 6210 11240
rect 6240 11210 6245 11240
rect 6205 11170 6245 11210
rect 6205 11140 6210 11170
rect 6240 11140 6245 11170
rect 6205 11135 6245 11140
rect 6405 11240 6445 11245
rect 6405 11210 6410 11240
rect 6440 11210 6445 11240
rect 6405 11170 6445 11210
rect 6405 11140 6410 11170
rect 6440 11140 6445 11170
rect 6405 11135 6445 11140
rect -195 11055 -155 11060
rect -195 11025 -190 11055
rect -160 11025 -155 11055
rect -195 10985 -155 11025
rect -195 10955 -190 10985
rect -160 10955 -155 10985
rect -195 10950 -155 10955
rect 5 11055 45 11060
rect 5 11025 10 11055
rect 40 11025 45 11055
rect 5 10985 45 11025
rect 5 10955 10 10985
rect 40 10955 45 10985
rect 5 10950 45 10955
rect 205 11055 245 11060
rect 205 11025 210 11055
rect 240 11025 245 11055
rect 205 10985 245 11025
rect 205 10955 210 10985
rect 240 10955 245 10985
rect 205 10950 245 10955
rect 405 11055 445 11060
rect 405 11025 410 11055
rect 440 11025 445 11055
rect 405 10985 445 11025
rect 405 10955 410 10985
rect 440 10955 445 10985
rect 405 10950 445 10955
rect 605 11055 645 11060
rect 605 11025 610 11055
rect 640 11025 645 11055
rect 605 10985 645 11025
rect 605 10955 610 10985
rect 640 10955 645 10985
rect 605 10950 645 10955
rect 805 11055 845 11060
rect 805 11025 810 11055
rect 840 11025 845 11055
rect 805 10985 845 11025
rect 805 10955 810 10985
rect 840 10955 845 10985
rect 805 10950 845 10955
rect 1005 11055 1045 11060
rect 1005 11025 1010 11055
rect 1040 11025 1045 11055
rect 1005 10985 1045 11025
rect 1005 10955 1010 10985
rect 1040 10955 1045 10985
rect 1005 10950 1045 10955
rect 1205 11055 1245 11060
rect 1205 11025 1210 11055
rect 1240 11025 1245 11055
rect 1205 10985 1245 11025
rect 1205 10955 1210 10985
rect 1240 10955 1245 10985
rect 1205 10950 1245 10955
rect 1405 11055 1445 11060
rect 1405 11025 1410 11055
rect 1440 11025 1445 11055
rect 1405 10985 1445 11025
rect 1405 10955 1410 10985
rect 1440 10955 1445 10985
rect 1405 10950 1445 10955
rect 1605 11055 1645 11060
rect 1605 11025 1610 11055
rect 1640 11025 1645 11055
rect 1605 10985 1645 11025
rect 1605 10955 1610 10985
rect 1640 10955 1645 10985
rect 1605 10950 1645 10955
rect 1805 11055 1845 11060
rect 1805 11025 1810 11055
rect 1840 11025 1845 11055
rect 1805 10985 1845 11025
rect 1805 10955 1810 10985
rect 1840 10955 1845 10985
rect 1805 10950 1845 10955
rect 2005 11055 2045 11060
rect 2005 11025 2010 11055
rect 2040 11025 2045 11055
rect 2005 10985 2045 11025
rect 2005 10955 2010 10985
rect 2040 10955 2045 10985
rect 2005 10950 2045 10955
rect 2205 11055 2245 11060
rect 2205 11025 2210 11055
rect 2240 11025 2245 11055
rect 2205 10985 2245 11025
rect 2205 10955 2210 10985
rect 2240 10955 2245 10985
rect 2205 10950 2245 10955
rect 2405 11055 2445 11060
rect 2405 11025 2410 11055
rect 2440 11025 2445 11055
rect 2405 10985 2445 11025
rect 2405 10955 2410 10985
rect 2440 10955 2445 10985
rect 2405 10950 2445 10955
rect 2605 11055 2645 11060
rect 2605 11025 2610 11055
rect 2640 11025 2645 11055
rect 2605 10985 2645 11025
rect 2605 10955 2610 10985
rect 2640 10955 2645 10985
rect 2605 10950 2645 10955
rect 2805 11055 2845 11060
rect 2805 11025 2810 11055
rect 2840 11025 2845 11055
rect 2805 10985 2845 11025
rect 2805 10955 2810 10985
rect 2840 10955 2845 10985
rect 2805 10950 2845 10955
rect 3005 11055 3045 11060
rect 3005 11025 3010 11055
rect 3040 11025 3045 11055
rect 3005 10985 3045 11025
rect 3005 10955 3010 10985
rect 3040 10955 3045 10985
rect 3005 10950 3045 10955
rect 3205 11055 3245 11060
rect 3205 11025 3210 11055
rect 3240 11025 3245 11055
rect 3205 10985 3245 11025
rect 3205 10955 3210 10985
rect 3240 10955 3245 10985
rect 3205 10950 3245 10955
rect 3405 11055 3445 11060
rect 3405 11025 3410 11055
rect 3440 11025 3445 11055
rect 3405 10985 3445 11025
rect 3405 10955 3410 10985
rect 3440 10955 3445 10985
rect 3405 10950 3445 10955
rect 3605 11055 3645 11060
rect 3605 11025 3610 11055
rect 3640 11025 3645 11055
rect 3605 10985 3645 11025
rect 3605 10955 3610 10985
rect 3640 10955 3645 10985
rect 3605 10950 3645 10955
rect 3805 11055 3845 11060
rect 3805 11025 3810 11055
rect 3840 11025 3845 11055
rect 3805 10985 3845 11025
rect 3805 10955 3810 10985
rect 3840 10955 3845 10985
rect 3805 10950 3845 10955
rect 4005 11055 4045 11060
rect 4005 11025 4010 11055
rect 4040 11025 4045 11055
rect 4005 10985 4045 11025
rect 4005 10955 4010 10985
rect 4040 10955 4045 10985
rect 4005 10950 4045 10955
rect 4205 11055 4245 11060
rect 4205 11025 4210 11055
rect 4240 11025 4245 11055
rect 4205 10985 4245 11025
rect 4205 10955 4210 10985
rect 4240 10955 4245 10985
rect 4205 10950 4245 10955
rect 4405 11055 4445 11060
rect 4405 11025 4410 11055
rect 4440 11025 4445 11055
rect 4405 10985 4445 11025
rect 4405 10955 4410 10985
rect 4440 10955 4445 10985
rect 4405 10950 4445 10955
rect 4605 11055 4645 11060
rect 4605 11025 4610 11055
rect 4640 11025 4645 11055
rect 4605 10985 4645 11025
rect 4605 10955 4610 10985
rect 4640 10955 4645 10985
rect 4605 10950 4645 10955
rect 4805 11055 4845 11060
rect 4805 11025 4810 11055
rect 4840 11025 4845 11055
rect 4805 10985 4845 11025
rect 4805 10955 4810 10985
rect 4840 10955 4845 10985
rect 4805 10950 4845 10955
rect 5005 11055 5045 11060
rect 5005 11025 5010 11055
rect 5040 11025 5045 11055
rect 5005 10985 5045 11025
rect 5005 10955 5010 10985
rect 5040 10955 5045 10985
rect 5005 10950 5045 10955
rect 5205 11055 5245 11060
rect 5205 11025 5210 11055
rect 5240 11025 5245 11055
rect 5205 10985 5245 11025
rect 5205 10955 5210 10985
rect 5240 10955 5245 10985
rect 5205 10950 5245 10955
rect 5405 11055 5445 11060
rect 5405 11025 5410 11055
rect 5440 11025 5445 11055
rect 5405 10985 5445 11025
rect 5405 10955 5410 10985
rect 5440 10955 5445 10985
rect 5405 10950 5445 10955
rect 5605 11055 5645 11060
rect 5605 11025 5610 11055
rect 5640 11025 5645 11055
rect 5605 10985 5645 11025
rect 5605 10955 5610 10985
rect 5640 10955 5645 10985
rect 5605 10950 5645 10955
rect 5805 11055 5845 11060
rect 5805 11025 5810 11055
rect 5840 11025 5845 11055
rect 5805 10985 5845 11025
rect 5805 10955 5810 10985
rect 5840 10955 5845 10985
rect 5805 10950 5845 10955
rect 6005 11055 6045 11060
rect 6005 11025 6010 11055
rect 6040 11025 6045 11055
rect 6005 10985 6045 11025
rect 6005 10955 6010 10985
rect 6040 10955 6045 10985
rect 6005 10950 6045 10955
rect 6205 11055 6245 11060
rect 6205 11025 6210 11055
rect 6240 11025 6245 11055
rect 6205 10985 6245 11025
rect 6205 10955 6210 10985
rect 6240 10955 6245 10985
rect 6205 10950 6245 10955
rect 6405 11055 6445 11060
rect 6405 11025 6410 11055
rect 6440 11025 6445 11055
rect 6405 10985 6445 11025
rect 6405 10955 6410 10985
rect 6440 10955 6445 10985
rect 6405 10950 6445 10955
rect -195 10870 -155 10875
rect -195 10840 -190 10870
rect -160 10840 -155 10870
rect -195 10800 -155 10840
rect -195 10770 -190 10800
rect -160 10770 -155 10800
rect -195 10765 -155 10770
rect 5 10870 45 10875
rect 5 10840 10 10870
rect 40 10840 45 10870
rect 5 10800 45 10840
rect 5 10770 10 10800
rect 40 10770 45 10800
rect 5 10765 45 10770
rect 205 10870 245 10875
rect 205 10840 210 10870
rect 240 10840 245 10870
rect 205 10800 245 10840
rect 205 10770 210 10800
rect 240 10770 245 10800
rect 205 10765 245 10770
rect 405 10870 445 10875
rect 405 10840 410 10870
rect 440 10840 445 10870
rect 405 10800 445 10840
rect 405 10770 410 10800
rect 440 10770 445 10800
rect 405 10765 445 10770
rect 605 10870 645 10875
rect 605 10840 610 10870
rect 640 10840 645 10870
rect 605 10800 645 10840
rect 605 10770 610 10800
rect 640 10770 645 10800
rect 605 10765 645 10770
rect 805 10870 845 10875
rect 805 10840 810 10870
rect 840 10840 845 10870
rect 805 10800 845 10840
rect 805 10770 810 10800
rect 840 10770 845 10800
rect 805 10765 845 10770
rect 1005 10870 1045 10875
rect 1005 10840 1010 10870
rect 1040 10840 1045 10870
rect 1005 10800 1045 10840
rect 1005 10770 1010 10800
rect 1040 10770 1045 10800
rect 1005 10765 1045 10770
rect 1205 10870 1245 10875
rect 1205 10840 1210 10870
rect 1240 10840 1245 10870
rect 1205 10800 1245 10840
rect 1205 10770 1210 10800
rect 1240 10770 1245 10800
rect 1205 10765 1245 10770
rect 1405 10870 1445 10875
rect 1405 10840 1410 10870
rect 1440 10840 1445 10870
rect 1405 10800 1445 10840
rect 1405 10770 1410 10800
rect 1440 10770 1445 10800
rect 1405 10765 1445 10770
rect 1605 10870 1645 10875
rect 1605 10840 1610 10870
rect 1640 10840 1645 10870
rect 1605 10800 1645 10840
rect 1605 10770 1610 10800
rect 1640 10770 1645 10800
rect 1605 10765 1645 10770
rect 1805 10870 1845 10875
rect 1805 10840 1810 10870
rect 1840 10840 1845 10870
rect 1805 10800 1845 10840
rect 1805 10770 1810 10800
rect 1840 10770 1845 10800
rect 1805 10765 1845 10770
rect 2005 10870 2045 10875
rect 2005 10840 2010 10870
rect 2040 10840 2045 10870
rect 2005 10800 2045 10840
rect 2005 10770 2010 10800
rect 2040 10770 2045 10800
rect 2005 10765 2045 10770
rect 2205 10870 2245 10875
rect 2205 10840 2210 10870
rect 2240 10840 2245 10870
rect 2205 10800 2245 10840
rect 2205 10770 2210 10800
rect 2240 10770 2245 10800
rect 2205 10765 2245 10770
rect 2405 10870 2445 10875
rect 2405 10840 2410 10870
rect 2440 10840 2445 10870
rect 2405 10800 2445 10840
rect 2405 10770 2410 10800
rect 2440 10770 2445 10800
rect 2405 10765 2445 10770
rect 2605 10870 2645 10875
rect 2605 10840 2610 10870
rect 2640 10840 2645 10870
rect 2605 10800 2645 10840
rect 2605 10770 2610 10800
rect 2640 10770 2645 10800
rect 2605 10765 2645 10770
rect 2805 10870 2845 10875
rect 2805 10840 2810 10870
rect 2840 10840 2845 10870
rect 2805 10800 2845 10840
rect 2805 10770 2810 10800
rect 2840 10770 2845 10800
rect 2805 10765 2845 10770
rect 3005 10870 3045 10875
rect 3005 10840 3010 10870
rect 3040 10840 3045 10870
rect 3005 10800 3045 10840
rect 3005 10770 3010 10800
rect 3040 10770 3045 10800
rect 3005 10765 3045 10770
rect 3205 10870 3245 10875
rect 3205 10840 3210 10870
rect 3240 10840 3245 10870
rect 3205 10800 3245 10840
rect 3205 10770 3210 10800
rect 3240 10770 3245 10800
rect 3205 10765 3245 10770
rect 3405 10870 3445 10875
rect 3405 10840 3410 10870
rect 3440 10840 3445 10870
rect 3405 10800 3445 10840
rect 3405 10770 3410 10800
rect 3440 10770 3445 10800
rect 3405 10765 3445 10770
rect 3605 10870 3645 10875
rect 3605 10840 3610 10870
rect 3640 10840 3645 10870
rect 3605 10800 3645 10840
rect 3605 10770 3610 10800
rect 3640 10770 3645 10800
rect 3605 10765 3645 10770
rect 3805 10870 3845 10875
rect 3805 10840 3810 10870
rect 3840 10840 3845 10870
rect 3805 10800 3845 10840
rect 3805 10770 3810 10800
rect 3840 10770 3845 10800
rect 3805 10765 3845 10770
rect 4005 10870 4045 10875
rect 4005 10840 4010 10870
rect 4040 10840 4045 10870
rect 4005 10800 4045 10840
rect 4005 10770 4010 10800
rect 4040 10770 4045 10800
rect 4005 10765 4045 10770
rect 4205 10870 4245 10875
rect 4205 10840 4210 10870
rect 4240 10840 4245 10870
rect 4205 10800 4245 10840
rect 4205 10770 4210 10800
rect 4240 10770 4245 10800
rect 4205 10765 4245 10770
rect 4405 10870 4445 10875
rect 4405 10840 4410 10870
rect 4440 10840 4445 10870
rect 4405 10800 4445 10840
rect 4405 10770 4410 10800
rect 4440 10770 4445 10800
rect 4405 10765 4445 10770
rect 4605 10870 4645 10875
rect 4605 10840 4610 10870
rect 4640 10840 4645 10870
rect 4605 10800 4645 10840
rect 4605 10770 4610 10800
rect 4640 10770 4645 10800
rect 4605 10765 4645 10770
rect 4805 10870 4845 10875
rect 4805 10840 4810 10870
rect 4840 10840 4845 10870
rect 4805 10800 4845 10840
rect 4805 10770 4810 10800
rect 4840 10770 4845 10800
rect 4805 10765 4845 10770
rect 5005 10870 5045 10875
rect 5005 10840 5010 10870
rect 5040 10840 5045 10870
rect 5005 10800 5045 10840
rect 5005 10770 5010 10800
rect 5040 10770 5045 10800
rect 5005 10765 5045 10770
rect 5205 10870 5245 10875
rect 5205 10840 5210 10870
rect 5240 10840 5245 10870
rect 5205 10800 5245 10840
rect 5205 10770 5210 10800
rect 5240 10770 5245 10800
rect 5205 10765 5245 10770
rect 5405 10870 5445 10875
rect 5405 10840 5410 10870
rect 5440 10840 5445 10870
rect 5405 10800 5445 10840
rect 5405 10770 5410 10800
rect 5440 10770 5445 10800
rect 5405 10765 5445 10770
rect 5605 10870 5645 10875
rect 5605 10840 5610 10870
rect 5640 10840 5645 10870
rect 5605 10800 5645 10840
rect 5605 10770 5610 10800
rect 5640 10770 5645 10800
rect 5605 10765 5645 10770
rect 5805 10870 5845 10875
rect 5805 10840 5810 10870
rect 5840 10840 5845 10870
rect 5805 10800 5845 10840
rect 5805 10770 5810 10800
rect 5840 10770 5845 10800
rect 5805 10765 5845 10770
rect 6005 10870 6045 10875
rect 6005 10840 6010 10870
rect 6040 10840 6045 10870
rect 6005 10800 6045 10840
rect 6005 10770 6010 10800
rect 6040 10770 6045 10800
rect 6005 10765 6045 10770
rect 6205 10870 6245 10875
rect 6205 10840 6210 10870
rect 6240 10840 6245 10870
rect 6205 10800 6245 10840
rect 6205 10770 6210 10800
rect 6240 10770 6245 10800
rect 6205 10765 6245 10770
rect 6405 10870 6445 10875
rect 6405 10840 6410 10870
rect 6440 10840 6445 10870
rect 6405 10800 6445 10840
rect 6405 10770 6410 10800
rect 6440 10770 6445 10800
rect 6405 10765 6445 10770
rect -195 10685 -155 10690
rect -195 10655 -190 10685
rect -160 10655 -155 10685
rect -195 10615 -155 10655
rect -195 10585 -190 10615
rect -160 10585 -155 10615
rect -195 10580 -155 10585
rect 5 10685 45 10690
rect 5 10655 10 10685
rect 40 10655 45 10685
rect 5 10615 45 10655
rect 5 10585 10 10615
rect 40 10585 45 10615
rect 5 10580 45 10585
rect 205 10685 245 10690
rect 205 10655 210 10685
rect 240 10655 245 10685
rect 205 10615 245 10655
rect 205 10585 210 10615
rect 240 10585 245 10615
rect 205 10580 245 10585
rect 405 10685 445 10690
rect 405 10655 410 10685
rect 440 10655 445 10685
rect 405 10615 445 10655
rect 405 10585 410 10615
rect 440 10585 445 10615
rect 405 10580 445 10585
rect 605 10685 645 10690
rect 605 10655 610 10685
rect 640 10655 645 10685
rect 605 10615 645 10655
rect 605 10585 610 10615
rect 640 10585 645 10615
rect 605 10580 645 10585
rect 805 10685 845 10690
rect 805 10655 810 10685
rect 840 10655 845 10685
rect 805 10615 845 10655
rect 805 10585 810 10615
rect 840 10585 845 10615
rect 805 10580 845 10585
rect 1005 10685 1045 10690
rect 1005 10655 1010 10685
rect 1040 10655 1045 10685
rect 1005 10615 1045 10655
rect 1005 10585 1010 10615
rect 1040 10585 1045 10615
rect 1005 10580 1045 10585
rect 1205 10685 1245 10690
rect 1205 10655 1210 10685
rect 1240 10655 1245 10685
rect 1205 10615 1245 10655
rect 1205 10585 1210 10615
rect 1240 10585 1245 10615
rect 1205 10580 1245 10585
rect 1405 10685 1445 10690
rect 1405 10655 1410 10685
rect 1440 10655 1445 10685
rect 1405 10615 1445 10655
rect 1405 10585 1410 10615
rect 1440 10585 1445 10615
rect 1405 10580 1445 10585
rect 1605 10685 1645 10690
rect 1605 10655 1610 10685
rect 1640 10655 1645 10685
rect 1605 10615 1645 10655
rect 1605 10585 1610 10615
rect 1640 10585 1645 10615
rect 1605 10580 1645 10585
rect 1805 10685 1845 10690
rect 1805 10655 1810 10685
rect 1840 10655 1845 10685
rect 1805 10615 1845 10655
rect 1805 10585 1810 10615
rect 1840 10585 1845 10615
rect 1805 10580 1845 10585
rect 2005 10685 2045 10690
rect 2005 10655 2010 10685
rect 2040 10655 2045 10685
rect 2005 10615 2045 10655
rect 2005 10585 2010 10615
rect 2040 10585 2045 10615
rect 2005 10580 2045 10585
rect 2205 10685 2245 10690
rect 2205 10655 2210 10685
rect 2240 10655 2245 10685
rect 2205 10615 2245 10655
rect 2205 10585 2210 10615
rect 2240 10585 2245 10615
rect 2205 10580 2245 10585
rect 2405 10685 2445 10690
rect 2405 10655 2410 10685
rect 2440 10655 2445 10685
rect 2405 10615 2445 10655
rect 2405 10585 2410 10615
rect 2440 10585 2445 10615
rect 2405 10580 2445 10585
rect 2605 10685 2645 10690
rect 2605 10655 2610 10685
rect 2640 10655 2645 10685
rect 2605 10615 2645 10655
rect 2605 10585 2610 10615
rect 2640 10585 2645 10615
rect 2605 10580 2645 10585
rect 2805 10685 2845 10690
rect 2805 10655 2810 10685
rect 2840 10655 2845 10685
rect 2805 10615 2845 10655
rect 2805 10585 2810 10615
rect 2840 10585 2845 10615
rect 2805 10580 2845 10585
rect 3005 10685 3045 10690
rect 3005 10655 3010 10685
rect 3040 10655 3045 10685
rect 3005 10615 3045 10655
rect 3005 10585 3010 10615
rect 3040 10585 3045 10615
rect 3005 10580 3045 10585
rect 3205 10685 3245 10690
rect 3205 10655 3210 10685
rect 3240 10655 3245 10685
rect 3205 10615 3245 10655
rect 3205 10585 3210 10615
rect 3240 10585 3245 10615
rect 3205 10580 3245 10585
rect 3405 10685 3445 10690
rect 3405 10655 3410 10685
rect 3440 10655 3445 10685
rect 3405 10615 3445 10655
rect 3405 10585 3410 10615
rect 3440 10585 3445 10615
rect 3405 10580 3445 10585
rect 3605 10685 3645 10690
rect 3605 10655 3610 10685
rect 3640 10655 3645 10685
rect 3605 10615 3645 10655
rect 3605 10585 3610 10615
rect 3640 10585 3645 10615
rect 3605 10580 3645 10585
rect 3805 10685 3845 10690
rect 3805 10655 3810 10685
rect 3840 10655 3845 10685
rect 3805 10615 3845 10655
rect 3805 10585 3810 10615
rect 3840 10585 3845 10615
rect 3805 10580 3845 10585
rect 4005 10685 4045 10690
rect 4005 10655 4010 10685
rect 4040 10655 4045 10685
rect 4005 10615 4045 10655
rect 4005 10585 4010 10615
rect 4040 10585 4045 10615
rect 4005 10580 4045 10585
rect 4205 10685 4245 10690
rect 4205 10655 4210 10685
rect 4240 10655 4245 10685
rect 4205 10615 4245 10655
rect 4205 10585 4210 10615
rect 4240 10585 4245 10615
rect 4205 10580 4245 10585
rect 4405 10685 4445 10690
rect 4405 10655 4410 10685
rect 4440 10655 4445 10685
rect 4405 10615 4445 10655
rect 4405 10585 4410 10615
rect 4440 10585 4445 10615
rect 4405 10580 4445 10585
rect 4605 10685 4645 10690
rect 4605 10655 4610 10685
rect 4640 10655 4645 10685
rect 4605 10615 4645 10655
rect 4605 10585 4610 10615
rect 4640 10585 4645 10615
rect 4605 10580 4645 10585
rect 4805 10685 4845 10690
rect 4805 10655 4810 10685
rect 4840 10655 4845 10685
rect 4805 10615 4845 10655
rect 4805 10585 4810 10615
rect 4840 10585 4845 10615
rect 4805 10580 4845 10585
rect 5005 10685 5045 10690
rect 5005 10655 5010 10685
rect 5040 10655 5045 10685
rect 5005 10615 5045 10655
rect 5005 10585 5010 10615
rect 5040 10585 5045 10615
rect 5005 10580 5045 10585
rect 5205 10685 5245 10690
rect 5205 10655 5210 10685
rect 5240 10655 5245 10685
rect 5205 10615 5245 10655
rect 5205 10585 5210 10615
rect 5240 10585 5245 10615
rect 5205 10580 5245 10585
rect 5405 10685 5445 10690
rect 5405 10655 5410 10685
rect 5440 10655 5445 10685
rect 5405 10615 5445 10655
rect 5405 10585 5410 10615
rect 5440 10585 5445 10615
rect 5405 10580 5445 10585
rect 5605 10685 5645 10690
rect 5605 10655 5610 10685
rect 5640 10655 5645 10685
rect 5605 10615 5645 10655
rect 5605 10585 5610 10615
rect 5640 10585 5645 10615
rect 5605 10580 5645 10585
rect 5805 10685 5845 10690
rect 5805 10655 5810 10685
rect 5840 10655 5845 10685
rect 5805 10615 5845 10655
rect 5805 10585 5810 10615
rect 5840 10585 5845 10615
rect 5805 10580 5845 10585
rect 6005 10685 6045 10690
rect 6005 10655 6010 10685
rect 6040 10655 6045 10685
rect 6005 10615 6045 10655
rect 6005 10585 6010 10615
rect 6040 10585 6045 10615
rect 6005 10580 6045 10585
rect 6205 10685 6245 10690
rect 6205 10655 6210 10685
rect 6240 10655 6245 10685
rect 6205 10615 6245 10655
rect 6205 10585 6210 10615
rect 6240 10585 6245 10615
rect 6205 10580 6245 10585
rect 6405 10685 6445 10690
rect 6405 10655 6410 10685
rect 6440 10655 6445 10685
rect 6405 10615 6445 10655
rect 6405 10585 6410 10615
rect 6440 10585 6445 10615
rect 6405 10580 6445 10585
rect -195 10500 -155 10505
rect -195 10470 -190 10500
rect -160 10470 -155 10500
rect -195 10430 -155 10470
rect -195 10400 -190 10430
rect -160 10400 -155 10430
rect -195 10395 -155 10400
rect 5 10500 45 10505
rect 5 10470 10 10500
rect 40 10470 45 10500
rect 5 10430 45 10470
rect 5 10400 10 10430
rect 40 10400 45 10430
rect 5 10395 45 10400
rect 205 10500 245 10505
rect 205 10470 210 10500
rect 240 10470 245 10500
rect 205 10430 245 10470
rect 205 10400 210 10430
rect 240 10400 245 10430
rect 205 10395 245 10400
rect 405 10500 445 10505
rect 405 10470 410 10500
rect 440 10470 445 10500
rect 405 10430 445 10470
rect 405 10400 410 10430
rect 440 10400 445 10430
rect 405 10395 445 10400
rect 605 10500 645 10505
rect 605 10470 610 10500
rect 640 10470 645 10500
rect 605 10430 645 10470
rect 605 10400 610 10430
rect 640 10400 645 10430
rect 605 10395 645 10400
rect 805 10500 845 10505
rect 805 10470 810 10500
rect 840 10470 845 10500
rect 805 10430 845 10470
rect 805 10400 810 10430
rect 840 10400 845 10430
rect 805 10395 845 10400
rect 1005 10500 1045 10505
rect 1005 10470 1010 10500
rect 1040 10470 1045 10500
rect 1005 10430 1045 10470
rect 1005 10400 1010 10430
rect 1040 10400 1045 10430
rect 1005 10395 1045 10400
rect 1205 10500 1245 10505
rect 1205 10470 1210 10500
rect 1240 10470 1245 10500
rect 1205 10430 1245 10470
rect 1205 10400 1210 10430
rect 1240 10400 1245 10430
rect 1205 10395 1245 10400
rect 1405 10500 1445 10505
rect 1405 10470 1410 10500
rect 1440 10470 1445 10500
rect 1405 10430 1445 10470
rect 1405 10400 1410 10430
rect 1440 10400 1445 10430
rect 1405 10395 1445 10400
rect 1605 10500 1645 10505
rect 1605 10470 1610 10500
rect 1640 10470 1645 10500
rect 1605 10430 1645 10470
rect 1605 10400 1610 10430
rect 1640 10400 1645 10430
rect 1605 10395 1645 10400
rect 1805 10500 1845 10505
rect 1805 10470 1810 10500
rect 1840 10470 1845 10500
rect 1805 10430 1845 10470
rect 1805 10400 1810 10430
rect 1840 10400 1845 10430
rect 1805 10395 1845 10400
rect 2005 10500 2045 10505
rect 2005 10470 2010 10500
rect 2040 10470 2045 10500
rect 2005 10430 2045 10470
rect 2005 10400 2010 10430
rect 2040 10400 2045 10430
rect 2005 10395 2045 10400
rect 2205 10500 2245 10505
rect 2205 10470 2210 10500
rect 2240 10470 2245 10500
rect 2205 10430 2245 10470
rect 2205 10400 2210 10430
rect 2240 10400 2245 10430
rect 2205 10395 2245 10400
rect 2405 10500 2445 10505
rect 2405 10470 2410 10500
rect 2440 10470 2445 10500
rect 2405 10430 2445 10470
rect 2405 10400 2410 10430
rect 2440 10400 2445 10430
rect 2405 10395 2445 10400
rect 2605 10500 2645 10505
rect 2605 10470 2610 10500
rect 2640 10470 2645 10500
rect 2605 10430 2645 10470
rect 2605 10400 2610 10430
rect 2640 10400 2645 10430
rect 2605 10395 2645 10400
rect 2805 10500 2845 10505
rect 2805 10470 2810 10500
rect 2840 10470 2845 10500
rect 2805 10430 2845 10470
rect 2805 10400 2810 10430
rect 2840 10400 2845 10430
rect 2805 10395 2845 10400
rect 3005 10500 3045 10505
rect 3005 10470 3010 10500
rect 3040 10470 3045 10500
rect 3005 10430 3045 10470
rect 3005 10400 3010 10430
rect 3040 10400 3045 10430
rect 3005 10395 3045 10400
rect 3205 10500 3245 10505
rect 3205 10470 3210 10500
rect 3240 10470 3245 10500
rect 3205 10430 3245 10470
rect 3205 10400 3210 10430
rect 3240 10400 3245 10430
rect 3205 10395 3245 10400
rect 3405 10500 3445 10505
rect 3405 10470 3410 10500
rect 3440 10470 3445 10500
rect 3405 10430 3445 10470
rect 3405 10400 3410 10430
rect 3440 10400 3445 10430
rect 3405 10395 3445 10400
rect 3605 10500 3645 10505
rect 3605 10470 3610 10500
rect 3640 10470 3645 10500
rect 3605 10430 3645 10470
rect 3605 10400 3610 10430
rect 3640 10400 3645 10430
rect 3605 10395 3645 10400
rect 3805 10500 3845 10505
rect 3805 10470 3810 10500
rect 3840 10470 3845 10500
rect 3805 10430 3845 10470
rect 3805 10400 3810 10430
rect 3840 10400 3845 10430
rect 3805 10395 3845 10400
rect 4005 10500 4045 10505
rect 4005 10470 4010 10500
rect 4040 10470 4045 10500
rect 4005 10430 4045 10470
rect 4005 10400 4010 10430
rect 4040 10400 4045 10430
rect 4005 10395 4045 10400
rect 4205 10500 4245 10505
rect 4205 10470 4210 10500
rect 4240 10470 4245 10500
rect 4205 10430 4245 10470
rect 4205 10400 4210 10430
rect 4240 10400 4245 10430
rect 4205 10395 4245 10400
rect 4405 10500 4445 10505
rect 4405 10470 4410 10500
rect 4440 10470 4445 10500
rect 4405 10430 4445 10470
rect 4405 10400 4410 10430
rect 4440 10400 4445 10430
rect 4405 10395 4445 10400
rect 4605 10500 4645 10505
rect 4605 10470 4610 10500
rect 4640 10470 4645 10500
rect 4605 10430 4645 10470
rect 4605 10400 4610 10430
rect 4640 10400 4645 10430
rect 4605 10395 4645 10400
rect 4805 10500 4845 10505
rect 4805 10470 4810 10500
rect 4840 10470 4845 10500
rect 4805 10430 4845 10470
rect 4805 10400 4810 10430
rect 4840 10400 4845 10430
rect 4805 10395 4845 10400
rect 5005 10500 5045 10505
rect 5005 10470 5010 10500
rect 5040 10470 5045 10500
rect 5005 10430 5045 10470
rect 5005 10400 5010 10430
rect 5040 10400 5045 10430
rect 5005 10395 5045 10400
rect 5205 10500 5245 10505
rect 5205 10470 5210 10500
rect 5240 10470 5245 10500
rect 5205 10430 5245 10470
rect 5205 10400 5210 10430
rect 5240 10400 5245 10430
rect 5205 10395 5245 10400
rect 5405 10500 5445 10505
rect 5405 10470 5410 10500
rect 5440 10470 5445 10500
rect 5405 10430 5445 10470
rect 5405 10400 5410 10430
rect 5440 10400 5445 10430
rect 5405 10395 5445 10400
rect 5605 10500 5645 10505
rect 5605 10470 5610 10500
rect 5640 10470 5645 10500
rect 5605 10430 5645 10470
rect 5605 10400 5610 10430
rect 5640 10400 5645 10430
rect 5605 10395 5645 10400
rect 5805 10500 5845 10505
rect 5805 10470 5810 10500
rect 5840 10470 5845 10500
rect 5805 10430 5845 10470
rect 5805 10400 5810 10430
rect 5840 10400 5845 10430
rect 5805 10395 5845 10400
rect 6005 10500 6045 10505
rect 6005 10470 6010 10500
rect 6040 10470 6045 10500
rect 6005 10430 6045 10470
rect 6005 10400 6010 10430
rect 6040 10400 6045 10430
rect 6005 10395 6045 10400
rect 6205 10500 6245 10505
rect 6205 10470 6210 10500
rect 6240 10470 6245 10500
rect 6205 10430 6245 10470
rect 6205 10400 6210 10430
rect 6240 10400 6245 10430
rect 6205 10395 6245 10400
rect 6405 10500 6445 10505
rect 6405 10470 6410 10500
rect 6440 10470 6445 10500
rect 6405 10430 6445 10470
rect 6405 10400 6410 10430
rect 6440 10400 6445 10430
rect 6405 10395 6445 10400
rect -195 10315 -155 10320
rect -195 10285 -190 10315
rect -160 10285 -155 10315
rect -195 10245 -155 10285
rect -195 10215 -190 10245
rect -160 10215 -155 10245
rect -195 10210 -155 10215
rect 5 10315 45 10320
rect 5 10285 10 10315
rect 40 10285 45 10315
rect 5 10245 45 10285
rect 5 10215 10 10245
rect 40 10215 45 10245
rect 5 10210 45 10215
rect 205 10315 245 10320
rect 205 10285 210 10315
rect 240 10285 245 10315
rect 205 10245 245 10285
rect 205 10215 210 10245
rect 240 10215 245 10245
rect 205 10210 245 10215
rect 405 10315 445 10320
rect 405 10285 410 10315
rect 440 10285 445 10315
rect 405 10245 445 10285
rect 405 10215 410 10245
rect 440 10215 445 10245
rect 405 10210 445 10215
rect 605 10315 645 10320
rect 605 10285 610 10315
rect 640 10285 645 10315
rect 605 10245 645 10285
rect 605 10215 610 10245
rect 640 10215 645 10245
rect 605 10210 645 10215
rect 805 10315 845 10320
rect 805 10285 810 10315
rect 840 10285 845 10315
rect 805 10245 845 10285
rect 805 10215 810 10245
rect 840 10215 845 10245
rect 805 10210 845 10215
rect 1005 10315 1045 10320
rect 1005 10285 1010 10315
rect 1040 10285 1045 10315
rect 1005 10245 1045 10285
rect 1005 10215 1010 10245
rect 1040 10215 1045 10245
rect 1005 10210 1045 10215
rect 1205 10315 1245 10320
rect 1205 10285 1210 10315
rect 1240 10285 1245 10315
rect 1205 10245 1245 10285
rect 1205 10215 1210 10245
rect 1240 10215 1245 10245
rect 1205 10210 1245 10215
rect 1405 10315 1445 10320
rect 1405 10285 1410 10315
rect 1440 10285 1445 10315
rect 1405 10245 1445 10285
rect 1405 10215 1410 10245
rect 1440 10215 1445 10245
rect 1405 10210 1445 10215
rect 1605 10315 1645 10320
rect 1605 10285 1610 10315
rect 1640 10285 1645 10315
rect 1605 10245 1645 10285
rect 1605 10215 1610 10245
rect 1640 10215 1645 10245
rect 1605 10210 1645 10215
rect 1805 10315 1845 10320
rect 1805 10285 1810 10315
rect 1840 10285 1845 10315
rect 1805 10245 1845 10285
rect 1805 10215 1810 10245
rect 1840 10215 1845 10245
rect 1805 10210 1845 10215
rect 2005 10315 2045 10320
rect 2005 10285 2010 10315
rect 2040 10285 2045 10315
rect 2005 10245 2045 10285
rect 2005 10215 2010 10245
rect 2040 10215 2045 10245
rect 2005 10210 2045 10215
rect 2205 10315 2245 10320
rect 2205 10285 2210 10315
rect 2240 10285 2245 10315
rect 2205 10245 2245 10285
rect 2205 10215 2210 10245
rect 2240 10215 2245 10245
rect 2205 10210 2245 10215
rect 2405 10315 2445 10320
rect 2405 10285 2410 10315
rect 2440 10285 2445 10315
rect 2405 10245 2445 10285
rect 2405 10215 2410 10245
rect 2440 10215 2445 10245
rect 2405 10210 2445 10215
rect 2605 10315 2645 10320
rect 2605 10285 2610 10315
rect 2640 10285 2645 10315
rect 2605 10245 2645 10285
rect 2605 10215 2610 10245
rect 2640 10215 2645 10245
rect 2605 10210 2645 10215
rect 2805 10315 2845 10320
rect 2805 10285 2810 10315
rect 2840 10285 2845 10315
rect 2805 10245 2845 10285
rect 2805 10215 2810 10245
rect 2840 10215 2845 10245
rect 2805 10210 2845 10215
rect 3005 10315 3045 10320
rect 3005 10285 3010 10315
rect 3040 10285 3045 10315
rect 3005 10245 3045 10285
rect 3005 10215 3010 10245
rect 3040 10215 3045 10245
rect 3005 10210 3045 10215
rect 3205 10315 3245 10320
rect 3205 10285 3210 10315
rect 3240 10285 3245 10315
rect 3205 10245 3245 10285
rect 3205 10215 3210 10245
rect 3240 10215 3245 10245
rect 3205 10210 3245 10215
rect 3405 10315 3445 10320
rect 3405 10285 3410 10315
rect 3440 10285 3445 10315
rect 3405 10245 3445 10285
rect 3405 10215 3410 10245
rect 3440 10215 3445 10245
rect 3405 10210 3445 10215
rect 3605 10315 3645 10320
rect 3605 10285 3610 10315
rect 3640 10285 3645 10315
rect 3605 10245 3645 10285
rect 3605 10215 3610 10245
rect 3640 10215 3645 10245
rect 3605 10210 3645 10215
rect 3805 10315 3845 10320
rect 3805 10285 3810 10315
rect 3840 10285 3845 10315
rect 3805 10245 3845 10285
rect 3805 10215 3810 10245
rect 3840 10215 3845 10245
rect 3805 10210 3845 10215
rect 4005 10315 4045 10320
rect 4005 10285 4010 10315
rect 4040 10285 4045 10315
rect 4005 10245 4045 10285
rect 4005 10215 4010 10245
rect 4040 10215 4045 10245
rect 4005 10210 4045 10215
rect 4205 10315 4245 10320
rect 4205 10285 4210 10315
rect 4240 10285 4245 10315
rect 4205 10245 4245 10285
rect 4205 10215 4210 10245
rect 4240 10215 4245 10245
rect 4205 10210 4245 10215
rect 4405 10315 4445 10320
rect 4405 10285 4410 10315
rect 4440 10285 4445 10315
rect 4405 10245 4445 10285
rect 4405 10215 4410 10245
rect 4440 10215 4445 10245
rect 4405 10210 4445 10215
rect 4605 10315 4645 10320
rect 4605 10285 4610 10315
rect 4640 10285 4645 10315
rect 4605 10245 4645 10285
rect 4605 10215 4610 10245
rect 4640 10215 4645 10245
rect 4605 10210 4645 10215
rect 4805 10315 4845 10320
rect 4805 10285 4810 10315
rect 4840 10285 4845 10315
rect 4805 10245 4845 10285
rect 4805 10215 4810 10245
rect 4840 10215 4845 10245
rect 4805 10210 4845 10215
rect 5005 10315 5045 10320
rect 5005 10285 5010 10315
rect 5040 10285 5045 10315
rect 5005 10245 5045 10285
rect 5005 10215 5010 10245
rect 5040 10215 5045 10245
rect 5005 10210 5045 10215
rect 5205 10315 5245 10320
rect 5205 10285 5210 10315
rect 5240 10285 5245 10315
rect 5205 10245 5245 10285
rect 5205 10215 5210 10245
rect 5240 10215 5245 10245
rect 5205 10210 5245 10215
rect 5405 10315 5445 10320
rect 5405 10285 5410 10315
rect 5440 10285 5445 10315
rect 5405 10245 5445 10285
rect 5405 10215 5410 10245
rect 5440 10215 5445 10245
rect 5405 10210 5445 10215
rect 5605 10315 5645 10320
rect 5605 10285 5610 10315
rect 5640 10285 5645 10315
rect 5605 10245 5645 10285
rect 5605 10215 5610 10245
rect 5640 10215 5645 10245
rect 5605 10210 5645 10215
rect 5805 10315 5845 10320
rect 5805 10285 5810 10315
rect 5840 10285 5845 10315
rect 5805 10245 5845 10285
rect 5805 10215 5810 10245
rect 5840 10215 5845 10245
rect 5805 10210 5845 10215
rect 6005 10315 6045 10320
rect 6005 10285 6010 10315
rect 6040 10285 6045 10315
rect 6005 10245 6045 10285
rect 6005 10215 6010 10245
rect 6040 10215 6045 10245
rect 6005 10210 6045 10215
rect 6205 10315 6245 10320
rect 6205 10285 6210 10315
rect 6240 10285 6245 10315
rect 6205 10245 6245 10285
rect 6205 10215 6210 10245
rect 6240 10215 6245 10245
rect 6205 10210 6245 10215
rect 6405 10315 6445 10320
rect 6405 10285 6410 10315
rect 6440 10285 6445 10315
rect 6405 10245 6445 10285
rect 6405 10215 6410 10245
rect 6440 10215 6445 10245
rect 6405 10210 6445 10215
rect -195 10130 -155 10135
rect -195 10100 -190 10130
rect -160 10100 -155 10130
rect -195 10060 -155 10100
rect -195 10030 -190 10060
rect -160 10030 -155 10060
rect -195 10025 -155 10030
rect 5 10130 45 10135
rect 5 10100 10 10130
rect 40 10100 45 10130
rect 5 10060 45 10100
rect 5 10030 10 10060
rect 40 10030 45 10060
rect 5 10025 45 10030
rect 205 10130 245 10135
rect 205 10100 210 10130
rect 240 10100 245 10130
rect 205 10060 245 10100
rect 205 10030 210 10060
rect 240 10030 245 10060
rect 205 10025 245 10030
rect 405 10130 445 10135
rect 405 10100 410 10130
rect 440 10100 445 10130
rect 405 10060 445 10100
rect 405 10030 410 10060
rect 440 10030 445 10060
rect 405 10025 445 10030
rect 605 10130 645 10135
rect 605 10100 610 10130
rect 640 10100 645 10130
rect 605 10060 645 10100
rect 605 10030 610 10060
rect 640 10030 645 10060
rect 605 10025 645 10030
rect 805 10130 845 10135
rect 805 10100 810 10130
rect 840 10100 845 10130
rect 805 10060 845 10100
rect 805 10030 810 10060
rect 840 10030 845 10060
rect 805 10025 845 10030
rect 1005 10130 1045 10135
rect 1005 10100 1010 10130
rect 1040 10100 1045 10130
rect 1005 10060 1045 10100
rect 1005 10030 1010 10060
rect 1040 10030 1045 10060
rect 1005 10025 1045 10030
rect 1205 10130 1245 10135
rect 1205 10100 1210 10130
rect 1240 10100 1245 10130
rect 1205 10060 1245 10100
rect 1205 10030 1210 10060
rect 1240 10030 1245 10060
rect 1205 10025 1245 10030
rect 1405 10130 1445 10135
rect 1405 10100 1410 10130
rect 1440 10100 1445 10130
rect 1405 10060 1445 10100
rect 1405 10030 1410 10060
rect 1440 10030 1445 10060
rect 1405 10025 1445 10030
rect 1605 10130 1645 10135
rect 1605 10100 1610 10130
rect 1640 10100 1645 10130
rect 1605 10060 1645 10100
rect 1605 10030 1610 10060
rect 1640 10030 1645 10060
rect 1605 10025 1645 10030
rect 1805 10130 1845 10135
rect 1805 10100 1810 10130
rect 1840 10100 1845 10130
rect 1805 10060 1845 10100
rect 1805 10030 1810 10060
rect 1840 10030 1845 10060
rect 1805 10025 1845 10030
rect 2005 10130 2045 10135
rect 2005 10100 2010 10130
rect 2040 10100 2045 10130
rect 2005 10060 2045 10100
rect 2005 10030 2010 10060
rect 2040 10030 2045 10060
rect 2005 10025 2045 10030
rect 2205 10130 2245 10135
rect 2205 10100 2210 10130
rect 2240 10100 2245 10130
rect 2205 10060 2245 10100
rect 2205 10030 2210 10060
rect 2240 10030 2245 10060
rect 2205 10025 2245 10030
rect 2405 10130 2445 10135
rect 2405 10100 2410 10130
rect 2440 10100 2445 10130
rect 2405 10060 2445 10100
rect 2405 10030 2410 10060
rect 2440 10030 2445 10060
rect 2405 10025 2445 10030
rect 2605 10130 2645 10135
rect 2605 10100 2610 10130
rect 2640 10100 2645 10130
rect 2605 10060 2645 10100
rect 2605 10030 2610 10060
rect 2640 10030 2645 10060
rect 2605 10025 2645 10030
rect 2805 10130 2845 10135
rect 2805 10100 2810 10130
rect 2840 10100 2845 10130
rect 2805 10060 2845 10100
rect 2805 10030 2810 10060
rect 2840 10030 2845 10060
rect 2805 10025 2845 10030
rect 3005 10130 3045 10135
rect 3005 10100 3010 10130
rect 3040 10100 3045 10130
rect 3005 10060 3045 10100
rect 3005 10030 3010 10060
rect 3040 10030 3045 10060
rect 3005 10025 3045 10030
rect 3205 10130 3245 10135
rect 3205 10100 3210 10130
rect 3240 10100 3245 10130
rect 3205 10060 3245 10100
rect 3205 10030 3210 10060
rect 3240 10030 3245 10060
rect 3205 10025 3245 10030
rect 3405 10130 3445 10135
rect 3405 10100 3410 10130
rect 3440 10100 3445 10130
rect 3405 10060 3445 10100
rect 3405 10030 3410 10060
rect 3440 10030 3445 10060
rect 3405 10025 3445 10030
rect 3605 10130 3645 10135
rect 3605 10100 3610 10130
rect 3640 10100 3645 10130
rect 3605 10060 3645 10100
rect 3605 10030 3610 10060
rect 3640 10030 3645 10060
rect 3605 10025 3645 10030
rect 3805 10130 3845 10135
rect 3805 10100 3810 10130
rect 3840 10100 3845 10130
rect 3805 10060 3845 10100
rect 3805 10030 3810 10060
rect 3840 10030 3845 10060
rect 3805 10025 3845 10030
rect 4005 10130 4045 10135
rect 4005 10100 4010 10130
rect 4040 10100 4045 10130
rect 4005 10060 4045 10100
rect 4005 10030 4010 10060
rect 4040 10030 4045 10060
rect 4005 10025 4045 10030
rect 4205 10130 4245 10135
rect 4205 10100 4210 10130
rect 4240 10100 4245 10130
rect 4205 10060 4245 10100
rect 4205 10030 4210 10060
rect 4240 10030 4245 10060
rect 4205 10025 4245 10030
rect 4405 10130 4445 10135
rect 4405 10100 4410 10130
rect 4440 10100 4445 10130
rect 4405 10060 4445 10100
rect 4405 10030 4410 10060
rect 4440 10030 4445 10060
rect 4405 10025 4445 10030
rect 4605 10130 4645 10135
rect 4605 10100 4610 10130
rect 4640 10100 4645 10130
rect 4605 10060 4645 10100
rect 4605 10030 4610 10060
rect 4640 10030 4645 10060
rect 4605 10025 4645 10030
rect 4805 10130 4845 10135
rect 4805 10100 4810 10130
rect 4840 10100 4845 10130
rect 4805 10060 4845 10100
rect 4805 10030 4810 10060
rect 4840 10030 4845 10060
rect 4805 10025 4845 10030
rect 5005 10130 5045 10135
rect 5005 10100 5010 10130
rect 5040 10100 5045 10130
rect 5005 10060 5045 10100
rect 5005 10030 5010 10060
rect 5040 10030 5045 10060
rect 5005 10025 5045 10030
rect 5205 10130 5245 10135
rect 5205 10100 5210 10130
rect 5240 10100 5245 10130
rect 5205 10060 5245 10100
rect 5205 10030 5210 10060
rect 5240 10030 5245 10060
rect 5205 10025 5245 10030
rect 5405 10130 5445 10135
rect 5405 10100 5410 10130
rect 5440 10100 5445 10130
rect 5405 10060 5445 10100
rect 5405 10030 5410 10060
rect 5440 10030 5445 10060
rect 5405 10025 5445 10030
rect 5605 10130 5645 10135
rect 5605 10100 5610 10130
rect 5640 10100 5645 10130
rect 5605 10060 5645 10100
rect 5605 10030 5610 10060
rect 5640 10030 5645 10060
rect 5605 10025 5645 10030
rect 5805 10130 5845 10135
rect 5805 10100 5810 10130
rect 5840 10100 5845 10130
rect 5805 10060 5845 10100
rect 5805 10030 5810 10060
rect 5840 10030 5845 10060
rect 5805 10025 5845 10030
rect 6005 10130 6045 10135
rect 6005 10100 6010 10130
rect 6040 10100 6045 10130
rect 6005 10060 6045 10100
rect 6005 10030 6010 10060
rect 6040 10030 6045 10060
rect 6005 10025 6045 10030
rect 6205 10130 6245 10135
rect 6205 10100 6210 10130
rect 6240 10100 6245 10130
rect 6205 10060 6245 10100
rect 6205 10030 6210 10060
rect 6240 10030 6245 10060
rect 6205 10025 6245 10030
rect 6405 10130 6445 10135
rect 6405 10100 6410 10130
rect 6440 10100 6445 10130
rect 6405 10060 6445 10100
rect 6405 10030 6410 10060
rect 6440 10030 6445 10060
rect 6405 10025 6445 10030
rect -195 9945 -155 9950
rect -195 9915 -190 9945
rect -160 9915 -155 9945
rect -195 9875 -155 9915
rect -195 9845 -190 9875
rect -160 9845 -155 9875
rect -195 9840 -155 9845
rect 5 9945 45 9950
rect 5 9915 10 9945
rect 40 9915 45 9945
rect 5 9875 45 9915
rect 5 9845 10 9875
rect 40 9845 45 9875
rect 5 9840 45 9845
rect 205 9945 245 9950
rect 205 9915 210 9945
rect 240 9915 245 9945
rect 205 9875 245 9915
rect 205 9845 210 9875
rect 240 9845 245 9875
rect 205 9840 245 9845
rect 405 9945 445 9950
rect 405 9915 410 9945
rect 440 9915 445 9945
rect 405 9875 445 9915
rect 405 9845 410 9875
rect 440 9845 445 9875
rect 405 9840 445 9845
rect 605 9945 645 9950
rect 605 9915 610 9945
rect 640 9915 645 9945
rect 605 9875 645 9915
rect 605 9845 610 9875
rect 640 9845 645 9875
rect 605 9840 645 9845
rect 805 9945 845 9950
rect 805 9915 810 9945
rect 840 9915 845 9945
rect 805 9875 845 9915
rect 805 9845 810 9875
rect 840 9845 845 9875
rect 805 9840 845 9845
rect 1005 9945 1045 9950
rect 1005 9915 1010 9945
rect 1040 9915 1045 9945
rect 1005 9875 1045 9915
rect 1005 9845 1010 9875
rect 1040 9845 1045 9875
rect 1005 9840 1045 9845
rect 1205 9945 1245 9950
rect 1205 9915 1210 9945
rect 1240 9915 1245 9945
rect 1205 9875 1245 9915
rect 1205 9845 1210 9875
rect 1240 9845 1245 9875
rect 1205 9840 1245 9845
rect 1405 9945 1445 9950
rect 1405 9915 1410 9945
rect 1440 9915 1445 9945
rect 1405 9875 1445 9915
rect 1405 9845 1410 9875
rect 1440 9845 1445 9875
rect 1405 9840 1445 9845
rect 1605 9945 1645 9950
rect 1605 9915 1610 9945
rect 1640 9915 1645 9945
rect 1605 9875 1645 9915
rect 1605 9845 1610 9875
rect 1640 9845 1645 9875
rect 1605 9840 1645 9845
rect 1805 9945 1845 9950
rect 1805 9915 1810 9945
rect 1840 9915 1845 9945
rect 1805 9875 1845 9915
rect 1805 9845 1810 9875
rect 1840 9845 1845 9875
rect 1805 9840 1845 9845
rect 2005 9945 2045 9950
rect 2005 9915 2010 9945
rect 2040 9915 2045 9945
rect 2005 9875 2045 9915
rect 2005 9845 2010 9875
rect 2040 9845 2045 9875
rect 2005 9840 2045 9845
rect 2205 9945 2245 9950
rect 2205 9915 2210 9945
rect 2240 9915 2245 9945
rect 2205 9875 2245 9915
rect 2205 9845 2210 9875
rect 2240 9845 2245 9875
rect 2205 9840 2245 9845
rect 2405 9945 2445 9950
rect 2405 9915 2410 9945
rect 2440 9915 2445 9945
rect 2405 9875 2445 9915
rect 2405 9845 2410 9875
rect 2440 9845 2445 9875
rect 2405 9840 2445 9845
rect 2605 9945 2645 9950
rect 2605 9915 2610 9945
rect 2640 9915 2645 9945
rect 2605 9875 2645 9915
rect 2605 9845 2610 9875
rect 2640 9845 2645 9875
rect 2605 9840 2645 9845
rect 2805 9945 2845 9950
rect 2805 9915 2810 9945
rect 2840 9915 2845 9945
rect 2805 9875 2845 9915
rect 2805 9845 2810 9875
rect 2840 9845 2845 9875
rect 2805 9840 2845 9845
rect 3005 9945 3045 9950
rect 3005 9915 3010 9945
rect 3040 9915 3045 9945
rect 3005 9875 3045 9915
rect 3005 9845 3010 9875
rect 3040 9845 3045 9875
rect 3005 9840 3045 9845
rect 3205 9945 3245 9950
rect 3205 9915 3210 9945
rect 3240 9915 3245 9945
rect 3205 9875 3245 9915
rect 3205 9845 3210 9875
rect 3240 9845 3245 9875
rect 3205 9840 3245 9845
rect 3405 9945 3445 9950
rect 3405 9915 3410 9945
rect 3440 9915 3445 9945
rect 3405 9875 3445 9915
rect 3405 9845 3410 9875
rect 3440 9845 3445 9875
rect 3405 9840 3445 9845
rect 3605 9945 3645 9950
rect 3605 9915 3610 9945
rect 3640 9915 3645 9945
rect 3605 9875 3645 9915
rect 3605 9845 3610 9875
rect 3640 9845 3645 9875
rect 3605 9840 3645 9845
rect 3805 9945 3845 9950
rect 3805 9915 3810 9945
rect 3840 9915 3845 9945
rect 3805 9875 3845 9915
rect 3805 9845 3810 9875
rect 3840 9845 3845 9875
rect 3805 9840 3845 9845
rect 4005 9945 4045 9950
rect 4005 9915 4010 9945
rect 4040 9915 4045 9945
rect 4005 9875 4045 9915
rect 4005 9845 4010 9875
rect 4040 9845 4045 9875
rect 4005 9840 4045 9845
rect 4205 9945 4245 9950
rect 4205 9915 4210 9945
rect 4240 9915 4245 9945
rect 4205 9875 4245 9915
rect 4205 9845 4210 9875
rect 4240 9845 4245 9875
rect 4205 9840 4245 9845
rect 4405 9945 4445 9950
rect 4405 9915 4410 9945
rect 4440 9915 4445 9945
rect 4405 9875 4445 9915
rect 4405 9845 4410 9875
rect 4440 9845 4445 9875
rect 4405 9840 4445 9845
rect 4605 9945 4645 9950
rect 4605 9915 4610 9945
rect 4640 9915 4645 9945
rect 4605 9875 4645 9915
rect 4605 9845 4610 9875
rect 4640 9845 4645 9875
rect 4605 9840 4645 9845
rect 4805 9945 4845 9950
rect 4805 9915 4810 9945
rect 4840 9915 4845 9945
rect 4805 9875 4845 9915
rect 4805 9845 4810 9875
rect 4840 9845 4845 9875
rect 4805 9840 4845 9845
rect 5005 9945 5045 9950
rect 5005 9915 5010 9945
rect 5040 9915 5045 9945
rect 5005 9875 5045 9915
rect 5005 9845 5010 9875
rect 5040 9845 5045 9875
rect 5005 9840 5045 9845
rect 5205 9945 5245 9950
rect 5205 9915 5210 9945
rect 5240 9915 5245 9945
rect 5205 9875 5245 9915
rect 5205 9845 5210 9875
rect 5240 9845 5245 9875
rect 5205 9840 5245 9845
rect 5405 9945 5445 9950
rect 5405 9915 5410 9945
rect 5440 9915 5445 9945
rect 5405 9875 5445 9915
rect 5405 9845 5410 9875
rect 5440 9845 5445 9875
rect 5405 9840 5445 9845
rect 5605 9945 5645 9950
rect 5605 9915 5610 9945
rect 5640 9915 5645 9945
rect 5605 9875 5645 9915
rect 5605 9845 5610 9875
rect 5640 9845 5645 9875
rect 5605 9840 5645 9845
rect 5805 9945 5845 9950
rect 5805 9915 5810 9945
rect 5840 9915 5845 9945
rect 5805 9875 5845 9915
rect 5805 9845 5810 9875
rect 5840 9845 5845 9875
rect 5805 9840 5845 9845
rect 6005 9945 6045 9950
rect 6005 9915 6010 9945
rect 6040 9915 6045 9945
rect 6005 9875 6045 9915
rect 6005 9845 6010 9875
rect 6040 9845 6045 9875
rect 6005 9840 6045 9845
rect 6205 9945 6245 9950
rect 6205 9915 6210 9945
rect 6240 9915 6245 9945
rect 6205 9875 6245 9915
rect 6205 9845 6210 9875
rect 6240 9845 6245 9875
rect 6205 9840 6245 9845
rect 6405 9945 6445 9950
rect 6405 9915 6410 9945
rect 6440 9915 6445 9945
rect 6405 9875 6445 9915
rect 6405 9845 6410 9875
rect 6440 9845 6445 9875
rect 6405 9840 6445 9845
rect -195 9760 -155 9765
rect -195 9730 -190 9760
rect -160 9730 -155 9760
rect -195 9690 -155 9730
rect -195 9660 -190 9690
rect -160 9660 -155 9690
rect -195 9655 -155 9660
rect 5 9760 45 9765
rect 5 9730 10 9760
rect 40 9730 45 9760
rect 5 9690 45 9730
rect 5 9660 10 9690
rect 40 9660 45 9690
rect 5 9655 45 9660
rect 205 9760 245 9765
rect 205 9730 210 9760
rect 240 9730 245 9760
rect 205 9690 245 9730
rect 205 9660 210 9690
rect 240 9660 245 9690
rect 205 9655 245 9660
rect 405 9760 445 9765
rect 405 9730 410 9760
rect 440 9730 445 9760
rect 405 9690 445 9730
rect 405 9660 410 9690
rect 440 9660 445 9690
rect 405 9655 445 9660
rect 605 9760 645 9765
rect 605 9730 610 9760
rect 640 9730 645 9760
rect 605 9690 645 9730
rect 605 9660 610 9690
rect 640 9660 645 9690
rect 605 9655 645 9660
rect 805 9760 845 9765
rect 805 9730 810 9760
rect 840 9730 845 9760
rect 805 9690 845 9730
rect 805 9660 810 9690
rect 840 9660 845 9690
rect 805 9655 845 9660
rect 1005 9760 1045 9765
rect 1005 9730 1010 9760
rect 1040 9730 1045 9760
rect 1005 9690 1045 9730
rect 1005 9660 1010 9690
rect 1040 9660 1045 9690
rect 1005 9655 1045 9660
rect 1205 9760 1245 9765
rect 1205 9730 1210 9760
rect 1240 9730 1245 9760
rect 1205 9690 1245 9730
rect 1205 9660 1210 9690
rect 1240 9660 1245 9690
rect 1205 9655 1245 9660
rect 1405 9760 1445 9765
rect 1405 9730 1410 9760
rect 1440 9730 1445 9760
rect 1405 9690 1445 9730
rect 1405 9660 1410 9690
rect 1440 9660 1445 9690
rect 1405 9655 1445 9660
rect 1605 9760 1645 9765
rect 1605 9730 1610 9760
rect 1640 9730 1645 9760
rect 1605 9690 1645 9730
rect 1605 9660 1610 9690
rect 1640 9660 1645 9690
rect 1605 9655 1645 9660
rect 1805 9760 1845 9765
rect 1805 9730 1810 9760
rect 1840 9730 1845 9760
rect 1805 9690 1845 9730
rect 1805 9660 1810 9690
rect 1840 9660 1845 9690
rect 1805 9655 1845 9660
rect 2005 9760 2045 9765
rect 2005 9730 2010 9760
rect 2040 9730 2045 9760
rect 2005 9690 2045 9730
rect 2005 9660 2010 9690
rect 2040 9660 2045 9690
rect 2005 9655 2045 9660
rect 2205 9760 2245 9765
rect 2205 9730 2210 9760
rect 2240 9730 2245 9760
rect 2205 9690 2245 9730
rect 2205 9660 2210 9690
rect 2240 9660 2245 9690
rect 2205 9655 2245 9660
rect 2405 9760 2445 9765
rect 2405 9730 2410 9760
rect 2440 9730 2445 9760
rect 2405 9690 2445 9730
rect 2405 9660 2410 9690
rect 2440 9660 2445 9690
rect 2405 9655 2445 9660
rect 2605 9760 2645 9765
rect 2605 9730 2610 9760
rect 2640 9730 2645 9760
rect 2605 9690 2645 9730
rect 2605 9660 2610 9690
rect 2640 9660 2645 9690
rect 2605 9655 2645 9660
rect 2805 9760 2845 9765
rect 2805 9730 2810 9760
rect 2840 9730 2845 9760
rect 2805 9690 2845 9730
rect 2805 9660 2810 9690
rect 2840 9660 2845 9690
rect 2805 9655 2845 9660
rect 3005 9760 3045 9765
rect 3005 9730 3010 9760
rect 3040 9730 3045 9760
rect 3005 9690 3045 9730
rect 3005 9660 3010 9690
rect 3040 9660 3045 9690
rect 3005 9655 3045 9660
rect 3205 9760 3245 9765
rect 3205 9730 3210 9760
rect 3240 9730 3245 9760
rect 3205 9690 3245 9730
rect 3205 9660 3210 9690
rect 3240 9660 3245 9690
rect 3205 9655 3245 9660
rect 3405 9760 3445 9765
rect 3405 9730 3410 9760
rect 3440 9730 3445 9760
rect 3405 9690 3445 9730
rect 3405 9660 3410 9690
rect 3440 9660 3445 9690
rect 3405 9655 3445 9660
rect 3605 9760 3645 9765
rect 3605 9730 3610 9760
rect 3640 9730 3645 9760
rect 3605 9690 3645 9730
rect 3605 9660 3610 9690
rect 3640 9660 3645 9690
rect 3605 9655 3645 9660
rect 3805 9760 3845 9765
rect 3805 9730 3810 9760
rect 3840 9730 3845 9760
rect 3805 9690 3845 9730
rect 3805 9660 3810 9690
rect 3840 9660 3845 9690
rect 3805 9655 3845 9660
rect 4005 9760 4045 9765
rect 4005 9730 4010 9760
rect 4040 9730 4045 9760
rect 4005 9690 4045 9730
rect 4005 9660 4010 9690
rect 4040 9660 4045 9690
rect 4005 9655 4045 9660
rect 4205 9760 4245 9765
rect 4205 9730 4210 9760
rect 4240 9730 4245 9760
rect 4205 9690 4245 9730
rect 4205 9660 4210 9690
rect 4240 9660 4245 9690
rect 4205 9655 4245 9660
rect 4405 9760 4445 9765
rect 4405 9730 4410 9760
rect 4440 9730 4445 9760
rect 4405 9690 4445 9730
rect 4405 9660 4410 9690
rect 4440 9660 4445 9690
rect 4405 9655 4445 9660
rect 4605 9760 4645 9765
rect 4605 9730 4610 9760
rect 4640 9730 4645 9760
rect 4605 9690 4645 9730
rect 4605 9660 4610 9690
rect 4640 9660 4645 9690
rect 4605 9655 4645 9660
rect 4805 9760 4845 9765
rect 4805 9730 4810 9760
rect 4840 9730 4845 9760
rect 4805 9690 4845 9730
rect 4805 9660 4810 9690
rect 4840 9660 4845 9690
rect 4805 9655 4845 9660
rect 5005 9760 5045 9765
rect 5005 9730 5010 9760
rect 5040 9730 5045 9760
rect 5005 9690 5045 9730
rect 5005 9660 5010 9690
rect 5040 9660 5045 9690
rect 5005 9655 5045 9660
rect 5205 9760 5245 9765
rect 5205 9730 5210 9760
rect 5240 9730 5245 9760
rect 5205 9690 5245 9730
rect 5205 9660 5210 9690
rect 5240 9660 5245 9690
rect 5205 9655 5245 9660
rect 5405 9760 5445 9765
rect 5405 9730 5410 9760
rect 5440 9730 5445 9760
rect 5405 9690 5445 9730
rect 5405 9660 5410 9690
rect 5440 9660 5445 9690
rect 5405 9655 5445 9660
rect 5605 9760 5645 9765
rect 5605 9730 5610 9760
rect 5640 9730 5645 9760
rect 5605 9690 5645 9730
rect 5605 9660 5610 9690
rect 5640 9660 5645 9690
rect 5605 9655 5645 9660
rect 5805 9760 5845 9765
rect 5805 9730 5810 9760
rect 5840 9730 5845 9760
rect 5805 9690 5845 9730
rect 5805 9660 5810 9690
rect 5840 9660 5845 9690
rect 5805 9655 5845 9660
rect 6005 9760 6045 9765
rect 6005 9730 6010 9760
rect 6040 9730 6045 9760
rect 6005 9690 6045 9730
rect 6005 9660 6010 9690
rect 6040 9660 6045 9690
rect 6005 9655 6045 9660
rect 6205 9760 6245 9765
rect 6205 9730 6210 9760
rect 6240 9730 6245 9760
rect 6205 9690 6245 9730
rect 6205 9660 6210 9690
rect 6240 9660 6245 9690
rect 6205 9655 6245 9660
rect 6405 9760 6445 9765
rect 6405 9730 6410 9760
rect 6440 9730 6445 9760
rect 6405 9690 6445 9730
rect 6405 9660 6410 9690
rect 6440 9660 6445 9690
rect 6405 9655 6445 9660
rect -195 9575 -155 9580
rect -195 9545 -190 9575
rect -160 9545 -155 9575
rect -195 9505 -155 9545
rect -195 9475 -190 9505
rect -160 9475 -155 9505
rect -195 9470 -155 9475
rect 5 9575 45 9580
rect 5 9545 10 9575
rect 40 9545 45 9575
rect 5 9505 45 9545
rect 5 9475 10 9505
rect 40 9475 45 9505
rect 5 9470 45 9475
rect 205 9575 245 9580
rect 205 9545 210 9575
rect 240 9545 245 9575
rect 205 9505 245 9545
rect 205 9475 210 9505
rect 240 9475 245 9505
rect 205 9470 245 9475
rect 405 9575 445 9580
rect 405 9545 410 9575
rect 440 9545 445 9575
rect 405 9505 445 9545
rect 405 9475 410 9505
rect 440 9475 445 9505
rect 405 9470 445 9475
rect 605 9575 645 9580
rect 605 9545 610 9575
rect 640 9545 645 9575
rect 605 9505 645 9545
rect 605 9475 610 9505
rect 640 9475 645 9505
rect 605 9470 645 9475
rect 805 9575 845 9580
rect 805 9545 810 9575
rect 840 9545 845 9575
rect 805 9505 845 9545
rect 805 9475 810 9505
rect 840 9475 845 9505
rect 805 9470 845 9475
rect 1005 9575 1045 9580
rect 1005 9545 1010 9575
rect 1040 9545 1045 9575
rect 1005 9505 1045 9545
rect 1005 9475 1010 9505
rect 1040 9475 1045 9505
rect 1005 9470 1045 9475
rect 1205 9575 1245 9580
rect 1205 9545 1210 9575
rect 1240 9545 1245 9575
rect 1205 9505 1245 9545
rect 1205 9475 1210 9505
rect 1240 9475 1245 9505
rect 1205 9470 1245 9475
rect 1405 9575 1445 9580
rect 1405 9545 1410 9575
rect 1440 9545 1445 9575
rect 1405 9505 1445 9545
rect 1405 9475 1410 9505
rect 1440 9475 1445 9505
rect 1405 9470 1445 9475
rect 1605 9575 1645 9580
rect 1605 9545 1610 9575
rect 1640 9545 1645 9575
rect 1605 9505 1645 9545
rect 1605 9475 1610 9505
rect 1640 9475 1645 9505
rect 1605 9470 1645 9475
rect 1805 9575 1845 9580
rect 1805 9545 1810 9575
rect 1840 9545 1845 9575
rect 1805 9505 1845 9545
rect 1805 9475 1810 9505
rect 1840 9475 1845 9505
rect 1805 9470 1845 9475
rect 2005 9575 2045 9580
rect 2005 9545 2010 9575
rect 2040 9545 2045 9575
rect 2005 9505 2045 9545
rect 2005 9475 2010 9505
rect 2040 9475 2045 9505
rect 2005 9470 2045 9475
rect 2205 9575 2245 9580
rect 2205 9545 2210 9575
rect 2240 9545 2245 9575
rect 2205 9505 2245 9545
rect 2205 9475 2210 9505
rect 2240 9475 2245 9505
rect 2205 9470 2245 9475
rect 2405 9575 2445 9580
rect 2405 9545 2410 9575
rect 2440 9545 2445 9575
rect 2405 9505 2445 9545
rect 2405 9475 2410 9505
rect 2440 9475 2445 9505
rect 2405 9470 2445 9475
rect 2605 9575 2645 9580
rect 2605 9545 2610 9575
rect 2640 9545 2645 9575
rect 2605 9505 2645 9545
rect 2605 9475 2610 9505
rect 2640 9475 2645 9505
rect 2605 9470 2645 9475
rect 2805 9575 2845 9580
rect 2805 9545 2810 9575
rect 2840 9545 2845 9575
rect 2805 9505 2845 9545
rect 2805 9475 2810 9505
rect 2840 9475 2845 9505
rect 2805 9470 2845 9475
rect 3005 9575 3045 9580
rect 3005 9545 3010 9575
rect 3040 9545 3045 9575
rect 3005 9505 3045 9545
rect 3005 9475 3010 9505
rect 3040 9475 3045 9505
rect 3005 9470 3045 9475
rect 3205 9575 3245 9580
rect 3205 9545 3210 9575
rect 3240 9545 3245 9575
rect 3205 9505 3245 9545
rect 3205 9475 3210 9505
rect 3240 9475 3245 9505
rect 3205 9470 3245 9475
rect 3405 9575 3445 9580
rect 3405 9545 3410 9575
rect 3440 9545 3445 9575
rect 3405 9505 3445 9545
rect 3405 9475 3410 9505
rect 3440 9475 3445 9505
rect 3405 9470 3445 9475
rect 3605 9575 3645 9580
rect 3605 9545 3610 9575
rect 3640 9545 3645 9575
rect 3605 9505 3645 9545
rect 3605 9475 3610 9505
rect 3640 9475 3645 9505
rect 3605 9470 3645 9475
rect 3805 9575 3845 9580
rect 3805 9545 3810 9575
rect 3840 9545 3845 9575
rect 3805 9505 3845 9545
rect 3805 9475 3810 9505
rect 3840 9475 3845 9505
rect 3805 9470 3845 9475
rect 4005 9575 4045 9580
rect 4005 9545 4010 9575
rect 4040 9545 4045 9575
rect 4005 9505 4045 9545
rect 4005 9475 4010 9505
rect 4040 9475 4045 9505
rect 4005 9470 4045 9475
rect 4205 9575 4245 9580
rect 4205 9545 4210 9575
rect 4240 9545 4245 9575
rect 4205 9505 4245 9545
rect 4205 9475 4210 9505
rect 4240 9475 4245 9505
rect 4205 9470 4245 9475
rect 4405 9575 4445 9580
rect 4405 9545 4410 9575
rect 4440 9545 4445 9575
rect 4405 9505 4445 9545
rect 4405 9475 4410 9505
rect 4440 9475 4445 9505
rect 4405 9470 4445 9475
rect 4605 9575 4645 9580
rect 4605 9545 4610 9575
rect 4640 9545 4645 9575
rect 4605 9505 4645 9545
rect 4605 9475 4610 9505
rect 4640 9475 4645 9505
rect 4605 9470 4645 9475
rect 4805 9575 4845 9580
rect 4805 9545 4810 9575
rect 4840 9545 4845 9575
rect 4805 9505 4845 9545
rect 4805 9475 4810 9505
rect 4840 9475 4845 9505
rect 4805 9470 4845 9475
rect 5005 9575 5045 9580
rect 5005 9545 5010 9575
rect 5040 9545 5045 9575
rect 5005 9505 5045 9545
rect 5005 9475 5010 9505
rect 5040 9475 5045 9505
rect 5005 9470 5045 9475
rect 5205 9575 5245 9580
rect 5205 9545 5210 9575
rect 5240 9545 5245 9575
rect 5205 9505 5245 9545
rect 5205 9475 5210 9505
rect 5240 9475 5245 9505
rect 5205 9470 5245 9475
rect 5405 9575 5445 9580
rect 5405 9545 5410 9575
rect 5440 9545 5445 9575
rect 5405 9505 5445 9545
rect 5405 9475 5410 9505
rect 5440 9475 5445 9505
rect 5405 9470 5445 9475
rect 5605 9575 5645 9580
rect 5605 9545 5610 9575
rect 5640 9545 5645 9575
rect 5605 9505 5645 9545
rect 5605 9475 5610 9505
rect 5640 9475 5645 9505
rect 5605 9470 5645 9475
rect 5805 9575 5845 9580
rect 5805 9545 5810 9575
rect 5840 9545 5845 9575
rect 5805 9505 5845 9545
rect 5805 9475 5810 9505
rect 5840 9475 5845 9505
rect 5805 9470 5845 9475
rect 6005 9575 6045 9580
rect 6005 9545 6010 9575
rect 6040 9545 6045 9575
rect 6005 9505 6045 9545
rect 6005 9475 6010 9505
rect 6040 9475 6045 9505
rect 6005 9470 6045 9475
rect 6205 9575 6245 9580
rect 6205 9545 6210 9575
rect 6240 9545 6245 9575
rect 6205 9505 6245 9545
rect 6205 9475 6210 9505
rect 6240 9475 6245 9505
rect 6205 9470 6245 9475
rect 6405 9575 6445 9580
rect 6405 9545 6410 9575
rect 6440 9545 6445 9575
rect 6405 9505 6445 9545
rect 6405 9475 6410 9505
rect 6440 9475 6445 9505
rect 6405 9470 6445 9475
rect -195 9390 -155 9395
rect -195 9360 -190 9390
rect -160 9360 -155 9390
rect -195 9320 -155 9360
rect -195 9290 -190 9320
rect -160 9290 -155 9320
rect -195 9285 -155 9290
rect 5 9390 45 9395
rect 5 9360 10 9390
rect 40 9360 45 9390
rect 5 9320 45 9360
rect 5 9290 10 9320
rect 40 9290 45 9320
rect 5 9285 45 9290
rect 205 9390 245 9395
rect 205 9360 210 9390
rect 240 9360 245 9390
rect 205 9320 245 9360
rect 205 9290 210 9320
rect 240 9290 245 9320
rect 205 9285 245 9290
rect 405 9390 445 9395
rect 405 9360 410 9390
rect 440 9360 445 9390
rect 405 9320 445 9360
rect 405 9290 410 9320
rect 440 9290 445 9320
rect 405 9285 445 9290
rect 605 9390 645 9395
rect 605 9360 610 9390
rect 640 9360 645 9390
rect 605 9320 645 9360
rect 605 9290 610 9320
rect 640 9290 645 9320
rect 605 9285 645 9290
rect 805 9390 845 9395
rect 805 9360 810 9390
rect 840 9360 845 9390
rect 805 9320 845 9360
rect 805 9290 810 9320
rect 840 9290 845 9320
rect 805 9285 845 9290
rect 1005 9390 1045 9395
rect 1005 9360 1010 9390
rect 1040 9360 1045 9390
rect 1005 9320 1045 9360
rect 1005 9290 1010 9320
rect 1040 9290 1045 9320
rect 1005 9285 1045 9290
rect 1205 9390 1245 9395
rect 1205 9360 1210 9390
rect 1240 9360 1245 9390
rect 1205 9320 1245 9360
rect 1205 9290 1210 9320
rect 1240 9290 1245 9320
rect 1205 9285 1245 9290
rect 1405 9390 1445 9395
rect 1405 9360 1410 9390
rect 1440 9360 1445 9390
rect 1405 9320 1445 9360
rect 1405 9290 1410 9320
rect 1440 9290 1445 9320
rect 1405 9285 1445 9290
rect 1605 9390 1645 9395
rect 1605 9360 1610 9390
rect 1640 9360 1645 9390
rect 1605 9320 1645 9360
rect 1605 9290 1610 9320
rect 1640 9290 1645 9320
rect 1605 9285 1645 9290
rect 1805 9390 1845 9395
rect 1805 9360 1810 9390
rect 1840 9360 1845 9390
rect 1805 9320 1845 9360
rect 1805 9290 1810 9320
rect 1840 9290 1845 9320
rect 1805 9285 1845 9290
rect 2005 9390 2045 9395
rect 2005 9360 2010 9390
rect 2040 9360 2045 9390
rect 2005 9320 2045 9360
rect 2005 9290 2010 9320
rect 2040 9290 2045 9320
rect 2005 9285 2045 9290
rect 2205 9390 2245 9395
rect 2205 9360 2210 9390
rect 2240 9360 2245 9390
rect 2205 9320 2245 9360
rect 2205 9290 2210 9320
rect 2240 9290 2245 9320
rect 2205 9285 2245 9290
rect 2405 9390 2445 9395
rect 2405 9360 2410 9390
rect 2440 9360 2445 9390
rect 2405 9320 2445 9360
rect 2405 9290 2410 9320
rect 2440 9290 2445 9320
rect 2405 9285 2445 9290
rect 2605 9390 2645 9395
rect 2605 9360 2610 9390
rect 2640 9360 2645 9390
rect 2605 9320 2645 9360
rect 2605 9290 2610 9320
rect 2640 9290 2645 9320
rect 2605 9285 2645 9290
rect 2805 9390 2845 9395
rect 2805 9360 2810 9390
rect 2840 9360 2845 9390
rect 2805 9320 2845 9360
rect 2805 9290 2810 9320
rect 2840 9290 2845 9320
rect 2805 9285 2845 9290
rect 3005 9390 3045 9395
rect 3005 9360 3010 9390
rect 3040 9360 3045 9390
rect 3005 9320 3045 9360
rect 3005 9290 3010 9320
rect 3040 9290 3045 9320
rect 3005 9285 3045 9290
rect 3205 9390 3245 9395
rect 3205 9360 3210 9390
rect 3240 9360 3245 9390
rect 3205 9320 3245 9360
rect 3205 9290 3210 9320
rect 3240 9290 3245 9320
rect 3205 9285 3245 9290
rect 3405 9390 3445 9395
rect 3405 9360 3410 9390
rect 3440 9360 3445 9390
rect 3405 9320 3445 9360
rect 3405 9290 3410 9320
rect 3440 9290 3445 9320
rect 3405 9285 3445 9290
rect 3605 9390 3645 9395
rect 3605 9360 3610 9390
rect 3640 9360 3645 9390
rect 3605 9320 3645 9360
rect 3605 9290 3610 9320
rect 3640 9290 3645 9320
rect 3605 9285 3645 9290
rect 3805 9390 3845 9395
rect 3805 9360 3810 9390
rect 3840 9360 3845 9390
rect 3805 9320 3845 9360
rect 3805 9290 3810 9320
rect 3840 9290 3845 9320
rect 3805 9285 3845 9290
rect 4005 9390 4045 9395
rect 4005 9360 4010 9390
rect 4040 9360 4045 9390
rect 4005 9320 4045 9360
rect 4005 9290 4010 9320
rect 4040 9290 4045 9320
rect 4005 9285 4045 9290
rect 4205 9390 4245 9395
rect 4205 9360 4210 9390
rect 4240 9360 4245 9390
rect 4205 9320 4245 9360
rect 4205 9290 4210 9320
rect 4240 9290 4245 9320
rect 4205 9285 4245 9290
rect 4405 9390 4445 9395
rect 4405 9360 4410 9390
rect 4440 9360 4445 9390
rect 4405 9320 4445 9360
rect 4405 9290 4410 9320
rect 4440 9290 4445 9320
rect 4405 9285 4445 9290
rect 4605 9390 4645 9395
rect 4605 9360 4610 9390
rect 4640 9360 4645 9390
rect 4605 9320 4645 9360
rect 4605 9290 4610 9320
rect 4640 9290 4645 9320
rect 4605 9285 4645 9290
rect 4805 9390 4845 9395
rect 4805 9360 4810 9390
rect 4840 9360 4845 9390
rect 4805 9320 4845 9360
rect 4805 9290 4810 9320
rect 4840 9290 4845 9320
rect 4805 9285 4845 9290
rect 5005 9390 5045 9395
rect 5005 9360 5010 9390
rect 5040 9360 5045 9390
rect 5005 9320 5045 9360
rect 5005 9290 5010 9320
rect 5040 9290 5045 9320
rect 5005 9285 5045 9290
rect 5205 9390 5245 9395
rect 5205 9360 5210 9390
rect 5240 9360 5245 9390
rect 5205 9320 5245 9360
rect 5205 9290 5210 9320
rect 5240 9290 5245 9320
rect 5205 9285 5245 9290
rect 5405 9390 5445 9395
rect 5405 9360 5410 9390
rect 5440 9360 5445 9390
rect 5405 9320 5445 9360
rect 5405 9290 5410 9320
rect 5440 9290 5445 9320
rect 5405 9285 5445 9290
rect 5605 9390 5645 9395
rect 5605 9360 5610 9390
rect 5640 9360 5645 9390
rect 5605 9320 5645 9360
rect 5605 9290 5610 9320
rect 5640 9290 5645 9320
rect 5605 9285 5645 9290
rect 5805 9390 5845 9395
rect 5805 9360 5810 9390
rect 5840 9360 5845 9390
rect 5805 9320 5845 9360
rect 5805 9290 5810 9320
rect 5840 9290 5845 9320
rect 5805 9285 5845 9290
rect 6005 9390 6045 9395
rect 6005 9360 6010 9390
rect 6040 9360 6045 9390
rect 6005 9320 6045 9360
rect 6005 9290 6010 9320
rect 6040 9290 6045 9320
rect 6005 9285 6045 9290
rect 6205 9390 6245 9395
rect 6205 9360 6210 9390
rect 6240 9360 6245 9390
rect 6205 9320 6245 9360
rect 6205 9290 6210 9320
rect 6240 9290 6245 9320
rect 6205 9285 6245 9290
rect 6405 9390 6445 9395
rect 6405 9360 6410 9390
rect 6440 9360 6445 9390
rect 6405 9320 6445 9360
rect 6405 9290 6410 9320
rect 6440 9290 6445 9320
rect 6405 9285 6445 9290
rect -195 9205 -155 9210
rect -195 9175 -190 9205
rect -160 9175 -155 9205
rect -195 9135 -155 9175
rect -195 9105 -190 9135
rect -160 9105 -155 9135
rect -195 9100 -155 9105
rect 5 9205 45 9210
rect 5 9175 10 9205
rect 40 9175 45 9205
rect 5 9135 45 9175
rect 5 9105 10 9135
rect 40 9105 45 9135
rect 5 9100 45 9105
rect 205 9205 245 9210
rect 205 9175 210 9205
rect 240 9175 245 9205
rect 205 9135 245 9175
rect 205 9105 210 9135
rect 240 9105 245 9135
rect 205 9100 245 9105
rect 405 9205 445 9210
rect 405 9175 410 9205
rect 440 9175 445 9205
rect 405 9135 445 9175
rect 405 9105 410 9135
rect 440 9105 445 9135
rect 405 9100 445 9105
rect 605 9205 645 9210
rect 605 9175 610 9205
rect 640 9175 645 9205
rect 605 9135 645 9175
rect 605 9105 610 9135
rect 640 9105 645 9135
rect 605 9100 645 9105
rect 805 9205 845 9210
rect 805 9175 810 9205
rect 840 9175 845 9205
rect 805 9135 845 9175
rect 805 9105 810 9135
rect 840 9105 845 9135
rect 805 9100 845 9105
rect 1005 9205 1045 9210
rect 1005 9175 1010 9205
rect 1040 9175 1045 9205
rect 1005 9135 1045 9175
rect 1005 9105 1010 9135
rect 1040 9105 1045 9135
rect 1005 9100 1045 9105
rect 1205 9205 1245 9210
rect 1205 9175 1210 9205
rect 1240 9175 1245 9205
rect 1205 9135 1245 9175
rect 1205 9105 1210 9135
rect 1240 9105 1245 9135
rect 1205 9100 1245 9105
rect 1405 9205 1445 9210
rect 1405 9175 1410 9205
rect 1440 9175 1445 9205
rect 1405 9135 1445 9175
rect 1405 9105 1410 9135
rect 1440 9105 1445 9135
rect 1405 9100 1445 9105
rect 1605 9205 1645 9210
rect 1605 9175 1610 9205
rect 1640 9175 1645 9205
rect 1605 9135 1645 9175
rect 1605 9105 1610 9135
rect 1640 9105 1645 9135
rect 1605 9100 1645 9105
rect 1805 9205 1845 9210
rect 1805 9175 1810 9205
rect 1840 9175 1845 9205
rect 1805 9135 1845 9175
rect 1805 9105 1810 9135
rect 1840 9105 1845 9135
rect 1805 9100 1845 9105
rect 2005 9205 2045 9210
rect 2005 9175 2010 9205
rect 2040 9175 2045 9205
rect 2005 9135 2045 9175
rect 2005 9105 2010 9135
rect 2040 9105 2045 9135
rect 2005 9100 2045 9105
rect 2205 9205 2245 9210
rect 2205 9175 2210 9205
rect 2240 9175 2245 9205
rect 2205 9135 2245 9175
rect 2205 9105 2210 9135
rect 2240 9105 2245 9135
rect 2205 9100 2245 9105
rect 2405 9205 2445 9210
rect 2405 9175 2410 9205
rect 2440 9175 2445 9205
rect 2405 9135 2445 9175
rect 2405 9105 2410 9135
rect 2440 9105 2445 9135
rect 2405 9100 2445 9105
rect 2605 9205 2645 9210
rect 2605 9175 2610 9205
rect 2640 9175 2645 9205
rect 2605 9135 2645 9175
rect 2605 9105 2610 9135
rect 2640 9105 2645 9135
rect 2605 9100 2645 9105
rect 2805 9205 2845 9210
rect 2805 9175 2810 9205
rect 2840 9175 2845 9205
rect 2805 9135 2845 9175
rect 2805 9105 2810 9135
rect 2840 9105 2845 9135
rect 2805 9100 2845 9105
rect 3005 9205 3045 9210
rect 3005 9175 3010 9205
rect 3040 9175 3045 9205
rect 3005 9135 3045 9175
rect 3005 9105 3010 9135
rect 3040 9105 3045 9135
rect 3005 9100 3045 9105
rect 3205 9205 3245 9210
rect 3205 9175 3210 9205
rect 3240 9175 3245 9205
rect 3205 9135 3245 9175
rect 3205 9105 3210 9135
rect 3240 9105 3245 9135
rect 3205 9100 3245 9105
rect 3405 9205 3445 9210
rect 3405 9175 3410 9205
rect 3440 9175 3445 9205
rect 3405 9135 3445 9175
rect 3405 9105 3410 9135
rect 3440 9105 3445 9135
rect 3405 9100 3445 9105
rect 3605 9205 3645 9210
rect 3605 9175 3610 9205
rect 3640 9175 3645 9205
rect 3605 9135 3645 9175
rect 3605 9105 3610 9135
rect 3640 9105 3645 9135
rect 3605 9100 3645 9105
rect 3805 9205 3845 9210
rect 3805 9175 3810 9205
rect 3840 9175 3845 9205
rect 3805 9135 3845 9175
rect 3805 9105 3810 9135
rect 3840 9105 3845 9135
rect 3805 9100 3845 9105
rect 4005 9205 4045 9210
rect 4005 9175 4010 9205
rect 4040 9175 4045 9205
rect 4005 9135 4045 9175
rect 4005 9105 4010 9135
rect 4040 9105 4045 9135
rect 4005 9100 4045 9105
rect 4205 9205 4245 9210
rect 4205 9175 4210 9205
rect 4240 9175 4245 9205
rect 4205 9135 4245 9175
rect 4205 9105 4210 9135
rect 4240 9105 4245 9135
rect 4205 9100 4245 9105
rect 4405 9205 4445 9210
rect 4405 9175 4410 9205
rect 4440 9175 4445 9205
rect 4405 9135 4445 9175
rect 4405 9105 4410 9135
rect 4440 9105 4445 9135
rect 4405 9100 4445 9105
rect 4605 9205 4645 9210
rect 4605 9175 4610 9205
rect 4640 9175 4645 9205
rect 4605 9135 4645 9175
rect 4605 9105 4610 9135
rect 4640 9105 4645 9135
rect 4605 9100 4645 9105
rect 4805 9205 4845 9210
rect 4805 9175 4810 9205
rect 4840 9175 4845 9205
rect 4805 9135 4845 9175
rect 4805 9105 4810 9135
rect 4840 9105 4845 9135
rect 4805 9100 4845 9105
rect 5005 9205 5045 9210
rect 5005 9175 5010 9205
rect 5040 9175 5045 9205
rect 5005 9135 5045 9175
rect 5005 9105 5010 9135
rect 5040 9105 5045 9135
rect 5005 9100 5045 9105
rect 5205 9205 5245 9210
rect 5205 9175 5210 9205
rect 5240 9175 5245 9205
rect 5205 9135 5245 9175
rect 5205 9105 5210 9135
rect 5240 9105 5245 9135
rect 5205 9100 5245 9105
rect 5405 9205 5445 9210
rect 5405 9175 5410 9205
rect 5440 9175 5445 9205
rect 5405 9135 5445 9175
rect 5405 9105 5410 9135
rect 5440 9105 5445 9135
rect 5405 9100 5445 9105
rect 5605 9205 5645 9210
rect 5605 9175 5610 9205
rect 5640 9175 5645 9205
rect 5605 9135 5645 9175
rect 5605 9105 5610 9135
rect 5640 9105 5645 9135
rect 5605 9100 5645 9105
rect 5805 9205 5845 9210
rect 5805 9175 5810 9205
rect 5840 9175 5845 9205
rect 5805 9135 5845 9175
rect 5805 9105 5810 9135
rect 5840 9105 5845 9135
rect 5805 9100 5845 9105
rect 6005 9205 6045 9210
rect 6005 9175 6010 9205
rect 6040 9175 6045 9205
rect 6005 9135 6045 9175
rect 6005 9105 6010 9135
rect 6040 9105 6045 9135
rect 6005 9100 6045 9105
rect 6205 9205 6245 9210
rect 6205 9175 6210 9205
rect 6240 9175 6245 9205
rect 6205 9135 6245 9175
rect 6205 9105 6210 9135
rect 6240 9105 6245 9135
rect 6205 9100 6245 9105
rect 6405 9205 6445 9210
rect 6405 9175 6410 9205
rect 6440 9175 6445 9205
rect 6405 9135 6445 9175
rect 6405 9105 6410 9135
rect 6440 9105 6445 9135
rect 6405 9100 6445 9105
rect -195 9020 -155 9025
rect -195 8990 -190 9020
rect -160 8990 -155 9020
rect -195 8950 -155 8990
rect -195 8920 -190 8950
rect -160 8920 -155 8950
rect -195 8915 -155 8920
rect 5 9020 45 9025
rect 5 8990 10 9020
rect 40 8990 45 9020
rect 5 8950 45 8990
rect 5 8920 10 8950
rect 40 8920 45 8950
rect 5 8915 45 8920
rect 205 9020 245 9025
rect 205 8990 210 9020
rect 240 8990 245 9020
rect 205 8950 245 8990
rect 205 8920 210 8950
rect 240 8920 245 8950
rect 205 8915 245 8920
rect 405 9020 445 9025
rect 405 8990 410 9020
rect 440 8990 445 9020
rect 405 8950 445 8990
rect 405 8920 410 8950
rect 440 8920 445 8950
rect 405 8915 445 8920
rect 605 9020 645 9025
rect 605 8990 610 9020
rect 640 8990 645 9020
rect 605 8950 645 8990
rect 605 8920 610 8950
rect 640 8920 645 8950
rect 605 8915 645 8920
rect 805 9020 845 9025
rect 805 8990 810 9020
rect 840 8990 845 9020
rect 805 8950 845 8990
rect 805 8920 810 8950
rect 840 8920 845 8950
rect 805 8915 845 8920
rect 1005 9020 1045 9025
rect 1005 8990 1010 9020
rect 1040 8990 1045 9020
rect 1005 8950 1045 8990
rect 1005 8920 1010 8950
rect 1040 8920 1045 8950
rect 1005 8915 1045 8920
rect 1205 9020 1245 9025
rect 1205 8990 1210 9020
rect 1240 8990 1245 9020
rect 1205 8950 1245 8990
rect 1205 8920 1210 8950
rect 1240 8920 1245 8950
rect 1205 8915 1245 8920
rect 1405 9020 1445 9025
rect 1405 8990 1410 9020
rect 1440 8990 1445 9020
rect 1405 8950 1445 8990
rect 1405 8920 1410 8950
rect 1440 8920 1445 8950
rect 1405 8915 1445 8920
rect 1605 9020 1645 9025
rect 1605 8990 1610 9020
rect 1640 8990 1645 9020
rect 1605 8950 1645 8990
rect 1605 8920 1610 8950
rect 1640 8920 1645 8950
rect 1605 8915 1645 8920
rect 1805 9020 1845 9025
rect 1805 8990 1810 9020
rect 1840 8990 1845 9020
rect 1805 8950 1845 8990
rect 1805 8920 1810 8950
rect 1840 8920 1845 8950
rect 1805 8915 1845 8920
rect 2005 9020 2045 9025
rect 2005 8990 2010 9020
rect 2040 8990 2045 9020
rect 2005 8950 2045 8990
rect 2005 8920 2010 8950
rect 2040 8920 2045 8950
rect 2005 8915 2045 8920
rect 2205 9020 2245 9025
rect 2205 8990 2210 9020
rect 2240 8990 2245 9020
rect 2205 8950 2245 8990
rect 2205 8920 2210 8950
rect 2240 8920 2245 8950
rect 2205 8915 2245 8920
rect 2405 9020 2445 9025
rect 2405 8990 2410 9020
rect 2440 8990 2445 9020
rect 2405 8950 2445 8990
rect 2405 8920 2410 8950
rect 2440 8920 2445 8950
rect 2405 8915 2445 8920
rect 2605 9020 2645 9025
rect 2605 8990 2610 9020
rect 2640 8990 2645 9020
rect 2605 8950 2645 8990
rect 2605 8920 2610 8950
rect 2640 8920 2645 8950
rect 2605 8915 2645 8920
rect 2805 9020 2845 9025
rect 2805 8990 2810 9020
rect 2840 8990 2845 9020
rect 2805 8950 2845 8990
rect 2805 8920 2810 8950
rect 2840 8920 2845 8950
rect 2805 8915 2845 8920
rect 3005 9020 3045 9025
rect 3005 8990 3010 9020
rect 3040 8990 3045 9020
rect 3005 8950 3045 8990
rect 3005 8920 3010 8950
rect 3040 8920 3045 8950
rect 3005 8915 3045 8920
rect 3205 9020 3245 9025
rect 3205 8990 3210 9020
rect 3240 8990 3245 9020
rect 3205 8950 3245 8990
rect 3205 8920 3210 8950
rect 3240 8920 3245 8950
rect 3205 8915 3245 8920
rect 3405 9020 3445 9025
rect 3405 8990 3410 9020
rect 3440 8990 3445 9020
rect 3405 8950 3445 8990
rect 3405 8920 3410 8950
rect 3440 8920 3445 8950
rect 3405 8915 3445 8920
rect 3605 9020 3645 9025
rect 3605 8990 3610 9020
rect 3640 8990 3645 9020
rect 3605 8950 3645 8990
rect 3605 8920 3610 8950
rect 3640 8920 3645 8950
rect 3605 8915 3645 8920
rect 3805 9020 3845 9025
rect 3805 8990 3810 9020
rect 3840 8990 3845 9020
rect 3805 8950 3845 8990
rect 3805 8920 3810 8950
rect 3840 8920 3845 8950
rect 3805 8915 3845 8920
rect 4005 9020 4045 9025
rect 4005 8990 4010 9020
rect 4040 8990 4045 9020
rect 4005 8950 4045 8990
rect 4005 8920 4010 8950
rect 4040 8920 4045 8950
rect 4005 8915 4045 8920
rect 4205 9020 4245 9025
rect 4205 8990 4210 9020
rect 4240 8990 4245 9020
rect 4205 8950 4245 8990
rect 4205 8920 4210 8950
rect 4240 8920 4245 8950
rect 4205 8915 4245 8920
rect 4405 9020 4445 9025
rect 4405 8990 4410 9020
rect 4440 8990 4445 9020
rect 4405 8950 4445 8990
rect 4405 8920 4410 8950
rect 4440 8920 4445 8950
rect 4405 8915 4445 8920
rect 4605 9020 4645 9025
rect 4605 8990 4610 9020
rect 4640 8990 4645 9020
rect 4605 8950 4645 8990
rect 4605 8920 4610 8950
rect 4640 8920 4645 8950
rect 4605 8915 4645 8920
rect 4805 9020 4845 9025
rect 4805 8990 4810 9020
rect 4840 8990 4845 9020
rect 4805 8950 4845 8990
rect 4805 8920 4810 8950
rect 4840 8920 4845 8950
rect 4805 8915 4845 8920
rect 5005 9020 5045 9025
rect 5005 8990 5010 9020
rect 5040 8990 5045 9020
rect 5005 8950 5045 8990
rect 5005 8920 5010 8950
rect 5040 8920 5045 8950
rect 5005 8915 5045 8920
rect 5205 9020 5245 9025
rect 5205 8990 5210 9020
rect 5240 8990 5245 9020
rect 5205 8950 5245 8990
rect 5205 8920 5210 8950
rect 5240 8920 5245 8950
rect 5205 8915 5245 8920
rect 5405 9020 5445 9025
rect 5405 8990 5410 9020
rect 5440 8990 5445 9020
rect 5405 8950 5445 8990
rect 5405 8920 5410 8950
rect 5440 8920 5445 8950
rect 5405 8915 5445 8920
rect 5605 9020 5645 9025
rect 5605 8990 5610 9020
rect 5640 8990 5645 9020
rect 5605 8950 5645 8990
rect 5605 8920 5610 8950
rect 5640 8920 5645 8950
rect 5605 8915 5645 8920
rect 5805 9020 5845 9025
rect 5805 8990 5810 9020
rect 5840 8990 5845 9020
rect 5805 8950 5845 8990
rect 5805 8920 5810 8950
rect 5840 8920 5845 8950
rect 5805 8915 5845 8920
rect 6005 9020 6045 9025
rect 6005 8990 6010 9020
rect 6040 8990 6045 9020
rect 6005 8950 6045 8990
rect 6005 8920 6010 8950
rect 6040 8920 6045 8950
rect 6005 8915 6045 8920
rect 6205 9020 6245 9025
rect 6205 8990 6210 9020
rect 6240 8990 6245 9020
rect 6205 8950 6245 8990
rect 6205 8920 6210 8950
rect 6240 8920 6245 8950
rect 6205 8915 6245 8920
rect 6405 9020 6445 9025
rect 6405 8990 6410 9020
rect 6440 8990 6445 9020
rect 6405 8950 6445 8990
rect 6405 8920 6410 8950
rect 6440 8920 6445 8950
rect 6405 8915 6445 8920
rect -195 8835 -155 8840
rect -195 8805 -190 8835
rect -160 8805 -155 8835
rect -195 8765 -155 8805
rect -195 8735 -190 8765
rect -160 8735 -155 8765
rect -195 8730 -155 8735
rect 5 8835 45 8840
rect 5 8805 10 8835
rect 40 8805 45 8835
rect 5 8765 45 8805
rect 5 8735 10 8765
rect 40 8735 45 8765
rect 5 8730 45 8735
rect 205 8835 245 8840
rect 205 8805 210 8835
rect 240 8805 245 8835
rect 205 8765 245 8805
rect 205 8735 210 8765
rect 240 8735 245 8765
rect 205 8730 245 8735
rect 405 8835 445 8840
rect 405 8805 410 8835
rect 440 8805 445 8835
rect 405 8765 445 8805
rect 405 8735 410 8765
rect 440 8735 445 8765
rect 405 8730 445 8735
rect 605 8835 645 8840
rect 605 8805 610 8835
rect 640 8805 645 8835
rect 605 8765 645 8805
rect 605 8735 610 8765
rect 640 8735 645 8765
rect 605 8730 645 8735
rect 805 8835 845 8840
rect 805 8805 810 8835
rect 840 8805 845 8835
rect 805 8765 845 8805
rect 805 8735 810 8765
rect 840 8735 845 8765
rect 805 8730 845 8735
rect 1005 8835 1045 8840
rect 1005 8805 1010 8835
rect 1040 8805 1045 8835
rect 1005 8765 1045 8805
rect 1005 8735 1010 8765
rect 1040 8735 1045 8765
rect 1005 8730 1045 8735
rect 1205 8835 1245 8840
rect 1205 8805 1210 8835
rect 1240 8805 1245 8835
rect 1205 8765 1245 8805
rect 1205 8735 1210 8765
rect 1240 8735 1245 8765
rect 1205 8730 1245 8735
rect 1405 8835 1445 8840
rect 1405 8805 1410 8835
rect 1440 8805 1445 8835
rect 1405 8765 1445 8805
rect 1405 8735 1410 8765
rect 1440 8735 1445 8765
rect 1405 8730 1445 8735
rect 1605 8835 1645 8840
rect 1605 8805 1610 8835
rect 1640 8805 1645 8835
rect 1605 8765 1645 8805
rect 1605 8735 1610 8765
rect 1640 8735 1645 8765
rect 1605 8730 1645 8735
rect 1805 8835 1845 8840
rect 1805 8805 1810 8835
rect 1840 8805 1845 8835
rect 1805 8765 1845 8805
rect 1805 8735 1810 8765
rect 1840 8735 1845 8765
rect 1805 8730 1845 8735
rect 2005 8835 2045 8840
rect 2005 8805 2010 8835
rect 2040 8805 2045 8835
rect 2005 8765 2045 8805
rect 2005 8735 2010 8765
rect 2040 8735 2045 8765
rect 2005 8730 2045 8735
rect 2205 8835 2245 8840
rect 2205 8805 2210 8835
rect 2240 8805 2245 8835
rect 2205 8765 2245 8805
rect 2205 8735 2210 8765
rect 2240 8735 2245 8765
rect 2205 8730 2245 8735
rect 2405 8835 2445 8840
rect 2405 8805 2410 8835
rect 2440 8805 2445 8835
rect 2405 8765 2445 8805
rect 2405 8735 2410 8765
rect 2440 8735 2445 8765
rect 2405 8730 2445 8735
rect 2605 8835 2645 8840
rect 2605 8805 2610 8835
rect 2640 8805 2645 8835
rect 2605 8765 2645 8805
rect 2605 8735 2610 8765
rect 2640 8735 2645 8765
rect 2605 8730 2645 8735
rect 2805 8835 2845 8840
rect 2805 8805 2810 8835
rect 2840 8805 2845 8835
rect 2805 8765 2845 8805
rect 2805 8735 2810 8765
rect 2840 8735 2845 8765
rect 2805 8730 2845 8735
rect 3005 8835 3045 8840
rect 3005 8805 3010 8835
rect 3040 8805 3045 8835
rect 3005 8765 3045 8805
rect 3005 8735 3010 8765
rect 3040 8735 3045 8765
rect 3005 8730 3045 8735
rect 3205 8835 3245 8840
rect 3205 8805 3210 8835
rect 3240 8805 3245 8835
rect 3205 8765 3245 8805
rect 3205 8735 3210 8765
rect 3240 8735 3245 8765
rect 3205 8730 3245 8735
rect 3405 8835 3445 8840
rect 3405 8805 3410 8835
rect 3440 8805 3445 8835
rect 3405 8765 3445 8805
rect 3405 8735 3410 8765
rect 3440 8735 3445 8765
rect 3405 8730 3445 8735
rect 3605 8835 3645 8840
rect 3605 8805 3610 8835
rect 3640 8805 3645 8835
rect 3605 8765 3645 8805
rect 3605 8735 3610 8765
rect 3640 8735 3645 8765
rect 3605 8730 3645 8735
rect 3805 8835 3845 8840
rect 3805 8805 3810 8835
rect 3840 8805 3845 8835
rect 3805 8765 3845 8805
rect 3805 8735 3810 8765
rect 3840 8735 3845 8765
rect 3805 8730 3845 8735
rect 4005 8835 4045 8840
rect 4005 8805 4010 8835
rect 4040 8805 4045 8835
rect 4005 8765 4045 8805
rect 4005 8735 4010 8765
rect 4040 8735 4045 8765
rect 4005 8730 4045 8735
rect 4205 8835 4245 8840
rect 4205 8805 4210 8835
rect 4240 8805 4245 8835
rect 4205 8765 4245 8805
rect 4205 8735 4210 8765
rect 4240 8735 4245 8765
rect 4205 8730 4245 8735
rect 4405 8835 4445 8840
rect 4405 8805 4410 8835
rect 4440 8805 4445 8835
rect 4405 8765 4445 8805
rect 4405 8735 4410 8765
rect 4440 8735 4445 8765
rect 4405 8730 4445 8735
rect 4605 8835 4645 8840
rect 4605 8805 4610 8835
rect 4640 8805 4645 8835
rect 4605 8765 4645 8805
rect 4605 8735 4610 8765
rect 4640 8735 4645 8765
rect 4605 8730 4645 8735
rect 4805 8835 4845 8840
rect 4805 8805 4810 8835
rect 4840 8805 4845 8835
rect 4805 8765 4845 8805
rect 4805 8735 4810 8765
rect 4840 8735 4845 8765
rect 4805 8730 4845 8735
rect 5005 8835 5045 8840
rect 5005 8805 5010 8835
rect 5040 8805 5045 8835
rect 5005 8765 5045 8805
rect 5005 8735 5010 8765
rect 5040 8735 5045 8765
rect 5005 8730 5045 8735
rect 5205 8835 5245 8840
rect 5205 8805 5210 8835
rect 5240 8805 5245 8835
rect 5205 8765 5245 8805
rect 5205 8735 5210 8765
rect 5240 8735 5245 8765
rect 5205 8730 5245 8735
rect 5405 8835 5445 8840
rect 5405 8805 5410 8835
rect 5440 8805 5445 8835
rect 5405 8765 5445 8805
rect 5405 8735 5410 8765
rect 5440 8735 5445 8765
rect 5405 8730 5445 8735
rect 5605 8835 5645 8840
rect 5605 8805 5610 8835
rect 5640 8805 5645 8835
rect 5605 8765 5645 8805
rect 5605 8735 5610 8765
rect 5640 8735 5645 8765
rect 5605 8730 5645 8735
rect 5805 8835 5845 8840
rect 5805 8805 5810 8835
rect 5840 8805 5845 8835
rect 5805 8765 5845 8805
rect 5805 8735 5810 8765
rect 5840 8735 5845 8765
rect 5805 8730 5845 8735
rect 6005 8835 6045 8840
rect 6005 8805 6010 8835
rect 6040 8805 6045 8835
rect 6005 8765 6045 8805
rect 6005 8735 6010 8765
rect 6040 8735 6045 8765
rect 6005 8730 6045 8735
rect 6205 8835 6245 8840
rect 6205 8805 6210 8835
rect 6240 8805 6245 8835
rect 6205 8765 6245 8805
rect 6205 8735 6210 8765
rect 6240 8735 6245 8765
rect 6205 8730 6245 8735
rect 6405 8835 6445 8840
rect 6405 8805 6410 8835
rect 6440 8805 6445 8835
rect 6405 8765 6445 8805
rect 6405 8735 6410 8765
rect 6440 8735 6445 8765
rect 6405 8730 6445 8735
rect -195 8650 -155 8655
rect -195 8620 -190 8650
rect -160 8620 -155 8650
rect -195 8580 -155 8620
rect -195 8550 -190 8580
rect -160 8550 -155 8580
rect -195 8545 -155 8550
rect 5 8650 45 8655
rect 5 8620 10 8650
rect 40 8620 45 8650
rect 5 8580 45 8620
rect 5 8550 10 8580
rect 40 8550 45 8580
rect 5 8545 45 8550
rect 205 8650 245 8655
rect 205 8620 210 8650
rect 240 8620 245 8650
rect 205 8580 245 8620
rect 205 8550 210 8580
rect 240 8550 245 8580
rect 205 8545 245 8550
rect 405 8650 445 8655
rect 405 8620 410 8650
rect 440 8620 445 8650
rect 405 8580 445 8620
rect 405 8550 410 8580
rect 440 8550 445 8580
rect 405 8545 445 8550
rect 605 8650 645 8655
rect 605 8620 610 8650
rect 640 8620 645 8650
rect 605 8580 645 8620
rect 605 8550 610 8580
rect 640 8550 645 8580
rect 605 8545 645 8550
rect 805 8650 845 8655
rect 805 8620 810 8650
rect 840 8620 845 8650
rect 805 8580 845 8620
rect 805 8550 810 8580
rect 840 8550 845 8580
rect 805 8545 845 8550
rect 1005 8650 1045 8655
rect 1005 8620 1010 8650
rect 1040 8620 1045 8650
rect 1005 8580 1045 8620
rect 1005 8550 1010 8580
rect 1040 8550 1045 8580
rect 1005 8545 1045 8550
rect 1205 8650 1245 8655
rect 1205 8620 1210 8650
rect 1240 8620 1245 8650
rect 1205 8580 1245 8620
rect 1205 8550 1210 8580
rect 1240 8550 1245 8580
rect 1205 8545 1245 8550
rect 1405 8650 1445 8655
rect 1405 8620 1410 8650
rect 1440 8620 1445 8650
rect 1405 8580 1445 8620
rect 1405 8550 1410 8580
rect 1440 8550 1445 8580
rect 1405 8545 1445 8550
rect 1605 8650 1645 8655
rect 1605 8620 1610 8650
rect 1640 8620 1645 8650
rect 1605 8580 1645 8620
rect 1605 8550 1610 8580
rect 1640 8550 1645 8580
rect 1605 8545 1645 8550
rect 1805 8650 1845 8655
rect 1805 8620 1810 8650
rect 1840 8620 1845 8650
rect 1805 8580 1845 8620
rect 1805 8550 1810 8580
rect 1840 8550 1845 8580
rect 1805 8545 1845 8550
rect 2005 8650 2045 8655
rect 2005 8620 2010 8650
rect 2040 8620 2045 8650
rect 2005 8580 2045 8620
rect 2005 8550 2010 8580
rect 2040 8550 2045 8580
rect 2005 8545 2045 8550
rect 2205 8650 2245 8655
rect 2205 8620 2210 8650
rect 2240 8620 2245 8650
rect 2205 8580 2245 8620
rect 2205 8550 2210 8580
rect 2240 8550 2245 8580
rect 2205 8545 2245 8550
rect 2405 8650 2445 8655
rect 2405 8620 2410 8650
rect 2440 8620 2445 8650
rect 2405 8580 2445 8620
rect 2405 8550 2410 8580
rect 2440 8550 2445 8580
rect 2405 8545 2445 8550
rect 2605 8650 2645 8655
rect 2605 8620 2610 8650
rect 2640 8620 2645 8650
rect 2605 8580 2645 8620
rect 2605 8550 2610 8580
rect 2640 8550 2645 8580
rect 2605 8545 2645 8550
rect 2805 8650 2845 8655
rect 2805 8620 2810 8650
rect 2840 8620 2845 8650
rect 2805 8580 2845 8620
rect 2805 8550 2810 8580
rect 2840 8550 2845 8580
rect 2805 8545 2845 8550
rect 3005 8650 3045 8655
rect 3005 8620 3010 8650
rect 3040 8620 3045 8650
rect 3005 8580 3045 8620
rect 3005 8550 3010 8580
rect 3040 8550 3045 8580
rect 3005 8545 3045 8550
rect 3205 8650 3245 8655
rect 3205 8620 3210 8650
rect 3240 8620 3245 8650
rect 3205 8580 3245 8620
rect 3205 8550 3210 8580
rect 3240 8550 3245 8580
rect 3205 8545 3245 8550
rect 3405 8650 3445 8655
rect 3405 8620 3410 8650
rect 3440 8620 3445 8650
rect 3405 8580 3445 8620
rect 3405 8550 3410 8580
rect 3440 8550 3445 8580
rect 3405 8545 3445 8550
rect 3605 8650 3645 8655
rect 3605 8620 3610 8650
rect 3640 8620 3645 8650
rect 3605 8580 3645 8620
rect 3605 8550 3610 8580
rect 3640 8550 3645 8580
rect 3605 8545 3645 8550
rect 3805 8650 3845 8655
rect 3805 8620 3810 8650
rect 3840 8620 3845 8650
rect 3805 8580 3845 8620
rect 3805 8550 3810 8580
rect 3840 8550 3845 8580
rect 3805 8545 3845 8550
rect 4005 8650 4045 8655
rect 4005 8620 4010 8650
rect 4040 8620 4045 8650
rect 4005 8580 4045 8620
rect 4005 8550 4010 8580
rect 4040 8550 4045 8580
rect 4005 8545 4045 8550
rect 4205 8650 4245 8655
rect 4205 8620 4210 8650
rect 4240 8620 4245 8650
rect 4205 8580 4245 8620
rect 4205 8550 4210 8580
rect 4240 8550 4245 8580
rect 4205 8545 4245 8550
rect 4405 8650 4445 8655
rect 4405 8620 4410 8650
rect 4440 8620 4445 8650
rect 4405 8580 4445 8620
rect 4405 8550 4410 8580
rect 4440 8550 4445 8580
rect 4405 8545 4445 8550
rect 4605 8650 4645 8655
rect 4605 8620 4610 8650
rect 4640 8620 4645 8650
rect 4605 8580 4645 8620
rect 4605 8550 4610 8580
rect 4640 8550 4645 8580
rect 4605 8545 4645 8550
rect 4805 8650 4845 8655
rect 4805 8620 4810 8650
rect 4840 8620 4845 8650
rect 4805 8580 4845 8620
rect 4805 8550 4810 8580
rect 4840 8550 4845 8580
rect 4805 8545 4845 8550
rect 5005 8650 5045 8655
rect 5005 8620 5010 8650
rect 5040 8620 5045 8650
rect 5005 8580 5045 8620
rect 5005 8550 5010 8580
rect 5040 8550 5045 8580
rect 5005 8545 5045 8550
rect 5205 8650 5245 8655
rect 5205 8620 5210 8650
rect 5240 8620 5245 8650
rect 5205 8580 5245 8620
rect 5205 8550 5210 8580
rect 5240 8550 5245 8580
rect 5205 8545 5245 8550
rect 5405 8650 5445 8655
rect 5405 8620 5410 8650
rect 5440 8620 5445 8650
rect 5405 8580 5445 8620
rect 5405 8550 5410 8580
rect 5440 8550 5445 8580
rect 5405 8545 5445 8550
rect 5605 8650 5645 8655
rect 5605 8620 5610 8650
rect 5640 8620 5645 8650
rect 5605 8580 5645 8620
rect 5605 8550 5610 8580
rect 5640 8550 5645 8580
rect 5605 8545 5645 8550
rect 5805 8650 5845 8655
rect 5805 8620 5810 8650
rect 5840 8620 5845 8650
rect 5805 8580 5845 8620
rect 5805 8550 5810 8580
rect 5840 8550 5845 8580
rect 5805 8545 5845 8550
rect 6005 8650 6045 8655
rect 6005 8620 6010 8650
rect 6040 8620 6045 8650
rect 6005 8580 6045 8620
rect 6005 8550 6010 8580
rect 6040 8550 6045 8580
rect 6005 8545 6045 8550
rect 6205 8650 6245 8655
rect 6205 8620 6210 8650
rect 6240 8620 6245 8650
rect 6205 8580 6245 8620
rect 6205 8550 6210 8580
rect 6240 8550 6245 8580
rect 6205 8545 6245 8550
rect 6405 8650 6445 8655
rect 6405 8620 6410 8650
rect 6440 8620 6445 8650
rect 6405 8580 6445 8620
rect 6405 8550 6410 8580
rect 6440 8550 6445 8580
rect 6405 8545 6445 8550
rect -195 8465 -155 8470
rect -195 8435 -190 8465
rect -160 8435 -155 8465
rect -195 8395 -155 8435
rect -195 8365 -190 8395
rect -160 8365 -155 8395
rect -195 8360 -155 8365
rect 5 8465 45 8470
rect 5 8435 10 8465
rect 40 8435 45 8465
rect 5 8395 45 8435
rect 5 8365 10 8395
rect 40 8365 45 8395
rect 5 8360 45 8365
rect 205 8465 245 8470
rect 205 8435 210 8465
rect 240 8435 245 8465
rect 205 8395 245 8435
rect 205 8365 210 8395
rect 240 8365 245 8395
rect 205 8360 245 8365
rect 405 8465 445 8470
rect 405 8435 410 8465
rect 440 8435 445 8465
rect 405 8395 445 8435
rect 405 8365 410 8395
rect 440 8365 445 8395
rect 405 8360 445 8365
rect 605 8465 645 8470
rect 605 8435 610 8465
rect 640 8435 645 8465
rect 605 8395 645 8435
rect 605 8365 610 8395
rect 640 8365 645 8395
rect 605 8360 645 8365
rect 805 8465 845 8470
rect 805 8435 810 8465
rect 840 8435 845 8465
rect 805 8395 845 8435
rect 805 8365 810 8395
rect 840 8365 845 8395
rect 805 8360 845 8365
rect 1005 8465 1045 8470
rect 1005 8435 1010 8465
rect 1040 8435 1045 8465
rect 1005 8395 1045 8435
rect 1005 8365 1010 8395
rect 1040 8365 1045 8395
rect 1005 8360 1045 8365
rect 1205 8465 1245 8470
rect 1205 8435 1210 8465
rect 1240 8435 1245 8465
rect 1205 8395 1245 8435
rect 1205 8365 1210 8395
rect 1240 8365 1245 8395
rect 1205 8360 1245 8365
rect 1405 8465 1445 8470
rect 1405 8435 1410 8465
rect 1440 8435 1445 8465
rect 1405 8395 1445 8435
rect 1405 8365 1410 8395
rect 1440 8365 1445 8395
rect 1405 8360 1445 8365
rect 1605 8465 1645 8470
rect 1605 8435 1610 8465
rect 1640 8435 1645 8465
rect 1605 8395 1645 8435
rect 1605 8365 1610 8395
rect 1640 8365 1645 8395
rect 1605 8360 1645 8365
rect 1805 8465 1845 8470
rect 1805 8435 1810 8465
rect 1840 8435 1845 8465
rect 1805 8395 1845 8435
rect 1805 8365 1810 8395
rect 1840 8365 1845 8395
rect 1805 8360 1845 8365
rect 2005 8465 2045 8470
rect 2005 8435 2010 8465
rect 2040 8435 2045 8465
rect 2005 8395 2045 8435
rect 2005 8365 2010 8395
rect 2040 8365 2045 8395
rect 2005 8360 2045 8365
rect 2205 8465 2245 8470
rect 2205 8435 2210 8465
rect 2240 8435 2245 8465
rect 2205 8395 2245 8435
rect 2205 8365 2210 8395
rect 2240 8365 2245 8395
rect 2205 8360 2245 8365
rect 2405 8465 2445 8470
rect 2405 8435 2410 8465
rect 2440 8435 2445 8465
rect 2405 8395 2445 8435
rect 2405 8365 2410 8395
rect 2440 8365 2445 8395
rect 2405 8360 2445 8365
rect 2605 8465 2645 8470
rect 2605 8435 2610 8465
rect 2640 8435 2645 8465
rect 2605 8395 2645 8435
rect 2605 8365 2610 8395
rect 2640 8365 2645 8395
rect 2605 8360 2645 8365
rect 2805 8465 2845 8470
rect 2805 8435 2810 8465
rect 2840 8435 2845 8465
rect 2805 8395 2845 8435
rect 2805 8365 2810 8395
rect 2840 8365 2845 8395
rect 2805 8360 2845 8365
rect 3005 8465 3045 8470
rect 3005 8435 3010 8465
rect 3040 8435 3045 8465
rect 3005 8395 3045 8435
rect 3005 8365 3010 8395
rect 3040 8365 3045 8395
rect 3005 8360 3045 8365
rect 3205 8465 3245 8470
rect 3205 8435 3210 8465
rect 3240 8435 3245 8465
rect 3205 8395 3245 8435
rect 3205 8365 3210 8395
rect 3240 8365 3245 8395
rect 3205 8360 3245 8365
rect 3405 8465 3445 8470
rect 3405 8435 3410 8465
rect 3440 8435 3445 8465
rect 3405 8395 3445 8435
rect 3405 8365 3410 8395
rect 3440 8365 3445 8395
rect 3405 8360 3445 8365
rect 3605 8465 3645 8470
rect 3605 8435 3610 8465
rect 3640 8435 3645 8465
rect 3605 8395 3645 8435
rect 3605 8365 3610 8395
rect 3640 8365 3645 8395
rect 3605 8360 3645 8365
rect 3805 8465 3845 8470
rect 3805 8435 3810 8465
rect 3840 8435 3845 8465
rect 3805 8395 3845 8435
rect 3805 8365 3810 8395
rect 3840 8365 3845 8395
rect 3805 8360 3845 8365
rect 4005 8465 4045 8470
rect 4005 8435 4010 8465
rect 4040 8435 4045 8465
rect 4005 8395 4045 8435
rect 4005 8365 4010 8395
rect 4040 8365 4045 8395
rect 4005 8360 4045 8365
rect 4205 8465 4245 8470
rect 4205 8435 4210 8465
rect 4240 8435 4245 8465
rect 4205 8395 4245 8435
rect 4205 8365 4210 8395
rect 4240 8365 4245 8395
rect 4205 8360 4245 8365
rect 4405 8465 4445 8470
rect 4405 8435 4410 8465
rect 4440 8435 4445 8465
rect 4405 8395 4445 8435
rect 4405 8365 4410 8395
rect 4440 8365 4445 8395
rect 4405 8360 4445 8365
rect 4605 8465 4645 8470
rect 4605 8435 4610 8465
rect 4640 8435 4645 8465
rect 4605 8395 4645 8435
rect 4605 8365 4610 8395
rect 4640 8365 4645 8395
rect 4605 8360 4645 8365
rect 4805 8465 4845 8470
rect 4805 8435 4810 8465
rect 4840 8435 4845 8465
rect 4805 8395 4845 8435
rect 4805 8365 4810 8395
rect 4840 8365 4845 8395
rect 4805 8360 4845 8365
rect 5005 8465 5045 8470
rect 5005 8435 5010 8465
rect 5040 8435 5045 8465
rect 5005 8395 5045 8435
rect 5005 8365 5010 8395
rect 5040 8365 5045 8395
rect 5005 8360 5045 8365
rect 5205 8465 5245 8470
rect 5205 8435 5210 8465
rect 5240 8435 5245 8465
rect 5205 8395 5245 8435
rect 5205 8365 5210 8395
rect 5240 8365 5245 8395
rect 5205 8360 5245 8365
rect 5405 8465 5445 8470
rect 5405 8435 5410 8465
rect 5440 8435 5445 8465
rect 5405 8395 5445 8435
rect 5405 8365 5410 8395
rect 5440 8365 5445 8395
rect 5405 8360 5445 8365
rect 5605 8465 5645 8470
rect 5605 8435 5610 8465
rect 5640 8435 5645 8465
rect 5605 8395 5645 8435
rect 5605 8365 5610 8395
rect 5640 8365 5645 8395
rect 5605 8360 5645 8365
rect 5805 8465 5845 8470
rect 5805 8435 5810 8465
rect 5840 8435 5845 8465
rect 5805 8395 5845 8435
rect 5805 8365 5810 8395
rect 5840 8365 5845 8395
rect 5805 8360 5845 8365
rect 6005 8465 6045 8470
rect 6005 8435 6010 8465
rect 6040 8435 6045 8465
rect 6005 8395 6045 8435
rect 6005 8365 6010 8395
rect 6040 8365 6045 8395
rect 6005 8360 6045 8365
rect 6205 8465 6245 8470
rect 6205 8435 6210 8465
rect 6240 8435 6245 8465
rect 6205 8395 6245 8435
rect 6205 8365 6210 8395
rect 6240 8365 6245 8395
rect 6205 8360 6245 8365
rect 6405 8465 6445 8470
rect 6405 8435 6410 8465
rect 6440 8435 6445 8465
rect 6405 8395 6445 8435
rect 6405 8365 6410 8395
rect 6440 8365 6445 8395
rect 6405 8360 6445 8365
rect -195 8280 -155 8285
rect -195 8250 -190 8280
rect -160 8250 -155 8280
rect -195 8210 -155 8250
rect -195 8180 -190 8210
rect -160 8180 -155 8210
rect -195 8175 -155 8180
rect 5 8280 45 8285
rect 5 8250 10 8280
rect 40 8250 45 8280
rect 5 8210 45 8250
rect 5 8180 10 8210
rect 40 8180 45 8210
rect 5 8175 45 8180
rect 205 8280 245 8285
rect 205 8250 210 8280
rect 240 8250 245 8280
rect 205 8210 245 8250
rect 205 8180 210 8210
rect 240 8180 245 8210
rect 205 8175 245 8180
rect 405 8280 445 8285
rect 405 8250 410 8280
rect 440 8250 445 8280
rect 405 8210 445 8250
rect 405 8180 410 8210
rect 440 8180 445 8210
rect 405 8175 445 8180
rect 605 8280 645 8285
rect 605 8250 610 8280
rect 640 8250 645 8280
rect 605 8210 645 8250
rect 605 8180 610 8210
rect 640 8180 645 8210
rect 605 8175 645 8180
rect 805 8280 845 8285
rect 805 8250 810 8280
rect 840 8250 845 8280
rect 805 8210 845 8250
rect 805 8180 810 8210
rect 840 8180 845 8210
rect 805 8175 845 8180
rect 1005 8280 1045 8285
rect 1005 8250 1010 8280
rect 1040 8250 1045 8280
rect 1005 8210 1045 8250
rect 1005 8180 1010 8210
rect 1040 8180 1045 8210
rect 1005 8175 1045 8180
rect 1205 8280 1245 8285
rect 1205 8250 1210 8280
rect 1240 8250 1245 8280
rect 1205 8210 1245 8250
rect 1205 8180 1210 8210
rect 1240 8180 1245 8210
rect 1205 8175 1245 8180
rect 1405 8280 1445 8285
rect 1405 8250 1410 8280
rect 1440 8250 1445 8280
rect 1405 8210 1445 8250
rect 1405 8180 1410 8210
rect 1440 8180 1445 8210
rect 1405 8175 1445 8180
rect 1605 8280 1645 8285
rect 1605 8250 1610 8280
rect 1640 8250 1645 8280
rect 1605 8210 1645 8250
rect 1605 8180 1610 8210
rect 1640 8180 1645 8210
rect 1605 8175 1645 8180
rect 1805 8280 1845 8285
rect 1805 8250 1810 8280
rect 1840 8250 1845 8280
rect 1805 8210 1845 8250
rect 1805 8180 1810 8210
rect 1840 8180 1845 8210
rect 1805 8175 1845 8180
rect 2005 8280 2045 8285
rect 2005 8250 2010 8280
rect 2040 8250 2045 8280
rect 2005 8210 2045 8250
rect 2005 8180 2010 8210
rect 2040 8180 2045 8210
rect 2005 8175 2045 8180
rect 2205 8280 2245 8285
rect 2205 8250 2210 8280
rect 2240 8250 2245 8280
rect 2205 8210 2245 8250
rect 2205 8180 2210 8210
rect 2240 8180 2245 8210
rect 2205 8175 2245 8180
rect 2405 8280 2445 8285
rect 2405 8250 2410 8280
rect 2440 8250 2445 8280
rect 2405 8210 2445 8250
rect 2405 8180 2410 8210
rect 2440 8180 2445 8210
rect 2405 8175 2445 8180
rect 2605 8280 2645 8285
rect 2605 8250 2610 8280
rect 2640 8250 2645 8280
rect 2605 8210 2645 8250
rect 2605 8180 2610 8210
rect 2640 8180 2645 8210
rect 2605 8175 2645 8180
rect 2805 8280 2845 8285
rect 2805 8250 2810 8280
rect 2840 8250 2845 8280
rect 2805 8210 2845 8250
rect 2805 8180 2810 8210
rect 2840 8180 2845 8210
rect 2805 8175 2845 8180
rect 3005 8280 3045 8285
rect 3005 8250 3010 8280
rect 3040 8250 3045 8280
rect 3005 8210 3045 8250
rect 3005 8180 3010 8210
rect 3040 8180 3045 8210
rect 3005 8175 3045 8180
rect 3205 8280 3245 8285
rect 3205 8250 3210 8280
rect 3240 8250 3245 8280
rect 3205 8210 3245 8250
rect 3205 8180 3210 8210
rect 3240 8180 3245 8210
rect 3205 8175 3245 8180
rect 3405 8280 3445 8285
rect 3405 8250 3410 8280
rect 3440 8250 3445 8280
rect 3405 8210 3445 8250
rect 3405 8180 3410 8210
rect 3440 8180 3445 8210
rect 3405 8175 3445 8180
rect 3605 8280 3645 8285
rect 3605 8250 3610 8280
rect 3640 8250 3645 8280
rect 3605 8210 3645 8250
rect 3605 8180 3610 8210
rect 3640 8180 3645 8210
rect 3605 8175 3645 8180
rect 3805 8280 3845 8285
rect 3805 8250 3810 8280
rect 3840 8250 3845 8280
rect 3805 8210 3845 8250
rect 3805 8180 3810 8210
rect 3840 8180 3845 8210
rect 3805 8175 3845 8180
rect 4005 8280 4045 8285
rect 4005 8250 4010 8280
rect 4040 8250 4045 8280
rect 4005 8210 4045 8250
rect 4005 8180 4010 8210
rect 4040 8180 4045 8210
rect 4005 8175 4045 8180
rect 4205 8280 4245 8285
rect 4205 8250 4210 8280
rect 4240 8250 4245 8280
rect 4205 8210 4245 8250
rect 4205 8180 4210 8210
rect 4240 8180 4245 8210
rect 4205 8175 4245 8180
rect 4405 8280 4445 8285
rect 4405 8250 4410 8280
rect 4440 8250 4445 8280
rect 4405 8210 4445 8250
rect 4405 8180 4410 8210
rect 4440 8180 4445 8210
rect 4405 8175 4445 8180
rect 4605 8280 4645 8285
rect 4605 8250 4610 8280
rect 4640 8250 4645 8280
rect 4605 8210 4645 8250
rect 4605 8180 4610 8210
rect 4640 8180 4645 8210
rect 4605 8175 4645 8180
rect 4805 8280 4845 8285
rect 4805 8250 4810 8280
rect 4840 8250 4845 8280
rect 4805 8210 4845 8250
rect 4805 8180 4810 8210
rect 4840 8180 4845 8210
rect 4805 8175 4845 8180
rect 5005 8280 5045 8285
rect 5005 8250 5010 8280
rect 5040 8250 5045 8280
rect 5005 8210 5045 8250
rect 5005 8180 5010 8210
rect 5040 8180 5045 8210
rect 5005 8175 5045 8180
rect 5205 8280 5245 8285
rect 5205 8250 5210 8280
rect 5240 8250 5245 8280
rect 5205 8210 5245 8250
rect 5205 8180 5210 8210
rect 5240 8180 5245 8210
rect 5205 8175 5245 8180
rect 5405 8280 5445 8285
rect 5405 8250 5410 8280
rect 5440 8250 5445 8280
rect 5405 8210 5445 8250
rect 5405 8180 5410 8210
rect 5440 8180 5445 8210
rect 5405 8175 5445 8180
rect 5605 8280 5645 8285
rect 5605 8250 5610 8280
rect 5640 8250 5645 8280
rect 5605 8210 5645 8250
rect 5605 8180 5610 8210
rect 5640 8180 5645 8210
rect 5605 8175 5645 8180
rect 5805 8280 5845 8285
rect 5805 8250 5810 8280
rect 5840 8250 5845 8280
rect 5805 8210 5845 8250
rect 5805 8180 5810 8210
rect 5840 8180 5845 8210
rect 5805 8175 5845 8180
rect 6005 8280 6045 8285
rect 6005 8250 6010 8280
rect 6040 8250 6045 8280
rect 6005 8210 6045 8250
rect 6005 8180 6010 8210
rect 6040 8180 6045 8210
rect 6005 8175 6045 8180
rect 6205 8280 6245 8285
rect 6205 8250 6210 8280
rect 6240 8250 6245 8280
rect 6205 8210 6245 8250
rect 6205 8180 6210 8210
rect 6240 8180 6245 8210
rect 6205 8175 6245 8180
rect 6405 8280 6445 8285
rect 6405 8250 6410 8280
rect 6440 8250 6445 8280
rect 6405 8210 6445 8250
rect 6405 8180 6410 8210
rect 6440 8180 6445 8210
rect 6405 8175 6445 8180
rect -195 8095 -155 8100
rect -195 8065 -190 8095
rect -160 8065 -155 8095
rect -195 8025 -155 8065
rect -195 7995 -190 8025
rect -160 7995 -155 8025
rect -195 7990 -155 7995
rect 5 8095 45 8100
rect 5 8065 10 8095
rect 40 8065 45 8095
rect 5 8025 45 8065
rect 5 7995 10 8025
rect 40 7995 45 8025
rect 5 7990 45 7995
rect 205 8095 245 8100
rect 205 8065 210 8095
rect 240 8065 245 8095
rect 205 8025 245 8065
rect 205 7995 210 8025
rect 240 7995 245 8025
rect 205 7990 245 7995
rect 405 8095 445 8100
rect 405 8065 410 8095
rect 440 8065 445 8095
rect 405 8025 445 8065
rect 405 7995 410 8025
rect 440 7995 445 8025
rect 405 7990 445 7995
rect 605 8095 645 8100
rect 605 8065 610 8095
rect 640 8065 645 8095
rect 605 8025 645 8065
rect 605 7995 610 8025
rect 640 7995 645 8025
rect 605 7990 645 7995
rect 805 8095 845 8100
rect 805 8065 810 8095
rect 840 8065 845 8095
rect 805 8025 845 8065
rect 805 7995 810 8025
rect 840 7995 845 8025
rect 805 7990 845 7995
rect 1005 8095 1045 8100
rect 1005 8065 1010 8095
rect 1040 8065 1045 8095
rect 1005 8025 1045 8065
rect 1005 7995 1010 8025
rect 1040 7995 1045 8025
rect 1005 7990 1045 7995
rect 1205 8095 1245 8100
rect 1205 8065 1210 8095
rect 1240 8065 1245 8095
rect 1205 8025 1245 8065
rect 1205 7995 1210 8025
rect 1240 7995 1245 8025
rect 1205 7990 1245 7995
rect 1405 8095 1445 8100
rect 1405 8065 1410 8095
rect 1440 8065 1445 8095
rect 1405 8025 1445 8065
rect 1405 7995 1410 8025
rect 1440 7995 1445 8025
rect 1405 7990 1445 7995
rect 1605 8095 1645 8100
rect 1605 8065 1610 8095
rect 1640 8065 1645 8095
rect 1605 8025 1645 8065
rect 1605 7995 1610 8025
rect 1640 7995 1645 8025
rect 1605 7990 1645 7995
rect 1805 8095 1845 8100
rect 1805 8065 1810 8095
rect 1840 8065 1845 8095
rect 1805 8025 1845 8065
rect 1805 7995 1810 8025
rect 1840 7995 1845 8025
rect 1805 7990 1845 7995
rect 2005 8095 2045 8100
rect 2005 8065 2010 8095
rect 2040 8065 2045 8095
rect 2005 8025 2045 8065
rect 2005 7995 2010 8025
rect 2040 7995 2045 8025
rect 2005 7990 2045 7995
rect 2205 8095 2245 8100
rect 2205 8065 2210 8095
rect 2240 8065 2245 8095
rect 2205 8025 2245 8065
rect 2205 7995 2210 8025
rect 2240 7995 2245 8025
rect 2205 7990 2245 7995
rect 2405 8095 2445 8100
rect 2405 8065 2410 8095
rect 2440 8065 2445 8095
rect 2405 8025 2445 8065
rect 2405 7995 2410 8025
rect 2440 7995 2445 8025
rect 2405 7990 2445 7995
rect 2605 8095 2645 8100
rect 2605 8065 2610 8095
rect 2640 8065 2645 8095
rect 2605 8025 2645 8065
rect 2605 7995 2610 8025
rect 2640 7995 2645 8025
rect 2605 7990 2645 7995
rect 2805 8095 2845 8100
rect 2805 8065 2810 8095
rect 2840 8065 2845 8095
rect 2805 8025 2845 8065
rect 2805 7995 2810 8025
rect 2840 7995 2845 8025
rect 2805 7990 2845 7995
rect 3005 8095 3045 8100
rect 3005 8065 3010 8095
rect 3040 8065 3045 8095
rect 3005 8025 3045 8065
rect 3005 7995 3010 8025
rect 3040 7995 3045 8025
rect 3005 7990 3045 7995
rect 3205 8095 3245 8100
rect 3205 8065 3210 8095
rect 3240 8065 3245 8095
rect 3205 8025 3245 8065
rect 3205 7995 3210 8025
rect 3240 7995 3245 8025
rect 3205 7990 3245 7995
rect 3405 8095 3445 8100
rect 3405 8065 3410 8095
rect 3440 8065 3445 8095
rect 3405 8025 3445 8065
rect 3405 7995 3410 8025
rect 3440 7995 3445 8025
rect 3405 7990 3445 7995
rect 3605 8095 3645 8100
rect 3605 8065 3610 8095
rect 3640 8065 3645 8095
rect 3605 8025 3645 8065
rect 3605 7995 3610 8025
rect 3640 7995 3645 8025
rect 3605 7990 3645 7995
rect 3805 8095 3845 8100
rect 3805 8065 3810 8095
rect 3840 8065 3845 8095
rect 3805 8025 3845 8065
rect 3805 7995 3810 8025
rect 3840 7995 3845 8025
rect 3805 7990 3845 7995
rect 4005 8095 4045 8100
rect 4005 8065 4010 8095
rect 4040 8065 4045 8095
rect 4005 8025 4045 8065
rect 4005 7995 4010 8025
rect 4040 7995 4045 8025
rect 4005 7990 4045 7995
rect 4205 8095 4245 8100
rect 4205 8065 4210 8095
rect 4240 8065 4245 8095
rect 4205 8025 4245 8065
rect 4205 7995 4210 8025
rect 4240 7995 4245 8025
rect 4205 7990 4245 7995
rect 4405 8095 4445 8100
rect 4405 8065 4410 8095
rect 4440 8065 4445 8095
rect 4405 8025 4445 8065
rect 4405 7995 4410 8025
rect 4440 7995 4445 8025
rect 4405 7990 4445 7995
rect 4605 8095 4645 8100
rect 4605 8065 4610 8095
rect 4640 8065 4645 8095
rect 4605 8025 4645 8065
rect 4605 7995 4610 8025
rect 4640 7995 4645 8025
rect 4605 7990 4645 7995
rect 4805 8095 4845 8100
rect 4805 8065 4810 8095
rect 4840 8065 4845 8095
rect 4805 8025 4845 8065
rect 4805 7995 4810 8025
rect 4840 7995 4845 8025
rect 4805 7990 4845 7995
rect 5005 8095 5045 8100
rect 5005 8065 5010 8095
rect 5040 8065 5045 8095
rect 5005 8025 5045 8065
rect 5005 7995 5010 8025
rect 5040 7995 5045 8025
rect 5005 7990 5045 7995
rect 5205 8095 5245 8100
rect 5205 8065 5210 8095
rect 5240 8065 5245 8095
rect 5205 8025 5245 8065
rect 5205 7995 5210 8025
rect 5240 7995 5245 8025
rect 5205 7990 5245 7995
rect 5405 8095 5445 8100
rect 5405 8065 5410 8095
rect 5440 8065 5445 8095
rect 5405 8025 5445 8065
rect 5405 7995 5410 8025
rect 5440 7995 5445 8025
rect 5405 7990 5445 7995
rect 5605 8095 5645 8100
rect 5605 8065 5610 8095
rect 5640 8065 5645 8095
rect 5605 8025 5645 8065
rect 5605 7995 5610 8025
rect 5640 7995 5645 8025
rect 5605 7990 5645 7995
rect 5805 8095 5845 8100
rect 5805 8065 5810 8095
rect 5840 8065 5845 8095
rect 5805 8025 5845 8065
rect 5805 7995 5810 8025
rect 5840 7995 5845 8025
rect 5805 7990 5845 7995
rect 6005 8095 6045 8100
rect 6005 8065 6010 8095
rect 6040 8065 6045 8095
rect 6005 8025 6045 8065
rect 6005 7995 6010 8025
rect 6040 7995 6045 8025
rect 6005 7990 6045 7995
rect 6205 8095 6245 8100
rect 6205 8065 6210 8095
rect 6240 8065 6245 8095
rect 6205 8025 6245 8065
rect 6205 7995 6210 8025
rect 6240 7995 6245 8025
rect 6205 7990 6245 7995
rect 6405 8095 6445 8100
rect 6405 8065 6410 8095
rect 6440 8065 6445 8095
rect 6405 8025 6445 8065
rect 6405 7995 6410 8025
rect 6440 7995 6445 8025
rect 6405 7990 6445 7995
rect -195 7910 -155 7915
rect -195 7880 -190 7910
rect -160 7880 -155 7910
rect -195 7840 -155 7880
rect -195 7810 -190 7840
rect -160 7810 -155 7840
rect -195 7805 -155 7810
rect 5 7910 45 7915
rect 5 7880 10 7910
rect 40 7880 45 7910
rect 5 7840 45 7880
rect 5 7810 10 7840
rect 40 7810 45 7840
rect 5 7805 45 7810
rect 205 7910 245 7915
rect 205 7880 210 7910
rect 240 7880 245 7910
rect 205 7840 245 7880
rect 205 7810 210 7840
rect 240 7810 245 7840
rect 205 7805 245 7810
rect 405 7910 445 7915
rect 405 7880 410 7910
rect 440 7880 445 7910
rect 405 7840 445 7880
rect 405 7810 410 7840
rect 440 7810 445 7840
rect 405 7805 445 7810
rect 605 7910 645 7915
rect 605 7880 610 7910
rect 640 7880 645 7910
rect 605 7840 645 7880
rect 605 7810 610 7840
rect 640 7810 645 7840
rect 605 7805 645 7810
rect 805 7910 845 7915
rect 805 7880 810 7910
rect 840 7880 845 7910
rect 805 7840 845 7880
rect 805 7810 810 7840
rect 840 7810 845 7840
rect 805 7805 845 7810
rect 1005 7910 1045 7915
rect 1005 7880 1010 7910
rect 1040 7880 1045 7910
rect 1005 7840 1045 7880
rect 1005 7810 1010 7840
rect 1040 7810 1045 7840
rect 1005 7805 1045 7810
rect 1205 7910 1245 7915
rect 1205 7880 1210 7910
rect 1240 7880 1245 7910
rect 1205 7840 1245 7880
rect 1205 7810 1210 7840
rect 1240 7810 1245 7840
rect 1205 7805 1245 7810
rect 1405 7910 1445 7915
rect 1405 7880 1410 7910
rect 1440 7880 1445 7910
rect 1405 7840 1445 7880
rect 1405 7810 1410 7840
rect 1440 7810 1445 7840
rect 1405 7805 1445 7810
rect 1605 7910 1645 7915
rect 1605 7880 1610 7910
rect 1640 7880 1645 7910
rect 1605 7840 1645 7880
rect 1605 7810 1610 7840
rect 1640 7810 1645 7840
rect 1605 7805 1645 7810
rect 1805 7910 1845 7915
rect 1805 7880 1810 7910
rect 1840 7880 1845 7910
rect 1805 7840 1845 7880
rect 1805 7810 1810 7840
rect 1840 7810 1845 7840
rect 1805 7805 1845 7810
rect 2005 7910 2045 7915
rect 2005 7880 2010 7910
rect 2040 7880 2045 7910
rect 2005 7840 2045 7880
rect 2005 7810 2010 7840
rect 2040 7810 2045 7840
rect 2005 7805 2045 7810
rect 2205 7910 2245 7915
rect 2205 7880 2210 7910
rect 2240 7880 2245 7910
rect 2205 7840 2245 7880
rect 2205 7810 2210 7840
rect 2240 7810 2245 7840
rect 2205 7805 2245 7810
rect 2405 7910 2445 7915
rect 2405 7880 2410 7910
rect 2440 7880 2445 7910
rect 2405 7840 2445 7880
rect 2405 7810 2410 7840
rect 2440 7810 2445 7840
rect 2405 7805 2445 7810
rect 2605 7910 2645 7915
rect 2605 7880 2610 7910
rect 2640 7880 2645 7910
rect 2605 7840 2645 7880
rect 2605 7810 2610 7840
rect 2640 7810 2645 7840
rect 2605 7805 2645 7810
rect 2805 7910 2845 7915
rect 2805 7880 2810 7910
rect 2840 7880 2845 7910
rect 2805 7840 2845 7880
rect 2805 7810 2810 7840
rect 2840 7810 2845 7840
rect 2805 7805 2845 7810
rect 3005 7910 3045 7915
rect 3005 7880 3010 7910
rect 3040 7880 3045 7910
rect 3005 7840 3045 7880
rect 3005 7810 3010 7840
rect 3040 7810 3045 7840
rect 3005 7805 3045 7810
rect 3205 7910 3245 7915
rect 3205 7880 3210 7910
rect 3240 7880 3245 7910
rect 3205 7840 3245 7880
rect 3205 7810 3210 7840
rect 3240 7810 3245 7840
rect 3205 7805 3245 7810
rect 3405 7910 3445 7915
rect 3405 7880 3410 7910
rect 3440 7880 3445 7910
rect 3405 7840 3445 7880
rect 3405 7810 3410 7840
rect 3440 7810 3445 7840
rect 3405 7805 3445 7810
rect 3605 7910 3645 7915
rect 3605 7880 3610 7910
rect 3640 7880 3645 7910
rect 3605 7840 3645 7880
rect 3605 7810 3610 7840
rect 3640 7810 3645 7840
rect 3605 7805 3645 7810
rect 3805 7910 3845 7915
rect 3805 7880 3810 7910
rect 3840 7880 3845 7910
rect 3805 7840 3845 7880
rect 3805 7810 3810 7840
rect 3840 7810 3845 7840
rect 3805 7805 3845 7810
rect 4005 7910 4045 7915
rect 4005 7880 4010 7910
rect 4040 7880 4045 7910
rect 4005 7840 4045 7880
rect 4005 7810 4010 7840
rect 4040 7810 4045 7840
rect 4005 7805 4045 7810
rect 4205 7910 4245 7915
rect 4205 7880 4210 7910
rect 4240 7880 4245 7910
rect 4205 7840 4245 7880
rect 4205 7810 4210 7840
rect 4240 7810 4245 7840
rect 4205 7805 4245 7810
rect 4405 7910 4445 7915
rect 4405 7880 4410 7910
rect 4440 7880 4445 7910
rect 4405 7840 4445 7880
rect 4405 7810 4410 7840
rect 4440 7810 4445 7840
rect 4405 7805 4445 7810
rect 4605 7910 4645 7915
rect 4605 7880 4610 7910
rect 4640 7880 4645 7910
rect 4605 7840 4645 7880
rect 4605 7810 4610 7840
rect 4640 7810 4645 7840
rect 4605 7805 4645 7810
rect 4805 7910 4845 7915
rect 4805 7880 4810 7910
rect 4840 7880 4845 7910
rect 4805 7840 4845 7880
rect 4805 7810 4810 7840
rect 4840 7810 4845 7840
rect 4805 7805 4845 7810
rect 5005 7910 5045 7915
rect 5005 7880 5010 7910
rect 5040 7880 5045 7910
rect 5005 7840 5045 7880
rect 5005 7810 5010 7840
rect 5040 7810 5045 7840
rect 5005 7805 5045 7810
rect 5205 7910 5245 7915
rect 5205 7880 5210 7910
rect 5240 7880 5245 7910
rect 5205 7840 5245 7880
rect 5205 7810 5210 7840
rect 5240 7810 5245 7840
rect 5205 7805 5245 7810
rect 5405 7910 5445 7915
rect 5405 7880 5410 7910
rect 5440 7880 5445 7910
rect 5405 7840 5445 7880
rect 5405 7810 5410 7840
rect 5440 7810 5445 7840
rect 5405 7805 5445 7810
rect 5605 7910 5645 7915
rect 5605 7880 5610 7910
rect 5640 7880 5645 7910
rect 5605 7840 5645 7880
rect 5605 7810 5610 7840
rect 5640 7810 5645 7840
rect 5605 7805 5645 7810
rect 5805 7910 5845 7915
rect 5805 7880 5810 7910
rect 5840 7880 5845 7910
rect 5805 7840 5845 7880
rect 5805 7810 5810 7840
rect 5840 7810 5845 7840
rect 5805 7805 5845 7810
rect 6005 7910 6045 7915
rect 6005 7880 6010 7910
rect 6040 7880 6045 7910
rect 6005 7840 6045 7880
rect 6005 7810 6010 7840
rect 6040 7810 6045 7840
rect 6005 7805 6045 7810
rect 6205 7910 6245 7915
rect 6205 7880 6210 7910
rect 6240 7880 6245 7910
rect 6205 7840 6245 7880
rect 6205 7810 6210 7840
rect 6240 7810 6245 7840
rect 6205 7805 6245 7810
rect 6405 7910 6445 7915
rect 6405 7880 6410 7910
rect 6440 7880 6445 7910
rect 6405 7840 6445 7880
rect 6405 7810 6410 7840
rect 6440 7810 6445 7840
rect 6405 7805 6445 7810
rect -195 7725 -155 7730
rect -195 7695 -190 7725
rect -160 7695 -155 7725
rect -195 7655 -155 7695
rect -195 7625 -190 7655
rect -160 7625 -155 7655
rect -195 7620 -155 7625
rect 5 7725 45 7730
rect 5 7695 10 7725
rect 40 7695 45 7725
rect 5 7655 45 7695
rect 5 7625 10 7655
rect 40 7625 45 7655
rect 5 7620 45 7625
rect 205 7725 245 7730
rect 205 7695 210 7725
rect 240 7695 245 7725
rect 205 7655 245 7695
rect 205 7625 210 7655
rect 240 7625 245 7655
rect 205 7620 245 7625
rect 405 7725 445 7730
rect 405 7695 410 7725
rect 440 7695 445 7725
rect 405 7655 445 7695
rect 405 7625 410 7655
rect 440 7625 445 7655
rect 405 7620 445 7625
rect 605 7725 645 7730
rect 605 7695 610 7725
rect 640 7695 645 7725
rect 605 7655 645 7695
rect 605 7625 610 7655
rect 640 7625 645 7655
rect 605 7620 645 7625
rect 805 7725 845 7730
rect 805 7695 810 7725
rect 840 7695 845 7725
rect 805 7655 845 7695
rect 805 7625 810 7655
rect 840 7625 845 7655
rect 805 7620 845 7625
rect 1005 7725 1045 7730
rect 1005 7695 1010 7725
rect 1040 7695 1045 7725
rect 1005 7655 1045 7695
rect 1005 7625 1010 7655
rect 1040 7625 1045 7655
rect 1005 7620 1045 7625
rect 1205 7725 1245 7730
rect 1205 7695 1210 7725
rect 1240 7695 1245 7725
rect 1205 7655 1245 7695
rect 1205 7625 1210 7655
rect 1240 7625 1245 7655
rect 1205 7620 1245 7625
rect 1405 7725 1445 7730
rect 1405 7695 1410 7725
rect 1440 7695 1445 7725
rect 1405 7655 1445 7695
rect 1405 7625 1410 7655
rect 1440 7625 1445 7655
rect 1405 7620 1445 7625
rect 1605 7725 1645 7730
rect 1605 7695 1610 7725
rect 1640 7695 1645 7725
rect 1605 7655 1645 7695
rect 1605 7625 1610 7655
rect 1640 7625 1645 7655
rect 1605 7620 1645 7625
rect 1805 7725 1845 7730
rect 1805 7695 1810 7725
rect 1840 7695 1845 7725
rect 1805 7655 1845 7695
rect 1805 7625 1810 7655
rect 1840 7625 1845 7655
rect 1805 7620 1845 7625
rect 2005 7725 2045 7730
rect 2005 7695 2010 7725
rect 2040 7695 2045 7725
rect 2005 7655 2045 7695
rect 2005 7625 2010 7655
rect 2040 7625 2045 7655
rect 2005 7620 2045 7625
rect 2205 7725 2245 7730
rect 2205 7695 2210 7725
rect 2240 7695 2245 7725
rect 2205 7655 2245 7695
rect 2205 7625 2210 7655
rect 2240 7625 2245 7655
rect 2205 7620 2245 7625
rect 2405 7725 2445 7730
rect 2405 7695 2410 7725
rect 2440 7695 2445 7725
rect 2405 7655 2445 7695
rect 2405 7625 2410 7655
rect 2440 7625 2445 7655
rect 2405 7620 2445 7625
rect 2605 7725 2645 7730
rect 2605 7695 2610 7725
rect 2640 7695 2645 7725
rect 2605 7655 2645 7695
rect 2605 7625 2610 7655
rect 2640 7625 2645 7655
rect 2605 7620 2645 7625
rect 2805 7725 2845 7730
rect 2805 7695 2810 7725
rect 2840 7695 2845 7725
rect 2805 7655 2845 7695
rect 2805 7625 2810 7655
rect 2840 7625 2845 7655
rect 2805 7620 2845 7625
rect 3005 7725 3045 7730
rect 3005 7695 3010 7725
rect 3040 7695 3045 7725
rect 3005 7655 3045 7695
rect 3005 7625 3010 7655
rect 3040 7625 3045 7655
rect 3005 7620 3045 7625
rect 3205 7725 3245 7730
rect 3205 7695 3210 7725
rect 3240 7695 3245 7725
rect 3205 7655 3245 7695
rect 3205 7625 3210 7655
rect 3240 7625 3245 7655
rect 3205 7620 3245 7625
rect 3405 7725 3445 7730
rect 3405 7695 3410 7725
rect 3440 7695 3445 7725
rect 3405 7655 3445 7695
rect 3405 7625 3410 7655
rect 3440 7625 3445 7655
rect 3405 7620 3445 7625
rect 3605 7725 3645 7730
rect 3605 7695 3610 7725
rect 3640 7695 3645 7725
rect 3605 7655 3645 7695
rect 3605 7625 3610 7655
rect 3640 7625 3645 7655
rect 3605 7620 3645 7625
rect 3805 7725 3845 7730
rect 3805 7695 3810 7725
rect 3840 7695 3845 7725
rect 3805 7655 3845 7695
rect 3805 7625 3810 7655
rect 3840 7625 3845 7655
rect 3805 7620 3845 7625
rect 4005 7725 4045 7730
rect 4005 7695 4010 7725
rect 4040 7695 4045 7725
rect 4005 7655 4045 7695
rect 4005 7625 4010 7655
rect 4040 7625 4045 7655
rect 4005 7620 4045 7625
rect 4205 7725 4245 7730
rect 4205 7695 4210 7725
rect 4240 7695 4245 7725
rect 4205 7655 4245 7695
rect 4205 7625 4210 7655
rect 4240 7625 4245 7655
rect 4205 7620 4245 7625
rect 4405 7725 4445 7730
rect 4405 7695 4410 7725
rect 4440 7695 4445 7725
rect 4405 7655 4445 7695
rect 4405 7625 4410 7655
rect 4440 7625 4445 7655
rect 4405 7620 4445 7625
rect 4605 7725 4645 7730
rect 4605 7695 4610 7725
rect 4640 7695 4645 7725
rect 4605 7655 4645 7695
rect 4605 7625 4610 7655
rect 4640 7625 4645 7655
rect 4605 7620 4645 7625
rect 4805 7725 4845 7730
rect 4805 7695 4810 7725
rect 4840 7695 4845 7725
rect 4805 7655 4845 7695
rect 4805 7625 4810 7655
rect 4840 7625 4845 7655
rect 4805 7620 4845 7625
rect 5005 7725 5045 7730
rect 5005 7695 5010 7725
rect 5040 7695 5045 7725
rect 5005 7655 5045 7695
rect 5005 7625 5010 7655
rect 5040 7625 5045 7655
rect 5005 7620 5045 7625
rect 5205 7725 5245 7730
rect 5205 7695 5210 7725
rect 5240 7695 5245 7725
rect 5205 7655 5245 7695
rect 5205 7625 5210 7655
rect 5240 7625 5245 7655
rect 5205 7620 5245 7625
rect 5405 7725 5445 7730
rect 5405 7695 5410 7725
rect 5440 7695 5445 7725
rect 5405 7655 5445 7695
rect 5405 7625 5410 7655
rect 5440 7625 5445 7655
rect 5405 7620 5445 7625
rect 5605 7725 5645 7730
rect 5605 7695 5610 7725
rect 5640 7695 5645 7725
rect 5605 7655 5645 7695
rect 5605 7625 5610 7655
rect 5640 7625 5645 7655
rect 5605 7620 5645 7625
rect 5805 7725 5845 7730
rect 5805 7695 5810 7725
rect 5840 7695 5845 7725
rect 5805 7655 5845 7695
rect 5805 7625 5810 7655
rect 5840 7625 5845 7655
rect 5805 7620 5845 7625
rect 6005 7725 6045 7730
rect 6005 7695 6010 7725
rect 6040 7695 6045 7725
rect 6005 7655 6045 7695
rect 6005 7625 6010 7655
rect 6040 7625 6045 7655
rect 6005 7620 6045 7625
rect 6205 7725 6245 7730
rect 6205 7695 6210 7725
rect 6240 7695 6245 7725
rect 6205 7655 6245 7695
rect 6205 7625 6210 7655
rect 6240 7625 6245 7655
rect 6205 7620 6245 7625
rect 6405 7725 6445 7730
rect 6405 7695 6410 7725
rect 6440 7695 6445 7725
rect 6405 7655 6445 7695
rect 6405 7625 6410 7655
rect 6440 7625 6445 7655
rect 6405 7620 6445 7625
rect -195 7540 -155 7545
rect -195 7510 -190 7540
rect -160 7510 -155 7540
rect -195 7470 -155 7510
rect -195 7440 -190 7470
rect -160 7440 -155 7470
rect -195 7435 -155 7440
rect 5 7540 45 7545
rect 5 7510 10 7540
rect 40 7510 45 7540
rect 5 7470 45 7510
rect 5 7440 10 7470
rect 40 7440 45 7470
rect 5 7435 45 7440
rect 205 7540 245 7545
rect 205 7510 210 7540
rect 240 7510 245 7540
rect 205 7470 245 7510
rect 205 7440 210 7470
rect 240 7440 245 7470
rect 205 7435 245 7440
rect 405 7540 445 7545
rect 405 7510 410 7540
rect 440 7510 445 7540
rect 405 7470 445 7510
rect 405 7440 410 7470
rect 440 7440 445 7470
rect 405 7435 445 7440
rect 605 7540 645 7545
rect 605 7510 610 7540
rect 640 7510 645 7540
rect 605 7470 645 7510
rect 605 7440 610 7470
rect 640 7440 645 7470
rect 605 7435 645 7440
rect 805 7540 845 7545
rect 805 7510 810 7540
rect 840 7510 845 7540
rect 805 7470 845 7510
rect 805 7440 810 7470
rect 840 7440 845 7470
rect 805 7435 845 7440
rect 1005 7540 1045 7545
rect 1005 7510 1010 7540
rect 1040 7510 1045 7540
rect 1005 7470 1045 7510
rect 1005 7440 1010 7470
rect 1040 7440 1045 7470
rect 1005 7435 1045 7440
rect 1205 7540 1245 7545
rect 1205 7510 1210 7540
rect 1240 7510 1245 7540
rect 1205 7470 1245 7510
rect 1205 7440 1210 7470
rect 1240 7440 1245 7470
rect 1205 7435 1245 7440
rect 1405 7540 1445 7545
rect 1405 7510 1410 7540
rect 1440 7510 1445 7540
rect 1405 7470 1445 7510
rect 1405 7440 1410 7470
rect 1440 7440 1445 7470
rect 1405 7435 1445 7440
rect 1605 7540 1645 7545
rect 1605 7510 1610 7540
rect 1640 7510 1645 7540
rect 1605 7470 1645 7510
rect 1605 7440 1610 7470
rect 1640 7440 1645 7470
rect 1605 7435 1645 7440
rect 1805 7540 1845 7545
rect 1805 7510 1810 7540
rect 1840 7510 1845 7540
rect 1805 7470 1845 7510
rect 1805 7440 1810 7470
rect 1840 7440 1845 7470
rect 1805 7435 1845 7440
rect 2005 7540 2045 7545
rect 2005 7510 2010 7540
rect 2040 7510 2045 7540
rect 2005 7470 2045 7510
rect 2005 7440 2010 7470
rect 2040 7440 2045 7470
rect 2005 7435 2045 7440
rect 2205 7540 2245 7545
rect 2205 7510 2210 7540
rect 2240 7510 2245 7540
rect 2205 7470 2245 7510
rect 2205 7440 2210 7470
rect 2240 7440 2245 7470
rect 2205 7435 2245 7440
rect 2405 7540 2445 7545
rect 2405 7510 2410 7540
rect 2440 7510 2445 7540
rect 2405 7470 2445 7510
rect 2405 7440 2410 7470
rect 2440 7440 2445 7470
rect 2405 7435 2445 7440
rect 2605 7540 2645 7545
rect 2605 7510 2610 7540
rect 2640 7510 2645 7540
rect 2605 7470 2645 7510
rect 2605 7440 2610 7470
rect 2640 7440 2645 7470
rect 2605 7435 2645 7440
rect 2805 7540 2845 7545
rect 2805 7510 2810 7540
rect 2840 7510 2845 7540
rect 2805 7470 2845 7510
rect 2805 7440 2810 7470
rect 2840 7440 2845 7470
rect 2805 7435 2845 7440
rect 3005 7540 3045 7545
rect 3005 7510 3010 7540
rect 3040 7510 3045 7540
rect 3005 7470 3045 7510
rect 3005 7440 3010 7470
rect 3040 7440 3045 7470
rect 3005 7435 3045 7440
rect 3205 7540 3245 7545
rect 3205 7510 3210 7540
rect 3240 7510 3245 7540
rect 3205 7470 3245 7510
rect 3205 7440 3210 7470
rect 3240 7440 3245 7470
rect 3205 7435 3245 7440
rect 3405 7540 3445 7545
rect 3405 7510 3410 7540
rect 3440 7510 3445 7540
rect 3405 7470 3445 7510
rect 3405 7440 3410 7470
rect 3440 7440 3445 7470
rect 3405 7435 3445 7440
rect 3605 7540 3645 7545
rect 3605 7510 3610 7540
rect 3640 7510 3645 7540
rect 3605 7470 3645 7510
rect 3605 7440 3610 7470
rect 3640 7440 3645 7470
rect 3605 7435 3645 7440
rect 3805 7540 3845 7545
rect 3805 7510 3810 7540
rect 3840 7510 3845 7540
rect 3805 7470 3845 7510
rect 3805 7440 3810 7470
rect 3840 7440 3845 7470
rect 3805 7435 3845 7440
rect 4005 7540 4045 7545
rect 4005 7510 4010 7540
rect 4040 7510 4045 7540
rect 4005 7470 4045 7510
rect 4005 7440 4010 7470
rect 4040 7440 4045 7470
rect 4005 7435 4045 7440
rect 4205 7540 4245 7545
rect 4205 7510 4210 7540
rect 4240 7510 4245 7540
rect 4205 7470 4245 7510
rect 4205 7440 4210 7470
rect 4240 7440 4245 7470
rect 4205 7435 4245 7440
rect 4405 7540 4445 7545
rect 4405 7510 4410 7540
rect 4440 7510 4445 7540
rect 4405 7470 4445 7510
rect 4405 7440 4410 7470
rect 4440 7440 4445 7470
rect 4405 7435 4445 7440
rect 4605 7540 4645 7545
rect 4605 7510 4610 7540
rect 4640 7510 4645 7540
rect 4605 7470 4645 7510
rect 4605 7440 4610 7470
rect 4640 7440 4645 7470
rect 4605 7435 4645 7440
rect 4805 7540 4845 7545
rect 4805 7510 4810 7540
rect 4840 7510 4845 7540
rect 4805 7470 4845 7510
rect 4805 7440 4810 7470
rect 4840 7440 4845 7470
rect 4805 7435 4845 7440
rect 5005 7540 5045 7545
rect 5005 7510 5010 7540
rect 5040 7510 5045 7540
rect 5005 7470 5045 7510
rect 5005 7440 5010 7470
rect 5040 7440 5045 7470
rect 5005 7435 5045 7440
rect 5205 7540 5245 7545
rect 5205 7510 5210 7540
rect 5240 7510 5245 7540
rect 5205 7470 5245 7510
rect 5205 7440 5210 7470
rect 5240 7440 5245 7470
rect 5205 7435 5245 7440
rect 5405 7540 5445 7545
rect 5405 7510 5410 7540
rect 5440 7510 5445 7540
rect 5405 7470 5445 7510
rect 5405 7440 5410 7470
rect 5440 7440 5445 7470
rect 5405 7435 5445 7440
rect 5605 7540 5645 7545
rect 5605 7510 5610 7540
rect 5640 7510 5645 7540
rect 5605 7470 5645 7510
rect 5605 7440 5610 7470
rect 5640 7440 5645 7470
rect 5605 7435 5645 7440
rect 5805 7540 5845 7545
rect 5805 7510 5810 7540
rect 5840 7510 5845 7540
rect 5805 7470 5845 7510
rect 5805 7440 5810 7470
rect 5840 7440 5845 7470
rect 5805 7435 5845 7440
rect 6005 7540 6045 7545
rect 6005 7510 6010 7540
rect 6040 7510 6045 7540
rect 6005 7470 6045 7510
rect 6005 7440 6010 7470
rect 6040 7440 6045 7470
rect 6005 7435 6045 7440
rect 6205 7540 6245 7545
rect 6205 7510 6210 7540
rect 6240 7510 6245 7540
rect 6205 7470 6245 7510
rect 6205 7440 6210 7470
rect 6240 7440 6245 7470
rect 6205 7435 6245 7440
rect 6405 7540 6445 7545
rect 6405 7510 6410 7540
rect 6440 7510 6445 7540
rect 6405 7470 6445 7510
rect 6405 7440 6410 7470
rect 6440 7440 6445 7470
rect 6405 7435 6445 7440
rect -195 7355 -155 7360
rect -195 7325 -190 7355
rect -160 7325 -155 7355
rect -195 7285 -155 7325
rect -195 7255 -190 7285
rect -160 7255 -155 7285
rect -195 7250 -155 7255
rect 5 7355 45 7360
rect 5 7325 10 7355
rect 40 7325 45 7355
rect 5 7285 45 7325
rect 5 7255 10 7285
rect 40 7255 45 7285
rect 5 7250 45 7255
rect 205 7355 245 7360
rect 205 7325 210 7355
rect 240 7325 245 7355
rect 205 7285 245 7325
rect 205 7255 210 7285
rect 240 7255 245 7285
rect 205 7250 245 7255
rect 405 7355 445 7360
rect 405 7325 410 7355
rect 440 7325 445 7355
rect 405 7285 445 7325
rect 405 7255 410 7285
rect 440 7255 445 7285
rect 405 7250 445 7255
rect 605 7355 645 7360
rect 605 7325 610 7355
rect 640 7325 645 7355
rect 605 7285 645 7325
rect 605 7255 610 7285
rect 640 7255 645 7285
rect 605 7250 645 7255
rect 805 7355 845 7360
rect 805 7325 810 7355
rect 840 7325 845 7355
rect 805 7285 845 7325
rect 805 7255 810 7285
rect 840 7255 845 7285
rect 805 7250 845 7255
rect 1005 7355 1045 7360
rect 1005 7325 1010 7355
rect 1040 7325 1045 7355
rect 1005 7285 1045 7325
rect 1005 7255 1010 7285
rect 1040 7255 1045 7285
rect 1005 7250 1045 7255
rect 1205 7355 1245 7360
rect 1205 7325 1210 7355
rect 1240 7325 1245 7355
rect 1205 7285 1245 7325
rect 1205 7255 1210 7285
rect 1240 7255 1245 7285
rect 1205 7250 1245 7255
rect 1405 7355 1445 7360
rect 1405 7325 1410 7355
rect 1440 7325 1445 7355
rect 1405 7285 1445 7325
rect 1405 7255 1410 7285
rect 1440 7255 1445 7285
rect 1405 7250 1445 7255
rect 1605 7355 1645 7360
rect 1605 7325 1610 7355
rect 1640 7325 1645 7355
rect 1605 7285 1645 7325
rect 1605 7255 1610 7285
rect 1640 7255 1645 7285
rect 1605 7250 1645 7255
rect 1805 7355 1845 7360
rect 1805 7325 1810 7355
rect 1840 7325 1845 7355
rect 1805 7285 1845 7325
rect 1805 7255 1810 7285
rect 1840 7255 1845 7285
rect 1805 7250 1845 7255
rect 2005 7355 2045 7360
rect 2005 7325 2010 7355
rect 2040 7325 2045 7355
rect 2005 7285 2045 7325
rect 2005 7255 2010 7285
rect 2040 7255 2045 7285
rect 2005 7250 2045 7255
rect 2205 7355 2245 7360
rect 2205 7325 2210 7355
rect 2240 7325 2245 7355
rect 2205 7285 2245 7325
rect 2205 7255 2210 7285
rect 2240 7255 2245 7285
rect 2205 7250 2245 7255
rect 2405 7355 2445 7360
rect 2405 7325 2410 7355
rect 2440 7325 2445 7355
rect 2405 7285 2445 7325
rect 2405 7255 2410 7285
rect 2440 7255 2445 7285
rect 2405 7250 2445 7255
rect 2605 7355 2645 7360
rect 2605 7325 2610 7355
rect 2640 7325 2645 7355
rect 2605 7285 2645 7325
rect 2605 7255 2610 7285
rect 2640 7255 2645 7285
rect 2605 7250 2645 7255
rect 2805 7355 2845 7360
rect 2805 7325 2810 7355
rect 2840 7325 2845 7355
rect 2805 7285 2845 7325
rect 2805 7255 2810 7285
rect 2840 7255 2845 7285
rect 2805 7250 2845 7255
rect 3005 7355 3045 7360
rect 3005 7325 3010 7355
rect 3040 7325 3045 7355
rect 3005 7285 3045 7325
rect 3005 7255 3010 7285
rect 3040 7255 3045 7285
rect 3005 7250 3045 7255
rect 3205 7355 3245 7360
rect 3205 7325 3210 7355
rect 3240 7325 3245 7355
rect 3205 7285 3245 7325
rect 3205 7255 3210 7285
rect 3240 7255 3245 7285
rect 3205 7250 3245 7255
rect 3405 7355 3445 7360
rect 3405 7325 3410 7355
rect 3440 7325 3445 7355
rect 3405 7285 3445 7325
rect 3405 7255 3410 7285
rect 3440 7255 3445 7285
rect 3405 7250 3445 7255
rect 3605 7355 3645 7360
rect 3605 7325 3610 7355
rect 3640 7325 3645 7355
rect 3605 7285 3645 7325
rect 3605 7255 3610 7285
rect 3640 7255 3645 7285
rect 3605 7250 3645 7255
rect 3805 7355 3845 7360
rect 3805 7325 3810 7355
rect 3840 7325 3845 7355
rect 3805 7285 3845 7325
rect 3805 7255 3810 7285
rect 3840 7255 3845 7285
rect 3805 7250 3845 7255
rect 4005 7355 4045 7360
rect 4005 7325 4010 7355
rect 4040 7325 4045 7355
rect 4005 7285 4045 7325
rect 4005 7255 4010 7285
rect 4040 7255 4045 7285
rect 4005 7250 4045 7255
rect 4205 7355 4245 7360
rect 4205 7325 4210 7355
rect 4240 7325 4245 7355
rect 4205 7285 4245 7325
rect 4205 7255 4210 7285
rect 4240 7255 4245 7285
rect 4205 7250 4245 7255
rect 4405 7355 4445 7360
rect 4405 7325 4410 7355
rect 4440 7325 4445 7355
rect 4405 7285 4445 7325
rect 4405 7255 4410 7285
rect 4440 7255 4445 7285
rect 4405 7250 4445 7255
rect 4605 7355 4645 7360
rect 4605 7325 4610 7355
rect 4640 7325 4645 7355
rect 4605 7285 4645 7325
rect 4605 7255 4610 7285
rect 4640 7255 4645 7285
rect 4605 7250 4645 7255
rect 4805 7355 4845 7360
rect 4805 7325 4810 7355
rect 4840 7325 4845 7355
rect 4805 7285 4845 7325
rect 4805 7255 4810 7285
rect 4840 7255 4845 7285
rect 4805 7250 4845 7255
rect 5005 7355 5045 7360
rect 5005 7325 5010 7355
rect 5040 7325 5045 7355
rect 5005 7285 5045 7325
rect 5005 7255 5010 7285
rect 5040 7255 5045 7285
rect 5005 7250 5045 7255
rect 5205 7355 5245 7360
rect 5205 7325 5210 7355
rect 5240 7325 5245 7355
rect 5205 7285 5245 7325
rect 5205 7255 5210 7285
rect 5240 7255 5245 7285
rect 5205 7250 5245 7255
rect 5405 7355 5445 7360
rect 5405 7325 5410 7355
rect 5440 7325 5445 7355
rect 5405 7285 5445 7325
rect 5405 7255 5410 7285
rect 5440 7255 5445 7285
rect 5405 7250 5445 7255
rect 5605 7355 5645 7360
rect 5605 7325 5610 7355
rect 5640 7325 5645 7355
rect 5605 7285 5645 7325
rect 5605 7255 5610 7285
rect 5640 7255 5645 7285
rect 5605 7250 5645 7255
rect 5805 7355 5845 7360
rect 5805 7325 5810 7355
rect 5840 7325 5845 7355
rect 5805 7285 5845 7325
rect 5805 7255 5810 7285
rect 5840 7255 5845 7285
rect 5805 7250 5845 7255
rect 6005 7355 6045 7360
rect 6005 7325 6010 7355
rect 6040 7325 6045 7355
rect 6005 7285 6045 7325
rect 6005 7255 6010 7285
rect 6040 7255 6045 7285
rect 6005 7250 6045 7255
rect 6205 7355 6245 7360
rect 6205 7325 6210 7355
rect 6240 7325 6245 7355
rect 6205 7285 6245 7325
rect 6205 7255 6210 7285
rect 6240 7255 6245 7285
rect 6205 7250 6245 7255
rect 6405 7355 6445 7360
rect 6405 7325 6410 7355
rect 6440 7325 6445 7355
rect 6405 7285 6445 7325
rect 6405 7255 6410 7285
rect 6440 7255 6445 7285
rect 6405 7250 6445 7255
rect -195 7170 -155 7175
rect -195 7140 -190 7170
rect -160 7140 -155 7170
rect -195 7100 -155 7140
rect -195 7070 -190 7100
rect -160 7070 -155 7100
rect -195 7065 -155 7070
rect 5 7170 45 7175
rect 5 7140 10 7170
rect 40 7140 45 7170
rect 5 7100 45 7140
rect 5 7070 10 7100
rect 40 7070 45 7100
rect 5 7065 45 7070
rect 205 7170 245 7175
rect 205 7140 210 7170
rect 240 7140 245 7170
rect 205 7100 245 7140
rect 205 7070 210 7100
rect 240 7070 245 7100
rect 205 7065 245 7070
rect 405 7170 445 7175
rect 405 7140 410 7170
rect 440 7140 445 7170
rect 405 7100 445 7140
rect 405 7070 410 7100
rect 440 7070 445 7100
rect 405 7065 445 7070
rect 605 7170 645 7175
rect 605 7140 610 7170
rect 640 7140 645 7170
rect 605 7100 645 7140
rect 605 7070 610 7100
rect 640 7070 645 7100
rect 605 7065 645 7070
rect 805 7170 845 7175
rect 805 7140 810 7170
rect 840 7140 845 7170
rect 805 7100 845 7140
rect 805 7070 810 7100
rect 840 7070 845 7100
rect 805 7065 845 7070
rect 1005 7170 1045 7175
rect 1005 7140 1010 7170
rect 1040 7140 1045 7170
rect 1005 7100 1045 7140
rect 1005 7070 1010 7100
rect 1040 7070 1045 7100
rect 1005 7065 1045 7070
rect 1205 7170 1245 7175
rect 1205 7140 1210 7170
rect 1240 7140 1245 7170
rect 1205 7100 1245 7140
rect 1205 7070 1210 7100
rect 1240 7070 1245 7100
rect 1205 7065 1245 7070
rect 1405 7170 1445 7175
rect 1405 7140 1410 7170
rect 1440 7140 1445 7170
rect 1405 7100 1445 7140
rect 1405 7070 1410 7100
rect 1440 7070 1445 7100
rect 1405 7065 1445 7070
rect 1605 7170 1645 7175
rect 1605 7140 1610 7170
rect 1640 7140 1645 7170
rect 1605 7100 1645 7140
rect 1605 7070 1610 7100
rect 1640 7070 1645 7100
rect 1605 7065 1645 7070
rect 1805 7170 1845 7175
rect 1805 7140 1810 7170
rect 1840 7140 1845 7170
rect 1805 7100 1845 7140
rect 1805 7070 1810 7100
rect 1840 7070 1845 7100
rect 1805 7065 1845 7070
rect 2005 7170 2045 7175
rect 2005 7140 2010 7170
rect 2040 7140 2045 7170
rect 2005 7100 2045 7140
rect 2005 7070 2010 7100
rect 2040 7070 2045 7100
rect 2005 7065 2045 7070
rect 2205 7170 2245 7175
rect 2205 7140 2210 7170
rect 2240 7140 2245 7170
rect 2205 7100 2245 7140
rect 2205 7070 2210 7100
rect 2240 7070 2245 7100
rect 2205 7065 2245 7070
rect 2405 7170 2445 7175
rect 2405 7140 2410 7170
rect 2440 7140 2445 7170
rect 2405 7100 2445 7140
rect 2405 7070 2410 7100
rect 2440 7070 2445 7100
rect 2405 7065 2445 7070
rect 2605 7170 2645 7175
rect 2605 7140 2610 7170
rect 2640 7140 2645 7170
rect 2605 7100 2645 7140
rect 2605 7070 2610 7100
rect 2640 7070 2645 7100
rect 2605 7065 2645 7070
rect 2805 7170 2845 7175
rect 2805 7140 2810 7170
rect 2840 7140 2845 7170
rect 2805 7100 2845 7140
rect 2805 7070 2810 7100
rect 2840 7070 2845 7100
rect 2805 7065 2845 7070
rect 3005 7170 3045 7175
rect 3005 7140 3010 7170
rect 3040 7140 3045 7170
rect 3005 7100 3045 7140
rect 3005 7070 3010 7100
rect 3040 7070 3045 7100
rect 3005 7065 3045 7070
rect 3205 7170 3245 7175
rect 3205 7140 3210 7170
rect 3240 7140 3245 7170
rect 3205 7100 3245 7140
rect 3205 7070 3210 7100
rect 3240 7070 3245 7100
rect 3205 7065 3245 7070
rect 3405 7170 3445 7175
rect 3405 7140 3410 7170
rect 3440 7140 3445 7170
rect 3405 7100 3445 7140
rect 3405 7070 3410 7100
rect 3440 7070 3445 7100
rect 3405 7065 3445 7070
rect 3605 7170 3645 7175
rect 3605 7140 3610 7170
rect 3640 7140 3645 7170
rect 3605 7100 3645 7140
rect 3605 7070 3610 7100
rect 3640 7070 3645 7100
rect 3605 7065 3645 7070
rect 3805 7170 3845 7175
rect 3805 7140 3810 7170
rect 3840 7140 3845 7170
rect 3805 7100 3845 7140
rect 3805 7070 3810 7100
rect 3840 7070 3845 7100
rect 3805 7065 3845 7070
rect 4005 7170 4045 7175
rect 4005 7140 4010 7170
rect 4040 7140 4045 7170
rect 4005 7100 4045 7140
rect 4005 7070 4010 7100
rect 4040 7070 4045 7100
rect 4005 7065 4045 7070
rect 4205 7170 4245 7175
rect 4205 7140 4210 7170
rect 4240 7140 4245 7170
rect 4205 7100 4245 7140
rect 4205 7070 4210 7100
rect 4240 7070 4245 7100
rect 4205 7065 4245 7070
rect 4405 7170 4445 7175
rect 4405 7140 4410 7170
rect 4440 7140 4445 7170
rect 4405 7100 4445 7140
rect 4405 7070 4410 7100
rect 4440 7070 4445 7100
rect 4405 7065 4445 7070
rect 4605 7170 4645 7175
rect 4605 7140 4610 7170
rect 4640 7140 4645 7170
rect 4605 7100 4645 7140
rect 4605 7070 4610 7100
rect 4640 7070 4645 7100
rect 4605 7065 4645 7070
rect 4805 7170 4845 7175
rect 4805 7140 4810 7170
rect 4840 7140 4845 7170
rect 4805 7100 4845 7140
rect 4805 7070 4810 7100
rect 4840 7070 4845 7100
rect 4805 7065 4845 7070
rect 5005 7170 5045 7175
rect 5005 7140 5010 7170
rect 5040 7140 5045 7170
rect 5005 7100 5045 7140
rect 5005 7070 5010 7100
rect 5040 7070 5045 7100
rect 5005 7065 5045 7070
rect 5205 7170 5245 7175
rect 5205 7140 5210 7170
rect 5240 7140 5245 7170
rect 5205 7100 5245 7140
rect 5205 7070 5210 7100
rect 5240 7070 5245 7100
rect 5205 7065 5245 7070
rect 5405 7170 5445 7175
rect 5405 7140 5410 7170
rect 5440 7140 5445 7170
rect 5405 7100 5445 7140
rect 5405 7070 5410 7100
rect 5440 7070 5445 7100
rect 5405 7065 5445 7070
rect 5605 7170 5645 7175
rect 5605 7140 5610 7170
rect 5640 7140 5645 7170
rect 5605 7100 5645 7140
rect 5605 7070 5610 7100
rect 5640 7070 5645 7100
rect 5605 7065 5645 7070
rect 5805 7170 5845 7175
rect 5805 7140 5810 7170
rect 5840 7140 5845 7170
rect 5805 7100 5845 7140
rect 5805 7070 5810 7100
rect 5840 7070 5845 7100
rect 5805 7065 5845 7070
rect 6005 7170 6045 7175
rect 6005 7140 6010 7170
rect 6040 7140 6045 7170
rect 6005 7100 6045 7140
rect 6005 7070 6010 7100
rect 6040 7070 6045 7100
rect 6005 7065 6045 7070
rect 6205 7170 6245 7175
rect 6205 7140 6210 7170
rect 6240 7140 6245 7170
rect 6205 7100 6245 7140
rect 6205 7070 6210 7100
rect 6240 7070 6245 7100
rect 6205 7065 6245 7070
rect 6405 7170 6445 7175
rect 6405 7140 6410 7170
rect 6440 7140 6445 7170
rect 6405 7100 6445 7140
rect 6405 7070 6410 7100
rect 6440 7070 6445 7100
rect 6405 7065 6445 7070
rect -195 6985 -155 6990
rect -195 6955 -190 6985
rect -160 6955 -155 6985
rect -195 6915 -155 6955
rect -195 6885 -190 6915
rect -160 6885 -155 6915
rect -195 6880 -155 6885
rect 5 6985 45 6990
rect 5 6955 10 6985
rect 40 6955 45 6985
rect 5 6915 45 6955
rect 5 6885 10 6915
rect 40 6885 45 6915
rect 5 6880 45 6885
rect 205 6985 245 6990
rect 205 6955 210 6985
rect 240 6955 245 6985
rect 205 6915 245 6955
rect 205 6885 210 6915
rect 240 6885 245 6915
rect 205 6880 245 6885
rect 405 6985 445 6990
rect 405 6955 410 6985
rect 440 6955 445 6985
rect 405 6915 445 6955
rect 405 6885 410 6915
rect 440 6885 445 6915
rect 405 6880 445 6885
rect 605 6985 645 6990
rect 605 6955 610 6985
rect 640 6955 645 6985
rect 605 6915 645 6955
rect 605 6885 610 6915
rect 640 6885 645 6915
rect 605 6880 645 6885
rect 805 6985 845 6990
rect 805 6955 810 6985
rect 840 6955 845 6985
rect 805 6915 845 6955
rect 805 6885 810 6915
rect 840 6885 845 6915
rect 805 6880 845 6885
rect 1005 6985 1045 6990
rect 1005 6955 1010 6985
rect 1040 6955 1045 6985
rect 1005 6915 1045 6955
rect 1005 6885 1010 6915
rect 1040 6885 1045 6915
rect 1005 6880 1045 6885
rect 1205 6985 1245 6990
rect 1205 6955 1210 6985
rect 1240 6955 1245 6985
rect 1205 6915 1245 6955
rect 1205 6885 1210 6915
rect 1240 6885 1245 6915
rect 1205 6880 1245 6885
rect 1405 6985 1445 6990
rect 1405 6955 1410 6985
rect 1440 6955 1445 6985
rect 1405 6915 1445 6955
rect 1405 6885 1410 6915
rect 1440 6885 1445 6915
rect 1405 6880 1445 6885
rect 1605 6985 1645 6990
rect 1605 6955 1610 6985
rect 1640 6955 1645 6985
rect 1605 6915 1645 6955
rect 1605 6885 1610 6915
rect 1640 6885 1645 6915
rect 1605 6880 1645 6885
rect 1805 6985 1845 6990
rect 1805 6955 1810 6985
rect 1840 6955 1845 6985
rect 1805 6915 1845 6955
rect 1805 6885 1810 6915
rect 1840 6885 1845 6915
rect 1805 6880 1845 6885
rect 2005 6985 2045 6990
rect 2005 6955 2010 6985
rect 2040 6955 2045 6985
rect 2005 6915 2045 6955
rect 2005 6885 2010 6915
rect 2040 6885 2045 6915
rect 2005 6880 2045 6885
rect 2205 6985 2245 6990
rect 2205 6955 2210 6985
rect 2240 6955 2245 6985
rect 2205 6915 2245 6955
rect 2205 6885 2210 6915
rect 2240 6885 2245 6915
rect 2205 6880 2245 6885
rect 2405 6985 2445 6990
rect 2405 6955 2410 6985
rect 2440 6955 2445 6985
rect 2405 6915 2445 6955
rect 2405 6885 2410 6915
rect 2440 6885 2445 6915
rect 2405 6880 2445 6885
rect 2605 6985 2645 6990
rect 2605 6955 2610 6985
rect 2640 6955 2645 6985
rect 2605 6915 2645 6955
rect 2605 6885 2610 6915
rect 2640 6885 2645 6915
rect 2605 6880 2645 6885
rect 2805 6985 2845 6990
rect 2805 6955 2810 6985
rect 2840 6955 2845 6985
rect 2805 6915 2845 6955
rect 2805 6885 2810 6915
rect 2840 6885 2845 6915
rect 2805 6880 2845 6885
rect 3005 6985 3045 6990
rect 3005 6955 3010 6985
rect 3040 6955 3045 6985
rect 3005 6915 3045 6955
rect 3005 6885 3010 6915
rect 3040 6885 3045 6915
rect 3005 6880 3045 6885
rect 3205 6985 3245 6990
rect 3205 6955 3210 6985
rect 3240 6955 3245 6985
rect 3205 6915 3245 6955
rect 3205 6885 3210 6915
rect 3240 6885 3245 6915
rect 3205 6880 3245 6885
rect 3405 6985 3445 6990
rect 3405 6955 3410 6985
rect 3440 6955 3445 6985
rect 3405 6915 3445 6955
rect 3405 6885 3410 6915
rect 3440 6885 3445 6915
rect 3405 6880 3445 6885
rect 3605 6985 3645 6990
rect 3605 6955 3610 6985
rect 3640 6955 3645 6985
rect 3605 6915 3645 6955
rect 3605 6885 3610 6915
rect 3640 6885 3645 6915
rect 3605 6880 3645 6885
rect 3805 6985 3845 6990
rect 3805 6955 3810 6985
rect 3840 6955 3845 6985
rect 3805 6915 3845 6955
rect 3805 6885 3810 6915
rect 3840 6885 3845 6915
rect 3805 6880 3845 6885
rect 4005 6985 4045 6990
rect 4005 6955 4010 6985
rect 4040 6955 4045 6985
rect 4005 6915 4045 6955
rect 4005 6885 4010 6915
rect 4040 6885 4045 6915
rect 4005 6880 4045 6885
rect 4205 6985 4245 6990
rect 4205 6955 4210 6985
rect 4240 6955 4245 6985
rect 4205 6915 4245 6955
rect 4205 6885 4210 6915
rect 4240 6885 4245 6915
rect 4205 6880 4245 6885
rect 4405 6985 4445 6990
rect 4405 6955 4410 6985
rect 4440 6955 4445 6985
rect 4405 6915 4445 6955
rect 4405 6885 4410 6915
rect 4440 6885 4445 6915
rect 4405 6880 4445 6885
rect 4605 6985 4645 6990
rect 4605 6955 4610 6985
rect 4640 6955 4645 6985
rect 4605 6915 4645 6955
rect 4605 6885 4610 6915
rect 4640 6885 4645 6915
rect 4605 6880 4645 6885
rect 4805 6985 4845 6990
rect 4805 6955 4810 6985
rect 4840 6955 4845 6985
rect 4805 6915 4845 6955
rect 4805 6885 4810 6915
rect 4840 6885 4845 6915
rect 4805 6880 4845 6885
rect 5005 6985 5045 6990
rect 5005 6955 5010 6985
rect 5040 6955 5045 6985
rect 5005 6915 5045 6955
rect 5005 6885 5010 6915
rect 5040 6885 5045 6915
rect 5005 6880 5045 6885
rect 5205 6985 5245 6990
rect 5205 6955 5210 6985
rect 5240 6955 5245 6985
rect 5205 6915 5245 6955
rect 5205 6885 5210 6915
rect 5240 6885 5245 6915
rect 5205 6880 5245 6885
rect 5405 6985 5445 6990
rect 5405 6955 5410 6985
rect 5440 6955 5445 6985
rect 5405 6915 5445 6955
rect 5405 6885 5410 6915
rect 5440 6885 5445 6915
rect 5405 6880 5445 6885
rect 5605 6985 5645 6990
rect 5605 6955 5610 6985
rect 5640 6955 5645 6985
rect 5605 6915 5645 6955
rect 5605 6885 5610 6915
rect 5640 6885 5645 6915
rect 5605 6880 5645 6885
rect 5805 6985 5845 6990
rect 5805 6955 5810 6985
rect 5840 6955 5845 6985
rect 5805 6915 5845 6955
rect 5805 6885 5810 6915
rect 5840 6885 5845 6915
rect 5805 6880 5845 6885
rect 6005 6985 6045 6990
rect 6005 6955 6010 6985
rect 6040 6955 6045 6985
rect 6005 6915 6045 6955
rect 6005 6885 6010 6915
rect 6040 6885 6045 6915
rect 6005 6880 6045 6885
rect 6205 6985 6245 6990
rect 6205 6955 6210 6985
rect 6240 6955 6245 6985
rect 6205 6915 6245 6955
rect 6205 6885 6210 6915
rect 6240 6885 6245 6915
rect 6205 6880 6245 6885
rect 6405 6985 6445 6990
rect 6405 6955 6410 6985
rect 6440 6955 6445 6985
rect 6405 6915 6445 6955
rect 6405 6885 6410 6915
rect 6440 6885 6445 6915
rect 6405 6880 6445 6885
rect -195 6800 -155 6805
rect -195 6770 -190 6800
rect -160 6770 -155 6800
rect -195 6730 -155 6770
rect -195 6700 -190 6730
rect -160 6700 -155 6730
rect -195 6695 -155 6700
rect 5 6800 45 6805
rect 5 6770 10 6800
rect 40 6770 45 6800
rect 5 6730 45 6770
rect 5 6700 10 6730
rect 40 6700 45 6730
rect 5 6695 45 6700
rect 205 6800 245 6805
rect 205 6770 210 6800
rect 240 6770 245 6800
rect 205 6730 245 6770
rect 205 6700 210 6730
rect 240 6700 245 6730
rect 205 6695 245 6700
rect 405 6800 445 6805
rect 405 6770 410 6800
rect 440 6770 445 6800
rect 405 6730 445 6770
rect 405 6700 410 6730
rect 440 6700 445 6730
rect 405 6695 445 6700
rect 605 6800 645 6805
rect 605 6770 610 6800
rect 640 6770 645 6800
rect 605 6730 645 6770
rect 605 6700 610 6730
rect 640 6700 645 6730
rect 605 6695 645 6700
rect 805 6800 845 6805
rect 805 6770 810 6800
rect 840 6770 845 6800
rect 805 6730 845 6770
rect 805 6700 810 6730
rect 840 6700 845 6730
rect 805 6695 845 6700
rect 1005 6800 1045 6805
rect 1005 6770 1010 6800
rect 1040 6770 1045 6800
rect 1005 6730 1045 6770
rect 1005 6700 1010 6730
rect 1040 6700 1045 6730
rect 1005 6695 1045 6700
rect 1205 6800 1245 6805
rect 1205 6770 1210 6800
rect 1240 6770 1245 6800
rect 1205 6730 1245 6770
rect 1205 6700 1210 6730
rect 1240 6700 1245 6730
rect 1205 6695 1245 6700
rect 1405 6800 1445 6805
rect 1405 6770 1410 6800
rect 1440 6770 1445 6800
rect 1405 6730 1445 6770
rect 1405 6700 1410 6730
rect 1440 6700 1445 6730
rect 1405 6695 1445 6700
rect 1605 6800 1645 6805
rect 1605 6770 1610 6800
rect 1640 6770 1645 6800
rect 1605 6730 1645 6770
rect 1605 6700 1610 6730
rect 1640 6700 1645 6730
rect 1605 6695 1645 6700
rect 1805 6800 1845 6805
rect 1805 6770 1810 6800
rect 1840 6770 1845 6800
rect 1805 6730 1845 6770
rect 1805 6700 1810 6730
rect 1840 6700 1845 6730
rect 1805 6695 1845 6700
rect 2005 6800 2045 6805
rect 2005 6770 2010 6800
rect 2040 6770 2045 6800
rect 2005 6730 2045 6770
rect 2005 6700 2010 6730
rect 2040 6700 2045 6730
rect 2005 6695 2045 6700
rect 2205 6800 2245 6805
rect 2205 6770 2210 6800
rect 2240 6770 2245 6800
rect 2205 6730 2245 6770
rect 2205 6700 2210 6730
rect 2240 6700 2245 6730
rect 2205 6695 2245 6700
rect 2405 6800 2445 6805
rect 2405 6770 2410 6800
rect 2440 6770 2445 6800
rect 2405 6730 2445 6770
rect 2405 6700 2410 6730
rect 2440 6700 2445 6730
rect 2405 6695 2445 6700
rect 2605 6800 2645 6805
rect 2605 6770 2610 6800
rect 2640 6770 2645 6800
rect 2605 6730 2645 6770
rect 2605 6700 2610 6730
rect 2640 6700 2645 6730
rect 2605 6695 2645 6700
rect 2805 6800 2845 6805
rect 2805 6770 2810 6800
rect 2840 6770 2845 6800
rect 2805 6730 2845 6770
rect 2805 6700 2810 6730
rect 2840 6700 2845 6730
rect 2805 6695 2845 6700
rect 3005 6800 3045 6805
rect 3005 6770 3010 6800
rect 3040 6770 3045 6800
rect 3005 6730 3045 6770
rect 3005 6700 3010 6730
rect 3040 6700 3045 6730
rect 3005 6695 3045 6700
rect 3205 6800 3245 6805
rect 3205 6770 3210 6800
rect 3240 6770 3245 6800
rect 3205 6730 3245 6770
rect 3205 6700 3210 6730
rect 3240 6700 3245 6730
rect 3205 6695 3245 6700
rect 3405 6800 3445 6805
rect 3405 6770 3410 6800
rect 3440 6770 3445 6800
rect 3405 6730 3445 6770
rect 3405 6700 3410 6730
rect 3440 6700 3445 6730
rect 3405 6695 3445 6700
rect 3605 6800 3645 6805
rect 3605 6770 3610 6800
rect 3640 6770 3645 6800
rect 3605 6730 3645 6770
rect 3605 6700 3610 6730
rect 3640 6700 3645 6730
rect 3605 6695 3645 6700
rect 3805 6800 3845 6805
rect 3805 6770 3810 6800
rect 3840 6770 3845 6800
rect 3805 6730 3845 6770
rect 3805 6700 3810 6730
rect 3840 6700 3845 6730
rect 3805 6695 3845 6700
rect 4005 6800 4045 6805
rect 4005 6770 4010 6800
rect 4040 6770 4045 6800
rect 4005 6730 4045 6770
rect 4005 6700 4010 6730
rect 4040 6700 4045 6730
rect 4005 6695 4045 6700
rect 4205 6800 4245 6805
rect 4205 6770 4210 6800
rect 4240 6770 4245 6800
rect 4205 6730 4245 6770
rect 4205 6700 4210 6730
rect 4240 6700 4245 6730
rect 4205 6695 4245 6700
rect 4405 6800 4445 6805
rect 4405 6770 4410 6800
rect 4440 6770 4445 6800
rect 4405 6730 4445 6770
rect 4405 6700 4410 6730
rect 4440 6700 4445 6730
rect 4405 6695 4445 6700
rect 4605 6800 4645 6805
rect 4605 6770 4610 6800
rect 4640 6770 4645 6800
rect 4605 6730 4645 6770
rect 4605 6700 4610 6730
rect 4640 6700 4645 6730
rect 4605 6695 4645 6700
rect 4805 6800 4845 6805
rect 4805 6770 4810 6800
rect 4840 6770 4845 6800
rect 4805 6730 4845 6770
rect 4805 6700 4810 6730
rect 4840 6700 4845 6730
rect 4805 6695 4845 6700
rect 5005 6800 5045 6805
rect 5005 6770 5010 6800
rect 5040 6770 5045 6800
rect 5005 6730 5045 6770
rect 5005 6700 5010 6730
rect 5040 6700 5045 6730
rect 5005 6695 5045 6700
rect 5205 6800 5245 6805
rect 5205 6770 5210 6800
rect 5240 6770 5245 6800
rect 5205 6730 5245 6770
rect 5205 6700 5210 6730
rect 5240 6700 5245 6730
rect 5205 6695 5245 6700
rect 5405 6800 5445 6805
rect 5405 6770 5410 6800
rect 5440 6770 5445 6800
rect 5405 6730 5445 6770
rect 5405 6700 5410 6730
rect 5440 6700 5445 6730
rect 5405 6695 5445 6700
rect 5605 6800 5645 6805
rect 5605 6770 5610 6800
rect 5640 6770 5645 6800
rect 5605 6730 5645 6770
rect 5605 6700 5610 6730
rect 5640 6700 5645 6730
rect 5605 6695 5645 6700
rect 5805 6800 5845 6805
rect 5805 6770 5810 6800
rect 5840 6770 5845 6800
rect 5805 6730 5845 6770
rect 5805 6700 5810 6730
rect 5840 6700 5845 6730
rect 5805 6695 5845 6700
rect 6005 6800 6045 6805
rect 6005 6770 6010 6800
rect 6040 6770 6045 6800
rect 6005 6730 6045 6770
rect 6005 6700 6010 6730
rect 6040 6700 6045 6730
rect 6005 6695 6045 6700
rect 6205 6800 6245 6805
rect 6205 6770 6210 6800
rect 6240 6770 6245 6800
rect 6205 6730 6245 6770
rect 6205 6700 6210 6730
rect 6240 6700 6245 6730
rect 6205 6695 6245 6700
rect 6405 6800 6445 6805
rect 6405 6770 6410 6800
rect 6440 6770 6445 6800
rect 6405 6730 6445 6770
rect 6405 6700 6410 6730
rect 6440 6700 6445 6730
rect 6405 6695 6445 6700
rect -195 6615 -155 6620
rect -195 6585 -190 6615
rect -160 6585 -155 6615
rect -195 6545 -155 6585
rect -195 6515 -190 6545
rect -160 6515 -155 6545
rect -195 6510 -155 6515
rect 5 6615 45 6620
rect 5 6585 10 6615
rect 40 6585 45 6615
rect 5 6545 45 6585
rect 5 6515 10 6545
rect 40 6515 45 6545
rect 5 6510 45 6515
rect 205 6615 245 6620
rect 205 6585 210 6615
rect 240 6585 245 6615
rect 205 6545 245 6585
rect 205 6515 210 6545
rect 240 6515 245 6545
rect 205 6510 245 6515
rect 405 6615 445 6620
rect 405 6585 410 6615
rect 440 6585 445 6615
rect 405 6545 445 6585
rect 405 6515 410 6545
rect 440 6515 445 6545
rect 405 6510 445 6515
rect 605 6615 645 6620
rect 605 6585 610 6615
rect 640 6585 645 6615
rect 605 6545 645 6585
rect 605 6515 610 6545
rect 640 6515 645 6545
rect 605 6510 645 6515
rect 805 6615 845 6620
rect 805 6585 810 6615
rect 840 6585 845 6615
rect 805 6545 845 6585
rect 805 6515 810 6545
rect 840 6515 845 6545
rect 805 6510 845 6515
rect 1005 6615 1045 6620
rect 1005 6585 1010 6615
rect 1040 6585 1045 6615
rect 1005 6545 1045 6585
rect 1005 6515 1010 6545
rect 1040 6515 1045 6545
rect 1005 6510 1045 6515
rect 1205 6615 1245 6620
rect 1205 6585 1210 6615
rect 1240 6585 1245 6615
rect 1205 6545 1245 6585
rect 1205 6515 1210 6545
rect 1240 6515 1245 6545
rect 1205 6510 1245 6515
rect 1405 6615 1445 6620
rect 1405 6585 1410 6615
rect 1440 6585 1445 6615
rect 1405 6545 1445 6585
rect 1405 6515 1410 6545
rect 1440 6515 1445 6545
rect 1405 6510 1445 6515
rect 1605 6615 1645 6620
rect 1605 6585 1610 6615
rect 1640 6585 1645 6615
rect 1605 6545 1645 6585
rect 1605 6515 1610 6545
rect 1640 6515 1645 6545
rect 1605 6510 1645 6515
rect 1805 6615 1845 6620
rect 1805 6585 1810 6615
rect 1840 6585 1845 6615
rect 1805 6545 1845 6585
rect 1805 6515 1810 6545
rect 1840 6515 1845 6545
rect 1805 6510 1845 6515
rect 2005 6615 2045 6620
rect 2005 6585 2010 6615
rect 2040 6585 2045 6615
rect 2005 6545 2045 6585
rect 2005 6515 2010 6545
rect 2040 6515 2045 6545
rect 2005 6510 2045 6515
rect 2205 6615 2245 6620
rect 2205 6585 2210 6615
rect 2240 6585 2245 6615
rect 2205 6545 2245 6585
rect 2205 6515 2210 6545
rect 2240 6515 2245 6545
rect 2205 6510 2245 6515
rect 2405 6615 2445 6620
rect 2405 6585 2410 6615
rect 2440 6585 2445 6615
rect 2405 6545 2445 6585
rect 2405 6515 2410 6545
rect 2440 6515 2445 6545
rect 2405 6510 2445 6515
rect 2605 6615 2645 6620
rect 2605 6585 2610 6615
rect 2640 6585 2645 6615
rect 2605 6545 2645 6585
rect 2605 6515 2610 6545
rect 2640 6515 2645 6545
rect 2605 6510 2645 6515
rect 2805 6615 2845 6620
rect 2805 6585 2810 6615
rect 2840 6585 2845 6615
rect 2805 6545 2845 6585
rect 2805 6515 2810 6545
rect 2840 6515 2845 6545
rect 2805 6510 2845 6515
rect 3005 6615 3045 6620
rect 3005 6585 3010 6615
rect 3040 6585 3045 6615
rect 3005 6545 3045 6585
rect 3005 6515 3010 6545
rect 3040 6515 3045 6545
rect 3005 6510 3045 6515
rect 3205 6615 3245 6620
rect 3205 6585 3210 6615
rect 3240 6585 3245 6615
rect 3205 6545 3245 6585
rect 3205 6515 3210 6545
rect 3240 6515 3245 6545
rect 3205 6510 3245 6515
rect 3405 6615 3445 6620
rect 3405 6585 3410 6615
rect 3440 6585 3445 6615
rect 3405 6545 3445 6585
rect 3405 6515 3410 6545
rect 3440 6515 3445 6545
rect 3405 6510 3445 6515
rect 3605 6615 3645 6620
rect 3605 6585 3610 6615
rect 3640 6585 3645 6615
rect 3605 6545 3645 6585
rect 3605 6515 3610 6545
rect 3640 6515 3645 6545
rect 3605 6510 3645 6515
rect 3805 6615 3845 6620
rect 3805 6585 3810 6615
rect 3840 6585 3845 6615
rect 3805 6545 3845 6585
rect 3805 6515 3810 6545
rect 3840 6515 3845 6545
rect 3805 6510 3845 6515
rect 4005 6615 4045 6620
rect 4005 6585 4010 6615
rect 4040 6585 4045 6615
rect 4005 6545 4045 6585
rect 4005 6515 4010 6545
rect 4040 6515 4045 6545
rect 4005 6510 4045 6515
rect 4205 6615 4245 6620
rect 4205 6585 4210 6615
rect 4240 6585 4245 6615
rect 4205 6545 4245 6585
rect 4205 6515 4210 6545
rect 4240 6515 4245 6545
rect 4205 6510 4245 6515
rect 4405 6615 4445 6620
rect 4405 6585 4410 6615
rect 4440 6585 4445 6615
rect 4405 6545 4445 6585
rect 4405 6515 4410 6545
rect 4440 6515 4445 6545
rect 4405 6510 4445 6515
rect 4605 6615 4645 6620
rect 4605 6585 4610 6615
rect 4640 6585 4645 6615
rect 4605 6545 4645 6585
rect 4605 6515 4610 6545
rect 4640 6515 4645 6545
rect 4605 6510 4645 6515
rect 4805 6615 4845 6620
rect 4805 6585 4810 6615
rect 4840 6585 4845 6615
rect 4805 6545 4845 6585
rect 4805 6515 4810 6545
rect 4840 6515 4845 6545
rect 4805 6510 4845 6515
rect 5005 6615 5045 6620
rect 5005 6585 5010 6615
rect 5040 6585 5045 6615
rect 5005 6545 5045 6585
rect 5005 6515 5010 6545
rect 5040 6515 5045 6545
rect 5005 6510 5045 6515
rect 5205 6615 5245 6620
rect 5205 6585 5210 6615
rect 5240 6585 5245 6615
rect 5205 6545 5245 6585
rect 5205 6515 5210 6545
rect 5240 6515 5245 6545
rect 5205 6510 5245 6515
rect 5405 6615 5445 6620
rect 5405 6585 5410 6615
rect 5440 6585 5445 6615
rect 5405 6545 5445 6585
rect 5405 6515 5410 6545
rect 5440 6515 5445 6545
rect 5405 6510 5445 6515
rect 5605 6615 5645 6620
rect 5605 6585 5610 6615
rect 5640 6585 5645 6615
rect 5605 6545 5645 6585
rect 5605 6515 5610 6545
rect 5640 6515 5645 6545
rect 5605 6510 5645 6515
rect 5805 6615 5845 6620
rect 5805 6585 5810 6615
rect 5840 6585 5845 6615
rect 5805 6545 5845 6585
rect 5805 6515 5810 6545
rect 5840 6515 5845 6545
rect 5805 6510 5845 6515
rect 6005 6615 6045 6620
rect 6005 6585 6010 6615
rect 6040 6585 6045 6615
rect 6005 6545 6045 6585
rect 6005 6515 6010 6545
rect 6040 6515 6045 6545
rect 6005 6510 6045 6515
rect 6205 6615 6245 6620
rect 6205 6585 6210 6615
rect 6240 6585 6245 6615
rect 6205 6545 6245 6585
rect 6205 6515 6210 6545
rect 6240 6515 6245 6545
rect 6205 6510 6245 6515
rect 6405 6615 6445 6620
rect 6405 6585 6410 6615
rect 6440 6585 6445 6615
rect 6405 6545 6445 6585
rect 6405 6515 6410 6545
rect 6440 6515 6445 6545
rect 6405 6510 6445 6515
rect -195 6430 -155 6435
rect -195 6400 -190 6430
rect -160 6400 -155 6430
rect -195 6360 -155 6400
rect -195 6330 -190 6360
rect -160 6330 -155 6360
rect -195 6325 -155 6330
rect 5 6430 45 6435
rect 5 6400 10 6430
rect 40 6400 45 6430
rect 5 6360 45 6400
rect 5 6330 10 6360
rect 40 6330 45 6360
rect 5 6325 45 6330
rect 205 6430 245 6435
rect 205 6400 210 6430
rect 240 6400 245 6430
rect 205 6360 245 6400
rect 205 6330 210 6360
rect 240 6330 245 6360
rect 205 6325 245 6330
rect 405 6430 445 6435
rect 405 6400 410 6430
rect 440 6400 445 6430
rect 405 6360 445 6400
rect 405 6330 410 6360
rect 440 6330 445 6360
rect 405 6325 445 6330
rect 605 6430 645 6435
rect 605 6400 610 6430
rect 640 6400 645 6430
rect 605 6360 645 6400
rect 605 6330 610 6360
rect 640 6330 645 6360
rect 605 6325 645 6330
rect 805 6430 845 6435
rect 805 6400 810 6430
rect 840 6400 845 6430
rect 805 6360 845 6400
rect 805 6330 810 6360
rect 840 6330 845 6360
rect 805 6325 845 6330
rect 1005 6430 1045 6435
rect 1005 6400 1010 6430
rect 1040 6400 1045 6430
rect 1005 6360 1045 6400
rect 1005 6330 1010 6360
rect 1040 6330 1045 6360
rect 1005 6325 1045 6330
rect 1205 6430 1245 6435
rect 1205 6400 1210 6430
rect 1240 6400 1245 6430
rect 1205 6360 1245 6400
rect 1205 6330 1210 6360
rect 1240 6330 1245 6360
rect 1205 6325 1245 6330
rect 1405 6430 1445 6435
rect 1405 6400 1410 6430
rect 1440 6400 1445 6430
rect 1405 6360 1445 6400
rect 1405 6330 1410 6360
rect 1440 6330 1445 6360
rect 1405 6325 1445 6330
rect 1605 6430 1645 6435
rect 1605 6400 1610 6430
rect 1640 6400 1645 6430
rect 1605 6360 1645 6400
rect 1605 6330 1610 6360
rect 1640 6330 1645 6360
rect 1605 6325 1645 6330
rect 1805 6430 1845 6435
rect 1805 6400 1810 6430
rect 1840 6400 1845 6430
rect 1805 6360 1845 6400
rect 1805 6330 1810 6360
rect 1840 6330 1845 6360
rect 1805 6325 1845 6330
rect 2005 6430 2045 6435
rect 2005 6400 2010 6430
rect 2040 6400 2045 6430
rect 2005 6360 2045 6400
rect 2005 6330 2010 6360
rect 2040 6330 2045 6360
rect 2005 6325 2045 6330
rect 2205 6430 2245 6435
rect 2205 6400 2210 6430
rect 2240 6400 2245 6430
rect 2205 6360 2245 6400
rect 2205 6330 2210 6360
rect 2240 6330 2245 6360
rect 2205 6325 2245 6330
rect 2405 6430 2445 6435
rect 2405 6400 2410 6430
rect 2440 6400 2445 6430
rect 2405 6360 2445 6400
rect 2405 6330 2410 6360
rect 2440 6330 2445 6360
rect 2405 6325 2445 6330
rect 2605 6430 2645 6435
rect 2605 6400 2610 6430
rect 2640 6400 2645 6430
rect 2605 6360 2645 6400
rect 2605 6330 2610 6360
rect 2640 6330 2645 6360
rect 2605 6325 2645 6330
rect 2805 6430 2845 6435
rect 2805 6400 2810 6430
rect 2840 6400 2845 6430
rect 2805 6360 2845 6400
rect 2805 6330 2810 6360
rect 2840 6330 2845 6360
rect 2805 6325 2845 6330
rect 3005 6430 3045 6435
rect 3005 6400 3010 6430
rect 3040 6400 3045 6430
rect 3005 6360 3045 6400
rect 3005 6330 3010 6360
rect 3040 6330 3045 6360
rect 3005 6325 3045 6330
rect 3205 6430 3245 6435
rect 3205 6400 3210 6430
rect 3240 6400 3245 6430
rect 3205 6360 3245 6400
rect 3205 6330 3210 6360
rect 3240 6330 3245 6360
rect 3205 6325 3245 6330
rect 3405 6430 3445 6435
rect 3405 6400 3410 6430
rect 3440 6400 3445 6430
rect 3405 6360 3445 6400
rect 3405 6330 3410 6360
rect 3440 6330 3445 6360
rect 3405 6325 3445 6330
rect 3605 6430 3645 6435
rect 3605 6400 3610 6430
rect 3640 6400 3645 6430
rect 3605 6360 3645 6400
rect 3605 6330 3610 6360
rect 3640 6330 3645 6360
rect 3605 6325 3645 6330
rect 3805 6430 3845 6435
rect 3805 6400 3810 6430
rect 3840 6400 3845 6430
rect 3805 6360 3845 6400
rect 3805 6330 3810 6360
rect 3840 6330 3845 6360
rect 3805 6325 3845 6330
rect 4005 6430 4045 6435
rect 4005 6400 4010 6430
rect 4040 6400 4045 6430
rect 4005 6360 4045 6400
rect 4005 6330 4010 6360
rect 4040 6330 4045 6360
rect 4005 6325 4045 6330
rect 4205 6430 4245 6435
rect 4205 6400 4210 6430
rect 4240 6400 4245 6430
rect 4205 6360 4245 6400
rect 4205 6330 4210 6360
rect 4240 6330 4245 6360
rect 4205 6325 4245 6330
rect 4405 6430 4445 6435
rect 4405 6400 4410 6430
rect 4440 6400 4445 6430
rect 4405 6360 4445 6400
rect 4405 6330 4410 6360
rect 4440 6330 4445 6360
rect 4405 6325 4445 6330
rect 4605 6430 4645 6435
rect 4605 6400 4610 6430
rect 4640 6400 4645 6430
rect 4605 6360 4645 6400
rect 4605 6330 4610 6360
rect 4640 6330 4645 6360
rect 4605 6325 4645 6330
rect 4805 6430 4845 6435
rect 4805 6400 4810 6430
rect 4840 6400 4845 6430
rect 4805 6360 4845 6400
rect 4805 6330 4810 6360
rect 4840 6330 4845 6360
rect 4805 6325 4845 6330
rect 5005 6430 5045 6435
rect 5005 6400 5010 6430
rect 5040 6400 5045 6430
rect 5005 6360 5045 6400
rect 5005 6330 5010 6360
rect 5040 6330 5045 6360
rect 5005 6325 5045 6330
rect 5205 6430 5245 6435
rect 5205 6400 5210 6430
rect 5240 6400 5245 6430
rect 5205 6360 5245 6400
rect 5205 6330 5210 6360
rect 5240 6330 5245 6360
rect 5205 6325 5245 6330
rect 5405 6430 5445 6435
rect 5405 6400 5410 6430
rect 5440 6400 5445 6430
rect 5405 6360 5445 6400
rect 5405 6330 5410 6360
rect 5440 6330 5445 6360
rect 5405 6325 5445 6330
rect 5605 6430 5645 6435
rect 5605 6400 5610 6430
rect 5640 6400 5645 6430
rect 5605 6360 5645 6400
rect 5605 6330 5610 6360
rect 5640 6330 5645 6360
rect 5605 6325 5645 6330
rect 5805 6430 5845 6435
rect 5805 6400 5810 6430
rect 5840 6400 5845 6430
rect 5805 6360 5845 6400
rect 5805 6330 5810 6360
rect 5840 6330 5845 6360
rect 5805 6325 5845 6330
rect 6005 6430 6045 6435
rect 6005 6400 6010 6430
rect 6040 6400 6045 6430
rect 6005 6360 6045 6400
rect 6005 6330 6010 6360
rect 6040 6330 6045 6360
rect 6005 6325 6045 6330
rect 6205 6430 6245 6435
rect 6205 6400 6210 6430
rect 6240 6400 6245 6430
rect 6205 6360 6245 6400
rect 6205 6330 6210 6360
rect 6240 6330 6245 6360
rect 6205 6325 6245 6330
rect 6405 6430 6445 6435
rect 6405 6400 6410 6430
rect 6440 6400 6445 6430
rect 6405 6360 6445 6400
rect 6405 6330 6410 6360
rect 6440 6330 6445 6360
rect 6405 6325 6445 6330
rect -195 6245 -155 6250
rect -195 6215 -190 6245
rect -160 6215 -155 6245
rect -195 6175 -155 6215
rect -195 6145 -190 6175
rect -160 6145 -155 6175
rect -195 6140 -155 6145
rect 5 6245 45 6250
rect 5 6215 10 6245
rect 40 6215 45 6245
rect 5 6175 45 6215
rect 5 6145 10 6175
rect 40 6145 45 6175
rect 5 6140 45 6145
rect 205 6245 245 6250
rect 205 6215 210 6245
rect 240 6215 245 6245
rect 205 6175 245 6215
rect 205 6145 210 6175
rect 240 6145 245 6175
rect 205 6140 245 6145
rect 405 6245 445 6250
rect 405 6215 410 6245
rect 440 6215 445 6245
rect 405 6175 445 6215
rect 405 6145 410 6175
rect 440 6145 445 6175
rect 405 6140 445 6145
rect 605 6245 645 6250
rect 605 6215 610 6245
rect 640 6215 645 6245
rect 605 6175 645 6215
rect 605 6145 610 6175
rect 640 6145 645 6175
rect 605 6140 645 6145
rect 805 6245 845 6250
rect 805 6215 810 6245
rect 840 6215 845 6245
rect 805 6175 845 6215
rect 805 6145 810 6175
rect 840 6145 845 6175
rect 805 6140 845 6145
rect 1005 6245 1045 6250
rect 1005 6215 1010 6245
rect 1040 6215 1045 6245
rect 1005 6175 1045 6215
rect 1005 6145 1010 6175
rect 1040 6145 1045 6175
rect 1005 6140 1045 6145
rect 1205 6245 1245 6250
rect 1205 6215 1210 6245
rect 1240 6215 1245 6245
rect 1205 6175 1245 6215
rect 1205 6145 1210 6175
rect 1240 6145 1245 6175
rect 1205 6140 1245 6145
rect 1405 6245 1445 6250
rect 1405 6215 1410 6245
rect 1440 6215 1445 6245
rect 1405 6175 1445 6215
rect 1405 6145 1410 6175
rect 1440 6145 1445 6175
rect 1405 6140 1445 6145
rect 1605 6245 1645 6250
rect 1605 6215 1610 6245
rect 1640 6215 1645 6245
rect 1605 6175 1645 6215
rect 1605 6145 1610 6175
rect 1640 6145 1645 6175
rect 1605 6140 1645 6145
rect 1805 6245 1845 6250
rect 1805 6215 1810 6245
rect 1840 6215 1845 6245
rect 1805 6175 1845 6215
rect 1805 6145 1810 6175
rect 1840 6145 1845 6175
rect 1805 6140 1845 6145
rect 2005 6245 2045 6250
rect 2005 6215 2010 6245
rect 2040 6215 2045 6245
rect 2005 6175 2045 6215
rect 2005 6145 2010 6175
rect 2040 6145 2045 6175
rect 2005 6140 2045 6145
rect 2205 6245 2245 6250
rect 2205 6215 2210 6245
rect 2240 6215 2245 6245
rect 2205 6175 2245 6215
rect 2205 6145 2210 6175
rect 2240 6145 2245 6175
rect 2205 6140 2245 6145
rect 2405 6245 2445 6250
rect 2405 6215 2410 6245
rect 2440 6215 2445 6245
rect 2405 6175 2445 6215
rect 2405 6145 2410 6175
rect 2440 6145 2445 6175
rect 2405 6140 2445 6145
rect 2605 6245 2645 6250
rect 2605 6215 2610 6245
rect 2640 6215 2645 6245
rect 2605 6175 2645 6215
rect 2605 6145 2610 6175
rect 2640 6145 2645 6175
rect 2605 6140 2645 6145
rect 2805 6245 2845 6250
rect 2805 6215 2810 6245
rect 2840 6215 2845 6245
rect 2805 6175 2845 6215
rect 2805 6145 2810 6175
rect 2840 6145 2845 6175
rect 2805 6140 2845 6145
rect 3005 6245 3045 6250
rect 3005 6215 3010 6245
rect 3040 6215 3045 6245
rect 3005 6175 3045 6215
rect 3005 6145 3010 6175
rect 3040 6145 3045 6175
rect 3005 6140 3045 6145
rect 3205 6245 3245 6250
rect 3205 6215 3210 6245
rect 3240 6215 3245 6245
rect 3205 6175 3245 6215
rect 3205 6145 3210 6175
rect 3240 6145 3245 6175
rect 3205 6140 3245 6145
rect 3405 6245 3445 6250
rect 3405 6215 3410 6245
rect 3440 6215 3445 6245
rect 3405 6175 3445 6215
rect 3405 6145 3410 6175
rect 3440 6145 3445 6175
rect 3405 6140 3445 6145
rect 3605 6245 3645 6250
rect 3605 6215 3610 6245
rect 3640 6215 3645 6245
rect 3605 6175 3645 6215
rect 3605 6145 3610 6175
rect 3640 6145 3645 6175
rect 3605 6140 3645 6145
rect 3805 6245 3845 6250
rect 3805 6215 3810 6245
rect 3840 6215 3845 6245
rect 3805 6175 3845 6215
rect 3805 6145 3810 6175
rect 3840 6145 3845 6175
rect 3805 6140 3845 6145
rect 4005 6245 4045 6250
rect 4005 6215 4010 6245
rect 4040 6215 4045 6245
rect 4005 6175 4045 6215
rect 4005 6145 4010 6175
rect 4040 6145 4045 6175
rect 4005 6140 4045 6145
rect 4205 6245 4245 6250
rect 4205 6215 4210 6245
rect 4240 6215 4245 6245
rect 4205 6175 4245 6215
rect 4205 6145 4210 6175
rect 4240 6145 4245 6175
rect 4205 6140 4245 6145
rect 4405 6245 4445 6250
rect 4405 6215 4410 6245
rect 4440 6215 4445 6245
rect 4405 6175 4445 6215
rect 4405 6145 4410 6175
rect 4440 6145 4445 6175
rect 4405 6140 4445 6145
rect 4605 6245 4645 6250
rect 4605 6215 4610 6245
rect 4640 6215 4645 6245
rect 4605 6175 4645 6215
rect 4605 6145 4610 6175
rect 4640 6145 4645 6175
rect 4605 6140 4645 6145
rect 4805 6245 4845 6250
rect 4805 6215 4810 6245
rect 4840 6215 4845 6245
rect 4805 6175 4845 6215
rect 4805 6145 4810 6175
rect 4840 6145 4845 6175
rect 4805 6140 4845 6145
rect 5005 6245 5045 6250
rect 5005 6215 5010 6245
rect 5040 6215 5045 6245
rect 5005 6175 5045 6215
rect 5005 6145 5010 6175
rect 5040 6145 5045 6175
rect 5005 6140 5045 6145
rect 5205 6245 5245 6250
rect 5205 6215 5210 6245
rect 5240 6215 5245 6245
rect 5205 6175 5245 6215
rect 5205 6145 5210 6175
rect 5240 6145 5245 6175
rect 5205 6140 5245 6145
rect 5405 6245 5445 6250
rect 5405 6215 5410 6245
rect 5440 6215 5445 6245
rect 5405 6175 5445 6215
rect 5405 6145 5410 6175
rect 5440 6145 5445 6175
rect 5405 6140 5445 6145
rect 5605 6245 5645 6250
rect 5605 6215 5610 6245
rect 5640 6215 5645 6245
rect 5605 6175 5645 6215
rect 5605 6145 5610 6175
rect 5640 6145 5645 6175
rect 5605 6140 5645 6145
rect 5805 6245 5845 6250
rect 5805 6215 5810 6245
rect 5840 6215 5845 6245
rect 5805 6175 5845 6215
rect 5805 6145 5810 6175
rect 5840 6145 5845 6175
rect 5805 6140 5845 6145
rect 6005 6245 6045 6250
rect 6005 6215 6010 6245
rect 6040 6215 6045 6245
rect 6005 6175 6045 6215
rect 6005 6145 6010 6175
rect 6040 6145 6045 6175
rect 6005 6140 6045 6145
rect 6205 6245 6245 6250
rect 6205 6215 6210 6245
rect 6240 6215 6245 6245
rect 6205 6175 6245 6215
rect 6205 6145 6210 6175
rect 6240 6145 6245 6175
rect 6205 6140 6245 6145
rect 6405 6245 6445 6250
rect 6405 6215 6410 6245
rect 6440 6215 6445 6245
rect 6405 6175 6445 6215
rect 6405 6145 6410 6175
rect 6440 6145 6445 6175
rect 6405 6140 6445 6145
rect -195 6060 -155 6065
rect -195 6030 -190 6060
rect -160 6030 -155 6060
rect -195 5990 -155 6030
rect -195 5960 -190 5990
rect -160 5960 -155 5990
rect -195 5955 -155 5960
rect 5 6060 45 6065
rect 5 6030 10 6060
rect 40 6030 45 6060
rect 5 5990 45 6030
rect 5 5960 10 5990
rect 40 5960 45 5990
rect 5 5955 45 5960
rect 205 6060 245 6065
rect 205 6030 210 6060
rect 240 6030 245 6060
rect 205 5990 245 6030
rect 205 5960 210 5990
rect 240 5960 245 5990
rect 205 5955 245 5960
rect 405 6060 445 6065
rect 405 6030 410 6060
rect 440 6030 445 6060
rect 405 5990 445 6030
rect 405 5960 410 5990
rect 440 5960 445 5990
rect 405 5955 445 5960
rect 605 6060 645 6065
rect 605 6030 610 6060
rect 640 6030 645 6060
rect 605 5990 645 6030
rect 605 5960 610 5990
rect 640 5960 645 5990
rect 605 5955 645 5960
rect 805 6060 845 6065
rect 805 6030 810 6060
rect 840 6030 845 6060
rect 805 5990 845 6030
rect 805 5960 810 5990
rect 840 5960 845 5990
rect 805 5955 845 5960
rect 1005 6060 1045 6065
rect 1005 6030 1010 6060
rect 1040 6030 1045 6060
rect 1005 5990 1045 6030
rect 1005 5960 1010 5990
rect 1040 5960 1045 5990
rect 1005 5955 1045 5960
rect 1205 6060 1245 6065
rect 1205 6030 1210 6060
rect 1240 6030 1245 6060
rect 1205 5990 1245 6030
rect 1205 5960 1210 5990
rect 1240 5960 1245 5990
rect 1205 5955 1245 5960
rect 1405 6060 1445 6065
rect 1405 6030 1410 6060
rect 1440 6030 1445 6060
rect 1405 5990 1445 6030
rect 1405 5960 1410 5990
rect 1440 5960 1445 5990
rect 1405 5955 1445 5960
rect 1605 6060 1645 6065
rect 1605 6030 1610 6060
rect 1640 6030 1645 6060
rect 1605 5990 1645 6030
rect 1605 5960 1610 5990
rect 1640 5960 1645 5990
rect 1605 5955 1645 5960
rect 1805 6060 1845 6065
rect 1805 6030 1810 6060
rect 1840 6030 1845 6060
rect 1805 5990 1845 6030
rect 1805 5960 1810 5990
rect 1840 5960 1845 5990
rect 1805 5955 1845 5960
rect 2005 6060 2045 6065
rect 2005 6030 2010 6060
rect 2040 6030 2045 6060
rect 2005 5990 2045 6030
rect 2005 5960 2010 5990
rect 2040 5960 2045 5990
rect 2005 5955 2045 5960
rect 2205 6060 2245 6065
rect 2205 6030 2210 6060
rect 2240 6030 2245 6060
rect 2205 5990 2245 6030
rect 2205 5960 2210 5990
rect 2240 5960 2245 5990
rect 2205 5955 2245 5960
rect 2405 6060 2445 6065
rect 2405 6030 2410 6060
rect 2440 6030 2445 6060
rect 2405 5990 2445 6030
rect 2405 5960 2410 5990
rect 2440 5960 2445 5990
rect 2405 5955 2445 5960
rect 2605 6060 2645 6065
rect 2605 6030 2610 6060
rect 2640 6030 2645 6060
rect 2605 5990 2645 6030
rect 2605 5960 2610 5990
rect 2640 5960 2645 5990
rect 2605 5955 2645 5960
rect 2805 6060 2845 6065
rect 2805 6030 2810 6060
rect 2840 6030 2845 6060
rect 2805 5990 2845 6030
rect 2805 5960 2810 5990
rect 2840 5960 2845 5990
rect 2805 5955 2845 5960
rect 3005 6060 3045 6065
rect 3005 6030 3010 6060
rect 3040 6030 3045 6060
rect 3005 5990 3045 6030
rect 3005 5960 3010 5990
rect 3040 5960 3045 5990
rect 3005 5955 3045 5960
rect 3205 6060 3245 6065
rect 3205 6030 3210 6060
rect 3240 6030 3245 6060
rect 3205 5990 3245 6030
rect 3205 5960 3210 5990
rect 3240 5960 3245 5990
rect 3205 5955 3245 5960
rect 3405 6060 3445 6065
rect 3405 6030 3410 6060
rect 3440 6030 3445 6060
rect 3405 5990 3445 6030
rect 3405 5960 3410 5990
rect 3440 5960 3445 5990
rect 3405 5955 3445 5960
rect 3605 6060 3645 6065
rect 3605 6030 3610 6060
rect 3640 6030 3645 6060
rect 3605 5990 3645 6030
rect 3605 5960 3610 5990
rect 3640 5960 3645 5990
rect 3605 5955 3645 5960
rect 3805 6060 3845 6065
rect 3805 6030 3810 6060
rect 3840 6030 3845 6060
rect 3805 5990 3845 6030
rect 3805 5960 3810 5990
rect 3840 5960 3845 5990
rect 3805 5955 3845 5960
rect 4005 6060 4045 6065
rect 4005 6030 4010 6060
rect 4040 6030 4045 6060
rect 4005 5990 4045 6030
rect 4005 5960 4010 5990
rect 4040 5960 4045 5990
rect 4005 5955 4045 5960
rect 4205 6060 4245 6065
rect 4205 6030 4210 6060
rect 4240 6030 4245 6060
rect 4205 5990 4245 6030
rect 4205 5960 4210 5990
rect 4240 5960 4245 5990
rect 4205 5955 4245 5960
rect 4405 6060 4445 6065
rect 4405 6030 4410 6060
rect 4440 6030 4445 6060
rect 4405 5990 4445 6030
rect 4405 5960 4410 5990
rect 4440 5960 4445 5990
rect 4405 5955 4445 5960
rect 4605 6060 4645 6065
rect 4605 6030 4610 6060
rect 4640 6030 4645 6060
rect 4605 5990 4645 6030
rect 4605 5960 4610 5990
rect 4640 5960 4645 5990
rect 4605 5955 4645 5960
rect 4805 6060 4845 6065
rect 4805 6030 4810 6060
rect 4840 6030 4845 6060
rect 4805 5990 4845 6030
rect 4805 5960 4810 5990
rect 4840 5960 4845 5990
rect 4805 5955 4845 5960
rect 5005 6060 5045 6065
rect 5005 6030 5010 6060
rect 5040 6030 5045 6060
rect 5005 5990 5045 6030
rect 5005 5960 5010 5990
rect 5040 5960 5045 5990
rect 5005 5955 5045 5960
rect 5205 6060 5245 6065
rect 5205 6030 5210 6060
rect 5240 6030 5245 6060
rect 5205 5990 5245 6030
rect 5205 5960 5210 5990
rect 5240 5960 5245 5990
rect 5205 5955 5245 5960
rect 5405 6060 5445 6065
rect 5405 6030 5410 6060
rect 5440 6030 5445 6060
rect 5405 5990 5445 6030
rect 5405 5960 5410 5990
rect 5440 5960 5445 5990
rect 5405 5955 5445 5960
rect 5605 6060 5645 6065
rect 5605 6030 5610 6060
rect 5640 6030 5645 6060
rect 5605 5990 5645 6030
rect 5605 5960 5610 5990
rect 5640 5960 5645 5990
rect 5605 5955 5645 5960
rect 5805 6060 5845 6065
rect 5805 6030 5810 6060
rect 5840 6030 5845 6060
rect 5805 5990 5845 6030
rect 5805 5960 5810 5990
rect 5840 5960 5845 5990
rect 5805 5955 5845 5960
rect 6005 6060 6045 6065
rect 6005 6030 6010 6060
rect 6040 6030 6045 6060
rect 6005 5990 6045 6030
rect 6005 5960 6010 5990
rect 6040 5960 6045 5990
rect 6005 5955 6045 5960
rect 6205 6060 6245 6065
rect 6205 6030 6210 6060
rect 6240 6030 6245 6060
rect 6205 5990 6245 6030
rect 6205 5960 6210 5990
rect 6240 5960 6245 5990
rect 6205 5955 6245 5960
rect 6405 6060 6445 6065
rect 6405 6030 6410 6060
rect 6440 6030 6445 6060
rect 6405 5990 6445 6030
rect 6405 5960 6410 5990
rect 6440 5960 6445 5990
rect 6405 5955 6445 5960
rect -195 5875 -155 5880
rect -195 5845 -190 5875
rect -160 5845 -155 5875
rect -195 5805 -155 5845
rect -195 5775 -190 5805
rect -160 5775 -155 5805
rect -195 5770 -155 5775
rect 5 5875 45 5880
rect 5 5845 10 5875
rect 40 5845 45 5875
rect 5 5805 45 5845
rect 5 5775 10 5805
rect 40 5775 45 5805
rect 5 5770 45 5775
rect 205 5875 245 5880
rect 205 5845 210 5875
rect 240 5845 245 5875
rect 205 5805 245 5845
rect 205 5775 210 5805
rect 240 5775 245 5805
rect 205 5770 245 5775
rect 405 5875 445 5880
rect 405 5845 410 5875
rect 440 5845 445 5875
rect 405 5805 445 5845
rect 405 5775 410 5805
rect 440 5775 445 5805
rect 405 5770 445 5775
rect 605 5875 645 5880
rect 605 5845 610 5875
rect 640 5845 645 5875
rect 605 5805 645 5845
rect 605 5775 610 5805
rect 640 5775 645 5805
rect 605 5770 645 5775
rect 805 5875 845 5880
rect 805 5845 810 5875
rect 840 5845 845 5875
rect 805 5805 845 5845
rect 805 5775 810 5805
rect 840 5775 845 5805
rect 805 5770 845 5775
rect 1005 5875 1045 5880
rect 1005 5845 1010 5875
rect 1040 5845 1045 5875
rect 1005 5805 1045 5845
rect 1005 5775 1010 5805
rect 1040 5775 1045 5805
rect 1005 5770 1045 5775
rect 1205 5875 1245 5880
rect 1205 5845 1210 5875
rect 1240 5845 1245 5875
rect 1205 5805 1245 5845
rect 1205 5775 1210 5805
rect 1240 5775 1245 5805
rect 1205 5770 1245 5775
rect 1405 5875 1445 5880
rect 1405 5845 1410 5875
rect 1440 5845 1445 5875
rect 1405 5805 1445 5845
rect 1405 5775 1410 5805
rect 1440 5775 1445 5805
rect 1405 5770 1445 5775
rect 1605 5875 1645 5880
rect 1605 5845 1610 5875
rect 1640 5845 1645 5875
rect 1605 5805 1645 5845
rect 1605 5775 1610 5805
rect 1640 5775 1645 5805
rect 1605 5770 1645 5775
rect 1805 5875 1845 5880
rect 1805 5845 1810 5875
rect 1840 5845 1845 5875
rect 1805 5805 1845 5845
rect 1805 5775 1810 5805
rect 1840 5775 1845 5805
rect 1805 5770 1845 5775
rect 2005 5875 2045 5880
rect 2005 5845 2010 5875
rect 2040 5845 2045 5875
rect 2005 5805 2045 5845
rect 2005 5775 2010 5805
rect 2040 5775 2045 5805
rect 2005 5770 2045 5775
rect 2205 5875 2245 5880
rect 2205 5845 2210 5875
rect 2240 5845 2245 5875
rect 2205 5805 2245 5845
rect 2205 5775 2210 5805
rect 2240 5775 2245 5805
rect 2205 5770 2245 5775
rect 2405 5875 2445 5880
rect 2405 5845 2410 5875
rect 2440 5845 2445 5875
rect 2405 5805 2445 5845
rect 2405 5775 2410 5805
rect 2440 5775 2445 5805
rect 2405 5770 2445 5775
rect 2605 5875 2645 5880
rect 2605 5845 2610 5875
rect 2640 5845 2645 5875
rect 2605 5805 2645 5845
rect 2605 5775 2610 5805
rect 2640 5775 2645 5805
rect 2605 5770 2645 5775
rect 2805 5875 2845 5880
rect 2805 5845 2810 5875
rect 2840 5845 2845 5875
rect 2805 5805 2845 5845
rect 2805 5775 2810 5805
rect 2840 5775 2845 5805
rect 2805 5770 2845 5775
rect 3005 5875 3045 5880
rect 3005 5845 3010 5875
rect 3040 5845 3045 5875
rect 3005 5805 3045 5845
rect 3005 5775 3010 5805
rect 3040 5775 3045 5805
rect 3005 5770 3045 5775
rect 3205 5875 3245 5880
rect 3205 5845 3210 5875
rect 3240 5845 3245 5875
rect 3205 5805 3245 5845
rect 3205 5775 3210 5805
rect 3240 5775 3245 5805
rect 3205 5770 3245 5775
rect 3405 5875 3445 5880
rect 3405 5845 3410 5875
rect 3440 5845 3445 5875
rect 3405 5805 3445 5845
rect 3405 5775 3410 5805
rect 3440 5775 3445 5805
rect 3405 5770 3445 5775
rect 3605 5875 3645 5880
rect 3605 5845 3610 5875
rect 3640 5845 3645 5875
rect 3605 5805 3645 5845
rect 3605 5775 3610 5805
rect 3640 5775 3645 5805
rect 3605 5770 3645 5775
rect 3805 5875 3845 5880
rect 3805 5845 3810 5875
rect 3840 5845 3845 5875
rect 3805 5805 3845 5845
rect 3805 5775 3810 5805
rect 3840 5775 3845 5805
rect 3805 5770 3845 5775
rect 4005 5875 4045 5880
rect 4005 5845 4010 5875
rect 4040 5845 4045 5875
rect 4005 5805 4045 5845
rect 4005 5775 4010 5805
rect 4040 5775 4045 5805
rect 4005 5770 4045 5775
rect 4205 5875 4245 5880
rect 4205 5845 4210 5875
rect 4240 5845 4245 5875
rect 4205 5805 4245 5845
rect 4205 5775 4210 5805
rect 4240 5775 4245 5805
rect 4205 5770 4245 5775
rect 4405 5875 4445 5880
rect 4405 5845 4410 5875
rect 4440 5845 4445 5875
rect 4405 5805 4445 5845
rect 4405 5775 4410 5805
rect 4440 5775 4445 5805
rect 4405 5770 4445 5775
rect 4605 5875 4645 5880
rect 4605 5845 4610 5875
rect 4640 5845 4645 5875
rect 4605 5805 4645 5845
rect 4605 5775 4610 5805
rect 4640 5775 4645 5805
rect 4605 5770 4645 5775
rect 4805 5875 4845 5880
rect 4805 5845 4810 5875
rect 4840 5845 4845 5875
rect 4805 5805 4845 5845
rect 4805 5775 4810 5805
rect 4840 5775 4845 5805
rect 4805 5770 4845 5775
rect 5005 5875 5045 5880
rect 5005 5845 5010 5875
rect 5040 5845 5045 5875
rect 5005 5805 5045 5845
rect 5005 5775 5010 5805
rect 5040 5775 5045 5805
rect 5005 5770 5045 5775
rect 5205 5875 5245 5880
rect 5205 5845 5210 5875
rect 5240 5845 5245 5875
rect 5205 5805 5245 5845
rect 5205 5775 5210 5805
rect 5240 5775 5245 5805
rect 5205 5770 5245 5775
rect 5405 5875 5445 5880
rect 5405 5845 5410 5875
rect 5440 5845 5445 5875
rect 5405 5805 5445 5845
rect 5405 5775 5410 5805
rect 5440 5775 5445 5805
rect 5405 5770 5445 5775
rect 5605 5875 5645 5880
rect 5605 5845 5610 5875
rect 5640 5845 5645 5875
rect 5605 5805 5645 5845
rect 5605 5775 5610 5805
rect 5640 5775 5645 5805
rect 5605 5770 5645 5775
rect 5805 5875 5845 5880
rect 5805 5845 5810 5875
rect 5840 5845 5845 5875
rect 5805 5805 5845 5845
rect 5805 5775 5810 5805
rect 5840 5775 5845 5805
rect 5805 5770 5845 5775
rect 6005 5875 6045 5880
rect 6005 5845 6010 5875
rect 6040 5845 6045 5875
rect 6005 5805 6045 5845
rect 6005 5775 6010 5805
rect 6040 5775 6045 5805
rect 6005 5770 6045 5775
rect 6205 5875 6245 5880
rect 6205 5845 6210 5875
rect 6240 5845 6245 5875
rect 6205 5805 6245 5845
rect 6205 5775 6210 5805
rect 6240 5775 6245 5805
rect 6205 5770 6245 5775
rect 6405 5875 6445 5880
rect 6405 5845 6410 5875
rect 6440 5845 6445 5875
rect 6405 5805 6445 5845
rect 6405 5775 6410 5805
rect 6440 5775 6445 5805
rect 6405 5770 6445 5775
rect -195 5690 -155 5695
rect -195 5660 -190 5690
rect -160 5660 -155 5690
rect -195 5620 -155 5660
rect -195 5590 -190 5620
rect -160 5590 -155 5620
rect -195 5585 -155 5590
rect 5 5690 45 5695
rect 5 5660 10 5690
rect 40 5660 45 5690
rect 5 5620 45 5660
rect 5 5590 10 5620
rect 40 5590 45 5620
rect 5 5585 45 5590
rect 205 5690 245 5695
rect 205 5660 210 5690
rect 240 5660 245 5690
rect 205 5620 245 5660
rect 205 5590 210 5620
rect 240 5590 245 5620
rect 205 5585 245 5590
rect 405 5690 445 5695
rect 405 5660 410 5690
rect 440 5660 445 5690
rect 405 5620 445 5660
rect 405 5590 410 5620
rect 440 5590 445 5620
rect 405 5585 445 5590
rect 605 5690 645 5695
rect 605 5660 610 5690
rect 640 5660 645 5690
rect 605 5620 645 5660
rect 605 5590 610 5620
rect 640 5590 645 5620
rect 605 5585 645 5590
rect 805 5690 845 5695
rect 805 5660 810 5690
rect 840 5660 845 5690
rect 805 5620 845 5660
rect 805 5590 810 5620
rect 840 5590 845 5620
rect 805 5585 845 5590
rect 1005 5690 1045 5695
rect 1005 5660 1010 5690
rect 1040 5660 1045 5690
rect 1005 5620 1045 5660
rect 1005 5590 1010 5620
rect 1040 5590 1045 5620
rect 1005 5585 1045 5590
rect 1205 5690 1245 5695
rect 1205 5660 1210 5690
rect 1240 5660 1245 5690
rect 1205 5620 1245 5660
rect 1205 5590 1210 5620
rect 1240 5590 1245 5620
rect 1205 5585 1245 5590
rect 1405 5690 1445 5695
rect 1405 5660 1410 5690
rect 1440 5660 1445 5690
rect 1405 5620 1445 5660
rect 1405 5590 1410 5620
rect 1440 5590 1445 5620
rect 1405 5585 1445 5590
rect 1605 5690 1645 5695
rect 1605 5660 1610 5690
rect 1640 5660 1645 5690
rect 1605 5620 1645 5660
rect 1605 5590 1610 5620
rect 1640 5590 1645 5620
rect 1605 5585 1645 5590
rect 1805 5690 1845 5695
rect 1805 5660 1810 5690
rect 1840 5660 1845 5690
rect 1805 5620 1845 5660
rect 1805 5590 1810 5620
rect 1840 5590 1845 5620
rect 1805 5585 1845 5590
rect 2005 5690 2045 5695
rect 2005 5660 2010 5690
rect 2040 5660 2045 5690
rect 2005 5620 2045 5660
rect 2005 5590 2010 5620
rect 2040 5590 2045 5620
rect 2005 5585 2045 5590
rect 2205 5690 2245 5695
rect 2205 5660 2210 5690
rect 2240 5660 2245 5690
rect 2205 5620 2245 5660
rect 2205 5590 2210 5620
rect 2240 5590 2245 5620
rect 2205 5585 2245 5590
rect 2405 5690 2445 5695
rect 2405 5660 2410 5690
rect 2440 5660 2445 5690
rect 2405 5620 2445 5660
rect 2405 5590 2410 5620
rect 2440 5590 2445 5620
rect 2405 5585 2445 5590
rect 2605 5690 2645 5695
rect 2605 5660 2610 5690
rect 2640 5660 2645 5690
rect 2605 5620 2645 5660
rect 2605 5590 2610 5620
rect 2640 5590 2645 5620
rect 2605 5585 2645 5590
rect 2805 5690 2845 5695
rect 2805 5660 2810 5690
rect 2840 5660 2845 5690
rect 2805 5620 2845 5660
rect 2805 5590 2810 5620
rect 2840 5590 2845 5620
rect 2805 5585 2845 5590
rect 3005 5690 3045 5695
rect 3005 5660 3010 5690
rect 3040 5660 3045 5690
rect 3005 5620 3045 5660
rect 3005 5590 3010 5620
rect 3040 5590 3045 5620
rect 3005 5585 3045 5590
rect 3205 5690 3245 5695
rect 3205 5660 3210 5690
rect 3240 5660 3245 5690
rect 3205 5620 3245 5660
rect 3205 5590 3210 5620
rect 3240 5590 3245 5620
rect 3205 5585 3245 5590
rect 3405 5690 3445 5695
rect 3405 5660 3410 5690
rect 3440 5660 3445 5690
rect 3405 5620 3445 5660
rect 3405 5590 3410 5620
rect 3440 5590 3445 5620
rect 3405 5585 3445 5590
rect 3605 5690 3645 5695
rect 3605 5660 3610 5690
rect 3640 5660 3645 5690
rect 3605 5620 3645 5660
rect 3605 5590 3610 5620
rect 3640 5590 3645 5620
rect 3605 5585 3645 5590
rect 3805 5690 3845 5695
rect 3805 5660 3810 5690
rect 3840 5660 3845 5690
rect 3805 5620 3845 5660
rect 3805 5590 3810 5620
rect 3840 5590 3845 5620
rect 3805 5585 3845 5590
rect 4005 5690 4045 5695
rect 4005 5660 4010 5690
rect 4040 5660 4045 5690
rect 4005 5620 4045 5660
rect 4005 5590 4010 5620
rect 4040 5590 4045 5620
rect 4005 5585 4045 5590
rect 4205 5690 4245 5695
rect 4205 5660 4210 5690
rect 4240 5660 4245 5690
rect 4205 5620 4245 5660
rect 4205 5590 4210 5620
rect 4240 5590 4245 5620
rect 4205 5585 4245 5590
rect 4405 5690 4445 5695
rect 4405 5660 4410 5690
rect 4440 5660 4445 5690
rect 4405 5620 4445 5660
rect 4405 5590 4410 5620
rect 4440 5590 4445 5620
rect 4405 5585 4445 5590
rect 4605 5690 4645 5695
rect 4605 5660 4610 5690
rect 4640 5660 4645 5690
rect 4605 5620 4645 5660
rect 4605 5590 4610 5620
rect 4640 5590 4645 5620
rect 4605 5585 4645 5590
rect 4805 5690 4845 5695
rect 4805 5660 4810 5690
rect 4840 5660 4845 5690
rect 4805 5620 4845 5660
rect 4805 5590 4810 5620
rect 4840 5590 4845 5620
rect 4805 5585 4845 5590
rect 5005 5690 5045 5695
rect 5005 5660 5010 5690
rect 5040 5660 5045 5690
rect 5005 5620 5045 5660
rect 5005 5590 5010 5620
rect 5040 5590 5045 5620
rect 5005 5585 5045 5590
rect 5205 5690 5245 5695
rect 5205 5660 5210 5690
rect 5240 5660 5245 5690
rect 5205 5620 5245 5660
rect 5205 5590 5210 5620
rect 5240 5590 5245 5620
rect 5205 5585 5245 5590
rect 5405 5690 5445 5695
rect 5405 5660 5410 5690
rect 5440 5660 5445 5690
rect 5405 5620 5445 5660
rect 5405 5590 5410 5620
rect 5440 5590 5445 5620
rect 5405 5585 5445 5590
rect 5605 5690 5645 5695
rect 5605 5660 5610 5690
rect 5640 5660 5645 5690
rect 5605 5620 5645 5660
rect 5605 5590 5610 5620
rect 5640 5590 5645 5620
rect 5605 5585 5645 5590
rect 5805 5690 5845 5695
rect 5805 5660 5810 5690
rect 5840 5660 5845 5690
rect 5805 5620 5845 5660
rect 5805 5590 5810 5620
rect 5840 5590 5845 5620
rect 5805 5585 5845 5590
rect 6005 5690 6045 5695
rect 6005 5660 6010 5690
rect 6040 5660 6045 5690
rect 6005 5620 6045 5660
rect 6005 5590 6010 5620
rect 6040 5590 6045 5620
rect 6005 5585 6045 5590
rect 6205 5690 6245 5695
rect 6205 5660 6210 5690
rect 6240 5660 6245 5690
rect 6205 5620 6245 5660
rect 6205 5590 6210 5620
rect 6240 5590 6245 5620
rect 6205 5585 6245 5590
rect 6405 5690 6445 5695
rect 6405 5660 6410 5690
rect 6440 5660 6445 5690
rect 6405 5620 6445 5660
rect 6405 5590 6410 5620
rect 6440 5590 6445 5620
rect 6405 5585 6445 5590
rect -195 5505 -155 5510
rect -195 5475 -190 5505
rect -160 5475 -155 5505
rect -195 5435 -155 5475
rect -195 5405 -190 5435
rect -160 5405 -155 5435
rect -195 5400 -155 5405
rect 5 5505 45 5510
rect 5 5475 10 5505
rect 40 5475 45 5505
rect 5 5435 45 5475
rect 5 5405 10 5435
rect 40 5405 45 5435
rect 5 5400 45 5405
rect 205 5505 245 5510
rect 205 5475 210 5505
rect 240 5475 245 5505
rect 205 5435 245 5475
rect 205 5405 210 5435
rect 240 5405 245 5435
rect 205 5400 245 5405
rect 405 5505 445 5510
rect 405 5475 410 5505
rect 440 5475 445 5505
rect 405 5435 445 5475
rect 405 5405 410 5435
rect 440 5405 445 5435
rect 405 5400 445 5405
rect 605 5505 645 5510
rect 605 5475 610 5505
rect 640 5475 645 5505
rect 605 5435 645 5475
rect 605 5405 610 5435
rect 640 5405 645 5435
rect 605 5400 645 5405
rect 805 5505 845 5510
rect 805 5475 810 5505
rect 840 5475 845 5505
rect 805 5435 845 5475
rect 805 5405 810 5435
rect 840 5405 845 5435
rect 805 5400 845 5405
rect 1005 5505 1045 5510
rect 1005 5475 1010 5505
rect 1040 5475 1045 5505
rect 1005 5435 1045 5475
rect 1005 5405 1010 5435
rect 1040 5405 1045 5435
rect 1005 5400 1045 5405
rect 1205 5505 1245 5510
rect 1205 5475 1210 5505
rect 1240 5475 1245 5505
rect 1205 5435 1245 5475
rect 1205 5405 1210 5435
rect 1240 5405 1245 5435
rect 1205 5400 1245 5405
rect 1405 5505 1445 5510
rect 1405 5475 1410 5505
rect 1440 5475 1445 5505
rect 1405 5435 1445 5475
rect 1405 5405 1410 5435
rect 1440 5405 1445 5435
rect 1405 5400 1445 5405
rect 1605 5505 1645 5510
rect 1605 5475 1610 5505
rect 1640 5475 1645 5505
rect 1605 5435 1645 5475
rect 1605 5405 1610 5435
rect 1640 5405 1645 5435
rect 1605 5400 1645 5405
rect 1805 5505 1845 5510
rect 1805 5475 1810 5505
rect 1840 5475 1845 5505
rect 1805 5435 1845 5475
rect 1805 5405 1810 5435
rect 1840 5405 1845 5435
rect 1805 5400 1845 5405
rect 2005 5505 2045 5510
rect 2005 5475 2010 5505
rect 2040 5475 2045 5505
rect 2005 5435 2045 5475
rect 2005 5405 2010 5435
rect 2040 5405 2045 5435
rect 2005 5400 2045 5405
rect 2205 5505 2245 5510
rect 2205 5475 2210 5505
rect 2240 5475 2245 5505
rect 2205 5435 2245 5475
rect 2205 5405 2210 5435
rect 2240 5405 2245 5435
rect 2205 5400 2245 5405
rect 2405 5505 2445 5510
rect 2405 5475 2410 5505
rect 2440 5475 2445 5505
rect 2405 5435 2445 5475
rect 2405 5405 2410 5435
rect 2440 5405 2445 5435
rect 2405 5400 2445 5405
rect 2605 5505 2645 5510
rect 2605 5475 2610 5505
rect 2640 5475 2645 5505
rect 2605 5435 2645 5475
rect 2605 5405 2610 5435
rect 2640 5405 2645 5435
rect 2605 5400 2645 5405
rect 2805 5505 2845 5510
rect 2805 5475 2810 5505
rect 2840 5475 2845 5505
rect 2805 5435 2845 5475
rect 2805 5405 2810 5435
rect 2840 5405 2845 5435
rect 2805 5400 2845 5405
rect 3005 5505 3045 5510
rect 3005 5475 3010 5505
rect 3040 5475 3045 5505
rect 3005 5435 3045 5475
rect 3005 5405 3010 5435
rect 3040 5405 3045 5435
rect 3005 5400 3045 5405
rect 3205 5505 3245 5510
rect 3205 5475 3210 5505
rect 3240 5475 3245 5505
rect 3205 5435 3245 5475
rect 3205 5405 3210 5435
rect 3240 5405 3245 5435
rect 3205 5400 3245 5405
rect 3405 5505 3445 5510
rect 3405 5475 3410 5505
rect 3440 5475 3445 5505
rect 3405 5435 3445 5475
rect 3405 5405 3410 5435
rect 3440 5405 3445 5435
rect 3405 5400 3445 5405
rect 3605 5505 3645 5510
rect 3605 5475 3610 5505
rect 3640 5475 3645 5505
rect 3605 5435 3645 5475
rect 3605 5405 3610 5435
rect 3640 5405 3645 5435
rect 3605 5400 3645 5405
rect 3805 5505 3845 5510
rect 3805 5475 3810 5505
rect 3840 5475 3845 5505
rect 3805 5435 3845 5475
rect 3805 5405 3810 5435
rect 3840 5405 3845 5435
rect 3805 5400 3845 5405
rect 4005 5505 4045 5510
rect 4005 5475 4010 5505
rect 4040 5475 4045 5505
rect 4005 5435 4045 5475
rect 4005 5405 4010 5435
rect 4040 5405 4045 5435
rect 4005 5400 4045 5405
rect 4205 5505 4245 5510
rect 4205 5475 4210 5505
rect 4240 5475 4245 5505
rect 4205 5435 4245 5475
rect 4205 5405 4210 5435
rect 4240 5405 4245 5435
rect 4205 5400 4245 5405
rect 4405 5505 4445 5510
rect 4405 5475 4410 5505
rect 4440 5475 4445 5505
rect 4405 5435 4445 5475
rect 4405 5405 4410 5435
rect 4440 5405 4445 5435
rect 4405 5400 4445 5405
rect 4605 5505 4645 5510
rect 4605 5475 4610 5505
rect 4640 5475 4645 5505
rect 4605 5435 4645 5475
rect 4605 5405 4610 5435
rect 4640 5405 4645 5435
rect 4605 5400 4645 5405
rect 4805 5505 4845 5510
rect 4805 5475 4810 5505
rect 4840 5475 4845 5505
rect 4805 5435 4845 5475
rect 4805 5405 4810 5435
rect 4840 5405 4845 5435
rect 4805 5400 4845 5405
rect 5005 5505 5045 5510
rect 5005 5475 5010 5505
rect 5040 5475 5045 5505
rect 5005 5435 5045 5475
rect 5005 5405 5010 5435
rect 5040 5405 5045 5435
rect 5005 5400 5045 5405
rect 5205 5505 5245 5510
rect 5205 5475 5210 5505
rect 5240 5475 5245 5505
rect 5205 5435 5245 5475
rect 5205 5405 5210 5435
rect 5240 5405 5245 5435
rect 5205 5400 5245 5405
rect 5405 5505 5445 5510
rect 5405 5475 5410 5505
rect 5440 5475 5445 5505
rect 5405 5435 5445 5475
rect 5405 5405 5410 5435
rect 5440 5405 5445 5435
rect 5405 5400 5445 5405
rect 5605 5505 5645 5510
rect 5605 5475 5610 5505
rect 5640 5475 5645 5505
rect 5605 5435 5645 5475
rect 5605 5405 5610 5435
rect 5640 5405 5645 5435
rect 5605 5400 5645 5405
rect 5805 5505 5845 5510
rect 5805 5475 5810 5505
rect 5840 5475 5845 5505
rect 5805 5435 5845 5475
rect 5805 5405 5810 5435
rect 5840 5405 5845 5435
rect 5805 5400 5845 5405
rect 6005 5505 6045 5510
rect 6005 5475 6010 5505
rect 6040 5475 6045 5505
rect 6005 5435 6045 5475
rect 6005 5405 6010 5435
rect 6040 5405 6045 5435
rect 6005 5400 6045 5405
rect 6205 5505 6245 5510
rect 6205 5475 6210 5505
rect 6240 5475 6245 5505
rect 6205 5435 6245 5475
rect 6205 5405 6210 5435
rect 6240 5405 6245 5435
rect 6205 5400 6245 5405
rect 6405 5505 6445 5510
rect 6405 5475 6410 5505
rect 6440 5475 6445 5505
rect 6405 5435 6445 5475
rect 6405 5405 6410 5435
rect 6440 5405 6445 5435
rect 6405 5400 6445 5405
rect -195 5320 -155 5325
rect -195 5290 -190 5320
rect -160 5290 -155 5320
rect -195 5250 -155 5290
rect -195 5220 -190 5250
rect -160 5220 -155 5250
rect -195 5215 -155 5220
rect 5 5320 45 5325
rect 5 5290 10 5320
rect 40 5290 45 5320
rect 5 5250 45 5290
rect 5 5220 10 5250
rect 40 5220 45 5250
rect 5 5215 45 5220
rect 205 5320 245 5325
rect 205 5290 210 5320
rect 240 5290 245 5320
rect 205 5250 245 5290
rect 205 5220 210 5250
rect 240 5220 245 5250
rect 205 5215 245 5220
rect 405 5320 445 5325
rect 405 5290 410 5320
rect 440 5290 445 5320
rect 405 5250 445 5290
rect 405 5220 410 5250
rect 440 5220 445 5250
rect 405 5215 445 5220
rect 605 5320 645 5325
rect 605 5290 610 5320
rect 640 5290 645 5320
rect 605 5250 645 5290
rect 605 5220 610 5250
rect 640 5220 645 5250
rect 605 5215 645 5220
rect 805 5320 845 5325
rect 805 5290 810 5320
rect 840 5290 845 5320
rect 805 5250 845 5290
rect 805 5220 810 5250
rect 840 5220 845 5250
rect 805 5215 845 5220
rect 1005 5320 1045 5325
rect 1005 5290 1010 5320
rect 1040 5290 1045 5320
rect 1005 5250 1045 5290
rect 1005 5220 1010 5250
rect 1040 5220 1045 5250
rect 1005 5215 1045 5220
rect 1205 5320 1245 5325
rect 1205 5290 1210 5320
rect 1240 5290 1245 5320
rect 1205 5250 1245 5290
rect 1205 5220 1210 5250
rect 1240 5220 1245 5250
rect 1205 5215 1245 5220
rect 1405 5320 1445 5325
rect 1405 5290 1410 5320
rect 1440 5290 1445 5320
rect 1405 5250 1445 5290
rect 1405 5220 1410 5250
rect 1440 5220 1445 5250
rect 1405 5215 1445 5220
rect 1605 5320 1645 5325
rect 1605 5290 1610 5320
rect 1640 5290 1645 5320
rect 1605 5250 1645 5290
rect 1605 5220 1610 5250
rect 1640 5220 1645 5250
rect 1605 5215 1645 5220
rect 1805 5320 1845 5325
rect 1805 5290 1810 5320
rect 1840 5290 1845 5320
rect 1805 5250 1845 5290
rect 1805 5220 1810 5250
rect 1840 5220 1845 5250
rect 1805 5215 1845 5220
rect 2005 5320 2045 5325
rect 2005 5290 2010 5320
rect 2040 5290 2045 5320
rect 2005 5250 2045 5290
rect 2005 5220 2010 5250
rect 2040 5220 2045 5250
rect 2005 5215 2045 5220
rect 2205 5320 2245 5325
rect 2205 5290 2210 5320
rect 2240 5290 2245 5320
rect 2205 5250 2245 5290
rect 2205 5220 2210 5250
rect 2240 5220 2245 5250
rect 2205 5215 2245 5220
rect 2405 5320 2445 5325
rect 2405 5290 2410 5320
rect 2440 5290 2445 5320
rect 2405 5250 2445 5290
rect 2405 5220 2410 5250
rect 2440 5220 2445 5250
rect 2405 5215 2445 5220
rect 2605 5320 2645 5325
rect 2605 5290 2610 5320
rect 2640 5290 2645 5320
rect 2605 5250 2645 5290
rect 2605 5220 2610 5250
rect 2640 5220 2645 5250
rect 2605 5215 2645 5220
rect 2805 5320 2845 5325
rect 2805 5290 2810 5320
rect 2840 5290 2845 5320
rect 2805 5250 2845 5290
rect 2805 5220 2810 5250
rect 2840 5220 2845 5250
rect 2805 5215 2845 5220
rect 3005 5320 3045 5325
rect 3005 5290 3010 5320
rect 3040 5290 3045 5320
rect 3005 5250 3045 5290
rect 3005 5220 3010 5250
rect 3040 5220 3045 5250
rect 3005 5215 3045 5220
rect 3205 5320 3245 5325
rect 3205 5290 3210 5320
rect 3240 5290 3245 5320
rect 3205 5250 3245 5290
rect 3205 5220 3210 5250
rect 3240 5220 3245 5250
rect 3205 5215 3245 5220
rect 3405 5320 3445 5325
rect 3405 5290 3410 5320
rect 3440 5290 3445 5320
rect 3405 5250 3445 5290
rect 3405 5220 3410 5250
rect 3440 5220 3445 5250
rect 3405 5215 3445 5220
rect 3605 5320 3645 5325
rect 3605 5290 3610 5320
rect 3640 5290 3645 5320
rect 3605 5250 3645 5290
rect 3605 5220 3610 5250
rect 3640 5220 3645 5250
rect 3605 5215 3645 5220
rect 3805 5320 3845 5325
rect 3805 5290 3810 5320
rect 3840 5290 3845 5320
rect 3805 5250 3845 5290
rect 3805 5220 3810 5250
rect 3840 5220 3845 5250
rect 3805 5215 3845 5220
rect 4005 5320 4045 5325
rect 4005 5290 4010 5320
rect 4040 5290 4045 5320
rect 4005 5250 4045 5290
rect 4005 5220 4010 5250
rect 4040 5220 4045 5250
rect 4005 5215 4045 5220
rect 4205 5320 4245 5325
rect 4205 5290 4210 5320
rect 4240 5290 4245 5320
rect 4205 5250 4245 5290
rect 4205 5220 4210 5250
rect 4240 5220 4245 5250
rect 4205 5215 4245 5220
rect 4405 5320 4445 5325
rect 4405 5290 4410 5320
rect 4440 5290 4445 5320
rect 4405 5250 4445 5290
rect 4405 5220 4410 5250
rect 4440 5220 4445 5250
rect 4405 5215 4445 5220
rect 4605 5320 4645 5325
rect 4605 5290 4610 5320
rect 4640 5290 4645 5320
rect 4605 5250 4645 5290
rect 4605 5220 4610 5250
rect 4640 5220 4645 5250
rect 4605 5215 4645 5220
rect 4805 5320 4845 5325
rect 4805 5290 4810 5320
rect 4840 5290 4845 5320
rect 4805 5250 4845 5290
rect 4805 5220 4810 5250
rect 4840 5220 4845 5250
rect 4805 5215 4845 5220
rect 5005 5320 5045 5325
rect 5005 5290 5010 5320
rect 5040 5290 5045 5320
rect 5005 5250 5045 5290
rect 5005 5220 5010 5250
rect 5040 5220 5045 5250
rect 5005 5215 5045 5220
rect 5205 5320 5245 5325
rect 5205 5290 5210 5320
rect 5240 5290 5245 5320
rect 5205 5250 5245 5290
rect 5205 5220 5210 5250
rect 5240 5220 5245 5250
rect 5205 5215 5245 5220
rect 5405 5320 5445 5325
rect 5405 5290 5410 5320
rect 5440 5290 5445 5320
rect 5405 5250 5445 5290
rect 5405 5220 5410 5250
rect 5440 5220 5445 5250
rect 5405 5215 5445 5220
rect 5605 5320 5645 5325
rect 5605 5290 5610 5320
rect 5640 5290 5645 5320
rect 5605 5250 5645 5290
rect 5605 5220 5610 5250
rect 5640 5220 5645 5250
rect 5605 5215 5645 5220
rect 5805 5320 5845 5325
rect 5805 5290 5810 5320
rect 5840 5290 5845 5320
rect 5805 5250 5845 5290
rect 5805 5220 5810 5250
rect 5840 5220 5845 5250
rect 5805 5215 5845 5220
rect 6005 5320 6045 5325
rect 6005 5290 6010 5320
rect 6040 5290 6045 5320
rect 6005 5250 6045 5290
rect 6005 5220 6010 5250
rect 6040 5220 6045 5250
rect 6005 5215 6045 5220
rect 6205 5320 6245 5325
rect 6205 5290 6210 5320
rect 6240 5290 6245 5320
rect 6205 5250 6245 5290
rect 6205 5220 6210 5250
rect 6240 5220 6245 5250
rect 6205 5215 6245 5220
rect 6405 5320 6445 5325
rect 6405 5290 6410 5320
rect 6440 5290 6445 5320
rect 6405 5250 6445 5290
rect 6405 5220 6410 5250
rect 6440 5220 6445 5250
rect 6405 5215 6445 5220
rect -195 5135 -155 5140
rect -195 5105 -190 5135
rect -160 5105 -155 5135
rect -195 5065 -155 5105
rect -195 5035 -190 5065
rect -160 5035 -155 5065
rect -195 5030 -155 5035
rect 5 5135 45 5140
rect 5 5105 10 5135
rect 40 5105 45 5135
rect 5 5065 45 5105
rect 5 5035 10 5065
rect 40 5035 45 5065
rect 5 5030 45 5035
rect 205 5135 245 5140
rect 205 5105 210 5135
rect 240 5105 245 5135
rect 205 5065 245 5105
rect 205 5035 210 5065
rect 240 5035 245 5065
rect 205 5030 245 5035
rect 405 5135 445 5140
rect 405 5105 410 5135
rect 440 5105 445 5135
rect 405 5065 445 5105
rect 405 5035 410 5065
rect 440 5035 445 5065
rect 405 5030 445 5035
rect 605 5135 645 5140
rect 605 5105 610 5135
rect 640 5105 645 5135
rect 605 5065 645 5105
rect 605 5035 610 5065
rect 640 5035 645 5065
rect 605 5030 645 5035
rect 805 5135 845 5140
rect 805 5105 810 5135
rect 840 5105 845 5135
rect 805 5065 845 5105
rect 805 5035 810 5065
rect 840 5035 845 5065
rect 805 5030 845 5035
rect 1005 5135 1045 5140
rect 1005 5105 1010 5135
rect 1040 5105 1045 5135
rect 1005 5065 1045 5105
rect 1005 5035 1010 5065
rect 1040 5035 1045 5065
rect 1005 5030 1045 5035
rect 1205 5135 1245 5140
rect 1205 5105 1210 5135
rect 1240 5105 1245 5135
rect 1205 5065 1245 5105
rect 1205 5035 1210 5065
rect 1240 5035 1245 5065
rect 1205 5030 1245 5035
rect 1405 5135 1445 5140
rect 1405 5105 1410 5135
rect 1440 5105 1445 5135
rect 1405 5065 1445 5105
rect 1405 5035 1410 5065
rect 1440 5035 1445 5065
rect 1405 5030 1445 5035
rect 1605 5135 1645 5140
rect 1605 5105 1610 5135
rect 1640 5105 1645 5135
rect 1605 5065 1645 5105
rect 1605 5035 1610 5065
rect 1640 5035 1645 5065
rect 1605 5030 1645 5035
rect 1805 5135 1845 5140
rect 1805 5105 1810 5135
rect 1840 5105 1845 5135
rect 1805 5065 1845 5105
rect 1805 5035 1810 5065
rect 1840 5035 1845 5065
rect 1805 5030 1845 5035
rect 2005 5135 2045 5140
rect 2005 5105 2010 5135
rect 2040 5105 2045 5135
rect 2005 5065 2045 5105
rect 2005 5035 2010 5065
rect 2040 5035 2045 5065
rect 2005 5030 2045 5035
rect 2205 5135 2245 5140
rect 2205 5105 2210 5135
rect 2240 5105 2245 5135
rect 2205 5065 2245 5105
rect 2205 5035 2210 5065
rect 2240 5035 2245 5065
rect 2205 5030 2245 5035
rect 2405 5135 2445 5140
rect 2405 5105 2410 5135
rect 2440 5105 2445 5135
rect 2405 5065 2445 5105
rect 2405 5035 2410 5065
rect 2440 5035 2445 5065
rect 2405 5030 2445 5035
rect 2605 5135 2645 5140
rect 2605 5105 2610 5135
rect 2640 5105 2645 5135
rect 2605 5065 2645 5105
rect 2605 5035 2610 5065
rect 2640 5035 2645 5065
rect 2605 5030 2645 5035
rect 2805 5135 2845 5140
rect 2805 5105 2810 5135
rect 2840 5105 2845 5135
rect 2805 5065 2845 5105
rect 2805 5035 2810 5065
rect 2840 5035 2845 5065
rect 2805 5030 2845 5035
rect 3005 5135 3045 5140
rect 3005 5105 3010 5135
rect 3040 5105 3045 5135
rect 3005 5065 3045 5105
rect 3005 5035 3010 5065
rect 3040 5035 3045 5065
rect 3005 5030 3045 5035
rect 3205 5135 3245 5140
rect 3205 5105 3210 5135
rect 3240 5105 3245 5135
rect 3205 5065 3245 5105
rect 3205 5035 3210 5065
rect 3240 5035 3245 5065
rect 3205 5030 3245 5035
rect 3405 5135 3445 5140
rect 3405 5105 3410 5135
rect 3440 5105 3445 5135
rect 3405 5065 3445 5105
rect 3405 5035 3410 5065
rect 3440 5035 3445 5065
rect 3405 5030 3445 5035
rect 3605 5135 3645 5140
rect 3605 5105 3610 5135
rect 3640 5105 3645 5135
rect 3605 5065 3645 5105
rect 3605 5035 3610 5065
rect 3640 5035 3645 5065
rect 3605 5030 3645 5035
rect 3805 5135 3845 5140
rect 3805 5105 3810 5135
rect 3840 5105 3845 5135
rect 3805 5065 3845 5105
rect 3805 5035 3810 5065
rect 3840 5035 3845 5065
rect 3805 5030 3845 5035
rect 4005 5135 4045 5140
rect 4005 5105 4010 5135
rect 4040 5105 4045 5135
rect 4005 5065 4045 5105
rect 4005 5035 4010 5065
rect 4040 5035 4045 5065
rect 4005 5030 4045 5035
rect 4205 5135 4245 5140
rect 4205 5105 4210 5135
rect 4240 5105 4245 5135
rect 4205 5065 4245 5105
rect 4205 5035 4210 5065
rect 4240 5035 4245 5065
rect 4205 5030 4245 5035
rect 4405 5135 4445 5140
rect 4405 5105 4410 5135
rect 4440 5105 4445 5135
rect 4405 5065 4445 5105
rect 4405 5035 4410 5065
rect 4440 5035 4445 5065
rect 4405 5030 4445 5035
rect 4605 5135 4645 5140
rect 4605 5105 4610 5135
rect 4640 5105 4645 5135
rect 4605 5065 4645 5105
rect 4605 5035 4610 5065
rect 4640 5035 4645 5065
rect 4605 5030 4645 5035
rect 4805 5135 4845 5140
rect 4805 5105 4810 5135
rect 4840 5105 4845 5135
rect 4805 5065 4845 5105
rect 4805 5035 4810 5065
rect 4840 5035 4845 5065
rect 4805 5030 4845 5035
rect 5005 5135 5045 5140
rect 5005 5105 5010 5135
rect 5040 5105 5045 5135
rect 5005 5065 5045 5105
rect 5005 5035 5010 5065
rect 5040 5035 5045 5065
rect 5005 5030 5045 5035
rect 5205 5135 5245 5140
rect 5205 5105 5210 5135
rect 5240 5105 5245 5135
rect 5205 5065 5245 5105
rect 5205 5035 5210 5065
rect 5240 5035 5245 5065
rect 5205 5030 5245 5035
rect 5405 5135 5445 5140
rect 5405 5105 5410 5135
rect 5440 5105 5445 5135
rect 5405 5065 5445 5105
rect 5405 5035 5410 5065
rect 5440 5035 5445 5065
rect 5405 5030 5445 5035
rect 5605 5135 5645 5140
rect 5605 5105 5610 5135
rect 5640 5105 5645 5135
rect 5605 5065 5645 5105
rect 5605 5035 5610 5065
rect 5640 5035 5645 5065
rect 5605 5030 5645 5035
rect 5805 5135 5845 5140
rect 5805 5105 5810 5135
rect 5840 5105 5845 5135
rect 5805 5065 5845 5105
rect 5805 5035 5810 5065
rect 5840 5035 5845 5065
rect 5805 5030 5845 5035
rect 6005 5135 6045 5140
rect 6005 5105 6010 5135
rect 6040 5105 6045 5135
rect 6005 5065 6045 5105
rect 6005 5035 6010 5065
rect 6040 5035 6045 5065
rect 6005 5030 6045 5035
rect 6205 5135 6245 5140
rect 6205 5105 6210 5135
rect 6240 5105 6245 5135
rect 6205 5065 6245 5105
rect 6205 5035 6210 5065
rect 6240 5035 6245 5065
rect 6205 5030 6245 5035
rect 6405 5135 6445 5140
rect 6405 5105 6410 5135
rect 6440 5105 6445 5135
rect 6405 5065 6445 5105
rect 6405 5035 6410 5065
rect 6440 5035 6445 5065
rect 6405 5030 6445 5035
rect -195 4950 -155 4955
rect -195 4920 -190 4950
rect -160 4920 -155 4950
rect -195 4880 -155 4920
rect -195 4850 -190 4880
rect -160 4850 -155 4880
rect -195 4845 -155 4850
rect 5 4950 45 4955
rect 5 4920 10 4950
rect 40 4920 45 4950
rect 5 4880 45 4920
rect 5 4850 10 4880
rect 40 4850 45 4880
rect 5 4845 45 4850
rect 205 4950 245 4955
rect 205 4920 210 4950
rect 240 4920 245 4950
rect 205 4880 245 4920
rect 205 4850 210 4880
rect 240 4850 245 4880
rect 205 4845 245 4850
rect 405 4950 445 4955
rect 405 4920 410 4950
rect 440 4920 445 4950
rect 405 4880 445 4920
rect 405 4850 410 4880
rect 440 4850 445 4880
rect 405 4845 445 4850
rect 605 4950 645 4955
rect 605 4920 610 4950
rect 640 4920 645 4950
rect 605 4880 645 4920
rect 605 4850 610 4880
rect 640 4850 645 4880
rect 605 4845 645 4850
rect 805 4950 845 4955
rect 805 4920 810 4950
rect 840 4920 845 4950
rect 805 4880 845 4920
rect 805 4850 810 4880
rect 840 4850 845 4880
rect 805 4845 845 4850
rect 1005 4950 1045 4955
rect 1005 4920 1010 4950
rect 1040 4920 1045 4950
rect 1005 4880 1045 4920
rect 1005 4850 1010 4880
rect 1040 4850 1045 4880
rect 1005 4845 1045 4850
rect 1205 4950 1245 4955
rect 1205 4920 1210 4950
rect 1240 4920 1245 4950
rect 1205 4880 1245 4920
rect 1205 4850 1210 4880
rect 1240 4850 1245 4880
rect 1205 4845 1245 4850
rect 1405 4950 1445 4955
rect 1405 4920 1410 4950
rect 1440 4920 1445 4950
rect 1405 4880 1445 4920
rect 1405 4850 1410 4880
rect 1440 4850 1445 4880
rect 1405 4845 1445 4850
rect 1605 4950 1645 4955
rect 1605 4920 1610 4950
rect 1640 4920 1645 4950
rect 1605 4880 1645 4920
rect 1605 4850 1610 4880
rect 1640 4850 1645 4880
rect 1605 4845 1645 4850
rect 1805 4950 1845 4955
rect 1805 4920 1810 4950
rect 1840 4920 1845 4950
rect 1805 4880 1845 4920
rect 1805 4850 1810 4880
rect 1840 4850 1845 4880
rect 1805 4845 1845 4850
rect 2005 4950 2045 4955
rect 2005 4920 2010 4950
rect 2040 4920 2045 4950
rect 2005 4880 2045 4920
rect 2005 4850 2010 4880
rect 2040 4850 2045 4880
rect 2005 4845 2045 4850
rect 2205 4950 2245 4955
rect 2205 4920 2210 4950
rect 2240 4920 2245 4950
rect 2205 4880 2245 4920
rect 2205 4850 2210 4880
rect 2240 4850 2245 4880
rect 2205 4845 2245 4850
rect 2405 4950 2445 4955
rect 2405 4920 2410 4950
rect 2440 4920 2445 4950
rect 2405 4880 2445 4920
rect 2405 4850 2410 4880
rect 2440 4850 2445 4880
rect 2405 4845 2445 4850
rect 2605 4950 2645 4955
rect 2605 4920 2610 4950
rect 2640 4920 2645 4950
rect 2605 4880 2645 4920
rect 2605 4850 2610 4880
rect 2640 4850 2645 4880
rect 2605 4845 2645 4850
rect 2805 4950 2845 4955
rect 2805 4920 2810 4950
rect 2840 4920 2845 4950
rect 2805 4880 2845 4920
rect 2805 4850 2810 4880
rect 2840 4850 2845 4880
rect 2805 4845 2845 4850
rect 3005 4950 3045 4955
rect 3005 4920 3010 4950
rect 3040 4920 3045 4950
rect 3005 4880 3045 4920
rect 3005 4850 3010 4880
rect 3040 4850 3045 4880
rect 3005 4845 3045 4850
rect 3205 4950 3245 4955
rect 3205 4920 3210 4950
rect 3240 4920 3245 4950
rect 3205 4880 3245 4920
rect 3205 4850 3210 4880
rect 3240 4850 3245 4880
rect 3205 4845 3245 4850
rect 3405 4950 3445 4955
rect 3405 4920 3410 4950
rect 3440 4920 3445 4950
rect 3405 4880 3445 4920
rect 3405 4850 3410 4880
rect 3440 4850 3445 4880
rect 3405 4845 3445 4850
rect 3605 4950 3645 4955
rect 3605 4920 3610 4950
rect 3640 4920 3645 4950
rect 3605 4880 3645 4920
rect 3605 4850 3610 4880
rect 3640 4850 3645 4880
rect 3605 4845 3645 4850
rect 3805 4950 3845 4955
rect 3805 4920 3810 4950
rect 3840 4920 3845 4950
rect 3805 4880 3845 4920
rect 3805 4850 3810 4880
rect 3840 4850 3845 4880
rect 3805 4845 3845 4850
rect 4005 4950 4045 4955
rect 4005 4920 4010 4950
rect 4040 4920 4045 4950
rect 4005 4880 4045 4920
rect 4005 4850 4010 4880
rect 4040 4850 4045 4880
rect 4005 4845 4045 4850
rect 4205 4950 4245 4955
rect 4205 4920 4210 4950
rect 4240 4920 4245 4950
rect 4205 4880 4245 4920
rect 4205 4850 4210 4880
rect 4240 4850 4245 4880
rect 4205 4845 4245 4850
rect 4405 4950 4445 4955
rect 4405 4920 4410 4950
rect 4440 4920 4445 4950
rect 4405 4880 4445 4920
rect 4405 4850 4410 4880
rect 4440 4850 4445 4880
rect 4405 4845 4445 4850
rect 4605 4950 4645 4955
rect 4605 4920 4610 4950
rect 4640 4920 4645 4950
rect 4605 4880 4645 4920
rect 4605 4850 4610 4880
rect 4640 4850 4645 4880
rect 4605 4845 4645 4850
rect 4805 4950 4845 4955
rect 4805 4920 4810 4950
rect 4840 4920 4845 4950
rect 4805 4880 4845 4920
rect 4805 4850 4810 4880
rect 4840 4850 4845 4880
rect 4805 4845 4845 4850
rect 5005 4950 5045 4955
rect 5005 4920 5010 4950
rect 5040 4920 5045 4950
rect 5005 4880 5045 4920
rect 5005 4850 5010 4880
rect 5040 4850 5045 4880
rect 5005 4845 5045 4850
rect 5205 4950 5245 4955
rect 5205 4920 5210 4950
rect 5240 4920 5245 4950
rect 5205 4880 5245 4920
rect 5205 4850 5210 4880
rect 5240 4850 5245 4880
rect 5205 4845 5245 4850
rect 5405 4950 5445 4955
rect 5405 4920 5410 4950
rect 5440 4920 5445 4950
rect 5405 4880 5445 4920
rect 5405 4850 5410 4880
rect 5440 4850 5445 4880
rect 5405 4845 5445 4850
rect 5605 4950 5645 4955
rect 5605 4920 5610 4950
rect 5640 4920 5645 4950
rect 5605 4880 5645 4920
rect 5605 4850 5610 4880
rect 5640 4850 5645 4880
rect 5605 4845 5645 4850
rect 5805 4950 5845 4955
rect 5805 4920 5810 4950
rect 5840 4920 5845 4950
rect 5805 4880 5845 4920
rect 5805 4850 5810 4880
rect 5840 4850 5845 4880
rect 5805 4845 5845 4850
rect 6005 4950 6045 4955
rect 6005 4920 6010 4950
rect 6040 4920 6045 4950
rect 6005 4880 6045 4920
rect 6005 4850 6010 4880
rect 6040 4850 6045 4880
rect 6005 4845 6045 4850
rect 6205 4950 6245 4955
rect 6205 4920 6210 4950
rect 6240 4920 6245 4950
rect 6205 4880 6245 4920
rect 6205 4850 6210 4880
rect 6240 4850 6245 4880
rect 6205 4845 6245 4850
rect 6405 4950 6445 4955
rect 6405 4920 6410 4950
rect 6440 4920 6445 4950
rect 6405 4880 6445 4920
rect 6405 4850 6410 4880
rect 6440 4850 6445 4880
rect 6405 4845 6445 4850
rect -195 4765 -155 4770
rect -195 4735 -190 4765
rect -160 4735 -155 4765
rect -195 4695 -155 4735
rect -195 4665 -190 4695
rect -160 4665 -155 4695
rect -195 4660 -155 4665
rect 5 4765 45 4770
rect 5 4735 10 4765
rect 40 4735 45 4765
rect 5 4695 45 4735
rect 5 4665 10 4695
rect 40 4665 45 4695
rect 5 4660 45 4665
rect 205 4765 245 4770
rect 205 4735 210 4765
rect 240 4735 245 4765
rect 205 4695 245 4735
rect 205 4665 210 4695
rect 240 4665 245 4695
rect 205 4660 245 4665
rect 405 4765 445 4770
rect 405 4735 410 4765
rect 440 4735 445 4765
rect 405 4695 445 4735
rect 405 4665 410 4695
rect 440 4665 445 4695
rect 405 4660 445 4665
rect 605 4765 645 4770
rect 605 4735 610 4765
rect 640 4735 645 4765
rect 605 4695 645 4735
rect 605 4665 610 4695
rect 640 4665 645 4695
rect 605 4660 645 4665
rect 805 4765 845 4770
rect 805 4735 810 4765
rect 840 4735 845 4765
rect 805 4695 845 4735
rect 805 4665 810 4695
rect 840 4665 845 4695
rect 805 4660 845 4665
rect 1005 4765 1045 4770
rect 1005 4735 1010 4765
rect 1040 4735 1045 4765
rect 1005 4695 1045 4735
rect 1005 4665 1010 4695
rect 1040 4665 1045 4695
rect 1005 4660 1045 4665
rect 1205 4765 1245 4770
rect 1205 4735 1210 4765
rect 1240 4735 1245 4765
rect 1205 4695 1245 4735
rect 1205 4665 1210 4695
rect 1240 4665 1245 4695
rect 1205 4660 1245 4665
rect 1405 4765 1445 4770
rect 1405 4735 1410 4765
rect 1440 4735 1445 4765
rect 1405 4695 1445 4735
rect 1405 4665 1410 4695
rect 1440 4665 1445 4695
rect 1405 4660 1445 4665
rect 1605 4765 1645 4770
rect 1605 4735 1610 4765
rect 1640 4735 1645 4765
rect 1605 4695 1645 4735
rect 1605 4665 1610 4695
rect 1640 4665 1645 4695
rect 1605 4660 1645 4665
rect 1805 4765 1845 4770
rect 1805 4735 1810 4765
rect 1840 4735 1845 4765
rect 1805 4695 1845 4735
rect 1805 4665 1810 4695
rect 1840 4665 1845 4695
rect 1805 4660 1845 4665
rect 2005 4765 2045 4770
rect 2005 4735 2010 4765
rect 2040 4735 2045 4765
rect 2005 4695 2045 4735
rect 2005 4665 2010 4695
rect 2040 4665 2045 4695
rect 2005 4660 2045 4665
rect 2205 4765 2245 4770
rect 2205 4735 2210 4765
rect 2240 4735 2245 4765
rect 2205 4695 2245 4735
rect 2205 4665 2210 4695
rect 2240 4665 2245 4695
rect 2205 4660 2245 4665
rect 2405 4765 2445 4770
rect 2405 4735 2410 4765
rect 2440 4735 2445 4765
rect 2405 4695 2445 4735
rect 2405 4665 2410 4695
rect 2440 4665 2445 4695
rect 2405 4660 2445 4665
rect 2605 4765 2645 4770
rect 2605 4735 2610 4765
rect 2640 4735 2645 4765
rect 2605 4695 2645 4735
rect 2605 4665 2610 4695
rect 2640 4665 2645 4695
rect 2605 4660 2645 4665
rect 2805 4765 2845 4770
rect 2805 4735 2810 4765
rect 2840 4735 2845 4765
rect 2805 4695 2845 4735
rect 2805 4665 2810 4695
rect 2840 4665 2845 4695
rect 2805 4660 2845 4665
rect 3005 4765 3045 4770
rect 3005 4735 3010 4765
rect 3040 4735 3045 4765
rect 3005 4695 3045 4735
rect 3005 4665 3010 4695
rect 3040 4665 3045 4695
rect 3005 4660 3045 4665
rect 3205 4765 3245 4770
rect 3205 4735 3210 4765
rect 3240 4735 3245 4765
rect 3205 4695 3245 4735
rect 3205 4665 3210 4695
rect 3240 4665 3245 4695
rect 3205 4660 3245 4665
rect 3405 4765 3445 4770
rect 3405 4735 3410 4765
rect 3440 4735 3445 4765
rect 3405 4695 3445 4735
rect 3405 4665 3410 4695
rect 3440 4665 3445 4695
rect 3405 4660 3445 4665
rect 3605 4765 3645 4770
rect 3605 4735 3610 4765
rect 3640 4735 3645 4765
rect 3605 4695 3645 4735
rect 3605 4665 3610 4695
rect 3640 4665 3645 4695
rect 3605 4660 3645 4665
rect 3805 4765 3845 4770
rect 3805 4735 3810 4765
rect 3840 4735 3845 4765
rect 3805 4695 3845 4735
rect 3805 4665 3810 4695
rect 3840 4665 3845 4695
rect 3805 4660 3845 4665
rect 4005 4765 4045 4770
rect 4005 4735 4010 4765
rect 4040 4735 4045 4765
rect 4005 4695 4045 4735
rect 4005 4665 4010 4695
rect 4040 4665 4045 4695
rect 4005 4660 4045 4665
rect 4205 4765 4245 4770
rect 4205 4735 4210 4765
rect 4240 4735 4245 4765
rect 4205 4695 4245 4735
rect 4205 4665 4210 4695
rect 4240 4665 4245 4695
rect 4205 4660 4245 4665
rect 4405 4765 4445 4770
rect 4405 4735 4410 4765
rect 4440 4735 4445 4765
rect 4405 4695 4445 4735
rect 4405 4665 4410 4695
rect 4440 4665 4445 4695
rect 4405 4660 4445 4665
rect 4605 4765 4645 4770
rect 4605 4735 4610 4765
rect 4640 4735 4645 4765
rect 4605 4695 4645 4735
rect 4605 4665 4610 4695
rect 4640 4665 4645 4695
rect 4605 4660 4645 4665
rect 4805 4765 4845 4770
rect 4805 4735 4810 4765
rect 4840 4735 4845 4765
rect 4805 4695 4845 4735
rect 4805 4665 4810 4695
rect 4840 4665 4845 4695
rect 4805 4660 4845 4665
rect 5005 4765 5045 4770
rect 5005 4735 5010 4765
rect 5040 4735 5045 4765
rect 5005 4695 5045 4735
rect 5005 4665 5010 4695
rect 5040 4665 5045 4695
rect 5005 4660 5045 4665
rect 5205 4765 5245 4770
rect 5205 4735 5210 4765
rect 5240 4735 5245 4765
rect 5205 4695 5245 4735
rect 5205 4665 5210 4695
rect 5240 4665 5245 4695
rect 5205 4660 5245 4665
rect 5405 4765 5445 4770
rect 5405 4735 5410 4765
rect 5440 4735 5445 4765
rect 5405 4695 5445 4735
rect 5405 4665 5410 4695
rect 5440 4665 5445 4695
rect 5405 4660 5445 4665
rect 5605 4765 5645 4770
rect 5605 4735 5610 4765
rect 5640 4735 5645 4765
rect 5605 4695 5645 4735
rect 5605 4665 5610 4695
rect 5640 4665 5645 4695
rect 5605 4660 5645 4665
rect 5805 4765 5845 4770
rect 5805 4735 5810 4765
rect 5840 4735 5845 4765
rect 5805 4695 5845 4735
rect 5805 4665 5810 4695
rect 5840 4665 5845 4695
rect 5805 4660 5845 4665
rect 6005 4765 6045 4770
rect 6005 4735 6010 4765
rect 6040 4735 6045 4765
rect 6005 4695 6045 4735
rect 6005 4665 6010 4695
rect 6040 4665 6045 4695
rect 6005 4660 6045 4665
rect 6205 4765 6245 4770
rect 6205 4735 6210 4765
rect 6240 4735 6245 4765
rect 6205 4695 6245 4735
rect 6205 4665 6210 4695
rect 6240 4665 6245 4695
rect 6205 4660 6245 4665
rect 6405 4765 6445 4770
rect 6405 4735 6410 4765
rect 6440 4735 6445 4765
rect 6405 4695 6445 4735
rect 6405 4665 6410 4695
rect 6440 4665 6445 4695
rect 6405 4660 6445 4665
rect -195 4580 -155 4585
rect -195 4550 -190 4580
rect -160 4550 -155 4580
rect -195 4510 -155 4550
rect -195 4480 -190 4510
rect -160 4480 -155 4510
rect -195 4475 -155 4480
rect 5 4580 45 4585
rect 5 4550 10 4580
rect 40 4550 45 4580
rect 5 4510 45 4550
rect 5 4480 10 4510
rect 40 4480 45 4510
rect 5 4475 45 4480
rect 205 4580 245 4585
rect 205 4550 210 4580
rect 240 4550 245 4580
rect 205 4510 245 4550
rect 205 4480 210 4510
rect 240 4480 245 4510
rect 205 4475 245 4480
rect 405 4580 445 4585
rect 405 4550 410 4580
rect 440 4550 445 4580
rect 405 4510 445 4550
rect 405 4480 410 4510
rect 440 4480 445 4510
rect 405 4475 445 4480
rect 605 4580 645 4585
rect 605 4550 610 4580
rect 640 4550 645 4580
rect 605 4510 645 4550
rect 605 4480 610 4510
rect 640 4480 645 4510
rect 605 4475 645 4480
rect 805 4580 845 4585
rect 805 4550 810 4580
rect 840 4550 845 4580
rect 805 4510 845 4550
rect 805 4480 810 4510
rect 840 4480 845 4510
rect 805 4475 845 4480
rect 1005 4580 1045 4585
rect 1005 4550 1010 4580
rect 1040 4550 1045 4580
rect 1005 4510 1045 4550
rect 1005 4480 1010 4510
rect 1040 4480 1045 4510
rect 1005 4475 1045 4480
rect 1205 4580 1245 4585
rect 1205 4550 1210 4580
rect 1240 4550 1245 4580
rect 1205 4510 1245 4550
rect 1205 4480 1210 4510
rect 1240 4480 1245 4510
rect 1205 4475 1245 4480
rect 1405 4580 1445 4585
rect 1405 4550 1410 4580
rect 1440 4550 1445 4580
rect 1405 4510 1445 4550
rect 1405 4480 1410 4510
rect 1440 4480 1445 4510
rect 1405 4475 1445 4480
rect 1605 4580 1645 4585
rect 1605 4550 1610 4580
rect 1640 4550 1645 4580
rect 1605 4510 1645 4550
rect 1605 4480 1610 4510
rect 1640 4480 1645 4510
rect 1605 4475 1645 4480
rect 1805 4580 1845 4585
rect 1805 4550 1810 4580
rect 1840 4550 1845 4580
rect 1805 4510 1845 4550
rect 1805 4480 1810 4510
rect 1840 4480 1845 4510
rect 1805 4475 1845 4480
rect 2005 4580 2045 4585
rect 2005 4550 2010 4580
rect 2040 4550 2045 4580
rect 2005 4510 2045 4550
rect 2005 4480 2010 4510
rect 2040 4480 2045 4510
rect 2005 4475 2045 4480
rect 2205 4580 2245 4585
rect 2205 4550 2210 4580
rect 2240 4550 2245 4580
rect 2205 4510 2245 4550
rect 2205 4480 2210 4510
rect 2240 4480 2245 4510
rect 2205 4475 2245 4480
rect 2405 4580 2445 4585
rect 2405 4550 2410 4580
rect 2440 4550 2445 4580
rect 2405 4510 2445 4550
rect 2405 4480 2410 4510
rect 2440 4480 2445 4510
rect 2405 4475 2445 4480
rect 2605 4580 2645 4585
rect 2605 4550 2610 4580
rect 2640 4550 2645 4580
rect 2605 4510 2645 4550
rect 2605 4480 2610 4510
rect 2640 4480 2645 4510
rect 2605 4475 2645 4480
rect 2805 4580 2845 4585
rect 2805 4550 2810 4580
rect 2840 4550 2845 4580
rect 2805 4510 2845 4550
rect 2805 4480 2810 4510
rect 2840 4480 2845 4510
rect 2805 4475 2845 4480
rect 3005 4580 3045 4585
rect 3005 4550 3010 4580
rect 3040 4550 3045 4580
rect 3005 4510 3045 4550
rect 3005 4480 3010 4510
rect 3040 4480 3045 4510
rect 3005 4475 3045 4480
rect 3205 4580 3245 4585
rect 3205 4550 3210 4580
rect 3240 4550 3245 4580
rect 3205 4510 3245 4550
rect 3205 4480 3210 4510
rect 3240 4480 3245 4510
rect 3205 4475 3245 4480
rect 3405 4580 3445 4585
rect 3405 4550 3410 4580
rect 3440 4550 3445 4580
rect 3405 4510 3445 4550
rect 3405 4480 3410 4510
rect 3440 4480 3445 4510
rect 3405 4475 3445 4480
rect 3605 4580 3645 4585
rect 3605 4550 3610 4580
rect 3640 4550 3645 4580
rect 3605 4510 3645 4550
rect 3605 4480 3610 4510
rect 3640 4480 3645 4510
rect 3605 4475 3645 4480
rect 3805 4580 3845 4585
rect 3805 4550 3810 4580
rect 3840 4550 3845 4580
rect 3805 4510 3845 4550
rect 3805 4480 3810 4510
rect 3840 4480 3845 4510
rect 3805 4475 3845 4480
rect 4005 4580 4045 4585
rect 4005 4550 4010 4580
rect 4040 4550 4045 4580
rect 4005 4510 4045 4550
rect 4005 4480 4010 4510
rect 4040 4480 4045 4510
rect 4005 4475 4045 4480
rect 4205 4580 4245 4585
rect 4205 4550 4210 4580
rect 4240 4550 4245 4580
rect 4205 4510 4245 4550
rect 4205 4480 4210 4510
rect 4240 4480 4245 4510
rect 4205 4475 4245 4480
rect 4405 4580 4445 4585
rect 4405 4550 4410 4580
rect 4440 4550 4445 4580
rect 4405 4510 4445 4550
rect 4405 4480 4410 4510
rect 4440 4480 4445 4510
rect 4405 4475 4445 4480
rect 4605 4580 4645 4585
rect 4605 4550 4610 4580
rect 4640 4550 4645 4580
rect 4605 4510 4645 4550
rect 4605 4480 4610 4510
rect 4640 4480 4645 4510
rect 4605 4475 4645 4480
rect 4805 4580 4845 4585
rect 4805 4550 4810 4580
rect 4840 4550 4845 4580
rect 4805 4510 4845 4550
rect 4805 4480 4810 4510
rect 4840 4480 4845 4510
rect 4805 4475 4845 4480
rect 5005 4580 5045 4585
rect 5005 4550 5010 4580
rect 5040 4550 5045 4580
rect 5005 4510 5045 4550
rect 5005 4480 5010 4510
rect 5040 4480 5045 4510
rect 5005 4475 5045 4480
rect 5205 4580 5245 4585
rect 5205 4550 5210 4580
rect 5240 4550 5245 4580
rect 5205 4510 5245 4550
rect 5205 4480 5210 4510
rect 5240 4480 5245 4510
rect 5205 4475 5245 4480
rect 5405 4580 5445 4585
rect 5405 4550 5410 4580
rect 5440 4550 5445 4580
rect 5405 4510 5445 4550
rect 5405 4480 5410 4510
rect 5440 4480 5445 4510
rect 5405 4475 5445 4480
rect 5605 4580 5645 4585
rect 5605 4550 5610 4580
rect 5640 4550 5645 4580
rect 5605 4510 5645 4550
rect 5605 4480 5610 4510
rect 5640 4480 5645 4510
rect 5605 4475 5645 4480
rect 5805 4580 5845 4585
rect 5805 4550 5810 4580
rect 5840 4550 5845 4580
rect 5805 4510 5845 4550
rect 5805 4480 5810 4510
rect 5840 4480 5845 4510
rect 5805 4475 5845 4480
rect 6005 4580 6045 4585
rect 6005 4550 6010 4580
rect 6040 4550 6045 4580
rect 6005 4510 6045 4550
rect 6005 4480 6010 4510
rect 6040 4480 6045 4510
rect 6005 4475 6045 4480
rect 6205 4580 6245 4585
rect 6205 4550 6210 4580
rect 6240 4550 6245 4580
rect 6205 4510 6245 4550
rect 6205 4480 6210 4510
rect 6240 4480 6245 4510
rect 6205 4475 6245 4480
rect 6405 4580 6445 4585
rect 6405 4550 6410 4580
rect 6440 4550 6445 4580
rect 6405 4510 6445 4550
rect 6405 4480 6410 4510
rect 6440 4480 6445 4510
rect 6405 4475 6445 4480
rect -195 4395 -155 4400
rect -195 4365 -190 4395
rect -160 4365 -155 4395
rect -195 4325 -155 4365
rect -195 4295 -190 4325
rect -160 4295 -155 4325
rect -195 4290 -155 4295
rect 5 4395 45 4400
rect 5 4365 10 4395
rect 40 4365 45 4395
rect 5 4325 45 4365
rect 5 4295 10 4325
rect 40 4295 45 4325
rect 5 4290 45 4295
rect 205 4395 245 4400
rect 205 4365 210 4395
rect 240 4365 245 4395
rect 205 4325 245 4365
rect 205 4295 210 4325
rect 240 4295 245 4325
rect 205 4290 245 4295
rect 405 4395 445 4400
rect 405 4365 410 4395
rect 440 4365 445 4395
rect 405 4325 445 4365
rect 405 4295 410 4325
rect 440 4295 445 4325
rect 405 4290 445 4295
rect 605 4395 645 4400
rect 605 4365 610 4395
rect 640 4365 645 4395
rect 605 4325 645 4365
rect 605 4295 610 4325
rect 640 4295 645 4325
rect 605 4290 645 4295
rect 805 4395 845 4400
rect 805 4365 810 4395
rect 840 4365 845 4395
rect 805 4325 845 4365
rect 805 4295 810 4325
rect 840 4295 845 4325
rect 805 4290 845 4295
rect 1005 4395 1045 4400
rect 1005 4365 1010 4395
rect 1040 4365 1045 4395
rect 1005 4325 1045 4365
rect 1005 4295 1010 4325
rect 1040 4295 1045 4325
rect 1005 4290 1045 4295
rect 1205 4395 1245 4400
rect 1205 4365 1210 4395
rect 1240 4365 1245 4395
rect 1205 4325 1245 4365
rect 1205 4295 1210 4325
rect 1240 4295 1245 4325
rect 1205 4290 1245 4295
rect 1405 4395 1445 4400
rect 1405 4365 1410 4395
rect 1440 4365 1445 4395
rect 1405 4325 1445 4365
rect 1405 4295 1410 4325
rect 1440 4295 1445 4325
rect 1405 4290 1445 4295
rect 1605 4395 1645 4400
rect 1605 4365 1610 4395
rect 1640 4365 1645 4395
rect 1605 4325 1645 4365
rect 1605 4295 1610 4325
rect 1640 4295 1645 4325
rect 1605 4290 1645 4295
rect 1805 4395 1845 4400
rect 1805 4365 1810 4395
rect 1840 4365 1845 4395
rect 1805 4325 1845 4365
rect 1805 4295 1810 4325
rect 1840 4295 1845 4325
rect 1805 4290 1845 4295
rect 2005 4395 2045 4400
rect 2005 4365 2010 4395
rect 2040 4365 2045 4395
rect 2005 4325 2045 4365
rect 2005 4295 2010 4325
rect 2040 4295 2045 4325
rect 2005 4290 2045 4295
rect 2205 4395 2245 4400
rect 2205 4365 2210 4395
rect 2240 4365 2245 4395
rect 2205 4325 2245 4365
rect 2205 4295 2210 4325
rect 2240 4295 2245 4325
rect 2205 4290 2245 4295
rect 2405 4395 2445 4400
rect 2405 4365 2410 4395
rect 2440 4365 2445 4395
rect 2405 4325 2445 4365
rect 2405 4295 2410 4325
rect 2440 4295 2445 4325
rect 2405 4290 2445 4295
rect 2605 4395 2645 4400
rect 2605 4365 2610 4395
rect 2640 4365 2645 4395
rect 2605 4325 2645 4365
rect 2605 4295 2610 4325
rect 2640 4295 2645 4325
rect 2605 4290 2645 4295
rect 2805 4395 2845 4400
rect 2805 4365 2810 4395
rect 2840 4365 2845 4395
rect 2805 4325 2845 4365
rect 2805 4295 2810 4325
rect 2840 4295 2845 4325
rect 2805 4290 2845 4295
rect 3005 4395 3045 4400
rect 3005 4365 3010 4395
rect 3040 4365 3045 4395
rect 3005 4325 3045 4365
rect 3005 4295 3010 4325
rect 3040 4295 3045 4325
rect 3005 4290 3045 4295
rect 3205 4395 3245 4400
rect 3205 4365 3210 4395
rect 3240 4365 3245 4395
rect 3205 4325 3245 4365
rect 3205 4295 3210 4325
rect 3240 4295 3245 4325
rect 3205 4290 3245 4295
rect 3405 4395 3445 4400
rect 3405 4365 3410 4395
rect 3440 4365 3445 4395
rect 3405 4325 3445 4365
rect 3405 4295 3410 4325
rect 3440 4295 3445 4325
rect 3405 4290 3445 4295
rect 3605 4395 3645 4400
rect 3605 4365 3610 4395
rect 3640 4365 3645 4395
rect 3605 4325 3645 4365
rect 3605 4295 3610 4325
rect 3640 4295 3645 4325
rect 3605 4290 3645 4295
rect 3805 4395 3845 4400
rect 3805 4365 3810 4395
rect 3840 4365 3845 4395
rect 3805 4325 3845 4365
rect 3805 4295 3810 4325
rect 3840 4295 3845 4325
rect 3805 4290 3845 4295
rect 4005 4395 4045 4400
rect 4005 4365 4010 4395
rect 4040 4365 4045 4395
rect 4005 4325 4045 4365
rect 4005 4295 4010 4325
rect 4040 4295 4045 4325
rect 4005 4290 4045 4295
rect 4205 4395 4245 4400
rect 4205 4365 4210 4395
rect 4240 4365 4245 4395
rect 4205 4325 4245 4365
rect 4205 4295 4210 4325
rect 4240 4295 4245 4325
rect 4205 4290 4245 4295
rect 4405 4395 4445 4400
rect 4405 4365 4410 4395
rect 4440 4365 4445 4395
rect 4405 4325 4445 4365
rect 4405 4295 4410 4325
rect 4440 4295 4445 4325
rect 4405 4290 4445 4295
rect 4605 4395 4645 4400
rect 4605 4365 4610 4395
rect 4640 4365 4645 4395
rect 4605 4325 4645 4365
rect 4605 4295 4610 4325
rect 4640 4295 4645 4325
rect 4605 4290 4645 4295
rect 4805 4395 4845 4400
rect 4805 4365 4810 4395
rect 4840 4365 4845 4395
rect 4805 4325 4845 4365
rect 4805 4295 4810 4325
rect 4840 4295 4845 4325
rect 4805 4290 4845 4295
rect 5005 4395 5045 4400
rect 5005 4365 5010 4395
rect 5040 4365 5045 4395
rect 5005 4325 5045 4365
rect 5005 4295 5010 4325
rect 5040 4295 5045 4325
rect 5005 4290 5045 4295
rect 5205 4395 5245 4400
rect 5205 4365 5210 4395
rect 5240 4365 5245 4395
rect 5205 4325 5245 4365
rect 5205 4295 5210 4325
rect 5240 4295 5245 4325
rect 5205 4290 5245 4295
rect 5405 4395 5445 4400
rect 5405 4365 5410 4395
rect 5440 4365 5445 4395
rect 5405 4325 5445 4365
rect 5405 4295 5410 4325
rect 5440 4295 5445 4325
rect 5405 4290 5445 4295
rect 5605 4395 5645 4400
rect 5605 4365 5610 4395
rect 5640 4365 5645 4395
rect 5605 4325 5645 4365
rect 5605 4295 5610 4325
rect 5640 4295 5645 4325
rect 5605 4290 5645 4295
rect 5805 4395 5845 4400
rect 5805 4365 5810 4395
rect 5840 4365 5845 4395
rect 5805 4325 5845 4365
rect 5805 4295 5810 4325
rect 5840 4295 5845 4325
rect 5805 4290 5845 4295
rect 6005 4395 6045 4400
rect 6005 4365 6010 4395
rect 6040 4365 6045 4395
rect 6005 4325 6045 4365
rect 6005 4295 6010 4325
rect 6040 4295 6045 4325
rect 6005 4290 6045 4295
rect 6205 4395 6245 4400
rect 6205 4365 6210 4395
rect 6240 4365 6245 4395
rect 6205 4325 6245 4365
rect 6205 4295 6210 4325
rect 6240 4295 6245 4325
rect 6205 4290 6245 4295
rect 6405 4395 6445 4400
rect 6405 4365 6410 4395
rect 6440 4365 6445 4395
rect 6405 4325 6445 4365
rect 6405 4295 6410 4325
rect 6440 4295 6445 4325
rect 6405 4290 6445 4295
rect -195 4210 -155 4215
rect -195 4180 -190 4210
rect -160 4180 -155 4210
rect -195 4140 -155 4180
rect -195 4110 -190 4140
rect -160 4110 -155 4140
rect -195 4105 -155 4110
rect 5 4210 45 4215
rect 5 4180 10 4210
rect 40 4180 45 4210
rect 5 4140 45 4180
rect 5 4110 10 4140
rect 40 4110 45 4140
rect 5 4105 45 4110
rect 205 4210 245 4215
rect 205 4180 210 4210
rect 240 4180 245 4210
rect 205 4140 245 4180
rect 205 4110 210 4140
rect 240 4110 245 4140
rect 205 4105 245 4110
rect 405 4210 445 4215
rect 405 4180 410 4210
rect 440 4180 445 4210
rect 405 4140 445 4180
rect 405 4110 410 4140
rect 440 4110 445 4140
rect 405 4105 445 4110
rect 605 4210 645 4215
rect 605 4180 610 4210
rect 640 4180 645 4210
rect 605 4140 645 4180
rect 605 4110 610 4140
rect 640 4110 645 4140
rect 605 4105 645 4110
rect 805 4210 845 4215
rect 805 4180 810 4210
rect 840 4180 845 4210
rect 805 4140 845 4180
rect 805 4110 810 4140
rect 840 4110 845 4140
rect 805 4105 845 4110
rect 1005 4210 1045 4215
rect 1005 4180 1010 4210
rect 1040 4180 1045 4210
rect 1005 4140 1045 4180
rect 1005 4110 1010 4140
rect 1040 4110 1045 4140
rect 1005 4105 1045 4110
rect 1205 4210 1245 4215
rect 1205 4180 1210 4210
rect 1240 4180 1245 4210
rect 1205 4140 1245 4180
rect 1205 4110 1210 4140
rect 1240 4110 1245 4140
rect 1205 4105 1245 4110
rect 1405 4210 1445 4215
rect 1405 4180 1410 4210
rect 1440 4180 1445 4210
rect 1405 4140 1445 4180
rect 1405 4110 1410 4140
rect 1440 4110 1445 4140
rect 1405 4105 1445 4110
rect 1605 4210 1645 4215
rect 1605 4180 1610 4210
rect 1640 4180 1645 4210
rect 1605 4140 1645 4180
rect 1605 4110 1610 4140
rect 1640 4110 1645 4140
rect 1605 4105 1645 4110
rect 1805 4210 1845 4215
rect 1805 4180 1810 4210
rect 1840 4180 1845 4210
rect 1805 4140 1845 4180
rect 1805 4110 1810 4140
rect 1840 4110 1845 4140
rect 1805 4105 1845 4110
rect 2005 4210 2045 4215
rect 2005 4180 2010 4210
rect 2040 4180 2045 4210
rect 2005 4140 2045 4180
rect 2005 4110 2010 4140
rect 2040 4110 2045 4140
rect 2005 4105 2045 4110
rect 2205 4210 2245 4215
rect 2205 4180 2210 4210
rect 2240 4180 2245 4210
rect 2205 4140 2245 4180
rect 2205 4110 2210 4140
rect 2240 4110 2245 4140
rect 2205 4105 2245 4110
rect 2405 4210 2445 4215
rect 2405 4180 2410 4210
rect 2440 4180 2445 4210
rect 2405 4140 2445 4180
rect 2405 4110 2410 4140
rect 2440 4110 2445 4140
rect 2405 4105 2445 4110
rect 2605 4210 2645 4215
rect 2605 4180 2610 4210
rect 2640 4180 2645 4210
rect 2605 4140 2645 4180
rect 2605 4110 2610 4140
rect 2640 4110 2645 4140
rect 2605 4105 2645 4110
rect 2805 4210 2845 4215
rect 2805 4180 2810 4210
rect 2840 4180 2845 4210
rect 2805 4140 2845 4180
rect 2805 4110 2810 4140
rect 2840 4110 2845 4140
rect 2805 4105 2845 4110
rect 3005 4210 3045 4215
rect 3005 4180 3010 4210
rect 3040 4180 3045 4210
rect 3005 4140 3045 4180
rect 3005 4110 3010 4140
rect 3040 4110 3045 4140
rect 3005 4105 3045 4110
rect 3205 4210 3245 4215
rect 3205 4180 3210 4210
rect 3240 4180 3245 4210
rect 3205 4140 3245 4180
rect 3205 4110 3210 4140
rect 3240 4110 3245 4140
rect 3205 4105 3245 4110
rect 3405 4210 3445 4215
rect 3405 4180 3410 4210
rect 3440 4180 3445 4210
rect 3405 4140 3445 4180
rect 3405 4110 3410 4140
rect 3440 4110 3445 4140
rect 3405 4105 3445 4110
rect 3605 4210 3645 4215
rect 3605 4180 3610 4210
rect 3640 4180 3645 4210
rect 3605 4140 3645 4180
rect 3605 4110 3610 4140
rect 3640 4110 3645 4140
rect 3605 4105 3645 4110
rect 3805 4210 3845 4215
rect 3805 4180 3810 4210
rect 3840 4180 3845 4210
rect 3805 4140 3845 4180
rect 3805 4110 3810 4140
rect 3840 4110 3845 4140
rect 3805 4105 3845 4110
rect 4005 4210 4045 4215
rect 4005 4180 4010 4210
rect 4040 4180 4045 4210
rect 4005 4140 4045 4180
rect 4005 4110 4010 4140
rect 4040 4110 4045 4140
rect 4005 4105 4045 4110
rect 4205 4210 4245 4215
rect 4205 4180 4210 4210
rect 4240 4180 4245 4210
rect 4205 4140 4245 4180
rect 4205 4110 4210 4140
rect 4240 4110 4245 4140
rect 4205 4105 4245 4110
rect 4405 4210 4445 4215
rect 4405 4180 4410 4210
rect 4440 4180 4445 4210
rect 4405 4140 4445 4180
rect 4405 4110 4410 4140
rect 4440 4110 4445 4140
rect 4405 4105 4445 4110
rect 4605 4210 4645 4215
rect 4605 4180 4610 4210
rect 4640 4180 4645 4210
rect 4605 4140 4645 4180
rect 4605 4110 4610 4140
rect 4640 4110 4645 4140
rect 4605 4105 4645 4110
rect 4805 4210 4845 4215
rect 4805 4180 4810 4210
rect 4840 4180 4845 4210
rect 4805 4140 4845 4180
rect 4805 4110 4810 4140
rect 4840 4110 4845 4140
rect 4805 4105 4845 4110
rect 5005 4210 5045 4215
rect 5005 4180 5010 4210
rect 5040 4180 5045 4210
rect 5005 4140 5045 4180
rect 5005 4110 5010 4140
rect 5040 4110 5045 4140
rect 5005 4105 5045 4110
rect 5205 4210 5245 4215
rect 5205 4180 5210 4210
rect 5240 4180 5245 4210
rect 5205 4140 5245 4180
rect 5205 4110 5210 4140
rect 5240 4110 5245 4140
rect 5205 4105 5245 4110
rect 5405 4210 5445 4215
rect 5405 4180 5410 4210
rect 5440 4180 5445 4210
rect 5405 4140 5445 4180
rect 5405 4110 5410 4140
rect 5440 4110 5445 4140
rect 5405 4105 5445 4110
rect 5605 4210 5645 4215
rect 5605 4180 5610 4210
rect 5640 4180 5645 4210
rect 5605 4140 5645 4180
rect 5605 4110 5610 4140
rect 5640 4110 5645 4140
rect 5605 4105 5645 4110
rect 5805 4210 5845 4215
rect 5805 4180 5810 4210
rect 5840 4180 5845 4210
rect 5805 4140 5845 4180
rect 5805 4110 5810 4140
rect 5840 4110 5845 4140
rect 5805 4105 5845 4110
rect 6005 4210 6045 4215
rect 6005 4180 6010 4210
rect 6040 4180 6045 4210
rect 6005 4140 6045 4180
rect 6005 4110 6010 4140
rect 6040 4110 6045 4140
rect 6005 4105 6045 4110
rect 6205 4210 6245 4215
rect 6205 4180 6210 4210
rect 6240 4180 6245 4210
rect 6205 4140 6245 4180
rect 6205 4110 6210 4140
rect 6240 4110 6245 4140
rect 6205 4105 6245 4110
rect 6405 4210 6445 4215
rect 6405 4180 6410 4210
rect 6440 4180 6445 4210
rect 6405 4140 6445 4180
rect 6405 4110 6410 4140
rect 6440 4110 6445 4140
rect 6405 4105 6445 4110
rect -195 4025 -155 4030
rect -195 3995 -190 4025
rect -160 3995 -155 4025
rect -195 3955 -155 3995
rect -195 3925 -190 3955
rect -160 3925 -155 3955
rect -195 3920 -155 3925
rect 5 4025 45 4030
rect 5 3995 10 4025
rect 40 3995 45 4025
rect 5 3955 45 3995
rect 5 3925 10 3955
rect 40 3925 45 3955
rect 5 3920 45 3925
rect 205 4025 245 4030
rect 205 3995 210 4025
rect 240 3995 245 4025
rect 205 3955 245 3995
rect 205 3925 210 3955
rect 240 3925 245 3955
rect 205 3920 245 3925
rect 405 4025 445 4030
rect 405 3995 410 4025
rect 440 3995 445 4025
rect 405 3955 445 3995
rect 405 3925 410 3955
rect 440 3925 445 3955
rect 405 3920 445 3925
rect 605 4025 645 4030
rect 605 3995 610 4025
rect 640 3995 645 4025
rect 605 3955 645 3995
rect 605 3925 610 3955
rect 640 3925 645 3955
rect 605 3920 645 3925
rect 805 4025 845 4030
rect 805 3995 810 4025
rect 840 3995 845 4025
rect 805 3955 845 3995
rect 805 3925 810 3955
rect 840 3925 845 3955
rect 805 3920 845 3925
rect 1005 4025 1045 4030
rect 1005 3995 1010 4025
rect 1040 3995 1045 4025
rect 1005 3955 1045 3995
rect 1005 3925 1010 3955
rect 1040 3925 1045 3955
rect 1005 3920 1045 3925
rect 1205 4025 1245 4030
rect 1205 3995 1210 4025
rect 1240 3995 1245 4025
rect 1205 3955 1245 3995
rect 1205 3925 1210 3955
rect 1240 3925 1245 3955
rect 1205 3920 1245 3925
rect 1405 4025 1445 4030
rect 1405 3995 1410 4025
rect 1440 3995 1445 4025
rect 1405 3955 1445 3995
rect 1405 3925 1410 3955
rect 1440 3925 1445 3955
rect 1405 3920 1445 3925
rect 1605 4025 1645 4030
rect 1605 3995 1610 4025
rect 1640 3995 1645 4025
rect 1605 3955 1645 3995
rect 1605 3925 1610 3955
rect 1640 3925 1645 3955
rect 1605 3920 1645 3925
rect 1805 4025 1845 4030
rect 1805 3995 1810 4025
rect 1840 3995 1845 4025
rect 1805 3955 1845 3995
rect 1805 3925 1810 3955
rect 1840 3925 1845 3955
rect 1805 3920 1845 3925
rect 2005 4025 2045 4030
rect 2005 3995 2010 4025
rect 2040 3995 2045 4025
rect 2005 3955 2045 3995
rect 2005 3925 2010 3955
rect 2040 3925 2045 3955
rect 2005 3920 2045 3925
rect 2205 4025 2245 4030
rect 2205 3995 2210 4025
rect 2240 3995 2245 4025
rect 2205 3955 2245 3995
rect 2205 3925 2210 3955
rect 2240 3925 2245 3955
rect 2205 3920 2245 3925
rect 2405 4025 2445 4030
rect 2405 3995 2410 4025
rect 2440 3995 2445 4025
rect 2405 3955 2445 3995
rect 2405 3925 2410 3955
rect 2440 3925 2445 3955
rect 2405 3920 2445 3925
rect 2605 4025 2645 4030
rect 2605 3995 2610 4025
rect 2640 3995 2645 4025
rect 2605 3955 2645 3995
rect 2605 3925 2610 3955
rect 2640 3925 2645 3955
rect 2605 3920 2645 3925
rect 2805 4025 2845 4030
rect 2805 3995 2810 4025
rect 2840 3995 2845 4025
rect 2805 3955 2845 3995
rect 2805 3925 2810 3955
rect 2840 3925 2845 3955
rect 2805 3920 2845 3925
rect 3005 4025 3045 4030
rect 3005 3995 3010 4025
rect 3040 3995 3045 4025
rect 3005 3955 3045 3995
rect 3005 3925 3010 3955
rect 3040 3925 3045 3955
rect 3005 3920 3045 3925
rect 3205 4025 3245 4030
rect 3205 3995 3210 4025
rect 3240 3995 3245 4025
rect 3205 3955 3245 3995
rect 3205 3925 3210 3955
rect 3240 3925 3245 3955
rect 3205 3920 3245 3925
rect 3405 4025 3445 4030
rect 3405 3995 3410 4025
rect 3440 3995 3445 4025
rect 3405 3955 3445 3995
rect 3405 3925 3410 3955
rect 3440 3925 3445 3955
rect 3405 3920 3445 3925
rect 3605 4025 3645 4030
rect 3605 3995 3610 4025
rect 3640 3995 3645 4025
rect 3605 3955 3645 3995
rect 3605 3925 3610 3955
rect 3640 3925 3645 3955
rect 3605 3920 3645 3925
rect 3805 4025 3845 4030
rect 3805 3995 3810 4025
rect 3840 3995 3845 4025
rect 3805 3955 3845 3995
rect 3805 3925 3810 3955
rect 3840 3925 3845 3955
rect 3805 3920 3845 3925
rect 4005 4025 4045 4030
rect 4005 3995 4010 4025
rect 4040 3995 4045 4025
rect 4005 3955 4045 3995
rect 4005 3925 4010 3955
rect 4040 3925 4045 3955
rect 4005 3920 4045 3925
rect 4205 4025 4245 4030
rect 4205 3995 4210 4025
rect 4240 3995 4245 4025
rect 4205 3955 4245 3995
rect 4205 3925 4210 3955
rect 4240 3925 4245 3955
rect 4205 3920 4245 3925
rect 4405 4025 4445 4030
rect 4405 3995 4410 4025
rect 4440 3995 4445 4025
rect 4405 3955 4445 3995
rect 4405 3925 4410 3955
rect 4440 3925 4445 3955
rect 4405 3920 4445 3925
rect 4605 4025 4645 4030
rect 4605 3995 4610 4025
rect 4640 3995 4645 4025
rect 4605 3955 4645 3995
rect 4605 3925 4610 3955
rect 4640 3925 4645 3955
rect 4605 3920 4645 3925
rect 4805 4025 4845 4030
rect 4805 3995 4810 4025
rect 4840 3995 4845 4025
rect 4805 3955 4845 3995
rect 4805 3925 4810 3955
rect 4840 3925 4845 3955
rect 4805 3920 4845 3925
rect 5005 4025 5045 4030
rect 5005 3995 5010 4025
rect 5040 3995 5045 4025
rect 5005 3955 5045 3995
rect 5005 3925 5010 3955
rect 5040 3925 5045 3955
rect 5005 3920 5045 3925
rect 5205 4025 5245 4030
rect 5205 3995 5210 4025
rect 5240 3995 5245 4025
rect 5205 3955 5245 3995
rect 5205 3925 5210 3955
rect 5240 3925 5245 3955
rect 5205 3920 5245 3925
rect 5405 4025 5445 4030
rect 5405 3995 5410 4025
rect 5440 3995 5445 4025
rect 5405 3955 5445 3995
rect 5405 3925 5410 3955
rect 5440 3925 5445 3955
rect 5405 3920 5445 3925
rect 5605 4025 5645 4030
rect 5605 3995 5610 4025
rect 5640 3995 5645 4025
rect 5605 3955 5645 3995
rect 5605 3925 5610 3955
rect 5640 3925 5645 3955
rect 5605 3920 5645 3925
rect 5805 4025 5845 4030
rect 5805 3995 5810 4025
rect 5840 3995 5845 4025
rect 5805 3955 5845 3995
rect 5805 3925 5810 3955
rect 5840 3925 5845 3955
rect 5805 3920 5845 3925
rect 6005 4025 6045 4030
rect 6005 3995 6010 4025
rect 6040 3995 6045 4025
rect 6005 3955 6045 3995
rect 6005 3925 6010 3955
rect 6040 3925 6045 3955
rect 6005 3920 6045 3925
rect 6205 4025 6245 4030
rect 6205 3995 6210 4025
rect 6240 3995 6245 4025
rect 6205 3955 6245 3995
rect 6205 3925 6210 3955
rect 6240 3925 6245 3955
rect 6205 3920 6245 3925
rect 6405 4025 6445 4030
rect 6405 3995 6410 4025
rect 6440 3995 6445 4025
rect 6405 3955 6445 3995
rect 6405 3925 6410 3955
rect 6440 3925 6445 3955
rect 6405 3920 6445 3925
rect -195 3840 -155 3845
rect -195 3810 -190 3840
rect -160 3810 -155 3840
rect -195 3770 -155 3810
rect -195 3740 -190 3770
rect -160 3740 -155 3770
rect -195 3735 -155 3740
rect 5 3840 45 3845
rect 5 3810 10 3840
rect 40 3810 45 3840
rect 5 3770 45 3810
rect 5 3740 10 3770
rect 40 3740 45 3770
rect 5 3735 45 3740
rect 205 3840 245 3845
rect 205 3810 210 3840
rect 240 3810 245 3840
rect 205 3770 245 3810
rect 205 3740 210 3770
rect 240 3740 245 3770
rect 205 3735 245 3740
rect 405 3840 445 3845
rect 405 3810 410 3840
rect 440 3810 445 3840
rect 405 3770 445 3810
rect 405 3740 410 3770
rect 440 3740 445 3770
rect 405 3735 445 3740
rect 605 3840 645 3845
rect 605 3810 610 3840
rect 640 3810 645 3840
rect 605 3770 645 3810
rect 605 3740 610 3770
rect 640 3740 645 3770
rect 605 3735 645 3740
rect 805 3840 845 3845
rect 805 3810 810 3840
rect 840 3810 845 3840
rect 805 3770 845 3810
rect 805 3740 810 3770
rect 840 3740 845 3770
rect 805 3735 845 3740
rect 1005 3840 1045 3845
rect 1005 3810 1010 3840
rect 1040 3810 1045 3840
rect 1005 3770 1045 3810
rect 1005 3740 1010 3770
rect 1040 3740 1045 3770
rect 1005 3735 1045 3740
rect 1205 3840 1245 3845
rect 1205 3810 1210 3840
rect 1240 3810 1245 3840
rect 1205 3770 1245 3810
rect 1205 3740 1210 3770
rect 1240 3740 1245 3770
rect 1205 3735 1245 3740
rect 1405 3840 1445 3845
rect 1405 3810 1410 3840
rect 1440 3810 1445 3840
rect 1405 3770 1445 3810
rect 1405 3740 1410 3770
rect 1440 3740 1445 3770
rect 1405 3735 1445 3740
rect 1605 3840 1645 3845
rect 1605 3810 1610 3840
rect 1640 3810 1645 3840
rect 1605 3770 1645 3810
rect 1605 3740 1610 3770
rect 1640 3740 1645 3770
rect 1605 3735 1645 3740
rect 1805 3840 1845 3845
rect 1805 3810 1810 3840
rect 1840 3810 1845 3840
rect 1805 3770 1845 3810
rect 1805 3740 1810 3770
rect 1840 3740 1845 3770
rect 1805 3735 1845 3740
rect 2005 3840 2045 3845
rect 2005 3810 2010 3840
rect 2040 3810 2045 3840
rect 2005 3770 2045 3810
rect 2005 3740 2010 3770
rect 2040 3740 2045 3770
rect 2005 3735 2045 3740
rect 2205 3840 2245 3845
rect 2205 3810 2210 3840
rect 2240 3810 2245 3840
rect 2205 3770 2245 3810
rect 2205 3740 2210 3770
rect 2240 3740 2245 3770
rect 2205 3735 2245 3740
rect 2405 3840 2445 3845
rect 2405 3810 2410 3840
rect 2440 3810 2445 3840
rect 2405 3770 2445 3810
rect 2405 3740 2410 3770
rect 2440 3740 2445 3770
rect 2405 3735 2445 3740
rect 2605 3840 2645 3845
rect 2605 3810 2610 3840
rect 2640 3810 2645 3840
rect 2605 3770 2645 3810
rect 2605 3740 2610 3770
rect 2640 3740 2645 3770
rect 2605 3735 2645 3740
rect 2805 3840 2845 3845
rect 2805 3810 2810 3840
rect 2840 3810 2845 3840
rect 2805 3770 2845 3810
rect 2805 3740 2810 3770
rect 2840 3740 2845 3770
rect 2805 3735 2845 3740
rect 3005 3840 3045 3845
rect 3005 3810 3010 3840
rect 3040 3810 3045 3840
rect 3005 3770 3045 3810
rect 3005 3740 3010 3770
rect 3040 3740 3045 3770
rect 3005 3735 3045 3740
rect 3205 3840 3245 3845
rect 3205 3810 3210 3840
rect 3240 3810 3245 3840
rect 3205 3770 3245 3810
rect 3205 3740 3210 3770
rect 3240 3740 3245 3770
rect 3205 3735 3245 3740
rect 3405 3840 3445 3845
rect 3405 3810 3410 3840
rect 3440 3810 3445 3840
rect 3405 3770 3445 3810
rect 3405 3740 3410 3770
rect 3440 3740 3445 3770
rect 3405 3735 3445 3740
rect 3605 3840 3645 3845
rect 3605 3810 3610 3840
rect 3640 3810 3645 3840
rect 3605 3770 3645 3810
rect 3605 3740 3610 3770
rect 3640 3740 3645 3770
rect 3605 3735 3645 3740
rect 3805 3840 3845 3845
rect 3805 3810 3810 3840
rect 3840 3810 3845 3840
rect 3805 3770 3845 3810
rect 3805 3740 3810 3770
rect 3840 3740 3845 3770
rect 3805 3735 3845 3740
rect 4005 3840 4045 3845
rect 4005 3810 4010 3840
rect 4040 3810 4045 3840
rect 4005 3770 4045 3810
rect 4005 3740 4010 3770
rect 4040 3740 4045 3770
rect 4005 3735 4045 3740
rect 4205 3840 4245 3845
rect 4205 3810 4210 3840
rect 4240 3810 4245 3840
rect 4205 3770 4245 3810
rect 4205 3740 4210 3770
rect 4240 3740 4245 3770
rect 4205 3735 4245 3740
rect 4405 3840 4445 3845
rect 4405 3810 4410 3840
rect 4440 3810 4445 3840
rect 4405 3770 4445 3810
rect 4405 3740 4410 3770
rect 4440 3740 4445 3770
rect 4405 3735 4445 3740
rect 4605 3840 4645 3845
rect 4605 3810 4610 3840
rect 4640 3810 4645 3840
rect 4605 3770 4645 3810
rect 4605 3740 4610 3770
rect 4640 3740 4645 3770
rect 4605 3735 4645 3740
rect 4805 3840 4845 3845
rect 4805 3810 4810 3840
rect 4840 3810 4845 3840
rect 4805 3770 4845 3810
rect 4805 3740 4810 3770
rect 4840 3740 4845 3770
rect 4805 3735 4845 3740
rect 5005 3840 5045 3845
rect 5005 3810 5010 3840
rect 5040 3810 5045 3840
rect 5005 3770 5045 3810
rect 5005 3740 5010 3770
rect 5040 3740 5045 3770
rect 5005 3735 5045 3740
rect 5205 3840 5245 3845
rect 5205 3810 5210 3840
rect 5240 3810 5245 3840
rect 5205 3770 5245 3810
rect 5205 3740 5210 3770
rect 5240 3740 5245 3770
rect 5205 3735 5245 3740
rect 5405 3840 5445 3845
rect 5405 3810 5410 3840
rect 5440 3810 5445 3840
rect 5405 3770 5445 3810
rect 5405 3740 5410 3770
rect 5440 3740 5445 3770
rect 5405 3735 5445 3740
rect 5605 3840 5645 3845
rect 5605 3810 5610 3840
rect 5640 3810 5645 3840
rect 5605 3770 5645 3810
rect 5605 3740 5610 3770
rect 5640 3740 5645 3770
rect 5605 3735 5645 3740
rect 5805 3840 5845 3845
rect 5805 3810 5810 3840
rect 5840 3810 5845 3840
rect 5805 3770 5845 3810
rect 5805 3740 5810 3770
rect 5840 3740 5845 3770
rect 5805 3735 5845 3740
rect 6005 3840 6045 3845
rect 6005 3810 6010 3840
rect 6040 3810 6045 3840
rect 6005 3770 6045 3810
rect 6005 3740 6010 3770
rect 6040 3740 6045 3770
rect 6005 3735 6045 3740
rect 6205 3840 6245 3845
rect 6205 3810 6210 3840
rect 6240 3810 6245 3840
rect 6205 3770 6245 3810
rect 6205 3740 6210 3770
rect 6240 3740 6245 3770
rect 6205 3735 6245 3740
rect 6405 3840 6445 3845
rect 6405 3810 6410 3840
rect 6440 3810 6445 3840
rect 6405 3770 6445 3810
rect 6405 3740 6410 3770
rect 6440 3740 6445 3770
rect 6405 3735 6445 3740
rect -195 3655 -155 3660
rect -195 3625 -190 3655
rect -160 3625 -155 3655
rect -195 3585 -155 3625
rect -195 3555 -190 3585
rect -160 3555 -155 3585
rect -195 3550 -155 3555
rect 5 3655 45 3660
rect 5 3625 10 3655
rect 40 3625 45 3655
rect 5 3585 45 3625
rect 5 3555 10 3585
rect 40 3555 45 3585
rect 5 3550 45 3555
rect 205 3655 245 3660
rect 205 3625 210 3655
rect 240 3625 245 3655
rect 205 3585 245 3625
rect 205 3555 210 3585
rect 240 3555 245 3585
rect 205 3550 245 3555
rect 405 3655 445 3660
rect 405 3625 410 3655
rect 440 3625 445 3655
rect 405 3585 445 3625
rect 405 3555 410 3585
rect 440 3555 445 3585
rect 405 3550 445 3555
rect 605 3655 645 3660
rect 605 3625 610 3655
rect 640 3625 645 3655
rect 605 3585 645 3625
rect 605 3555 610 3585
rect 640 3555 645 3585
rect 605 3550 645 3555
rect 805 3655 845 3660
rect 805 3625 810 3655
rect 840 3625 845 3655
rect 805 3585 845 3625
rect 805 3555 810 3585
rect 840 3555 845 3585
rect 805 3550 845 3555
rect 1005 3655 1045 3660
rect 1005 3625 1010 3655
rect 1040 3625 1045 3655
rect 1005 3585 1045 3625
rect 1005 3555 1010 3585
rect 1040 3555 1045 3585
rect 1005 3550 1045 3555
rect 1205 3655 1245 3660
rect 1205 3625 1210 3655
rect 1240 3625 1245 3655
rect 1205 3585 1245 3625
rect 1205 3555 1210 3585
rect 1240 3555 1245 3585
rect 1205 3550 1245 3555
rect 1405 3655 1445 3660
rect 1405 3625 1410 3655
rect 1440 3625 1445 3655
rect 1405 3585 1445 3625
rect 1405 3555 1410 3585
rect 1440 3555 1445 3585
rect 1405 3550 1445 3555
rect 1605 3655 1645 3660
rect 1605 3625 1610 3655
rect 1640 3625 1645 3655
rect 1605 3585 1645 3625
rect 1605 3555 1610 3585
rect 1640 3555 1645 3585
rect 1605 3550 1645 3555
rect 1805 3655 1845 3660
rect 1805 3625 1810 3655
rect 1840 3625 1845 3655
rect 1805 3585 1845 3625
rect 1805 3555 1810 3585
rect 1840 3555 1845 3585
rect 1805 3550 1845 3555
rect 2005 3655 2045 3660
rect 2005 3625 2010 3655
rect 2040 3625 2045 3655
rect 2005 3585 2045 3625
rect 2005 3555 2010 3585
rect 2040 3555 2045 3585
rect 2005 3550 2045 3555
rect 2205 3655 2245 3660
rect 2205 3625 2210 3655
rect 2240 3625 2245 3655
rect 2205 3585 2245 3625
rect 2205 3555 2210 3585
rect 2240 3555 2245 3585
rect 2205 3550 2245 3555
rect 2405 3655 2445 3660
rect 2405 3625 2410 3655
rect 2440 3625 2445 3655
rect 2405 3585 2445 3625
rect 2405 3555 2410 3585
rect 2440 3555 2445 3585
rect 2405 3550 2445 3555
rect 2605 3655 2645 3660
rect 2605 3625 2610 3655
rect 2640 3625 2645 3655
rect 2605 3585 2645 3625
rect 2605 3555 2610 3585
rect 2640 3555 2645 3585
rect 2605 3550 2645 3555
rect 2805 3655 2845 3660
rect 2805 3625 2810 3655
rect 2840 3625 2845 3655
rect 2805 3585 2845 3625
rect 2805 3555 2810 3585
rect 2840 3555 2845 3585
rect 2805 3550 2845 3555
rect 3005 3655 3045 3660
rect 3005 3625 3010 3655
rect 3040 3625 3045 3655
rect 3005 3585 3045 3625
rect 3005 3555 3010 3585
rect 3040 3555 3045 3585
rect 3005 3550 3045 3555
rect 3205 3655 3245 3660
rect 3205 3625 3210 3655
rect 3240 3625 3245 3655
rect 3205 3585 3245 3625
rect 3205 3555 3210 3585
rect 3240 3555 3245 3585
rect 3205 3550 3245 3555
rect 3405 3655 3445 3660
rect 3405 3625 3410 3655
rect 3440 3625 3445 3655
rect 3405 3585 3445 3625
rect 3405 3555 3410 3585
rect 3440 3555 3445 3585
rect 3405 3550 3445 3555
rect 3605 3655 3645 3660
rect 3605 3625 3610 3655
rect 3640 3625 3645 3655
rect 3605 3585 3645 3625
rect 3605 3555 3610 3585
rect 3640 3555 3645 3585
rect 3605 3550 3645 3555
rect 3805 3655 3845 3660
rect 3805 3625 3810 3655
rect 3840 3625 3845 3655
rect 3805 3585 3845 3625
rect 3805 3555 3810 3585
rect 3840 3555 3845 3585
rect 3805 3550 3845 3555
rect 4005 3655 4045 3660
rect 4005 3625 4010 3655
rect 4040 3625 4045 3655
rect 4005 3585 4045 3625
rect 4005 3555 4010 3585
rect 4040 3555 4045 3585
rect 4005 3550 4045 3555
rect 4205 3655 4245 3660
rect 4205 3625 4210 3655
rect 4240 3625 4245 3655
rect 4205 3585 4245 3625
rect 4205 3555 4210 3585
rect 4240 3555 4245 3585
rect 4205 3550 4245 3555
rect 4405 3655 4445 3660
rect 4405 3625 4410 3655
rect 4440 3625 4445 3655
rect 4405 3585 4445 3625
rect 4405 3555 4410 3585
rect 4440 3555 4445 3585
rect 4405 3550 4445 3555
rect 4605 3655 4645 3660
rect 4605 3625 4610 3655
rect 4640 3625 4645 3655
rect 4605 3585 4645 3625
rect 4605 3555 4610 3585
rect 4640 3555 4645 3585
rect 4605 3550 4645 3555
rect 4805 3655 4845 3660
rect 4805 3625 4810 3655
rect 4840 3625 4845 3655
rect 4805 3585 4845 3625
rect 4805 3555 4810 3585
rect 4840 3555 4845 3585
rect 4805 3550 4845 3555
rect 5005 3655 5045 3660
rect 5005 3625 5010 3655
rect 5040 3625 5045 3655
rect 5005 3585 5045 3625
rect 5005 3555 5010 3585
rect 5040 3555 5045 3585
rect 5005 3550 5045 3555
rect 5205 3655 5245 3660
rect 5205 3625 5210 3655
rect 5240 3625 5245 3655
rect 5205 3585 5245 3625
rect 5205 3555 5210 3585
rect 5240 3555 5245 3585
rect 5205 3550 5245 3555
rect 5405 3655 5445 3660
rect 5405 3625 5410 3655
rect 5440 3625 5445 3655
rect 5405 3585 5445 3625
rect 5405 3555 5410 3585
rect 5440 3555 5445 3585
rect 5405 3550 5445 3555
rect 5605 3655 5645 3660
rect 5605 3625 5610 3655
rect 5640 3625 5645 3655
rect 5605 3585 5645 3625
rect 5605 3555 5610 3585
rect 5640 3555 5645 3585
rect 5605 3550 5645 3555
rect 5805 3655 5845 3660
rect 5805 3625 5810 3655
rect 5840 3625 5845 3655
rect 5805 3585 5845 3625
rect 5805 3555 5810 3585
rect 5840 3555 5845 3585
rect 5805 3550 5845 3555
rect 6005 3655 6045 3660
rect 6005 3625 6010 3655
rect 6040 3625 6045 3655
rect 6005 3585 6045 3625
rect 6005 3555 6010 3585
rect 6040 3555 6045 3585
rect 6005 3550 6045 3555
rect 6205 3655 6245 3660
rect 6205 3625 6210 3655
rect 6240 3625 6245 3655
rect 6205 3585 6245 3625
rect 6205 3555 6210 3585
rect 6240 3555 6245 3585
rect 6205 3550 6245 3555
rect 6405 3655 6445 3660
rect 6405 3625 6410 3655
rect 6440 3625 6445 3655
rect 6405 3585 6445 3625
rect 6405 3555 6410 3585
rect 6440 3555 6445 3585
rect 6405 3550 6445 3555
rect -195 3470 -155 3475
rect -195 3440 -190 3470
rect -160 3440 -155 3470
rect -195 3400 -155 3440
rect -195 3370 -190 3400
rect -160 3370 -155 3400
rect -195 3365 -155 3370
rect 5 3470 45 3475
rect 5 3440 10 3470
rect 40 3440 45 3470
rect 5 3400 45 3440
rect 5 3370 10 3400
rect 40 3370 45 3400
rect 5 3365 45 3370
rect 205 3470 245 3475
rect 205 3440 210 3470
rect 240 3440 245 3470
rect 205 3400 245 3440
rect 205 3370 210 3400
rect 240 3370 245 3400
rect 205 3365 245 3370
rect 405 3470 445 3475
rect 405 3440 410 3470
rect 440 3440 445 3470
rect 405 3400 445 3440
rect 405 3370 410 3400
rect 440 3370 445 3400
rect 405 3365 445 3370
rect 605 3470 645 3475
rect 605 3440 610 3470
rect 640 3440 645 3470
rect 605 3400 645 3440
rect 605 3370 610 3400
rect 640 3370 645 3400
rect 605 3365 645 3370
rect 805 3470 845 3475
rect 805 3440 810 3470
rect 840 3440 845 3470
rect 805 3400 845 3440
rect 805 3370 810 3400
rect 840 3370 845 3400
rect 805 3365 845 3370
rect 1005 3470 1045 3475
rect 1005 3440 1010 3470
rect 1040 3440 1045 3470
rect 1005 3400 1045 3440
rect 1005 3370 1010 3400
rect 1040 3370 1045 3400
rect 1005 3365 1045 3370
rect 1205 3470 1245 3475
rect 1205 3440 1210 3470
rect 1240 3440 1245 3470
rect 1205 3400 1245 3440
rect 1205 3370 1210 3400
rect 1240 3370 1245 3400
rect 1205 3365 1245 3370
rect 1405 3470 1445 3475
rect 1405 3440 1410 3470
rect 1440 3440 1445 3470
rect 1405 3400 1445 3440
rect 1405 3370 1410 3400
rect 1440 3370 1445 3400
rect 1405 3365 1445 3370
rect 1605 3470 1645 3475
rect 1605 3440 1610 3470
rect 1640 3440 1645 3470
rect 1605 3400 1645 3440
rect 1605 3370 1610 3400
rect 1640 3370 1645 3400
rect 1605 3365 1645 3370
rect 1805 3470 1845 3475
rect 1805 3440 1810 3470
rect 1840 3440 1845 3470
rect 1805 3400 1845 3440
rect 1805 3370 1810 3400
rect 1840 3370 1845 3400
rect 1805 3365 1845 3370
rect 2005 3470 2045 3475
rect 2005 3440 2010 3470
rect 2040 3440 2045 3470
rect 2005 3400 2045 3440
rect 2005 3370 2010 3400
rect 2040 3370 2045 3400
rect 2005 3365 2045 3370
rect 2205 3470 2245 3475
rect 2205 3440 2210 3470
rect 2240 3440 2245 3470
rect 2205 3400 2245 3440
rect 2205 3370 2210 3400
rect 2240 3370 2245 3400
rect 2205 3365 2245 3370
rect 2405 3470 2445 3475
rect 2405 3440 2410 3470
rect 2440 3440 2445 3470
rect 2405 3400 2445 3440
rect 2405 3370 2410 3400
rect 2440 3370 2445 3400
rect 2405 3365 2445 3370
rect 2605 3470 2645 3475
rect 2605 3440 2610 3470
rect 2640 3440 2645 3470
rect 2605 3400 2645 3440
rect 2605 3370 2610 3400
rect 2640 3370 2645 3400
rect 2605 3365 2645 3370
rect 2805 3470 2845 3475
rect 2805 3440 2810 3470
rect 2840 3440 2845 3470
rect 2805 3400 2845 3440
rect 2805 3370 2810 3400
rect 2840 3370 2845 3400
rect 2805 3365 2845 3370
rect 3005 3470 3045 3475
rect 3005 3440 3010 3470
rect 3040 3440 3045 3470
rect 3005 3400 3045 3440
rect 3005 3370 3010 3400
rect 3040 3370 3045 3400
rect 3005 3365 3045 3370
rect 3205 3470 3245 3475
rect 3205 3440 3210 3470
rect 3240 3440 3245 3470
rect 3205 3400 3245 3440
rect 3205 3370 3210 3400
rect 3240 3370 3245 3400
rect 3205 3365 3245 3370
rect 3405 3470 3445 3475
rect 3405 3440 3410 3470
rect 3440 3440 3445 3470
rect 3405 3400 3445 3440
rect 3405 3370 3410 3400
rect 3440 3370 3445 3400
rect 3405 3365 3445 3370
rect 3605 3470 3645 3475
rect 3605 3440 3610 3470
rect 3640 3440 3645 3470
rect 3605 3400 3645 3440
rect 3605 3370 3610 3400
rect 3640 3370 3645 3400
rect 3605 3365 3645 3370
rect 3805 3470 3845 3475
rect 3805 3440 3810 3470
rect 3840 3440 3845 3470
rect 3805 3400 3845 3440
rect 3805 3370 3810 3400
rect 3840 3370 3845 3400
rect 3805 3365 3845 3370
rect 4005 3470 4045 3475
rect 4005 3440 4010 3470
rect 4040 3440 4045 3470
rect 4005 3400 4045 3440
rect 4005 3370 4010 3400
rect 4040 3370 4045 3400
rect 4005 3365 4045 3370
rect 4205 3470 4245 3475
rect 4205 3440 4210 3470
rect 4240 3440 4245 3470
rect 4205 3400 4245 3440
rect 4205 3370 4210 3400
rect 4240 3370 4245 3400
rect 4205 3365 4245 3370
rect 4405 3470 4445 3475
rect 4405 3440 4410 3470
rect 4440 3440 4445 3470
rect 4405 3400 4445 3440
rect 4405 3370 4410 3400
rect 4440 3370 4445 3400
rect 4405 3365 4445 3370
rect 4605 3470 4645 3475
rect 4605 3440 4610 3470
rect 4640 3440 4645 3470
rect 4605 3400 4645 3440
rect 4605 3370 4610 3400
rect 4640 3370 4645 3400
rect 4605 3365 4645 3370
rect 4805 3470 4845 3475
rect 4805 3440 4810 3470
rect 4840 3440 4845 3470
rect 4805 3400 4845 3440
rect 4805 3370 4810 3400
rect 4840 3370 4845 3400
rect 4805 3365 4845 3370
rect 5005 3470 5045 3475
rect 5005 3440 5010 3470
rect 5040 3440 5045 3470
rect 5005 3400 5045 3440
rect 5005 3370 5010 3400
rect 5040 3370 5045 3400
rect 5005 3365 5045 3370
rect 5205 3470 5245 3475
rect 5205 3440 5210 3470
rect 5240 3440 5245 3470
rect 5205 3400 5245 3440
rect 5205 3370 5210 3400
rect 5240 3370 5245 3400
rect 5205 3365 5245 3370
rect 5405 3470 5445 3475
rect 5405 3440 5410 3470
rect 5440 3440 5445 3470
rect 5405 3400 5445 3440
rect 5405 3370 5410 3400
rect 5440 3370 5445 3400
rect 5405 3365 5445 3370
rect 5605 3470 5645 3475
rect 5605 3440 5610 3470
rect 5640 3440 5645 3470
rect 5605 3400 5645 3440
rect 5605 3370 5610 3400
rect 5640 3370 5645 3400
rect 5605 3365 5645 3370
rect 5805 3470 5845 3475
rect 5805 3440 5810 3470
rect 5840 3440 5845 3470
rect 5805 3400 5845 3440
rect 5805 3370 5810 3400
rect 5840 3370 5845 3400
rect 5805 3365 5845 3370
rect 6005 3470 6045 3475
rect 6005 3440 6010 3470
rect 6040 3440 6045 3470
rect 6005 3400 6045 3440
rect 6005 3370 6010 3400
rect 6040 3370 6045 3400
rect 6005 3365 6045 3370
rect 6205 3470 6245 3475
rect 6205 3440 6210 3470
rect 6240 3440 6245 3470
rect 6205 3400 6245 3440
rect 6205 3370 6210 3400
rect 6240 3370 6245 3400
rect 6205 3365 6245 3370
rect 6405 3470 6445 3475
rect 6405 3440 6410 3470
rect 6440 3440 6445 3470
rect 6405 3400 6445 3440
rect 6405 3370 6410 3400
rect 6440 3370 6445 3400
rect 6405 3365 6445 3370
rect -195 3285 -155 3290
rect -195 3255 -190 3285
rect -160 3255 -155 3285
rect -195 3215 -155 3255
rect -195 3185 -190 3215
rect -160 3185 -155 3215
rect -195 3180 -155 3185
rect 5 3285 45 3290
rect 5 3255 10 3285
rect 40 3255 45 3285
rect 5 3215 45 3255
rect 5 3185 10 3215
rect 40 3185 45 3215
rect 5 3180 45 3185
rect 205 3285 245 3290
rect 205 3255 210 3285
rect 240 3255 245 3285
rect 205 3215 245 3255
rect 205 3185 210 3215
rect 240 3185 245 3215
rect 205 3180 245 3185
rect 405 3285 445 3290
rect 405 3255 410 3285
rect 440 3255 445 3285
rect 405 3215 445 3255
rect 405 3185 410 3215
rect 440 3185 445 3215
rect 405 3180 445 3185
rect 605 3285 645 3290
rect 605 3255 610 3285
rect 640 3255 645 3285
rect 605 3215 645 3255
rect 605 3185 610 3215
rect 640 3185 645 3215
rect 605 3180 645 3185
rect 805 3285 845 3290
rect 805 3255 810 3285
rect 840 3255 845 3285
rect 805 3215 845 3255
rect 805 3185 810 3215
rect 840 3185 845 3215
rect 805 3180 845 3185
rect 1005 3285 1045 3290
rect 1005 3255 1010 3285
rect 1040 3255 1045 3285
rect 1005 3215 1045 3255
rect 1005 3185 1010 3215
rect 1040 3185 1045 3215
rect 1005 3180 1045 3185
rect 1205 3285 1245 3290
rect 1205 3255 1210 3285
rect 1240 3255 1245 3285
rect 1205 3215 1245 3255
rect 1205 3185 1210 3215
rect 1240 3185 1245 3215
rect 1205 3180 1245 3185
rect 1405 3285 1445 3290
rect 1405 3255 1410 3285
rect 1440 3255 1445 3285
rect 1405 3215 1445 3255
rect 1405 3185 1410 3215
rect 1440 3185 1445 3215
rect 1405 3180 1445 3185
rect 1605 3285 1645 3290
rect 1605 3255 1610 3285
rect 1640 3255 1645 3285
rect 1605 3215 1645 3255
rect 1605 3185 1610 3215
rect 1640 3185 1645 3215
rect 1605 3180 1645 3185
rect 1805 3285 1845 3290
rect 1805 3255 1810 3285
rect 1840 3255 1845 3285
rect 1805 3215 1845 3255
rect 1805 3185 1810 3215
rect 1840 3185 1845 3215
rect 1805 3180 1845 3185
rect 2005 3285 2045 3290
rect 2005 3255 2010 3285
rect 2040 3255 2045 3285
rect 2005 3215 2045 3255
rect 2005 3185 2010 3215
rect 2040 3185 2045 3215
rect 2005 3180 2045 3185
rect 2205 3285 2245 3290
rect 2205 3255 2210 3285
rect 2240 3255 2245 3285
rect 2205 3215 2245 3255
rect 2205 3185 2210 3215
rect 2240 3185 2245 3215
rect 2205 3180 2245 3185
rect 2405 3285 2445 3290
rect 2405 3255 2410 3285
rect 2440 3255 2445 3285
rect 2405 3215 2445 3255
rect 2405 3185 2410 3215
rect 2440 3185 2445 3215
rect 2405 3180 2445 3185
rect 2605 3285 2645 3290
rect 2605 3255 2610 3285
rect 2640 3255 2645 3285
rect 2605 3215 2645 3255
rect 2605 3185 2610 3215
rect 2640 3185 2645 3215
rect 2605 3180 2645 3185
rect 2805 3285 2845 3290
rect 2805 3255 2810 3285
rect 2840 3255 2845 3285
rect 2805 3215 2845 3255
rect 2805 3185 2810 3215
rect 2840 3185 2845 3215
rect 2805 3180 2845 3185
rect 3005 3285 3045 3290
rect 3005 3255 3010 3285
rect 3040 3255 3045 3285
rect 3005 3215 3045 3255
rect 3005 3185 3010 3215
rect 3040 3185 3045 3215
rect 3005 3180 3045 3185
rect 3205 3285 3245 3290
rect 3205 3255 3210 3285
rect 3240 3255 3245 3285
rect 3205 3215 3245 3255
rect 3205 3185 3210 3215
rect 3240 3185 3245 3215
rect 3205 3180 3245 3185
rect 3405 3285 3445 3290
rect 3405 3255 3410 3285
rect 3440 3255 3445 3285
rect 3405 3215 3445 3255
rect 3405 3185 3410 3215
rect 3440 3185 3445 3215
rect 3405 3180 3445 3185
rect 3605 3285 3645 3290
rect 3605 3255 3610 3285
rect 3640 3255 3645 3285
rect 3605 3215 3645 3255
rect 3605 3185 3610 3215
rect 3640 3185 3645 3215
rect 3605 3180 3645 3185
rect 3805 3285 3845 3290
rect 3805 3255 3810 3285
rect 3840 3255 3845 3285
rect 3805 3215 3845 3255
rect 3805 3185 3810 3215
rect 3840 3185 3845 3215
rect 3805 3180 3845 3185
rect 4005 3285 4045 3290
rect 4005 3255 4010 3285
rect 4040 3255 4045 3285
rect 4005 3215 4045 3255
rect 4005 3185 4010 3215
rect 4040 3185 4045 3215
rect 4005 3180 4045 3185
rect 4205 3285 4245 3290
rect 4205 3255 4210 3285
rect 4240 3255 4245 3285
rect 4205 3215 4245 3255
rect 4205 3185 4210 3215
rect 4240 3185 4245 3215
rect 4205 3180 4245 3185
rect 4405 3285 4445 3290
rect 4405 3255 4410 3285
rect 4440 3255 4445 3285
rect 4405 3215 4445 3255
rect 4405 3185 4410 3215
rect 4440 3185 4445 3215
rect 4405 3180 4445 3185
rect 4605 3285 4645 3290
rect 4605 3255 4610 3285
rect 4640 3255 4645 3285
rect 4605 3215 4645 3255
rect 4605 3185 4610 3215
rect 4640 3185 4645 3215
rect 4605 3180 4645 3185
rect 4805 3285 4845 3290
rect 4805 3255 4810 3285
rect 4840 3255 4845 3285
rect 4805 3215 4845 3255
rect 4805 3185 4810 3215
rect 4840 3185 4845 3215
rect 4805 3180 4845 3185
rect 5005 3285 5045 3290
rect 5005 3255 5010 3285
rect 5040 3255 5045 3285
rect 5005 3215 5045 3255
rect 5005 3185 5010 3215
rect 5040 3185 5045 3215
rect 5005 3180 5045 3185
rect 5205 3285 5245 3290
rect 5205 3255 5210 3285
rect 5240 3255 5245 3285
rect 5205 3215 5245 3255
rect 5205 3185 5210 3215
rect 5240 3185 5245 3215
rect 5205 3180 5245 3185
rect 5405 3285 5445 3290
rect 5405 3255 5410 3285
rect 5440 3255 5445 3285
rect 5405 3215 5445 3255
rect 5405 3185 5410 3215
rect 5440 3185 5445 3215
rect 5405 3180 5445 3185
rect 5605 3285 5645 3290
rect 5605 3255 5610 3285
rect 5640 3255 5645 3285
rect 5605 3215 5645 3255
rect 5605 3185 5610 3215
rect 5640 3185 5645 3215
rect 5605 3180 5645 3185
rect 5805 3285 5845 3290
rect 5805 3255 5810 3285
rect 5840 3255 5845 3285
rect 5805 3215 5845 3255
rect 5805 3185 5810 3215
rect 5840 3185 5845 3215
rect 5805 3180 5845 3185
rect 6005 3285 6045 3290
rect 6005 3255 6010 3285
rect 6040 3255 6045 3285
rect 6005 3215 6045 3255
rect 6005 3185 6010 3215
rect 6040 3185 6045 3215
rect 6005 3180 6045 3185
rect 6205 3285 6245 3290
rect 6205 3255 6210 3285
rect 6240 3255 6245 3285
rect 6205 3215 6245 3255
rect 6205 3185 6210 3215
rect 6240 3185 6245 3215
rect 6205 3180 6245 3185
rect 6405 3285 6445 3290
rect 6405 3255 6410 3285
rect 6440 3255 6445 3285
rect 6405 3215 6445 3255
rect 6405 3185 6410 3215
rect 6440 3185 6445 3215
rect 6405 3180 6445 3185
rect -195 3100 -155 3105
rect -195 3070 -190 3100
rect -160 3070 -155 3100
rect -195 3030 -155 3070
rect -195 3000 -190 3030
rect -160 3000 -155 3030
rect -195 2995 -155 3000
rect 5 3100 45 3105
rect 5 3070 10 3100
rect 40 3070 45 3100
rect 5 3030 45 3070
rect 5 3000 10 3030
rect 40 3000 45 3030
rect 5 2995 45 3000
rect 205 3100 245 3105
rect 205 3070 210 3100
rect 240 3070 245 3100
rect 205 3030 245 3070
rect 205 3000 210 3030
rect 240 3000 245 3030
rect 205 2995 245 3000
rect 405 3100 445 3105
rect 405 3070 410 3100
rect 440 3070 445 3100
rect 405 3030 445 3070
rect 405 3000 410 3030
rect 440 3000 445 3030
rect 405 2995 445 3000
rect 605 3100 645 3105
rect 605 3070 610 3100
rect 640 3070 645 3100
rect 605 3030 645 3070
rect 605 3000 610 3030
rect 640 3000 645 3030
rect 605 2995 645 3000
rect 805 3100 845 3105
rect 805 3070 810 3100
rect 840 3070 845 3100
rect 805 3030 845 3070
rect 805 3000 810 3030
rect 840 3000 845 3030
rect 805 2995 845 3000
rect 1005 3100 1045 3105
rect 1005 3070 1010 3100
rect 1040 3070 1045 3100
rect 1005 3030 1045 3070
rect 1005 3000 1010 3030
rect 1040 3000 1045 3030
rect 1005 2995 1045 3000
rect 1205 3100 1245 3105
rect 1205 3070 1210 3100
rect 1240 3070 1245 3100
rect 1205 3030 1245 3070
rect 1205 3000 1210 3030
rect 1240 3000 1245 3030
rect 1205 2995 1245 3000
rect 1405 3100 1445 3105
rect 1405 3070 1410 3100
rect 1440 3070 1445 3100
rect 1405 3030 1445 3070
rect 1405 3000 1410 3030
rect 1440 3000 1445 3030
rect 1405 2995 1445 3000
rect 1605 3100 1645 3105
rect 1605 3070 1610 3100
rect 1640 3070 1645 3100
rect 1605 3030 1645 3070
rect 1605 3000 1610 3030
rect 1640 3000 1645 3030
rect 1605 2995 1645 3000
rect 1805 3100 1845 3105
rect 1805 3070 1810 3100
rect 1840 3070 1845 3100
rect 1805 3030 1845 3070
rect 1805 3000 1810 3030
rect 1840 3000 1845 3030
rect 1805 2995 1845 3000
rect 2005 3100 2045 3105
rect 2005 3070 2010 3100
rect 2040 3070 2045 3100
rect 2005 3030 2045 3070
rect 2005 3000 2010 3030
rect 2040 3000 2045 3030
rect 2005 2995 2045 3000
rect 2205 3100 2245 3105
rect 2205 3070 2210 3100
rect 2240 3070 2245 3100
rect 2205 3030 2245 3070
rect 2205 3000 2210 3030
rect 2240 3000 2245 3030
rect 2205 2995 2245 3000
rect 2405 3100 2445 3105
rect 2405 3070 2410 3100
rect 2440 3070 2445 3100
rect 2405 3030 2445 3070
rect 2405 3000 2410 3030
rect 2440 3000 2445 3030
rect 2405 2995 2445 3000
rect 2605 3100 2645 3105
rect 2605 3070 2610 3100
rect 2640 3070 2645 3100
rect 2605 3030 2645 3070
rect 2605 3000 2610 3030
rect 2640 3000 2645 3030
rect 2605 2995 2645 3000
rect 2805 3100 2845 3105
rect 2805 3070 2810 3100
rect 2840 3070 2845 3100
rect 2805 3030 2845 3070
rect 2805 3000 2810 3030
rect 2840 3000 2845 3030
rect 2805 2995 2845 3000
rect 3005 3100 3045 3105
rect 3005 3070 3010 3100
rect 3040 3070 3045 3100
rect 3005 3030 3045 3070
rect 3005 3000 3010 3030
rect 3040 3000 3045 3030
rect 3005 2995 3045 3000
rect 3205 3100 3245 3105
rect 3205 3070 3210 3100
rect 3240 3070 3245 3100
rect 3205 3030 3245 3070
rect 3205 3000 3210 3030
rect 3240 3000 3245 3030
rect 3205 2995 3245 3000
rect 3405 3100 3445 3105
rect 3405 3070 3410 3100
rect 3440 3070 3445 3100
rect 3405 3030 3445 3070
rect 3405 3000 3410 3030
rect 3440 3000 3445 3030
rect 3405 2995 3445 3000
rect 3605 3100 3645 3105
rect 3605 3070 3610 3100
rect 3640 3070 3645 3100
rect 3605 3030 3645 3070
rect 3605 3000 3610 3030
rect 3640 3000 3645 3030
rect 3605 2995 3645 3000
rect 3805 3100 3845 3105
rect 3805 3070 3810 3100
rect 3840 3070 3845 3100
rect 3805 3030 3845 3070
rect 3805 3000 3810 3030
rect 3840 3000 3845 3030
rect 3805 2995 3845 3000
rect 4005 3100 4045 3105
rect 4005 3070 4010 3100
rect 4040 3070 4045 3100
rect 4005 3030 4045 3070
rect 4005 3000 4010 3030
rect 4040 3000 4045 3030
rect 4005 2995 4045 3000
rect 4205 3100 4245 3105
rect 4205 3070 4210 3100
rect 4240 3070 4245 3100
rect 4205 3030 4245 3070
rect 4205 3000 4210 3030
rect 4240 3000 4245 3030
rect 4205 2995 4245 3000
rect 4405 3100 4445 3105
rect 4405 3070 4410 3100
rect 4440 3070 4445 3100
rect 4405 3030 4445 3070
rect 4405 3000 4410 3030
rect 4440 3000 4445 3030
rect 4405 2995 4445 3000
rect 4605 3100 4645 3105
rect 4605 3070 4610 3100
rect 4640 3070 4645 3100
rect 4605 3030 4645 3070
rect 4605 3000 4610 3030
rect 4640 3000 4645 3030
rect 4605 2995 4645 3000
rect 4805 3100 4845 3105
rect 4805 3070 4810 3100
rect 4840 3070 4845 3100
rect 4805 3030 4845 3070
rect 4805 3000 4810 3030
rect 4840 3000 4845 3030
rect 4805 2995 4845 3000
rect 5005 3100 5045 3105
rect 5005 3070 5010 3100
rect 5040 3070 5045 3100
rect 5005 3030 5045 3070
rect 5005 3000 5010 3030
rect 5040 3000 5045 3030
rect 5005 2995 5045 3000
rect 5205 3100 5245 3105
rect 5205 3070 5210 3100
rect 5240 3070 5245 3100
rect 5205 3030 5245 3070
rect 5205 3000 5210 3030
rect 5240 3000 5245 3030
rect 5205 2995 5245 3000
rect 5405 3100 5445 3105
rect 5405 3070 5410 3100
rect 5440 3070 5445 3100
rect 5405 3030 5445 3070
rect 5405 3000 5410 3030
rect 5440 3000 5445 3030
rect 5405 2995 5445 3000
rect 5605 3100 5645 3105
rect 5605 3070 5610 3100
rect 5640 3070 5645 3100
rect 5605 3030 5645 3070
rect 5605 3000 5610 3030
rect 5640 3000 5645 3030
rect 5605 2995 5645 3000
rect 5805 3100 5845 3105
rect 5805 3070 5810 3100
rect 5840 3070 5845 3100
rect 5805 3030 5845 3070
rect 5805 3000 5810 3030
rect 5840 3000 5845 3030
rect 5805 2995 5845 3000
rect 6005 3100 6045 3105
rect 6005 3070 6010 3100
rect 6040 3070 6045 3100
rect 6005 3030 6045 3070
rect 6005 3000 6010 3030
rect 6040 3000 6045 3030
rect 6005 2995 6045 3000
rect 6205 3100 6245 3105
rect 6205 3070 6210 3100
rect 6240 3070 6245 3100
rect 6205 3030 6245 3070
rect 6205 3000 6210 3030
rect 6240 3000 6245 3030
rect 6205 2995 6245 3000
rect 6405 3100 6445 3105
rect 6405 3070 6410 3100
rect 6440 3070 6445 3100
rect 6405 3030 6445 3070
rect 6405 3000 6410 3030
rect 6440 3000 6445 3030
rect 6405 2995 6445 3000
rect -195 2915 -155 2920
rect -195 2885 -190 2915
rect -160 2885 -155 2915
rect -195 2845 -155 2885
rect -195 2815 -190 2845
rect -160 2815 -155 2845
rect -195 2810 -155 2815
rect 5 2915 45 2920
rect 5 2885 10 2915
rect 40 2885 45 2915
rect 5 2845 45 2885
rect 5 2815 10 2845
rect 40 2815 45 2845
rect 5 2810 45 2815
rect 205 2915 245 2920
rect 205 2885 210 2915
rect 240 2885 245 2915
rect 205 2845 245 2885
rect 205 2815 210 2845
rect 240 2815 245 2845
rect 205 2810 245 2815
rect 405 2915 445 2920
rect 405 2885 410 2915
rect 440 2885 445 2915
rect 405 2845 445 2885
rect 405 2815 410 2845
rect 440 2815 445 2845
rect 405 2810 445 2815
rect 605 2915 645 2920
rect 605 2885 610 2915
rect 640 2885 645 2915
rect 605 2845 645 2885
rect 605 2815 610 2845
rect 640 2815 645 2845
rect 605 2810 645 2815
rect 805 2915 845 2920
rect 805 2885 810 2915
rect 840 2885 845 2915
rect 805 2845 845 2885
rect 805 2815 810 2845
rect 840 2815 845 2845
rect 805 2810 845 2815
rect 1005 2915 1045 2920
rect 1005 2885 1010 2915
rect 1040 2885 1045 2915
rect 1005 2845 1045 2885
rect 1005 2815 1010 2845
rect 1040 2815 1045 2845
rect 1005 2810 1045 2815
rect 1205 2915 1245 2920
rect 1205 2885 1210 2915
rect 1240 2885 1245 2915
rect 1205 2845 1245 2885
rect 1205 2815 1210 2845
rect 1240 2815 1245 2845
rect 1205 2810 1245 2815
rect 1405 2915 1445 2920
rect 1405 2885 1410 2915
rect 1440 2885 1445 2915
rect 1405 2845 1445 2885
rect 1405 2815 1410 2845
rect 1440 2815 1445 2845
rect 1405 2810 1445 2815
rect 1605 2915 1645 2920
rect 1605 2885 1610 2915
rect 1640 2885 1645 2915
rect 1605 2845 1645 2885
rect 1605 2815 1610 2845
rect 1640 2815 1645 2845
rect 1605 2810 1645 2815
rect 1805 2915 1845 2920
rect 1805 2885 1810 2915
rect 1840 2885 1845 2915
rect 1805 2845 1845 2885
rect 1805 2815 1810 2845
rect 1840 2815 1845 2845
rect 1805 2810 1845 2815
rect 2005 2915 2045 2920
rect 2005 2885 2010 2915
rect 2040 2885 2045 2915
rect 2005 2845 2045 2885
rect 2005 2815 2010 2845
rect 2040 2815 2045 2845
rect 2005 2810 2045 2815
rect 2205 2915 2245 2920
rect 2205 2885 2210 2915
rect 2240 2885 2245 2915
rect 2205 2845 2245 2885
rect 2205 2815 2210 2845
rect 2240 2815 2245 2845
rect 2205 2810 2245 2815
rect 2405 2915 2445 2920
rect 2405 2885 2410 2915
rect 2440 2885 2445 2915
rect 2405 2845 2445 2885
rect 2405 2815 2410 2845
rect 2440 2815 2445 2845
rect 2405 2810 2445 2815
rect 2605 2915 2645 2920
rect 2605 2885 2610 2915
rect 2640 2885 2645 2915
rect 2605 2845 2645 2885
rect 2605 2815 2610 2845
rect 2640 2815 2645 2845
rect 2605 2810 2645 2815
rect 2805 2915 2845 2920
rect 2805 2885 2810 2915
rect 2840 2885 2845 2915
rect 2805 2845 2845 2885
rect 2805 2815 2810 2845
rect 2840 2815 2845 2845
rect 2805 2810 2845 2815
rect 3005 2915 3045 2920
rect 3005 2885 3010 2915
rect 3040 2885 3045 2915
rect 3005 2845 3045 2885
rect 3005 2815 3010 2845
rect 3040 2815 3045 2845
rect 3005 2810 3045 2815
rect 3205 2915 3245 2920
rect 3205 2885 3210 2915
rect 3240 2885 3245 2915
rect 3205 2845 3245 2885
rect 3205 2815 3210 2845
rect 3240 2815 3245 2845
rect 3205 2810 3245 2815
rect 3405 2915 3445 2920
rect 3405 2885 3410 2915
rect 3440 2885 3445 2915
rect 3405 2845 3445 2885
rect 3405 2815 3410 2845
rect 3440 2815 3445 2845
rect 3405 2810 3445 2815
rect 3605 2915 3645 2920
rect 3605 2885 3610 2915
rect 3640 2885 3645 2915
rect 3605 2845 3645 2885
rect 3605 2815 3610 2845
rect 3640 2815 3645 2845
rect 3605 2810 3645 2815
rect 3805 2915 3845 2920
rect 3805 2885 3810 2915
rect 3840 2885 3845 2915
rect 3805 2845 3845 2885
rect 3805 2815 3810 2845
rect 3840 2815 3845 2845
rect 3805 2810 3845 2815
rect 4005 2915 4045 2920
rect 4005 2885 4010 2915
rect 4040 2885 4045 2915
rect 4005 2845 4045 2885
rect 4005 2815 4010 2845
rect 4040 2815 4045 2845
rect 4005 2810 4045 2815
rect 4205 2915 4245 2920
rect 4205 2885 4210 2915
rect 4240 2885 4245 2915
rect 4205 2845 4245 2885
rect 4205 2815 4210 2845
rect 4240 2815 4245 2845
rect 4205 2810 4245 2815
rect 4405 2915 4445 2920
rect 4405 2885 4410 2915
rect 4440 2885 4445 2915
rect 4405 2845 4445 2885
rect 4405 2815 4410 2845
rect 4440 2815 4445 2845
rect 4405 2810 4445 2815
rect 4605 2915 4645 2920
rect 4605 2885 4610 2915
rect 4640 2885 4645 2915
rect 4605 2845 4645 2885
rect 4605 2815 4610 2845
rect 4640 2815 4645 2845
rect 4605 2810 4645 2815
rect 4805 2915 4845 2920
rect 4805 2885 4810 2915
rect 4840 2885 4845 2915
rect 4805 2845 4845 2885
rect 4805 2815 4810 2845
rect 4840 2815 4845 2845
rect 4805 2810 4845 2815
rect 5005 2915 5045 2920
rect 5005 2885 5010 2915
rect 5040 2885 5045 2915
rect 5005 2845 5045 2885
rect 5005 2815 5010 2845
rect 5040 2815 5045 2845
rect 5005 2810 5045 2815
rect 5205 2915 5245 2920
rect 5205 2885 5210 2915
rect 5240 2885 5245 2915
rect 5205 2845 5245 2885
rect 5205 2815 5210 2845
rect 5240 2815 5245 2845
rect 5205 2810 5245 2815
rect 5405 2915 5445 2920
rect 5405 2885 5410 2915
rect 5440 2885 5445 2915
rect 5405 2845 5445 2885
rect 5405 2815 5410 2845
rect 5440 2815 5445 2845
rect 5405 2810 5445 2815
rect 5605 2915 5645 2920
rect 5605 2885 5610 2915
rect 5640 2885 5645 2915
rect 5605 2845 5645 2885
rect 5605 2815 5610 2845
rect 5640 2815 5645 2845
rect 5605 2810 5645 2815
rect 5805 2915 5845 2920
rect 5805 2885 5810 2915
rect 5840 2885 5845 2915
rect 5805 2845 5845 2885
rect 5805 2815 5810 2845
rect 5840 2815 5845 2845
rect 5805 2810 5845 2815
rect 6005 2915 6045 2920
rect 6005 2885 6010 2915
rect 6040 2885 6045 2915
rect 6005 2845 6045 2885
rect 6005 2815 6010 2845
rect 6040 2815 6045 2845
rect 6005 2810 6045 2815
rect 6205 2915 6245 2920
rect 6205 2885 6210 2915
rect 6240 2885 6245 2915
rect 6205 2845 6245 2885
rect 6205 2815 6210 2845
rect 6240 2815 6245 2845
rect 6205 2810 6245 2815
rect 6405 2915 6445 2920
rect 6405 2885 6410 2915
rect 6440 2885 6445 2915
rect 6405 2845 6445 2885
rect 6405 2815 6410 2845
rect 6440 2815 6445 2845
rect 6405 2810 6445 2815
rect -195 2730 -155 2735
rect -195 2700 -190 2730
rect -160 2700 -155 2730
rect -195 2660 -155 2700
rect -195 2630 -190 2660
rect -160 2630 -155 2660
rect -195 2625 -155 2630
rect 5 2730 45 2735
rect 5 2700 10 2730
rect 40 2700 45 2730
rect 5 2660 45 2700
rect 5 2630 10 2660
rect 40 2630 45 2660
rect 5 2625 45 2630
rect 205 2730 245 2735
rect 205 2700 210 2730
rect 240 2700 245 2730
rect 205 2660 245 2700
rect 205 2630 210 2660
rect 240 2630 245 2660
rect 205 2625 245 2630
rect 405 2730 445 2735
rect 405 2700 410 2730
rect 440 2700 445 2730
rect 405 2660 445 2700
rect 405 2630 410 2660
rect 440 2630 445 2660
rect 405 2625 445 2630
rect 605 2730 645 2735
rect 605 2700 610 2730
rect 640 2700 645 2730
rect 605 2660 645 2700
rect 605 2630 610 2660
rect 640 2630 645 2660
rect 605 2625 645 2630
rect 805 2730 845 2735
rect 805 2700 810 2730
rect 840 2700 845 2730
rect 805 2660 845 2700
rect 805 2630 810 2660
rect 840 2630 845 2660
rect 805 2625 845 2630
rect 1005 2730 1045 2735
rect 1005 2700 1010 2730
rect 1040 2700 1045 2730
rect 1005 2660 1045 2700
rect 1005 2630 1010 2660
rect 1040 2630 1045 2660
rect 1005 2625 1045 2630
rect 1205 2730 1245 2735
rect 1205 2700 1210 2730
rect 1240 2700 1245 2730
rect 1205 2660 1245 2700
rect 1205 2630 1210 2660
rect 1240 2630 1245 2660
rect 1205 2625 1245 2630
rect 1405 2730 1445 2735
rect 1405 2700 1410 2730
rect 1440 2700 1445 2730
rect 1405 2660 1445 2700
rect 1405 2630 1410 2660
rect 1440 2630 1445 2660
rect 1405 2625 1445 2630
rect 1605 2730 1645 2735
rect 1605 2700 1610 2730
rect 1640 2700 1645 2730
rect 1605 2660 1645 2700
rect 1605 2630 1610 2660
rect 1640 2630 1645 2660
rect 1605 2625 1645 2630
rect 1805 2730 1845 2735
rect 1805 2700 1810 2730
rect 1840 2700 1845 2730
rect 1805 2660 1845 2700
rect 1805 2630 1810 2660
rect 1840 2630 1845 2660
rect 1805 2625 1845 2630
rect 2005 2730 2045 2735
rect 2005 2700 2010 2730
rect 2040 2700 2045 2730
rect 2005 2660 2045 2700
rect 2005 2630 2010 2660
rect 2040 2630 2045 2660
rect 2005 2625 2045 2630
rect 2205 2730 2245 2735
rect 2205 2700 2210 2730
rect 2240 2700 2245 2730
rect 2205 2660 2245 2700
rect 2205 2630 2210 2660
rect 2240 2630 2245 2660
rect 2205 2625 2245 2630
rect 2405 2730 2445 2735
rect 2405 2700 2410 2730
rect 2440 2700 2445 2730
rect 2405 2660 2445 2700
rect 2405 2630 2410 2660
rect 2440 2630 2445 2660
rect 2405 2625 2445 2630
rect 2605 2730 2645 2735
rect 2605 2700 2610 2730
rect 2640 2700 2645 2730
rect 2605 2660 2645 2700
rect 2605 2630 2610 2660
rect 2640 2630 2645 2660
rect 2605 2625 2645 2630
rect 2805 2730 2845 2735
rect 2805 2700 2810 2730
rect 2840 2700 2845 2730
rect 2805 2660 2845 2700
rect 2805 2630 2810 2660
rect 2840 2630 2845 2660
rect 2805 2625 2845 2630
rect 3005 2730 3045 2735
rect 3005 2700 3010 2730
rect 3040 2700 3045 2730
rect 3005 2660 3045 2700
rect 3005 2630 3010 2660
rect 3040 2630 3045 2660
rect 3005 2625 3045 2630
rect 3205 2730 3245 2735
rect 3205 2700 3210 2730
rect 3240 2700 3245 2730
rect 3205 2660 3245 2700
rect 3205 2630 3210 2660
rect 3240 2630 3245 2660
rect 3205 2625 3245 2630
rect 3405 2730 3445 2735
rect 3405 2700 3410 2730
rect 3440 2700 3445 2730
rect 3405 2660 3445 2700
rect 3405 2630 3410 2660
rect 3440 2630 3445 2660
rect 3405 2625 3445 2630
rect 3605 2730 3645 2735
rect 3605 2700 3610 2730
rect 3640 2700 3645 2730
rect 3605 2660 3645 2700
rect 3605 2630 3610 2660
rect 3640 2630 3645 2660
rect 3605 2625 3645 2630
rect 3805 2730 3845 2735
rect 3805 2700 3810 2730
rect 3840 2700 3845 2730
rect 3805 2660 3845 2700
rect 3805 2630 3810 2660
rect 3840 2630 3845 2660
rect 3805 2625 3845 2630
rect 4005 2730 4045 2735
rect 4005 2700 4010 2730
rect 4040 2700 4045 2730
rect 4005 2660 4045 2700
rect 4005 2630 4010 2660
rect 4040 2630 4045 2660
rect 4005 2625 4045 2630
rect 4205 2730 4245 2735
rect 4205 2700 4210 2730
rect 4240 2700 4245 2730
rect 4205 2660 4245 2700
rect 4205 2630 4210 2660
rect 4240 2630 4245 2660
rect 4205 2625 4245 2630
rect 4405 2730 4445 2735
rect 4405 2700 4410 2730
rect 4440 2700 4445 2730
rect 4405 2660 4445 2700
rect 4405 2630 4410 2660
rect 4440 2630 4445 2660
rect 4405 2625 4445 2630
rect 4605 2730 4645 2735
rect 4605 2700 4610 2730
rect 4640 2700 4645 2730
rect 4605 2660 4645 2700
rect 4605 2630 4610 2660
rect 4640 2630 4645 2660
rect 4605 2625 4645 2630
rect 4805 2730 4845 2735
rect 4805 2700 4810 2730
rect 4840 2700 4845 2730
rect 4805 2660 4845 2700
rect 4805 2630 4810 2660
rect 4840 2630 4845 2660
rect 4805 2625 4845 2630
rect 5005 2730 5045 2735
rect 5005 2700 5010 2730
rect 5040 2700 5045 2730
rect 5005 2660 5045 2700
rect 5005 2630 5010 2660
rect 5040 2630 5045 2660
rect 5005 2625 5045 2630
rect 5205 2730 5245 2735
rect 5205 2700 5210 2730
rect 5240 2700 5245 2730
rect 5205 2660 5245 2700
rect 5205 2630 5210 2660
rect 5240 2630 5245 2660
rect 5205 2625 5245 2630
rect 5405 2730 5445 2735
rect 5405 2700 5410 2730
rect 5440 2700 5445 2730
rect 5405 2660 5445 2700
rect 5405 2630 5410 2660
rect 5440 2630 5445 2660
rect 5405 2625 5445 2630
rect 5605 2730 5645 2735
rect 5605 2700 5610 2730
rect 5640 2700 5645 2730
rect 5605 2660 5645 2700
rect 5605 2630 5610 2660
rect 5640 2630 5645 2660
rect 5605 2625 5645 2630
rect 5805 2730 5845 2735
rect 5805 2700 5810 2730
rect 5840 2700 5845 2730
rect 5805 2660 5845 2700
rect 5805 2630 5810 2660
rect 5840 2630 5845 2660
rect 5805 2625 5845 2630
rect 6005 2730 6045 2735
rect 6005 2700 6010 2730
rect 6040 2700 6045 2730
rect 6005 2660 6045 2700
rect 6005 2630 6010 2660
rect 6040 2630 6045 2660
rect 6005 2625 6045 2630
rect 6205 2730 6245 2735
rect 6205 2700 6210 2730
rect 6240 2700 6245 2730
rect 6205 2660 6245 2700
rect 6205 2630 6210 2660
rect 6240 2630 6245 2660
rect 6205 2625 6245 2630
rect 6405 2730 6445 2735
rect 6405 2700 6410 2730
rect 6440 2700 6445 2730
rect 6405 2660 6445 2700
rect 6405 2630 6410 2660
rect 6440 2630 6445 2660
rect 6405 2625 6445 2630
rect -195 2545 -155 2550
rect -195 2515 -190 2545
rect -160 2515 -155 2545
rect -195 2475 -155 2515
rect -195 2445 -190 2475
rect -160 2445 -155 2475
rect -195 2440 -155 2445
rect 5 2545 45 2550
rect 5 2515 10 2545
rect 40 2515 45 2545
rect 5 2475 45 2515
rect 5 2445 10 2475
rect 40 2445 45 2475
rect 5 2440 45 2445
rect 205 2545 245 2550
rect 205 2515 210 2545
rect 240 2515 245 2545
rect 205 2475 245 2515
rect 205 2445 210 2475
rect 240 2445 245 2475
rect 205 2440 245 2445
rect 405 2545 445 2550
rect 405 2515 410 2545
rect 440 2515 445 2545
rect 405 2475 445 2515
rect 405 2445 410 2475
rect 440 2445 445 2475
rect 405 2440 445 2445
rect 605 2545 645 2550
rect 605 2515 610 2545
rect 640 2515 645 2545
rect 605 2475 645 2515
rect 605 2445 610 2475
rect 640 2445 645 2475
rect 605 2440 645 2445
rect 805 2545 845 2550
rect 805 2515 810 2545
rect 840 2515 845 2545
rect 805 2475 845 2515
rect 805 2445 810 2475
rect 840 2445 845 2475
rect 805 2440 845 2445
rect 1005 2545 1045 2550
rect 1005 2515 1010 2545
rect 1040 2515 1045 2545
rect 1005 2475 1045 2515
rect 1005 2445 1010 2475
rect 1040 2445 1045 2475
rect 1005 2440 1045 2445
rect 1205 2545 1245 2550
rect 1205 2515 1210 2545
rect 1240 2515 1245 2545
rect 1205 2475 1245 2515
rect 1205 2445 1210 2475
rect 1240 2445 1245 2475
rect 1205 2440 1245 2445
rect 1405 2545 1445 2550
rect 1405 2515 1410 2545
rect 1440 2515 1445 2545
rect 1405 2475 1445 2515
rect 1405 2445 1410 2475
rect 1440 2445 1445 2475
rect 1405 2440 1445 2445
rect 1605 2545 1645 2550
rect 1605 2515 1610 2545
rect 1640 2515 1645 2545
rect 1605 2475 1645 2515
rect 1605 2445 1610 2475
rect 1640 2445 1645 2475
rect 1605 2440 1645 2445
rect 1805 2545 1845 2550
rect 1805 2515 1810 2545
rect 1840 2515 1845 2545
rect 1805 2475 1845 2515
rect 1805 2445 1810 2475
rect 1840 2445 1845 2475
rect 1805 2440 1845 2445
rect 2005 2545 2045 2550
rect 2005 2515 2010 2545
rect 2040 2515 2045 2545
rect 2005 2475 2045 2515
rect 2005 2445 2010 2475
rect 2040 2445 2045 2475
rect 2005 2440 2045 2445
rect 2205 2545 2245 2550
rect 2205 2515 2210 2545
rect 2240 2515 2245 2545
rect 2205 2475 2245 2515
rect 2205 2445 2210 2475
rect 2240 2445 2245 2475
rect 2205 2440 2245 2445
rect 2405 2545 2445 2550
rect 2405 2515 2410 2545
rect 2440 2515 2445 2545
rect 2405 2475 2445 2515
rect 2405 2445 2410 2475
rect 2440 2445 2445 2475
rect 2405 2440 2445 2445
rect 2605 2545 2645 2550
rect 2605 2515 2610 2545
rect 2640 2515 2645 2545
rect 2605 2475 2645 2515
rect 2605 2445 2610 2475
rect 2640 2445 2645 2475
rect 2605 2440 2645 2445
rect 2805 2545 2845 2550
rect 2805 2515 2810 2545
rect 2840 2515 2845 2545
rect 2805 2475 2845 2515
rect 2805 2445 2810 2475
rect 2840 2445 2845 2475
rect 2805 2440 2845 2445
rect 3005 2545 3045 2550
rect 3005 2515 3010 2545
rect 3040 2515 3045 2545
rect 3005 2475 3045 2515
rect 3005 2445 3010 2475
rect 3040 2445 3045 2475
rect 3005 2440 3045 2445
rect 3205 2545 3245 2550
rect 3205 2515 3210 2545
rect 3240 2515 3245 2545
rect 3205 2475 3245 2515
rect 3205 2445 3210 2475
rect 3240 2445 3245 2475
rect 3205 2440 3245 2445
rect 3405 2545 3445 2550
rect 3405 2515 3410 2545
rect 3440 2515 3445 2545
rect 3405 2475 3445 2515
rect 3405 2445 3410 2475
rect 3440 2445 3445 2475
rect 3405 2440 3445 2445
rect 3605 2545 3645 2550
rect 3605 2515 3610 2545
rect 3640 2515 3645 2545
rect 3605 2475 3645 2515
rect 3605 2445 3610 2475
rect 3640 2445 3645 2475
rect 3605 2440 3645 2445
rect 3805 2545 3845 2550
rect 3805 2515 3810 2545
rect 3840 2515 3845 2545
rect 3805 2475 3845 2515
rect 3805 2445 3810 2475
rect 3840 2445 3845 2475
rect 3805 2440 3845 2445
rect 4005 2545 4045 2550
rect 4005 2515 4010 2545
rect 4040 2515 4045 2545
rect 4005 2475 4045 2515
rect 4005 2445 4010 2475
rect 4040 2445 4045 2475
rect 4005 2440 4045 2445
rect 4205 2545 4245 2550
rect 4205 2515 4210 2545
rect 4240 2515 4245 2545
rect 4205 2475 4245 2515
rect 4205 2445 4210 2475
rect 4240 2445 4245 2475
rect 4205 2440 4245 2445
rect 4405 2545 4445 2550
rect 4405 2515 4410 2545
rect 4440 2515 4445 2545
rect 4405 2475 4445 2515
rect 4405 2445 4410 2475
rect 4440 2445 4445 2475
rect 4405 2440 4445 2445
rect 4605 2545 4645 2550
rect 4605 2515 4610 2545
rect 4640 2515 4645 2545
rect 4605 2475 4645 2515
rect 4605 2445 4610 2475
rect 4640 2445 4645 2475
rect 4605 2440 4645 2445
rect 4805 2545 4845 2550
rect 4805 2515 4810 2545
rect 4840 2515 4845 2545
rect 4805 2475 4845 2515
rect 4805 2445 4810 2475
rect 4840 2445 4845 2475
rect 4805 2440 4845 2445
rect 5005 2545 5045 2550
rect 5005 2515 5010 2545
rect 5040 2515 5045 2545
rect 5005 2475 5045 2515
rect 5005 2445 5010 2475
rect 5040 2445 5045 2475
rect 5005 2440 5045 2445
rect 5205 2545 5245 2550
rect 5205 2515 5210 2545
rect 5240 2515 5245 2545
rect 5205 2475 5245 2515
rect 5205 2445 5210 2475
rect 5240 2445 5245 2475
rect 5205 2440 5245 2445
rect 5405 2545 5445 2550
rect 5405 2515 5410 2545
rect 5440 2515 5445 2545
rect 5405 2475 5445 2515
rect 5405 2445 5410 2475
rect 5440 2445 5445 2475
rect 5405 2440 5445 2445
rect 5605 2545 5645 2550
rect 5605 2515 5610 2545
rect 5640 2515 5645 2545
rect 5605 2475 5645 2515
rect 5605 2445 5610 2475
rect 5640 2445 5645 2475
rect 5605 2440 5645 2445
rect 5805 2545 5845 2550
rect 5805 2515 5810 2545
rect 5840 2515 5845 2545
rect 5805 2475 5845 2515
rect 5805 2445 5810 2475
rect 5840 2445 5845 2475
rect 5805 2440 5845 2445
rect 6005 2545 6045 2550
rect 6005 2515 6010 2545
rect 6040 2515 6045 2545
rect 6005 2475 6045 2515
rect 6005 2445 6010 2475
rect 6040 2445 6045 2475
rect 6005 2440 6045 2445
rect 6205 2545 6245 2550
rect 6205 2515 6210 2545
rect 6240 2515 6245 2545
rect 6205 2475 6245 2515
rect 6205 2445 6210 2475
rect 6240 2445 6245 2475
rect 6205 2440 6245 2445
rect 6405 2545 6445 2550
rect 6405 2515 6410 2545
rect 6440 2515 6445 2545
rect 6405 2475 6445 2515
rect 6405 2445 6410 2475
rect 6440 2445 6445 2475
rect 6405 2440 6445 2445
rect -195 2360 -155 2365
rect -195 2330 -190 2360
rect -160 2330 -155 2360
rect -195 2290 -155 2330
rect -195 2260 -190 2290
rect -160 2260 -155 2290
rect -195 2255 -155 2260
rect 5 2360 45 2365
rect 5 2330 10 2360
rect 40 2330 45 2360
rect 5 2290 45 2330
rect 5 2260 10 2290
rect 40 2260 45 2290
rect 5 2255 45 2260
rect 205 2360 245 2365
rect 205 2330 210 2360
rect 240 2330 245 2360
rect 205 2290 245 2330
rect 205 2260 210 2290
rect 240 2260 245 2290
rect 205 2255 245 2260
rect 405 2360 445 2365
rect 405 2330 410 2360
rect 440 2330 445 2360
rect 405 2290 445 2330
rect 405 2260 410 2290
rect 440 2260 445 2290
rect 405 2255 445 2260
rect 605 2360 645 2365
rect 605 2330 610 2360
rect 640 2330 645 2360
rect 605 2290 645 2330
rect 605 2260 610 2290
rect 640 2260 645 2290
rect 605 2255 645 2260
rect 805 2360 845 2365
rect 805 2330 810 2360
rect 840 2330 845 2360
rect 805 2290 845 2330
rect 805 2260 810 2290
rect 840 2260 845 2290
rect 805 2255 845 2260
rect 1005 2360 1045 2365
rect 1005 2330 1010 2360
rect 1040 2330 1045 2360
rect 1005 2290 1045 2330
rect 1005 2260 1010 2290
rect 1040 2260 1045 2290
rect 1005 2255 1045 2260
rect 1205 2360 1245 2365
rect 1205 2330 1210 2360
rect 1240 2330 1245 2360
rect 1205 2290 1245 2330
rect 1205 2260 1210 2290
rect 1240 2260 1245 2290
rect 1205 2255 1245 2260
rect 1405 2360 1445 2365
rect 1405 2330 1410 2360
rect 1440 2330 1445 2360
rect 1405 2290 1445 2330
rect 1405 2260 1410 2290
rect 1440 2260 1445 2290
rect 1405 2255 1445 2260
rect 1605 2360 1645 2365
rect 1605 2330 1610 2360
rect 1640 2330 1645 2360
rect 1605 2290 1645 2330
rect 1605 2260 1610 2290
rect 1640 2260 1645 2290
rect 1605 2255 1645 2260
rect 1805 2360 1845 2365
rect 1805 2330 1810 2360
rect 1840 2330 1845 2360
rect 1805 2290 1845 2330
rect 1805 2260 1810 2290
rect 1840 2260 1845 2290
rect 1805 2255 1845 2260
rect 2005 2360 2045 2365
rect 2005 2330 2010 2360
rect 2040 2330 2045 2360
rect 2005 2290 2045 2330
rect 2005 2260 2010 2290
rect 2040 2260 2045 2290
rect 2005 2255 2045 2260
rect 2205 2360 2245 2365
rect 2205 2330 2210 2360
rect 2240 2330 2245 2360
rect 2205 2290 2245 2330
rect 2205 2260 2210 2290
rect 2240 2260 2245 2290
rect 2205 2255 2245 2260
rect 2405 2360 2445 2365
rect 2405 2330 2410 2360
rect 2440 2330 2445 2360
rect 2405 2290 2445 2330
rect 2405 2260 2410 2290
rect 2440 2260 2445 2290
rect 2405 2255 2445 2260
rect 2605 2360 2645 2365
rect 2605 2330 2610 2360
rect 2640 2330 2645 2360
rect 2605 2290 2645 2330
rect 2605 2260 2610 2290
rect 2640 2260 2645 2290
rect 2605 2255 2645 2260
rect 2805 2360 2845 2365
rect 2805 2330 2810 2360
rect 2840 2330 2845 2360
rect 2805 2290 2845 2330
rect 2805 2260 2810 2290
rect 2840 2260 2845 2290
rect 2805 2255 2845 2260
rect 3005 2360 3045 2365
rect 3005 2330 3010 2360
rect 3040 2330 3045 2360
rect 3005 2290 3045 2330
rect 3005 2260 3010 2290
rect 3040 2260 3045 2290
rect 3005 2255 3045 2260
rect 3205 2360 3245 2365
rect 3205 2330 3210 2360
rect 3240 2330 3245 2360
rect 3205 2290 3245 2330
rect 3205 2260 3210 2290
rect 3240 2260 3245 2290
rect 3205 2255 3245 2260
rect 3405 2360 3445 2365
rect 3405 2330 3410 2360
rect 3440 2330 3445 2360
rect 3405 2290 3445 2330
rect 3405 2260 3410 2290
rect 3440 2260 3445 2290
rect 3405 2255 3445 2260
rect 3605 2360 3645 2365
rect 3605 2330 3610 2360
rect 3640 2330 3645 2360
rect 3605 2290 3645 2330
rect 3605 2260 3610 2290
rect 3640 2260 3645 2290
rect 3605 2255 3645 2260
rect 3805 2360 3845 2365
rect 3805 2330 3810 2360
rect 3840 2330 3845 2360
rect 3805 2290 3845 2330
rect 3805 2260 3810 2290
rect 3840 2260 3845 2290
rect 3805 2255 3845 2260
rect 4005 2360 4045 2365
rect 4005 2330 4010 2360
rect 4040 2330 4045 2360
rect 4005 2290 4045 2330
rect 4005 2260 4010 2290
rect 4040 2260 4045 2290
rect 4005 2255 4045 2260
rect 4205 2360 4245 2365
rect 4205 2330 4210 2360
rect 4240 2330 4245 2360
rect 4205 2290 4245 2330
rect 4205 2260 4210 2290
rect 4240 2260 4245 2290
rect 4205 2255 4245 2260
rect 4405 2360 4445 2365
rect 4405 2330 4410 2360
rect 4440 2330 4445 2360
rect 4405 2290 4445 2330
rect 4405 2260 4410 2290
rect 4440 2260 4445 2290
rect 4405 2255 4445 2260
rect 4605 2360 4645 2365
rect 4605 2330 4610 2360
rect 4640 2330 4645 2360
rect 4605 2290 4645 2330
rect 4605 2260 4610 2290
rect 4640 2260 4645 2290
rect 4605 2255 4645 2260
rect 4805 2360 4845 2365
rect 4805 2330 4810 2360
rect 4840 2330 4845 2360
rect 4805 2290 4845 2330
rect 4805 2260 4810 2290
rect 4840 2260 4845 2290
rect 4805 2255 4845 2260
rect 5005 2360 5045 2365
rect 5005 2330 5010 2360
rect 5040 2330 5045 2360
rect 5005 2290 5045 2330
rect 5005 2260 5010 2290
rect 5040 2260 5045 2290
rect 5005 2255 5045 2260
rect 5205 2360 5245 2365
rect 5205 2330 5210 2360
rect 5240 2330 5245 2360
rect 5205 2290 5245 2330
rect 5205 2260 5210 2290
rect 5240 2260 5245 2290
rect 5205 2255 5245 2260
rect 5405 2360 5445 2365
rect 5405 2330 5410 2360
rect 5440 2330 5445 2360
rect 5405 2290 5445 2330
rect 5405 2260 5410 2290
rect 5440 2260 5445 2290
rect 5405 2255 5445 2260
rect 5605 2360 5645 2365
rect 5605 2330 5610 2360
rect 5640 2330 5645 2360
rect 5605 2290 5645 2330
rect 5605 2260 5610 2290
rect 5640 2260 5645 2290
rect 5605 2255 5645 2260
rect 5805 2360 5845 2365
rect 5805 2330 5810 2360
rect 5840 2330 5845 2360
rect 5805 2290 5845 2330
rect 5805 2260 5810 2290
rect 5840 2260 5845 2290
rect 5805 2255 5845 2260
rect 6005 2360 6045 2365
rect 6005 2330 6010 2360
rect 6040 2330 6045 2360
rect 6005 2290 6045 2330
rect 6005 2260 6010 2290
rect 6040 2260 6045 2290
rect 6005 2255 6045 2260
rect 6205 2360 6245 2365
rect 6205 2330 6210 2360
rect 6240 2330 6245 2360
rect 6205 2290 6245 2330
rect 6205 2260 6210 2290
rect 6240 2260 6245 2290
rect 6205 2255 6245 2260
rect 6405 2360 6445 2365
rect 6405 2330 6410 2360
rect 6440 2330 6445 2360
rect 6405 2290 6445 2330
rect 6405 2260 6410 2290
rect 6440 2260 6445 2290
rect 6405 2255 6445 2260
rect -195 2175 -155 2180
rect -195 2145 -190 2175
rect -160 2145 -155 2175
rect -195 2105 -155 2145
rect -195 2075 -190 2105
rect -160 2075 -155 2105
rect -195 2070 -155 2075
rect 5 2175 45 2180
rect 5 2145 10 2175
rect 40 2145 45 2175
rect 5 2105 45 2145
rect 5 2075 10 2105
rect 40 2075 45 2105
rect 5 2070 45 2075
rect 205 2175 245 2180
rect 205 2145 210 2175
rect 240 2145 245 2175
rect 205 2105 245 2145
rect 205 2075 210 2105
rect 240 2075 245 2105
rect 205 2070 245 2075
rect 405 2175 445 2180
rect 405 2145 410 2175
rect 440 2145 445 2175
rect 405 2105 445 2145
rect 405 2075 410 2105
rect 440 2075 445 2105
rect 405 2070 445 2075
rect 605 2175 645 2180
rect 605 2145 610 2175
rect 640 2145 645 2175
rect 605 2105 645 2145
rect 605 2075 610 2105
rect 640 2075 645 2105
rect 605 2070 645 2075
rect 805 2175 845 2180
rect 805 2145 810 2175
rect 840 2145 845 2175
rect 805 2105 845 2145
rect 805 2075 810 2105
rect 840 2075 845 2105
rect 805 2070 845 2075
rect 1005 2175 1045 2180
rect 1005 2145 1010 2175
rect 1040 2145 1045 2175
rect 1005 2105 1045 2145
rect 1005 2075 1010 2105
rect 1040 2075 1045 2105
rect 1005 2070 1045 2075
rect 1205 2175 1245 2180
rect 1205 2145 1210 2175
rect 1240 2145 1245 2175
rect 1205 2105 1245 2145
rect 1205 2075 1210 2105
rect 1240 2075 1245 2105
rect 1205 2070 1245 2075
rect 1405 2175 1445 2180
rect 1405 2145 1410 2175
rect 1440 2145 1445 2175
rect 1405 2105 1445 2145
rect 1405 2075 1410 2105
rect 1440 2075 1445 2105
rect 1405 2070 1445 2075
rect 1605 2175 1645 2180
rect 1605 2145 1610 2175
rect 1640 2145 1645 2175
rect 1605 2105 1645 2145
rect 1605 2075 1610 2105
rect 1640 2075 1645 2105
rect 1605 2070 1645 2075
rect 1805 2175 1845 2180
rect 1805 2145 1810 2175
rect 1840 2145 1845 2175
rect 1805 2105 1845 2145
rect 1805 2075 1810 2105
rect 1840 2075 1845 2105
rect 1805 2070 1845 2075
rect 2005 2175 2045 2180
rect 2005 2145 2010 2175
rect 2040 2145 2045 2175
rect 2005 2105 2045 2145
rect 2005 2075 2010 2105
rect 2040 2075 2045 2105
rect 2005 2070 2045 2075
rect 2205 2175 2245 2180
rect 2205 2145 2210 2175
rect 2240 2145 2245 2175
rect 2205 2105 2245 2145
rect 2205 2075 2210 2105
rect 2240 2075 2245 2105
rect 2205 2070 2245 2075
rect 2405 2175 2445 2180
rect 2405 2145 2410 2175
rect 2440 2145 2445 2175
rect 2405 2105 2445 2145
rect 2405 2075 2410 2105
rect 2440 2075 2445 2105
rect 2405 2070 2445 2075
rect 2605 2175 2645 2180
rect 2605 2145 2610 2175
rect 2640 2145 2645 2175
rect 2605 2105 2645 2145
rect 2605 2075 2610 2105
rect 2640 2075 2645 2105
rect 2605 2070 2645 2075
rect 2805 2175 2845 2180
rect 2805 2145 2810 2175
rect 2840 2145 2845 2175
rect 2805 2105 2845 2145
rect 2805 2075 2810 2105
rect 2840 2075 2845 2105
rect 2805 2070 2845 2075
rect 3005 2175 3045 2180
rect 3005 2145 3010 2175
rect 3040 2145 3045 2175
rect 3005 2105 3045 2145
rect 3005 2075 3010 2105
rect 3040 2075 3045 2105
rect 3005 2070 3045 2075
rect 3205 2175 3245 2180
rect 3205 2145 3210 2175
rect 3240 2145 3245 2175
rect 3205 2105 3245 2145
rect 3205 2075 3210 2105
rect 3240 2075 3245 2105
rect 3205 2070 3245 2075
rect 3405 2175 3445 2180
rect 3405 2145 3410 2175
rect 3440 2145 3445 2175
rect 3405 2105 3445 2145
rect 3405 2075 3410 2105
rect 3440 2075 3445 2105
rect 3405 2070 3445 2075
rect 3605 2175 3645 2180
rect 3605 2145 3610 2175
rect 3640 2145 3645 2175
rect 3605 2105 3645 2145
rect 3605 2075 3610 2105
rect 3640 2075 3645 2105
rect 3605 2070 3645 2075
rect 3805 2175 3845 2180
rect 3805 2145 3810 2175
rect 3840 2145 3845 2175
rect 3805 2105 3845 2145
rect 3805 2075 3810 2105
rect 3840 2075 3845 2105
rect 3805 2070 3845 2075
rect 4005 2175 4045 2180
rect 4005 2145 4010 2175
rect 4040 2145 4045 2175
rect 4005 2105 4045 2145
rect 4005 2075 4010 2105
rect 4040 2075 4045 2105
rect 4005 2070 4045 2075
rect 4205 2175 4245 2180
rect 4205 2145 4210 2175
rect 4240 2145 4245 2175
rect 4205 2105 4245 2145
rect 4205 2075 4210 2105
rect 4240 2075 4245 2105
rect 4205 2070 4245 2075
rect 4405 2175 4445 2180
rect 4405 2145 4410 2175
rect 4440 2145 4445 2175
rect 4405 2105 4445 2145
rect 4405 2075 4410 2105
rect 4440 2075 4445 2105
rect 4405 2070 4445 2075
rect 4605 2175 4645 2180
rect 4605 2145 4610 2175
rect 4640 2145 4645 2175
rect 4605 2105 4645 2145
rect 4605 2075 4610 2105
rect 4640 2075 4645 2105
rect 4605 2070 4645 2075
rect 4805 2175 4845 2180
rect 4805 2145 4810 2175
rect 4840 2145 4845 2175
rect 4805 2105 4845 2145
rect 4805 2075 4810 2105
rect 4840 2075 4845 2105
rect 4805 2070 4845 2075
rect 5005 2175 5045 2180
rect 5005 2145 5010 2175
rect 5040 2145 5045 2175
rect 5005 2105 5045 2145
rect 5005 2075 5010 2105
rect 5040 2075 5045 2105
rect 5005 2070 5045 2075
rect 5205 2175 5245 2180
rect 5205 2145 5210 2175
rect 5240 2145 5245 2175
rect 5205 2105 5245 2145
rect 5205 2075 5210 2105
rect 5240 2075 5245 2105
rect 5205 2070 5245 2075
rect 5405 2175 5445 2180
rect 5405 2145 5410 2175
rect 5440 2145 5445 2175
rect 5405 2105 5445 2145
rect 5405 2075 5410 2105
rect 5440 2075 5445 2105
rect 5405 2070 5445 2075
rect 5605 2175 5645 2180
rect 5605 2145 5610 2175
rect 5640 2145 5645 2175
rect 5605 2105 5645 2145
rect 5605 2075 5610 2105
rect 5640 2075 5645 2105
rect 5605 2070 5645 2075
rect 5805 2175 5845 2180
rect 5805 2145 5810 2175
rect 5840 2145 5845 2175
rect 5805 2105 5845 2145
rect 5805 2075 5810 2105
rect 5840 2075 5845 2105
rect 5805 2070 5845 2075
rect 6005 2175 6045 2180
rect 6005 2145 6010 2175
rect 6040 2145 6045 2175
rect 6005 2105 6045 2145
rect 6005 2075 6010 2105
rect 6040 2075 6045 2105
rect 6005 2070 6045 2075
rect 6205 2175 6245 2180
rect 6205 2145 6210 2175
rect 6240 2145 6245 2175
rect 6205 2105 6245 2145
rect 6205 2075 6210 2105
rect 6240 2075 6245 2105
rect 6205 2070 6245 2075
rect 6405 2175 6445 2180
rect 6405 2145 6410 2175
rect 6440 2145 6445 2175
rect 6405 2105 6445 2145
rect 6405 2075 6410 2105
rect 6440 2075 6445 2105
rect 6405 2070 6445 2075
rect -195 1990 -155 1995
rect -195 1960 -190 1990
rect -160 1960 -155 1990
rect -195 1920 -155 1960
rect -195 1890 -190 1920
rect -160 1890 -155 1920
rect -195 1885 -155 1890
rect 5 1990 45 1995
rect 5 1960 10 1990
rect 40 1960 45 1990
rect 5 1920 45 1960
rect 5 1890 10 1920
rect 40 1890 45 1920
rect 5 1885 45 1890
rect 205 1990 245 1995
rect 205 1960 210 1990
rect 240 1960 245 1990
rect 205 1920 245 1960
rect 205 1890 210 1920
rect 240 1890 245 1920
rect 205 1885 245 1890
rect 405 1990 445 1995
rect 405 1960 410 1990
rect 440 1960 445 1990
rect 405 1920 445 1960
rect 405 1890 410 1920
rect 440 1890 445 1920
rect 405 1885 445 1890
rect 605 1990 645 1995
rect 605 1960 610 1990
rect 640 1960 645 1990
rect 605 1920 645 1960
rect 605 1890 610 1920
rect 640 1890 645 1920
rect 605 1885 645 1890
rect 805 1990 845 1995
rect 805 1960 810 1990
rect 840 1960 845 1990
rect 805 1920 845 1960
rect 805 1890 810 1920
rect 840 1890 845 1920
rect 805 1885 845 1890
rect 1005 1990 1045 1995
rect 1005 1960 1010 1990
rect 1040 1960 1045 1990
rect 1005 1920 1045 1960
rect 1005 1890 1010 1920
rect 1040 1890 1045 1920
rect 1005 1885 1045 1890
rect 1205 1990 1245 1995
rect 1205 1960 1210 1990
rect 1240 1960 1245 1990
rect 1205 1920 1245 1960
rect 1205 1890 1210 1920
rect 1240 1890 1245 1920
rect 1205 1885 1245 1890
rect 1405 1990 1445 1995
rect 1405 1960 1410 1990
rect 1440 1960 1445 1990
rect 1405 1920 1445 1960
rect 1405 1890 1410 1920
rect 1440 1890 1445 1920
rect 1405 1885 1445 1890
rect 1605 1990 1645 1995
rect 1605 1960 1610 1990
rect 1640 1960 1645 1990
rect 1605 1920 1645 1960
rect 1605 1890 1610 1920
rect 1640 1890 1645 1920
rect 1605 1885 1645 1890
rect 1805 1990 1845 1995
rect 1805 1960 1810 1990
rect 1840 1960 1845 1990
rect 1805 1920 1845 1960
rect 1805 1890 1810 1920
rect 1840 1890 1845 1920
rect 1805 1885 1845 1890
rect 2005 1990 2045 1995
rect 2005 1960 2010 1990
rect 2040 1960 2045 1990
rect 2005 1920 2045 1960
rect 2005 1890 2010 1920
rect 2040 1890 2045 1920
rect 2005 1885 2045 1890
rect 2205 1990 2245 1995
rect 2205 1960 2210 1990
rect 2240 1960 2245 1990
rect 2205 1920 2245 1960
rect 2205 1890 2210 1920
rect 2240 1890 2245 1920
rect 2205 1885 2245 1890
rect 2405 1990 2445 1995
rect 2405 1960 2410 1990
rect 2440 1960 2445 1990
rect 2405 1920 2445 1960
rect 2405 1890 2410 1920
rect 2440 1890 2445 1920
rect 2405 1885 2445 1890
rect 2605 1990 2645 1995
rect 2605 1960 2610 1990
rect 2640 1960 2645 1990
rect 2605 1920 2645 1960
rect 2605 1890 2610 1920
rect 2640 1890 2645 1920
rect 2605 1885 2645 1890
rect 2805 1990 2845 1995
rect 2805 1960 2810 1990
rect 2840 1960 2845 1990
rect 2805 1920 2845 1960
rect 2805 1890 2810 1920
rect 2840 1890 2845 1920
rect 2805 1885 2845 1890
rect 3005 1990 3045 1995
rect 3005 1960 3010 1990
rect 3040 1960 3045 1990
rect 3005 1920 3045 1960
rect 3005 1890 3010 1920
rect 3040 1890 3045 1920
rect 3005 1885 3045 1890
rect 3205 1990 3245 1995
rect 3205 1960 3210 1990
rect 3240 1960 3245 1990
rect 3205 1920 3245 1960
rect 3205 1890 3210 1920
rect 3240 1890 3245 1920
rect 3205 1885 3245 1890
rect 3405 1990 3445 1995
rect 3405 1960 3410 1990
rect 3440 1960 3445 1990
rect 3405 1920 3445 1960
rect 3405 1890 3410 1920
rect 3440 1890 3445 1920
rect 3405 1885 3445 1890
rect 3605 1990 3645 1995
rect 3605 1960 3610 1990
rect 3640 1960 3645 1990
rect 3605 1920 3645 1960
rect 3605 1890 3610 1920
rect 3640 1890 3645 1920
rect 3605 1885 3645 1890
rect 3805 1990 3845 1995
rect 3805 1960 3810 1990
rect 3840 1960 3845 1990
rect 3805 1920 3845 1960
rect 3805 1890 3810 1920
rect 3840 1890 3845 1920
rect 3805 1885 3845 1890
rect 4005 1990 4045 1995
rect 4005 1960 4010 1990
rect 4040 1960 4045 1990
rect 4005 1920 4045 1960
rect 4005 1890 4010 1920
rect 4040 1890 4045 1920
rect 4005 1885 4045 1890
rect 4205 1990 4245 1995
rect 4205 1960 4210 1990
rect 4240 1960 4245 1990
rect 4205 1920 4245 1960
rect 4205 1890 4210 1920
rect 4240 1890 4245 1920
rect 4205 1885 4245 1890
rect 4405 1990 4445 1995
rect 4405 1960 4410 1990
rect 4440 1960 4445 1990
rect 4405 1920 4445 1960
rect 4405 1890 4410 1920
rect 4440 1890 4445 1920
rect 4405 1885 4445 1890
rect 4605 1990 4645 1995
rect 4605 1960 4610 1990
rect 4640 1960 4645 1990
rect 4605 1920 4645 1960
rect 4605 1890 4610 1920
rect 4640 1890 4645 1920
rect 4605 1885 4645 1890
rect 4805 1990 4845 1995
rect 4805 1960 4810 1990
rect 4840 1960 4845 1990
rect 4805 1920 4845 1960
rect 4805 1890 4810 1920
rect 4840 1890 4845 1920
rect 4805 1885 4845 1890
rect 5005 1990 5045 1995
rect 5005 1960 5010 1990
rect 5040 1960 5045 1990
rect 5005 1920 5045 1960
rect 5005 1890 5010 1920
rect 5040 1890 5045 1920
rect 5005 1885 5045 1890
rect 5205 1990 5245 1995
rect 5205 1960 5210 1990
rect 5240 1960 5245 1990
rect 5205 1920 5245 1960
rect 5205 1890 5210 1920
rect 5240 1890 5245 1920
rect 5205 1885 5245 1890
rect 5405 1990 5445 1995
rect 5405 1960 5410 1990
rect 5440 1960 5445 1990
rect 5405 1920 5445 1960
rect 5405 1890 5410 1920
rect 5440 1890 5445 1920
rect 5405 1885 5445 1890
rect 5605 1990 5645 1995
rect 5605 1960 5610 1990
rect 5640 1960 5645 1990
rect 5605 1920 5645 1960
rect 5605 1890 5610 1920
rect 5640 1890 5645 1920
rect 5605 1885 5645 1890
rect 5805 1990 5845 1995
rect 5805 1960 5810 1990
rect 5840 1960 5845 1990
rect 5805 1920 5845 1960
rect 5805 1890 5810 1920
rect 5840 1890 5845 1920
rect 5805 1885 5845 1890
rect 6005 1990 6045 1995
rect 6005 1960 6010 1990
rect 6040 1960 6045 1990
rect 6005 1920 6045 1960
rect 6005 1890 6010 1920
rect 6040 1890 6045 1920
rect 6005 1885 6045 1890
rect 6205 1990 6245 1995
rect 6205 1960 6210 1990
rect 6240 1960 6245 1990
rect 6205 1920 6245 1960
rect 6205 1890 6210 1920
rect 6240 1890 6245 1920
rect 6205 1885 6245 1890
rect 6405 1990 6445 1995
rect 6405 1960 6410 1990
rect 6440 1960 6445 1990
rect 6405 1920 6445 1960
rect 6405 1890 6410 1920
rect 6440 1890 6445 1920
rect 6405 1885 6445 1890
rect -195 1805 -155 1810
rect -195 1775 -190 1805
rect -160 1775 -155 1805
rect -195 1735 -155 1775
rect -195 1705 -190 1735
rect -160 1705 -155 1735
rect -195 1700 -155 1705
rect 5 1805 45 1810
rect 5 1775 10 1805
rect 40 1775 45 1805
rect 5 1735 45 1775
rect 5 1705 10 1735
rect 40 1705 45 1735
rect 5 1700 45 1705
rect 205 1805 245 1810
rect 205 1775 210 1805
rect 240 1775 245 1805
rect 205 1735 245 1775
rect 205 1705 210 1735
rect 240 1705 245 1735
rect 205 1700 245 1705
rect 405 1805 445 1810
rect 405 1775 410 1805
rect 440 1775 445 1805
rect 405 1735 445 1775
rect 405 1705 410 1735
rect 440 1705 445 1735
rect 405 1700 445 1705
rect 605 1805 645 1810
rect 605 1775 610 1805
rect 640 1775 645 1805
rect 605 1735 645 1775
rect 605 1705 610 1735
rect 640 1705 645 1735
rect 605 1700 645 1705
rect 805 1805 845 1810
rect 805 1775 810 1805
rect 840 1775 845 1805
rect 805 1735 845 1775
rect 805 1705 810 1735
rect 840 1705 845 1735
rect 805 1700 845 1705
rect 1005 1805 1045 1810
rect 1005 1775 1010 1805
rect 1040 1775 1045 1805
rect 1005 1735 1045 1775
rect 1005 1705 1010 1735
rect 1040 1705 1045 1735
rect 1005 1700 1045 1705
rect 1205 1805 1245 1810
rect 1205 1775 1210 1805
rect 1240 1775 1245 1805
rect 1205 1735 1245 1775
rect 1205 1705 1210 1735
rect 1240 1705 1245 1735
rect 1205 1700 1245 1705
rect 1405 1805 1445 1810
rect 1405 1775 1410 1805
rect 1440 1775 1445 1805
rect 1405 1735 1445 1775
rect 1405 1705 1410 1735
rect 1440 1705 1445 1735
rect 1405 1700 1445 1705
rect 1605 1805 1645 1810
rect 1605 1775 1610 1805
rect 1640 1775 1645 1805
rect 1605 1735 1645 1775
rect 1605 1705 1610 1735
rect 1640 1705 1645 1735
rect 1605 1700 1645 1705
rect 1805 1805 1845 1810
rect 1805 1775 1810 1805
rect 1840 1775 1845 1805
rect 1805 1735 1845 1775
rect 1805 1705 1810 1735
rect 1840 1705 1845 1735
rect 1805 1700 1845 1705
rect 2005 1805 2045 1810
rect 2005 1775 2010 1805
rect 2040 1775 2045 1805
rect 2005 1735 2045 1775
rect 2005 1705 2010 1735
rect 2040 1705 2045 1735
rect 2005 1700 2045 1705
rect 2205 1805 2245 1810
rect 2205 1775 2210 1805
rect 2240 1775 2245 1805
rect 2205 1735 2245 1775
rect 2205 1705 2210 1735
rect 2240 1705 2245 1735
rect 2205 1700 2245 1705
rect 2405 1805 2445 1810
rect 2405 1775 2410 1805
rect 2440 1775 2445 1805
rect 2405 1735 2445 1775
rect 2405 1705 2410 1735
rect 2440 1705 2445 1735
rect 2405 1700 2445 1705
rect 2605 1805 2645 1810
rect 2605 1775 2610 1805
rect 2640 1775 2645 1805
rect 2605 1735 2645 1775
rect 2605 1705 2610 1735
rect 2640 1705 2645 1735
rect 2605 1700 2645 1705
rect 2805 1805 2845 1810
rect 2805 1775 2810 1805
rect 2840 1775 2845 1805
rect 2805 1735 2845 1775
rect 2805 1705 2810 1735
rect 2840 1705 2845 1735
rect 2805 1700 2845 1705
rect 3005 1805 3045 1810
rect 3005 1775 3010 1805
rect 3040 1775 3045 1805
rect 3005 1735 3045 1775
rect 3005 1705 3010 1735
rect 3040 1705 3045 1735
rect 3005 1700 3045 1705
rect 3205 1805 3245 1810
rect 3205 1775 3210 1805
rect 3240 1775 3245 1805
rect 3205 1735 3245 1775
rect 3205 1705 3210 1735
rect 3240 1705 3245 1735
rect 3205 1700 3245 1705
rect 3405 1805 3445 1810
rect 3405 1775 3410 1805
rect 3440 1775 3445 1805
rect 3405 1735 3445 1775
rect 3405 1705 3410 1735
rect 3440 1705 3445 1735
rect 3405 1700 3445 1705
rect 3605 1805 3645 1810
rect 3605 1775 3610 1805
rect 3640 1775 3645 1805
rect 3605 1735 3645 1775
rect 3605 1705 3610 1735
rect 3640 1705 3645 1735
rect 3605 1700 3645 1705
rect 3805 1805 3845 1810
rect 3805 1775 3810 1805
rect 3840 1775 3845 1805
rect 3805 1735 3845 1775
rect 3805 1705 3810 1735
rect 3840 1705 3845 1735
rect 3805 1700 3845 1705
rect 4005 1805 4045 1810
rect 4005 1775 4010 1805
rect 4040 1775 4045 1805
rect 4005 1735 4045 1775
rect 4005 1705 4010 1735
rect 4040 1705 4045 1735
rect 4005 1700 4045 1705
rect 4205 1805 4245 1810
rect 4205 1775 4210 1805
rect 4240 1775 4245 1805
rect 4205 1735 4245 1775
rect 4205 1705 4210 1735
rect 4240 1705 4245 1735
rect 4205 1700 4245 1705
rect 4405 1805 4445 1810
rect 4405 1775 4410 1805
rect 4440 1775 4445 1805
rect 4405 1735 4445 1775
rect 4405 1705 4410 1735
rect 4440 1705 4445 1735
rect 4405 1700 4445 1705
rect 4605 1805 4645 1810
rect 4605 1775 4610 1805
rect 4640 1775 4645 1805
rect 4605 1735 4645 1775
rect 4605 1705 4610 1735
rect 4640 1705 4645 1735
rect 4605 1700 4645 1705
rect 4805 1805 4845 1810
rect 4805 1775 4810 1805
rect 4840 1775 4845 1805
rect 4805 1735 4845 1775
rect 4805 1705 4810 1735
rect 4840 1705 4845 1735
rect 4805 1700 4845 1705
rect 5005 1805 5045 1810
rect 5005 1775 5010 1805
rect 5040 1775 5045 1805
rect 5005 1735 5045 1775
rect 5005 1705 5010 1735
rect 5040 1705 5045 1735
rect 5005 1700 5045 1705
rect 5205 1805 5245 1810
rect 5205 1775 5210 1805
rect 5240 1775 5245 1805
rect 5205 1735 5245 1775
rect 5205 1705 5210 1735
rect 5240 1705 5245 1735
rect 5205 1700 5245 1705
rect 5405 1805 5445 1810
rect 5405 1775 5410 1805
rect 5440 1775 5445 1805
rect 5405 1735 5445 1775
rect 5405 1705 5410 1735
rect 5440 1705 5445 1735
rect 5405 1700 5445 1705
rect 5605 1805 5645 1810
rect 5605 1775 5610 1805
rect 5640 1775 5645 1805
rect 5605 1735 5645 1775
rect 5605 1705 5610 1735
rect 5640 1705 5645 1735
rect 5605 1700 5645 1705
rect 5805 1805 5845 1810
rect 5805 1775 5810 1805
rect 5840 1775 5845 1805
rect 5805 1735 5845 1775
rect 5805 1705 5810 1735
rect 5840 1705 5845 1735
rect 5805 1700 5845 1705
rect 6005 1805 6045 1810
rect 6005 1775 6010 1805
rect 6040 1775 6045 1805
rect 6005 1735 6045 1775
rect 6005 1705 6010 1735
rect 6040 1705 6045 1735
rect 6005 1700 6045 1705
rect 6205 1805 6245 1810
rect 6205 1775 6210 1805
rect 6240 1775 6245 1805
rect 6205 1735 6245 1775
rect 6205 1705 6210 1735
rect 6240 1705 6245 1735
rect 6205 1700 6245 1705
rect 6405 1805 6445 1810
rect 6405 1775 6410 1805
rect 6440 1775 6445 1805
rect 6405 1735 6445 1775
rect 6405 1705 6410 1735
rect 6440 1705 6445 1735
rect 6405 1700 6445 1705
rect -195 1620 -155 1625
rect -195 1590 -190 1620
rect -160 1590 -155 1620
rect -195 1550 -155 1590
rect -195 1520 -190 1550
rect -160 1520 -155 1550
rect -195 1515 -155 1520
rect 5 1620 45 1625
rect 5 1590 10 1620
rect 40 1590 45 1620
rect 5 1550 45 1590
rect 5 1520 10 1550
rect 40 1520 45 1550
rect 5 1515 45 1520
rect 205 1620 245 1625
rect 205 1590 210 1620
rect 240 1590 245 1620
rect 205 1550 245 1590
rect 205 1520 210 1550
rect 240 1520 245 1550
rect 205 1515 245 1520
rect 405 1620 445 1625
rect 405 1590 410 1620
rect 440 1590 445 1620
rect 405 1550 445 1590
rect 405 1520 410 1550
rect 440 1520 445 1550
rect 405 1515 445 1520
rect 605 1620 645 1625
rect 605 1590 610 1620
rect 640 1590 645 1620
rect 605 1550 645 1590
rect 605 1520 610 1550
rect 640 1520 645 1550
rect 605 1515 645 1520
rect 805 1620 845 1625
rect 805 1590 810 1620
rect 840 1590 845 1620
rect 805 1550 845 1590
rect 805 1520 810 1550
rect 840 1520 845 1550
rect 805 1515 845 1520
rect 1005 1620 1045 1625
rect 1005 1590 1010 1620
rect 1040 1590 1045 1620
rect 1005 1550 1045 1590
rect 1005 1520 1010 1550
rect 1040 1520 1045 1550
rect 1005 1515 1045 1520
rect 1205 1620 1245 1625
rect 1205 1590 1210 1620
rect 1240 1590 1245 1620
rect 1205 1550 1245 1590
rect 1205 1520 1210 1550
rect 1240 1520 1245 1550
rect 1205 1515 1245 1520
rect 1405 1620 1445 1625
rect 1405 1590 1410 1620
rect 1440 1590 1445 1620
rect 1405 1550 1445 1590
rect 1405 1520 1410 1550
rect 1440 1520 1445 1550
rect 1405 1515 1445 1520
rect 1605 1620 1645 1625
rect 1605 1590 1610 1620
rect 1640 1590 1645 1620
rect 1605 1550 1645 1590
rect 1605 1520 1610 1550
rect 1640 1520 1645 1550
rect 1605 1515 1645 1520
rect 1805 1620 1845 1625
rect 1805 1590 1810 1620
rect 1840 1590 1845 1620
rect 1805 1550 1845 1590
rect 1805 1520 1810 1550
rect 1840 1520 1845 1550
rect 1805 1515 1845 1520
rect 2005 1620 2045 1625
rect 2005 1590 2010 1620
rect 2040 1590 2045 1620
rect 2005 1550 2045 1590
rect 2005 1520 2010 1550
rect 2040 1520 2045 1550
rect 2005 1515 2045 1520
rect 2205 1620 2245 1625
rect 2205 1590 2210 1620
rect 2240 1590 2245 1620
rect 2205 1550 2245 1590
rect 2205 1520 2210 1550
rect 2240 1520 2245 1550
rect 2205 1515 2245 1520
rect 2405 1620 2445 1625
rect 2405 1590 2410 1620
rect 2440 1590 2445 1620
rect 2405 1550 2445 1590
rect 2405 1520 2410 1550
rect 2440 1520 2445 1550
rect 2405 1515 2445 1520
rect 2605 1620 2645 1625
rect 2605 1590 2610 1620
rect 2640 1590 2645 1620
rect 2605 1550 2645 1590
rect 2605 1520 2610 1550
rect 2640 1520 2645 1550
rect 2605 1515 2645 1520
rect 2805 1620 2845 1625
rect 2805 1590 2810 1620
rect 2840 1590 2845 1620
rect 2805 1550 2845 1590
rect 2805 1520 2810 1550
rect 2840 1520 2845 1550
rect 2805 1515 2845 1520
rect 3005 1620 3045 1625
rect 3005 1590 3010 1620
rect 3040 1590 3045 1620
rect 3005 1550 3045 1590
rect 3005 1520 3010 1550
rect 3040 1520 3045 1550
rect 3005 1515 3045 1520
rect 3205 1620 3245 1625
rect 3205 1590 3210 1620
rect 3240 1590 3245 1620
rect 3205 1550 3245 1590
rect 3205 1520 3210 1550
rect 3240 1520 3245 1550
rect 3205 1515 3245 1520
rect 3405 1620 3445 1625
rect 3405 1590 3410 1620
rect 3440 1590 3445 1620
rect 3405 1550 3445 1590
rect 3405 1520 3410 1550
rect 3440 1520 3445 1550
rect 3405 1515 3445 1520
rect 3605 1620 3645 1625
rect 3605 1590 3610 1620
rect 3640 1590 3645 1620
rect 3605 1550 3645 1590
rect 3605 1520 3610 1550
rect 3640 1520 3645 1550
rect 3605 1515 3645 1520
rect 3805 1620 3845 1625
rect 3805 1590 3810 1620
rect 3840 1590 3845 1620
rect 3805 1550 3845 1590
rect 3805 1520 3810 1550
rect 3840 1520 3845 1550
rect 3805 1515 3845 1520
rect 4005 1620 4045 1625
rect 4005 1590 4010 1620
rect 4040 1590 4045 1620
rect 4005 1550 4045 1590
rect 4005 1520 4010 1550
rect 4040 1520 4045 1550
rect 4005 1515 4045 1520
rect 4205 1620 4245 1625
rect 4205 1590 4210 1620
rect 4240 1590 4245 1620
rect 4205 1550 4245 1590
rect 4205 1520 4210 1550
rect 4240 1520 4245 1550
rect 4205 1515 4245 1520
rect 4405 1620 4445 1625
rect 4405 1590 4410 1620
rect 4440 1590 4445 1620
rect 4405 1550 4445 1590
rect 4405 1520 4410 1550
rect 4440 1520 4445 1550
rect 4405 1515 4445 1520
rect 4605 1620 4645 1625
rect 4605 1590 4610 1620
rect 4640 1590 4645 1620
rect 4605 1550 4645 1590
rect 4605 1520 4610 1550
rect 4640 1520 4645 1550
rect 4605 1515 4645 1520
rect 4805 1620 4845 1625
rect 4805 1590 4810 1620
rect 4840 1590 4845 1620
rect 4805 1550 4845 1590
rect 4805 1520 4810 1550
rect 4840 1520 4845 1550
rect 4805 1515 4845 1520
rect 5005 1620 5045 1625
rect 5005 1590 5010 1620
rect 5040 1590 5045 1620
rect 5005 1550 5045 1590
rect 5005 1520 5010 1550
rect 5040 1520 5045 1550
rect 5005 1515 5045 1520
rect 5205 1620 5245 1625
rect 5205 1590 5210 1620
rect 5240 1590 5245 1620
rect 5205 1550 5245 1590
rect 5205 1520 5210 1550
rect 5240 1520 5245 1550
rect 5205 1515 5245 1520
rect 5405 1620 5445 1625
rect 5405 1590 5410 1620
rect 5440 1590 5445 1620
rect 5405 1550 5445 1590
rect 5405 1520 5410 1550
rect 5440 1520 5445 1550
rect 5405 1515 5445 1520
rect 5605 1620 5645 1625
rect 5605 1590 5610 1620
rect 5640 1590 5645 1620
rect 5605 1550 5645 1590
rect 5605 1520 5610 1550
rect 5640 1520 5645 1550
rect 5605 1515 5645 1520
rect 5805 1620 5845 1625
rect 5805 1590 5810 1620
rect 5840 1590 5845 1620
rect 5805 1550 5845 1590
rect 5805 1520 5810 1550
rect 5840 1520 5845 1550
rect 5805 1515 5845 1520
rect 6005 1620 6045 1625
rect 6005 1590 6010 1620
rect 6040 1590 6045 1620
rect 6005 1550 6045 1590
rect 6005 1520 6010 1550
rect 6040 1520 6045 1550
rect 6005 1515 6045 1520
rect 6205 1620 6245 1625
rect 6205 1590 6210 1620
rect 6240 1590 6245 1620
rect 6205 1550 6245 1590
rect 6205 1520 6210 1550
rect 6240 1520 6245 1550
rect 6205 1515 6245 1520
rect 6405 1620 6445 1625
rect 6405 1590 6410 1620
rect 6440 1590 6445 1620
rect 6405 1550 6445 1590
rect 6405 1520 6410 1550
rect 6440 1520 6445 1550
rect 6405 1515 6445 1520
rect -195 1435 -155 1440
rect -195 1405 -190 1435
rect -160 1405 -155 1435
rect -195 1365 -155 1405
rect -195 1335 -190 1365
rect -160 1335 -155 1365
rect -195 1330 -155 1335
rect 5 1435 45 1440
rect 5 1405 10 1435
rect 40 1405 45 1435
rect 5 1365 45 1405
rect 5 1335 10 1365
rect 40 1335 45 1365
rect 5 1330 45 1335
rect 205 1435 245 1440
rect 205 1405 210 1435
rect 240 1405 245 1435
rect 205 1365 245 1405
rect 205 1335 210 1365
rect 240 1335 245 1365
rect 205 1330 245 1335
rect 405 1435 445 1440
rect 405 1405 410 1435
rect 440 1405 445 1435
rect 405 1365 445 1405
rect 405 1335 410 1365
rect 440 1335 445 1365
rect 405 1330 445 1335
rect 605 1435 645 1440
rect 605 1405 610 1435
rect 640 1405 645 1435
rect 605 1365 645 1405
rect 605 1335 610 1365
rect 640 1335 645 1365
rect 605 1330 645 1335
rect 805 1435 845 1440
rect 805 1405 810 1435
rect 840 1405 845 1435
rect 805 1365 845 1405
rect 805 1335 810 1365
rect 840 1335 845 1365
rect 805 1330 845 1335
rect 1005 1435 1045 1440
rect 1005 1405 1010 1435
rect 1040 1405 1045 1435
rect 1005 1365 1045 1405
rect 1005 1335 1010 1365
rect 1040 1335 1045 1365
rect 1005 1330 1045 1335
rect 1205 1435 1245 1440
rect 1205 1405 1210 1435
rect 1240 1405 1245 1435
rect 1205 1365 1245 1405
rect 1205 1335 1210 1365
rect 1240 1335 1245 1365
rect 1205 1330 1245 1335
rect 1405 1435 1445 1440
rect 1405 1405 1410 1435
rect 1440 1405 1445 1435
rect 1405 1365 1445 1405
rect 1405 1335 1410 1365
rect 1440 1335 1445 1365
rect 1405 1330 1445 1335
rect 1605 1435 1645 1440
rect 1605 1405 1610 1435
rect 1640 1405 1645 1435
rect 1605 1365 1645 1405
rect 1605 1335 1610 1365
rect 1640 1335 1645 1365
rect 1605 1330 1645 1335
rect 1805 1435 1845 1440
rect 1805 1405 1810 1435
rect 1840 1405 1845 1435
rect 1805 1365 1845 1405
rect 1805 1335 1810 1365
rect 1840 1335 1845 1365
rect 1805 1330 1845 1335
rect 2005 1435 2045 1440
rect 2005 1405 2010 1435
rect 2040 1405 2045 1435
rect 2005 1365 2045 1405
rect 2005 1335 2010 1365
rect 2040 1335 2045 1365
rect 2005 1330 2045 1335
rect 2205 1435 2245 1440
rect 2205 1405 2210 1435
rect 2240 1405 2245 1435
rect 2205 1365 2245 1405
rect 2205 1335 2210 1365
rect 2240 1335 2245 1365
rect 2205 1330 2245 1335
rect 2405 1435 2445 1440
rect 2405 1405 2410 1435
rect 2440 1405 2445 1435
rect 2405 1365 2445 1405
rect 2405 1335 2410 1365
rect 2440 1335 2445 1365
rect 2405 1330 2445 1335
rect 2605 1435 2645 1440
rect 2605 1405 2610 1435
rect 2640 1405 2645 1435
rect 2605 1365 2645 1405
rect 2605 1335 2610 1365
rect 2640 1335 2645 1365
rect 2605 1330 2645 1335
rect 2805 1435 2845 1440
rect 2805 1405 2810 1435
rect 2840 1405 2845 1435
rect 2805 1365 2845 1405
rect 2805 1335 2810 1365
rect 2840 1335 2845 1365
rect 2805 1330 2845 1335
rect 3005 1435 3045 1440
rect 3005 1405 3010 1435
rect 3040 1405 3045 1435
rect 3005 1365 3045 1405
rect 3005 1335 3010 1365
rect 3040 1335 3045 1365
rect 3005 1330 3045 1335
rect 3205 1435 3245 1440
rect 3205 1405 3210 1435
rect 3240 1405 3245 1435
rect 3205 1365 3245 1405
rect 3205 1335 3210 1365
rect 3240 1335 3245 1365
rect 3205 1330 3245 1335
rect 3405 1435 3445 1440
rect 3405 1405 3410 1435
rect 3440 1405 3445 1435
rect 3405 1365 3445 1405
rect 3405 1335 3410 1365
rect 3440 1335 3445 1365
rect 3405 1330 3445 1335
rect 3605 1435 3645 1440
rect 3605 1405 3610 1435
rect 3640 1405 3645 1435
rect 3605 1365 3645 1405
rect 3605 1335 3610 1365
rect 3640 1335 3645 1365
rect 3605 1330 3645 1335
rect 3805 1435 3845 1440
rect 3805 1405 3810 1435
rect 3840 1405 3845 1435
rect 3805 1365 3845 1405
rect 3805 1335 3810 1365
rect 3840 1335 3845 1365
rect 3805 1330 3845 1335
rect 4005 1435 4045 1440
rect 4005 1405 4010 1435
rect 4040 1405 4045 1435
rect 4005 1365 4045 1405
rect 4005 1335 4010 1365
rect 4040 1335 4045 1365
rect 4005 1330 4045 1335
rect 4205 1435 4245 1440
rect 4205 1405 4210 1435
rect 4240 1405 4245 1435
rect 4205 1365 4245 1405
rect 4205 1335 4210 1365
rect 4240 1335 4245 1365
rect 4205 1330 4245 1335
rect 4405 1435 4445 1440
rect 4405 1405 4410 1435
rect 4440 1405 4445 1435
rect 4405 1365 4445 1405
rect 4405 1335 4410 1365
rect 4440 1335 4445 1365
rect 4405 1330 4445 1335
rect 4605 1435 4645 1440
rect 4605 1405 4610 1435
rect 4640 1405 4645 1435
rect 4605 1365 4645 1405
rect 4605 1335 4610 1365
rect 4640 1335 4645 1365
rect 4605 1330 4645 1335
rect 4805 1435 4845 1440
rect 4805 1405 4810 1435
rect 4840 1405 4845 1435
rect 4805 1365 4845 1405
rect 4805 1335 4810 1365
rect 4840 1335 4845 1365
rect 4805 1330 4845 1335
rect 5005 1435 5045 1440
rect 5005 1405 5010 1435
rect 5040 1405 5045 1435
rect 5005 1365 5045 1405
rect 5005 1335 5010 1365
rect 5040 1335 5045 1365
rect 5005 1330 5045 1335
rect 5205 1435 5245 1440
rect 5205 1405 5210 1435
rect 5240 1405 5245 1435
rect 5205 1365 5245 1405
rect 5205 1335 5210 1365
rect 5240 1335 5245 1365
rect 5205 1330 5245 1335
rect 5405 1435 5445 1440
rect 5405 1405 5410 1435
rect 5440 1405 5445 1435
rect 5405 1365 5445 1405
rect 5405 1335 5410 1365
rect 5440 1335 5445 1365
rect 5405 1330 5445 1335
rect 5605 1435 5645 1440
rect 5605 1405 5610 1435
rect 5640 1405 5645 1435
rect 5605 1365 5645 1405
rect 5605 1335 5610 1365
rect 5640 1335 5645 1365
rect 5605 1330 5645 1335
rect 5805 1435 5845 1440
rect 5805 1405 5810 1435
rect 5840 1405 5845 1435
rect 5805 1365 5845 1405
rect 5805 1335 5810 1365
rect 5840 1335 5845 1365
rect 5805 1330 5845 1335
rect 6005 1435 6045 1440
rect 6005 1405 6010 1435
rect 6040 1405 6045 1435
rect 6005 1365 6045 1405
rect 6005 1335 6010 1365
rect 6040 1335 6045 1365
rect 6005 1330 6045 1335
rect 6205 1435 6245 1440
rect 6205 1405 6210 1435
rect 6240 1405 6245 1435
rect 6205 1365 6245 1405
rect 6205 1335 6210 1365
rect 6240 1335 6245 1365
rect 6205 1330 6245 1335
rect 6405 1435 6445 1440
rect 6405 1405 6410 1435
rect 6440 1405 6445 1435
rect 6405 1365 6445 1405
rect 6405 1335 6410 1365
rect 6440 1335 6445 1365
rect 6405 1330 6445 1335
rect -195 1250 -155 1255
rect -195 1220 -190 1250
rect -160 1220 -155 1250
rect -195 1180 -155 1220
rect -195 1150 -190 1180
rect -160 1150 -155 1180
rect -195 1145 -155 1150
rect 5 1250 45 1255
rect 5 1220 10 1250
rect 40 1220 45 1250
rect 5 1180 45 1220
rect 5 1150 10 1180
rect 40 1150 45 1180
rect 5 1145 45 1150
rect 205 1250 245 1255
rect 205 1220 210 1250
rect 240 1220 245 1250
rect 205 1180 245 1220
rect 205 1150 210 1180
rect 240 1150 245 1180
rect 205 1145 245 1150
rect 405 1250 445 1255
rect 405 1220 410 1250
rect 440 1220 445 1250
rect 405 1180 445 1220
rect 405 1150 410 1180
rect 440 1150 445 1180
rect 405 1145 445 1150
rect 605 1250 645 1255
rect 605 1220 610 1250
rect 640 1220 645 1250
rect 605 1180 645 1220
rect 605 1150 610 1180
rect 640 1150 645 1180
rect 605 1145 645 1150
rect 805 1250 845 1255
rect 805 1220 810 1250
rect 840 1220 845 1250
rect 805 1180 845 1220
rect 805 1150 810 1180
rect 840 1150 845 1180
rect 805 1145 845 1150
rect 1005 1250 1045 1255
rect 1005 1220 1010 1250
rect 1040 1220 1045 1250
rect 1005 1180 1045 1220
rect 1005 1150 1010 1180
rect 1040 1150 1045 1180
rect 1005 1145 1045 1150
rect 1205 1250 1245 1255
rect 1205 1220 1210 1250
rect 1240 1220 1245 1250
rect 1205 1180 1245 1220
rect 1205 1150 1210 1180
rect 1240 1150 1245 1180
rect 1205 1145 1245 1150
rect 1405 1250 1445 1255
rect 1405 1220 1410 1250
rect 1440 1220 1445 1250
rect 1405 1180 1445 1220
rect 1405 1150 1410 1180
rect 1440 1150 1445 1180
rect 1405 1145 1445 1150
rect 1605 1250 1645 1255
rect 1605 1220 1610 1250
rect 1640 1220 1645 1250
rect 1605 1180 1645 1220
rect 1605 1150 1610 1180
rect 1640 1150 1645 1180
rect 1605 1145 1645 1150
rect 1805 1250 1845 1255
rect 1805 1220 1810 1250
rect 1840 1220 1845 1250
rect 1805 1180 1845 1220
rect 1805 1150 1810 1180
rect 1840 1150 1845 1180
rect 1805 1145 1845 1150
rect 2005 1250 2045 1255
rect 2005 1220 2010 1250
rect 2040 1220 2045 1250
rect 2005 1180 2045 1220
rect 2005 1150 2010 1180
rect 2040 1150 2045 1180
rect 2005 1145 2045 1150
rect 2205 1250 2245 1255
rect 2205 1220 2210 1250
rect 2240 1220 2245 1250
rect 2205 1180 2245 1220
rect 2205 1150 2210 1180
rect 2240 1150 2245 1180
rect 2205 1145 2245 1150
rect 2405 1250 2445 1255
rect 2405 1220 2410 1250
rect 2440 1220 2445 1250
rect 2405 1180 2445 1220
rect 2405 1150 2410 1180
rect 2440 1150 2445 1180
rect 2405 1145 2445 1150
rect 2605 1250 2645 1255
rect 2605 1220 2610 1250
rect 2640 1220 2645 1250
rect 2605 1180 2645 1220
rect 2605 1150 2610 1180
rect 2640 1150 2645 1180
rect 2605 1145 2645 1150
rect 2805 1250 2845 1255
rect 2805 1220 2810 1250
rect 2840 1220 2845 1250
rect 2805 1180 2845 1220
rect 2805 1150 2810 1180
rect 2840 1150 2845 1180
rect 2805 1145 2845 1150
rect 3005 1250 3045 1255
rect 3005 1220 3010 1250
rect 3040 1220 3045 1250
rect 3005 1180 3045 1220
rect 3005 1150 3010 1180
rect 3040 1150 3045 1180
rect 3005 1145 3045 1150
rect 3205 1250 3245 1255
rect 3205 1220 3210 1250
rect 3240 1220 3245 1250
rect 3205 1180 3245 1220
rect 3205 1150 3210 1180
rect 3240 1150 3245 1180
rect 3205 1145 3245 1150
rect 3405 1250 3445 1255
rect 3405 1220 3410 1250
rect 3440 1220 3445 1250
rect 3405 1180 3445 1220
rect 3405 1150 3410 1180
rect 3440 1150 3445 1180
rect 3405 1145 3445 1150
rect 3605 1250 3645 1255
rect 3605 1220 3610 1250
rect 3640 1220 3645 1250
rect 3605 1180 3645 1220
rect 3605 1150 3610 1180
rect 3640 1150 3645 1180
rect 3605 1145 3645 1150
rect 3805 1250 3845 1255
rect 3805 1220 3810 1250
rect 3840 1220 3845 1250
rect 3805 1180 3845 1220
rect 3805 1150 3810 1180
rect 3840 1150 3845 1180
rect 3805 1145 3845 1150
rect 4005 1250 4045 1255
rect 4005 1220 4010 1250
rect 4040 1220 4045 1250
rect 4005 1180 4045 1220
rect 4005 1150 4010 1180
rect 4040 1150 4045 1180
rect 4005 1145 4045 1150
rect 4205 1250 4245 1255
rect 4205 1220 4210 1250
rect 4240 1220 4245 1250
rect 4205 1180 4245 1220
rect 4205 1150 4210 1180
rect 4240 1150 4245 1180
rect 4205 1145 4245 1150
rect 4405 1250 4445 1255
rect 4405 1220 4410 1250
rect 4440 1220 4445 1250
rect 4405 1180 4445 1220
rect 4405 1150 4410 1180
rect 4440 1150 4445 1180
rect 4405 1145 4445 1150
rect 4605 1250 4645 1255
rect 4605 1220 4610 1250
rect 4640 1220 4645 1250
rect 4605 1180 4645 1220
rect 4605 1150 4610 1180
rect 4640 1150 4645 1180
rect 4605 1145 4645 1150
rect 4805 1250 4845 1255
rect 4805 1220 4810 1250
rect 4840 1220 4845 1250
rect 4805 1180 4845 1220
rect 4805 1150 4810 1180
rect 4840 1150 4845 1180
rect 4805 1145 4845 1150
rect 5005 1250 5045 1255
rect 5005 1220 5010 1250
rect 5040 1220 5045 1250
rect 5005 1180 5045 1220
rect 5005 1150 5010 1180
rect 5040 1150 5045 1180
rect 5005 1145 5045 1150
rect 5205 1250 5245 1255
rect 5205 1220 5210 1250
rect 5240 1220 5245 1250
rect 5205 1180 5245 1220
rect 5205 1150 5210 1180
rect 5240 1150 5245 1180
rect 5205 1145 5245 1150
rect 5405 1250 5445 1255
rect 5405 1220 5410 1250
rect 5440 1220 5445 1250
rect 5405 1180 5445 1220
rect 5405 1150 5410 1180
rect 5440 1150 5445 1180
rect 5405 1145 5445 1150
rect 5605 1250 5645 1255
rect 5605 1220 5610 1250
rect 5640 1220 5645 1250
rect 5605 1180 5645 1220
rect 5605 1150 5610 1180
rect 5640 1150 5645 1180
rect 5605 1145 5645 1150
rect 5805 1250 5845 1255
rect 5805 1220 5810 1250
rect 5840 1220 5845 1250
rect 5805 1180 5845 1220
rect 5805 1150 5810 1180
rect 5840 1150 5845 1180
rect 5805 1145 5845 1150
rect 6005 1250 6045 1255
rect 6005 1220 6010 1250
rect 6040 1220 6045 1250
rect 6005 1180 6045 1220
rect 6005 1150 6010 1180
rect 6040 1150 6045 1180
rect 6005 1145 6045 1150
rect 6205 1250 6245 1255
rect 6205 1220 6210 1250
rect 6240 1220 6245 1250
rect 6205 1180 6245 1220
rect 6205 1150 6210 1180
rect 6240 1150 6245 1180
rect 6205 1145 6245 1150
rect 6405 1250 6445 1255
rect 6405 1220 6410 1250
rect 6440 1220 6445 1250
rect 6405 1180 6445 1220
rect 6405 1150 6410 1180
rect 6440 1150 6445 1180
rect 6405 1145 6445 1150
rect -195 1065 -155 1070
rect -195 1035 -190 1065
rect -160 1035 -155 1065
rect -195 995 -155 1035
rect -195 965 -190 995
rect -160 965 -155 995
rect -195 960 -155 965
rect 5 1065 45 1070
rect 5 1035 10 1065
rect 40 1035 45 1065
rect 5 995 45 1035
rect 5 965 10 995
rect 40 965 45 995
rect 5 960 45 965
rect 205 1065 245 1070
rect 205 1035 210 1065
rect 240 1035 245 1065
rect 205 995 245 1035
rect 205 965 210 995
rect 240 965 245 995
rect 205 960 245 965
rect 405 1065 445 1070
rect 405 1035 410 1065
rect 440 1035 445 1065
rect 405 995 445 1035
rect 405 965 410 995
rect 440 965 445 995
rect 405 960 445 965
rect 605 1065 645 1070
rect 605 1035 610 1065
rect 640 1035 645 1065
rect 605 995 645 1035
rect 605 965 610 995
rect 640 965 645 995
rect 605 960 645 965
rect 805 1065 845 1070
rect 805 1035 810 1065
rect 840 1035 845 1065
rect 805 995 845 1035
rect 805 965 810 995
rect 840 965 845 995
rect 805 960 845 965
rect 1005 1065 1045 1070
rect 1005 1035 1010 1065
rect 1040 1035 1045 1065
rect 1005 995 1045 1035
rect 1005 965 1010 995
rect 1040 965 1045 995
rect 1005 960 1045 965
rect 1205 1065 1245 1070
rect 1205 1035 1210 1065
rect 1240 1035 1245 1065
rect 1205 995 1245 1035
rect 1205 965 1210 995
rect 1240 965 1245 995
rect 1205 960 1245 965
rect 1405 1065 1445 1070
rect 1405 1035 1410 1065
rect 1440 1035 1445 1065
rect 1405 995 1445 1035
rect 1405 965 1410 995
rect 1440 965 1445 995
rect 1405 960 1445 965
rect 1605 1065 1645 1070
rect 1605 1035 1610 1065
rect 1640 1035 1645 1065
rect 1605 995 1645 1035
rect 1605 965 1610 995
rect 1640 965 1645 995
rect 1605 960 1645 965
rect 1805 1065 1845 1070
rect 1805 1035 1810 1065
rect 1840 1035 1845 1065
rect 1805 995 1845 1035
rect 1805 965 1810 995
rect 1840 965 1845 995
rect 1805 960 1845 965
rect 2005 1065 2045 1070
rect 2005 1035 2010 1065
rect 2040 1035 2045 1065
rect 2005 995 2045 1035
rect 2005 965 2010 995
rect 2040 965 2045 995
rect 2005 960 2045 965
rect 2205 1065 2245 1070
rect 2205 1035 2210 1065
rect 2240 1035 2245 1065
rect 2205 995 2245 1035
rect 2205 965 2210 995
rect 2240 965 2245 995
rect 2205 960 2245 965
rect 2405 1065 2445 1070
rect 2405 1035 2410 1065
rect 2440 1035 2445 1065
rect 2405 995 2445 1035
rect 2405 965 2410 995
rect 2440 965 2445 995
rect 2405 960 2445 965
rect 2605 1065 2645 1070
rect 2605 1035 2610 1065
rect 2640 1035 2645 1065
rect 2605 995 2645 1035
rect 2605 965 2610 995
rect 2640 965 2645 995
rect 2605 960 2645 965
rect 2805 1065 2845 1070
rect 2805 1035 2810 1065
rect 2840 1035 2845 1065
rect 2805 995 2845 1035
rect 2805 965 2810 995
rect 2840 965 2845 995
rect 2805 960 2845 965
rect 3005 1065 3045 1070
rect 3005 1035 3010 1065
rect 3040 1035 3045 1065
rect 3005 995 3045 1035
rect 3005 965 3010 995
rect 3040 965 3045 995
rect 3005 960 3045 965
rect 3205 1065 3245 1070
rect 3205 1035 3210 1065
rect 3240 1035 3245 1065
rect 3205 995 3245 1035
rect 3205 965 3210 995
rect 3240 965 3245 995
rect 3205 960 3245 965
rect 3405 1065 3445 1070
rect 3405 1035 3410 1065
rect 3440 1035 3445 1065
rect 3405 995 3445 1035
rect 3405 965 3410 995
rect 3440 965 3445 995
rect 3405 960 3445 965
rect 3605 1065 3645 1070
rect 3605 1035 3610 1065
rect 3640 1035 3645 1065
rect 3605 995 3645 1035
rect 3605 965 3610 995
rect 3640 965 3645 995
rect 3605 960 3645 965
rect 3805 1065 3845 1070
rect 3805 1035 3810 1065
rect 3840 1035 3845 1065
rect 3805 995 3845 1035
rect 3805 965 3810 995
rect 3840 965 3845 995
rect 3805 960 3845 965
rect 4005 1065 4045 1070
rect 4005 1035 4010 1065
rect 4040 1035 4045 1065
rect 4005 995 4045 1035
rect 4005 965 4010 995
rect 4040 965 4045 995
rect 4005 960 4045 965
rect 4205 1065 4245 1070
rect 4205 1035 4210 1065
rect 4240 1035 4245 1065
rect 4205 995 4245 1035
rect 4205 965 4210 995
rect 4240 965 4245 995
rect 4205 960 4245 965
rect 4405 1065 4445 1070
rect 4405 1035 4410 1065
rect 4440 1035 4445 1065
rect 4405 995 4445 1035
rect 4405 965 4410 995
rect 4440 965 4445 995
rect 4405 960 4445 965
rect 4605 1065 4645 1070
rect 4605 1035 4610 1065
rect 4640 1035 4645 1065
rect 4605 995 4645 1035
rect 4605 965 4610 995
rect 4640 965 4645 995
rect 4605 960 4645 965
rect 4805 1065 4845 1070
rect 4805 1035 4810 1065
rect 4840 1035 4845 1065
rect 4805 995 4845 1035
rect 4805 965 4810 995
rect 4840 965 4845 995
rect 4805 960 4845 965
rect 5005 1065 5045 1070
rect 5005 1035 5010 1065
rect 5040 1035 5045 1065
rect 5005 995 5045 1035
rect 5005 965 5010 995
rect 5040 965 5045 995
rect 5005 960 5045 965
rect 5205 1065 5245 1070
rect 5205 1035 5210 1065
rect 5240 1035 5245 1065
rect 5205 995 5245 1035
rect 5205 965 5210 995
rect 5240 965 5245 995
rect 5205 960 5245 965
rect 5405 1065 5445 1070
rect 5405 1035 5410 1065
rect 5440 1035 5445 1065
rect 5405 995 5445 1035
rect 5405 965 5410 995
rect 5440 965 5445 995
rect 5405 960 5445 965
rect 5605 1065 5645 1070
rect 5605 1035 5610 1065
rect 5640 1035 5645 1065
rect 5605 995 5645 1035
rect 5605 965 5610 995
rect 5640 965 5645 995
rect 5605 960 5645 965
rect 5805 1065 5845 1070
rect 5805 1035 5810 1065
rect 5840 1035 5845 1065
rect 5805 995 5845 1035
rect 5805 965 5810 995
rect 5840 965 5845 995
rect 5805 960 5845 965
rect 6005 1065 6045 1070
rect 6005 1035 6010 1065
rect 6040 1035 6045 1065
rect 6005 995 6045 1035
rect 6005 965 6010 995
rect 6040 965 6045 995
rect 6005 960 6045 965
rect 6205 1065 6245 1070
rect 6205 1035 6210 1065
rect 6240 1035 6245 1065
rect 6205 995 6245 1035
rect 6205 965 6210 995
rect 6240 965 6245 995
rect 6205 960 6245 965
rect 6405 1065 6445 1070
rect 6405 1035 6410 1065
rect 6440 1035 6445 1065
rect 6405 995 6445 1035
rect 6405 965 6410 995
rect 6440 965 6445 995
rect 6405 960 6445 965
rect -195 880 -155 885
rect -195 850 -190 880
rect -160 850 -155 880
rect -195 810 -155 850
rect -195 780 -190 810
rect -160 780 -155 810
rect -195 775 -155 780
rect 5 880 45 885
rect 5 850 10 880
rect 40 850 45 880
rect 5 810 45 850
rect 5 780 10 810
rect 40 780 45 810
rect 5 775 45 780
rect 205 880 245 885
rect 205 850 210 880
rect 240 850 245 880
rect 205 810 245 850
rect 205 780 210 810
rect 240 780 245 810
rect 205 775 245 780
rect 405 880 445 885
rect 405 850 410 880
rect 440 850 445 880
rect 405 810 445 850
rect 405 780 410 810
rect 440 780 445 810
rect 405 775 445 780
rect 605 880 645 885
rect 605 850 610 880
rect 640 850 645 880
rect 605 810 645 850
rect 605 780 610 810
rect 640 780 645 810
rect 605 775 645 780
rect 805 880 845 885
rect 805 850 810 880
rect 840 850 845 880
rect 805 810 845 850
rect 805 780 810 810
rect 840 780 845 810
rect 805 775 845 780
rect 1005 880 1045 885
rect 1005 850 1010 880
rect 1040 850 1045 880
rect 1005 810 1045 850
rect 1005 780 1010 810
rect 1040 780 1045 810
rect 1005 775 1045 780
rect 1205 880 1245 885
rect 1205 850 1210 880
rect 1240 850 1245 880
rect 1205 810 1245 850
rect 1205 780 1210 810
rect 1240 780 1245 810
rect 1205 775 1245 780
rect 1405 880 1445 885
rect 1405 850 1410 880
rect 1440 850 1445 880
rect 1405 810 1445 850
rect 1405 780 1410 810
rect 1440 780 1445 810
rect 1405 775 1445 780
rect 1605 880 1645 885
rect 1605 850 1610 880
rect 1640 850 1645 880
rect 1605 810 1645 850
rect 1605 780 1610 810
rect 1640 780 1645 810
rect 1605 775 1645 780
rect 1805 880 1845 885
rect 1805 850 1810 880
rect 1840 850 1845 880
rect 1805 810 1845 850
rect 1805 780 1810 810
rect 1840 780 1845 810
rect 1805 775 1845 780
rect 2005 880 2045 885
rect 2005 850 2010 880
rect 2040 850 2045 880
rect 2005 810 2045 850
rect 2005 780 2010 810
rect 2040 780 2045 810
rect 2005 775 2045 780
rect 2205 880 2245 885
rect 2205 850 2210 880
rect 2240 850 2245 880
rect 2205 810 2245 850
rect 2205 780 2210 810
rect 2240 780 2245 810
rect 2205 775 2245 780
rect 2405 880 2445 885
rect 2405 850 2410 880
rect 2440 850 2445 880
rect 2405 810 2445 850
rect 2405 780 2410 810
rect 2440 780 2445 810
rect 2405 775 2445 780
rect 2605 880 2645 885
rect 2605 850 2610 880
rect 2640 850 2645 880
rect 2605 810 2645 850
rect 2605 780 2610 810
rect 2640 780 2645 810
rect 2605 775 2645 780
rect 2805 880 2845 885
rect 2805 850 2810 880
rect 2840 850 2845 880
rect 2805 810 2845 850
rect 2805 780 2810 810
rect 2840 780 2845 810
rect 2805 775 2845 780
rect 3005 880 3045 885
rect 3005 850 3010 880
rect 3040 850 3045 880
rect 3005 810 3045 850
rect 3005 780 3010 810
rect 3040 780 3045 810
rect 3005 775 3045 780
rect 3205 880 3245 885
rect 3205 850 3210 880
rect 3240 850 3245 880
rect 3205 810 3245 850
rect 3205 780 3210 810
rect 3240 780 3245 810
rect 3205 775 3245 780
rect 3405 880 3445 885
rect 3405 850 3410 880
rect 3440 850 3445 880
rect 3405 810 3445 850
rect 3405 780 3410 810
rect 3440 780 3445 810
rect 3405 775 3445 780
rect 3605 880 3645 885
rect 3605 850 3610 880
rect 3640 850 3645 880
rect 3605 810 3645 850
rect 3605 780 3610 810
rect 3640 780 3645 810
rect 3605 775 3645 780
rect 3805 880 3845 885
rect 3805 850 3810 880
rect 3840 850 3845 880
rect 3805 810 3845 850
rect 3805 780 3810 810
rect 3840 780 3845 810
rect 3805 775 3845 780
rect 4005 880 4045 885
rect 4005 850 4010 880
rect 4040 850 4045 880
rect 4005 810 4045 850
rect 4005 780 4010 810
rect 4040 780 4045 810
rect 4005 775 4045 780
rect 4205 880 4245 885
rect 4205 850 4210 880
rect 4240 850 4245 880
rect 4205 810 4245 850
rect 4205 780 4210 810
rect 4240 780 4245 810
rect 4205 775 4245 780
rect 4405 880 4445 885
rect 4405 850 4410 880
rect 4440 850 4445 880
rect 4405 810 4445 850
rect 4405 780 4410 810
rect 4440 780 4445 810
rect 4405 775 4445 780
rect 4605 880 4645 885
rect 4605 850 4610 880
rect 4640 850 4645 880
rect 4605 810 4645 850
rect 4605 780 4610 810
rect 4640 780 4645 810
rect 4605 775 4645 780
rect 4805 880 4845 885
rect 4805 850 4810 880
rect 4840 850 4845 880
rect 4805 810 4845 850
rect 4805 780 4810 810
rect 4840 780 4845 810
rect 4805 775 4845 780
rect 5005 880 5045 885
rect 5005 850 5010 880
rect 5040 850 5045 880
rect 5005 810 5045 850
rect 5005 780 5010 810
rect 5040 780 5045 810
rect 5005 775 5045 780
rect 5205 880 5245 885
rect 5205 850 5210 880
rect 5240 850 5245 880
rect 5205 810 5245 850
rect 5205 780 5210 810
rect 5240 780 5245 810
rect 5205 775 5245 780
rect 5405 880 5445 885
rect 5405 850 5410 880
rect 5440 850 5445 880
rect 5405 810 5445 850
rect 5405 780 5410 810
rect 5440 780 5445 810
rect 5405 775 5445 780
rect 5605 880 5645 885
rect 5605 850 5610 880
rect 5640 850 5645 880
rect 5605 810 5645 850
rect 5605 780 5610 810
rect 5640 780 5645 810
rect 5605 775 5645 780
rect 5805 880 5845 885
rect 5805 850 5810 880
rect 5840 850 5845 880
rect 5805 810 5845 850
rect 5805 780 5810 810
rect 5840 780 5845 810
rect 5805 775 5845 780
rect 6005 880 6045 885
rect 6005 850 6010 880
rect 6040 850 6045 880
rect 6005 810 6045 850
rect 6005 780 6010 810
rect 6040 780 6045 810
rect 6005 775 6045 780
rect 6205 880 6245 885
rect 6205 850 6210 880
rect 6240 850 6245 880
rect 6205 810 6245 850
rect 6205 780 6210 810
rect 6240 780 6245 810
rect 6205 775 6245 780
rect 6405 880 6445 885
rect 6405 850 6410 880
rect 6440 850 6445 880
rect 6405 810 6445 850
rect 6405 780 6410 810
rect 6440 780 6445 810
rect 6405 775 6445 780
rect -195 695 -155 700
rect -195 665 -190 695
rect -160 665 -155 695
rect -195 625 -155 665
rect -195 595 -190 625
rect -160 595 -155 625
rect -195 590 -155 595
rect 5 695 45 700
rect 5 665 10 695
rect 40 665 45 695
rect 5 625 45 665
rect 5 595 10 625
rect 40 595 45 625
rect 5 590 45 595
rect 205 695 245 700
rect 205 665 210 695
rect 240 665 245 695
rect 205 625 245 665
rect 205 595 210 625
rect 240 595 245 625
rect 205 590 245 595
rect 405 695 445 700
rect 405 665 410 695
rect 440 665 445 695
rect 405 625 445 665
rect 405 595 410 625
rect 440 595 445 625
rect 405 590 445 595
rect 605 695 645 700
rect 605 665 610 695
rect 640 665 645 695
rect 605 625 645 665
rect 605 595 610 625
rect 640 595 645 625
rect 605 590 645 595
rect 805 695 845 700
rect 805 665 810 695
rect 840 665 845 695
rect 805 625 845 665
rect 805 595 810 625
rect 840 595 845 625
rect 805 590 845 595
rect 1005 695 1045 700
rect 1005 665 1010 695
rect 1040 665 1045 695
rect 1005 625 1045 665
rect 1005 595 1010 625
rect 1040 595 1045 625
rect 1005 590 1045 595
rect 1205 695 1245 700
rect 1205 665 1210 695
rect 1240 665 1245 695
rect 1205 625 1245 665
rect 1205 595 1210 625
rect 1240 595 1245 625
rect 1205 590 1245 595
rect 1405 695 1445 700
rect 1405 665 1410 695
rect 1440 665 1445 695
rect 1405 625 1445 665
rect 1405 595 1410 625
rect 1440 595 1445 625
rect 1405 590 1445 595
rect 1605 695 1645 700
rect 1605 665 1610 695
rect 1640 665 1645 695
rect 1605 625 1645 665
rect 1605 595 1610 625
rect 1640 595 1645 625
rect 1605 590 1645 595
rect 1805 695 1845 700
rect 1805 665 1810 695
rect 1840 665 1845 695
rect 1805 625 1845 665
rect 1805 595 1810 625
rect 1840 595 1845 625
rect 1805 590 1845 595
rect 2005 695 2045 700
rect 2005 665 2010 695
rect 2040 665 2045 695
rect 2005 625 2045 665
rect 2005 595 2010 625
rect 2040 595 2045 625
rect 2005 590 2045 595
rect 2205 695 2245 700
rect 2205 665 2210 695
rect 2240 665 2245 695
rect 2205 625 2245 665
rect 2205 595 2210 625
rect 2240 595 2245 625
rect 2205 590 2245 595
rect 2405 695 2445 700
rect 2405 665 2410 695
rect 2440 665 2445 695
rect 2405 625 2445 665
rect 2405 595 2410 625
rect 2440 595 2445 625
rect 2405 590 2445 595
rect 2605 695 2645 700
rect 2605 665 2610 695
rect 2640 665 2645 695
rect 2605 625 2645 665
rect 2605 595 2610 625
rect 2640 595 2645 625
rect 2605 590 2645 595
rect 2805 695 2845 700
rect 2805 665 2810 695
rect 2840 665 2845 695
rect 2805 625 2845 665
rect 2805 595 2810 625
rect 2840 595 2845 625
rect 2805 590 2845 595
rect 3005 695 3045 700
rect 3005 665 3010 695
rect 3040 665 3045 695
rect 3005 625 3045 665
rect 3005 595 3010 625
rect 3040 595 3045 625
rect 3005 590 3045 595
rect 3205 695 3245 700
rect 3205 665 3210 695
rect 3240 665 3245 695
rect 3205 625 3245 665
rect 3205 595 3210 625
rect 3240 595 3245 625
rect 3205 590 3245 595
rect 3405 695 3445 700
rect 3405 665 3410 695
rect 3440 665 3445 695
rect 3405 625 3445 665
rect 3405 595 3410 625
rect 3440 595 3445 625
rect 3405 590 3445 595
rect 3605 695 3645 700
rect 3605 665 3610 695
rect 3640 665 3645 695
rect 3605 625 3645 665
rect 3605 595 3610 625
rect 3640 595 3645 625
rect 3605 590 3645 595
rect 3805 695 3845 700
rect 3805 665 3810 695
rect 3840 665 3845 695
rect 3805 625 3845 665
rect 3805 595 3810 625
rect 3840 595 3845 625
rect 3805 590 3845 595
rect 4005 695 4045 700
rect 4005 665 4010 695
rect 4040 665 4045 695
rect 4005 625 4045 665
rect 4005 595 4010 625
rect 4040 595 4045 625
rect 4005 590 4045 595
rect 4205 695 4245 700
rect 4205 665 4210 695
rect 4240 665 4245 695
rect 4205 625 4245 665
rect 4205 595 4210 625
rect 4240 595 4245 625
rect 4205 590 4245 595
rect 4405 695 4445 700
rect 4405 665 4410 695
rect 4440 665 4445 695
rect 4405 625 4445 665
rect 4405 595 4410 625
rect 4440 595 4445 625
rect 4405 590 4445 595
rect 4605 695 4645 700
rect 4605 665 4610 695
rect 4640 665 4645 695
rect 4605 625 4645 665
rect 4605 595 4610 625
rect 4640 595 4645 625
rect 4605 590 4645 595
rect 4805 695 4845 700
rect 4805 665 4810 695
rect 4840 665 4845 695
rect 4805 625 4845 665
rect 4805 595 4810 625
rect 4840 595 4845 625
rect 4805 590 4845 595
rect 5005 695 5045 700
rect 5005 665 5010 695
rect 5040 665 5045 695
rect 5005 625 5045 665
rect 5005 595 5010 625
rect 5040 595 5045 625
rect 5005 590 5045 595
rect 5205 695 5245 700
rect 5205 665 5210 695
rect 5240 665 5245 695
rect 5205 625 5245 665
rect 5205 595 5210 625
rect 5240 595 5245 625
rect 5205 590 5245 595
rect 5405 695 5445 700
rect 5405 665 5410 695
rect 5440 665 5445 695
rect 5405 625 5445 665
rect 5405 595 5410 625
rect 5440 595 5445 625
rect 5405 590 5445 595
rect 5605 695 5645 700
rect 5605 665 5610 695
rect 5640 665 5645 695
rect 5605 625 5645 665
rect 5605 595 5610 625
rect 5640 595 5645 625
rect 5605 590 5645 595
rect 5805 695 5845 700
rect 5805 665 5810 695
rect 5840 665 5845 695
rect 5805 625 5845 665
rect 5805 595 5810 625
rect 5840 595 5845 625
rect 5805 590 5845 595
rect 6005 695 6045 700
rect 6005 665 6010 695
rect 6040 665 6045 695
rect 6005 625 6045 665
rect 6005 595 6010 625
rect 6040 595 6045 625
rect 6005 590 6045 595
rect 6205 695 6245 700
rect 6205 665 6210 695
rect 6240 665 6245 695
rect 6205 625 6245 665
rect 6205 595 6210 625
rect 6240 595 6245 625
rect 6205 590 6245 595
rect 6405 695 6445 700
rect 6405 665 6410 695
rect 6440 665 6445 695
rect 6405 625 6445 665
rect 6405 595 6410 625
rect 6440 595 6445 625
rect 6405 590 6445 595
rect -195 510 -155 515
rect -195 480 -190 510
rect -160 480 -155 510
rect -195 440 -155 480
rect -195 410 -190 440
rect -160 410 -155 440
rect -195 405 -155 410
rect 5 510 45 515
rect 5 480 10 510
rect 40 480 45 510
rect 5 440 45 480
rect 5 410 10 440
rect 40 410 45 440
rect 5 405 45 410
rect 205 510 245 515
rect 205 480 210 510
rect 240 480 245 510
rect 205 440 245 480
rect 205 410 210 440
rect 240 410 245 440
rect 205 405 245 410
rect 405 510 445 515
rect 405 480 410 510
rect 440 480 445 510
rect 405 440 445 480
rect 405 410 410 440
rect 440 410 445 440
rect 405 405 445 410
rect 605 510 645 515
rect 605 480 610 510
rect 640 480 645 510
rect 605 440 645 480
rect 605 410 610 440
rect 640 410 645 440
rect 605 405 645 410
rect 805 510 845 515
rect 805 480 810 510
rect 840 480 845 510
rect 805 440 845 480
rect 805 410 810 440
rect 840 410 845 440
rect 805 405 845 410
rect 1005 510 1045 515
rect 1005 480 1010 510
rect 1040 480 1045 510
rect 1005 440 1045 480
rect 1005 410 1010 440
rect 1040 410 1045 440
rect 1005 405 1045 410
rect 1205 510 1245 515
rect 1205 480 1210 510
rect 1240 480 1245 510
rect 1205 440 1245 480
rect 1205 410 1210 440
rect 1240 410 1245 440
rect 1205 405 1245 410
rect 1405 510 1445 515
rect 1405 480 1410 510
rect 1440 480 1445 510
rect 1405 440 1445 480
rect 1405 410 1410 440
rect 1440 410 1445 440
rect 1405 405 1445 410
rect 1605 510 1645 515
rect 1605 480 1610 510
rect 1640 480 1645 510
rect 1605 440 1645 480
rect 1605 410 1610 440
rect 1640 410 1645 440
rect 1605 405 1645 410
rect 1805 510 1845 515
rect 1805 480 1810 510
rect 1840 480 1845 510
rect 1805 440 1845 480
rect 1805 410 1810 440
rect 1840 410 1845 440
rect 1805 405 1845 410
rect 2005 510 2045 515
rect 2005 480 2010 510
rect 2040 480 2045 510
rect 2005 440 2045 480
rect 2005 410 2010 440
rect 2040 410 2045 440
rect 2005 405 2045 410
rect 2205 510 2245 515
rect 2205 480 2210 510
rect 2240 480 2245 510
rect 2205 440 2245 480
rect 2205 410 2210 440
rect 2240 410 2245 440
rect 2205 405 2245 410
rect 2405 510 2445 515
rect 2405 480 2410 510
rect 2440 480 2445 510
rect 2405 440 2445 480
rect 2405 410 2410 440
rect 2440 410 2445 440
rect 2405 405 2445 410
rect 2605 510 2645 515
rect 2605 480 2610 510
rect 2640 480 2645 510
rect 2605 440 2645 480
rect 2605 410 2610 440
rect 2640 410 2645 440
rect 2605 405 2645 410
rect 2805 510 2845 515
rect 2805 480 2810 510
rect 2840 480 2845 510
rect 2805 440 2845 480
rect 2805 410 2810 440
rect 2840 410 2845 440
rect 2805 405 2845 410
rect 3005 510 3045 515
rect 3005 480 3010 510
rect 3040 480 3045 510
rect 3005 440 3045 480
rect 3005 410 3010 440
rect 3040 410 3045 440
rect 3005 405 3045 410
rect 3205 510 3245 515
rect 3205 480 3210 510
rect 3240 480 3245 510
rect 3205 440 3245 480
rect 3205 410 3210 440
rect 3240 410 3245 440
rect 3205 405 3245 410
rect 3405 510 3445 515
rect 3405 480 3410 510
rect 3440 480 3445 510
rect 3405 440 3445 480
rect 3405 410 3410 440
rect 3440 410 3445 440
rect 3405 405 3445 410
rect 3605 510 3645 515
rect 3605 480 3610 510
rect 3640 480 3645 510
rect 3605 440 3645 480
rect 3605 410 3610 440
rect 3640 410 3645 440
rect 3605 405 3645 410
rect 3805 510 3845 515
rect 3805 480 3810 510
rect 3840 480 3845 510
rect 3805 440 3845 480
rect 3805 410 3810 440
rect 3840 410 3845 440
rect 3805 405 3845 410
rect 4005 510 4045 515
rect 4005 480 4010 510
rect 4040 480 4045 510
rect 4005 440 4045 480
rect 4005 410 4010 440
rect 4040 410 4045 440
rect 4005 405 4045 410
rect 4205 510 4245 515
rect 4205 480 4210 510
rect 4240 480 4245 510
rect 4205 440 4245 480
rect 4205 410 4210 440
rect 4240 410 4245 440
rect 4205 405 4245 410
rect 4405 510 4445 515
rect 4405 480 4410 510
rect 4440 480 4445 510
rect 4405 440 4445 480
rect 4405 410 4410 440
rect 4440 410 4445 440
rect 4405 405 4445 410
rect 4605 510 4645 515
rect 4605 480 4610 510
rect 4640 480 4645 510
rect 4605 440 4645 480
rect 4605 410 4610 440
rect 4640 410 4645 440
rect 4605 405 4645 410
rect 4805 510 4845 515
rect 4805 480 4810 510
rect 4840 480 4845 510
rect 4805 440 4845 480
rect 4805 410 4810 440
rect 4840 410 4845 440
rect 4805 405 4845 410
rect 5005 510 5045 515
rect 5005 480 5010 510
rect 5040 480 5045 510
rect 5005 440 5045 480
rect 5005 410 5010 440
rect 5040 410 5045 440
rect 5005 405 5045 410
rect 5205 510 5245 515
rect 5205 480 5210 510
rect 5240 480 5245 510
rect 5205 440 5245 480
rect 5205 410 5210 440
rect 5240 410 5245 440
rect 5205 405 5245 410
rect 5405 510 5445 515
rect 5405 480 5410 510
rect 5440 480 5445 510
rect 5405 440 5445 480
rect 5405 410 5410 440
rect 5440 410 5445 440
rect 5405 405 5445 410
rect 5605 510 5645 515
rect 5605 480 5610 510
rect 5640 480 5645 510
rect 5605 440 5645 480
rect 5605 410 5610 440
rect 5640 410 5645 440
rect 5605 405 5645 410
rect 5805 510 5845 515
rect 5805 480 5810 510
rect 5840 480 5845 510
rect 5805 440 5845 480
rect 5805 410 5810 440
rect 5840 410 5845 440
rect 5805 405 5845 410
rect 6005 510 6045 515
rect 6005 480 6010 510
rect 6040 480 6045 510
rect 6005 440 6045 480
rect 6005 410 6010 440
rect 6040 410 6045 440
rect 6005 405 6045 410
rect 6205 510 6245 515
rect 6205 480 6210 510
rect 6240 480 6245 510
rect 6205 440 6245 480
rect 6205 410 6210 440
rect 6240 410 6245 440
rect 6205 405 6245 410
rect 6405 510 6445 515
rect 6405 480 6410 510
rect 6440 480 6445 510
rect 6405 440 6445 480
rect 6405 410 6410 440
rect 6440 410 6445 440
rect 6405 405 6445 410
rect -195 325 -155 330
rect -195 295 -190 325
rect -160 295 -155 325
rect -195 255 -155 295
rect -195 225 -190 255
rect -160 225 -155 255
rect -195 220 -155 225
rect 5 325 45 330
rect 5 295 10 325
rect 40 295 45 325
rect 5 255 45 295
rect 5 225 10 255
rect 40 225 45 255
rect 5 220 45 225
rect 205 325 245 330
rect 205 295 210 325
rect 240 295 245 325
rect 205 255 245 295
rect 205 225 210 255
rect 240 225 245 255
rect 205 220 245 225
rect 405 325 445 330
rect 405 295 410 325
rect 440 295 445 325
rect 405 255 445 295
rect 405 225 410 255
rect 440 225 445 255
rect 405 220 445 225
rect 605 325 645 330
rect 605 295 610 325
rect 640 295 645 325
rect 605 255 645 295
rect 605 225 610 255
rect 640 225 645 255
rect 605 220 645 225
rect 805 325 845 330
rect 805 295 810 325
rect 840 295 845 325
rect 805 255 845 295
rect 805 225 810 255
rect 840 225 845 255
rect 805 220 845 225
rect 1005 325 1045 330
rect 1005 295 1010 325
rect 1040 295 1045 325
rect 1005 255 1045 295
rect 1005 225 1010 255
rect 1040 225 1045 255
rect 1005 220 1045 225
rect 1205 325 1245 330
rect 1205 295 1210 325
rect 1240 295 1245 325
rect 1205 255 1245 295
rect 1205 225 1210 255
rect 1240 225 1245 255
rect 1205 220 1245 225
rect 1405 325 1445 330
rect 1405 295 1410 325
rect 1440 295 1445 325
rect 1405 255 1445 295
rect 1405 225 1410 255
rect 1440 225 1445 255
rect 1405 220 1445 225
rect 1605 325 1645 330
rect 1605 295 1610 325
rect 1640 295 1645 325
rect 1605 255 1645 295
rect 1605 225 1610 255
rect 1640 225 1645 255
rect 1605 220 1645 225
rect 1805 325 1845 330
rect 1805 295 1810 325
rect 1840 295 1845 325
rect 1805 255 1845 295
rect 1805 225 1810 255
rect 1840 225 1845 255
rect 1805 220 1845 225
rect 2005 325 2045 330
rect 2005 295 2010 325
rect 2040 295 2045 325
rect 2005 255 2045 295
rect 2005 225 2010 255
rect 2040 225 2045 255
rect 2005 220 2045 225
rect 2205 325 2245 330
rect 2205 295 2210 325
rect 2240 295 2245 325
rect 2205 255 2245 295
rect 2205 225 2210 255
rect 2240 225 2245 255
rect 2205 220 2245 225
rect 2405 325 2445 330
rect 2405 295 2410 325
rect 2440 295 2445 325
rect 2405 255 2445 295
rect 2405 225 2410 255
rect 2440 225 2445 255
rect 2405 220 2445 225
rect 2605 325 2645 330
rect 2605 295 2610 325
rect 2640 295 2645 325
rect 2605 255 2645 295
rect 2605 225 2610 255
rect 2640 225 2645 255
rect 2605 220 2645 225
rect 2805 325 2845 330
rect 2805 295 2810 325
rect 2840 295 2845 325
rect 2805 255 2845 295
rect 2805 225 2810 255
rect 2840 225 2845 255
rect 2805 220 2845 225
rect 3005 325 3045 330
rect 3005 295 3010 325
rect 3040 295 3045 325
rect 3005 255 3045 295
rect 3005 225 3010 255
rect 3040 225 3045 255
rect 3005 220 3045 225
rect 3205 325 3245 330
rect 3205 295 3210 325
rect 3240 295 3245 325
rect 3205 255 3245 295
rect 3205 225 3210 255
rect 3240 225 3245 255
rect 3205 220 3245 225
rect 3405 325 3445 330
rect 3405 295 3410 325
rect 3440 295 3445 325
rect 3405 255 3445 295
rect 3405 225 3410 255
rect 3440 225 3445 255
rect 3405 220 3445 225
rect 3605 325 3645 330
rect 3605 295 3610 325
rect 3640 295 3645 325
rect 3605 255 3645 295
rect 3605 225 3610 255
rect 3640 225 3645 255
rect 3605 220 3645 225
rect 3805 325 3845 330
rect 3805 295 3810 325
rect 3840 295 3845 325
rect 3805 255 3845 295
rect 3805 225 3810 255
rect 3840 225 3845 255
rect 3805 220 3845 225
rect 4005 325 4045 330
rect 4005 295 4010 325
rect 4040 295 4045 325
rect 4005 255 4045 295
rect 4005 225 4010 255
rect 4040 225 4045 255
rect 4005 220 4045 225
rect 4205 325 4245 330
rect 4205 295 4210 325
rect 4240 295 4245 325
rect 4205 255 4245 295
rect 4205 225 4210 255
rect 4240 225 4245 255
rect 4205 220 4245 225
rect 4405 325 4445 330
rect 4405 295 4410 325
rect 4440 295 4445 325
rect 4405 255 4445 295
rect 4405 225 4410 255
rect 4440 225 4445 255
rect 4405 220 4445 225
rect 4605 325 4645 330
rect 4605 295 4610 325
rect 4640 295 4645 325
rect 4605 255 4645 295
rect 4605 225 4610 255
rect 4640 225 4645 255
rect 4605 220 4645 225
rect 4805 325 4845 330
rect 4805 295 4810 325
rect 4840 295 4845 325
rect 4805 255 4845 295
rect 4805 225 4810 255
rect 4840 225 4845 255
rect 4805 220 4845 225
rect 5005 325 5045 330
rect 5005 295 5010 325
rect 5040 295 5045 325
rect 5005 255 5045 295
rect 5005 225 5010 255
rect 5040 225 5045 255
rect 5005 220 5045 225
rect 5205 325 5245 330
rect 5205 295 5210 325
rect 5240 295 5245 325
rect 5205 255 5245 295
rect 5205 225 5210 255
rect 5240 225 5245 255
rect 5205 220 5245 225
rect 5405 325 5445 330
rect 5405 295 5410 325
rect 5440 295 5445 325
rect 5405 255 5445 295
rect 5405 225 5410 255
rect 5440 225 5445 255
rect 5405 220 5445 225
rect 5605 325 5645 330
rect 5605 295 5610 325
rect 5640 295 5645 325
rect 5605 255 5645 295
rect 5605 225 5610 255
rect 5640 225 5645 255
rect 5605 220 5645 225
rect 5805 325 5845 330
rect 5805 295 5810 325
rect 5840 295 5845 325
rect 5805 255 5845 295
rect 5805 225 5810 255
rect 5840 225 5845 255
rect 5805 220 5845 225
rect 6005 325 6045 330
rect 6005 295 6010 325
rect 6040 295 6045 325
rect 6005 255 6045 295
rect 6005 225 6010 255
rect 6040 225 6045 255
rect 6005 220 6045 225
rect 6205 325 6245 330
rect 6205 295 6210 325
rect 6240 295 6245 325
rect 6205 255 6245 295
rect 6205 225 6210 255
rect 6240 225 6245 255
rect 6205 220 6245 225
rect 6405 325 6445 330
rect 6405 295 6410 325
rect 6440 295 6445 325
rect 6405 255 6445 295
rect 6405 225 6410 255
rect 6440 225 6445 255
rect 6405 220 6445 225
rect -195 140 -155 145
rect -195 110 -190 140
rect -160 110 -155 140
rect -195 70 -155 110
rect -195 40 -190 70
rect -160 40 -155 70
rect -195 35 -155 40
rect 5 140 45 145
rect 5 110 10 140
rect 40 110 45 140
rect 5 70 45 110
rect 5 40 10 70
rect 40 40 45 70
rect 5 35 45 40
rect 205 140 245 145
rect 205 110 210 140
rect 240 110 245 140
rect 205 70 245 110
rect 205 40 210 70
rect 240 40 245 70
rect 205 35 245 40
rect 405 140 445 145
rect 405 110 410 140
rect 440 110 445 140
rect 405 70 445 110
rect 405 40 410 70
rect 440 40 445 70
rect 405 35 445 40
rect 605 140 645 145
rect 605 110 610 140
rect 640 110 645 140
rect 605 70 645 110
rect 605 40 610 70
rect 640 40 645 70
rect 605 35 645 40
rect 805 140 845 145
rect 805 110 810 140
rect 840 110 845 140
rect 805 70 845 110
rect 805 40 810 70
rect 840 40 845 70
rect 805 35 845 40
rect 1005 140 1045 145
rect 1005 110 1010 140
rect 1040 110 1045 140
rect 1005 70 1045 110
rect 1005 40 1010 70
rect 1040 40 1045 70
rect 1005 35 1045 40
rect 1205 140 1245 145
rect 1205 110 1210 140
rect 1240 110 1245 140
rect 1205 70 1245 110
rect 1205 40 1210 70
rect 1240 40 1245 70
rect 1205 35 1245 40
rect 1405 140 1445 145
rect 1405 110 1410 140
rect 1440 110 1445 140
rect 1405 70 1445 110
rect 1405 40 1410 70
rect 1440 40 1445 70
rect 1405 35 1445 40
rect 1605 140 1645 145
rect 1605 110 1610 140
rect 1640 110 1645 140
rect 1605 70 1645 110
rect 1605 40 1610 70
rect 1640 40 1645 70
rect 1605 35 1645 40
rect 1805 140 1845 145
rect 1805 110 1810 140
rect 1840 110 1845 140
rect 1805 70 1845 110
rect 1805 40 1810 70
rect 1840 40 1845 70
rect 1805 35 1845 40
rect 2005 140 2045 145
rect 2005 110 2010 140
rect 2040 110 2045 140
rect 2005 70 2045 110
rect 2005 40 2010 70
rect 2040 40 2045 70
rect 2005 35 2045 40
rect 2205 140 2245 145
rect 2205 110 2210 140
rect 2240 110 2245 140
rect 2205 70 2245 110
rect 2205 40 2210 70
rect 2240 40 2245 70
rect 2205 35 2245 40
rect 2405 140 2445 145
rect 2405 110 2410 140
rect 2440 110 2445 140
rect 2405 70 2445 110
rect 2405 40 2410 70
rect 2440 40 2445 70
rect 2405 35 2445 40
rect 2605 140 2645 145
rect 2605 110 2610 140
rect 2640 110 2645 140
rect 2605 70 2645 110
rect 2605 40 2610 70
rect 2640 40 2645 70
rect 2605 35 2645 40
rect 2805 140 2845 145
rect 2805 110 2810 140
rect 2840 110 2845 140
rect 2805 70 2845 110
rect 2805 40 2810 70
rect 2840 40 2845 70
rect 2805 35 2845 40
rect 3005 140 3045 145
rect 3005 110 3010 140
rect 3040 110 3045 140
rect 3005 70 3045 110
rect 3005 40 3010 70
rect 3040 40 3045 70
rect 3005 35 3045 40
rect 3205 140 3245 145
rect 3205 110 3210 140
rect 3240 110 3245 140
rect 3205 70 3245 110
rect 3205 40 3210 70
rect 3240 40 3245 70
rect 3205 35 3245 40
rect 3405 140 3445 145
rect 3405 110 3410 140
rect 3440 110 3445 140
rect 3405 70 3445 110
rect 3405 40 3410 70
rect 3440 40 3445 70
rect 3405 35 3445 40
rect 3605 140 3645 145
rect 3605 110 3610 140
rect 3640 110 3645 140
rect 3605 70 3645 110
rect 3605 40 3610 70
rect 3640 40 3645 70
rect 3605 35 3645 40
rect 3805 140 3845 145
rect 3805 110 3810 140
rect 3840 110 3845 140
rect 3805 70 3845 110
rect 3805 40 3810 70
rect 3840 40 3845 70
rect 3805 35 3845 40
rect 4005 140 4045 145
rect 4005 110 4010 140
rect 4040 110 4045 140
rect 4005 70 4045 110
rect 4005 40 4010 70
rect 4040 40 4045 70
rect 4005 35 4045 40
rect 4205 140 4245 145
rect 4205 110 4210 140
rect 4240 110 4245 140
rect 4205 70 4245 110
rect 4205 40 4210 70
rect 4240 40 4245 70
rect 4205 35 4245 40
rect 4405 140 4445 145
rect 4405 110 4410 140
rect 4440 110 4445 140
rect 4405 70 4445 110
rect 4405 40 4410 70
rect 4440 40 4445 70
rect 4405 35 4445 40
rect 4605 140 4645 145
rect 4605 110 4610 140
rect 4640 110 4645 140
rect 4605 70 4645 110
rect 4605 40 4610 70
rect 4640 40 4645 70
rect 4605 35 4645 40
rect 4805 140 4845 145
rect 4805 110 4810 140
rect 4840 110 4845 140
rect 4805 70 4845 110
rect 4805 40 4810 70
rect 4840 40 4845 70
rect 4805 35 4845 40
rect 5005 140 5045 145
rect 5005 110 5010 140
rect 5040 110 5045 140
rect 5005 70 5045 110
rect 5005 40 5010 70
rect 5040 40 5045 70
rect 5005 35 5045 40
rect 5205 140 5245 145
rect 5205 110 5210 140
rect 5240 110 5245 140
rect 5205 70 5245 110
rect 5205 40 5210 70
rect 5240 40 5245 70
rect 5205 35 5245 40
rect 5405 140 5445 145
rect 5405 110 5410 140
rect 5440 110 5445 140
rect 5405 70 5445 110
rect 5405 40 5410 70
rect 5440 40 5445 70
rect 5405 35 5445 40
rect 5605 140 5645 145
rect 5605 110 5610 140
rect 5640 110 5645 140
rect 5605 70 5645 110
rect 5605 40 5610 70
rect 5640 40 5645 70
rect 5605 35 5645 40
rect 5805 140 5845 145
rect 5805 110 5810 140
rect 5840 110 5845 140
rect 5805 70 5845 110
rect 5805 40 5810 70
rect 5840 40 5845 70
rect 5805 35 5845 40
rect 6005 140 6045 145
rect 6005 110 6010 140
rect 6040 110 6045 140
rect 6005 70 6045 110
rect 6005 40 6010 70
rect 6040 40 6045 70
rect 6005 35 6045 40
rect 6205 140 6245 145
rect 6205 110 6210 140
rect 6240 110 6245 140
rect 6205 70 6245 110
rect 6205 40 6210 70
rect 6240 40 6245 70
rect 6205 35 6245 40
rect 6405 140 6445 145
rect 6405 110 6410 140
rect 6440 110 6445 140
rect 6405 70 6445 110
rect 6405 40 6410 70
rect 6440 40 6445 70
rect 6405 35 6445 40
rect -195 -45 -155 -40
rect -195 -75 -190 -45
rect -160 -75 -155 -45
rect -195 -115 -155 -75
rect -195 -145 -190 -115
rect -160 -145 -155 -115
rect -195 -150 -155 -145
rect 5 -45 45 -40
rect 5 -75 10 -45
rect 40 -75 45 -45
rect 5 -115 45 -75
rect 5 -145 10 -115
rect 40 -145 45 -115
rect 5 -150 45 -145
rect 205 -45 245 -40
rect 205 -75 210 -45
rect 240 -75 245 -45
rect 205 -115 245 -75
rect 205 -145 210 -115
rect 240 -145 245 -115
rect 205 -150 245 -145
rect 405 -45 445 -40
rect 405 -75 410 -45
rect 440 -75 445 -45
rect 405 -115 445 -75
rect 405 -145 410 -115
rect 440 -145 445 -115
rect 405 -150 445 -145
rect 605 -45 645 -40
rect 605 -75 610 -45
rect 640 -75 645 -45
rect 605 -115 645 -75
rect 605 -145 610 -115
rect 640 -145 645 -115
rect 605 -150 645 -145
rect 805 -45 845 -40
rect 805 -75 810 -45
rect 840 -75 845 -45
rect 805 -115 845 -75
rect 805 -145 810 -115
rect 840 -145 845 -115
rect 805 -150 845 -145
rect 1005 -45 1045 -40
rect 1005 -75 1010 -45
rect 1040 -75 1045 -45
rect 1005 -115 1045 -75
rect 1005 -145 1010 -115
rect 1040 -145 1045 -115
rect 1005 -150 1045 -145
rect 1205 -45 1245 -40
rect 1205 -75 1210 -45
rect 1240 -75 1245 -45
rect 1205 -115 1245 -75
rect 1205 -145 1210 -115
rect 1240 -145 1245 -115
rect 1205 -150 1245 -145
rect 1405 -45 1445 -40
rect 1405 -75 1410 -45
rect 1440 -75 1445 -45
rect 1405 -115 1445 -75
rect 1405 -145 1410 -115
rect 1440 -145 1445 -115
rect 1405 -150 1445 -145
rect 1605 -45 1645 -40
rect 1605 -75 1610 -45
rect 1640 -75 1645 -45
rect 1605 -115 1645 -75
rect 1605 -145 1610 -115
rect 1640 -145 1645 -115
rect 1605 -150 1645 -145
rect 1805 -45 1845 -40
rect 1805 -75 1810 -45
rect 1840 -75 1845 -45
rect 1805 -115 1845 -75
rect 1805 -145 1810 -115
rect 1840 -145 1845 -115
rect 1805 -150 1845 -145
rect 2005 -45 2045 -40
rect 2005 -75 2010 -45
rect 2040 -75 2045 -45
rect 2005 -115 2045 -75
rect 2005 -145 2010 -115
rect 2040 -145 2045 -115
rect 2005 -150 2045 -145
rect 2205 -45 2245 -40
rect 2205 -75 2210 -45
rect 2240 -75 2245 -45
rect 2205 -115 2245 -75
rect 2205 -145 2210 -115
rect 2240 -145 2245 -115
rect 2205 -150 2245 -145
rect 2405 -45 2445 -40
rect 2405 -75 2410 -45
rect 2440 -75 2445 -45
rect 2405 -115 2445 -75
rect 2405 -145 2410 -115
rect 2440 -145 2445 -115
rect 2405 -150 2445 -145
rect 2605 -45 2645 -40
rect 2605 -75 2610 -45
rect 2640 -75 2645 -45
rect 2605 -115 2645 -75
rect 2605 -145 2610 -115
rect 2640 -145 2645 -115
rect 2605 -150 2645 -145
rect 2805 -45 2845 -40
rect 2805 -75 2810 -45
rect 2840 -75 2845 -45
rect 2805 -115 2845 -75
rect 2805 -145 2810 -115
rect 2840 -145 2845 -115
rect 2805 -150 2845 -145
rect 3005 -45 3045 -40
rect 3005 -75 3010 -45
rect 3040 -75 3045 -45
rect 3005 -115 3045 -75
rect 3005 -145 3010 -115
rect 3040 -145 3045 -115
rect 3005 -150 3045 -145
rect 3205 -45 3245 -40
rect 3205 -75 3210 -45
rect 3240 -75 3245 -45
rect 3205 -115 3245 -75
rect 3205 -145 3210 -115
rect 3240 -145 3245 -115
rect 3205 -150 3245 -145
rect 3405 -45 3445 -40
rect 3405 -75 3410 -45
rect 3440 -75 3445 -45
rect 3405 -115 3445 -75
rect 3405 -145 3410 -115
rect 3440 -145 3445 -115
rect 3405 -150 3445 -145
rect 3605 -45 3645 -40
rect 3605 -75 3610 -45
rect 3640 -75 3645 -45
rect 3605 -115 3645 -75
rect 3605 -145 3610 -115
rect 3640 -145 3645 -115
rect 3605 -150 3645 -145
rect 3805 -45 3845 -40
rect 3805 -75 3810 -45
rect 3840 -75 3845 -45
rect 3805 -115 3845 -75
rect 3805 -145 3810 -115
rect 3840 -145 3845 -115
rect 3805 -150 3845 -145
rect 4005 -45 4045 -40
rect 4005 -75 4010 -45
rect 4040 -75 4045 -45
rect 4005 -115 4045 -75
rect 4005 -145 4010 -115
rect 4040 -145 4045 -115
rect 4005 -150 4045 -145
rect 4205 -45 4245 -40
rect 4205 -75 4210 -45
rect 4240 -75 4245 -45
rect 4205 -115 4245 -75
rect 4205 -145 4210 -115
rect 4240 -145 4245 -115
rect 4205 -150 4245 -145
rect 4405 -45 4445 -40
rect 4405 -75 4410 -45
rect 4440 -75 4445 -45
rect 4405 -115 4445 -75
rect 4405 -145 4410 -115
rect 4440 -145 4445 -115
rect 4405 -150 4445 -145
rect 4605 -45 4645 -40
rect 4605 -75 4610 -45
rect 4640 -75 4645 -45
rect 4605 -115 4645 -75
rect 4605 -145 4610 -115
rect 4640 -145 4645 -115
rect 4605 -150 4645 -145
rect 4805 -45 4845 -40
rect 4805 -75 4810 -45
rect 4840 -75 4845 -45
rect 4805 -115 4845 -75
rect 4805 -145 4810 -115
rect 4840 -145 4845 -115
rect 4805 -150 4845 -145
rect 5005 -45 5045 -40
rect 5005 -75 5010 -45
rect 5040 -75 5045 -45
rect 5005 -115 5045 -75
rect 5005 -145 5010 -115
rect 5040 -145 5045 -115
rect 5005 -150 5045 -145
rect 5205 -45 5245 -40
rect 5205 -75 5210 -45
rect 5240 -75 5245 -45
rect 5205 -115 5245 -75
rect 5205 -145 5210 -115
rect 5240 -145 5245 -115
rect 5205 -150 5245 -145
rect 5405 -45 5445 -40
rect 5405 -75 5410 -45
rect 5440 -75 5445 -45
rect 5405 -115 5445 -75
rect 5405 -145 5410 -115
rect 5440 -145 5445 -115
rect 5405 -150 5445 -145
rect 5605 -45 5645 -40
rect 5605 -75 5610 -45
rect 5640 -75 5645 -45
rect 5605 -115 5645 -75
rect 5605 -145 5610 -115
rect 5640 -145 5645 -115
rect 5605 -150 5645 -145
rect 5805 -45 5845 -40
rect 5805 -75 5810 -45
rect 5840 -75 5845 -45
rect 5805 -115 5845 -75
rect 5805 -145 5810 -115
rect 5840 -145 5845 -115
rect 5805 -150 5845 -145
rect 6005 -45 6045 -40
rect 6005 -75 6010 -45
rect 6040 -75 6045 -45
rect 6005 -115 6045 -75
rect 6005 -145 6010 -115
rect 6040 -145 6045 -115
rect 6005 -150 6045 -145
rect 6205 -45 6245 -40
rect 6205 -75 6210 -45
rect 6240 -75 6245 -45
rect 6205 -115 6245 -75
rect 6205 -145 6210 -115
rect 6240 -145 6245 -115
rect 6205 -150 6245 -145
rect 6405 -45 6445 -40
rect 6405 -75 6410 -45
rect 6440 -75 6445 -45
rect 6405 -115 6445 -75
rect 6405 -145 6410 -115
rect 6440 -145 6445 -115
rect 6405 -150 6445 -145
<< via2 >>
rect -140 12060 -110 12090
rect -90 12060 -60 12090
rect 6460 12035 6490 12065
rect 6510 12035 6540 12065
rect -190 11950 -160 11980
rect -190 11880 -160 11910
rect 10 11950 40 11980
rect 10 11880 40 11910
rect 210 11950 240 11980
rect 210 11880 240 11910
rect 410 11950 440 11980
rect 410 11880 440 11910
rect 610 11950 640 11980
rect 610 11880 640 11910
rect 810 11950 840 11980
rect 810 11880 840 11910
rect 1010 11950 1040 11980
rect 1010 11880 1040 11910
rect 1210 11950 1240 11980
rect 1210 11880 1240 11910
rect 1410 11950 1440 11980
rect 1410 11880 1440 11910
rect 1610 11950 1640 11980
rect 1610 11880 1640 11910
rect 1810 11950 1840 11980
rect 1810 11880 1840 11910
rect 2010 11950 2040 11980
rect 2010 11880 2040 11910
rect 2210 11950 2240 11980
rect 2210 11880 2240 11910
rect 2410 11950 2440 11980
rect 2410 11880 2440 11910
rect 2610 11950 2640 11980
rect 2610 11880 2640 11910
rect 2810 11950 2840 11980
rect 2810 11880 2840 11910
rect 3010 11950 3040 11980
rect 3010 11880 3040 11910
rect 3210 11950 3240 11980
rect 3210 11880 3240 11910
rect 3410 11950 3440 11980
rect 3410 11880 3440 11910
rect 3610 11950 3640 11980
rect 3610 11880 3640 11910
rect 3810 11950 3840 11980
rect 3810 11880 3840 11910
rect 4010 11950 4040 11980
rect 4010 11880 4040 11910
rect 4210 11950 4240 11980
rect 4210 11880 4240 11910
rect 4410 11950 4440 11980
rect 4410 11880 4440 11910
rect 4610 11950 4640 11980
rect 4610 11880 4640 11910
rect 4810 11950 4840 11980
rect 4810 11880 4840 11910
rect 5010 11950 5040 11980
rect 5010 11880 5040 11910
rect 5210 11950 5240 11980
rect 5210 11880 5240 11910
rect 5410 11950 5440 11980
rect 5410 11880 5440 11910
rect 5610 11950 5640 11980
rect 5610 11880 5640 11910
rect 5810 11950 5840 11980
rect 5810 11880 5840 11910
rect 6010 11950 6040 11980
rect 6010 11880 6040 11910
rect 6210 11950 6240 11980
rect 6210 11880 6240 11910
rect 6410 11950 6440 11980
rect 6410 11880 6440 11910
rect -190 11765 -160 11795
rect -190 11695 -160 11725
rect 10 11765 40 11795
rect 10 11695 40 11725
rect 210 11765 240 11795
rect 210 11695 240 11725
rect 410 11765 440 11795
rect 410 11695 440 11725
rect 610 11765 640 11795
rect 610 11695 640 11725
rect 810 11765 840 11795
rect 810 11695 840 11725
rect 1010 11765 1040 11795
rect 1010 11695 1040 11725
rect 1210 11765 1240 11795
rect 1210 11695 1240 11725
rect 1410 11765 1440 11795
rect 1410 11695 1440 11725
rect 1610 11765 1640 11795
rect 1610 11695 1640 11725
rect 1810 11765 1840 11795
rect 1810 11695 1840 11725
rect 2010 11765 2040 11795
rect 2010 11695 2040 11725
rect 2210 11765 2240 11795
rect 2210 11695 2240 11725
rect 2410 11765 2440 11795
rect 2410 11695 2440 11725
rect 2610 11765 2640 11795
rect 2610 11695 2640 11725
rect 2810 11765 2840 11795
rect 2810 11695 2840 11725
rect 3010 11765 3040 11795
rect 3010 11695 3040 11725
rect 3210 11765 3240 11795
rect 3210 11695 3240 11725
rect 3410 11765 3440 11795
rect 3410 11695 3440 11725
rect 3610 11765 3640 11795
rect 3610 11695 3640 11725
rect 3810 11765 3840 11795
rect 3810 11695 3840 11725
rect 4010 11765 4040 11795
rect 4010 11695 4040 11725
rect 4210 11765 4240 11795
rect 4210 11695 4240 11725
rect 4410 11765 4440 11795
rect 4410 11695 4440 11725
rect 4610 11765 4640 11795
rect 4610 11695 4640 11725
rect 4810 11765 4840 11795
rect 4810 11695 4840 11725
rect 5010 11765 5040 11795
rect 5010 11695 5040 11725
rect 5210 11765 5240 11795
rect 5210 11695 5240 11725
rect 5410 11765 5440 11795
rect 5410 11695 5440 11725
rect 5610 11765 5640 11795
rect 5610 11695 5640 11725
rect 5810 11765 5840 11795
rect 5810 11695 5840 11725
rect 6010 11765 6040 11795
rect 6010 11695 6040 11725
rect 6210 11765 6240 11795
rect 6210 11695 6240 11725
rect 6410 11765 6440 11795
rect 6410 11695 6440 11725
rect -190 11580 -160 11610
rect -190 11510 -160 11540
rect 10 11580 40 11610
rect 10 11510 40 11540
rect 210 11580 240 11610
rect 210 11510 240 11540
rect 410 11580 440 11610
rect 410 11510 440 11540
rect 610 11580 640 11610
rect 610 11510 640 11540
rect 810 11580 840 11610
rect 810 11510 840 11540
rect 1010 11580 1040 11610
rect 1010 11510 1040 11540
rect 1210 11580 1240 11610
rect 1210 11510 1240 11540
rect 1410 11580 1440 11610
rect 1410 11510 1440 11540
rect 1610 11580 1640 11610
rect 1610 11510 1640 11540
rect 1810 11580 1840 11610
rect 1810 11510 1840 11540
rect 2010 11580 2040 11610
rect 2010 11510 2040 11540
rect 2210 11580 2240 11610
rect 2210 11510 2240 11540
rect 2410 11580 2440 11610
rect 2410 11510 2440 11540
rect 2610 11580 2640 11610
rect 2610 11510 2640 11540
rect 2810 11580 2840 11610
rect 2810 11510 2840 11540
rect 3010 11580 3040 11610
rect 3010 11510 3040 11540
rect 3210 11580 3240 11610
rect 3210 11510 3240 11540
rect 3410 11580 3440 11610
rect 3410 11510 3440 11540
rect 3610 11580 3640 11610
rect 3610 11510 3640 11540
rect 3810 11580 3840 11610
rect 3810 11510 3840 11540
rect 4010 11580 4040 11610
rect 4010 11510 4040 11540
rect 4210 11580 4240 11610
rect 4210 11510 4240 11540
rect 4410 11580 4440 11610
rect 4410 11510 4440 11540
rect 4610 11580 4640 11610
rect 4610 11510 4640 11540
rect 4810 11580 4840 11610
rect 4810 11510 4840 11540
rect 5010 11580 5040 11610
rect 5010 11510 5040 11540
rect 5210 11580 5240 11610
rect 5210 11510 5240 11540
rect 5410 11580 5440 11610
rect 5410 11510 5440 11540
rect 5610 11580 5640 11610
rect 5610 11510 5640 11540
rect 5810 11580 5840 11610
rect 5810 11510 5840 11540
rect 6010 11580 6040 11610
rect 6010 11510 6040 11540
rect 6210 11580 6240 11610
rect 6210 11510 6240 11540
rect 6410 11580 6440 11610
rect 6410 11510 6440 11540
rect -190 11395 -160 11425
rect -190 11325 -160 11355
rect 10 11395 40 11425
rect 10 11325 40 11355
rect 210 11395 240 11425
rect 210 11325 240 11355
rect 410 11395 440 11425
rect 410 11325 440 11355
rect 610 11395 640 11425
rect 610 11325 640 11355
rect 810 11395 840 11425
rect 810 11325 840 11355
rect 1010 11395 1040 11425
rect 1010 11325 1040 11355
rect 1210 11395 1240 11425
rect 1210 11325 1240 11355
rect 1410 11395 1440 11425
rect 1410 11325 1440 11355
rect 1610 11395 1640 11425
rect 1610 11325 1640 11355
rect 1810 11395 1840 11425
rect 1810 11325 1840 11355
rect 2010 11395 2040 11425
rect 2010 11325 2040 11355
rect 2210 11395 2240 11425
rect 2210 11325 2240 11355
rect 2410 11395 2440 11425
rect 2410 11325 2440 11355
rect 2610 11395 2640 11425
rect 2610 11325 2640 11355
rect 2810 11395 2840 11425
rect 2810 11325 2840 11355
rect 3010 11395 3040 11425
rect 3010 11325 3040 11355
rect 3210 11395 3240 11425
rect 3210 11325 3240 11355
rect 3410 11395 3440 11425
rect 3410 11325 3440 11355
rect 3610 11395 3640 11425
rect 3610 11325 3640 11355
rect 3810 11395 3840 11425
rect 3810 11325 3840 11355
rect 4010 11395 4040 11425
rect 4010 11325 4040 11355
rect 4210 11395 4240 11425
rect 4210 11325 4240 11355
rect 4410 11395 4440 11425
rect 4410 11325 4440 11355
rect 4610 11395 4640 11425
rect 4610 11325 4640 11355
rect 4810 11395 4840 11425
rect 4810 11325 4840 11355
rect 5010 11395 5040 11425
rect 5010 11325 5040 11355
rect 5210 11395 5240 11425
rect 5210 11325 5240 11355
rect 5410 11395 5440 11425
rect 5410 11325 5440 11355
rect 5610 11395 5640 11425
rect 5610 11325 5640 11355
rect 5810 11395 5840 11425
rect 5810 11325 5840 11355
rect 6010 11395 6040 11425
rect 6010 11325 6040 11355
rect 6210 11395 6240 11425
rect 6210 11325 6240 11355
rect 6410 11395 6440 11425
rect 6410 11325 6440 11355
rect -190 11210 -160 11240
rect -190 11140 -160 11170
rect 10 11210 40 11240
rect 10 11140 40 11170
rect 210 11210 240 11240
rect 210 11140 240 11170
rect 410 11210 440 11240
rect 410 11140 440 11170
rect 610 11210 640 11240
rect 610 11140 640 11170
rect 810 11210 840 11240
rect 810 11140 840 11170
rect 1010 11210 1040 11240
rect 1010 11140 1040 11170
rect 1210 11210 1240 11240
rect 1210 11140 1240 11170
rect 1410 11210 1440 11240
rect 1410 11140 1440 11170
rect 1610 11210 1640 11240
rect 1610 11140 1640 11170
rect 1810 11210 1840 11240
rect 1810 11140 1840 11170
rect 2010 11210 2040 11240
rect 2010 11140 2040 11170
rect 2210 11210 2240 11240
rect 2210 11140 2240 11170
rect 2410 11210 2440 11240
rect 2410 11140 2440 11170
rect 2610 11210 2640 11240
rect 2610 11140 2640 11170
rect 2810 11210 2840 11240
rect 2810 11140 2840 11170
rect 3010 11210 3040 11240
rect 3010 11140 3040 11170
rect 3210 11210 3240 11240
rect 3210 11140 3240 11170
rect 3410 11210 3440 11240
rect 3410 11140 3440 11170
rect 3610 11210 3640 11240
rect 3610 11140 3640 11170
rect 3810 11210 3840 11240
rect 3810 11140 3840 11170
rect 4010 11210 4040 11240
rect 4010 11140 4040 11170
rect 4210 11210 4240 11240
rect 4210 11140 4240 11170
rect 4410 11210 4440 11240
rect 4410 11140 4440 11170
rect 4610 11210 4640 11240
rect 4610 11140 4640 11170
rect 4810 11210 4840 11240
rect 4810 11140 4840 11170
rect 5010 11210 5040 11240
rect 5010 11140 5040 11170
rect 5210 11210 5240 11240
rect 5210 11140 5240 11170
rect 5410 11210 5440 11240
rect 5410 11140 5440 11170
rect 5610 11210 5640 11240
rect 5610 11140 5640 11170
rect 5810 11210 5840 11240
rect 5810 11140 5840 11170
rect 6010 11210 6040 11240
rect 6010 11140 6040 11170
rect 6210 11210 6240 11240
rect 6210 11140 6240 11170
rect 6410 11210 6440 11240
rect 6410 11140 6440 11170
rect -190 11025 -160 11055
rect -190 10955 -160 10985
rect 10 11025 40 11055
rect 10 10955 40 10985
rect 210 11025 240 11055
rect 210 10955 240 10985
rect 410 11025 440 11055
rect 410 10955 440 10985
rect 610 11025 640 11055
rect 610 10955 640 10985
rect 810 11025 840 11055
rect 810 10955 840 10985
rect 1010 11025 1040 11055
rect 1010 10955 1040 10985
rect 1210 11025 1240 11055
rect 1210 10955 1240 10985
rect 1410 11025 1440 11055
rect 1410 10955 1440 10985
rect 1610 11025 1640 11055
rect 1610 10955 1640 10985
rect 1810 11025 1840 11055
rect 1810 10955 1840 10985
rect 2010 11025 2040 11055
rect 2010 10955 2040 10985
rect 2210 11025 2240 11055
rect 2210 10955 2240 10985
rect 2410 11025 2440 11055
rect 2410 10955 2440 10985
rect 2610 11025 2640 11055
rect 2610 10955 2640 10985
rect 2810 11025 2840 11055
rect 2810 10955 2840 10985
rect 3010 11025 3040 11055
rect 3010 10955 3040 10985
rect 3210 11025 3240 11055
rect 3210 10955 3240 10985
rect 3410 11025 3440 11055
rect 3410 10955 3440 10985
rect 3610 11025 3640 11055
rect 3610 10955 3640 10985
rect 3810 11025 3840 11055
rect 3810 10955 3840 10985
rect 4010 11025 4040 11055
rect 4010 10955 4040 10985
rect 4210 11025 4240 11055
rect 4210 10955 4240 10985
rect 4410 11025 4440 11055
rect 4410 10955 4440 10985
rect 4610 11025 4640 11055
rect 4610 10955 4640 10985
rect 4810 11025 4840 11055
rect 4810 10955 4840 10985
rect 5010 11025 5040 11055
rect 5010 10955 5040 10985
rect 5210 11025 5240 11055
rect 5210 10955 5240 10985
rect 5410 11025 5440 11055
rect 5410 10955 5440 10985
rect 5610 11025 5640 11055
rect 5610 10955 5640 10985
rect 5810 11025 5840 11055
rect 5810 10955 5840 10985
rect 6010 11025 6040 11055
rect 6010 10955 6040 10985
rect 6210 11025 6240 11055
rect 6210 10955 6240 10985
rect 6410 11025 6440 11055
rect 6410 10955 6440 10985
rect -190 10840 -160 10870
rect -190 10770 -160 10800
rect 10 10840 40 10870
rect 10 10770 40 10800
rect 210 10840 240 10870
rect 210 10770 240 10800
rect 410 10840 440 10870
rect 410 10770 440 10800
rect 610 10840 640 10870
rect 610 10770 640 10800
rect 810 10840 840 10870
rect 810 10770 840 10800
rect 1010 10840 1040 10870
rect 1010 10770 1040 10800
rect 1210 10840 1240 10870
rect 1210 10770 1240 10800
rect 1410 10840 1440 10870
rect 1410 10770 1440 10800
rect 1610 10840 1640 10870
rect 1610 10770 1640 10800
rect 1810 10840 1840 10870
rect 1810 10770 1840 10800
rect 2010 10840 2040 10870
rect 2010 10770 2040 10800
rect 2210 10840 2240 10870
rect 2210 10770 2240 10800
rect 2410 10840 2440 10870
rect 2410 10770 2440 10800
rect 2610 10840 2640 10870
rect 2610 10770 2640 10800
rect 2810 10840 2840 10870
rect 2810 10770 2840 10800
rect 3010 10840 3040 10870
rect 3010 10770 3040 10800
rect 3210 10840 3240 10870
rect 3210 10770 3240 10800
rect 3410 10840 3440 10870
rect 3410 10770 3440 10800
rect 3610 10840 3640 10870
rect 3610 10770 3640 10800
rect 3810 10840 3840 10870
rect 3810 10770 3840 10800
rect 4010 10840 4040 10870
rect 4010 10770 4040 10800
rect 4210 10840 4240 10870
rect 4210 10770 4240 10800
rect 4410 10840 4440 10870
rect 4410 10770 4440 10800
rect 4610 10840 4640 10870
rect 4610 10770 4640 10800
rect 4810 10840 4840 10870
rect 4810 10770 4840 10800
rect 5010 10840 5040 10870
rect 5010 10770 5040 10800
rect 5210 10840 5240 10870
rect 5210 10770 5240 10800
rect 5410 10840 5440 10870
rect 5410 10770 5440 10800
rect 5610 10840 5640 10870
rect 5610 10770 5640 10800
rect 5810 10840 5840 10870
rect 5810 10770 5840 10800
rect 6010 10840 6040 10870
rect 6010 10770 6040 10800
rect 6210 10840 6240 10870
rect 6210 10770 6240 10800
rect 6410 10840 6440 10870
rect 6410 10770 6440 10800
rect -190 10655 -160 10685
rect -190 10585 -160 10615
rect 10 10655 40 10685
rect 10 10585 40 10615
rect 210 10655 240 10685
rect 210 10585 240 10615
rect 410 10655 440 10685
rect 410 10585 440 10615
rect 610 10655 640 10685
rect 610 10585 640 10615
rect 810 10655 840 10685
rect 810 10585 840 10615
rect 1010 10655 1040 10685
rect 1010 10585 1040 10615
rect 1210 10655 1240 10685
rect 1210 10585 1240 10615
rect 1410 10655 1440 10685
rect 1410 10585 1440 10615
rect 1610 10655 1640 10685
rect 1610 10585 1640 10615
rect 1810 10655 1840 10685
rect 1810 10585 1840 10615
rect 2010 10655 2040 10685
rect 2010 10585 2040 10615
rect 2210 10655 2240 10685
rect 2210 10585 2240 10615
rect 2410 10655 2440 10685
rect 2410 10585 2440 10615
rect 2610 10655 2640 10685
rect 2610 10585 2640 10615
rect 2810 10655 2840 10685
rect 2810 10585 2840 10615
rect 3010 10655 3040 10685
rect 3010 10585 3040 10615
rect 3210 10655 3240 10685
rect 3210 10585 3240 10615
rect 3410 10655 3440 10685
rect 3410 10585 3440 10615
rect 3610 10655 3640 10685
rect 3610 10585 3640 10615
rect 3810 10655 3840 10685
rect 3810 10585 3840 10615
rect 4010 10655 4040 10685
rect 4010 10585 4040 10615
rect 4210 10655 4240 10685
rect 4210 10585 4240 10615
rect 4410 10655 4440 10685
rect 4410 10585 4440 10615
rect 4610 10655 4640 10685
rect 4610 10585 4640 10615
rect 4810 10655 4840 10685
rect 4810 10585 4840 10615
rect 5010 10655 5040 10685
rect 5010 10585 5040 10615
rect 5210 10655 5240 10685
rect 5210 10585 5240 10615
rect 5410 10655 5440 10685
rect 5410 10585 5440 10615
rect 5610 10655 5640 10685
rect 5610 10585 5640 10615
rect 5810 10655 5840 10685
rect 5810 10585 5840 10615
rect 6010 10655 6040 10685
rect 6010 10585 6040 10615
rect 6210 10655 6240 10685
rect 6210 10585 6240 10615
rect 6410 10655 6440 10685
rect 6410 10585 6440 10615
rect -190 10470 -160 10500
rect -190 10400 -160 10430
rect 10 10470 40 10500
rect 10 10400 40 10430
rect 210 10470 240 10500
rect 210 10400 240 10430
rect 410 10470 440 10500
rect 410 10400 440 10430
rect 610 10470 640 10500
rect 610 10400 640 10430
rect 810 10470 840 10500
rect 810 10400 840 10430
rect 1010 10470 1040 10500
rect 1010 10400 1040 10430
rect 1210 10470 1240 10500
rect 1210 10400 1240 10430
rect 1410 10470 1440 10500
rect 1410 10400 1440 10430
rect 1610 10470 1640 10500
rect 1610 10400 1640 10430
rect 1810 10470 1840 10500
rect 1810 10400 1840 10430
rect 2010 10470 2040 10500
rect 2010 10400 2040 10430
rect 2210 10470 2240 10500
rect 2210 10400 2240 10430
rect 2410 10470 2440 10500
rect 2410 10400 2440 10430
rect 2610 10470 2640 10500
rect 2610 10400 2640 10430
rect 2810 10470 2840 10500
rect 2810 10400 2840 10430
rect 3010 10470 3040 10500
rect 3010 10400 3040 10430
rect 3210 10470 3240 10500
rect 3210 10400 3240 10430
rect 3410 10470 3440 10500
rect 3410 10400 3440 10430
rect 3610 10470 3640 10500
rect 3610 10400 3640 10430
rect 3810 10470 3840 10500
rect 3810 10400 3840 10430
rect 4010 10470 4040 10500
rect 4010 10400 4040 10430
rect 4210 10470 4240 10500
rect 4210 10400 4240 10430
rect 4410 10470 4440 10500
rect 4410 10400 4440 10430
rect 4610 10470 4640 10500
rect 4610 10400 4640 10430
rect 4810 10470 4840 10500
rect 4810 10400 4840 10430
rect 5010 10470 5040 10500
rect 5010 10400 5040 10430
rect 5210 10470 5240 10500
rect 5210 10400 5240 10430
rect 5410 10470 5440 10500
rect 5410 10400 5440 10430
rect 5610 10470 5640 10500
rect 5610 10400 5640 10430
rect 5810 10470 5840 10500
rect 5810 10400 5840 10430
rect 6010 10470 6040 10500
rect 6010 10400 6040 10430
rect 6210 10470 6240 10500
rect 6210 10400 6240 10430
rect 6410 10470 6440 10500
rect 6410 10400 6440 10430
rect -190 10285 -160 10315
rect -190 10215 -160 10245
rect 10 10285 40 10315
rect 10 10215 40 10245
rect 210 10285 240 10315
rect 210 10215 240 10245
rect 410 10285 440 10315
rect 410 10215 440 10245
rect 610 10285 640 10315
rect 610 10215 640 10245
rect 810 10285 840 10315
rect 810 10215 840 10245
rect 1010 10285 1040 10315
rect 1010 10215 1040 10245
rect 1210 10285 1240 10315
rect 1210 10215 1240 10245
rect 1410 10285 1440 10315
rect 1410 10215 1440 10245
rect 1610 10285 1640 10315
rect 1610 10215 1640 10245
rect 1810 10285 1840 10315
rect 1810 10215 1840 10245
rect 2010 10285 2040 10315
rect 2010 10215 2040 10245
rect 2210 10285 2240 10315
rect 2210 10215 2240 10245
rect 2410 10285 2440 10315
rect 2410 10215 2440 10245
rect 2610 10285 2640 10315
rect 2610 10215 2640 10245
rect 2810 10285 2840 10315
rect 2810 10215 2840 10245
rect 3010 10285 3040 10315
rect 3010 10215 3040 10245
rect 3210 10285 3240 10315
rect 3210 10215 3240 10245
rect 3410 10285 3440 10315
rect 3410 10215 3440 10245
rect 3610 10285 3640 10315
rect 3610 10215 3640 10245
rect 3810 10285 3840 10315
rect 3810 10215 3840 10245
rect 4010 10285 4040 10315
rect 4010 10215 4040 10245
rect 4210 10285 4240 10315
rect 4210 10215 4240 10245
rect 4410 10285 4440 10315
rect 4410 10215 4440 10245
rect 4610 10285 4640 10315
rect 4610 10215 4640 10245
rect 4810 10285 4840 10315
rect 4810 10215 4840 10245
rect 5010 10285 5040 10315
rect 5010 10215 5040 10245
rect 5210 10285 5240 10315
rect 5210 10215 5240 10245
rect 5410 10285 5440 10315
rect 5410 10215 5440 10245
rect 5610 10285 5640 10315
rect 5610 10215 5640 10245
rect 5810 10285 5840 10315
rect 5810 10215 5840 10245
rect 6010 10285 6040 10315
rect 6010 10215 6040 10245
rect 6210 10285 6240 10315
rect 6210 10215 6240 10245
rect 6410 10285 6440 10315
rect 6410 10215 6440 10245
rect -190 10100 -160 10130
rect -190 10030 -160 10060
rect 10 10100 40 10130
rect 10 10030 40 10060
rect 210 10100 240 10130
rect 210 10030 240 10060
rect 410 10100 440 10130
rect 410 10030 440 10060
rect 610 10100 640 10130
rect 610 10030 640 10060
rect 810 10100 840 10130
rect 810 10030 840 10060
rect 1010 10100 1040 10130
rect 1010 10030 1040 10060
rect 1210 10100 1240 10130
rect 1210 10030 1240 10060
rect 1410 10100 1440 10130
rect 1410 10030 1440 10060
rect 1610 10100 1640 10130
rect 1610 10030 1640 10060
rect 1810 10100 1840 10130
rect 1810 10030 1840 10060
rect 2010 10100 2040 10130
rect 2010 10030 2040 10060
rect 2210 10100 2240 10130
rect 2210 10030 2240 10060
rect 2410 10100 2440 10130
rect 2410 10030 2440 10060
rect 2610 10100 2640 10130
rect 2610 10030 2640 10060
rect 2810 10100 2840 10130
rect 2810 10030 2840 10060
rect 3010 10100 3040 10130
rect 3010 10030 3040 10060
rect 3210 10100 3240 10130
rect 3210 10030 3240 10060
rect 3410 10100 3440 10130
rect 3410 10030 3440 10060
rect 3610 10100 3640 10130
rect 3610 10030 3640 10060
rect 3810 10100 3840 10130
rect 3810 10030 3840 10060
rect 4010 10100 4040 10130
rect 4010 10030 4040 10060
rect 4210 10100 4240 10130
rect 4210 10030 4240 10060
rect 4410 10100 4440 10130
rect 4410 10030 4440 10060
rect 4610 10100 4640 10130
rect 4610 10030 4640 10060
rect 4810 10100 4840 10130
rect 4810 10030 4840 10060
rect 5010 10100 5040 10130
rect 5010 10030 5040 10060
rect 5210 10100 5240 10130
rect 5210 10030 5240 10060
rect 5410 10100 5440 10130
rect 5410 10030 5440 10060
rect 5610 10100 5640 10130
rect 5610 10030 5640 10060
rect 5810 10100 5840 10130
rect 5810 10030 5840 10060
rect 6010 10100 6040 10130
rect 6010 10030 6040 10060
rect 6210 10100 6240 10130
rect 6210 10030 6240 10060
rect 6410 10100 6440 10130
rect 6410 10030 6440 10060
rect -190 9915 -160 9945
rect -190 9845 -160 9875
rect 10 9915 40 9945
rect 10 9845 40 9875
rect 210 9915 240 9945
rect 210 9845 240 9875
rect 410 9915 440 9945
rect 410 9845 440 9875
rect 610 9915 640 9945
rect 610 9845 640 9875
rect 810 9915 840 9945
rect 810 9845 840 9875
rect 1010 9915 1040 9945
rect 1010 9845 1040 9875
rect 1210 9915 1240 9945
rect 1210 9845 1240 9875
rect 1410 9915 1440 9945
rect 1410 9845 1440 9875
rect 1610 9915 1640 9945
rect 1610 9845 1640 9875
rect 1810 9915 1840 9945
rect 1810 9845 1840 9875
rect 2010 9915 2040 9945
rect 2010 9845 2040 9875
rect 2210 9915 2240 9945
rect 2210 9845 2240 9875
rect 2410 9915 2440 9945
rect 2410 9845 2440 9875
rect 2610 9915 2640 9945
rect 2610 9845 2640 9875
rect 2810 9915 2840 9945
rect 2810 9845 2840 9875
rect 3010 9915 3040 9945
rect 3010 9845 3040 9875
rect 3210 9915 3240 9945
rect 3210 9845 3240 9875
rect 3410 9915 3440 9945
rect 3410 9845 3440 9875
rect 3610 9915 3640 9945
rect 3610 9845 3640 9875
rect 3810 9915 3840 9945
rect 3810 9845 3840 9875
rect 4010 9915 4040 9945
rect 4010 9845 4040 9875
rect 4210 9915 4240 9945
rect 4210 9845 4240 9875
rect 4410 9915 4440 9945
rect 4410 9845 4440 9875
rect 4610 9915 4640 9945
rect 4610 9845 4640 9875
rect 4810 9915 4840 9945
rect 4810 9845 4840 9875
rect 5010 9915 5040 9945
rect 5010 9845 5040 9875
rect 5210 9915 5240 9945
rect 5210 9845 5240 9875
rect 5410 9915 5440 9945
rect 5410 9845 5440 9875
rect 5610 9915 5640 9945
rect 5610 9845 5640 9875
rect 5810 9915 5840 9945
rect 5810 9845 5840 9875
rect 6010 9915 6040 9945
rect 6010 9845 6040 9875
rect 6210 9915 6240 9945
rect 6210 9845 6240 9875
rect 6410 9915 6440 9945
rect 6410 9845 6440 9875
rect -190 9730 -160 9760
rect -190 9660 -160 9690
rect 10 9730 40 9760
rect 10 9660 40 9690
rect 210 9730 240 9760
rect 210 9660 240 9690
rect 410 9730 440 9760
rect 410 9660 440 9690
rect 610 9730 640 9760
rect 610 9660 640 9690
rect 810 9730 840 9760
rect 810 9660 840 9690
rect 1010 9730 1040 9760
rect 1010 9660 1040 9690
rect 1210 9730 1240 9760
rect 1210 9660 1240 9690
rect 1410 9730 1440 9760
rect 1410 9660 1440 9690
rect 1610 9730 1640 9760
rect 1610 9660 1640 9690
rect 1810 9730 1840 9760
rect 1810 9660 1840 9690
rect 2010 9730 2040 9760
rect 2010 9660 2040 9690
rect 2210 9730 2240 9760
rect 2210 9660 2240 9690
rect 2410 9730 2440 9760
rect 2410 9660 2440 9690
rect 2610 9730 2640 9760
rect 2610 9660 2640 9690
rect 2810 9730 2840 9760
rect 2810 9660 2840 9690
rect 3010 9730 3040 9760
rect 3010 9660 3040 9690
rect 3210 9730 3240 9760
rect 3210 9660 3240 9690
rect 3410 9730 3440 9760
rect 3410 9660 3440 9690
rect 3610 9730 3640 9760
rect 3610 9660 3640 9690
rect 3810 9730 3840 9760
rect 3810 9660 3840 9690
rect 4010 9730 4040 9760
rect 4010 9660 4040 9690
rect 4210 9730 4240 9760
rect 4210 9660 4240 9690
rect 4410 9730 4440 9760
rect 4410 9660 4440 9690
rect 4610 9730 4640 9760
rect 4610 9660 4640 9690
rect 4810 9730 4840 9760
rect 4810 9660 4840 9690
rect 5010 9730 5040 9760
rect 5010 9660 5040 9690
rect 5210 9730 5240 9760
rect 5210 9660 5240 9690
rect 5410 9730 5440 9760
rect 5410 9660 5440 9690
rect 5610 9730 5640 9760
rect 5610 9660 5640 9690
rect 5810 9730 5840 9760
rect 5810 9660 5840 9690
rect 6010 9730 6040 9760
rect 6010 9660 6040 9690
rect 6210 9730 6240 9760
rect 6210 9660 6240 9690
rect 6410 9730 6440 9760
rect 6410 9660 6440 9690
rect -190 9545 -160 9575
rect -190 9475 -160 9505
rect 10 9545 40 9575
rect 10 9475 40 9505
rect 210 9545 240 9575
rect 210 9475 240 9505
rect 410 9545 440 9575
rect 410 9475 440 9505
rect 610 9545 640 9575
rect 610 9475 640 9505
rect 810 9545 840 9575
rect 810 9475 840 9505
rect 1010 9545 1040 9575
rect 1010 9475 1040 9505
rect 1210 9545 1240 9575
rect 1210 9475 1240 9505
rect 1410 9545 1440 9575
rect 1410 9475 1440 9505
rect 1610 9545 1640 9575
rect 1610 9475 1640 9505
rect 1810 9545 1840 9575
rect 1810 9475 1840 9505
rect 2010 9545 2040 9575
rect 2010 9475 2040 9505
rect 2210 9545 2240 9575
rect 2210 9475 2240 9505
rect 2410 9545 2440 9575
rect 2410 9475 2440 9505
rect 2610 9545 2640 9575
rect 2610 9475 2640 9505
rect 2810 9545 2840 9575
rect 2810 9475 2840 9505
rect 3010 9545 3040 9575
rect 3010 9475 3040 9505
rect 3210 9545 3240 9575
rect 3210 9475 3240 9505
rect 3410 9545 3440 9575
rect 3410 9475 3440 9505
rect 3610 9545 3640 9575
rect 3610 9475 3640 9505
rect 3810 9545 3840 9575
rect 3810 9475 3840 9505
rect 4010 9545 4040 9575
rect 4010 9475 4040 9505
rect 4210 9545 4240 9575
rect 4210 9475 4240 9505
rect 4410 9545 4440 9575
rect 4410 9475 4440 9505
rect 4610 9545 4640 9575
rect 4610 9475 4640 9505
rect 4810 9545 4840 9575
rect 4810 9475 4840 9505
rect 5010 9545 5040 9575
rect 5010 9475 5040 9505
rect 5210 9545 5240 9575
rect 5210 9475 5240 9505
rect 5410 9545 5440 9575
rect 5410 9475 5440 9505
rect 5610 9545 5640 9575
rect 5610 9475 5640 9505
rect 5810 9545 5840 9575
rect 5810 9475 5840 9505
rect 6010 9545 6040 9575
rect 6010 9475 6040 9505
rect 6210 9545 6240 9575
rect 6210 9475 6240 9505
rect 6410 9545 6440 9575
rect 6410 9475 6440 9505
rect -190 9360 -160 9390
rect -190 9290 -160 9320
rect 10 9360 40 9390
rect 10 9290 40 9320
rect 210 9360 240 9390
rect 210 9290 240 9320
rect 410 9360 440 9390
rect 410 9290 440 9320
rect 610 9360 640 9390
rect 610 9290 640 9320
rect 810 9360 840 9390
rect 810 9290 840 9320
rect 1010 9360 1040 9390
rect 1010 9290 1040 9320
rect 1210 9360 1240 9390
rect 1210 9290 1240 9320
rect 1410 9360 1440 9390
rect 1410 9290 1440 9320
rect 1610 9360 1640 9390
rect 1610 9290 1640 9320
rect 1810 9360 1840 9390
rect 1810 9290 1840 9320
rect 2010 9360 2040 9390
rect 2010 9290 2040 9320
rect 2210 9360 2240 9390
rect 2210 9290 2240 9320
rect 2410 9360 2440 9390
rect 2410 9290 2440 9320
rect 2610 9360 2640 9390
rect 2610 9290 2640 9320
rect 2810 9360 2840 9390
rect 2810 9290 2840 9320
rect 3010 9360 3040 9390
rect 3010 9290 3040 9320
rect 3210 9360 3240 9390
rect 3210 9290 3240 9320
rect 3410 9360 3440 9390
rect 3410 9290 3440 9320
rect 3610 9360 3640 9390
rect 3610 9290 3640 9320
rect 3810 9360 3840 9390
rect 3810 9290 3840 9320
rect 4010 9360 4040 9390
rect 4010 9290 4040 9320
rect 4210 9360 4240 9390
rect 4210 9290 4240 9320
rect 4410 9360 4440 9390
rect 4410 9290 4440 9320
rect 4610 9360 4640 9390
rect 4610 9290 4640 9320
rect 4810 9360 4840 9390
rect 4810 9290 4840 9320
rect 5010 9360 5040 9390
rect 5010 9290 5040 9320
rect 5210 9360 5240 9390
rect 5210 9290 5240 9320
rect 5410 9360 5440 9390
rect 5410 9290 5440 9320
rect 5610 9360 5640 9390
rect 5610 9290 5640 9320
rect 5810 9360 5840 9390
rect 5810 9290 5840 9320
rect 6010 9360 6040 9390
rect 6010 9290 6040 9320
rect 6210 9360 6240 9390
rect 6210 9290 6240 9320
rect 6410 9360 6440 9390
rect 6410 9290 6440 9320
rect -190 9175 -160 9205
rect -190 9105 -160 9135
rect 10 9175 40 9205
rect 10 9105 40 9135
rect 210 9175 240 9205
rect 210 9105 240 9135
rect 410 9175 440 9205
rect 410 9105 440 9135
rect 610 9175 640 9205
rect 610 9105 640 9135
rect 810 9175 840 9205
rect 810 9105 840 9135
rect 1010 9175 1040 9205
rect 1010 9105 1040 9135
rect 1210 9175 1240 9205
rect 1210 9105 1240 9135
rect 1410 9175 1440 9205
rect 1410 9105 1440 9135
rect 1610 9175 1640 9205
rect 1610 9105 1640 9135
rect 1810 9175 1840 9205
rect 1810 9105 1840 9135
rect 2010 9175 2040 9205
rect 2010 9105 2040 9135
rect 2210 9175 2240 9205
rect 2210 9105 2240 9135
rect 2410 9175 2440 9205
rect 2410 9105 2440 9135
rect 2610 9175 2640 9205
rect 2610 9105 2640 9135
rect 2810 9175 2840 9205
rect 2810 9105 2840 9135
rect 3010 9175 3040 9205
rect 3010 9105 3040 9135
rect 3210 9175 3240 9205
rect 3210 9105 3240 9135
rect 3410 9175 3440 9205
rect 3410 9105 3440 9135
rect 3610 9175 3640 9205
rect 3610 9105 3640 9135
rect 3810 9175 3840 9205
rect 3810 9105 3840 9135
rect 4010 9175 4040 9205
rect 4010 9105 4040 9135
rect 4210 9175 4240 9205
rect 4210 9105 4240 9135
rect 4410 9175 4440 9205
rect 4410 9105 4440 9135
rect 4610 9175 4640 9205
rect 4610 9105 4640 9135
rect 4810 9175 4840 9205
rect 4810 9105 4840 9135
rect 5010 9175 5040 9205
rect 5010 9105 5040 9135
rect 5210 9175 5240 9205
rect 5210 9105 5240 9135
rect 5410 9175 5440 9205
rect 5410 9105 5440 9135
rect 5610 9175 5640 9205
rect 5610 9105 5640 9135
rect 5810 9175 5840 9205
rect 5810 9105 5840 9135
rect 6010 9175 6040 9205
rect 6010 9105 6040 9135
rect 6210 9175 6240 9205
rect 6210 9105 6240 9135
rect 6410 9175 6440 9205
rect 6410 9105 6440 9135
rect -190 8990 -160 9020
rect -190 8920 -160 8950
rect 10 8990 40 9020
rect 10 8920 40 8950
rect 210 8990 240 9020
rect 210 8920 240 8950
rect 410 8990 440 9020
rect 410 8920 440 8950
rect 610 8990 640 9020
rect 610 8920 640 8950
rect 810 8990 840 9020
rect 810 8920 840 8950
rect 1010 8990 1040 9020
rect 1010 8920 1040 8950
rect 1210 8990 1240 9020
rect 1210 8920 1240 8950
rect 1410 8990 1440 9020
rect 1410 8920 1440 8950
rect 1610 8990 1640 9020
rect 1610 8920 1640 8950
rect 1810 8990 1840 9020
rect 1810 8920 1840 8950
rect 2010 8990 2040 9020
rect 2010 8920 2040 8950
rect 2210 8990 2240 9020
rect 2210 8920 2240 8950
rect 2410 8990 2440 9020
rect 2410 8920 2440 8950
rect 2610 8990 2640 9020
rect 2610 8920 2640 8950
rect 2810 8990 2840 9020
rect 2810 8920 2840 8950
rect 3010 8990 3040 9020
rect 3010 8920 3040 8950
rect 3210 8990 3240 9020
rect 3210 8920 3240 8950
rect 3410 8990 3440 9020
rect 3410 8920 3440 8950
rect 3610 8990 3640 9020
rect 3610 8920 3640 8950
rect 3810 8990 3840 9020
rect 3810 8920 3840 8950
rect 4010 8990 4040 9020
rect 4010 8920 4040 8950
rect 4210 8990 4240 9020
rect 4210 8920 4240 8950
rect 4410 8990 4440 9020
rect 4410 8920 4440 8950
rect 4610 8990 4640 9020
rect 4610 8920 4640 8950
rect 4810 8990 4840 9020
rect 4810 8920 4840 8950
rect 5010 8990 5040 9020
rect 5010 8920 5040 8950
rect 5210 8990 5240 9020
rect 5210 8920 5240 8950
rect 5410 8990 5440 9020
rect 5410 8920 5440 8950
rect 5610 8990 5640 9020
rect 5610 8920 5640 8950
rect 5810 8990 5840 9020
rect 5810 8920 5840 8950
rect 6010 8990 6040 9020
rect 6010 8920 6040 8950
rect 6210 8990 6240 9020
rect 6210 8920 6240 8950
rect 6410 8990 6440 9020
rect 6410 8920 6440 8950
rect -190 8805 -160 8835
rect -190 8735 -160 8765
rect 10 8805 40 8835
rect 10 8735 40 8765
rect 210 8805 240 8835
rect 210 8735 240 8765
rect 410 8805 440 8835
rect 410 8735 440 8765
rect 610 8805 640 8835
rect 610 8735 640 8765
rect 810 8805 840 8835
rect 810 8735 840 8765
rect 1010 8805 1040 8835
rect 1010 8735 1040 8765
rect 1210 8805 1240 8835
rect 1210 8735 1240 8765
rect 1410 8805 1440 8835
rect 1410 8735 1440 8765
rect 1610 8805 1640 8835
rect 1610 8735 1640 8765
rect 1810 8805 1840 8835
rect 1810 8735 1840 8765
rect 2010 8805 2040 8835
rect 2010 8735 2040 8765
rect 2210 8805 2240 8835
rect 2210 8735 2240 8765
rect 2410 8805 2440 8835
rect 2410 8735 2440 8765
rect 2610 8805 2640 8835
rect 2610 8735 2640 8765
rect 2810 8805 2840 8835
rect 2810 8735 2840 8765
rect 3010 8805 3040 8835
rect 3010 8735 3040 8765
rect 3210 8805 3240 8835
rect 3210 8735 3240 8765
rect 3410 8805 3440 8835
rect 3410 8735 3440 8765
rect 3610 8805 3640 8835
rect 3610 8735 3640 8765
rect 3810 8805 3840 8835
rect 3810 8735 3840 8765
rect 4010 8805 4040 8835
rect 4010 8735 4040 8765
rect 4210 8805 4240 8835
rect 4210 8735 4240 8765
rect 4410 8805 4440 8835
rect 4410 8735 4440 8765
rect 4610 8805 4640 8835
rect 4610 8735 4640 8765
rect 4810 8805 4840 8835
rect 4810 8735 4840 8765
rect 5010 8805 5040 8835
rect 5010 8735 5040 8765
rect 5210 8805 5240 8835
rect 5210 8735 5240 8765
rect 5410 8805 5440 8835
rect 5410 8735 5440 8765
rect 5610 8805 5640 8835
rect 5610 8735 5640 8765
rect 5810 8805 5840 8835
rect 5810 8735 5840 8765
rect 6010 8805 6040 8835
rect 6010 8735 6040 8765
rect 6210 8805 6240 8835
rect 6210 8735 6240 8765
rect 6410 8805 6440 8835
rect 6410 8735 6440 8765
rect -190 8620 -160 8650
rect -190 8550 -160 8580
rect 10 8620 40 8650
rect 10 8550 40 8580
rect 210 8620 240 8650
rect 210 8550 240 8580
rect 410 8620 440 8650
rect 410 8550 440 8580
rect 610 8620 640 8650
rect 610 8550 640 8580
rect 810 8620 840 8650
rect 810 8550 840 8580
rect 1010 8620 1040 8650
rect 1010 8550 1040 8580
rect 1210 8620 1240 8650
rect 1210 8550 1240 8580
rect 1410 8620 1440 8650
rect 1410 8550 1440 8580
rect 1610 8620 1640 8650
rect 1610 8550 1640 8580
rect 1810 8620 1840 8650
rect 1810 8550 1840 8580
rect 2010 8620 2040 8650
rect 2010 8550 2040 8580
rect 2210 8620 2240 8650
rect 2210 8550 2240 8580
rect 2410 8620 2440 8650
rect 2410 8550 2440 8580
rect 2610 8620 2640 8650
rect 2610 8550 2640 8580
rect 2810 8620 2840 8650
rect 2810 8550 2840 8580
rect 3010 8620 3040 8650
rect 3010 8550 3040 8580
rect 3210 8620 3240 8650
rect 3210 8550 3240 8580
rect 3410 8620 3440 8650
rect 3410 8550 3440 8580
rect 3610 8620 3640 8650
rect 3610 8550 3640 8580
rect 3810 8620 3840 8650
rect 3810 8550 3840 8580
rect 4010 8620 4040 8650
rect 4010 8550 4040 8580
rect 4210 8620 4240 8650
rect 4210 8550 4240 8580
rect 4410 8620 4440 8650
rect 4410 8550 4440 8580
rect 4610 8620 4640 8650
rect 4610 8550 4640 8580
rect 4810 8620 4840 8650
rect 4810 8550 4840 8580
rect 5010 8620 5040 8650
rect 5010 8550 5040 8580
rect 5210 8620 5240 8650
rect 5210 8550 5240 8580
rect 5410 8620 5440 8650
rect 5410 8550 5440 8580
rect 5610 8620 5640 8650
rect 5610 8550 5640 8580
rect 5810 8620 5840 8650
rect 5810 8550 5840 8580
rect 6010 8620 6040 8650
rect 6010 8550 6040 8580
rect 6210 8620 6240 8650
rect 6210 8550 6240 8580
rect 6410 8620 6440 8650
rect 6410 8550 6440 8580
rect -190 8435 -160 8465
rect -190 8365 -160 8395
rect 10 8435 40 8465
rect 10 8365 40 8395
rect 210 8435 240 8465
rect 210 8365 240 8395
rect 410 8435 440 8465
rect 410 8365 440 8395
rect 610 8435 640 8465
rect 610 8365 640 8395
rect 810 8435 840 8465
rect 810 8365 840 8395
rect 1010 8435 1040 8465
rect 1010 8365 1040 8395
rect 1210 8435 1240 8465
rect 1210 8365 1240 8395
rect 1410 8435 1440 8465
rect 1410 8365 1440 8395
rect 1610 8435 1640 8465
rect 1610 8365 1640 8395
rect 1810 8435 1840 8465
rect 1810 8365 1840 8395
rect 2010 8435 2040 8465
rect 2010 8365 2040 8395
rect 2210 8435 2240 8465
rect 2210 8365 2240 8395
rect 2410 8435 2440 8465
rect 2410 8365 2440 8395
rect 2610 8435 2640 8465
rect 2610 8365 2640 8395
rect 2810 8435 2840 8465
rect 2810 8365 2840 8395
rect 3010 8435 3040 8465
rect 3010 8365 3040 8395
rect 3210 8435 3240 8465
rect 3210 8365 3240 8395
rect 3410 8435 3440 8465
rect 3410 8365 3440 8395
rect 3610 8435 3640 8465
rect 3610 8365 3640 8395
rect 3810 8435 3840 8465
rect 3810 8365 3840 8395
rect 4010 8435 4040 8465
rect 4010 8365 4040 8395
rect 4210 8435 4240 8465
rect 4210 8365 4240 8395
rect 4410 8435 4440 8465
rect 4410 8365 4440 8395
rect 4610 8435 4640 8465
rect 4610 8365 4640 8395
rect 4810 8435 4840 8465
rect 4810 8365 4840 8395
rect 5010 8435 5040 8465
rect 5010 8365 5040 8395
rect 5210 8435 5240 8465
rect 5210 8365 5240 8395
rect 5410 8435 5440 8465
rect 5410 8365 5440 8395
rect 5610 8435 5640 8465
rect 5610 8365 5640 8395
rect 5810 8435 5840 8465
rect 5810 8365 5840 8395
rect 6010 8435 6040 8465
rect 6010 8365 6040 8395
rect 6210 8435 6240 8465
rect 6210 8365 6240 8395
rect 6410 8435 6440 8465
rect 6410 8365 6440 8395
rect -190 8250 -160 8280
rect -190 8180 -160 8210
rect 10 8250 40 8280
rect 10 8180 40 8210
rect 210 8250 240 8280
rect 210 8180 240 8210
rect 410 8250 440 8280
rect 410 8180 440 8210
rect 610 8250 640 8280
rect 610 8180 640 8210
rect 810 8250 840 8280
rect 810 8180 840 8210
rect 1010 8250 1040 8280
rect 1010 8180 1040 8210
rect 1210 8250 1240 8280
rect 1210 8180 1240 8210
rect 1410 8250 1440 8280
rect 1410 8180 1440 8210
rect 1610 8250 1640 8280
rect 1610 8180 1640 8210
rect 1810 8250 1840 8280
rect 1810 8180 1840 8210
rect 2010 8250 2040 8280
rect 2010 8180 2040 8210
rect 2210 8250 2240 8280
rect 2210 8180 2240 8210
rect 2410 8250 2440 8280
rect 2410 8180 2440 8210
rect 2610 8250 2640 8280
rect 2610 8180 2640 8210
rect 2810 8250 2840 8280
rect 2810 8180 2840 8210
rect 3010 8250 3040 8280
rect 3010 8180 3040 8210
rect 3210 8250 3240 8280
rect 3210 8180 3240 8210
rect 3410 8250 3440 8280
rect 3410 8180 3440 8210
rect 3610 8250 3640 8280
rect 3610 8180 3640 8210
rect 3810 8250 3840 8280
rect 3810 8180 3840 8210
rect 4010 8250 4040 8280
rect 4010 8180 4040 8210
rect 4210 8250 4240 8280
rect 4210 8180 4240 8210
rect 4410 8250 4440 8280
rect 4410 8180 4440 8210
rect 4610 8250 4640 8280
rect 4610 8180 4640 8210
rect 4810 8250 4840 8280
rect 4810 8180 4840 8210
rect 5010 8250 5040 8280
rect 5010 8180 5040 8210
rect 5210 8250 5240 8280
rect 5210 8180 5240 8210
rect 5410 8250 5440 8280
rect 5410 8180 5440 8210
rect 5610 8250 5640 8280
rect 5610 8180 5640 8210
rect 5810 8250 5840 8280
rect 5810 8180 5840 8210
rect 6010 8250 6040 8280
rect 6010 8180 6040 8210
rect 6210 8250 6240 8280
rect 6210 8180 6240 8210
rect 6410 8250 6440 8280
rect 6410 8180 6440 8210
rect -190 8065 -160 8095
rect -190 7995 -160 8025
rect 10 8065 40 8095
rect 10 7995 40 8025
rect 210 8065 240 8095
rect 210 7995 240 8025
rect 410 8065 440 8095
rect 410 7995 440 8025
rect 610 8065 640 8095
rect 610 7995 640 8025
rect 810 8065 840 8095
rect 810 7995 840 8025
rect 1010 8065 1040 8095
rect 1010 7995 1040 8025
rect 1210 8065 1240 8095
rect 1210 7995 1240 8025
rect 1410 8065 1440 8095
rect 1410 7995 1440 8025
rect 1610 8065 1640 8095
rect 1610 7995 1640 8025
rect 1810 8065 1840 8095
rect 1810 7995 1840 8025
rect 2010 8065 2040 8095
rect 2010 7995 2040 8025
rect 2210 8065 2240 8095
rect 2210 7995 2240 8025
rect 2410 8065 2440 8095
rect 2410 7995 2440 8025
rect 2610 8065 2640 8095
rect 2610 7995 2640 8025
rect 2810 8065 2840 8095
rect 2810 7995 2840 8025
rect 3010 8065 3040 8095
rect 3010 7995 3040 8025
rect 3210 8065 3240 8095
rect 3210 7995 3240 8025
rect 3410 8065 3440 8095
rect 3410 7995 3440 8025
rect 3610 8065 3640 8095
rect 3610 7995 3640 8025
rect 3810 8065 3840 8095
rect 3810 7995 3840 8025
rect 4010 8065 4040 8095
rect 4010 7995 4040 8025
rect 4210 8065 4240 8095
rect 4210 7995 4240 8025
rect 4410 8065 4440 8095
rect 4410 7995 4440 8025
rect 4610 8065 4640 8095
rect 4610 7995 4640 8025
rect 4810 8065 4840 8095
rect 4810 7995 4840 8025
rect 5010 8065 5040 8095
rect 5010 7995 5040 8025
rect 5210 8065 5240 8095
rect 5210 7995 5240 8025
rect 5410 8065 5440 8095
rect 5410 7995 5440 8025
rect 5610 8065 5640 8095
rect 5610 7995 5640 8025
rect 5810 8065 5840 8095
rect 5810 7995 5840 8025
rect 6010 8065 6040 8095
rect 6010 7995 6040 8025
rect 6210 8065 6240 8095
rect 6210 7995 6240 8025
rect 6410 8065 6440 8095
rect 6410 7995 6440 8025
rect -190 7880 -160 7910
rect -190 7810 -160 7840
rect 10 7880 40 7910
rect 10 7810 40 7840
rect 210 7880 240 7910
rect 210 7810 240 7840
rect 410 7880 440 7910
rect 410 7810 440 7840
rect 610 7880 640 7910
rect 610 7810 640 7840
rect 810 7880 840 7910
rect 810 7810 840 7840
rect 1010 7880 1040 7910
rect 1010 7810 1040 7840
rect 1210 7880 1240 7910
rect 1210 7810 1240 7840
rect 1410 7880 1440 7910
rect 1410 7810 1440 7840
rect 1610 7880 1640 7910
rect 1610 7810 1640 7840
rect 1810 7880 1840 7910
rect 1810 7810 1840 7840
rect 2010 7880 2040 7910
rect 2010 7810 2040 7840
rect 2210 7880 2240 7910
rect 2210 7810 2240 7840
rect 2410 7880 2440 7910
rect 2410 7810 2440 7840
rect 2610 7880 2640 7910
rect 2610 7810 2640 7840
rect 2810 7880 2840 7910
rect 2810 7810 2840 7840
rect 3010 7880 3040 7910
rect 3010 7810 3040 7840
rect 3210 7880 3240 7910
rect 3210 7810 3240 7840
rect 3410 7880 3440 7910
rect 3410 7810 3440 7840
rect 3610 7880 3640 7910
rect 3610 7810 3640 7840
rect 3810 7880 3840 7910
rect 3810 7810 3840 7840
rect 4010 7880 4040 7910
rect 4010 7810 4040 7840
rect 4210 7880 4240 7910
rect 4210 7810 4240 7840
rect 4410 7880 4440 7910
rect 4410 7810 4440 7840
rect 4610 7880 4640 7910
rect 4610 7810 4640 7840
rect 4810 7880 4840 7910
rect 4810 7810 4840 7840
rect 5010 7880 5040 7910
rect 5010 7810 5040 7840
rect 5210 7880 5240 7910
rect 5210 7810 5240 7840
rect 5410 7880 5440 7910
rect 5410 7810 5440 7840
rect 5610 7880 5640 7910
rect 5610 7810 5640 7840
rect 5810 7880 5840 7910
rect 5810 7810 5840 7840
rect 6010 7880 6040 7910
rect 6010 7810 6040 7840
rect 6210 7880 6240 7910
rect 6210 7810 6240 7840
rect 6410 7880 6440 7910
rect 6410 7810 6440 7840
rect -190 7695 -160 7725
rect -190 7625 -160 7655
rect 10 7695 40 7725
rect 10 7625 40 7655
rect 210 7695 240 7725
rect 210 7625 240 7655
rect 410 7695 440 7725
rect 410 7625 440 7655
rect 610 7695 640 7725
rect 610 7625 640 7655
rect 810 7695 840 7725
rect 810 7625 840 7655
rect 1010 7695 1040 7725
rect 1010 7625 1040 7655
rect 1210 7695 1240 7725
rect 1210 7625 1240 7655
rect 1410 7695 1440 7725
rect 1410 7625 1440 7655
rect 1610 7695 1640 7725
rect 1610 7625 1640 7655
rect 1810 7695 1840 7725
rect 1810 7625 1840 7655
rect 2010 7695 2040 7725
rect 2010 7625 2040 7655
rect 2210 7695 2240 7725
rect 2210 7625 2240 7655
rect 2410 7695 2440 7725
rect 2410 7625 2440 7655
rect 2610 7695 2640 7725
rect 2610 7625 2640 7655
rect 2810 7695 2840 7725
rect 2810 7625 2840 7655
rect 3010 7695 3040 7725
rect 3010 7625 3040 7655
rect 3210 7695 3240 7725
rect 3210 7625 3240 7655
rect 3410 7695 3440 7725
rect 3410 7625 3440 7655
rect 3610 7695 3640 7725
rect 3610 7625 3640 7655
rect 3810 7695 3840 7725
rect 3810 7625 3840 7655
rect 4010 7695 4040 7725
rect 4010 7625 4040 7655
rect 4210 7695 4240 7725
rect 4210 7625 4240 7655
rect 4410 7695 4440 7725
rect 4410 7625 4440 7655
rect 4610 7695 4640 7725
rect 4610 7625 4640 7655
rect 4810 7695 4840 7725
rect 4810 7625 4840 7655
rect 5010 7695 5040 7725
rect 5010 7625 5040 7655
rect 5210 7695 5240 7725
rect 5210 7625 5240 7655
rect 5410 7695 5440 7725
rect 5410 7625 5440 7655
rect 5610 7695 5640 7725
rect 5610 7625 5640 7655
rect 5810 7695 5840 7725
rect 5810 7625 5840 7655
rect 6010 7695 6040 7725
rect 6010 7625 6040 7655
rect 6210 7695 6240 7725
rect 6210 7625 6240 7655
rect 6410 7695 6440 7725
rect 6410 7625 6440 7655
rect -190 7510 -160 7540
rect -190 7440 -160 7470
rect 10 7510 40 7540
rect 10 7440 40 7470
rect 210 7510 240 7540
rect 210 7440 240 7470
rect 410 7510 440 7540
rect 410 7440 440 7470
rect 610 7510 640 7540
rect 610 7440 640 7470
rect 810 7510 840 7540
rect 810 7440 840 7470
rect 1010 7510 1040 7540
rect 1010 7440 1040 7470
rect 1210 7510 1240 7540
rect 1210 7440 1240 7470
rect 1410 7510 1440 7540
rect 1410 7440 1440 7470
rect 1610 7510 1640 7540
rect 1610 7440 1640 7470
rect 1810 7510 1840 7540
rect 1810 7440 1840 7470
rect 2010 7510 2040 7540
rect 2010 7440 2040 7470
rect 2210 7510 2240 7540
rect 2210 7440 2240 7470
rect 2410 7510 2440 7540
rect 2410 7440 2440 7470
rect 2610 7510 2640 7540
rect 2610 7440 2640 7470
rect 2810 7510 2840 7540
rect 2810 7440 2840 7470
rect 3010 7510 3040 7540
rect 3010 7440 3040 7470
rect 3210 7510 3240 7540
rect 3210 7440 3240 7470
rect 3410 7510 3440 7540
rect 3410 7440 3440 7470
rect 3610 7510 3640 7540
rect 3610 7440 3640 7470
rect 3810 7510 3840 7540
rect 3810 7440 3840 7470
rect 4010 7510 4040 7540
rect 4010 7440 4040 7470
rect 4210 7510 4240 7540
rect 4210 7440 4240 7470
rect 4410 7510 4440 7540
rect 4410 7440 4440 7470
rect 4610 7510 4640 7540
rect 4610 7440 4640 7470
rect 4810 7510 4840 7540
rect 4810 7440 4840 7470
rect 5010 7510 5040 7540
rect 5010 7440 5040 7470
rect 5210 7510 5240 7540
rect 5210 7440 5240 7470
rect 5410 7510 5440 7540
rect 5410 7440 5440 7470
rect 5610 7510 5640 7540
rect 5610 7440 5640 7470
rect 5810 7510 5840 7540
rect 5810 7440 5840 7470
rect 6010 7510 6040 7540
rect 6010 7440 6040 7470
rect 6210 7510 6240 7540
rect 6210 7440 6240 7470
rect 6410 7510 6440 7540
rect 6410 7440 6440 7470
rect -190 7325 -160 7355
rect -190 7255 -160 7285
rect 10 7325 40 7355
rect 10 7255 40 7285
rect 210 7325 240 7355
rect 210 7255 240 7285
rect 410 7325 440 7355
rect 410 7255 440 7285
rect 610 7325 640 7355
rect 610 7255 640 7285
rect 810 7325 840 7355
rect 810 7255 840 7285
rect 1010 7325 1040 7355
rect 1010 7255 1040 7285
rect 1210 7325 1240 7355
rect 1210 7255 1240 7285
rect 1410 7325 1440 7355
rect 1410 7255 1440 7285
rect 1610 7325 1640 7355
rect 1610 7255 1640 7285
rect 1810 7325 1840 7355
rect 1810 7255 1840 7285
rect 2010 7325 2040 7355
rect 2010 7255 2040 7285
rect 2210 7325 2240 7355
rect 2210 7255 2240 7285
rect 2410 7325 2440 7355
rect 2410 7255 2440 7285
rect 2610 7325 2640 7355
rect 2610 7255 2640 7285
rect 2810 7325 2840 7355
rect 2810 7255 2840 7285
rect 3010 7325 3040 7355
rect 3010 7255 3040 7285
rect 3210 7325 3240 7355
rect 3210 7255 3240 7285
rect 3410 7325 3440 7355
rect 3410 7255 3440 7285
rect 3610 7325 3640 7355
rect 3610 7255 3640 7285
rect 3810 7325 3840 7355
rect 3810 7255 3840 7285
rect 4010 7325 4040 7355
rect 4010 7255 4040 7285
rect 4210 7325 4240 7355
rect 4210 7255 4240 7285
rect 4410 7325 4440 7355
rect 4410 7255 4440 7285
rect 4610 7325 4640 7355
rect 4610 7255 4640 7285
rect 4810 7325 4840 7355
rect 4810 7255 4840 7285
rect 5010 7325 5040 7355
rect 5010 7255 5040 7285
rect 5210 7325 5240 7355
rect 5210 7255 5240 7285
rect 5410 7325 5440 7355
rect 5410 7255 5440 7285
rect 5610 7325 5640 7355
rect 5610 7255 5640 7285
rect 5810 7325 5840 7355
rect 5810 7255 5840 7285
rect 6010 7325 6040 7355
rect 6010 7255 6040 7285
rect 6210 7325 6240 7355
rect 6210 7255 6240 7285
rect 6410 7325 6440 7355
rect 6410 7255 6440 7285
rect -190 7140 -160 7170
rect -190 7070 -160 7100
rect 10 7140 40 7170
rect 10 7070 40 7100
rect 210 7140 240 7170
rect 210 7070 240 7100
rect 410 7140 440 7170
rect 410 7070 440 7100
rect 610 7140 640 7170
rect 610 7070 640 7100
rect 810 7140 840 7170
rect 810 7070 840 7100
rect 1010 7140 1040 7170
rect 1010 7070 1040 7100
rect 1210 7140 1240 7170
rect 1210 7070 1240 7100
rect 1410 7140 1440 7170
rect 1410 7070 1440 7100
rect 1610 7140 1640 7170
rect 1610 7070 1640 7100
rect 1810 7140 1840 7170
rect 1810 7070 1840 7100
rect 2010 7140 2040 7170
rect 2010 7070 2040 7100
rect 2210 7140 2240 7170
rect 2210 7070 2240 7100
rect 2410 7140 2440 7170
rect 2410 7070 2440 7100
rect 2610 7140 2640 7170
rect 2610 7070 2640 7100
rect 2810 7140 2840 7170
rect 2810 7070 2840 7100
rect 3010 7140 3040 7170
rect 3010 7070 3040 7100
rect 3210 7140 3240 7170
rect 3210 7070 3240 7100
rect 3410 7140 3440 7170
rect 3410 7070 3440 7100
rect 3610 7140 3640 7170
rect 3610 7070 3640 7100
rect 3810 7140 3840 7170
rect 3810 7070 3840 7100
rect 4010 7140 4040 7170
rect 4010 7070 4040 7100
rect 4210 7140 4240 7170
rect 4210 7070 4240 7100
rect 4410 7140 4440 7170
rect 4410 7070 4440 7100
rect 4610 7140 4640 7170
rect 4610 7070 4640 7100
rect 4810 7140 4840 7170
rect 4810 7070 4840 7100
rect 5010 7140 5040 7170
rect 5010 7070 5040 7100
rect 5210 7140 5240 7170
rect 5210 7070 5240 7100
rect 5410 7140 5440 7170
rect 5410 7070 5440 7100
rect 5610 7140 5640 7170
rect 5610 7070 5640 7100
rect 5810 7140 5840 7170
rect 5810 7070 5840 7100
rect 6010 7140 6040 7170
rect 6010 7070 6040 7100
rect 6210 7140 6240 7170
rect 6210 7070 6240 7100
rect 6410 7140 6440 7170
rect 6410 7070 6440 7100
rect -190 6955 -160 6985
rect -190 6885 -160 6915
rect 10 6955 40 6985
rect 10 6885 40 6915
rect 210 6955 240 6985
rect 210 6885 240 6915
rect 410 6955 440 6985
rect 410 6885 440 6915
rect 610 6955 640 6985
rect 610 6885 640 6915
rect 810 6955 840 6985
rect 810 6885 840 6915
rect 1010 6955 1040 6985
rect 1010 6885 1040 6915
rect 1210 6955 1240 6985
rect 1210 6885 1240 6915
rect 1410 6955 1440 6985
rect 1410 6885 1440 6915
rect 1610 6955 1640 6985
rect 1610 6885 1640 6915
rect 1810 6955 1840 6985
rect 1810 6885 1840 6915
rect 2010 6955 2040 6985
rect 2010 6885 2040 6915
rect 2210 6955 2240 6985
rect 2210 6885 2240 6915
rect 2410 6955 2440 6985
rect 2410 6885 2440 6915
rect 2610 6955 2640 6985
rect 2610 6885 2640 6915
rect 2810 6955 2840 6985
rect 2810 6885 2840 6915
rect 3010 6955 3040 6985
rect 3010 6885 3040 6915
rect 3210 6955 3240 6985
rect 3210 6885 3240 6915
rect 3410 6955 3440 6985
rect 3410 6885 3440 6915
rect 3610 6955 3640 6985
rect 3610 6885 3640 6915
rect 3810 6955 3840 6985
rect 3810 6885 3840 6915
rect 4010 6955 4040 6985
rect 4010 6885 4040 6915
rect 4210 6955 4240 6985
rect 4210 6885 4240 6915
rect 4410 6955 4440 6985
rect 4410 6885 4440 6915
rect 4610 6955 4640 6985
rect 4610 6885 4640 6915
rect 4810 6955 4840 6985
rect 4810 6885 4840 6915
rect 5010 6955 5040 6985
rect 5010 6885 5040 6915
rect 5210 6955 5240 6985
rect 5210 6885 5240 6915
rect 5410 6955 5440 6985
rect 5410 6885 5440 6915
rect 5610 6955 5640 6985
rect 5610 6885 5640 6915
rect 5810 6955 5840 6985
rect 5810 6885 5840 6915
rect 6010 6955 6040 6985
rect 6010 6885 6040 6915
rect 6210 6955 6240 6985
rect 6210 6885 6240 6915
rect 6410 6955 6440 6985
rect 6410 6885 6440 6915
rect -190 6770 -160 6800
rect -190 6700 -160 6730
rect 10 6770 40 6800
rect 10 6700 40 6730
rect 210 6770 240 6800
rect 210 6700 240 6730
rect 410 6770 440 6800
rect 410 6700 440 6730
rect 610 6770 640 6800
rect 610 6700 640 6730
rect 810 6770 840 6800
rect 810 6700 840 6730
rect 1010 6770 1040 6800
rect 1010 6700 1040 6730
rect 1210 6770 1240 6800
rect 1210 6700 1240 6730
rect 1410 6770 1440 6800
rect 1410 6700 1440 6730
rect 1610 6770 1640 6800
rect 1610 6700 1640 6730
rect 1810 6770 1840 6800
rect 1810 6700 1840 6730
rect 2010 6770 2040 6800
rect 2010 6700 2040 6730
rect 2210 6770 2240 6800
rect 2210 6700 2240 6730
rect 2410 6770 2440 6800
rect 2410 6700 2440 6730
rect 2610 6770 2640 6800
rect 2610 6700 2640 6730
rect 2810 6770 2840 6800
rect 2810 6700 2840 6730
rect 3010 6770 3040 6800
rect 3010 6700 3040 6730
rect 3210 6770 3240 6800
rect 3210 6700 3240 6730
rect 3410 6770 3440 6800
rect 3410 6700 3440 6730
rect 3610 6770 3640 6800
rect 3610 6700 3640 6730
rect 3810 6770 3840 6800
rect 3810 6700 3840 6730
rect 4010 6770 4040 6800
rect 4010 6700 4040 6730
rect 4210 6770 4240 6800
rect 4210 6700 4240 6730
rect 4410 6770 4440 6800
rect 4410 6700 4440 6730
rect 4610 6770 4640 6800
rect 4610 6700 4640 6730
rect 4810 6770 4840 6800
rect 4810 6700 4840 6730
rect 5010 6770 5040 6800
rect 5010 6700 5040 6730
rect 5210 6770 5240 6800
rect 5210 6700 5240 6730
rect 5410 6770 5440 6800
rect 5410 6700 5440 6730
rect 5610 6770 5640 6800
rect 5610 6700 5640 6730
rect 5810 6770 5840 6800
rect 5810 6700 5840 6730
rect 6010 6770 6040 6800
rect 6010 6700 6040 6730
rect 6210 6770 6240 6800
rect 6210 6700 6240 6730
rect 6410 6770 6440 6800
rect 6410 6700 6440 6730
rect -190 6585 -160 6615
rect -190 6515 -160 6545
rect 10 6585 40 6615
rect 10 6515 40 6545
rect 210 6585 240 6615
rect 210 6515 240 6545
rect 410 6585 440 6615
rect 410 6515 440 6545
rect 610 6585 640 6615
rect 610 6515 640 6545
rect 810 6585 840 6615
rect 810 6515 840 6545
rect 1010 6585 1040 6615
rect 1010 6515 1040 6545
rect 1210 6585 1240 6615
rect 1210 6515 1240 6545
rect 1410 6585 1440 6615
rect 1410 6515 1440 6545
rect 1610 6585 1640 6615
rect 1610 6515 1640 6545
rect 1810 6585 1840 6615
rect 1810 6515 1840 6545
rect 2010 6585 2040 6615
rect 2010 6515 2040 6545
rect 2210 6585 2240 6615
rect 2210 6515 2240 6545
rect 2410 6585 2440 6615
rect 2410 6515 2440 6545
rect 2610 6585 2640 6615
rect 2610 6515 2640 6545
rect 2810 6585 2840 6615
rect 2810 6515 2840 6545
rect 3010 6585 3040 6615
rect 3010 6515 3040 6545
rect 3210 6585 3240 6615
rect 3210 6515 3240 6545
rect 3410 6585 3440 6615
rect 3410 6515 3440 6545
rect 3610 6585 3640 6615
rect 3610 6515 3640 6545
rect 3810 6585 3840 6615
rect 3810 6515 3840 6545
rect 4010 6585 4040 6615
rect 4010 6515 4040 6545
rect 4210 6585 4240 6615
rect 4210 6515 4240 6545
rect 4410 6585 4440 6615
rect 4410 6515 4440 6545
rect 4610 6585 4640 6615
rect 4610 6515 4640 6545
rect 4810 6585 4840 6615
rect 4810 6515 4840 6545
rect 5010 6585 5040 6615
rect 5010 6515 5040 6545
rect 5210 6585 5240 6615
rect 5210 6515 5240 6545
rect 5410 6585 5440 6615
rect 5410 6515 5440 6545
rect 5610 6585 5640 6615
rect 5610 6515 5640 6545
rect 5810 6585 5840 6615
rect 5810 6515 5840 6545
rect 6010 6585 6040 6615
rect 6010 6515 6040 6545
rect 6210 6585 6240 6615
rect 6210 6515 6240 6545
rect 6410 6585 6440 6615
rect 6410 6515 6440 6545
rect -190 6400 -160 6430
rect -190 6330 -160 6360
rect 10 6400 40 6430
rect 10 6330 40 6360
rect 210 6400 240 6430
rect 210 6330 240 6360
rect 410 6400 440 6430
rect 410 6330 440 6360
rect 610 6400 640 6430
rect 610 6330 640 6360
rect 810 6400 840 6430
rect 810 6330 840 6360
rect 1010 6400 1040 6430
rect 1010 6330 1040 6360
rect 1210 6400 1240 6430
rect 1210 6330 1240 6360
rect 1410 6400 1440 6430
rect 1410 6330 1440 6360
rect 1610 6400 1640 6430
rect 1610 6330 1640 6360
rect 1810 6400 1840 6430
rect 1810 6330 1840 6360
rect 2010 6400 2040 6430
rect 2010 6330 2040 6360
rect 2210 6400 2240 6430
rect 2210 6330 2240 6360
rect 2410 6400 2440 6430
rect 2410 6330 2440 6360
rect 2610 6400 2640 6430
rect 2610 6330 2640 6360
rect 2810 6400 2840 6430
rect 2810 6330 2840 6360
rect 3010 6400 3040 6430
rect 3010 6330 3040 6360
rect 3210 6400 3240 6430
rect 3210 6330 3240 6360
rect 3410 6400 3440 6430
rect 3410 6330 3440 6360
rect 3610 6400 3640 6430
rect 3610 6330 3640 6360
rect 3810 6400 3840 6430
rect 3810 6330 3840 6360
rect 4010 6400 4040 6430
rect 4010 6330 4040 6360
rect 4210 6400 4240 6430
rect 4210 6330 4240 6360
rect 4410 6400 4440 6430
rect 4410 6330 4440 6360
rect 4610 6400 4640 6430
rect 4610 6330 4640 6360
rect 4810 6400 4840 6430
rect 4810 6330 4840 6360
rect 5010 6400 5040 6430
rect 5010 6330 5040 6360
rect 5210 6400 5240 6430
rect 5210 6330 5240 6360
rect 5410 6400 5440 6430
rect 5410 6330 5440 6360
rect 5610 6400 5640 6430
rect 5610 6330 5640 6360
rect 5810 6400 5840 6430
rect 5810 6330 5840 6360
rect 6010 6400 6040 6430
rect 6010 6330 6040 6360
rect 6210 6400 6240 6430
rect 6210 6330 6240 6360
rect 6410 6400 6440 6430
rect 6410 6330 6440 6360
rect -190 6215 -160 6245
rect -190 6145 -160 6175
rect 10 6215 40 6245
rect 10 6145 40 6175
rect 210 6215 240 6245
rect 210 6145 240 6175
rect 410 6215 440 6245
rect 410 6145 440 6175
rect 610 6215 640 6245
rect 610 6145 640 6175
rect 810 6215 840 6245
rect 810 6145 840 6175
rect 1010 6215 1040 6245
rect 1010 6145 1040 6175
rect 1210 6215 1240 6245
rect 1210 6145 1240 6175
rect 1410 6215 1440 6245
rect 1410 6145 1440 6175
rect 1610 6215 1640 6245
rect 1610 6145 1640 6175
rect 1810 6215 1840 6245
rect 1810 6145 1840 6175
rect 2010 6215 2040 6245
rect 2010 6145 2040 6175
rect 2210 6215 2240 6245
rect 2210 6145 2240 6175
rect 2410 6215 2440 6245
rect 2410 6145 2440 6175
rect 2610 6215 2640 6245
rect 2610 6145 2640 6175
rect 2810 6215 2840 6245
rect 2810 6145 2840 6175
rect 3010 6215 3040 6245
rect 3010 6145 3040 6175
rect 3210 6215 3240 6245
rect 3210 6145 3240 6175
rect 3410 6215 3440 6245
rect 3410 6145 3440 6175
rect 3610 6215 3640 6245
rect 3610 6145 3640 6175
rect 3810 6215 3840 6245
rect 3810 6145 3840 6175
rect 4010 6215 4040 6245
rect 4010 6145 4040 6175
rect 4210 6215 4240 6245
rect 4210 6145 4240 6175
rect 4410 6215 4440 6245
rect 4410 6145 4440 6175
rect 4610 6215 4640 6245
rect 4610 6145 4640 6175
rect 4810 6215 4840 6245
rect 4810 6145 4840 6175
rect 5010 6215 5040 6245
rect 5010 6145 5040 6175
rect 5210 6215 5240 6245
rect 5210 6145 5240 6175
rect 5410 6215 5440 6245
rect 5410 6145 5440 6175
rect 5610 6215 5640 6245
rect 5610 6145 5640 6175
rect 5810 6215 5840 6245
rect 5810 6145 5840 6175
rect 6010 6215 6040 6245
rect 6010 6145 6040 6175
rect 6210 6215 6240 6245
rect 6210 6145 6240 6175
rect 6410 6215 6440 6245
rect 6410 6145 6440 6175
rect -190 6030 -160 6060
rect -190 5960 -160 5990
rect 10 6030 40 6060
rect 10 5960 40 5990
rect 210 6030 240 6060
rect 210 5960 240 5990
rect 410 6030 440 6060
rect 410 5960 440 5990
rect 610 6030 640 6060
rect 610 5960 640 5990
rect 810 6030 840 6060
rect 810 5960 840 5990
rect 1010 6030 1040 6060
rect 1010 5960 1040 5990
rect 1210 6030 1240 6060
rect 1210 5960 1240 5990
rect 1410 6030 1440 6060
rect 1410 5960 1440 5990
rect 1610 6030 1640 6060
rect 1610 5960 1640 5990
rect 1810 6030 1840 6060
rect 1810 5960 1840 5990
rect 2010 6030 2040 6060
rect 2010 5960 2040 5990
rect 2210 6030 2240 6060
rect 2210 5960 2240 5990
rect 2410 6030 2440 6060
rect 2410 5960 2440 5990
rect 2610 6030 2640 6060
rect 2610 5960 2640 5990
rect 2810 6030 2840 6060
rect 2810 5960 2840 5990
rect 3010 6030 3040 6060
rect 3010 5960 3040 5990
rect 3210 6030 3240 6060
rect 3210 5960 3240 5990
rect 3410 6030 3440 6060
rect 3410 5960 3440 5990
rect 3610 6030 3640 6060
rect 3610 5960 3640 5990
rect 3810 6030 3840 6060
rect 3810 5960 3840 5990
rect 4010 6030 4040 6060
rect 4010 5960 4040 5990
rect 4210 6030 4240 6060
rect 4210 5960 4240 5990
rect 4410 6030 4440 6060
rect 4410 5960 4440 5990
rect 4610 6030 4640 6060
rect 4610 5960 4640 5990
rect 4810 6030 4840 6060
rect 4810 5960 4840 5990
rect 5010 6030 5040 6060
rect 5010 5960 5040 5990
rect 5210 6030 5240 6060
rect 5210 5960 5240 5990
rect 5410 6030 5440 6060
rect 5410 5960 5440 5990
rect 5610 6030 5640 6060
rect 5610 5960 5640 5990
rect 5810 6030 5840 6060
rect 5810 5960 5840 5990
rect 6010 6030 6040 6060
rect 6010 5960 6040 5990
rect 6210 6030 6240 6060
rect 6210 5960 6240 5990
rect 6410 6030 6440 6060
rect 6410 5960 6440 5990
rect -190 5845 -160 5875
rect -190 5775 -160 5805
rect 10 5845 40 5875
rect 10 5775 40 5805
rect 210 5845 240 5875
rect 210 5775 240 5805
rect 410 5845 440 5875
rect 410 5775 440 5805
rect 610 5845 640 5875
rect 610 5775 640 5805
rect 810 5845 840 5875
rect 810 5775 840 5805
rect 1010 5845 1040 5875
rect 1010 5775 1040 5805
rect 1210 5845 1240 5875
rect 1210 5775 1240 5805
rect 1410 5845 1440 5875
rect 1410 5775 1440 5805
rect 1610 5845 1640 5875
rect 1610 5775 1640 5805
rect 1810 5845 1840 5875
rect 1810 5775 1840 5805
rect 2010 5845 2040 5875
rect 2010 5775 2040 5805
rect 2210 5845 2240 5875
rect 2210 5775 2240 5805
rect 2410 5845 2440 5875
rect 2410 5775 2440 5805
rect 2610 5845 2640 5875
rect 2610 5775 2640 5805
rect 2810 5845 2840 5875
rect 2810 5775 2840 5805
rect 3010 5845 3040 5875
rect 3010 5775 3040 5805
rect 3210 5845 3240 5875
rect 3210 5775 3240 5805
rect 3410 5845 3440 5875
rect 3410 5775 3440 5805
rect 3610 5845 3640 5875
rect 3610 5775 3640 5805
rect 3810 5845 3840 5875
rect 3810 5775 3840 5805
rect 4010 5845 4040 5875
rect 4010 5775 4040 5805
rect 4210 5845 4240 5875
rect 4210 5775 4240 5805
rect 4410 5845 4440 5875
rect 4410 5775 4440 5805
rect 4610 5845 4640 5875
rect 4610 5775 4640 5805
rect 4810 5845 4840 5875
rect 4810 5775 4840 5805
rect 5010 5845 5040 5875
rect 5010 5775 5040 5805
rect 5210 5845 5240 5875
rect 5210 5775 5240 5805
rect 5410 5845 5440 5875
rect 5410 5775 5440 5805
rect 5610 5845 5640 5875
rect 5610 5775 5640 5805
rect 5810 5845 5840 5875
rect 5810 5775 5840 5805
rect 6010 5845 6040 5875
rect 6010 5775 6040 5805
rect 6210 5845 6240 5875
rect 6210 5775 6240 5805
rect 6410 5845 6440 5875
rect 6410 5775 6440 5805
rect -190 5660 -160 5690
rect -190 5590 -160 5620
rect 10 5660 40 5690
rect 10 5590 40 5620
rect 210 5660 240 5690
rect 210 5590 240 5620
rect 410 5660 440 5690
rect 410 5590 440 5620
rect 610 5660 640 5690
rect 610 5590 640 5620
rect 810 5660 840 5690
rect 810 5590 840 5620
rect 1010 5660 1040 5690
rect 1010 5590 1040 5620
rect 1210 5660 1240 5690
rect 1210 5590 1240 5620
rect 1410 5660 1440 5690
rect 1410 5590 1440 5620
rect 1610 5660 1640 5690
rect 1610 5590 1640 5620
rect 1810 5660 1840 5690
rect 1810 5590 1840 5620
rect 2010 5660 2040 5690
rect 2010 5590 2040 5620
rect 2210 5660 2240 5690
rect 2210 5590 2240 5620
rect 2410 5660 2440 5690
rect 2410 5590 2440 5620
rect 2610 5660 2640 5690
rect 2610 5590 2640 5620
rect 2810 5660 2840 5690
rect 2810 5590 2840 5620
rect 3010 5660 3040 5690
rect 3010 5590 3040 5620
rect 3210 5660 3240 5690
rect 3210 5590 3240 5620
rect 3410 5660 3440 5690
rect 3410 5590 3440 5620
rect 3610 5660 3640 5690
rect 3610 5590 3640 5620
rect 3810 5660 3840 5690
rect 3810 5590 3840 5620
rect 4010 5660 4040 5690
rect 4010 5590 4040 5620
rect 4210 5660 4240 5690
rect 4210 5590 4240 5620
rect 4410 5660 4440 5690
rect 4410 5590 4440 5620
rect 4610 5660 4640 5690
rect 4610 5590 4640 5620
rect 4810 5660 4840 5690
rect 4810 5590 4840 5620
rect 5010 5660 5040 5690
rect 5010 5590 5040 5620
rect 5210 5660 5240 5690
rect 5210 5590 5240 5620
rect 5410 5660 5440 5690
rect 5410 5590 5440 5620
rect 5610 5660 5640 5690
rect 5610 5590 5640 5620
rect 5810 5660 5840 5690
rect 5810 5590 5840 5620
rect 6010 5660 6040 5690
rect 6010 5590 6040 5620
rect 6210 5660 6240 5690
rect 6210 5590 6240 5620
rect 6410 5660 6440 5690
rect 6410 5590 6440 5620
rect -190 5475 -160 5505
rect -190 5405 -160 5435
rect 10 5475 40 5505
rect 10 5405 40 5435
rect 210 5475 240 5505
rect 210 5405 240 5435
rect 410 5475 440 5505
rect 410 5405 440 5435
rect 610 5475 640 5505
rect 610 5405 640 5435
rect 810 5475 840 5505
rect 810 5405 840 5435
rect 1010 5475 1040 5505
rect 1010 5405 1040 5435
rect 1210 5475 1240 5505
rect 1210 5405 1240 5435
rect 1410 5475 1440 5505
rect 1410 5405 1440 5435
rect 1610 5475 1640 5505
rect 1610 5405 1640 5435
rect 1810 5475 1840 5505
rect 1810 5405 1840 5435
rect 2010 5475 2040 5505
rect 2010 5405 2040 5435
rect 2210 5475 2240 5505
rect 2210 5405 2240 5435
rect 2410 5475 2440 5505
rect 2410 5405 2440 5435
rect 2610 5475 2640 5505
rect 2610 5405 2640 5435
rect 2810 5475 2840 5505
rect 2810 5405 2840 5435
rect 3010 5475 3040 5505
rect 3010 5405 3040 5435
rect 3210 5475 3240 5505
rect 3210 5405 3240 5435
rect 3410 5475 3440 5505
rect 3410 5405 3440 5435
rect 3610 5475 3640 5505
rect 3610 5405 3640 5435
rect 3810 5475 3840 5505
rect 3810 5405 3840 5435
rect 4010 5475 4040 5505
rect 4010 5405 4040 5435
rect 4210 5475 4240 5505
rect 4210 5405 4240 5435
rect 4410 5475 4440 5505
rect 4410 5405 4440 5435
rect 4610 5475 4640 5505
rect 4610 5405 4640 5435
rect 4810 5475 4840 5505
rect 4810 5405 4840 5435
rect 5010 5475 5040 5505
rect 5010 5405 5040 5435
rect 5210 5475 5240 5505
rect 5210 5405 5240 5435
rect 5410 5475 5440 5505
rect 5410 5405 5440 5435
rect 5610 5475 5640 5505
rect 5610 5405 5640 5435
rect 5810 5475 5840 5505
rect 5810 5405 5840 5435
rect 6010 5475 6040 5505
rect 6010 5405 6040 5435
rect 6210 5475 6240 5505
rect 6210 5405 6240 5435
rect 6410 5475 6440 5505
rect 6410 5405 6440 5435
rect -190 5290 -160 5320
rect -190 5220 -160 5250
rect 10 5290 40 5320
rect 10 5220 40 5250
rect 210 5290 240 5320
rect 210 5220 240 5250
rect 410 5290 440 5320
rect 410 5220 440 5250
rect 610 5290 640 5320
rect 610 5220 640 5250
rect 810 5290 840 5320
rect 810 5220 840 5250
rect 1010 5290 1040 5320
rect 1010 5220 1040 5250
rect 1210 5290 1240 5320
rect 1210 5220 1240 5250
rect 1410 5290 1440 5320
rect 1410 5220 1440 5250
rect 1610 5290 1640 5320
rect 1610 5220 1640 5250
rect 1810 5290 1840 5320
rect 1810 5220 1840 5250
rect 2010 5290 2040 5320
rect 2010 5220 2040 5250
rect 2210 5290 2240 5320
rect 2210 5220 2240 5250
rect 2410 5290 2440 5320
rect 2410 5220 2440 5250
rect 2610 5290 2640 5320
rect 2610 5220 2640 5250
rect 2810 5290 2840 5320
rect 2810 5220 2840 5250
rect 3010 5290 3040 5320
rect 3010 5220 3040 5250
rect 3210 5290 3240 5320
rect 3210 5220 3240 5250
rect 3410 5290 3440 5320
rect 3410 5220 3440 5250
rect 3610 5290 3640 5320
rect 3610 5220 3640 5250
rect 3810 5290 3840 5320
rect 3810 5220 3840 5250
rect 4010 5290 4040 5320
rect 4010 5220 4040 5250
rect 4210 5290 4240 5320
rect 4210 5220 4240 5250
rect 4410 5290 4440 5320
rect 4410 5220 4440 5250
rect 4610 5290 4640 5320
rect 4610 5220 4640 5250
rect 4810 5290 4840 5320
rect 4810 5220 4840 5250
rect 5010 5290 5040 5320
rect 5010 5220 5040 5250
rect 5210 5290 5240 5320
rect 5210 5220 5240 5250
rect 5410 5290 5440 5320
rect 5410 5220 5440 5250
rect 5610 5290 5640 5320
rect 5610 5220 5640 5250
rect 5810 5290 5840 5320
rect 5810 5220 5840 5250
rect 6010 5290 6040 5320
rect 6010 5220 6040 5250
rect 6210 5290 6240 5320
rect 6210 5220 6240 5250
rect 6410 5290 6440 5320
rect 6410 5220 6440 5250
rect -190 5105 -160 5135
rect -190 5035 -160 5065
rect 10 5105 40 5135
rect 10 5035 40 5065
rect 210 5105 240 5135
rect 210 5035 240 5065
rect 410 5105 440 5135
rect 410 5035 440 5065
rect 610 5105 640 5135
rect 610 5035 640 5065
rect 810 5105 840 5135
rect 810 5035 840 5065
rect 1010 5105 1040 5135
rect 1010 5035 1040 5065
rect 1210 5105 1240 5135
rect 1210 5035 1240 5065
rect 1410 5105 1440 5135
rect 1410 5035 1440 5065
rect 1610 5105 1640 5135
rect 1610 5035 1640 5065
rect 1810 5105 1840 5135
rect 1810 5035 1840 5065
rect 2010 5105 2040 5135
rect 2010 5035 2040 5065
rect 2210 5105 2240 5135
rect 2210 5035 2240 5065
rect 2410 5105 2440 5135
rect 2410 5035 2440 5065
rect 2610 5105 2640 5135
rect 2610 5035 2640 5065
rect 2810 5105 2840 5135
rect 2810 5035 2840 5065
rect 3010 5105 3040 5135
rect 3010 5035 3040 5065
rect 3210 5105 3240 5135
rect 3210 5035 3240 5065
rect 3410 5105 3440 5135
rect 3410 5035 3440 5065
rect 3610 5105 3640 5135
rect 3610 5035 3640 5065
rect 3810 5105 3840 5135
rect 3810 5035 3840 5065
rect 4010 5105 4040 5135
rect 4010 5035 4040 5065
rect 4210 5105 4240 5135
rect 4210 5035 4240 5065
rect 4410 5105 4440 5135
rect 4410 5035 4440 5065
rect 4610 5105 4640 5135
rect 4610 5035 4640 5065
rect 4810 5105 4840 5135
rect 4810 5035 4840 5065
rect 5010 5105 5040 5135
rect 5010 5035 5040 5065
rect 5210 5105 5240 5135
rect 5210 5035 5240 5065
rect 5410 5105 5440 5135
rect 5410 5035 5440 5065
rect 5610 5105 5640 5135
rect 5610 5035 5640 5065
rect 5810 5105 5840 5135
rect 5810 5035 5840 5065
rect 6010 5105 6040 5135
rect 6010 5035 6040 5065
rect 6210 5105 6240 5135
rect 6210 5035 6240 5065
rect 6410 5105 6440 5135
rect 6410 5035 6440 5065
rect -190 4920 -160 4950
rect -190 4850 -160 4880
rect 10 4920 40 4950
rect 10 4850 40 4880
rect 210 4920 240 4950
rect 210 4850 240 4880
rect 410 4920 440 4950
rect 410 4850 440 4880
rect 610 4920 640 4950
rect 610 4850 640 4880
rect 810 4920 840 4950
rect 810 4850 840 4880
rect 1010 4920 1040 4950
rect 1010 4850 1040 4880
rect 1210 4920 1240 4950
rect 1210 4850 1240 4880
rect 1410 4920 1440 4950
rect 1410 4850 1440 4880
rect 1610 4920 1640 4950
rect 1610 4850 1640 4880
rect 1810 4920 1840 4950
rect 1810 4850 1840 4880
rect 2010 4920 2040 4950
rect 2010 4850 2040 4880
rect 2210 4920 2240 4950
rect 2210 4850 2240 4880
rect 2410 4920 2440 4950
rect 2410 4850 2440 4880
rect 2610 4920 2640 4950
rect 2610 4850 2640 4880
rect 2810 4920 2840 4950
rect 2810 4850 2840 4880
rect 3010 4920 3040 4950
rect 3010 4850 3040 4880
rect 3210 4920 3240 4950
rect 3210 4850 3240 4880
rect 3410 4920 3440 4950
rect 3410 4850 3440 4880
rect 3610 4920 3640 4950
rect 3610 4850 3640 4880
rect 3810 4920 3840 4950
rect 3810 4850 3840 4880
rect 4010 4920 4040 4950
rect 4010 4850 4040 4880
rect 4210 4920 4240 4950
rect 4210 4850 4240 4880
rect 4410 4920 4440 4950
rect 4410 4850 4440 4880
rect 4610 4920 4640 4950
rect 4610 4850 4640 4880
rect 4810 4920 4840 4950
rect 4810 4850 4840 4880
rect 5010 4920 5040 4950
rect 5010 4850 5040 4880
rect 5210 4920 5240 4950
rect 5210 4850 5240 4880
rect 5410 4920 5440 4950
rect 5410 4850 5440 4880
rect 5610 4920 5640 4950
rect 5610 4850 5640 4880
rect 5810 4920 5840 4950
rect 5810 4850 5840 4880
rect 6010 4920 6040 4950
rect 6010 4850 6040 4880
rect 6210 4920 6240 4950
rect 6210 4850 6240 4880
rect 6410 4920 6440 4950
rect 6410 4850 6440 4880
rect -190 4735 -160 4765
rect -190 4665 -160 4695
rect 10 4735 40 4765
rect 10 4665 40 4695
rect 210 4735 240 4765
rect 210 4665 240 4695
rect 410 4735 440 4765
rect 410 4665 440 4695
rect 610 4735 640 4765
rect 610 4665 640 4695
rect 810 4735 840 4765
rect 810 4665 840 4695
rect 1010 4735 1040 4765
rect 1010 4665 1040 4695
rect 1210 4735 1240 4765
rect 1210 4665 1240 4695
rect 1410 4735 1440 4765
rect 1410 4665 1440 4695
rect 1610 4735 1640 4765
rect 1610 4665 1640 4695
rect 1810 4735 1840 4765
rect 1810 4665 1840 4695
rect 2010 4735 2040 4765
rect 2010 4665 2040 4695
rect 2210 4735 2240 4765
rect 2210 4665 2240 4695
rect 2410 4735 2440 4765
rect 2410 4665 2440 4695
rect 2610 4735 2640 4765
rect 2610 4665 2640 4695
rect 2810 4735 2840 4765
rect 2810 4665 2840 4695
rect 3010 4735 3040 4765
rect 3010 4665 3040 4695
rect 3210 4735 3240 4765
rect 3210 4665 3240 4695
rect 3410 4735 3440 4765
rect 3410 4665 3440 4695
rect 3610 4735 3640 4765
rect 3610 4665 3640 4695
rect 3810 4735 3840 4765
rect 3810 4665 3840 4695
rect 4010 4735 4040 4765
rect 4010 4665 4040 4695
rect 4210 4735 4240 4765
rect 4210 4665 4240 4695
rect 4410 4735 4440 4765
rect 4410 4665 4440 4695
rect 4610 4735 4640 4765
rect 4610 4665 4640 4695
rect 4810 4735 4840 4765
rect 4810 4665 4840 4695
rect 5010 4735 5040 4765
rect 5010 4665 5040 4695
rect 5210 4735 5240 4765
rect 5210 4665 5240 4695
rect 5410 4735 5440 4765
rect 5410 4665 5440 4695
rect 5610 4735 5640 4765
rect 5610 4665 5640 4695
rect 5810 4735 5840 4765
rect 5810 4665 5840 4695
rect 6010 4735 6040 4765
rect 6010 4665 6040 4695
rect 6210 4735 6240 4765
rect 6210 4665 6240 4695
rect 6410 4735 6440 4765
rect 6410 4665 6440 4695
rect -190 4550 -160 4580
rect -190 4480 -160 4510
rect 10 4550 40 4580
rect 10 4480 40 4510
rect 210 4550 240 4580
rect 210 4480 240 4510
rect 410 4550 440 4580
rect 410 4480 440 4510
rect 610 4550 640 4580
rect 610 4480 640 4510
rect 810 4550 840 4580
rect 810 4480 840 4510
rect 1010 4550 1040 4580
rect 1010 4480 1040 4510
rect 1210 4550 1240 4580
rect 1210 4480 1240 4510
rect 1410 4550 1440 4580
rect 1410 4480 1440 4510
rect 1610 4550 1640 4580
rect 1610 4480 1640 4510
rect 1810 4550 1840 4580
rect 1810 4480 1840 4510
rect 2010 4550 2040 4580
rect 2010 4480 2040 4510
rect 2210 4550 2240 4580
rect 2210 4480 2240 4510
rect 2410 4550 2440 4580
rect 2410 4480 2440 4510
rect 2610 4550 2640 4580
rect 2610 4480 2640 4510
rect 2810 4550 2840 4580
rect 2810 4480 2840 4510
rect 3010 4550 3040 4580
rect 3010 4480 3040 4510
rect 3210 4550 3240 4580
rect 3210 4480 3240 4510
rect 3410 4550 3440 4580
rect 3410 4480 3440 4510
rect 3610 4550 3640 4580
rect 3610 4480 3640 4510
rect 3810 4550 3840 4580
rect 3810 4480 3840 4510
rect 4010 4550 4040 4580
rect 4010 4480 4040 4510
rect 4210 4550 4240 4580
rect 4210 4480 4240 4510
rect 4410 4550 4440 4580
rect 4410 4480 4440 4510
rect 4610 4550 4640 4580
rect 4610 4480 4640 4510
rect 4810 4550 4840 4580
rect 4810 4480 4840 4510
rect 5010 4550 5040 4580
rect 5010 4480 5040 4510
rect 5210 4550 5240 4580
rect 5210 4480 5240 4510
rect 5410 4550 5440 4580
rect 5410 4480 5440 4510
rect 5610 4550 5640 4580
rect 5610 4480 5640 4510
rect 5810 4550 5840 4580
rect 5810 4480 5840 4510
rect 6010 4550 6040 4580
rect 6010 4480 6040 4510
rect 6210 4550 6240 4580
rect 6210 4480 6240 4510
rect 6410 4550 6440 4580
rect 6410 4480 6440 4510
rect -190 4365 -160 4395
rect -190 4295 -160 4325
rect 10 4365 40 4395
rect 10 4295 40 4325
rect 210 4365 240 4395
rect 210 4295 240 4325
rect 410 4365 440 4395
rect 410 4295 440 4325
rect 610 4365 640 4395
rect 610 4295 640 4325
rect 810 4365 840 4395
rect 810 4295 840 4325
rect 1010 4365 1040 4395
rect 1010 4295 1040 4325
rect 1210 4365 1240 4395
rect 1210 4295 1240 4325
rect 1410 4365 1440 4395
rect 1410 4295 1440 4325
rect 1610 4365 1640 4395
rect 1610 4295 1640 4325
rect 1810 4365 1840 4395
rect 1810 4295 1840 4325
rect 2010 4365 2040 4395
rect 2010 4295 2040 4325
rect 2210 4365 2240 4395
rect 2210 4295 2240 4325
rect 2410 4365 2440 4395
rect 2410 4295 2440 4325
rect 2610 4365 2640 4395
rect 2610 4295 2640 4325
rect 2810 4365 2840 4395
rect 2810 4295 2840 4325
rect 3010 4365 3040 4395
rect 3010 4295 3040 4325
rect 3210 4365 3240 4395
rect 3210 4295 3240 4325
rect 3410 4365 3440 4395
rect 3410 4295 3440 4325
rect 3610 4365 3640 4395
rect 3610 4295 3640 4325
rect 3810 4365 3840 4395
rect 3810 4295 3840 4325
rect 4010 4365 4040 4395
rect 4010 4295 4040 4325
rect 4210 4365 4240 4395
rect 4210 4295 4240 4325
rect 4410 4365 4440 4395
rect 4410 4295 4440 4325
rect 4610 4365 4640 4395
rect 4610 4295 4640 4325
rect 4810 4365 4840 4395
rect 4810 4295 4840 4325
rect 5010 4365 5040 4395
rect 5010 4295 5040 4325
rect 5210 4365 5240 4395
rect 5210 4295 5240 4325
rect 5410 4365 5440 4395
rect 5410 4295 5440 4325
rect 5610 4365 5640 4395
rect 5610 4295 5640 4325
rect 5810 4365 5840 4395
rect 5810 4295 5840 4325
rect 6010 4365 6040 4395
rect 6010 4295 6040 4325
rect 6210 4365 6240 4395
rect 6210 4295 6240 4325
rect 6410 4365 6440 4395
rect 6410 4295 6440 4325
rect -190 4180 -160 4210
rect -190 4110 -160 4140
rect 10 4180 40 4210
rect 10 4110 40 4140
rect 210 4180 240 4210
rect 210 4110 240 4140
rect 410 4180 440 4210
rect 410 4110 440 4140
rect 610 4180 640 4210
rect 610 4110 640 4140
rect 810 4180 840 4210
rect 810 4110 840 4140
rect 1010 4180 1040 4210
rect 1010 4110 1040 4140
rect 1210 4180 1240 4210
rect 1210 4110 1240 4140
rect 1410 4180 1440 4210
rect 1410 4110 1440 4140
rect 1610 4180 1640 4210
rect 1610 4110 1640 4140
rect 1810 4180 1840 4210
rect 1810 4110 1840 4140
rect 2010 4180 2040 4210
rect 2010 4110 2040 4140
rect 2210 4180 2240 4210
rect 2210 4110 2240 4140
rect 2410 4180 2440 4210
rect 2410 4110 2440 4140
rect 2610 4180 2640 4210
rect 2610 4110 2640 4140
rect 2810 4180 2840 4210
rect 2810 4110 2840 4140
rect 3010 4180 3040 4210
rect 3010 4110 3040 4140
rect 3210 4180 3240 4210
rect 3210 4110 3240 4140
rect 3410 4180 3440 4210
rect 3410 4110 3440 4140
rect 3610 4180 3640 4210
rect 3610 4110 3640 4140
rect 3810 4180 3840 4210
rect 3810 4110 3840 4140
rect 4010 4180 4040 4210
rect 4010 4110 4040 4140
rect 4210 4180 4240 4210
rect 4210 4110 4240 4140
rect 4410 4180 4440 4210
rect 4410 4110 4440 4140
rect 4610 4180 4640 4210
rect 4610 4110 4640 4140
rect 4810 4180 4840 4210
rect 4810 4110 4840 4140
rect 5010 4180 5040 4210
rect 5010 4110 5040 4140
rect 5210 4180 5240 4210
rect 5210 4110 5240 4140
rect 5410 4180 5440 4210
rect 5410 4110 5440 4140
rect 5610 4180 5640 4210
rect 5610 4110 5640 4140
rect 5810 4180 5840 4210
rect 5810 4110 5840 4140
rect 6010 4180 6040 4210
rect 6010 4110 6040 4140
rect 6210 4180 6240 4210
rect 6210 4110 6240 4140
rect 6410 4180 6440 4210
rect 6410 4110 6440 4140
rect -190 3995 -160 4025
rect -190 3925 -160 3955
rect 10 3995 40 4025
rect 10 3925 40 3955
rect 210 3995 240 4025
rect 210 3925 240 3955
rect 410 3995 440 4025
rect 410 3925 440 3955
rect 610 3995 640 4025
rect 610 3925 640 3955
rect 810 3995 840 4025
rect 810 3925 840 3955
rect 1010 3995 1040 4025
rect 1010 3925 1040 3955
rect 1210 3995 1240 4025
rect 1210 3925 1240 3955
rect 1410 3995 1440 4025
rect 1410 3925 1440 3955
rect 1610 3995 1640 4025
rect 1610 3925 1640 3955
rect 1810 3995 1840 4025
rect 1810 3925 1840 3955
rect 2010 3995 2040 4025
rect 2010 3925 2040 3955
rect 2210 3995 2240 4025
rect 2210 3925 2240 3955
rect 2410 3995 2440 4025
rect 2410 3925 2440 3955
rect 2610 3995 2640 4025
rect 2610 3925 2640 3955
rect 2810 3995 2840 4025
rect 2810 3925 2840 3955
rect 3010 3995 3040 4025
rect 3010 3925 3040 3955
rect 3210 3995 3240 4025
rect 3210 3925 3240 3955
rect 3410 3995 3440 4025
rect 3410 3925 3440 3955
rect 3610 3995 3640 4025
rect 3610 3925 3640 3955
rect 3810 3995 3840 4025
rect 3810 3925 3840 3955
rect 4010 3995 4040 4025
rect 4010 3925 4040 3955
rect 4210 3995 4240 4025
rect 4210 3925 4240 3955
rect 4410 3995 4440 4025
rect 4410 3925 4440 3955
rect 4610 3995 4640 4025
rect 4610 3925 4640 3955
rect 4810 3995 4840 4025
rect 4810 3925 4840 3955
rect 5010 3995 5040 4025
rect 5010 3925 5040 3955
rect 5210 3995 5240 4025
rect 5210 3925 5240 3955
rect 5410 3995 5440 4025
rect 5410 3925 5440 3955
rect 5610 3995 5640 4025
rect 5610 3925 5640 3955
rect 5810 3995 5840 4025
rect 5810 3925 5840 3955
rect 6010 3995 6040 4025
rect 6010 3925 6040 3955
rect 6210 3995 6240 4025
rect 6210 3925 6240 3955
rect 6410 3995 6440 4025
rect 6410 3925 6440 3955
rect -190 3810 -160 3840
rect -190 3740 -160 3770
rect 10 3810 40 3840
rect 10 3740 40 3770
rect 210 3810 240 3840
rect 210 3740 240 3770
rect 410 3810 440 3840
rect 410 3740 440 3770
rect 610 3810 640 3840
rect 610 3740 640 3770
rect 810 3810 840 3840
rect 810 3740 840 3770
rect 1010 3810 1040 3840
rect 1010 3740 1040 3770
rect 1210 3810 1240 3840
rect 1210 3740 1240 3770
rect 1410 3810 1440 3840
rect 1410 3740 1440 3770
rect 1610 3810 1640 3840
rect 1610 3740 1640 3770
rect 1810 3810 1840 3840
rect 1810 3740 1840 3770
rect 2010 3810 2040 3840
rect 2010 3740 2040 3770
rect 2210 3810 2240 3840
rect 2210 3740 2240 3770
rect 2410 3810 2440 3840
rect 2410 3740 2440 3770
rect 2610 3810 2640 3840
rect 2610 3740 2640 3770
rect 2810 3810 2840 3840
rect 2810 3740 2840 3770
rect 3010 3810 3040 3840
rect 3010 3740 3040 3770
rect 3210 3810 3240 3840
rect 3210 3740 3240 3770
rect 3410 3810 3440 3840
rect 3410 3740 3440 3770
rect 3610 3810 3640 3840
rect 3610 3740 3640 3770
rect 3810 3810 3840 3840
rect 3810 3740 3840 3770
rect 4010 3810 4040 3840
rect 4010 3740 4040 3770
rect 4210 3810 4240 3840
rect 4210 3740 4240 3770
rect 4410 3810 4440 3840
rect 4410 3740 4440 3770
rect 4610 3810 4640 3840
rect 4610 3740 4640 3770
rect 4810 3810 4840 3840
rect 4810 3740 4840 3770
rect 5010 3810 5040 3840
rect 5010 3740 5040 3770
rect 5210 3810 5240 3840
rect 5210 3740 5240 3770
rect 5410 3810 5440 3840
rect 5410 3740 5440 3770
rect 5610 3810 5640 3840
rect 5610 3740 5640 3770
rect 5810 3810 5840 3840
rect 5810 3740 5840 3770
rect 6010 3810 6040 3840
rect 6010 3740 6040 3770
rect 6210 3810 6240 3840
rect 6210 3740 6240 3770
rect 6410 3810 6440 3840
rect 6410 3740 6440 3770
rect -190 3625 -160 3655
rect -190 3555 -160 3585
rect 10 3625 40 3655
rect 10 3555 40 3585
rect 210 3625 240 3655
rect 210 3555 240 3585
rect 410 3625 440 3655
rect 410 3555 440 3585
rect 610 3625 640 3655
rect 610 3555 640 3585
rect 810 3625 840 3655
rect 810 3555 840 3585
rect 1010 3625 1040 3655
rect 1010 3555 1040 3585
rect 1210 3625 1240 3655
rect 1210 3555 1240 3585
rect 1410 3625 1440 3655
rect 1410 3555 1440 3585
rect 1610 3625 1640 3655
rect 1610 3555 1640 3585
rect 1810 3625 1840 3655
rect 1810 3555 1840 3585
rect 2010 3625 2040 3655
rect 2010 3555 2040 3585
rect 2210 3625 2240 3655
rect 2210 3555 2240 3585
rect 2410 3625 2440 3655
rect 2410 3555 2440 3585
rect 2610 3625 2640 3655
rect 2610 3555 2640 3585
rect 2810 3625 2840 3655
rect 2810 3555 2840 3585
rect 3010 3625 3040 3655
rect 3010 3555 3040 3585
rect 3210 3625 3240 3655
rect 3210 3555 3240 3585
rect 3410 3625 3440 3655
rect 3410 3555 3440 3585
rect 3610 3625 3640 3655
rect 3610 3555 3640 3585
rect 3810 3625 3840 3655
rect 3810 3555 3840 3585
rect 4010 3625 4040 3655
rect 4010 3555 4040 3585
rect 4210 3625 4240 3655
rect 4210 3555 4240 3585
rect 4410 3625 4440 3655
rect 4410 3555 4440 3585
rect 4610 3625 4640 3655
rect 4610 3555 4640 3585
rect 4810 3625 4840 3655
rect 4810 3555 4840 3585
rect 5010 3625 5040 3655
rect 5010 3555 5040 3585
rect 5210 3625 5240 3655
rect 5210 3555 5240 3585
rect 5410 3625 5440 3655
rect 5410 3555 5440 3585
rect 5610 3625 5640 3655
rect 5610 3555 5640 3585
rect 5810 3625 5840 3655
rect 5810 3555 5840 3585
rect 6010 3625 6040 3655
rect 6010 3555 6040 3585
rect 6210 3625 6240 3655
rect 6210 3555 6240 3585
rect 6410 3625 6440 3655
rect 6410 3555 6440 3585
rect -190 3440 -160 3470
rect -190 3370 -160 3400
rect 10 3440 40 3470
rect 10 3370 40 3400
rect 210 3440 240 3470
rect 210 3370 240 3400
rect 410 3440 440 3470
rect 410 3370 440 3400
rect 610 3440 640 3470
rect 610 3370 640 3400
rect 810 3440 840 3470
rect 810 3370 840 3400
rect 1010 3440 1040 3470
rect 1010 3370 1040 3400
rect 1210 3440 1240 3470
rect 1210 3370 1240 3400
rect 1410 3440 1440 3470
rect 1410 3370 1440 3400
rect 1610 3440 1640 3470
rect 1610 3370 1640 3400
rect 1810 3440 1840 3470
rect 1810 3370 1840 3400
rect 2010 3440 2040 3470
rect 2010 3370 2040 3400
rect 2210 3440 2240 3470
rect 2210 3370 2240 3400
rect 2410 3440 2440 3470
rect 2410 3370 2440 3400
rect 2610 3440 2640 3470
rect 2610 3370 2640 3400
rect 2810 3440 2840 3470
rect 2810 3370 2840 3400
rect 3010 3440 3040 3470
rect 3010 3370 3040 3400
rect 3210 3440 3240 3470
rect 3210 3370 3240 3400
rect 3410 3440 3440 3470
rect 3410 3370 3440 3400
rect 3610 3440 3640 3470
rect 3610 3370 3640 3400
rect 3810 3440 3840 3470
rect 3810 3370 3840 3400
rect 4010 3440 4040 3470
rect 4010 3370 4040 3400
rect 4210 3440 4240 3470
rect 4210 3370 4240 3400
rect 4410 3440 4440 3470
rect 4410 3370 4440 3400
rect 4610 3440 4640 3470
rect 4610 3370 4640 3400
rect 4810 3440 4840 3470
rect 4810 3370 4840 3400
rect 5010 3440 5040 3470
rect 5010 3370 5040 3400
rect 5210 3440 5240 3470
rect 5210 3370 5240 3400
rect 5410 3440 5440 3470
rect 5410 3370 5440 3400
rect 5610 3440 5640 3470
rect 5610 3370 5640 3400
rect 5810 3440 5840 3470
rect 5810 3370 5840 3400
rect 6010 3440 6040 3470
rect 6010 3370 6040 3400
rect 6210 3440 6240 3470
rect 6210 3370 6240 3400
rect 6410 3440 6440 3470
rect 6410 3370 6440 3400
rect -190 3255 -160 3285
rect -190 3185 -160 3215
rect 10 3255 40 3285
rect 10 3185 40 3215
rect 210 3255 240 3285
rect 210 3185 240 3215
rect 410 3255 440 3285
rect 410 3185 440 3215
rect 610 3255 640 3285
rect 610 3185 640 3215
rect 810 3255 840 3285
rect 810 3185 840 3215
rect 1010 3255 1040 3285
rect 1010 3185 1040 3215
rect 1210 3255 1240 3285
rect 1210 3185 1240 3215
rect 1410 3255 1440 3285
rect 1410 3185 1440 3215
rect 1610 3255 1640 3285
rect 1610 3185 1640 3215
rect 1810 3255 1840 3285
rect 1810 3185 1840 3215
rect 2010 3255 2040 3285
rect 2010 3185 2040 3215
rect 2210 3255 2240 3285
rect 2210 3185 2240 3215
rect 2410 3255 2440 3285
rect 2410 3185 2440 3215
rect 2610 3255 2640 3285
rect 2610 3185 2640 3215
rect 2810 3255 2840 3285
rect 2810 3185 2840 3215
rect 3010 3255 3040 3285
rect 3010 3185 3040 3215
rect 3210 3255 3240 3285
rect 3210 3185 3240 3215
rect 3410 3255 3440 3285
rect 3410 3185 3440 3215
rect 3610 3255 3640 3285
rect 3610 3185 3640 3215
rect 3810 3255 3840 3285
rect 3810 3185 3840 3215
rect 4010 3255 4040 3285
rect 4010 3185 4040 3215
rect 4210 3255 4240 3285
rect 4210 3185 4240 3215
rect 4410 3255 4440 3285
rect 4410 3185 4440 3215
rect 4610 3255 4640 3285
rect 4610 3185 4640 3215
rect 4810 3255 4840 3285
rect 4810 3185 4840 3215
rect 5010 3255 5040 3285
rect 5010 3185 5040 3215
rect 5210 3255 5240 3285
rect 5210 3185 5240 3215
rect 5410 3255 5440 3285
rect 5410 3185 5440 3215
rect 5610 3255 5640 3285
rect 5610 3185 5640 3215
rect 5810 3255 5840 3285
rect 5810 3185 5840 3215
rect 6010 3255 6040 3285
rect 6010 3185 6040 3215
rect 6210 3255 6240 3285
rect 6210 3185 6240 3215
rect 6410 3255 6440 3285
rect 6410 3185 6440 3215
rect -190 3070 -160 3100
rect -190 3000 -160 3030
rect 10 3070 40 3100
rect 10 3000 40 3030
rect 210 3070 240 3100
rect 210 3000 240 3030
rect 410 3070 440 3100
rect 410 3000 440 3030
rect 610 3070 640 3100
rect 610 3000 640 3030
rect 810 3070 840 3100
rect 810 3000 840 3030
rect 1010 3070 1040 3100
rect 1010 3000 1040 3030
rect 1210 3070 1240 3100
rect 1210 3000 1240 3030
rect 1410 3070 1440 3100
rect 1410 3000 1440 3030
rect 1610 3070 1640 3100
rect 1610 3000 1640 3030
rect 1810 3070 1840 3100
rect 1810 3000 1840 3030
rect 2010 3070 2040 3100
rect 2010 3000 2040 3030
rect 2210 3070 2240 3100
rect 2210 3000 2240 3030
rect 2410 3070 2440 3100
rect 2410 3000 2440 3030
rect 2610 3070 2640 3100
rect 2610 3000 2640 3030
rect 2810 3070 2840 3100
rect 2810 3000 2840 3030
rect 3010 3070 3040 3100
rect 3010 3000 3040 3030
rect 3210 3070 3240 3100
rect 3210 3000 3240 3030
rect 3410 3070 3440 3100
rect 3410 3000 3440 3030
rect 3610 3070 3640 3100
rect 3610 3000 3640 3030
rect 3810 3070 3840 3100
rect 3810 3000 3840 3030
rect 4010 3070 4040 3100
rect 4010 3000 4040 3030
rect 4210 3070 4240 3100
rect 4210 3000 4240 3030
rect 4410 3070 4440 3100
rect 4410 3000 4440 3030
rect 4610 3070 4640 3100
rect 4610 3000 4640 3030
rect 4810 3070 4840 3100
rect 4810 3000 4840 3030
rect 5010 3070 5040 3100
rect 5010 3000 5040 3030
rect 5210 3070 5240 3100
rect 5210 3000 5240 3030
rect 5410 3070 5440 3100
rect 5410 3000 5440 3030
rect 5610 3070 5640 3100
rect 5610 3000 5640 3030
rect 5810 3070 5840 3100
rect 5810 3000 5840 3030
rect 6010 3070 6040 3100
rect 6010 3000 6040 3030
rect 6210 3070 6240 3100
rect 6210 3000 6240 3030
rect 6410 3070 6440 3100
rect 6410 3000 6440 3030
rect -190 2885 -160 2915
rect -190 2815 -160 2845
rect 10 2885 40 2915
rect 10 2815 40 2845
rect 210 2885 240 2915
rect 210 2815 240 2845
rect 410 2885 440 2915
rect 410 2815 440 2845
rect 610 2885 640 2915
rect 610 2815 640 2845
rect 810 2885 840 2915
rect 810 2815 840 2845
rect 1010 2885 1040 2915
rect 1010 2815 1040 2845
rect 1210 2885 1240 2915
rect 1210 2815 1240 2845
rect 1410 2885 1440 2915
rect 1410 2815 1440 2845
rect 1610 2885 1640 2915
rect 1610 2815 1640 2845
rect 1810 2885 1840 2915
rect 1810 2815 1840 2845
rect 2010 2885 2040 2915
rect 2010 2815 2040 2845
rect 2210 2885 2240 2915
rect 2210 2815 2240 2845
rect 2410 2885 2440 2915
rect 2410 2815 2440 2845
rect 2610 2885 2640 2915
rect 2610 2815 2640 2845
rect 2810 2885 2840 2915
rect 2810 2815 2840 2845
rect 3010 2885 3040 2915
rect 3010 2815 3040 2845
rect 3210 2885 3240 2915
rect 3210 2815 3240 2845
rect 3410 2885 3440 2915
rect 3410 2815 3440 2845
rect 3610 2885 3640 2915
rect 3610 2815 3640 2845
rect 3810 2885 3840 2915
rect 3810 2815 3840 2845
rect 4010 2885 4040 2915
rect 4010 2815 4040 2845
rect 4210 2885 4240 2915
rect 4210 2815 4240 2845
rect 4410 2885 4440 2915
rect 4410 2815 4440 2845
rect 4610 2885 4640 2915
rect 4610 2815 4640 2845
rect 4810 2885 4840 2915
rect 4810 2815 4840 2845
rect 5010 2885 5040 2915
rect 5010 2815 5040 2845
rect 5210 2885 5240 2915
rect 5210 2815 5240 2845
rect 5410 2885 5440 2915
rect 5410 2815 5440 2845
rect 5610 2885 5640 2915
rect 5610 2815 5640 2845
rect 5810 2885 5840 2915
rect 5810 2815 5840 2845
rect 6010 2885 6040 2915
rect 6010 2815 6040 2845
rect 6210 2885 6240 2915
rect 6210 2815 6240 2845
rect 6410 2885 6440 2915
rect 6410 2815 6440 2845
rect -190 2700 -160 2730
rect -190 2630 -160 2660
rect 10 2700 40 2730
rect 10 2630 40 2660
rect 210 2700 240 2730
rect 210 2630 240 2660
rect 410 2700 440 2730
rect 410 2630 440 2660
rect 610 2700 640 2730
rect 610 2630 640 2660
rect 810 2700 840 2730
rect 810 2630 840 2660
rect 1010 2700 1040 2730
rect 1010 2630 1040 2660
rect 1210 2700 1240 2730
rect 1210 2630 1240 2660
rect 1410 2700 1440 2730
rect 1410 2630 1440 2660
rect 1610 2700 1640 2730
rect 1610 2630 1640 2660
rect 1810 2700 1840 2730
rect 1810 2630 1840 2660
rect 2010 2700 2040 2730
rect 2010 2630 2040 2660
rect 2210 2700 2240 2730
rect 2210 2630 2240 2660
rect 2410 2700 2440 2730
rect 2410 2630 2440 2660
rect 2610 2700 2640 2730
rect 2610 2630 2640 2660
rect 2810 2700 2840 2730
rect 2810 2630 2840 2660
rect 3010 2700 3040 2730
rect 3010 2630 3040 2660
rect 3210 2700 3240 2730
rect 3210 2630 3240 2660
rect 3410 2700 3440 2730
rect 3410 2630 3440 2660
rect 3610 2700 3640 2730
rect 3610 2630 3640 2660
rect 3810 2700 3840 2730
rect 3810 2630 3840 2660
rect 4010 2700 4040 2730
rect 4010 2630 4040 2660
rect 4210 2700 4240 2730
rect 4210 2630 4240 2660
rect 4410 2700 4440 2730
rect 4410 2630 4440 2660
rect 4610 2700 4640 2730
rect 4610 2630 4640 2660
rect 4810 2700 4840 2730
rect 4810 2630 4840 2660
rect 5010 2700 5040 2730
rect 5010 2630 5040 2660
rect 5210 2700 5240 2730
rect 5210 2630 5240 2660
rect 5410 2700 5440 2730
rect 5410 2630 5440 2660
rect 5610 2700 5640 2730
rect 5610 2630 5640 2660
rect 5810 2700 5840 2730
rect 5810 2630 5840 2660
rect 6010 2700 6040 2730
rect 6010 2630 6040 2660
rect 6210 2700 6240 2730
rect 6210 2630 6240 2660
rect 6410 2700 6440 2730
rect 6410 2630 6440 2660
rect -190 2515 -160 2545
rect -190 2445 -160 2475
rect 10 2515 40 2545
rect 10 2445 40 2475
rect 210 2515 240 2545
rect 210 2445 240 2475
rect 410 2515 440 2545
rect 410 2445 440 2475
rect 610 2515 640 2545
rect 610 2445 640 2475
rect 810 2515 840 2545
rect 810 2445 840 2475
rect 1010 2515 1040 2545
rect 1010 2445 1040 2475
rect 1210 2515 1240 2545
rect 1210 2445 1240 2475
rect 1410 2515 1440 2545
rect 1410 2445 1440 2475
rect 1610 2515 1640 2545
rect 1610 2445 1640 2475
rect 1810 2515 1840 2545
rect 1810 2445 1840 2475
rect 2010 2515 2040 2545
rect 2010 2445 2040 2475
rect 2210 2515 2240 2545
rect 2210 2445 2240 2475
rect 2410 2515 2440 2545
rect 2410 2445 2440 2475
rect 2610 2515 2640 2545
rect 2610 2445 2640 2475
rect 2810 2515 2840 2545
rect 2810 2445 2840 2475
rect 3010 2515 3040 2545
rect 3010 2445 3040 2475
rect 3210 2515 3240 2545
rect 3210 2445 3240 2475
rect 3410 2515 3440 2545
rect 3410 2445 3440 2475
rect 3610 2515 3640 2545
rect 3610 2445 3640 2475
rect 3810 2515 3840 2545
rect 3810 2445 3840 2475
rect 4010 2515 4040 2545
rect 4010 2445 4040 2475
rect 4210 2515 4240 2545
rect 4210 2445 4240 2475
rect 4410 2515 4440 2545
rect 4410 2445 4440 2475
rect 4610 2515 4640 2545
rect 4610 2445 4640 2475
rect 4810 2515 4840 2545
rect 4810 2445 4840 2475
rect 5010 2515 5040 2545
rect 5010 2445 5040 2475
rect 5210 2515 5240 2545
rect 5210 2445 5240 2475
rect 5410 2515 5440 2545
rect 5410 2445 5440 2475
rect 5610 2515 5640 2545
rect 5610 2445 5640 2475
rect 5810 2515 5840 2545
rect 5810 2445 5840 2475
rect 6010 2515 6040 2545
rect 6010 2445 6040 2475
rect 6210 2515 6240 2545
rect 6210 2445 6240 2475
rect 6410 2515 6440 2545
rect 6410 2445 6440 2475
rect -190 2330 -160 2360
rect -190 2260 -160 2290
rect 10 2330 40 2360
rect 10 2260 40 2290
rect 210 2330 240 2360
rect 210 2260 240 2290
rect 410 2330 440 2360
rect 410 2260 440 2290
rect 610 2330 640 2360
rect 610 2260 640 2290
rect 810 2330 840 2360
rect 810 2260 840 2290
rect 1010 2330 1040 2360
rect 1010 2260 1040 2290
rect 1210 2330 1240 2360
rect 1210 2260 1240 2290
rect 1410 2330 1440 2360
rect 1410 2260 1440 2290
rect 1610 2330 1640 2360
rect 1610 2260 1640 2290
rect 1810 2330 1840 2360
rect 1810 2260 1840 2290
rect 2010 2330 2040 2360
rect 2010 2260 2040 2290
rect 2210 2330 2240 2360
rect 2210 2260 2240 2290
rect 2410 2330 2440 2360
rect 2410 2260 2440 2290
rect 2610 2330 2640 2360
rect 2610 2260 2640 2290
rect 2810 2330 2840 2360
rect 2810 2260 2840 2290
rect 3010 2330 3040 2360
rect 3010 2260 3040 2290
rect 3210 2330 3240 2360
rect 3210 2260 3240 2290
rect 3410 2330 3440 2360
rect 3410 2260 3440 2290
rect 3610 2330 3640 2360
rect 3610 2260 3640 2290
rect 3810 2330 3840 2360
rect 3810 2260 3840 2290
rect 4010 2330 4040 2360
rect 4010 2260 4040 2290
rect 4210 2330 4240 2360
rect 4210 2260 4240 2290
rect 4410 2330 4440 2360
rect 4410 2260 4440 2290
rect 4610 2330 4640 2360
rect 4610 2260 4640 2290
rect 4810 2330 4840 2360
rect 4810 2260 4840 2290
rect 5010 2330 5040 2360
rect 5010 2260 5040 2290
rect 5210 2330 5240 2360
rect 5210 2260 5240 2290
rect 5410 2330 5440 2360
rect 5410 2260 5440 2290
rect 5610 2330 5640 2360
rect 5610 2260 5640 2290
rect 5810 2330 5840 2360
rect 5810 2260 5840 2290
rect 6010 2330 6040 2360
rect 6010 2260 6040 2290
rect 6210 2330 6240 2360
rect 6210 2260 6240 2290
rect 6410 2330 6440 2360
rect 6410 2260 6440 2290
rect -190 2145 -160 2175
rect -190 2075 -160 2105
rect 10 2145 40 2175
rect 10 2075 40 2105
rect 210 2145 240 2175
rect 210 2075 240 2105
rect 410 2145 440 2175
rect 410 2075 440 2105
rect 610 2145 640 2175
rect 610 2075 640 2105
rect 810 2145 840 2175
rect 810 2075 840 2105
rect 1010 2145 1040 2175
rect 1010 2075 1040 2105
rect 1210 2145 1240 2175
rect 1210 2075 1240 2105
rect 1410 2145 1440 2175
rect 1410 2075 1440 2105
rect 1610 2145 1640 2175
rect 1610 2075 1640 2105
rect 1810 2145 1840 2175
rect 1810 2075 1840 2105
rect 2010 2145 2040 2175
rect 2010 2075 2040 2105
rect 2210 2145 2240 2175
rect 2210 2075 2240 2105
rect 2410 2145 2440 2175
rect 2410 2075 2440 2105
rect 2610 2145 2640 2175
rect 2610 2075 2640 2105
rect 2810 2145 2840 2175
rect 2810 2075 2840 2105
rect 3010 2145 3040 2175
rect 3010 2075 3040 2105
rect 3210 2145 3240 2175
rect 3210 2075 3240 2105
rect 3410 2145 3440 2175
rect 3410 2075 3440 2105
rect 3610 2145 3640 2175
rect 3610 2075 3640 2105
rect 3810 2145 3840 2175
rect 3810 2075 3840 2105
rect 4010 2145 4040 2175
rect 4010 2075 4040 2105
rect 4210 2145 4240 2175
rect 4210 2075 4240 2105
rect 4410 2145 4440 2175
rect 4410 2075 4440 2105
rect 4610 2145 4640 2175
rect 4610 2075 4640 2105
rect 4810 2145 4840 2175
rect 4810 2075 4840 2105
rect 5010 2145 5040 2175
rect 5010 2075 5040 2105
rect 5210 2145 5240 2175
rect 5210 2075 5240 2105
rect 5410 2145 5440 2175
rect 5410 2075 5440 2105
rect 5610 2145 5640 2175
rect 5610 2075 5640 2105
rect 5810 2145 5840 2175
rect 5810 2075 5840 2105
rect 6010 2145 6040 2175
rect 6010 2075 6040 2105
rect 6210 2145 6240 2175
rect 6210 2075 6240 2105
rect 6410 2145 6440 2175
rect 6410 2075 6440 2105
rect -190 1960 -160 1990
rect -190 1890 -160 1920
rect 10 1960 40 1990
rect 10 1890 40 1920
rect 210 1960 240 1990
rect 210 1890 240 1920
rect 410 1960 440 1990
rect 410 1890 440 1920
rect 610 1960 640 1990
rect 610 1890 640 1920
rect 810 1960 840 1990
rect 810 1890 840 1920
rect 1010 1960 1040 1990
rect 1010 1890 1040 1920
rect 1210 1960 1240 1990
rect 1210 1890 1240 1920
rect 1410 1960 1440 1990
rect 1410 1890 1440 1920
rect 1610 1960 1640 1990
rect 1610 1890 1640 1920
rect 1810 1960 1840 1990
rect 1810 1890 1840 1920
rect 2010 1960 2040 1990
rect 2010 1890 2040 1920
rect 2210 1960 2240 1990
rect 2210 1890 2240 1920
rect 2410 1960 2440 1990
rect 2410 1890 2440 1920
rect 2610 1960 2640 1990
rect 2610 1890 2640 1920
rect 2810 1960 2840 1990
rect 2810 1890 2840 1920
rect 3010 1960 3040 1990
rect 3010 1890 3040 1920
rect 3210 1960 3240 1990
rect 3210 1890 3240 1920
rect 3410 1960 3440 1990
rect 3410 1890 3440 1920
rect 3610 1960 3640 1990
rect 3610 1890 3640 1920
rect 3810 1960 3840 1990
rect 3810 1890 3840 1920
rect 4010 1960 4040 1990
rect 4010 1890 4040 1920
rect 4210 1960 4240 1990
rect 4210 1890 4240 1920
rect 4410 1960 4440 1990
rect 4410 1890 4440 1920
rect 4610 1960 4640 1990
rect 4610 1890 4640 1920
rect 4810 1960 4840 1990
rect 4810 1890 4840 1920
rect 5010 1960 5040 1990
rect 5010 1890 5040 1920
rect 5210 1960 5240 1990
rect 5210 1890 5240 1920
rect 5410 1960 5440 1990
rect 5410 1890 5440 1920
rect 5610 1960 5640 1990
rect 5610 1890 5640 1920
rect 5810 1960 5840 1990
rect 5810 1890 5840 1920
rect 6010 1960 6040 1990
rect 6010 1890 6040 1920
rect 6210 1960 6240 1990
rect 6210 1890 6240 1920
rect 6410 1960 6440 1990
rect 6410 1890 6440 1920
rect -190 1775 -160 1805
rect -190 1705 -160 1735
rect 10 1775 40 1805
rect 10 1705 40 1735
rect 210 1775 240 1805
rect 210 1705 240 1735
rect 410 1775 440 1805
rect 410 1705 440 1735
rect 610 1775 640 1805
rect 610 1705 640 1735
rect 810 1775 840 1805
rect 810 1705 840 1735
rect 1010 1775 1040 1805
rect 1010 1705 1040 1735
rect 1210 1775 1240 1805
rect 1210 1705 1240 1735
rect 1410 1775 1440 1805
rect 1410 1705 1440 1735
rect 1610 1775 1640 1805
rect 1610 1705 1640 1735
rect 1810 1775 1840 1805
rect 1810 1705 1840 1735
rect 2010 1775 2040 1805
rect 2010 1705 2040 1735
rect 2210 1775 2240 1805
rect 2210 1705 2240 1735
rect 2410 1775 2440 1805
rect 2410 1705 2440 1735
rect 2610 1775 2640 1805
rect 2610 1705 2640 1735
rect 2810 1775 2840 1805
rect 2810 1705 2840 1735
rect 3010 1775 3040 1805
rect 3010 1705 3040 1735
rect 3210 1775 3240 1805
rect 3210 1705 3240 1735
rect 3410 1775 3440 1805
rect 3410 1705 3440 1735
rect 3610 1775 3640 1805
rect 3610 1705 3640 1735
rect 3810 1775 3840 1805
rect 3810 1705 3840 1735
rect 4010 1775 4040 1805
rect 4010 1705 4040 1735
rect 4210 1775 4240 1805
rect 4210 1705 4240 1735
rect 4410 1775 4440 1805
rect 4410 1705 4440 1735
rect 4610 1775 4640 1805
rect 4610 1705 4640 1735
rect 4810 1775 4840 1805
rect 4810 1705 4840 1735
rect 5010 1775 5040 1805
rect 5010 1705 5040 1735
rect 5210 1775 5240 1805
rect 5210 1705 5240 1735
rect 5410 1775 5440 1805
rect 5410 1705 5440 1735
rect 5610 1775 5640 1805
rect 5610 1705 5640 1735
rect 5810 1775 5840 1805
rect 5810 1705 5840 1735
rect 6010 1775 6040 1805
rect 6010 1705 6040 1735
rect 6210 1775 6240 1805
rect 6210 1705 6240 1735
rect 6410 1775 6440 1805
rect 6410 1705 6440 1735
rect -190 1590 -160 1620
rect -190 1520 -160 1550
rect 10 1590 40 1620
rect 10 1520 40 1550
rect 210 1590 240 1620
rect 210 1520 240 1550
rect 410 1590 440 1620
rect 410 1520 440 1550
rect 610 1590 640 1620
rect 610 1520 640 1550
rect 810 1590 840 1620
rect 810 1520 840 1550
rect 1010 1590 1040 1620
rect 1010 1520 1040 1550
rect 1210 1590 1240 1620
rect 1210 1520 1240 1550
rect 1410 1590 1440 1620
rect 1410 1520 1440 1550
rect 1610 1590 1640 1620
rect 1610 1520 1640 1550
rect 1810 1590 1840 1620
rect 1810 1520 1840 1550
rect 2010 1590 2040 1620
rect 2010 1520 2040 1550
rect 2210 1590 2240 1620
rect 2210 1520 2240 1550
rect 2410 1590 2440 1620
rect 2410 1520 2440 1550
rect 2610 1590 2640 1620
rect 2610 1520 2640 1550
rect 2810 1590 2840 1620
rect 2810 1520 2840 1550
rect 3010 1590 3040 1620
rect 3010 1520 3040 1550
rect 3210 1590 3240 1620
rect 3210 1520 3240 1550
rect 3410 1590 3440 1620
rect 3410 1520 3440 1550
rect 3610 1590 3640 1620
rect 3610 1520 3640 1550
rect 3810 1590 3840 1620
rect 3810 1520 3840 1550
rect 4010 1590 4040 1620
rect 4010 1520 4040 1550
rect 4210 1590 4240 1620
rect 4210 1520 4240 1550
rect 4410 1590 4440 1620
rect 4410 1520 4440 1550
rect 4610 1590 4640 1620
rect 4610 1520 4640 1550
rect 4810 1590 4840 1620
rect 4810 1520 4840 1550
rect 5010 1590 5040 1620
rect 5010 1520 5040 1550
rect 5210 1590 5240 1620
rect 5210 1520 5240 1550
rect 5410 1590 5440 1620
rect 5410 1520 5440 1550
rect 5610 1590 5640 1620
rect 5610 1520 5640 1550
rect 5810 1590 5840 1620
rect 5810 1520 5840 1550
rect 6010 1590 6040 1620
rect 6010 1520 6040 1550
rect 6210 1590 6240 1620
rect 6210 1520 6240 1550
rect 6410 1590 6440 1620
rect 6410 1520 6440 1550
rect -190 1405 -160 1435
rect -190 1335 -160 1365
rect 10 1405 40 1435
rect 10 1335 40 1365
rect 210 1405 240 1435
rect 210 1335 240 1365
rect 410 1405 440 1435
rect 410 1335 440 1365
rect 610 1405 640 1435
rect 610 1335 640 1365
rect 810 1405 840 1435
rect 810 1335 840 1365
rect 1010 1405 1040 1435
rect 1010 1335 1040 1365
rect 1210 1405 1240 1435
rect 1210 1335 1240 1365
rect 1410 1405 1440 1435
rect 1410 1335 1440 1365
rect 1610 1405 1640 1435
rect 1610 1335 1640 1365
rect 1810 1405 1840 1435
rect 1810 1335 1840 1365
rect 2010 1405 2040 1435
rect 2010 1335 2040 1365
rect 2210 1405 2240 1435
rect 2210 1335 2240 1365
rect 2410 1405 2440 1435
rect 2410 1335 2440 1365
rect 2610 1405 2640 1435
rect 2610 1335 2640 1365
rect 2810 1405 2840 1435
rect 2810 1335 2840 1365
rect 3010 1405 3040 1435
rect 3010 1335 3040 1365
rect 3210 1405 3240 1435
rect 3210 1335 3240 1365
rect 3410 1405 3440 1435
rect 3410 1335 3440 1365
rect 3610 1405 3640 1435
rect 3610 1335 3640 1365
rect 3810 1405 3840 1435
rect 3810 1335 3840 1365
rect 4010 1405 4040 1435
rect 4010 1335 4040 1365
rect 4210 1405 4240 1435
rect 4210 1335 4240 1365
rect 4410 1405 4440 1435
rect 4410 1335 4440 1365
rect 4610 1405 4640 1435
rect 4610 1335 4640 1365
rect 4810 1405 4840 1435
rect 4810 1335 4840 1365
rect 5010 1405 5040 1435
rect 5010 1335 5040 1365
rect 5210 1405 5240 1435
rect 5210 1335 5240 1365
rect 5410 1405 5440 1435
rect 5410 1335 5440 1365
rect 5610 1405 5640 1435
rect 5610 1335 5640 1365
rect 5810 1405 5840 1435
rect 5810 1335 5840 1365
rect 6010 1405 6040 1435
rect 6010 1335 6040 1365
rect 6210 1405 6240 1435
rect 6210 1335 6240 1365
rect 6410 1405 6440 1435
rect 6410 1335 6440 1365
rect -190 1220 -160 1250
rect -190 1150 -160 1180
rect 10 1220 40 1250
rect 10 1150 40 1180
rect 210 1220 240 1250
rect 210 1150 240 1180
rect 410 1220 440 1250
rect 410 1150 440 1180
rect 610 1220 640 1250
rect 610 1150 640 1180
rect 810 1220 840 1250
rect 810 1150 840 1180
rect 1010 1220 1040 1250
rect 1010 1150 1040 1180
rect 1210 1220 1240 1250
rect 1210 1150 1240 1180
rect 1410 1220 1440 1250
rect 1410 1150 1440 1180
rect 1610 1220 1640 1250
rect 1610 1150 1640 1180
rect 1810 1220 1840 1250
rect 1810 1150 1840 1180
rect 2010 1220 2040 1250
rect 2010 1150 2040 1180
rect 2210 1220 2240 1250
rect 2210 1150 2240 1180
rect 2410 1220 2440 1250
rect 2410 1150 2440 1180
rect 2610 1220 2640 1250
rect 2610 1150 2640 1180
rect 2810 1220 2840 1250
rect 2810 1150 2840 1180
rect 3010 1220 3040 1250
rect 3010 1150 3040 1180
rect 3210 1220 3240 1250
rect 3210 1150 3240 1180
rect 3410 1220 3440 1250
rect 3410 1150 3440 1180
rect 3610 1220 3640 1250
rect 3610 1150 3640 1180
rect 3810 1220 3840 1250
rect 3810 1150 3840 1180
rect 4010 1220 4040 1250
rect 4010 1150 4040 1180
rect 4210 1220 4240 1250
rect 4210 1150 4240 1180
rect 4410 1220 4440 1250
rect 4410 1150 4440 1180
rect 4610 1220 4640 1250
rect 4610 1150 4640 1180
rect 4810 1220 4840 1250
rect 4810 1150 4840 1180
rect 5010 1220 5040 1250
rect 5010 1150 5040 1180
rect 5210 1220 5240 1250
rect 5210 1150 5240 1180
rect 5410 1220 5440 1250
rect 5410 1150 5440 1180
rect 5610 1220 5640 1250
rect 5610 1150 5640 1180
rect 5810 1220 5840 1250
rect 5810 1150 5840 1180
rect 6010 1220 6040 1250
rect 6010 1150 6040 1180
rect 6210 1220 6240 1250
rect 6210 1150 6240 1180
rect 6410 1220 6440 1250
rect 6410 1150 6440 1180
rect -190 1035 -160 1065
rect -190 965 -160 995
rect 10 1035 40 1065
rect 10 965 40 995
rect 210 1035 240 1065
rect 210 965 240 995
rect 410 1035 440 1065
rect 410 965 440 995
rect 610 1035 640 1065
rect 610 965 640 995
rect 810 1035 840 1065
rect 810 965 840 995
rect 1010 1035 1040 1065
rect 1010 965 1040 995
rect 1210 1035 1240 1065
rect 1210 965 1240 995
rect 1410 1035 1440 1065
rect 1410 965 1440 995
rect 1610 1035 1640 1065
rect 1610 965 1640 995
rect 1810 1035 1840 1065
rect 1810 965 1840 995
rect 2010 1035 2040 1065
rect 2010 965 2040 995
rect 2210 1035 2240 1065
rect 2210 965 2240 995
rect 2410 1035 2440 1065
rect 2410 965 2440 995
rect 2610 1035 2640 1065
rect 2610 965 2640 995
rect 2810 1035 2840 1065
rect 2810 965 2840 995
rect 3010 1035 3040 1065
rect 3010 965 3040 995
rect 3210 1035 3240 1065
rect 3210 965 3240 995
rect 3410 1035 3440 1065
rect 3410 965 3440 995
rect 3610 1035 3640 1065
rect 3610 965 3640 995
rect 3810 1035 3840 1065
rect 3810 965 3840 995
rect 4010 1035 4040 1065
rect 4010 965 4040 995
rect 4210 1035 4240 1065
rect 4210 965 4240 995
rect 4410 1035 4440 1065
rect 4410 965 4440 995
rect 4610 1035 4640 1065
rect 4610 965 4640 995
rect 4810 1035 4840 1065
rect 4810 965 4840 995
rect 5010 1035 5040 1065
rect 5010 965 5040 995
rect 5210 1035 5240 1065
rect 5210 965 5240 995
rect 5410 1035 5440 1065
rect 5410 965 5440 995
rect 5610 1035 5640 1065
rect 5610 965 5640 995
rect 5810 1035 5840 1065
rect 5810 965 5840 995
rect 6010 1035 6040 1065
rect 6010 965 6040 995
rect 6210 1035 6240 1065
rect 6210 965 6240 995
rect 6410 1035 6440 1065
rect 6410 965 6440 995
rect -190 850 -160 880
rect -190 780 -160 810
rect 10 850 40 880
rect 10 780 40 810
rect 210 850 240 880
rect 210 780 240 810
rect 410 850 440 880
rect 410 780 440 810
rect 610 850 640 880
rect 610 780 640 810
rect 810 850 840 880
rect 810 780 840 810
rect 1010 850 1040 880
rect 1010 780 1040 810
rect 1210 850 1240 880
rect 1210 780 1240 810
rect 1410 850 1440 880
rect 1410 780 1440 810
rect 1610 850 1640 880
rect 1610 780 1640 810
rect 1810 850 1840 880
rect 1810 780 1840 810
rect 2010 850 2040 880
rect 2010 780 2040 810
rect 2210 850 2240 880
rect 2210 780 2240 810
rect 2410 850 2440 880
rect 2410 780 2440 810
rect 2610 850 2640 880
rect 2610 780 2640 810
rect 2810 850 2840 880
rect 2810 780 2840 810
rect 3010 850 3040 880
rect 3010 780 3040 810
rect 3210 850 3240 880
rect 3210 780 3240 810
rect 3410 850 3440 880
rect 3410 780 3440 810
rect 3610 850 3640 880
rect 3610 780 3640 810
rect 3810 850 3840 880
rect 3810 780 3840 810
rect 4010 850 4040 880
rect 4010 780 4040 810
rect 4210 850 4240 880
rect 4210 780 4240 810
rect 4410 850 4440 880
rect 4410 780 4440 810
rect 4610 850 4640 880
rect 4610 780 4640 810
rect 4810 850 4840 880
rect 4810 780 4840 810
rect 5010 850 5040 880
rect 5010 780 5040 810
rect 5210 850 5240 880
rect 5210 780 5240 810
rect 5410 850 5440 880
rect 5410 780 5440 810
rect 5610 850 5640 880
rect 5610 780 5640 810
rect 5810 850 5840 880
rect 5810 780 5840 810
rect 6010 850 6040 880
rect 6010 780 6040 810
rect 6210 850 6240 880
rect 6210 780 6240 810
rect 6410 850 6440 880
rect 6410 780 6440 810
rect -190 665 -160 695
rect -190 595 -160 625
rect 10 665 40 695
rect 10 595 40 625
rect 210 665 240 695
rect 210 595 240 625
rect 410 665 440 695
rect 410 595 440 625
rect 610 665 640 695
rect 610 595 640 625
rect 810 665 840 695
rect 810 595 840 625
rect 1010 665 1040 695
rect 1010 595 1040 625
rect 1210 665 1240 695
rect 1210 595 1240 625
rect 1410 665 1440 695
rect 1410 595 1440 625
rect 1610 665 1640 695
rect 1610 595 1640 625
rect 1810 665 1840 695
rect 1810 595 1840 625
rect 2010 665 2040 695
rect 2010 595 2040 625
rect 2210 665 2240 695
rect 2210 595 2240 625
rect 2410 665 2440 695
rect 2410 595 2440 625
rect 2610 665 2640 695
rect 2610 595 2640 625
rect 2810 665 2840 695
rect 2810 595 2840 625
rect 3010 665 3040 695
rect 3010 595 3040 625
rect 3210 665 3240 695
rect 3210 595 3240 625
rect 3410 665 3440 695
rect 3410 595 3440 625
rect 3610 665 3640 695
rect 3610 595 3640 625
rect 3810 665 3840 695
rect 3810 595 3840 625
rect 4010 665 4040 695
rect 4010 595 4040 625
rect 4210 665 4240 695
rect 4210 595 4240 625
rect 4410 665 4440 695
rect 4410 595 4440 625
rect 4610 665 4640 695
rect 4610 595 4640 625
rect 4810 665 4840 695
rect 4810 595 4840 625
rect 5010 665 5040 695
rect 5010 595 5040 625
rect 5210 665 5240 695
rect 5210 595 5240 625
rect 5410 665 5440 695
rect 5410 595 5440 625
rect 5610 665 5640 695
rect 5610 595 5640 625
rect 5810 665 5840 695
rect 5810 595 5840 625
rect 6010 665 6040 695
rect 6010 595 6040 625
rect 6210 665 6240 695
rect 6210 595 6240 625
rect 6410 665 6440 695
rect 6410 595 6440 625
rect -190 480 -160 510
rect -190 410 -160 440
rect 10 480 40 510
rect 10 410 40 440
rect 210 480 240 510
rect 210 410 240 440
rect 410 480 440 510
rect 410 410 440 440
rect 610 480 640 510
rect 610 410 640 440
rect 810 480 840 510
rect 810 410 840 440
rect 1010 480 1040 510
rect 1010 410 1040 440
rect 1210 480 1240 510
rect 1210 410 1240 440
rect 1410 480 1440 510
rect 1410 410 1440 440
rect 1610 480 1640 510
rect 1610 410 1640 440
rect 1810 480 1840 510
rect 1810 410 1840 440
rect 2010 480 2040 510
rect 2010 410 2040 440
rect 2210 480 2240 510
rect 2210 410 2240 440
rect 2410 480 2440 510
rect 2410 410 2440 440
rect 2610 480 2640 510
rect 2610 410 2640 440
rect 2810 480 2840 510
rect 2810 410 2840 440
rect 3010 480 3040 510
rect 3010 410 3040 440
rect 3210 480 3240 510
rect 3210 410 3240 440
rect 3410 480 3440 510
rect 3410 410 3440 440
rect 3610 480 3640 510
rect 3610 410 3640 440
rect 3810 480 3840 510
rect 3810 410 3840 440
rect 4010 480 4040 510
rect 4010 410 4040 440
rect 4210 480 4240 510
rect 4210 410 4240 440
rect 4410 480 4440 510
rect 4410 410 4440 440
rect 4610 480 4640 510
rect 4610 410 4640 440
rect 4810 480 4840 510
rect 4810 410 4840 440
rect 5010 480 5040 510
rect 5010 410 5040 440
rect 5210 480 5240 510
rect 5210 410 5240 440
rect 5410 480 5440 510
rect 5410 410 5440 440
rect 5610 480 5640 510
rect 5610 410 5640 440
rect 5810 480 5840 510
rect 5810 410 5840 440
rect 6010 480 6040 510
rect 6010 410 6040 440
rect 6210 480 6240 510
rect 6210 410 6240 440
rect 6410 480 6440 510
rect 6410 410 6440 440
rect -190 295 -160 325
rect -190 225 -160 255
rect 10 295 40 325
rect 10 225 40 255
rect 210 295 240 325
rect 210 225 240 255
rect 410 295 440 325
rect 410 225 440 255
rect 610 295 640 325
rect 610 225 640 255
rect 810 295 840 325
rect 810 225 840 255
rect 1010 295 1040 325
rect 1010 225 1040 255
rect 1210 295 1240 325
rect 1210 225 1240 255
rect 1410 295 1440 325
rect 1410 225 1440 255
rect 1610 295 1640 325
rect 1610 225 1640 255
rect 1810 295 1840 325
rect 1810 225 1840 255
rect 2010 295 2040 325
rect 2010 225 2040 255
rect 2210 295 2240 325
rect 2210 225 2240 255
rect 2410 295 2440 325
rect 2410 225 2440 255
rect 2610 295 2640 325
rect 2610 225 2640 255
rect 2810 295 2840 325
rect 2810 225 2840 255
rect 3010 295 3040 325
rect 3010 225 3040 255
rect 3210 295 3240 325
rect 3210 225 3240 255
rect 3410 295 3440 325
rect 3410 225 3440 255
rect 3610 295 3640 325
rect 3610 225 3640 255
rect 3810 295 3840 325
rect 3810 225 3840 255
rect 4010 295 4040 325
rect 4010 225 4040 255
rect 4210 295 4240 325
rect 4210 225 4240 255
rect 4410 295 4440 325
rect 4410 225 4440 255
rect 4610 295 4640 325
rect 4610 225 4640 255
rect 4810 295 4840 325
rect 4810 225 4840 255
rect 5010 295 5040 325
rect 5010 225 5040 255
rect 5210 295 5240 325
rect 5210 225 5240 255
rect 5410 295 5440 325
rect 5410 225 5440 255
rect 5610 295 5640 325
rect 5610 225 5640 255
rect 5810 295 5840 325
rect 5810 225 5840 255
rect 6010 295 6040 325
rect 6010 225 6040 255
rect 6210 295 6240 325
rect 6210 225 6240 255
rect 6410 295 6440 325
rect 6410 225 6440 255
rect -190 110 -160 140
rect -190 40 -160 70
rect 10 110 40 140
rect 10 40 40 70
rect 210 110 240 140
rect 210 40 240 70
rect 410 110 440 140
rect 410 40 440 70
rect 610 110 640 140
rect 610 40 640 70
rect 810 110 840 140
rect 810 40 840 70
rect 1010 110 1040 140
rect 1010 40 1040 70
rect 1210 110 1240 140
rect 1210 40 1240 70
rect 1410 110 1440 140
rect 1410 40 1440 70
rect 1610 110 1640 140
rect 1610 40 1640 70
rect 1810 110 1840 140
rect 1810 40 1840 70
rect 2010 110 2040 140
rect 2010 40 2040 70
rect 2210 110 2240 140
rect 2210 40 2240 70
rect 2410 110 2440 140
rect 2410 40 2440 70
rect 2610 110 2640 140
rect 2610 40 2640 70
rect 2810 110 2840 140
rect 2810 40 2840 70
rect 3010 110 3040 140
rect 3010 40 3040 70
rect 3210 110 3240 140
rect 3210 40 3240 70
rect 3410 110 3440 140
rect 3410 40 3440 70
rect 3610 110 3640 140
rect 3610 40 3640 70
rect 3810 110 3840 140
rect 3810 40 3840 70
rect 4010 110 4040 140
rect 4010 40 4040 70
rect 4210 110 4240 140
rect 4210 40 4240 70
rect 4410 110 4440 140
rect 4410 40 4440 70
rect 4610 110 4640 140
rect 4610 40 4640 70
rect 4810 110 4840 140
rect 4810 40 4840 70
rect 5010 110 5040 140
rect 5010 40 5040 70
rect 5210 110 5240 140
rect 5210 40 5240 70
rect 5410 110 5440 140
rect 5410 40 5440 70
rect 5610 110 5640 140
rect 5610 40 5640 70
rect 5810 110 5840 140
rect 5810 40 5840 70
rect 6010 110 6040 140
rect 6010 40 6040 70
rect 6210 110 6240 140
rect 6210 40 6240 70
rect 6410 110 6440 140
rect 6410 40 6440 70
rect -190 -75 -160 -45
rect -190 -145 -160 -115
rect 10 -75 40 -45
rect 10 -145 40 -115
rect 210 -75 240 -45
rect 210 -145 240 -115
rect 410 -75 440 -45
rect 410 -145 440 -115
rect 610 -75 640 -45
rect 610 -145 640 -115
rect 810 -75 840 -45
rect 810 -145 840 -115
rect 1010 -75 1040 -45
rect 1010 -145 1040 -115
rect 1210 -75 1240 -45
rect 1210 -145 1240 -115
rect 1410 -75 1440 -45
rect 1410 -145 1440 -115
rect 1610 -75 1640 -45
rect 1610 -145 1640 -115
rect 1810 -75 1840 -45
rect 1810 -145 1840 -115
rect 2010 -75 2040 -45
rect 2010 -145 2040 -115
rect 2210 -75 2240 -45
rect 2210 -145 2240 -115
rect 2410 -75 2440 -45
rect 2410 -145 2440 -115
rect 2610 -75 2640 -45
rect 2610 -145 2640 -115
rect 2810 -75 2840 -45
rect 2810 -145 2840 -115
rect 3010 -75 3040 -45
rect 3010 -145 3040 -115
rect 3210 -75 3240 -45
rect 3210 -145 3240 -115
rect 3410 -75 3440 -45
rect 3410 -145 3440 -115
rect 3610 -75 3640 -45
rect 3610 -145 3640 -115
rect 3810 -75 3840 -45
rect 3810 -145 3840 -115
rect 4010 -75 4040 -45
rect 4010 -145 4040 -115
rect 4210 -75 4240 -45
rect 4210 -145 4240 -115
rect 4410 -75 4440 -45
rect 4410 -145 4440 -115
rect 4610 -75 4640 -45
rect 4610 -145 4640 -115
rect 4810 -75 4840 -45
rect 4810 -145 4840 -115
rect 5010 -75 5040 -45
rect 5010 -145 5040 -115
rect 5210 -75 5240 -45
rect 5210 -145 5240 -115
rect 5410 -75 5440 -45
rect 5410 -145 5440 -115
rect 5610 -75 5640 -45
rect 5610 -145 5640 -115
rect 5810 -75 5840 -45
rect 5810 -145 5840 -115
rect 6010 -75 6040 -45
rect 6010 -145 6040 -115
rect 6210 -75 6240 -45
rect 6210 -145 6240 -115
rect 6410 -75 6440 -45
rect 6410 -145 6440 -115
<< metal3 >>
rect -150 12055 -145 12095
rect -105 12055 -95 12095
rect -55 12055 -50 12095
rect 6450 12030 6455 12070
rect 6495 12030 6505 12070
rect 6545 12030 6550 12070
rect -200 11980 -30 12000
rect -200 11950 -190 11980
rect -160 11950 -30 11980
rect -200 11910 -30 11950
rect -200 11880 -190 11910
rect -160 11880 -30 11910
rect -200 11860 -30 11880
rect 0 11980 170 12000
rect 0 11950 10 11980
rect 40 11950 170 11980
rect 0 11910 170 11950
rect 0 11880 10 11910
rect 40 11880 170 11910
rect 0 11860 170 11880
rect 200 11980 370 12000
rect 200 11950 210 11980
rect 240 11950 370 11980
rect 200 11910 370 11950
rect 200 11880 210 11910
rect 240 11880 370 11910
rect 200 11860 370 11880
rect 400 11980 570 12000
rect 400 11950 410 11980
rect 440 11950 570 11980
rect 400 11910 570 11950
rect 400 11880 410 11910
rect 440 11880 570 11910
rect 400 11860 570 11880
rect 600 11980 770 12000
rect 600 11950 610 11980
rect 640 11950 770 11980
rect 600 11910 770 11950
rect 600 11880 610 11910
rect 640 11880 770 11910
rect 600 11860 770 11880
rect 800 11980 970 12000
rect 800 11950 810 11980
rect 840 11950 970 11980
rect 800 11910 970 11950
rect 800 11880 810 11910
rect 840 11880 970 11910
rect 800 11860 970 11880
rect 1000 11980 1170 12000
rect 1000 11950 1010 11980
rect 1040 11950 1170 11980
rect 1000 11910 1170 11950
rect 1000 11880 1010 11910
rect 1040 11880 1170 11910
rect 1000 11860 1170 11880
rect 1200 11980 1370 12000
rect 1200 11950 1210 11980
rect 1240 11950 1370 11980
rect 1200 11910 1370 11950
rect 1200 11880 1210 11910
rect 1240 11880 1370 11910
rect 1200 11860 1370 11880
rect 1400 11980 1570 12000
rect 1400 11950 1410 11980
rect 1440 11950 1570 11980
rect 1400 11910 1570 11950
rect 1400 11880 1410 11910
rect 1440 11880 1570 11910
rect 1400 11860 1570 11880
rect 1600 11980 1770 12000
rect 1600 11950 1610 11980
rect 1640 11950 1770 11980
rect 1600 11910 1770 11950
rect 1600 11880 1610 11910
rect 1640 11880 1770 11910
rect 1600 11860 1770 11880
rect 1800 11980 1970 12000
rect 1800 11950 1810 11980
rect 1840 11950 1970 11980
rect 1800 11910 1970 11950
rect 1800 11880 1810 11910
rect 1840 11880 1970 11910
rect 1800 11860 1970 11880
rect 2000 11980 2170 12000
rect 2000 11950 2010 11980
rect 2040 11950 2170 11980
rect 2000 11910 2170 11950
rect 2000 11880 2010 11910
rect 2040 11880 2170 11910
rect 2000 11860 2170 11880
rect 2200 11980 2370 12000
rect 2200 11950 2210 11980
rect 2240 11950 2370 11980
rect 2200 11910 2370 11950
rect 2200 11880 2210 11910
rect 2240 11880 2370 11910
rect 2200 11860 2370 11880
rect 2400 11980 2570 12000
rect 2400 11950 2410 11980
rect 2440 11950 2570 11980
rect 2400 11910 2570 11950
rect 2400 11880 2410 11910
rect 2440 11880 2570 11910
rect 2400 11860 2570 11880
rect 2600 11980 2770 12000
rect 2600 11950 2610 11980
rect 2640 11950 2770 11980
rect 2600 11910 2770 11950
rect 2600 11880 2610 11910
rect 2640 11880 2770 11910
rect 2600 11860 2770 11880
rect 2800 11980 2970 12000
rect 2800 11950 2810 11980
rect 2840 11950 2970 11980
rect 2800 11910 2970 11950
rect 2800 11880 2810 11910
rect 2840 11880 2970 11910
rect 2800 11860 2970 11880
rect 3000 11980 3170 12000
rect 3000 11950 3010 11980
rect 3040 11950 3170 11980
rect 3000 11910 3170 11950
rect 3000 11880 3010 11910
rect 3040 11880 3170 11910
rect 3000 11860 3170 11880
rect 3200 11980 3370 12000
rect 3200 11950 3210 11980
rect 3240 11950 3370 11980
rect 3200 11910 3370 11950
rect 3200 11880 3210 11910
rect 3240 11880 3370 11910
rect 3200 11860 3370 11880
rect 3400 11980 3570 12000
rect 3400 11950 3410 11980
rect 3440 11950 3570 11980
rect 3400 11910 3570 11950
rect 3400 11880 3410 11910
rect 3440 11880 3570 11910
rect 3400 11860 3570 11880
rect 3600 11980 3770 12000
rect 3600 11950 3610 11980
rect 3640 11950 3770 11980
rect 3600 11910 3770 11950
rect 3600 11880 3610 11910
rect 3640 11880 3770 11910
rect 3600 11860 3770 11880
rect 3800 11980 3970 12000
rect 3800 11950 3810 11980
rect 3840 11950 3970 11980
rect 3800 11910 3970 11950
rect 3800 11880 3810 11910
rect 3840 11880 3970 11910
rect 3800 11860 3970 11880
rect 4000 11980 4170 12000
rect 4000 11950 4010 11980
rect 4040 11950 4170 11980
rect 4000 11910 4170 11950
rect 4000 11880 4010 11910
rect 4040 11880 4170 11910
rect 4000 11860 4170 11880
rect 4200 11980 4370 12000
rect 4200 11950 4210 11980
rect 4240 11950 4370 11980
rect 4200 11910 4370 11950
rect 4200 11880 4210 11910
rect 4240 11880 4370 11910
rect 4200 11860 4370 11880
rect 4400 11980 4570 12000
rect 4400 11950 4410 11980
rect 4440 11950 4570 11980
rect 4400 11910 4570 11950
rect 4400 11880 4410 11910
rect 4440 11880 4570 11910
rect 4400 11860 4570 11880
rect 4600 11980 4770 12000
rect 4600 11950 4610 11980
rect 4640 11950 4770 11980
rect 4600 11910 4770 11950
rect 4600 11880 4610 11910
rect 4640 11880 4770 11910
rect 4600 11860 4770 11880
rect 4800 11980 4970 12000
rect 4800 11950 4810 11980
rect 4840 11950 4970 11980
rect 4800 11910 4970 11950
rect 4800 11880 4810 11910
rect 4840 11880 4970 11910
rect 4800 11860 4970 11880
rect 5000 11980 5170 12000
rect 5000 11950 5010 11980
rect 5040 11950 5170 11980
rect 5000 11910 5170 11950
rect 5000 11880 5010 11910
rect 5040 11880 5170 11910
rect 5000 11860 5170 11880
rect 5200 11980 5370 12000
rect 5200 11950 5210 11980
rect 5240 11950 5370 11980
rect 5200 11910 5370 11950
rect 5200 11880 5210 11910
rect 5240 11880 5370 11910
rect 5200 11860 5370 11880
rect 5400 11980 5570 12000
rect 5400 11950 5410 11980
rect 5440 11950 5570 11980
rect 5400 11910 5570 11950
rect 5400 11880 5410 11910
rect 5440 11880 5570 11910
rect 5400 11860 5570 11880
rect 5600 11980 5770 12000
rect 5600 11950 5610 11980
rect 5640 11950 5770 11980
rect 5600 11910 5770 11950
rect 5600 11880 5610 11910
rect 5640 11880 5770 11910
rect 5600 11860 5770 11880
rect 5800 11980 5970 12000
rect 5800 11950 5810 11980
rect 5840 11950 5970 11980
rect 5800 11910 5970 11950
rect 5800 11880 5810 11910
rect 5840 11880 5970 11910
rect 5800 11860 5970 11880
rect 6000 11980 6170 12000
rect 6000 11950 6010 11980
rect 6040 11950 6170 11980
rect 6000 11910 6170 11950
rect 6000 11880 6010 11910
rect 6040 11880 6170 11910
rect 6000 11860 6170 11880
rect 6200 11980 6370 12000
rect 6200 11950 6210 11980
rect 6240 11950 6370 11980
rect 6200 11910 6370 11950
rect 6200 11880 6210 11910
rect 6240 11880 6370 11910
rect 6200 11860 6370 11880
rect 6400 11980 6570 12000
rect 6400 11950 6410 11980
rect 6440 11950 6570 11980
rect 6400 11910 6570 11950
rect 6400 11880 6410 11910
rect 6440 11880 6570 11910
rect 6400 11860 6570 11880
rect -200 11795 -30 11815
rect -200 11765 -190 11795
rect -160 11765 -30 11795
rect -200 11725 -30 11765
rect -200 11695 -190 11725
rect -160 11695 -30 11725
rect -200 11675 -30 11695
rect 0 11795 170 11815
rect 0 11765 10 11795
rect 40 11765 170 11795
rect 0 11725 170 11765
rect 0 11695 10 11725
rect 40 11695 170 11725
rect 0 11675 170 11695
rect 200 11795 370 11815
rect 200 11765 210 11795
rect 240 11765 370 11795
rect 200 11725 370 11765
rect 200 11695 210 11725
rect 240 11695 370 11725
rect 200 11675 370 11695
rect 400 11795 570 11815
rect 400 11765 410 11795
rect 440 11765 570 11795
rect 400 11725 570 11765
rect 400 11695 410 11725
rect 440 11695 570 11725
rect 400 11675 570 11695
rect 600 11795 770 11815
rect 600 11765 610 11795
rect 640 11765 770 11795
rect 600 11725 770 11765
rect 600 11695 610 11725
rect 640 11695 770 11725
rect 600 11675 770 11695
rect 800 11795 970 11815
rect 800 11765 810 11795
rect 840 11765 970 11795
rect 800 11725 970 11765
rect 800 11695 810 11725
rect 840 11695 970 11725
rect 800 11675 970 11695
rect 1000 11795 1170 11815
rect 1000 11765 1010 11795
rect 1040 11765 1170 11795
rect 1000 11725 1170 11765
rect 1000 11695 1010 11725
rect 1040 11695 1170 11725
rect 1000 11675 1170 11695
rect 1200 11795 1370 11815
rect 1200 11765 1210 11795
rect 1240 11765 1370 11795
rect 1200 11725 1370 11765
rect 1200 11695 1210 11725
rect 1240 11695 1370 11725
rect 1200 11675 1370 11695
rect 1400 11795 1570 11815
rect 1400 11765 1410 11795
rect 1440 11765 1570 11795
rect 1400 11725 1570 11765
rect 1400 11695 1410 11725
rect 1440 11695 1570 11725
rect 1400 11675 1570 11695
rect 1600 11795 1770 11815
rect 1600 11765 1610 11795
rect 1640 11765 1770 11795
rect 1600 11725 1770 11765
rect 1600 11695 1610 11725
rect 1640 11695 1770 11725
rect 1600 11675 1770 11695
rect 1800 11795 1970 11815
rect 1800 11765 1810 11795
rect 1840 11765 1970 11795
rect 1800 11725 1970 11765
rect 1800 11695 1810 11725
rect 1840 11695 1970 11725
rect 1800 11675 1970 11695
rect 2000 11795 2170 11815
rect 2000 11765 2010 11795
rect 2040 11765 2170 11795
rect 2000 11725 2170 11765
rect 2000 11695 2010 11725
rect 2040 11695 2170 11725
rect 2000 11675 2170 11695
rect 2200 11795 2370 11815
rect 2200 11765 2210 11795
rect 2240 11765 2370 11795
rect 2200 11725 2370 11765
rect 2200 11695 2210 11725
rect 2240 11695 2370 11725
rect 2200 11675 2370 11695
rect 2400 11795 2570 11815
rect 2400 11765 2410 11795
rect 2440 11765 2570 11795
rect 2400 11725 2570 11765
rect 2400 11695 2410 11725
rect 2440 11695 2570 11725
rect 2400 11675 2570 11695
rect 2600 11795 2770 11815
rect 2600 11765 2610 11795
rect 2640 11765 2770 11795
rect 2600 11725 2770 11765
rect 2600 11695 2610 11725
rect 2640 11695 2770 11725
rect 2600 11675 2770 11695
rect 2800 11795 2970 11815
rect 2800 11765 2810 11795
rect 2840 11765 2970 11795
rect 2800 11725 2970 11765
rect 2800 11695 2810 11725
rect 2840 11695 2970 11725
rect 2800 11675 2970 11695
rect 3000 11795 3170 11815
rect 3000 11765 3010 11795
rect 3040 11765 3170 11795
rect 3000 11725 3170 11765
rect 3000 11695 3010 11725
rect 3040 11695 3170 11725
rect 3000 11675 3170 11695
rect 3200 11795 3370 11815
rect 3200 11765 3210 11795
rect 3240 11765 3370 11795
rect 3200 11725 3370 11765
rect 3200 11695 3210 11725
rect 3240 11695 3370 11725
rect 3200 11675 3370 11695
rect 3400 11795 3570 11815
rect 3400 11765 3410 11795
rect 3440 11765 3570 11795
rect 3400 11725 3570 11765
rect 3400 11695 3410 11725
rect 3440 11695 3570 11725
rect 3400 11675 3570 11695
rect 3600 11795 3770 11815
rect 3600 11765 3610 11795
rect 3640 11765 3770 11795
rect 3600 11725 3770 11765
rect 3600 11695 3610 11725
rect 3640 11695 3770 11725
rect 3600 11675 3770 11695
rect 3800 11795 3970 11815
rect 3800 11765 3810 11795
rect 3840 11765 3970 11795
rect 3800 11725 3970 11765
rect 3800 11695 3810 11725
rect 3840 11695 3970 11725
rect 3800 11675 3970 11695
rect 4000 11795 4170 11815
rect 4000 11765 4010 11795
rect 4040 11765 4170 11795
rect 4000 11725 4170 11765
rect 4000 11695 4010 11725
rect 4040 11695 4170 11725
rect 4000 11675 4170 11695
rect 4200 11795 4370 11815
rect 4200 11765 4210 11795
rect 4240 11765 4370 11795
rect 4200 11725 4370 11765
rect 4200 11695 4210 11725
rect 4240 11695 4370 11725
rect 4200 11675 4370 11695
rect 4400 11795 4570 11815
rect 4400 11765 4410 11795
rect 4440 11765 4570 11795
rect 4400 11725 4570 11765
rect 4400 11695 4410 11725
rect 4440 11695 4570 11725
rect 4400 11675 4570 11695
rect 4600 11795 4770 11815
rect 4600 11765 4610 11795
rect 4640 11765 4770 11795
rect 4600 11725 4770 11765
rect 4600 11695 4610 11725
rect 4640 11695 4770 11725
rect 4600 11675 4770 11695
rect 4800 11795 4970 11815
rect 4800 11765 4810 11795
rect 4840 11765 4970 11795
rect 4800 11725 4970 11765
rect 4800 11695 4810 11725
rect 4840 11695 4970 11725
rect 4800 11675 4970 11695
rect 5000 11795 5170 11815
rect 5000 11765 5010 11795
rect 5040 11765 5170 11795
rect 5000 11725 5170 11765
rect 5000 11695 5010 11725
rect 5040 11695 5170 11725
rect 5000 11675 5170 11695
rect 5200 11795 5370 11815
rect 5200 11765 5210 11795
rect 5240 11765 5370 11795
rect 5200 11725 5370 11765
rect 5200 11695 5210 11725
rect 5240 11695 5370 11725
rect 5200 11675 5370 11695
rect 5400 11795 5570 11815
rect 5400 11765 5410 11795
rect 5440 11765 5570 11795
rect 5400 11725 5570 11765
rect 5400 11695 5410 11725
rect 5440 11695 5570 11725
rect 5400 11675 5570 11695
rect 5600 11795 5770 11815
rect 5600 11765 5610 11795
rect 5640 11765 5770 11795
rect 5600 11725 5770 11765
rect 5600 11695 5610 11725
rect 5640 11695 5770 11725
rect 5600 11675 5770 11695
rect 5800 11795 5970 11815
rect 5800 11765 5810 11795
rect 5840 11765 5970 11795
rect 5800 11725 5970 11765
rect 5800 11695 5810 11725
rect 5840 11695 5970 11725
rect 5800 11675 5970 11695
rect 6000 11795 6170 11815
rect 6000 11765 6010 11795
rect 6040 11765 6170 11795
rect 6000 11725 6170 11765
rect 6000 11695 6010 11725
rect 6040 11695 6170 11725
rect 6000 11675 6170 11695
rect 6200 11795 6370 11815
rect 6200 11765 6210 11795
rect 6240 11765 6370 11795
rect 6200 11725 6370 11765
rect 6200 11695 6210 11725
rect 6240 11695 6370 11725
rect 6200 11675 6370 11695
rect 6400 11795 6570 11815
rect 6400 11765 6410 11795
rect 6440 11765 6570 11795
rect 6400 11725 6570 11765
rect 6400 11695 6410 11725
rect 6440 11695 6570 11725
rect 6400 11675 6570 11695
rect -200 11610 -30 11630
rect -200 11580 -190 11610
rect -160 11580 -30 11610
rect -200 11540 -30 11580
rect -200 11510 -190 11540
rect -160 11510 -30 11540
rect -200 11490 -30 11510
rect 0 11610 170 11630
rect 0 11580 10 11610
rect 40 11580 170 11610
rect 0 11540 170 11580
rect 0 11510 10 11540
rect 40 11510 170 11540
rect 0 11490 170 11510
rect 200 11610 370 11630
rect 200 11580 210 11610
rect 240 11580 370 11610
rect 200 11540 370 11580
rect 200 11510 210 11540
rect 240 11510 370 11540
rect 200 11490 370 11510
rect 400 11610 570 11630
rect 400 11580 410 11610
rect 440 11580 570 11610
rect 400 11540 570 11580
rect 400 11510 410 11540
rect 440 11510 570 11540
rect 400 11490 570 11510
rect 600 11610 770 11630
rect 600 11580 610 11610
rect 640 11580 770 11610
rect 600 11540 770 11580
rect 600 11510 610 11540
rect 640 11510 770 11540
rect 600 11490 770 11510
rect 800 11610 970 11630
rect 800 11580 810 11610
rect 840 11580 970 11610
rect 800 11540 970 11580
rect 800 11510 810 11540
rect 840 11510 970 11540
rect 800 11490 970 11510
rect 1000 11610 1170 11630
rect 1000 11580 1010 11610
rect 1040 11580 1170 11610
rect 1000 11540 1170 11580
rect 1000 11510 1010 11540
rect 1040 11510 1170 11540
rect 1000 11490 1170 11510
rect 1200 11610 1370 11630
rect 1200 11580 1210 11610
rect 1240 11580 1370 11610
rect 1200 11540 1370 11580
rect 1200 11510 1210 11540
rect 1240 11510 1370 11540
rect 1200 11490 1370 11510
rect 1400 11610 1570 11630
rect 1400 11580 1410 11610
rect 1440 11580 1570 11610
rect 1400 11540 1570 11580
rect 1400 11510 1410 11540
rect 1440 11510 1570 11540
rect 1400 11490 1570 11510
rect 1600 11610 1770 11630
rect 1600 11580 1610 11610
rect 1640 11580 1770 11610
rect 1600 11540 1770 11580
rect 1600 11510 1610 11540
rect 1640 11510 1770 11540
rect 1600 11490 1770 11510
rect 1800 11610 1970 11630
rect 1800 11580 1810 11610
rect 1840 11580 1970 11610
rect 1800 11540 1970 11580
rect 1800 11510 1810 11540
rect 1840 11510 1970 11540
rect 1800 11490 1970 11510
rect 2000 11610 2170 11630
rect 2000 11580 2010 11610
rect 2040 11580 2170 11610
rect 2000 11540 2170 11580
rect 2000 11510 2010 11540
rect 2040 11510 2170 11540
rect 2000 11490 2170 11510
rect 2200 11610 2370 11630
rect 2200 11580 2210 11610
rect 2240 11580 2370 11610
rect 2200 11540 2370 11580
rect 2200 11510 2210 11540
rect 2240 11510 2370 11540
rect 2200 11490 2370 11510
rect 2400 11610 2570 11630
rect 2400 11580 2410 11610
rect 2440 11580 2570 11610
rect 2400 11540 2570 11580
rect 2400 11510 2410 11540
rect 2440 11510 2570 11540
rect 2400 11490 2570 11510
rect 2600 11610 2770 11630
rect 2600 11580 2610 11610
rect 2640 11580 2770 11610
rect 2600 11540 2770 11580
rect 2600 11510 2610 11540
rect 2640 11510 2770 11540
rect 2600 11490 2770 11510
rect 2800 11610 2970 11630
rect 2800 11580 2810 11610
rect 2840 11580 2970 11610
rect 2800 11540 2970 11580
rect 2800 11510 2810 11540
rect 2840 11510 2970 11540
rect 2800 11490 2970 11510
rect 3000 11610 3170 11630
rect 3000 11580 3010 11610
rect 3040 11580 3170 11610
rect 3000 11540 3170 11580
rect 3000 11510 3010 11540
rect 3040 11510 3170 11540
rect 3000 11490 3170 11510
rect 3200 11610 3370 11630
rect 3200 11580 3210 11610
rect 3240 11580 3370 11610
rect 3200 11540 3370 11580
rect 3200 11510 3210 11540
rect 3240 11510 3370 11540
rect 3200 11490 3370 11510
rect 3400 11610 3570 11630
rect 3400 11580 3410 11610
rect 3440 11580 3570 11610
rect 3400 11540 3570 11580
rect 3400 11510 3410 11540
rect 3440 11510 3570 11540
rect 3400 11490 3570 11510
rect 3600 11610 3770 11630
rect 3600 11580 3610 11610
rect 3640 11580 3770 11610
rect 3600 11540 3770 11580
rect 3600 11510 3610 11540
rect 3640 11510 3770 11540
rect 3600 11490 3770 11510
rect 3800 11610 3970 11630
rect 3800 11580 3810 11610
rect 3840 11580 3970 11610
rect 3800 11540 3970 11580
rect 3800 11510 3810 11540
rect 3840 11510 3970 11540
rect 3800 11490 3970 11510
rect 4000 11610 4170 11630
rect 4000 11580 4010 11610
rect 4040 11580 4170 11610
rect 4000 11540 4170 11580
rect 4000 11510 4010 11540
rect 4040 11510 4170 11540
rect 4000 11490 4170 11510
rect 4200 11610 4370 11630
rect 4200 11580 4210 11610
rect 4240 11580 4370 11610
rect 4200 11540 4370 11580
rect 4200 11510 4210 11540
rect 4240 11510 4370 11540
rect 4200 11490 4370 11510
rect 4400 11610 4570 11630
rect 4400 11580 4410 11610
rect 4440 11580 4570 11610
rect 4400 11540 4570 11580
rect 4400 11510 4410 11540
rect 4440 11510 4570 11540
rect 4400 11490 4570 11510
rect 4600 11610 4770 11630
rect 4600 11580 4610 11610
rect 4640 11580 4770 11610
rect 4600 11540 4770 11580
rect 4600 11510 4610 11540
rect 4640 11510 4770 11540
rect 4600 11490 4770 11510
rect 4800 11610 4970 11630
rect 4800 11580 4810 11610
rect 4840 11580 4970 11610
rect 4800 11540 4970 11580
rect 4800 11510 4810 11540
rect 4840 11510 4970 11540
rect 4800 11490 4970 11510
rect 5000 11610 5170 11630
rect 5000 11580 5010 11610
rect 5040 11580 5170 11610
rect 5000 11540 5170 11580
rect 5000 11510 5010 11540
rect 5040 11510 5170 11540
rect 5000 11490 5170 11510
rect 5200 11610 5370 11630
rect 5200 11580 5210 11610
rect 5240 11580 5370 11610
rect 5200 11540 5370 11580
rect 5200 11510 5210 11540
rect 5240 11510 5370 11540
rect 5200 11490 5370 11510
rect 5400 11610 5570 11630
rect 5400 11580 5410 11610
rect 5440 11580 5570 11610
rect 5400 11540 5570 11580
rect 5400 11510 5410 11540
rect 5440 11510 5570 11540
rect 5400 11490 5570 11510
rect 5600 11610 5770 11630
rect 5600 11580 5610 11610
rect 5640 11580 5770 11610
rect 5600 11540 5770 11580
rect 5600 11510 5610 11540
rect 5640 11510 5770 11540
rect 5600 11490 5770 11510
rect 5800 11610 5970 11630
rect 5800 11580 5810 11610
rect 5840 11580 5970 11610
rect 5800 11540 5970 11580
rect 5800 11510 5810 11540
rect 5840 11510 5970 11540
rect 5800 11490 5970 11510
rect 6000 11610 6170 11630
rect 6000 11580 6010 11610
rect 6040 11580 6170 11610
rect 6000 11540 6170 11580
rect 6000 11510 6010 11540
rect 6040 11510 6170 11540
rect 6000 11490 6170 11510
rect 6200 11610 6370 11630
rect 6200 11580 6210 11610
rect 6240 11580 6370 11610
rect 6200 11540 6370 11580
rect 6200 11510 6210 11540
rect 6240 11510 6370 11540
rect 6200 11490 6370 11510
rect 6400 11610 6570 11630
rect 6400 11580 6410 11610
rect 6440 11580 6570 11610
rect 6400 11540 6570 11580
rect 6400 11510 6410 11540
rect 6440 11510 6570 11540
rect 6400 11490 6570 11510
rect -200 11425 -30 11445
rect -200 11395 -190 11425
rect -160 11395 -30 11425
rect -200 11355 -30 11395
rect -200 11325 -190 11355
rect -160 11325 -30 11355
rect -200 11305 -30 11325
rect 0 11425 170 11445
rect 0 11395 10 11425
rect 40 11395 170 11425
rect 0 11355 170 11395
rect 0 11325 10 11355
rect 40 11325 170 11355
rect 0 11305 170 11325
rect 200 11425 370 11445
rect 200 11395 210 11425
rect 240 11395 370 11425
rect 200 11355 370 11395
rect 200 11325 210 11355
rect 240 11325 370 11355
rect 200 11305 370 11325
rect 400 11425 570 11445
rect 400 11395 410 11425
rect 440 11395 570 11425
rect 400 11355 570 11395
rect 400 11325 410 11355
rect 440 11325 570 11355
rect 400 11305 570 11325
rect 600 11425 770 11445
rect 600 11395 610 11425
rect 640 11395 770 11425
rect 600 11355 770 11395
rect 600 11325 610 11355
rect 640 11325 770 11355
rect 600 11305 770 11325
rect 800 11425 970 11445
rect 800 11395 810 11425
rect 840 11395 970 11425
rect 800 11355 970 11395
rect 800 11325 810 11355
rect 840 11325 970 11355
rect 800 11305 970 11325
rect 1000 11425 1170 11445
rect 1000 11395 1010 11425
rect 1040 11395 1170 11425
rect 1000 11355 1170 11395
rect 1000 11325 1010 11355
rect 1040 11325 1170 11355
rect 1000 11305 1170 11325
rect 1200 11425 1370 11445
rect 1200 11395 1210 11425
rect 1240 11395 1370 11425
rect 1200 11355 1370 11395
rect 1200 11325 1210 11355
rect 1240 11325 1370 11355
rect 1200 11305 1370 11325
rect 1400 11425 1570 11445
rect 1400 11395 1410 11425
rect 1440 11395 1570 11425
rect 1400 11355 1570 11395
rect 1400 11325 1410 11355
rect 1440 11325 1570 11355
rect 1400 11305 1570 11325
rect 1600 11425 1770 11445
rect 1600 11395 1610 11425
rect 1640 11395 1770 11425
rect 1600 11355 1770 11395
rect 1600 11325 1610 11355
rect 1640 11325 1770 11355
rect 1600 11305 1770 11325
rect 1800 11425 1970 11445
rect 1800 11395 1810 11425
rect 1840 11395 1970 11425
rect 1800 11355 1970 11395
rect 1800 11325 1810 11355
rect 1840 11325 1970 11355
rect 1800 11305 1970 11325
rect 2000 11425 2170 11445
rect 2000 11395 2010 11425
rect 2040 11395 2170 11425
rect 2000 11355 2170 11395
rect 2000 11325 2010 11355
rect 2040 11325 2170 11355
rect 2000 11305 2170 11325
rect 2200 11425 2370 11445
rect 2200 11395 2210 11425
rect 2240 11395 2370 11425
rect 2200 11355 2370 11395
rect 2200 11325 2210 11355
rect 2240 11325 2370 11355
rect 2200 11305 2370 11325
rect 2400 11425 2570 11445
rect 2400 11395 2410 11425
rect 2440 11395 2570 11425
rect 2400 11355 2570 11395
rect 2400 11325 2410 11355
rect 2440 11325 2570 11355
rect 2400 11305 2570 11325
rect 2600 11425 2770 11445
rect 2600 11395 2610 11425
rect 2640 11395 2770 11425
rect 2600 11355 2770 11395
rect 2600 11325 2610 11355
rect 2640 11325 2770 11355
rect 2600 11305 2770 11325
rect 2800 11425 2970 11445
rect 2800 11395 2810 11425
rect 2840 11395 2970 11425
rect 2800 11355 2970 11395
rect 2800 11325 2810 11355
rect 2840 11325 2970 11355
rect 2800 11305 2970 11325
rect 3000 11425 3170 11445
rect 3000 11395 3010 11425
rect 3040 11395 3170 11425
rect 3000 11355 3170 11395
rect 3000 11325 3010 11355
rect 3040 11325 3170 11355
rect 3000 11305 3170 11325
rect 3200 11425 3370 11445
rect 3200 11395 3210 11425
rect 3240 11395 3370 11425
rect 3200 11355 3370 11395
rect 3200 11325 3210 11355
rect 3240 11325 3370 11355
rect 3200 11305 3370 11325
rect 3400 11425 3570 11445
rect 3400 11395 3410 11425
rect 3440 11395 3570 11425
rect 3400 11355 3570 11395
rect 3400 11325 3410 11355
rect 3440 11325 3570 11355
rect 3400 11305 3570 11325
rect 3600 11425 3770 11445
rect 3600 11395 3610 11425
rect 3640 11395 3770 11425
rect 3600 11355 3770 11395
rect 3600 11325 3610 11355
rect 3640 11325 3770 11355
rect 3600 11305 3770 11325
rect 3800 11425 3970 11445
rect 3800 11395 3810 11425
rect 3840 11395 3970 11425
rect 3800 11355 3970 11395
rect 3800 11325 3810 11355
rect 3840 11325 3970 11355
rect 3800 11305 3970 11325
rect 4000 11425 4170 11445
rect 4000 11395 4010 11425
rect 4040 11395 4170 11425
rect 4000 11355 4170 11395
rect 4000 11325 4010 11355
rect 4040 11325 4170 11355
rect 4000 11305 4170 11325
rect 4200 11425 4370 11445
rect 4200 11395 4210 11425
rect 4240 11395 4370 11425
rect 4200 11355 4370 11395
rect 4200 11325 4210 11355
rect 4240 11325 4370 11355
rect 4200 11305 4370 11325
rect 4400 11425 4570 11445
rect 4400 11395 4410 11425
rect 4440 11395 4570 11425
rect 4400 11355 4570 11395
rect 4400 11325 4410 11355
rect 4440 11325 4570 11355
rect 4400 11305 4570 11325
rect 4600 11425 4770 11445
rect 4600 11395 4610 11425
rect 4640 11395 4770 11425
rect 4600 11355 4770 11395
rect 4600 11325 4610 11355
rect 4640 11325 4770 11355
rect 4600 11305 4770 11325
rect 4800 11425 4970 11445
rect 4800 11395 4810 11425
rect 4840 11395 4970 11425
rect 4800 11355 4970 11395
rect 4800 11325 4810 11355
rect 4840 11325 4970 11355
rect 4800 11305 4970 11325
rect 5000 11425 5170 11445
rect 5000 11395 5010 11425
rect 5040 11395 5170 11425
rect 5000 11355 5170 11395
rect 5000 11325 5010 11355
rect 5040 11325 5170 11355
rect 5000 11305 5170 11325
rect 5200 11425 5370 11445
rect 5200 11395 5210 11425
rect 5240 11395 5370 11425
rect 5200 11355 5370 11395
rect 5200 11325 5210 11355
rect 5240 11325 5370 11355
rect 5200 11305 5370 11325
rect 5400 11425 5570 11445
rect 5400 11395 5410 11425
rect 5440 11395 5570 11425
rect 5400 11355 5570 11395
rect 5400 11325 5410 11355
rect 5440 11325 5570 11355
rect 5400 11305 5570 11325
rect 5600 11425 5770 11445
rect 5600 11395 5610 11425
rect 5640 11395 5770 11425
rect 5600 11355 5770 11395
rect 5600 11325 5610 11355
rect 5640 11325 5770 11355
rect 5600 11305 5770 11325
rect 5800 11425 5970 11445
rect 5800 11395 5810 11425
rect 5840 11395 5970 11425
rect 5800 11355 5970 11395
rect 5800 11325 5810 11355
rect 5840 11325 5970 11355
rect 5800 11305 5970 11325
rect 6000 11425 6170 11445
rect 6000 11395 6010 11425
rect 6040 11395 6170 11425
rect 6000 11355 6170 11395
rect 6000 11325 6010 11355
rect 6040 11325 6170 11355
rect 6000 11305 6170 11325
rect 6200 11425 6370 11445
rect 6200 11395 6210 11425
rect 6240 11395 6370 11425
rect 6200 11355 6370 11395
rect 6200 11325 6210 11355
rect 6240 11325 6370 11355
rect 6200 11305 6370 11325
rect 6400 11425 6570 11445
rect 6400 11395 6410 11425
rect 6440 11395 6570 11425
rect 6400 11355 6570 11395
rect 6400 11325 6410 11355
rect 6440 11325 6570 11355
rect 6400 11305 6570 11325
rect -200 11240 -30 11260
rect -200 11210 -190 11240
rect -160 11210 -30 11240
rect -200 11170 -30 11210
rect -200 11140 -190 11170
rect -160 11140 -30 11170
rect -200 11120 -30 11140
rect 0 11240 170 11260
rect 0 11210 10 11240
rect 40 11210 170 11240
rect 0 11170 170 11210
rect 0 11140 10 11170
rect 40 11140 170 11170
rect 0 11120 170 11140
rect 200 11240 370 11260
rect 200 11210 210 11240
rect 240 11210 370 11240
rect 200 11170 370 11210
rect 200 11140 210 11170
rect 240 11140 370 11170
rect 200 11120 370 11140
rect 400 11240 570 11260
rect 400 11210 410 11240
rect 440 11210 570 11240
rect 400 11170 570 11210
rect 400 11140 410 11170
rect 440 11140 570 11170
rect 400 11120 570 11140
rect 600 11240 770 11260
rect 600 11210 610 11240
rect 640 11210 770 11240
rect 600 11170 770 11210
rect 600 11140 610 11170
rect 640 11140 770 11170
rect 600 11120 770 11140
rect 800 11240 970 11260
rect 800 11210 810 11240
rect 840 11210 970 11240
rect 800 11170 970 11210
rect 800 11140 810 11170
rect 840 11140 970 11170
rect 800 11120 970 11140
rect 1000 11240 1170 11260
rect 1000 11210 1010 11240
rect 1040 11210 1170 11240
rect 1000 11170 1170 11210
rect 1000 11140 1010 11170
rect 1040 11140 1170 11170
rect 1000 11120 1170 11140
rect 1200 11240 1370 11260
rect 1200 11210 1210 11240
rect 1240 11210 1370 11240
rect 1200 11170 1370 11210
rect 1200 11140 1210 11170
rect 1240 11140 1370 11170
rect 1200 11120 1370 11140
rect 1400 11240 1570 11260
rect 1400 11210 1410 11240
rect 1440 11210 1570 11240
rect 1400 11170 1570 11210
rect 1400 11140 1410 11170
rect 1440 11140 1570 11170
rect 1400 11120 1570 11140
rect 1600 11240 1770 11260
rect 1600 11210 1610 11240
rect 1640 11210 1770 11240
rect 1600 11170 1770 11210
rect 1600 11140 1610 11170
rect 1640 11140 1770 11170
rect 1600 11120 1770 11140
rect 1800 11240 1970 11260
rect 1800 11210 1810 11240
rect 1840 11210 1970 11240
rect 1800 11170 1970 11210
rect 1800 11140 1810 11170
rect 1840 11140 1970 11170
rect 1800 11120 1970 11140
rect 2000 11240 2170 11260
rect 2000 11210 2010 11240
rect 2040 11210 2170 11240
rect 2000 11170 2170 11210
rect 2000 11140 2010 11170
rect 2040 11140 2170 11170
rect 2000 11120 2170 11140
rect 2200 11240 2370 11260
rect 2200 11210 2210 11240
rect 2240 11210 2370 11240
rect 2200 11170 2370 11210
rect 2200 11140 2210 11170
rect 2240 11140 2370 11170
rect 2200 11120 2370 11140
rect 2400 11240 2570 11260
rect 2400 11210 2410 11240
rect 2440 11210 2570 11240
rect 2400 11170 2570 11210
rect 2400 11140 2410 11170
rect 2440 11140 2570 11170
rect 2400 11120 2570 11140
rect 2600 11240 2770 11260
rect 2600 11210 2610 11240
rect 2640 11210 2770 11240
rect 2600 11170 2770 11210
rect 2600 11140 2610 11170
rect 2640 11140 2770 11170
rect 2600 11120 2770 11140
rect 2800 11240 2970 11260
rect 2800 11210 2810 11240
rect 2840 11210 2970 11240
rect 2800 11170 2970 11210
rect 2800 11140 2810 11170
rect 2840 11140 2970 11170
rect 2800 11120 2970 11140
rect 3000 11240 3170 11260
rect 3000 11210 3010 11240
rect 3040 11210 3170 11240
rect 3000 11170 3170 11210
rect 3000 11140 3010 11170
rect 3040 11140 3170 11170
rect 3000 11120 3170 11140
rect 3200 11240 3370 11260
rect 3200 11210 3210 11240
rect 3240 11210 3370 11240
rect 3200 11170 3370 11210
rect 3200 11140 3210 11170
rect 3240 11140 3370 11170
rect 3200 11120 3370 11140
rect 3400 11240 3570 11260
rect 3400 11210 3410 11240
rect 3440 11210 3570 11240
rect 3400 11170 3570 11210
rect 3400 11140 3410 11170
rect 3440 11140 3570 11170
rect 3400 11120 3570 11140
rect 3600 11240 3770 11260
rect 3600 11210 3610 11240
rect 3640 11210 3770 11240
rect 3600 11170 3770 11210
rect 3600 11140 3610 11170
rect 3640 11140 3770 11170
rect 3600 11120 3770 11140
rect 3800 11240 3970 11260
rect 3800 11210 3810 11240
rect 3840 11210 3970 11240
rect 3800 11170 3970 11210
rect 3800 11140 3810 11170
rect 3840 11140 3970 11170
rect 3800 11120 3970 11140
rect 4000 11240 4170 11260
rect 4000 11210 4010 11240
rect 4040 11210 4170 11240
rect 4000 11170 4170 11210
rect 4000 11140 4010 11170
rect 4040 11140 4170 11170
rect 4000 11120 4170 11140
rect 4200 11240 4370 11260
rect 4200 11210 4210 11240
rect 4240 11210 4370 11240
rect 4200 11170 4370 11210
rect 4200 11140 4210 11170
rect 4240 11140 4370 11170
rect 4200 11120 4370 11140
rect 4400 11240 4570 11260
rect 4400 11210 4410 11240
rect 4440 11210 4570 11240
rect 4400 11170 4570 11210
rect 4400 11140 4410 11170
rect 4440 11140 4570 11170
rect 4400 11120 4570 11140
rect 4600 11240 4770 11260
rect 4600 11210 4610 11240
rect 4640 11210 4770 11240
rect 4600 11170 4770 11210
rect 4600 11140 4610 11170
rect 4640 11140 4770 11170
rect 4600 11120 4770 11140
rect 4800 11240 4970 11260
rect 4800 11210 4810 11240
rect 4840 11210 4970 11240
rect 4800 11170 4970 11210
rect 4800 11140 4810 11170
rect 4840 11140 4970 11170
rect 4800 11120 4970 11140
rect 5000 11240 5170 11260
rect 5000 11210 5010 11240
rect 5040 11210 5170 11240
rect 5000 11170 5170 11210
rect 5000 11140 5010 11170
rect 5040 11140 5170 11170
rect 5000 11120 5170 11140
rect 5200 11240 5370 11260
rect 5200 11210 5210 11240
rect 5240 11210 5370 11240
rect 5200 11170 5370 11210
rect 5200 11140 5210 11170
rect 5240 11140 5370 11170
rect 5200 11120 5370 11140
rect 5400 11240 5570 11260
rect 5400 11210 5410 11240
rect 5440 11210 5570 11240
rect 5400 11170 5570 11210
rect 5400 11140 5410 11170
rect 5440 11140 5570 11170
rect 5400 11120 5570 11140
rect 5600 11240 5770 11260
rect 5600 11210 5610 11240
rect 5640 11210 5770 11240
rect 5600 11170 5770 11210
rect 5600 11140 5610 11170
rect 5640 11140 5770 11170
rect 5600 11120 5770 11140
rect 5800 11240 5970 11260
rect 5800 11210 5810 11240
rect 5840 11210 5970 11240
rect 5800 11170 5970 11210
rect 5800 11140 5810 11170
rect 5840 11140 5970 11170
rect 5800 11120 5970 11140
rect 6000 11240 6170 11260
rect 6000 11210 6010 11240
rect 6040 11210 6170 11240
rect 6000 11170 6170 11210
rect 6000 11140 6010 11170
rect 6040 11140 6170 11170
rect 6000 11120 6170 11140
rect 6200 11240 6370 11260
rect 6200 11210 6210 11240
rect 6240 11210 6370 11240
rect 6200 11170 6370 11210
rect 6200 11140 6210 11170
rect 6240 11140 6370 11170
rect 6200 11120 6370 11140
rect 6400 11240 6570 11260
rect 6400 11210 6410 11240
rect 6440 11210 6570 11240
rect 6400 11170 6570 11210
rect 6400 11140 6410 11170
rect 6440 11140 6570 11170
rect 6400 11120 6570 11140
rect -200 11055 -30 11075
rect -200 11025 -190 11055
rect -160 11025 -30 11055
rect -200 10985 -30 11025
rect -200 10955 -190 10985
rect -160 10955 -30 10985
rect -200 10935 -30 10955
rect 0 11055 170 11075
rect 0 11025 10 11055
rect 40 11025 170 11055
rect 0 10985 170 11025
rect 0 10955 10 10985
rect 40 10955 170 10985
rect 0 10935 170 10955
rect 200 11055 370 11075
rect 200 11025 210 11055
rect 240 11025 370 11055
rect 200 10985 370 11025
rect 200 10955 210 10985
rect 240 10955 370 10985
rect 200 10935 370 10955
rect 400 11055 570 11075
rect 400 11025 410 11055
rect 440 11025 570 11055
rect 400 10985 570 11025
rect 400 10955 410 10985
rect 440 10955 570 10985
rect 400 10935 570 10955
rect 600 11055 770 11075
rect 600 11025 610 11055
rect 640 11025 770 11055
rect 600 10985 770 11025
rect 600 10955 610 10985
rect 640 10955 770 10985
rect 600 10935 770 10955
rect 800 11055 970 11075
rect 800 11025 810 11055
rect 840 11025 970 11055
rect 800 10985 970 11025
rect 800 10955 810 10985
rect 840 10955 970 10985
rect 800 10935 970 10955
rect 1000 11055 1170 11075
rect 1000 11025 1010 11055
rect 1040 11025 1170 11055
rect 1000 10985 1170 11025
rect 1000 10955 1010 10985
rect 1040 10955 1170 10985
rect 1000 10935 1170 10955
rect 1200 11055 1370 11075
rect 1200 11025 1210 11055
rect 1240 11025 1370 11055
rect 1200 10985 1370 11025
rect 1200 10955 1210 10985
rect 1240 10955 1370 10985
rect 1200 10935 1370 10955
rect 1400 11055 1570 11075
rect 1400 11025 1410 11055
rect 1440 11025 1570 11055
rect 1400 10985 1570 11025
rect 1400 10955 1410 10985
rect 1440 10955 1570 10985
rect 1400 10935 1570 10955
rect 1600 11055 1770 11075
rect 1600 11025 1610 11055
rect 1640 11025 1770 11055
rect 1600 10985 1770 11025
rect 1600 10955 1610 10985
rect 1640 10955 1770 10985
rect 1600 10935 1770 10955
rect 1800 11055 1970 11075
rect 1800 11025 1810 11055
rect 1840 11025 1970 11055
rect 1800 10985 1970 11025
rect 1800 10955 1810 10985
rect 1840 10955 1970 10985
rect 1800 10935 1970 10955
rect 2000 11055 2170 11075
rect 2000 11025 2010 11055
rect 2040 11025 2170 11055
rect 2000 10985 2170 11025
rect 2000 10955 2010 10985
rect 2040 10955 2170 10985
rect 2000 10935 2170 10955
rect 2200 11055 2370 11075
rect 2200 11025 2210 11055
rect 2240 11025 2370 11055
rect 2200 10985 2370 11025
rect 2200 10955 2210 10985
rect 2240 10955 2370 10985
rect 2200 10935 2370 10955
rect 2400 11055 2570 11075
rect 2400 11025 2410 11055
rect 2440 11025 2570 11055
rect 2400 10985 2570 11025
rect 2400 10955 2410 10985
rect 2440 10955 2570 10985
rect 2400 10935 2570 10955
rect 2600 11055 2770 11075
rect 2600 11025 2610 11055
rect 2640 11025 2770 11055
rect 2600 10985 2770 11025
rect 2600 10955 2610 10985
rect 2640 10955 2770 10985
rect 2600 10935 2770 10955
rect 2800 11055 2970 11075
rect 2800 11025 2810 11055
rect 2840 11025 2970 11055
rect 2800 10985 2970 11025
rect 2800 10955 2810 10985
rect 2840 10955 2970 10985
rect 2800 10935 2970 10955
rect 3000 11055 3170 11075
rect 3000 11025 3010 11055
rect 3040 11025 3170 11055
rect 3000 10985 3170 11025
rect 3000 10955 3010 10985
rect 3040 10955 3170 10985
rect 3000 10935 3170 10955
rect 3200 11055 3370 11075
rect 3200 11025 3210 11055
rect 3240 11025 3370 11055
rect 3200 10985 3370 11025
rect 3200 10955 3210 10985
rect 3240 10955 3370 10985
rect 3200 10935 3370 10955
rect 3400 11055 3570 11075
rect 3400 11025 3410 11055
rect 3440 11025 3570 11055
rect 3400 10985 3570 11025
rect 3400 10955 3410 10985
rect 3440 10955 3570 10985
rect 3400 10935 3570 10955
rect 3600 11055 3770 11075
rect 3600 11025 3610 11055
rect 3640 11025 3770 11055
rect 3600 10985 3770 11025
rect 3600 10955 3610 10985
rect 3640 10955 3770 10985
rect 3600 10935 3770 10955
rect 3800 11055 3970 11075
rect 3800 11025 3810 11055
rect 3840 11025 3970 11055
rect 3800 10985 3970 11025
rect 3800 10955 3810 10985
rect 3840 10955 3970 10985
rect 3800 10935 3970 10955
rect 4000 11055 4170 11075
rect 4000 11025 4010 11055
rect 4040 11025 4170 11055
rect 4000 10985 4170 11025
rect 4000 10955 4010 10985
rect 4040 10955 4170 10985
rect 4000 10935 4170 10955
rect 4200 11055 4370 11075
rect 4200 11025 4210 11055
rect 4240 11025 4370 11055
rect 4200 10985 4370 11025
rect 4200 10955 4210 10985
rect 4240 10955 4370 10985
rect 4200 10935 4370 10955
rect 4400 11055 4570 11075
rect 4400 11025 4410 11055
rect 4440 11025 4570 11055
rect 4400 10985 4570 11025
rect 4400 10955 4410 10985
rect 4440 10955 4570 10985
rect 4400 10935 4570 10955
rect 4600 11055 4770 11075
rect 4600 11025 4610 11055
rect 4640 11025 4770 11055
rect 4600 10985 4770 11025
rect 4600 10955 4610 10985
rect 4640 10955 4770 10985
rect 4600 10935 4770 10955
rect 4800 11055 4970 11075
rect 4800 11025 4810 11055
rect 4840 11025 4970 11055
rect 4800 10985 4970 11025
rect 4800 10955 4810 10985
rect 4840 10955 4970 10985
rect 4800 10935 4970 10955
rect 5000 11055 5170 11075
rect 5000 11025 5010 11055
rect 5040 11025 5170 11055
rect 5000 10985 5170 11025
rect 5000 10955 5010 10985
rect 5040 10955 5170 10985
rect 5000 10935 5170 10955
rect 5200 11055 5370 11075
rect 5200 11025 5210 11055
rect 5240 11025 5370 11055
rect 5200 10985 5370 11025
rect 5200 10955 5210 10985
rect 5240 10955 5370 10985
rect 5200 10935 5370 10955
rect 5400 11055 5570 11075
rect 5400 11025 5410 11055
rect 5440 11025 5570 11055
rect 5400 10985 5570 11025
rect 5400 10955 5410 10985
rect 5440 10955 5570 10985
rect 5400 10935 5570 10955
rect 5600 11055 5770 11075
rect 5600 11025 5610 11055
rect 5640 11025 5770 11055
rect 5600 10985 5770 11025
rect 5600 10955 5610 10985
rect 5640 10955 5770 10985
rect 5600 10935 5770 10955
rect 5800 11055 5970 11075
rect 5800 11025 5810 11055
rect 5840 11025 5970 11055
rect 5800 10985 5970 11025
rect 5800 10955 5810 10985
rect 5840 10955 5970 10985
rect 5800 10935 5970 10955
rect 6000 11055 6170 11075
rect 6000 11025 6010 11055
rect 6040 11025 6170 11055
rect 6000 10985 6170 11025
rect 6000 10955 6010 10985
rect 6040 10955 6170 10985
rect 6000 10935 6170 10955
rect 6200 11055 6370 11075
rect 6200 11025 6210 11055
rect 6240 11025 6370 11055
rect 6200 10985 6370 11025
rect 6200 10955 6210 10985
rect 6240 10955 6370 10985
rect 6200 10935 6370 10955
rect 6400 11055 6570 11075
rect 6400 11025 6410 11055
rect 6440 11025 6570 11055
rect 6400 10985 6570 11025
rect 6400 10955 6410 10985
rect 6440 10955 6570 10985
rect 6400 10935 6570 10955
rect -200 10870 -30 10890
rect -200 10840 -190 10870
rect -160 10840 -30 10870
rect -200 10800 -30 10840
rect -200 10770 -190 10800
rect -160 10770 -30 10800
rect -200 10750 -30 10770
rect 0 10870 170 10890
rect 0 10840 10 10870
rect 40 10840 170 10870
rect 0 10800 170 10840
rect 0 10770 10 10800
rect 40 10770 170 10800
rect 0 10750 170 10770
rect 200 10870 370 10890
rect 200 10840 210 10870
rect 240 10840 370 10870
rect 200 10800 370 10840
rect 200 10770 210 10800
rect 240 10770 370 10800
rect 200 10750 370 10770
rect 400 10870 570 10890
rect 400 10840 410 10870
rect 440 10840 570 10870
rect 400 10800 570 10840
rect 400 10770 410 10800
rect 440 10770 570 10800
rect 400 10750 570 10770
rect 600 10870 770 10890
rect 600 10840 610 10870
rect 640 10840 770 10870
rect 600 10800 770 10840
rect 600 10770 610 10800
rect 640 10770 770 10800
rect 600 10750 770 10770
rect 800 10870 970 10890
rect 800 10840 810 10870
rect 840 10840 970 10870
rect 800 10800 970 10840
rect 800 10770 810 10800
rect 840 10770 970 10800
rect 800 10750 970 10770
rect 1000 10870 1170 10890
rect 1000 10840 1010 10870
rect 1040 10840 1170 10870
rect 1000 10800 1170 10840
rect 1000 10770 1010 10800
rect 1040 10770 1170 10800
rect 1000 10750 1170 10770
rect 1200 10870 1370 10890
rect 1200 10840 1210 10870
rect 1240 10840 1370 10870
rect 1200 10800 1370 10840
rect 1200 10770 1210 10800
rect 1240 10770 1370 10800
rect 1200 10750 1370 10770
rect 1400 10870 1570 10890
rect 1400 10840 1410 10870
rect 1440 10840 1570 10870
rect 1400 10800 1570 10840
rect 1400 10770 1410 10800
rect 1440 10770 1570 10800
rect 1400 10750 1570 10770
rect 1600 10870 1770 10890
rect 1600 10840 1610 10870
rect 1640 10840 1770 10870
rect 1600 10800 1770 10840
rect 1600 10770 1610 10800
rect 1640 10770 1770 10800
rect 1600 10750 1770 10770
rect 1800 10870 1970 10890
rect 1800 10840 1810 10870
rect 1840 10840 1970 10870
rect 1800 10800 1970 10840
rect 1800 10770 1810 10800
rect 1840 10770 1970 10800
rect 1800 10750 1970 10770
rect 2000 10870 2170 10890
rect 2000 10840 2010 10870
rect 2040 10840 2170 10870
rect 2000 10800 2170 10840
rect 2000 10770 2010 10800
rect 2040 10770 2170 10800
rect 2000 10750 2170 10770
rect 2200 10870 2370 10890
rect 2200 10840 2210 10870
rect 2240 10840 2370 10870
rect 2200 10800 2370 10840
rect 2200 10770 2210 10800
rect 2240 10770 2370 10800
rect 2200 10750 2370 10770
rect 2400 10870 2570 10890
rect 2400 10840 2410 10870
rect 2440 10840 2570 10870
rect 2400 10800 2570 10840
rect 2400 10770 2410 10800
rect 2440 10770 2570 10800
rect 2400 10750 2570 10770
rect 2600 10870 2770 10890
rect 2600 10840 2610 10870
rect 2640 10840 2770 10870
rect 2600 10800 2770 10840
rect 2600 10770 2610 10800
rect 2640 10770 2770 10800
rect 2600 10750 2770 10770
rect 2800 10870 2970 10890
rect 2800 10840 2810 10870
rect 2840 10840 2970 10870
rect 2800 10800 2970 10840
rect 2800 10770 2810 10800
rect 2840 10770 2970 10800
rect 2800 10750 2970 10770
rect 3000 10870 3170 10890
rect 3000 10840 3010 10870
rect 3040 10840 3170 10870
rect 3000 10800 3170 10840
rect 3000 10770 3010 10800
rect 3040 10770 3170 10800
rect 3000 10750 3170 10770
rect 3200 10870 3370 10890
rect 3200 10840 3210 10870
rect 3240 10840 3370 10870
rect 3200 10800 3370 10840
rect 3200 10770 3210 10800
rect 3240 10770 3370 10800
rect 3200 10750 3370 10770
rect 3400 10870 3570 10890
rect 3400 10840 3410 10870
rect 3440 10840 3570 10870
rect 3400 10800 3570 10840
rect 3400 10770 3410 10800
rect 3440 10770 3570 10800
rect 3400 10750 3570 10770
rect 3600 10870 3770 10890
rect 3600 10840 3610 10870
rect 3640 10840 3770 10870
rect 3600 10800 3770 10840
rect 3600 10770 3610 10800
rect 3640 10770 3770 10800
rect 3600 10750 3770 10770
rect 3800 10870 3970 10890
rect 3800 10840 3810 10870
rect 3840 10840 3970 10870
rect 3800 10800 3970 10840
rect 3800 10770 3810 10800
rect 3840 10770 3970 10800
rect 3800 10750 3970 10770
rect 4000 10870 4170 10890
rect 4000 10840 4010 10870
rect 4040 10840 4170 10870
rect 4000 10800 4170 10840
rect 4000 10770 4010 10800
rect 4040 10770 4170 10800
rect 4000 10750 4170 10770
rect 4200 10870 4370 10890
rect 4200 10840 4210 10870
rect 4240 10840 4370 10870
rect 4200 10800 4370 10840
rect 4200 10770 4210 10800
rect 4240 10770 4370 10800
rect 4200 10750 4370 10770
rect 4400 10870 4570 10890
rect 4400 10840 4410 10870
rect 4440 10840 4570 10870
rect 4400 10800 4570 10840
rect 4400 10770 4410 10800
rect 4440 10770 4570 10800
rect 4400 10750 4570 10770
rect 4600 10870 4770 10890
rect 4600 10840 4610 10870
rect 4640 10840 4770 10870
rect 4600 10800 4770 10840
rect 4600 10770 4610 10800
rect 4640 10770 4770 10800
rect 4600 10750 4770 10770
rect 4800 10870 4970 10890
rect 4800 10840 4810 10870
rect 4840 10840 4970 10870
rect 4800 10800 4970 10840
rect 4800 10770 4810 10800
rect 4840 10770 4970 10800
rect 4800 10750 4970 10770
rect 5000 10870 5170 10890
rect 5000 10840 5010 10870
rect 5040 10840 5170 10870
rect 5000 10800 5170 10840
rect 5000 10770 5010 10800
rect 5040 10770 5170 10800
rect 5000 10750 5170 10770
rect 5200 10870 5370 10890
rect 5200 10840 5210 10870
rect 5240 10840 5370 10870
rect 5200 10800 5370 10840
rect 5200 10770 5210 10800
rect 5240 10770 5370 10800
rect 5200 10750 5370 10770
rect 5400 10870 5570 10890
rect 5400 10840 5410 10870
rect 5440 10840 5570 10870
rect 5400 10800 5570 10840
rect 5400 10770 5410 10800
rect 5440 10770 5570 10800
rect 5400 10750 5570 10770
rect 5600 10870 5770 10890
rect 5600 10840 5610 10870
rect 5640 10840 5770 10870
rect 5600 10800 5770 10840
rect 5600 10770 5610 10800
rect 5640 10770 5770 10800
rect 5600 10750 5770 10770
rect 5800 10870 5970 10890
rect 5800 10840 5810 10870
rect 5840 10840 5970 10870
rect 5800 10800 5970 10840
rect 5800 10770 5810 10800
rect 5840 10770 5970 10800
rect 5800 10750 5970 10770
rect 6000 10870 6170 10890
rect 6000 10840 6010 10870
rect 6040 10840 6170 10870
rect 6000 10800 6170 10840
rect 6000 10770 6010 10800
rect 6040 10770 6170 10800
rect 6000 10750 6170 10770
rect 6200 10870 6370 10890
rect 6200 10840 6210 10870
rect 6240 10840 6370 10870
rect 6200 10800 6370 10840
rect 6200 10770 6210 10800
rect 6240 10770 6370 10800
rect 6200 10750 6370 10770
rect 6400 10870 6570 10890
rect 6400 10840 6410 10870
rect 6440 10840 6570 10870
rect 6400 10800 6570 10840
rect 6400 10770 6410 10800
rect 6440 10770 6570 10800
rect 6400 10750 6570 10770
rect -200 10685 -30 10705
rect -200 10655 -190 10685
rect -160 10655 -30 10685
rect -200 10615 -30 10655
rect -200 10585 -190 10615
rect -160 10585 -30 10615
rect -200 10565 -30 10585
rect 0 10685 170 10705
rect 0 10655 10 10685
rect 40 10655 170 10685
rect 0 10615 170 10655
rect 0 10585 10 10615
rect 40 10585 170 10615
rect 0 10565 170 10585
rect 200 10685 370 10705
rect 200 10655 210 10685
rect 240 10655 370 10685
rect 200 10615 370 10655
rect 200 10585 210 10615
rect 240 10585 370 10615
rect 200 10565 370 10585
rect 400 10685 570 10705
rect 400 10655 410 10685
rect 440 10655 570 10685
rect 400 10615 570 10655
rect 400 10585 410 10615
rect 440 10585 570 10615
rect 400 10565 570 10585
rect 600 10685 770 10705
rect 600 10655 610 10685
rect 640 10655 770 10685
rect 600 10615 770 10655
rect 600 10585 610 10615
rect 640 10585 770 10615
rect 600 10565 770 10585
rect 800 10685 970 10705
rect 800 10655 810 10685
rect 840 10655 970 10685
rect 800 10615 970 10655
rect 800 10585 810 10615
rect 840 10585 970 10615
rect 800 10565 970 10585
rect 1000 10685 1170 10705
rect 1000 10655 1010 10685
rect 1040 10655 1170 10685
rect 1000 10615 1170 10655
rect 1000 10585 1010 10615
rect 1040 10585 1170 10615
rect 1000 10565 1170 10585
rect 1200 10685 1370 10705
rect 1200 10655 1210 10685
rect 1240 10655 1370 10685
rect 1200 10615 1370 10655
rect 1200 10585 1210 10615
rect 1240 10585 1370 10615
rect 1200 10565 1370 10585
rect 1400 10685 1570 10705
rect 1400 10655 1410 10685
rect 1440 10655 1570 10685
rect 1400 10615 1570 10655
rect 1400 10585 1410 10615
rect 1440 10585 1570 10615
rect 1400 10565 1570 10585
rect 1600 10685 1770 10705
rect 1600 10655 1610 10685
rect 1640 10655 1770 10685
rect 1600 10615 1770 10655
rect 1600 10585 1610 10615
rect 1640 10585 1770 10615
rect 1600 10565 1770 10585
rect 1800 10685 1970 10705
rect 1800 10655 1810 10685
rect 1840 10655 1970 10685
rect 1800 10615 1970 10655
rect 1800 10585 1810 10615
rect 1840 10585 1970 10615
rect 1800 10565 1970 10585
rect 2000 10685 2170 10705
rect 2000 10655 2010 10685
rect 2040 10655 2170 10685
rect 2000 10615 2170 10655
rect 2000 10585 2010 10615
rect 2040 10585 2170 10615
rect 2000 10565 2170 10585
rect 2200 10685 2370 10705
rect 2200 10655 2210 10685
rect 2240 10655 2370 10685
rect 2200 10615 2370 10655
rect 2200 10585 2210 10615
rect 2240 10585 2370 10615
rect 2200 10565 2370 10585
rect 2400 10685 2570 10705
rect 2400 10655 2410 10685
rect 2440 10655 2570 10685
rect 2400 10615 2570 10655
rect 2400 10585 2410 10615
rect 2440 10585 2570 10615
rect 2400 10565 2570 10585
rect 2600 10685 2770 10705
rect 2600 10655 2610 10685
rect 2640 10655 2770 10685
rect 2600 10615 2770 10655
rect 2600 10585 2610 10615
rect 2640 10585 2770 10615
rect 2600 10565 2770 10585
rect 2800 10685 2970 10705
rect 2800 10655 2810 10685
rect 2840 10655 2970 10685
rect 2800 10615 2970 10655
rect 2800 10585 2810 10615
rect 2840 10585 2970 10615
rect 2800 10565 2970 10585
rect 3000 10685 3170 10705
rect 3000 10655 3010 10685
rect 3040 10655 3170 10685
rect 3000 10615 3170 10655
rect 3000 10585 3010 10615
rect 3040 10585 3170 10615
rect 3000 10565 3170 10585
rect 3200 10685 3370 10705
rect 3200 10655 3210 10685
rect 3240 10655 3370 10685
rect 3200 10615 3370 10655
rect 3200 10585 3210 10615
rect 3240 10585 3370 10615
rect 3200 10565 3370 10585
rect 3400 10685 3570 10705
rect 3400 10655 3410 10685
rect 3440 10655 3570 10685
rect 3400 10615 3570 10655
rect 3400 10585 3410 10615
rect 3440 10585 3570 10615
rect 3400 10565 3570 10585
rect 3600 10685 3770 10705
rect 3600 10655 3610 10685
rect 3640 10655 3770 10685
rect 3600 10615 3770 10655
rect 3600 10585 3610 10615
rect 3640 10585 3770 10615
rect 3600 10565 3770 10585
rect 3800 10685 3970 10705
rect 3800 10655 3810 10685
rect 3840 10655 3970 10685
rect 3800 10615 3970 10655
rect 3800 10585 3810 10615
rect 3840 10585 3970 10615
rect 3800 10565 3970 10585
rect 4000 10685 4170 10705
rect 4000 10655 4010 10685
rect 4040 10655 4170 10685
rect 4000 10615 4170 10655
rect 4000 10585 4010 10615
rect 4040 10585 4170 10615
rect 4000 10565 4170 10585
rect 4200 10685 4370 10705
rect 4200 10655 4210 10685
rect 4240 10655 4370 10685
rect 4200 10615 4370 10655
rect 4200 10585 4210 10615
rect 4240 10585 4370 10615
rect 4200 10565 4370 10585
rect 4400 10685 4570 10705
rect 4400 10655 4410 10685
rect 4440 10655 4570 10685
rect 4400 10615 4570 10655
rect 4400 10585 4410 10615
rect 4440 10585 4570 10615
rect 4400 10565 4570 10585
rect 4600 10685 4770 10705
rect 4600 10655 4610 10685
rect 4640 10655 4770 10685
rect 4600 10615 4770 10655
rect 4600 10585 4610 10615
rect 4640 10585 4770 10615
rect 4600 10565 4770 10585
rect 4800 10685 4970 10705
rect 4800 10655 4810 10685
rect 4840 10655 4970 10685
rect 4800 10615 4970 10655
rect 4800 10585 4810 10615
rect 4840 10585 4970 10615
rect 4800 10565 4970 10585
rect 5000 10685 5170 10705
rect 5000 10655 5010 10685
rect 5040 10655 5170 10685
rect 5000 10615 5170 10655
rect 5000 10585 5010 10615
rect 5040 10585 5170 10615
rect 5000 10565 5170 10585
rect 5200 10685 5370 10705
rect 5200 10655 5210 10685
rect 5240 10655 5370 10685
rect 5200 10615 5370 10655
rect 5200 10585 5210 10615
rect 5240 10585 5370 10615
rect 5200 10565 5370 10585
rect 5400 10685 5570 10705
rect 5400 10655 5410 10685
rect 5440 10655 5570 10685
rect 5400 10615 5570 10655
rect 5400 10585 5410 10615
rect 5440 10585 5570 10615
rect 5400 10565 5570 10585
rect 5600 10685 5770 10705
rect 5600 10655 5610 10685
rect 5640 10655 5770 10685
rect 5600 10615 5770 10655
rect 5600 10585 5610 10615
rect 5640 10585 5770 10615
rect 5600 10565 5770 10585
rect 5800 10685 5970 10705
rect 5800 10655 5810 10685
rect 5840 10655 5970 10685
rect 5800 10615 5970 10655
rect 5800 10585 5810 10615
rect 5840 10585 5970 10615
rect 5800 10565 5970 10585
rect 6000 10685 6170 10705
rect 6000 10655 6010 10685
rect 6040 10655 6170 10685
rect 6000 10615 6170 10655
rect 6000 10585 6010 10615
rect 6040 10585 6170 10615
rect 6000 10565 6170 10585
rect 6200 10685 6370 10705
rect 6200 10655 6210 10685
rect 6240 10655 6370 10685
rect 6200 10615 6370 10655
rect 6200 10585 6210 10615
rect 6240 10585 6370 10615
rect 6200 10565 6370 10585
rect 6400 10685 6570 10705
rect 6400 10655 6410 10685
rect 6440 10655 6570 10685
rect 6400 10615 6570 10655
rect 6400 10585 6410 10615
rect 6440 10585 6570 10615
rect 6400 10565 6570 10585
rect -200 10500 -30 10520
rect -200 10470 -190 10500
rect -160 10470 -30 10500
rect -200 10430 -30 10470
rect -200 10400 -190 10430
rect -160 10400 -30 10430
rect -200 10380 -30 10400
rect 0 10500 170 10520
rect 0 10470 10 10500
rect 40 10470 170 10500
rect 0 10430 170 10470
rect 0 10400 10 10430
rect 40 10400 170 10430
rect 0 10380 170 10400
rect 200 10500 370 10520
rect 200 10470 210 10500
rect 240 10470 370 10500
rect 200 10430 370 10470
rect 200 10400 210 10430
rect 240 10400 370 10430
rect 200 10380 370 10400
rect 400 10500 570 10520
rect 400 10470 410 10500
rect 440 10470 570 10500
rect 400 10430 570 10470
rect 400 10400 410 10430
rect 440 10400 570 10430
rect 400 10380 570 10400
rect 600 10500 770 10520
rect 600 10470 610 10500
rect 640 10470 770 10500
rect 600 10430 770 10470
rect 600 10400 610 10430
rect 640 10400 770 10430
rect 600 10380 770 10400
rect 800 10500 970 10520
rect 800 10470 810 10500
rect 840 10470 970 10500
rect 800 10430 970 10470
rect 800 10400 810 10430
rect 840 10400 970 10430
rect 800 10380 970 10400
rect 1000 10500 1170 10520
rect 1000 10470 1010 10500
rect 1040 10470 1170 10500
rect 1000 10430 1170 10470
rect 1000 10400 1010 10430
rect 1040 10400 1170 10430
rect 1000 10380 1170 10400
rect 1200 10500 1370 10520
rect 1200 10470 1210 10500
rect 1240 10470 1370 10500
rect 1200 10430 1370 10470
rect 1200 10400 1210 10430
rect 1240 10400 1370 10430
rect 1200 10380 1370 10400
rect 1400 10500 1570 10520
rect 1400 10470 1410 10500
rect 1440 10470 1570 10500
rect 1400 10430 1570 10470
rect 1400 10400 1410 10430
rect 1440 10400 1570 10430
rect 1400 10380 1570 10400
rect 1600 10500 1770 10520
rect 1600 10470 1610 10500
rect 1640 10470 1770 10500
rect 1600 10430 1770 10470
rect 1600 10400 1610 10430
rect 1640 10400 1770 10430
rect 1600 10380 1770 10400
rect 1800 10500 1970 10520
rect 1800 10470 1810 10500
rect 1840 10470 1970 10500
rect 1800 10430 1970 10470
rect 1800 10400 1810 10430
rect 1840 10400 1970 10430
rect 1800 10380 1970 10400
rect 2000 10500 2170 10520
rect 2000 10470 2010 10500
rect 2040 10470 2170 10500
rect 2000 10430 2170 10470
rect 2000 10400 2010 10430
rect 2040 10400 2170 10430
rect 2000 10380 2170 10400
rect 2200 10500 2370 10520
rect 2200 10470 2210 10500
rect 2240 10470 2370 10500
rect 2200 10430 2370 10470
rect 2200 10400 2210 10430
rect 2240 10400 2370 10430
rect 2200 10380 2370 10400
rect 2400 10500 2570 10520
rect 2400 10470 2410 10500
rect 2440 10470 2570 10500
rect 2400 10430 2570 10470
rect 2400 10400 2410 10430
rect 2440 10400 2570 10430
rect 2400 10380 2570 10400
rect 2600 10500 2770 10520
rect 2600 10470 2610 10500
rect 2640 10470 2770 10500
rect 2600 10430 2770 10470
rect 2600 10400 2610 10430
rect 2640 10400 2770 10430
rect 2600 10380 2770 10400
rect 2800 10500 2970 10520
rect 2800 10470 2810 10500
rect 2840 10470 2970 10500
rect 2800 10430 2970 10470
rect 2800 10400 2810 10430
rect 2840 10400 2970 10430
rect 2800 10380 2970 10400
rect 3000 10500 3170 10520
rect 3000 10470 3010 10500
rect 3040 10470 3170 10500
rect 3000 10430 3170 10470
rect 3000 10400 3010 10430
rect 3040 10400 3170 10430
rect 3000 10380 3170 10400
rect 3200 10500 3370 10520
rect 3200 10470 3210 10500
rect 3240 10470 3370 10500
rect 3200 10430 3370 10470
rect 3200 10400 3210 10430
rect 3240 10400 3370 10430
rect 3200 10380 3370 10400
rect 3400 10500 3570 10520
rect 3400 10470 3410 10500
rect 3440 10470 3570 10500
rect 3400 10430 3570 10470
rect 3400 10400 3410 10430
rect 3440 10400 3570 10430
rect 3400 10380 3570 10400
rect 3600 10500 3770 10520
rect 3600 10470 3610 10500
rect 3640 10470 3770 10500
rect 3600 10430 3770 10470
rect 3600 10400 3610 10430
rect 3640 10400 3770 10430
rect 3600 10380 3770 10400
rect 3800 10500 3970 10520
rect 3800 10470 3810 10500
rect 3840 10470 3970 10500
rect 3800 10430 3970 10470
rect 3800 10400 3810 10430
rect 3840 10400 3970 10430
rect 3800 10380 3970 10400
rect 4000 10500 4170 10520
rect 4000 10470 4010 10500
rect 4040 10470 4170 10500
rect 4000 10430 4170 10470
rect 4000 10400 4010 10430
rect 4040 10400 4170 10430
rect 4000 10380 4170 10400
rect 4200 10500 4370 10520
rect 4200 10470 4210 10500
rect 4240 10470 4370 10500
rect 4200 10430 4370 10470
rect 4200 10400 4210 10430
rect 4240 10400 4370 10430
rect 4200 10380 4370 10400
rect 4400 10500 4570 10520
rect 4400 10470 4410 10500
rect 4440 10470 4570 10500
rect 4400 10430 4570 10470
rect 4400 10400 4410 10430
rect 4440 10400 4570 10430
rect 4400 10380 4570 10400
rect 4600 10500 4770 10520
rect 4600 10470 4610 10500
rect 4640 10470 4770 10500
rect 4600 10430 4770 10470
rect 4600 10400 4610 10430
rect 4640 10400 4770 10430
rect 4600 10380 4770 10400
rect 4800 10500 4970 10520
rect 4800 10470 4810 10500
rect 4840 10470 4970 10500
rect 4800 10430 4970 10470
rect 4800 10400 4810 10430
rect 4840 10400 4970 10430
rect 4800 10380 4970 10400
rect 5000 10500 5170 10520
rect 5000 10470 5010 10500
rect 5040 10470 5170 10500
rect 5000 10430 5170 10470
rect 5000 10400 5010 10430
rect 5040 10400 5170 10430
rect 5000 10380 5170 10400
rect 5200 10500 5370 10520
rect 5200 10470 5210 10500
rect 5240 10470 5370 10500
rect 5200 10430 5370 10470
rect 5200 10400 5210 10430
rect 5240 10400 5370 10430
rect 5200 10380 5370 10400
rect 5400 10500 5570 10520
rect 5400 10470 5410 10500
rect 5440 10470 5570 10500
rect 5400 10430 5570 10470
rect 5400 10400 5410 10430
rect 5440 10400 5570 10430
rect 5400 10380 5570 10400
rect 5600 10500 5770 10520
rect 5600 10470 5610 10500
rect 5640 10470 5770 10500
rect 5600 10430 5770 10470
rect 5600 10400 5610 10430
rect 5640 10400 5770 10430
rect 5600 10380 5770 10400
rect 5800 10500 5970 10520
rect 5800 10470 5810 10500
rect 5840 10470 5970 10500
rect 5800 10430 5970 10470
rect 5800 10400 5810 10430
rect 5840 10400 5970 10430
rect 5800 10380 5970 10400
rect 6000 10500 6170 10520
rect 6000 10470 6010 10500
rect 6040 10470 6170 10500
rect 6000 10430 6170 10470
rect 6000 10400 6010 10430
rect 6040 10400 6170 10430
rect 6000 10380 6170 10400
rect 6200 10500 6370 10520
rect 6200 10470 6210 10500
rect 6240 10470 6370 10500
rect 6200 10430 6370 10470
rect 6200 10400 6210 10430
rect 6240 10400 6370 10430
rect 6200 10380 6370 10400
rect 6400 10500 6570 10520
rect 6400 10470 6410 10500
rect 6440 10470 6570 10500
rect 6400 10430 6570 10470
rect 6400 10400 6410 10430
rect 6440 10400 6570 10430
rect 6400 10380 6570 10400
rect -200 10315 -30 10335
rect -200 10285 -190 10315
rect -160 10285 -30 10315
rect -200 10245 -30 10285
rect -200 10215 -190 10245
rect -160 10215 -30 10245
rect -200 10195 -30 10215
rect 0 10315 170 10335
rect 0 10285 10 10315
rect 40 10285 170 10315
rect 0 10245 170 10285
rect 0 10215 10 10245
rect 40 10215 170 10245
rect 0 10195 170 10215
rect 200 10315 370 10335
rect 200 10285 210 10315
rect 240 10285 370 10315
rect 200 10245 370 10285
rect 200 10215 210 10245
rect 240 10215 370 10245
rect 200 10195 370 10215
rect 400 10315 570 10335
rect 400 10285 410 10315
rect 440 10285 570 10315
rect 400 10245 570 10285
rect 400 10215 410 10245
rect 440 10215 570 10245
rect 400 10195 570 10215
rect 600 10315 770 10335
rect 600 10285 610 10315
rect 640 10285 770 10315
rect 600 10245 770 10285
rect 600 10215 610 10245
rect 640 10215 770 10245
rect 600 10195 770 10215
rect 800 10315 970 10335
rect 800 10285 810 10315
rect 840 10285 970 10315
rect 800 10245 970 10285
rect 800 10215 810 10245
rect 840 10215 970 10245
rect 800 10195 970 10215
rect 1000 10315 1170 10335
rect 1000 10285 1010 10315
rect 1040 10285 1170 10315
rect 1000 10245 1170 10285
rect 1000 10215 1010 10245
rect 1040 10215 1170 10245
rect 1000 10195 1170 10215
rect 1200 10315 1370 10335
rect 1200 10285 1210 10315
rect 1240 10285 1370 10315
rect 1200 10245 1370 10285
rect 1200 10215 1210 10245
rect 1240 10215 1370 10245
rect 1200 10195 1370 10215
rect 1400 10315 1570 10335
rect 1400 10285 1410 10315
rect 1440 10285 1570 10315
rect 1400 10245 1570 10285
rect 1400 10215 1410 10245
rect 1440 10215 1570 10245
rect 1400 10195 1570 10215
rect 1600 10315 1770 10335
rect 1600 10285 1610 10315
rect 1640 10285 1770 10315
rect 1600 10245 1770 10285
rect 1600 10215 1610 10245
rect 1640 10215 1770 10245
rect 1600 10195 1770 10215
rect 1800 10315 1970 10335
rect 1800 10285 1810 10315
rect 1840 10285 1970 10315
rect 1800 10245 1970 10285
rect 1800 10215 1810 10245
rect 1840 10215 1970 10245
rect 1800 10195 1970 10215
rect 2000 10315 2170 10335
rect 2000 10285 2010 10315
rect 2040 10285 2170 10315
rect 2000 10245 2170 10285
rect 2000 10215 2010 10245
rect 2040 10215 2170 10245
rect 2000 10195 2170 10215
rect 2200 10315 2370 10335
rect 2200 10285 2210 10315
rect 2240 10285 2370 10315
rect 2200 10245 2370 10285
rect 2200 10215 2210 10245
rect 2240 10215 2370 10245
rect 2200 10195 2370 10215
rect 2400 10315 2570 10335
rect 2400 10285 2410 10315
rect 2440 10285 2570 10315
rect 2400 10245 2570 10285
rect 2400 10215 2410 10245
rect 2440 10215 2570 10245
rect 2400 10195 2570 10215
rect 2600 10315 2770 10335
rect 2600 10285 2610 10315
rect 2640 10285 2770 10315
rect 2600 10245 2770 10285
rect 2600 10215 2610 10245
rect 2640 10215 2770 10245
rect 2600 10195 2770 10215
rect 2800 10315 2970 10335
rect 2800 10285 2810 10315
rect 2840 10285 2970 10315
rect 2800 10245 2970 10285
rect 2800 10215 2810 10245
rect 2840 10215 2970 10245
rect 2800 10195 2970 10215
rect 3000 10315 3170 10335
rect 3000 10285 3010 10315
rect 3040 10285 3170 10315
rect 3000 10245 3170 10285
rect 3000 10215 3010 10245
rect 3040 10215 3170 10245
rect 3000 10195 3170 10215
rect 3200 10315 3370 10335
rect 3200 10285 3210 10315
rect 3240 10285 3370 10315
rect 3200 10245 3370 10285
rect 3200 10215 3210 10245
rect 3240 10215 3370 10245
rect 3200 10195 3370 10215
rect 3400 10315 3570 10335
rect 3400 10285 3410 10315
rect 3440 10285 3570 10315
rect 3400 10245 3570 10285
rect 3400 10215 3410 10245
rect 3440 10215 3570 10245
rect 3400 10195 3570 10215
rect 3600 10315 3770 10335
rect 3600 10285 3610 10315
rect 3640 10285 3770 10315
rect 3600 10245 3770 10285
rect 3600 10215 3610 10245
rect 3640 10215 3770 10245
rect 3600 10195 3770 10215
rect 3800 10315 3970 10335
rect 3800 10285 3810 10315
rect 3840 10285 3970 10315
rect 3800 10245 3970 10285
rect 3800 10215 3810 10245
rect 3840 10215 3970 10245
rect 3800 10195 3970 10215
rect 4000 10315 4170 10335
rect 4000 10285 4010 10315
rect 4040 10285 4170 10315
rect 4000 10245 4170 10285
rect 4000 10215 4010 10245
rect 4040 10215 4170 10245
rect 4000 10195 4170 10215
rect 4200 10315 4370 10335
rect 4200 10285 4210 10315
rect 4240 10285 4370 10315
rect 4200 10245 4370 10285
rect 4200 10215 4210 10245
rect 4240 10215 4370 10245
rect 4200 10195 4370 10215
rect 4400 10315 4570 10335
rect 4400 10285 4410 10315
rect 4440 10285 4570 10315
rect 4400 10245 4570 10285
rect 4400 10215 4410 10245
rect 4440 10215 4570 10245
rect 4400 10195 4570 10215
rect 4600 10315 4770 10335
rect 4600 10285 4610 10315
rect 4640 10285 4770 10315
rect 4600 10245 4770 10285
rect 4600 10215 4610 10245
rect 4640 10215 4770 10245
rect 4600 10195 4770 10215
rect 4800 10315 4970 10335
rect 4800 10285 4810 10315
rect 4840 10285 4970 10315
rect 4800 10245 4970 10285
rect 4800 10215 4810 10245
rect 4840 10215 4970 10245
rect 4800 10195 4970 10215
rect 5000 10315 5170 10335
rect 5000 10285 5010 10315
rect 5040 10285 5170 10315
rect 5000 10245 5170 10285
rect 5000 10215 5010 10245
rect 5040 10215 5170 10245
rect 5000 10195 5170 10215
rect 5200 10315 5370 10335
rect 5200 10285 5210 10315
rect 5240 10285 5370 10315
rect 5200 10245 5370 10285
rect 5200 10215 5210 10245
rect 5240 10215 5370 10245
rect 5200 10195 5370 10215
rect 5400 10315 5570 10335
rect 5400 10285 5410 10315
rect 5440 10285 5570 10315
rect 5400 10245 5570 10285
rect 5400 10215 5410 10245
rect 5440 10215 5570 10245
rect 5400 10195 5570 10215
rect 5600 10315 5770 10335
rect 5600 10285 5610 10315
rect 5640 10285 5770 10315
rect 5600 10245 5770 10285
rect 5600 10215 5610 10245
rect 5640 10215 5770 10245
rect 5600 10195 5770 10215
rect 5800 10315 5970 10335
rect 5800 10285 5810 10315
rect 5840 10285 5970 10315
rect 5800 10245 5970 10285
rect 5800 10215 5810 10245
rect 5840 10215 5970 10245
rect 5800 10195 5970 10215
rect 6000 10315 6170 10335
rect 6000 10285 6010 10315
rect 6040 10285 6170 10315
rect 6000 10245 6170 10285
rect 6000 10215 6010 10245
rect 6040 10215 6170 10245
rect 6000 10195 6170 10215
rect 6200 10315 6370 10335
rect 6200 10285 6210 10315
rect 6240 10285 6370 10315
rect 6200 10245 6370 10285
rect 6200 10215 6210 10245
rect 6240 10215 6370 10245
rect 6200 10195 6370 10215
rect 6400 10315 6570 10335
rect 6400 10285 6410 10315
rect 6440 10285 6570 10315
rect 6400 10245 6570 10285
rect 6400 10215 6410 10245
rect 6440 10215 6570 10245
rect 6400 10195 6570 10215
rect -200 10130 -30 10150
rect -200 10100 -190 10130
rect -160 10100 -30 10130
rect -200 10060 -30 10100
rect -200 10030 -190 10060
rect -160 10030 -30 10060
rect -200 10010 -30 10030
rect 0 10130 170 10150
rect 0 10100 10 10130
rect 40 10100 170 10130
rect 0 10060 170 10100
rect 0 10030 10 10060
rect 40 10030 170 10060
rect 0 10010 170 10030
rect 200 10130 370 10150
rect 200 10100 210 10130
rect 240 10100 370 10130
rect 200 10060 370 10100
rect 200 10030 210 10060
rect 240 10030 370 10060
rect 200 10010 370 10030
rect 400 10130 570 10150
rect 400 10100 410 10130
rect 440 10100 570 10130
rect 400 10060 570 10100
rect 400 10030 410 10060
rect 440 10030 570 10060
rect 400 10010 570 10030
rect 600 10130 770 10150
rect 600 10100 610 10130
rect 640 10100 770 10130
rect 600 10060 770 10100
rect 600 10030 610 10060
rect 640 10030 770 10060
rect 600 10010 770 10030
rect 800 10130 970 10150
rect 800 10100 810 10130
rect 840 10100 970 10130
rect 800 10060 970 10100
rect 800 10030 810 10060
rect 840 10030 970 10060
rect 800 10010 970 10030
rect 1000 10130 1170 10150
rect 1000 10100 1010 10130
rect 1040 10100 1170 10130
rect 1000 10060 1170 10100
rect 1000 10030 1010 10060
rect 1040 10030 1170 10060
rect 1000 10010 1170 10030
rect 1200 10130 1370 10150
rect 1200 10100 1210 10130
rect 1240 10100 1370 10130
rect 1200 10060 1370 10100
rect 1200 10030 1210 10060
rect 1240 10030 1370 10060
rect 1200 10010 1370 10030
rect 1400 10130 1570 10150
rect 1400 10100 1410 10130
rect 1440 10100 1570 10130
rect 1400 10060 1570 10100
rect 1400 10030 1410 10060
rect 1440 10030 1570 10060
rect 1400 10010 1570 10030
rect 1600 10130 1770 10150
rect 1600 10100 1610 10130
rect 1640 10100 1770 10130
rect 1600 10060 1770 10100
rect 1600 10030 1610 10060
rect 1640 10030 1770 10060
rect 1600 10010 1770 10030
rect 1800 10130 1970 10150
rect 1800 10100 1810 10130
rect 1840 10100 1970 10130
rect 1800 10060 1970 10100
rect 1800 10030 1810 10060
rect 1840 10030 1970 10060
rect 1800 10010 1970 10030
rect 2000 10130 2170 10150
rect 2000 10100 2010 10130
rect 2040 10100 2170 10130
rect 2000 10060 2170 10100
rect 2000 10030 2010 10060
rect 2040 10030 2170 10060
rect 2000 10010 2170 10030
rect 2200 10130 2370 10150
rect 2200 10100 2210 10130
rect 2240 10100 2370 10130
rect 2200 10060 2370 10100
rect 2200 10030 2210 10060
rect 2240 10030 2370 10060
rect 2200 10010 2370 10030
rect 2400 10130 2570 10150
rect 2400 10100 2410 10130
rect 2440 10100 2570 10130
rect 2400 10060 2570 10100
rect 2400 10030 2410 10060
rect 2440 10030 2570 10060
rect 2400 10010 2570 10030
rect 2600 10130 2770 10150
rect 2600 10100 2610 10130
rect 2640 10100 2770 10130
rect 2600 10060 2770 10100
rect 2600 10030 2610 10060
rect 2640 10030 2770 10060
rect 2600 10010 2770 10030
rect 2800 10130 2970 10150
rect 2800 10100 2810 10130
rect 2840 10100 2970 10130
rect 2800 10060 2970 10100
rect 2800 10030 2810 10060
rect 2840 10030 2970 10060
rect 2800 10010 2970 10030
rect 3000 10130 3170 10150
rect 3000 10100 3010 10130
rect 3040 10100 3170 10130
rect 3000 10060 3170 10100
rect 3000 10030 3010 10060
rect 3040 10030 3170 10060
rect 3000 10010 3170 10030
rect 3200 10130 3370 10150
rect 3200 10100 3210 10130
rect 3240 10100 3370 10130
rect 3200 10060 3370 10100
rect 3200 10030 3210 10060
rect 3240 10030 3370 10060
rect 3200 10010 3370 10030
rect 3400 10130 3570 10150
rect 3400 10100 3410 10130
rect 3440 10100 3570 10130
rect 3400 10060 3570 10100
rect 3400 10030 3410 10060
rect 3440 10030 3570 10060
rect 3400 10010 3570 10030
rect 3600 10130 3770 10150
rect 3600 10100 3610 10130
rect 3640 10100 3770 10130
rect 3600 10060 3770 10100
rect 3600 10030 3610 10060
rect 3640 10030 3770 10060
rect 3600 10010 3770 10030
rect 3800 10130 3970 10150
rect 3800 10100 3810 10130
rect 3840 10100 3970 10130
rect 3800 10060 3970 10100
rect 3800 10030 3810 10060
rect 3840 10030 3970 10060
rect 3800 10010 3970 10030
rect 4000 10130 4170 10150
rect 4000 10100 4010 10130
rect 4040 10100 4170 10130
rect 4000 10060 4170 10100
rect 4000 10030 4010 10060
rect 4040 10030 4170 10060
rect 4000 10010 4170 10030
rect 4200 10130 4370 10150
rect 4200 10100 4210 10130
rect 4240 10100 4370 10130
rect 4200 10060 4370 10100
rect 4200 10030 4210 10060
rect 4240 10030 4370 10060
rect 4200 10010 4370 10030
rect 4400 10130 4570 10150
rect 4400 10100 4410 10130
rect 4440 10100 4570 10130
rect 4400 10060 4570 10100
rect 4400 10030 4410 10060
rect 4440 10030 4570 10060
rect 4400 10010 4570 10030
rect 4600 10130 4770 10150
rect 4600 10100 4610 10130
rect 4640 10100 4770 10130
rect 4600 10060 4770 10100
rect 4600 10030 4610 10060
rect 4640 10030 4770 10060
rect 4600 10010 4770 10030
rect 4800 10130 4970 10150
rect 4800 10100 4810 10130
rect 4840 10100 4970 10130
rect 4800 10060 4970 10100
rect 4800 10030 4810 10060
rect 4840 10030 4970 10060
rect 4800 10010 4970 10030
rect 5000 10130 5170 10150
rect 5000 10100 5010 10130
rect 5040 10100 5170 10130
rect 5000 10060 5170 10100
rect 5000 10030 5010 10060
rect 5040 10030 5170 10060
rect 5000 10010 5170 10030
rect 5200 10130 5370 10150
rect 5200 10100 5210 10130
rect 5240 10100 5370 10130
rect 5200 10060 5370 10100
rect 5200 10030 5210 10060
rect 5240 10030 5370 10060
rect 5200 10010 5370 10030
rect 5400 10130 5570 10150
rect 5400 10100 5410 10130
rect 5440 10100 5570 10130
rect 5400 10060 5570 10100
rect 5400 10030 5410 10060
rect 5440 10030 5570 10060
rect 5400 10010 5570 10030
rect 5600 10130 5770 10150
rect 5600 10100 5610 10130
rect 5640 10100 5770 10130
rect 5600 10060 5770 10100
rect 5600 10030 5610 10060
rect 5640 10030 5770 10060
rect 5600 10010 5770 10030
rect 5800 10130 5970 10150
rect 5800 10100 5810 10130
rect 5840 10100 5970 10130
rect 5800 10060 5970 10100
rect 5800 10030 5810 10060
rect 5840 10030 5970 10060
rect 5800 10010 5970 10030
rect 6000 10130 6170 10150
rect 6000 10100 6010 10130
rect 6040 10100 6170 10130
rect 6000 10060 6170 10100
rect 6000 10030 6010 10060
rect 6040 10030 6170 10060
rect 6000 10010 6170 10030
rect 6200 10130 6370 10150
rect 6200 10100 6210 10130
rect 6240 10100 6370 10130
rect 6200 10060 6370 10100
rect 6200 10030 6210 10060
rect 6240 10030 6370 10060
rect 6200 10010 6370 10030
rect 6400 10130 6570 10150
rect 6400 10100 6410 10130
rect 6440 10100 6570 10130
rect 6400 10060 6570 10100
rect 6400 10030 6410 10060
rect 6440 10030 6570 10060
rect 6400 10010 6570 10030
rect -200 9945 -30 9965
rect -200 9915 -190 9945
rect -160 9915 -30 9945
rect -200 9875 -30 9915
rect -200 9845 -190 9875
rect -160 9845 -30 9875
rect -200 9825 -30 9845
rect 0 9945 170 9965
rect 0 9915 10 9945
rect 40 9915 170 9945
rect 0 9875 170 9915
rect 0 9845 10 9875
rect 40 9845 170 9875
rect 0 9825 170 9845
rect 200 9945 370 9965
rect 200 9915 210 9945
rect 240 9915 370 9945
rect 200 9875 370 9915
rect 200 9845 210 9875
rect 240 9845 370 9875
rect 200 9825 370 9845
rect 400 9945 570 9965
rect 400 9915 410 9945
rect 440 9915 570 9945
rect 400 9875 570 9915
rect 400 9845 410 9875
rect 440 9845 570 9875
rect 400 9825 570 9845
rect 600 9945 770 9965
rect 600 9915 610 9945
rect 640 9915 770 9945
rect 600 9875 770 9915
rect 600 9845 610 9875
rect 640 9845 770 9875
rect 600 9825 770 9845
rect 800 9945 970 9965
rect 800 9915 810 9945
rect 840 9915 970 9945
rect 800 9875 970 9915
rect 800 9845 810 9875
rect 840 9845 970 9875
rect 800 9825 970 9845
rect 1000 9945 1170 9965
rect 1000 9915 1010 9945
rect 1040 9915 1170 9945
rect 1000 9875 1170 9915
rect 1000 9845 1010 9875
rect 1040 9845 1170 9875
rect 1000 9825 1170 9845
rect 1200 9945 1370 9965
rect 1200 9915 1210 9945
rect 1240 9915 1370 9945
rect 1200 9875 1370 9915
rect 1200 9845 1210 9875
rect 1240 9845 1370 9875
rect 1200 9825 1370 9845
rect 1400 9945 1570 9965
rect 1400 9915 1410 9945
rect 1440 9915 1570 9945
rect 1400 9875 1570 9915
rect 1400 9845 1410 9875
rect 1440 9845 1570 9875
rect 1400 9825 1570 9845
rect 1600 9945 1770 9965
rect 1600 9915 1610 9945
rect 1640 9915 1770 9945
rect 1600 9875 1770 9915
rect 1600 9845 1610 9875
rect 1640 9845 1770 9875
rect 1600 9825 1770 9845
rect 1800 9945 1970 9965
rect 1800 9915 1810 9945
rect 1840 9915 1970 9945
rect 1800 9875 1970 9915
rect 1800 9845 1810 9875
rect 1840 9845 1970 9875
rect 1800 9825 1970 9845
rect 2000 9945 2170 9965
rect 2000 9915 2010 9945
rect 2040 9915 2170 9945
rect 2000 9875 2170 9915
rect 2000 9845 2010 9875
rect 2040 9845 2170 9875
rect 2000 9825 2170 9845
rect 2200 9945 2370 9965
rect 2200 9915 2210 9945
rect 2240 9915 2370 9945
rect 2200 9875 2370 9915
rect 2200 9845 2210 9875
rect 2240 9845 2370 9875
rect 2200 9825 2370 9845
rect 2400 9945 2570 9965
rect 2400 9915 2410 9945
rect 2440 9915 2570 9945
rect 2400 9875 2570 9915
rect 2400 9845 2410 9875
rect 2440 9845 2570 9875
rect 2400 9825 2570 9845
rect 2600 9945 2770 9965
rect 2600 9915 2610 9945
rect 2640 9915 2770 9945
rect 2600 9875 2770 9915
rect 2600 9845 2610 9875
rect 2640 9845 2770 9875
rect 2600 9825 2770 9845
rect 2800 9945 2970 9965
rect 2800 9915 2810 9945
rect 2840 9915 2970 9945
rect 2800 9875 2970 9915
rect 2800 9845 2810 9875
rect 2840 9845 2970 9875
rect 2800 9825 2970 9845
rect 3000 9945 3170 9965
rect 3000 9915 3010 9945
rect 3040 9915 3170 9945
rect 3000 9875 3170 9915
rect 3000 9845 3010 9875
rect 3040 9845 3170 9875
rect 3000 9825 3170 9845
rect 3200 9945 3370 9965
rect 3200 9915 3210 9945
rect 3240 9915 3370 9945
rect 3200 9875 3370 9915
rect 3200 9845 3210 9875
rect 3240 9845 3370 9875
rect 3200 9825 3370 9845
rect 3400 9945 3570 9965
rect 3400 9915 3410 9945
rect 3440 9915 3570 9945
rect 3400 9875 3570 9915
rect 3400 9845 3410 9875
rect 3440 9845 3570 9875
rect 3400 9825 3570 9845
rect 3600 9945 3770 9965
rect 3600 9915 3610 9945
rect 3640 9915 3770 9945
rect 3600 9875 3770 9915
rect 3600 9845 3610 9875
rect 3640 9845 3770 9875
rect 3600 9825 3770 9845
rect 3800 9945 3970 9965
rect 3800 9915 3810 9945
rect 3840 9915 3970 9945
rect 3800 9875 3970 9915
rect 3800 9845 3810 9875
rect 3840 9845 3970 9875
rect 3800 9825 3970 9845
rect 4000 9945 4170 9965
rect 4000 9915 4010 9945
rect 4040 9915 4170 9945
rect 4000 9875 4170 9915
rect 4000 9845 4010 9875
rect 4040 9845 4170 9875
rect 4000 9825 4170 9845
rect 4200 9945 4370 9965
rect 4200 9915 4210 9945
rect 4240 9915 4370 9945
rect 4200 9875 4370 9915
rect 4200 9845 4210 9875
rect 4240 9845 4370 9875
rect 4200 9825 4370 9845
rect 4400 9945 4570 9965
rect 4400 9915 4410 9945
rect 4440 9915 4570 9945
rect 4400 9875 4570 9915
rect 4400 9845 4410 9875
rect 4440 9845 4570 9875
rect 4400 9825 4570 9845
rect 4600 9945 4770 9965
rect 4600 9915 4610 9945
rect 4640 9915 4770 9945
rect 4600 9875 4770 9915
rect 4600 9845 4610 9875
rect 4640 9845 4770 9875
rect 4600 9825 4770 9845
rect 4800 9945 4970 9965
rect 4800 9915 4810 9945
rect 4840 9915 4970 9945
rect 4800 9875 4970 9915
rect 4800 9845 4810 9875
rect 4840 9845 4970 9875
rect 4800 9825 4970 9845
rect 5000 9945 5170 9965
rect 5000 9915 5010 9945
rect 5040 9915 5170 9945
rect 5000 9875 5170 9915
rect 5000 9845 5010 9875
rect 5040 9845 5170 9875
rect 5000 9825 5170 9845
rect 5200 9945 5370 9965
rect 5200 9915 5210 9945
rect 5240 9915 5370 9945
rect 5200 9875 5370 9915
rect 5200 9845 5210 9875
rect 5240 9845 5370 9875
rect 5200 9825 5370 9845
rect 5400 9945 5570 9965
rect 5400 9915 5410 9945
rect 5440 9915 5570 9945
rect 5400 9875 5570 9915
rect 5400 9845 5410 9875
rect 5440 9845 5570 9875
rect 5400 9825 5570 9845
rect 5600 9945 5770 9965
rect 5600 9915 5610 9945
rect 5640 9915 5770 9945
rect 5600 9875 5770 9915
rect 5600 9845 5610 9875
rect 5640 9845 5770 9875
rect 5600 9825 5770 9845
rect 5800 9945 5970 9965
rect 5800 9915 5810 9945
rect 5840 9915 5970 9945
rect 5800 9875 5970 9915
rect 5800 9845 5810 9875
rect 5840 9845 5970 9875
rect 5800 9825 5970 9845
rect 6000 9945 6170 9965
rect 6000 9915 6010 9945
rect 6040 9915 6170 9945
rect 6000 9875 6170 9915
rect 6000 9845 6010 9875
rect 6040 9845 6170 9875
rect 6000 9825 6170 9845
rect 6200 9945 6370 9965
rect 6200 9915 6210 9945
rect 6240 9915 6370 9945
rect 6200 9875 6370 9915
rect 6200 9845 6210 9875
rect 6240 9845 6370 9875
rect 6200 9825 6370 9845
rect 6400 9945 6570 9965
rect 6400 9915 6410 9945
rect 6440 9915 6570 9945
rect 6400 9875 6570 9915
rect 6400 9845 6410 9875
rect 6440 9845 6570 9875
rect 6400 9825 6570 9845
rect -200 9760 -30 9780
rect -200 9730 -190 9760
rect -160 9730 -30 9760
rect -200 9690 -30 9730
rect -200 9660 -190 9690
rect -160 9660 -30 9690
rect -200 9640 -30 9660
rect 0 9760 170 9780
rect 0 9730 10 9760
rect 40 9730 170 9760
rect 0 9690 170 9730
rect 0 9660 10 9690
rect 40 9660 170 9690
rect 0 9640 170 9660
rect 200 9760 370 9780
rect 200 9730 210 9760
rect 240 9730 370 9760
rect 200 9690 370 9730
rect 200 9660 210 9690
rect 240 9660 370 9690
rect 200 9640 370 9660
rect 400 9760 570 9780
rect 400 9730 410 9760
rect 440 9730 570 9760
rect 400 9690 570 9730
rect 400 9660 410 9690
rect 440 9660 570 9690
rect 400 9640 570 9660
rect 600 9760 770 9780
rect 600 9730 610 9760
rect 640 9730 770 9760
rect 600 9690 770 9730
rect 600 9660 610 9690
rect 640 9660 770 9690
rect 600 9640 770 9660
rect 800 9760 970 9780
rect 800 9730 810 9760
rect 840 9730 970 9760
rect 800 9690 970 9730
rect 800 9660 810 9690
rect 840 9660 970 9690
rect 800 9640 970 9660
rect 1000 9760 1170 9780
rect 1000 9730 1010 9760
rect 1040 9730 1170 9760
rect 1000 9690 1170 9730
rect 1000 9660 1010 9690
rect 1040 9660 1170 9690
rect 1000 9640 1170 9660
rect 1200 9760 1370 9780
rect 1200 9730 1210 9760
rect 1240 9730 1370 9760
rect 1200 9690 1370 9730
rect 1200 9660 1210 9690
rect 1240 9660 1370 9690
rect 1200 9640 1370 9660
rect 1400 9760 1570 9780
rect 1400 9730 1410 9760
rect 1440 9730 1570 9760
rect 1400 9690 1570 9730
rect 1400 9660 1410 9690
rect 1440 9660 1570 9690
rect 1400 9640 1570 9660
rect 1600 9760 1770 9780
rect 1600 9730 1610 9760
rect 1640 9730 1770 9760
rect 1600 9690 1770 9730
rect 1600 9660 1610 9690
rect 1640 9660 1770 9690
rect 1600 9640 1770 9660
rect 1800 9760 1970 9780
rect 1800 9730 1810 9760
rect 1840 9730 1970 9760
rect 1800 9690 1970 9730
rect 1800 9660 1810 9690
rect 1840 9660 1970 9690
rect 1800 9640 1970 9660
rect 2000 9760 2170 9780
rect 2000 9730 2010 9760
rect 2040 9730 2170 9760
rect 2000 9690 2170 9730
rect 2000 9660 2010 9690
rect 2040 9660 2170 9690
rect 2000 9640 2170 9660
rect 2200 9760 2370 9780
rect 2200 9730 2210 9760
rect 2240 9730 2370 9760
rect 2200 9690 2370 9730
rect 2200 9660 2210 9690
rect 2240 9660 2370 9690
rect 2200 9640 2370 9660
rect 2400 9760 2570 9780
rect 2400 9730 2410 9760
rect 2440 9730 2570 9760
rect 2400 9690 2570 9730
rect 2400 9660 2410 9690
rect 2440 9660 2570 9690
rect 2400 9640 2570 9660
rect 2600 9760 2770 9780
rect 2600 9730 2610 9760
rect 2640 9730 2770 9760
rect 2600 9690 2770 9730
rect 2600 9660 2610 9690
rect 2640 9660 2770 9690
rect 2600 9640 2770 9660
rect 2800 9760 2970 9780
rect 2800 9730 2810 9760
rect 2840 9730 2970 9760
rect 2800 9690 2970 9730
rect 2800 9660 2810 9690
rect 2840 9660 2970 9690
rect 2800 9640 2970 9660
rect 3000 9760 3170 9780
rect 3000 9730 3010 9760
rect 3040 9730 3170 9760
rect 3000 9690 3170 9730
rect 3000 9660 3010 9690
rect 3040 9660 3170 9690
rect 3000 9640 3170 9660
rect 3200 9760 3370 9780
rect 3200 9730 3210 9760
rect 3240 9730 3370 9760
rect 3200 9690 3370 9730
rect 3200 9660 3210 9690
rect 3240 9660 3370 9690
rect 3200 9640 3370 9660
rect 3400 9760 3570 9780
rect 3400 9730 3410 9760
rect 3440 9730 3570 9760
rect 3400 9690 3570 9730
rect 3400 9660 3410 9690
rect 3440 9660 3570 9690
rect 3400 9640 3570 9660
rect 3600 9760 3770 9780
rect 3600 9730 3610 9760
rect 3640 9730 3770 9760
rect 3600 9690 3770 9730
rect 3600 9660 3610 9690
rect 3640 9660 3770 9690
rect 3600 9640 3770 9660
rect 3800 9760 3970 9780
rect 3800 9730 3810 9760
rect 3840 9730 3970 9760
rect 3800 9690 3970 9730
rect 3800 9660 3810 9690
rect 3840 9660 3970 9690
rect 3800 9640 3970 9660
rect 4000 9760 4170 9780
rect 4000 9730 4010 9760
rect 4040 9730 4170 9760
rect 4000 9690 4170 9730
rect 4000 9660 4010 9690
rect 4040 9660 4170 9690
rect 4000 9640 4170 9660
rect 4200 9760 4370 9780
rect 4200 9730 4210 9760
rect 4240 9730 4370 9760
rect 4200 9690 4370 9730
rect 4200 9660 4210 9690
rect 4240 9660 4370 9690
rect 4200 9640 4370 9660
rect 4400 9760 4570 9780
rect 4400 9730 4410 9760
rect 4440 9730 4570 9760
rect 4400 9690 4570 9730
rect 4400 9660 4410 9690
rect 4440 9660 4570 9690
rect 4400 9640 4570 9660
rect 4600 9760 4770 9780
rect 4600 9730 4610 9760
rect 4640 9730 4770 9760
rect 4600 9690 4770 9730
rect 4600 9660 4610 9690
rect 4640 9660 4770 9690
rect 4600 9640 4770 9660
rect 4800 9760 4970 9780
rect 4800 9730 4810 9760
rect 4840 9730 4970 9760
rect 4800 9690 4970 9730
rect 4800 9660 4810 9690
rect 4840 9660 4970 9690
rect 4800 9640 4970 9660
rect 5000 9760 5170 9780
rect 5000 9730 5010 9760
rect 5040 9730 5170 9760
rect 5000 9690 5170 9730
rect 5000 9660 5010 9690
rect 5040 9660 5170 9690
rect 5000 9640 5170 9660
rect 5200 9760 5370 9780
rect 5200 9730 5210 9760
rect 5240 9730 5370 9760
rect 5200 9690 5370 9730
rect 5200 9660 5210 9690
rect 5240 9660 5370 9690
rect 5200 9640 5370 9660
rect 5400 9760 5570 9780
rect 5400 9730 5410 9760
rect 5440 9730 5570 9760
rect 5400 9690 5570 9730
rect 5400 9660 5410 9690
rect 5440 9660 5570 9690
rect 5400 9640 5570 9660
rect 5600 9760 5770 9780
rect 5600 9730 5610 9760
rect 5640 9730 5770 9760
rect 5600 9690 5770 9730
rect 5600 9660 5610 9690
rect 5640 9660 5770 9690
rect 5600 9640 5770 9660
rect 5800 9760 5970 9780
rect 5800 9730 5810 9760
rect 5840 9730 5970 9760
rect 5800 9690 5970 9730
rect 5800 9660 5810 9690
rect 5840 9660 5970 9690
rect 5800 9640 5970 9660
rect 6000 9760 6170 9780
rect 6000 9730 6010 9760
rect 6040 9730 6170 9760
rect 6000 9690 6170 9730
rect 6000 9660 6010 9690
rect 6040 9660 6170 9690
rect 6000 9640 6170 9660
rect 6200 9760 6370 9780
rect 6200 9730 6210 9760
rect 6240 9730 6370 9760
rect 6200 9690 6370 9730
rect 6200 9660 6210 9690
rect 6240 9660 6370 9690
rect 6200 9640 6370 9660
rect 6400 9760 6570 9780
rect 6400 9730 6410 9760
rect 6440 9730 6570 9760
rect 6400 9690 6570 9730
rect 6400 9660 6410 9690
rect 6440 9660 6570 9690
rect 6400 9640 6570 9660
rect -200 9575 -30 9595
rect -200 9545 -190 9575
rect -160 9545 -30 9575
rect -200 9505 -30 9545
rect -200 9475 -190 9505
rect -160 9475 -30 9505
rect -200 9455 -30 9475
rect 0 9575 170 9595
rect 0 9545 10 9575
rect 40 9545 170 9575
rect 0 9505 170 9545
rect 0 9475 10 9505
rect 40 9475 170 9505
rect 0 9455 170 9475
rect 200 9575 370 9595
rect 200 9545 210 9575
rect 240 9545 370 9575
rect 200 9505 370 9545
rect 200 9475 210 9505
rect 240 9475 370 9505
rect 200 9455 370 9475
rect 400 9575 570 9595
rect 400 9545 410 9575
rect 440 9545 570 9575
rect 400 9505 570 9545
rect 400 9475 410 9505
rect 440 9475 570 9505
rect 400 9455 570 9475
rect 600 9575 770 9595
rect 600 9545 610 9575
rect 640 9545 770 9575
rect 600 9505 770 9545
rect 600 9475 610 9505
rect 640 9475 770 9505
rect 600 9455 770 9475
rect 800 9575 970 9595
rect 800 9545 810 9575
rect 840 9545 970 9575
rect 800 9505 970 9545
rect 800 9475 810 9505
rect 840 9475 970 9505
rect 800 9455 970 9475
rect 1000 9575 1170 9595
rect 1000 9545 1010 9575
rect 1040 9545 1170 9575
rect 1000 9505 1170 9545
rect 1000 9475 1010 9505
rect 1040 9475 1170 9505
rect 1000 9455 1170 9475
rect 1200 9575 1370 9595
rect 1200 9545 1210 9575
rect 1240 9545 1370 9575
rect 1200 9505 1370 9545
rect 1200 9475 1210 9505
rect 1240 9475 1370 9505
rect 1200 9455 1370 9475
rect 1400 9575 1570 9595
rect 1400 9545 1410 9575
rect 1440 9545 1570 9575
rect 1400 9505 1570 9545
rect 1400 9475 1410 9505
rect 1440 9475 1570 9505
rect 1400 9455 1570 9475
rect 1600 9575 1770 9595
rect 1600 9545 1610 9575
rect 1640 9545 1770 9575
rect 1600 9505 1770 9545
rect 1600 9475 1610 9505
rect 1640 9475 1770 9505
rect 1600 9455 1770 9475
rect 1800 9575 1970 9595
rect 1800 9545 1810 9575
rect 1840 9545 1970 9575
rect 1800 9505 1970 9545
rect 1800 9475 1810 9505
rect 1840 9475 1970 9505
rect 1800 9455 1970 9475
rect 2000 9575 2170 9595
rect 2000 9545 2010 9575
rect 2040 9545 2170 9575
rect 2000 9505 2170 9545
rect 2000 9475 2010 9505
rect 2040 9475 2170 9505
rect 2000 9455 2170 9475
rect 2200 9575 2370 9595
rect 2200 9545 2210 9575
rect 2240 9545 2370 9575
rect 2200 9505 2370 9545
rect 2200 9475 2210 9505
rect 2240 9475 2370 9505
rect 2200 9455 2370 9475
rect 2400 9575 2570 9595
rect 2400 9545 2410 9575
rect 2440 9545 2570 9575
rect 2400 9505 2570 9545
rect 2400 9475 2410 9505
rect 2440 9475 2570 9505
rect 2400 9455 2570 9475
rect 2600 9575 2770 9595
rect 2600 9545 2610 9575
rect 2640 9545 2770 9575
rect 2600 9505 2770 9545
rect 2600 9475 2610 9505
rect 2640 9475 2770 9505
rect 2600 9455 2770 9475
rect 2800 9575 2970 9595
rect 2800 9545 2810 9575
rect 2840 9545 2970 9575
rect 2800 9505 2970 9545
rect 2800 9475 2810 9505
rect 2840 9475 2970 9505
rect 2800 9455 2970 9475
rect 3000 9575 3170 9595
rect 3000 9545 3010 9575
rect 3040 9545 3170 9575
rect 3000 9505 3170 9545
rect 3000 9475 3010 9505
rect 3040 9475 3170 9505
rect 3000 9455 3170 9475
rect 3200 9575 3370 9595
rect 3200 9545 3210 9575
rect 3240 9545 3370 9575
rect 3200 9505 3370 9545
rect 3200 9475 3210 9505
rect 3240 9475 3370 9505
rect 3200 9455 3370 9475
rect 3400 9575 3570 9595
rect 3400 9545 3410 9575
rect 3440 9545 3570 9575
rect 3400 9505 3570 9545
rect 3400 9475 3410 9505
rect 3440 9475 3570 9505
rect 3400 9455 3570 9475
rect 3600 9575 3770 9595
rect 3600 9545 3610 9575
rect 3640 9545 3770 9575
rect 3600 9505 3770 9545
rect 3600 9475 3610 9505
rect 3640 9475 3770 9505
rect 3600 9455 3770 9475
rect 3800 9575 3970 9595
rect 3800 9545 3810 9575
rect 3840 9545 3970 9575
rect 3800 9505 3970 9545
rect 3800 9475 3810 9505
rect 3840 9475 3970 9505
rect 3800 9455 3970 9475
rect 4000 9575 4170 9595
rect 4000 9545 4010 9575
rect 4040 9545 4170 9575
rect 4000 9505 4170 9545
rect 4000 9475 4010 9505
rect 4040 9475 4170 9505
rect 4000 9455 4170 9475
rect 4200 9575 4370 9595
rect 4200 9545 4210 9575
rect 4240 9545 4370 9575
rect 4200 9505 4370 9545
rect 4200 9475 4210 9505
rect 4240 9475 4370 9505
rect 4200 9455 4370 9475
rect 4400 9575 4570 9595
rect 4400 9545 4410 9575
rect 4440 9545 4570 9575
rect 4400 9505 4570 9545
rect 4400 9475 4410 9505
rect 4440 9475 4570 9505
rect 4400 9455 4570 9475
rect 4600 9575 4770 9595
rect 4600 9545 4610 9575
rect 4640 9545 4770 9575
rect 4600 9505 4770 9545
rect 4600 9475 4610 9505
rect 4640 9475 4770 9505
rect 4600 9455 4770 9475
rect 4800 9575 4970 9595
rect 4800 9545 4810 9575
rect 4840 9545 4970 9575
rect 4800 9505 4970 9545
rect 4800 9475 4810 9505
rect 4840 9475 4970 9505
rect 4800 9455 4970 9475
rect 5000 9575 5170 9595
rect 5000 9545 5010 9575
rect 5040 9545 5170 9575
rect 5000 9505 5170 9545
rect 5000 9475 5010 9505
rect 5040 9475 5170 9505
rect 5000 9455 5170 9475
rect 5200 9575 5370 9595
rect 5200 9545 5210 9575
rect 5240 9545 5370 9575
rect 5200 9505 5370 9545
rect 5200 9475 5210 9505
rect 5240 9475 5370 9505
rect 5200 9455 5370 9475
rect 5400 9575 5570 9595
rect 5400 9545 5410 9575
rect 5440 9545 5570 9575
rect 5400 9505 5570 9545
rect 5400 9475 5410 9505
rect 5440 9475 5570 9505
rect 5400 9455 5570 9475
rect 5600 9575 5770 9595
rect 5600 9545 5610 9575
rect 5640 9545 5770 9575
rect 5600 9505 5770 9545
rect 5600 9475 5610 9505
rect 5640 9475 5770 9505
rect 5600 9455 5770 9475
rect 5800 9575 5970 9595
rect 5800 9545 5810 9575
rect 5840 9545 5970 9575
rect 5800 9505 5970 9545
rect 5800 9475 5810 9505
rect 5840 9475 5970 9505
rect 5800 9455 5970 9475
rect 6000 9575 6170 9595
rect 6000 9545 6010 9575
rect 6040 9545 6170 9575
rect 6000 9505 6170 9545
rect 6000 9475 6010 9505
rect 6040 9475 6170 9505
rect 6000 9455 6170 9475
rect 6200 9575 6370 9595
rect 6200 9545 6210 9575
rect 6240 9545 6370 9575
rect 6200 9505 6370 9545
rect 6200 9475 6210 9505
rect 6240 9475 6370 9505
rect 6200 9455 6370 9475
rect 6400 9575 6570 9595
rect 6400 9545 6410 9575
rect 6440 9545 6570 9575
rect 6400 9505 6570 9545
rect 6400 9475 6410 9505
rect 6440 9475 6570 9505
rect 6400 9455 6570 9475
rect -200 9390 -30 9410
rect -200 9360 -190 9390
rect -160 9360 -30 9390
rect -200 9320 -30 9360
rect -200 9290 -190 9320
rect -160 9290 -30 9320
rect -200 9270 -30 9290
rect 0 9390 170 9410
rect 0 9360 10 9390
rect 40 9360 170 9390
rect 0 9320 170 9360
rect 0 9290 10 9320
rect 40 9290 170 9320
rect 0 9270 170 9290
rect 200 9390 370 9410
rect 200 9360 210 9390
rect 240 9360 370 9390
rect 200 9320 370 9360
rect 200 9290 210 9320
rect 240 9290 370 9320
rect 200 9270 370 9290
rect 400 9390 570 9410
rect 400 9360 410 9390
rect 440 9360 570 9390
rect 400 9320 570 9360
rect 400 9290 410 9320
rect 440 9290 570 9320
rect 400 9270 570 9290
rect 600 9390 770 9410
rect 600 9360 610 9390
rect 640 9360 770 9390
rect 600 9320 770 9360
rect 600 9290 610 9320
rect 640 9290 770 9320
rect 600 9270 770 9290
rect 800 9390 970 9410
rect 800 9360 810 9390
rect 840 9360 970 9390
rect 800 9320 970 9360
rect 800 9290 810 9320
rect 840 9290 970 9320
rect 800 9270 970 9290
rect 1000 9390 1170 9410
rect 1000 9360 1010 9390
rect 1040 9360 1170 9390
rect 1000 9320 1170 9360
rect 1000 9290 1010 9320
rect 1040 9290 1170 9320
rect 1000 9270 1170 9290
rect 1200 9390 1370 9410
rect 1200 9360 1210 9390
rect 1240 9360 1370 9390
rect 1200 9320 1370 9360
rect 1200 9290 1210 9320
rect 1240 9290 1370 9320
rect 1200 9270 1370 9290
rect 1400 9390 1570 9410
rect 1400 9360 1410 9390
rect 1440 9360 1570 9390
rect 1400 9320 1570 9360
rect 1400 9290 1410 9320
rect 1440 9290 1570 9320
rect 1400 9270 1570 9290
rect 1600 9390 1770 9410
rect 1600 9360 1610 9390
rect 1640 9360 1770 9390
rect 1600 9320 1770 9360
rect 1600 9290 1610 9320
rect 1640 9290 1770 9320
rect 1600 9270 1770 9290
rect 1800 9390 1970 9410
rect 1800 9360 1810 9390
rect 1840 9360 1970 9390
rect 1800 9320 1970 9360
rect 1800 9290 1810 9320
rect 1840 9290 1970 9320
rect 1800 9270 1970 9290
rect 2000 9390 2170 9410
rect 2000 9360 2010 9390
rect 2040 9360 2170 9390
rect 2000 9320 2170 9360
rect 2000 9290 2010 9320
rect 2040 9290 2170 9320
rect 2000 9270 2170 9290
rect 2200 9390 2370 9410
rect 2200 9360 2210 9390
rect 2240 9360 2370 9390
rect 2200 9320 2370 9360
rect 2200 9290 2210 9320
rect 2240 9290 2370 9320
rect 2200 9270 2370 9290
rect 2400 9390 2570 9410
rect 2400 9360 2410 9390
rect 2440 9360 2570 9390
rect 2400 9320 2570 9360
rect 2400 9290 2410 9320
rect 2440 9290 2570 9320
rect 2400 9270 2570 9290
rect 2600 9390 2770 9410
rect 2600 9360 2610 9390
rect 2640 9360 2770 9390
rect 2600 9320 2770 9360
rect 2600 9290 2610 9320
rect 2640 9290 2770 9320
rect 2600 9270 2770 9290
rect 2800 9390 2970 9410
rect 2800 9360 2810 9390
rect 2840 9360 2970 9390
rect 2800 9320 2970 9360
rect 2800 9290 2810 9320
rect 2840 9290 2970 9320
rect 2800 9270 2970 9290
rect 3000 9390 3170 9410
rect 3000 9360 3010 9390
rect 3040 9360 3170 9390
rect 3000 9320 3170 9360
rect 3000 9290 3010 9320
rect 3040 9290 3170 9320
rect 3000 9270 3170 9290
rect 3200 9390 3370 9410
rect 3200 9360 3210 9390
rect 3240 9360 3370 9390
rect 3200 9320 3370 9360
rect 3200 9290 3210 9320
rect 3240 9290 3370 9320
rect 3200 9270 3370 9290
rect 3400 9390 3570 9410
rect 3400 9360 3410 9390
rect 3440 9360 3570 9390
rect 3400 9320 3570 9360
rect 3400 9290 3410 9320
rect 3440 9290 3570 9320
rect 3400 9270 3570 9290
rect 3600 9390 3770 9410
rect 3600 9360 3610 9390
rect 3640 9360 3770 9390
rect 3600 9320 3770 9360
rect 3600 9290 3610 9320
rect 3640 9290 3770 9320
rect 3600 9270 3770 9290
rect 3800 9390 3970 9410
rect 3800 9360 3810 9390
rect 3840 9360 3970 9390
rect 3800 9320 3970 9360
rect 3800 9290 3810 9320
rect 3840 9290 3970 9320
rect 3800 9270 3970 9290
rect 4000 9390 4170 9410
rect 4000 9360 4010 9390
rect 4040 9360 4170 9390
rect 4000 9320 4170 9360
rect 4000 9290 4010 9320
rect 4040 9290 4170 9320
rect 4000 9270 4170 9290
rect 4200 9390 4370 9410
rect 4200 9360 4210 9390
rect 4240 9360 4370 9390
rect 4200 9320 4370 9360
rect 4200 9290 4210 9320
rect 4240 9290 4370 9320
rect 4200 9270 4370 9290
rect 4400 9390 4570 9410
rect 4400 9360 4410 9390
rect 4440 9360 4570 9390
rect 4400 9320 4570 9360
rect 4400 9290 4410 9320
rect 4440 9290 4570 9320
rect 4400 9270 4570 9290
rect 4600 9390 4770 9410
rect 4600 9360 4610 9390
rect 4640 9360 4770 9390
rect 4600 9320 4770 9360
rect 4600 9290 4610 9320
rect 4640 9290 4770 9320
rect 4600 9270 4770 9290
rect 4800 9390 4970 9410
rect 4800 9360 4810 9390
rect 4840 9360 4970 9390
rect 4800 9320 4970 9360
rect 4800 9290 4810 9320
rect 4840 9290 4970 9320
rect 4800 9270 4970 9290
rect 5000 9390 5170 9410
rect 5000 9360 5010 9390
rect 5040 9360 5170 9390
rect 5000 9320 5170 9360
rect 5000 9290 5010 9320
rect 5040 9290 5170 9320
rect 5000 9270 5170 9290
rect 5200 9390 5370 9410
rect 5200 9360 5210 9390
rect 5240 9360 5370 9390
rect 5200 9320 5370 9360
rect 5200 9290 5210 9320
rect 5240 9290 5370 9320
rect 5200 9270 5370 9290
rect 5400 9390 5570 9410
rect 5400 9360 5410 9390
rect 5440 9360 5570 9390
rect 5400 9320 5570 9360
rect 5400 9290 5410 9320
rect 5440 9290 5570 9320
rect 5400 9270 5570 9290
rect 5600 9390 5770 9410
rect 5600 9360 5610 9390
rect 5640 9360 5770 9390
rect 5600 9320 5770 9360
rect 5600 9290 5610 9320
rect 5640 9290 5770 9320
rect 5600 9270 5770 9290
rect 5800 9390 5970 9410
rect 5800 9360 5810 9390
rect 5840 9360 5970 9390
rect 5800 9320 5970 9360
rect 5800 9290 5810 9320
rect 5840 9290 5970 9320
rect 5800 9270 5970 9290
rect 6000 9390 6170 9410
rect 6000 9360 6010 9390
rect 6040 9360 6170 9390
rect 6000 9320 6170 9360
rect 6000 9290 6010 9320
rect 6040 9290 6170 9320
rect 6000 9270 6170 9290
rect 6200 9390 6370 9410
rect 6200 9360 6210 9390
rect 6240 9360 6370 9390
rect 6200 9320 6370 9360
rect 6200 9290 6210 9320
rect 6240 9290 6370 9320
rect 6200 9270 6370 9290
rect 6400 9390 6570 9410
rect 6400 9360 6410 9390
rect 6440 9360 6570 9390
rect 6400 9320 6570 9360
rect 6400 9290 6410 9320
rect 6440 9290 6570 9320
rect 6400 9270 6570 9290
rect -200 9205 -30 9225
rect -200 9175 -190 9205
rect -160 9175 -30 9205
rect -200 9135 -30 9175
rect -200 9105 -190 9135
rect -160 9105 -30 9135
rect -200 9085 -30 9105
rect 0 9205 170 9225
rect 0 9175 10 9205
rect 40 9175 170 9205
rect 0 9135 170 9175
rect 0 9105 10 9135
rect 40 9105 170 9135
rect 0 9085 170 9105
rect 200 9205 370 9225
rect 200 9175 210 9205
rect 240 9175 370 9205
rect 200 9135 370 9175
rect 200 9105 210 9135
rect 240 9105 370 9135
rect 200 9085 370 9105
rect 400 9205 570 9225
rect 400 9175 410 9205
rect 440 9175 570 9205
rect 400 9135 570 9175
rect 400 9105 410 9135
rect 440 9105 570 9135
rect 400 9085 570 9105
rect 600 9205 770 9225
rect 600 9175 610 9205
rect 640 9175 770 9205
rect 600 9135 770 9175
rect 600 9105 610 9135
rect 640 9105 770 9135
rect 600 9085 770 9105
rect 800 9205 970 9225
rect 800 9175 810 9205
rect 840 9175 970 9205
rect 800 9135 970 9175
rect 800 9105 810 9135
rect 840 9105 970 9135
rect 800 9085 970 9105
rect 1000 9205 1170 9225
rect 1000 9175 1010 9205
rect 1040 9175 1170 9205
rect 1000 9135 1170 9175
rect 1000 9105 1010 9135
rect 1040 9105 1170 9135
rect 1000 9085 1170 9105
rect 1200 9205 1370 9225
rect 1200 9175 1210 9205
rect 1240 9175 1370 9205
rect 1200 9135 1370 9175
rect 1200 9105 1210 9135
rect 1240 9105 1370 9135
rect 1200 9085 1370 9105
rect 1400 9205 1570 9225
rect 1400 9175 1410 9205
rect 1440 9175 1570 9205
rect 1400 9135 1570 9175
rect 1400 9105 1410 9135
rect 1440 9105 1570 9135
rect 1400 9085 1570 9105
rect 1600 9205 1770 9225
rect 1600 9175 1610 9205
rect 1640 9175 1770 9205
rect 1600 9135 1770 9175
rect 1600 9105 1610 9135
rect 1640 9105 1770 9135
rect 1600 9085 1770 9105
rect 1800 9205 1970 9225
rect 1800 9175 1810 9205
rect 1840 9175 1970 9205
rect 1800 9135 1970 9175
rect 1800 9105 1810 9135
rect 1840 9105 1970 9135
rect 1800 9085 1970 9105
rect 2000 9205 2170 9225
rect 2000 9175 2010 9205
rect 2040 9175 2170 9205
rect 2000 9135 2170 9175
rect 2000 9105 2010 9135
rect 2040 9105 2170 9135
rect 2000 9085 2170 9105
rect 2200 9205 2370 9225
rect 2200 9175 2210 9205
rect 2240 9175 2370 9205
rect 2200 9135 2370 9175
rect 2200 9105 2210 9135
rect 2240 9105 2370 9135
rect 2200 9085 2370 9105
rect 2400 9205 2570 9225
rect 2400 9175 2410 9205
rect 2440 9175 2570 9205
rect 2400 9135 2570 9175
rect 2400 9105 2410 9135
rect 2440 9105 2570 9135
rect 2400 9085 2570 9105
rect 2600 9205 2770 9225
rect 2600 9175 2610 9205
rect 2640 9175 2770 9205
rect 2600 9135 2770 9175
rect 2600 9105 2610 9135
rect 2640 9105 2770 9135
rect 2600 9085 2770 9105
rect 2800 9205 2970 9225
rect 2800 9175 2810 9205
rect 2840 9175 2970 9205
rect 2800 9135 2970 9175
rect 2800 9105 2810 9135
rect 2840 9105 2970 9135
rect 2800 9085 2970 9105
rect 3000 9205 3170 9225
rect 3000 9175 3010 9205
rect 3040 9175 3170 9205
rect 3000 9135 3170 9175
rect 3000 9105 3010 9135
rect 3040 9105 3170 9135
rect 3000 9085 3170 9105
rect 3200 9205 3370 9225
rect 3200 9175 3210 9205
rect 3240 9175 3370 9205
rect 3200 9135 3370 9175
rect 3200 9105 3210 9135
rect 3240 9105 3370 9135
rect 3200 9085 3370 9105
rect 3400 9205 3570 9225
rect 3400 9175 3410 9205
rect 3440 9175 3570 9205
rect 3400 9135 3570 9175
rect 3400 9105 3410 9135
rect 3440 9105 3570 9135
rect 3400 9085 3570 9105
rect 3600 9205 3770 9225
rect 3600 9175 3610 9205
rect 3640 9175 3770 9205
rect 3600 9135 3770 9175
rect 3600 9105 3610 9135
rect 3640 9105 3770 9135
rect 3600 9085 3770 9105
rect 3800 9205 3970 9225
rect 3800 9175 3810 9205
rect 3840 9175 3970 9205
rect 3800 9135 3970 9175
rect 3800 9105 3810 9135
rect 3840 9105 3970 9135
rect 3800 9085 3970 9105
rect 4000 9205 4170 9225
rect 4000 9175 4010 9205
rect 4040 9175 4170 9205
rect 4000 9135 4170 9175
rect 4000 9105 4010 9135
rect 4040 9105 4170 9135
rect 4000 9085 4170 9105
rect 4200 9205 4370 9225
rect 4200 9175 4210 9205
rect 4240 9175 4370 9205
rect 4200 9135 4370 9175
rect 4200 9105 4210 9135
rect 4240 9105 4370 9135
rect 4200 9085 4370 9105
rect 4400 9205 4570 9225
rect 4400 9175 4410 9205
rect 4440 9175 4570 9205
rect 4400 9135 4570 9175
rect 4400 9105 4410 9135
rect 4440 9105 4570 9135
rect 4400 9085 4570 9105
rect 4600 9205 4770 9225
rect 4600 9175 4610 9205
rect 4640 9175 4770 9205
rect 4600 9135 4770 9175
rect 4600 9105 4610 9135
rect 4640 9105 4770 9135
rect 4600 9085 4770 9105
rect 4800 9205 4970 9225
rect 4800 9175 4810 9205
rect 4840 9175 4970 9205
rect 4800 9135 4970 9175
rect 4800 9105 4810 9135
rect 4840 9105 4970 9135
rect 4800 9085 4970 9105
rect 5000 9205 5170 9225
rect 5000 9175 5010 9205
rect 5040 9175 5170 9205
rect 5000 9135 5170 9175
rect 5000 9105 5010 9135
rect 5040 9105 5170 9135
rect 5000 9085 5170 9105
rect 5200 9205 5370 9225
rect 5200 9175 5210 9205
rect 5240 9175 5370 9205
rect 5200 9135 5370 9175
rect 5200 9105 5210 9135
rect 5240 9105 5370 9135
rect 5200 9085 5370 9105
rect 5400 9205 5570 9225
rect 5400 9175 5410 9205
rect 5440 9175 5570 9205
rect 5400 9135 5570 9175
rect 5400 9105 5410 9135
rect 5440 9105 5570 9135
rect 5400 9085 5570 9105
rect 5600 9205 5770 9225
rect 5600 9175 5610 9205
rect 5640 9175 5770 9205
rect 5600 9135 5770 9175
rect 5600 9105 5610 9135
rect 5640 9105 5770 9135
rect 5600 9085 5770 9105
rect 5800 9205 5970 9225
rect 5800 9175 5810 9205
rect 5840 9175 5970 9205
rect 5800 9135 5970 9175
rect 5800 9105 5810 9135
rect 5840 9105 5970 9135
rect 5800 9085 5970 9105
rect 6000 9205 6170 9225
rect 6000 9175 6010 9205
rect 6040 9175 6170 9205
rect 6000 9135 6170 9175
rect 6000 9105 6010 9135
rect 6040 9105 6170 9135
rect 6000 9085 6170 9105
rect 6200 9205 6370 9225
rect 6200 9175 6210 9205
rect 6240 9175 6370 9205
rect 6200 9135 6370 9175
rect 6200 9105 6210 9135
rect 6240 9105 6370 9135
rect 6200 9085 6370 9105
rect 6400 9205 6570 9225
rect 6400 9175 6410 9205
rect 6440 9175 6570 9205
rect 6400 9135 6570 9175
rect 6400 9105 6410 9135
rect 6440 9105 6570 9135
rect 6400 9085 6570 9105
rect -200 9020 -30 9040
rect -200 8990 -190 9020
rect -160 8990 -30 9020
rect -200 8950 -30 8990
rect -200 8920 -190 8950
rect -160 8920 -30 8950
rect -200 8900 -30 8920
rect 0 9020 170 9040
rect 0 8990 10 9020
rect 40 8990 170 9020
rect 0 8950 170 8990
rect 0 8920 10 8950
rect 40 8920 170 8950
rect 0 8900 170 8920
rect 200 9020 370 9040
rect 200 8990 210 9020
rect 240 8990 370 9020
rect 200 8950 370 8990
rect 200 8920 210 8950
rect 240 8920 370 8950
rect 200 8900 370 8920
rect 400 9020 570 9040
rect 400 8990 410 9020
rect 440 8990 570 9020
rect 400 8950 570 8990
rect 400 8920 410 8950
rect 440 8920 570 8950
rect 400 8900 570 8920
rect 600 9020 770 9040
rect 600 8990 610 9020
rect 640 8990 770 9020
rect 600 8950 770 8990
rect 600 8920 610 8950
rect 640 8920 770 8950
rect 600 8900 770 8920
rect 800 9020 970 9040
rect 800 8990 810 9020
rect 840 8990 970 9020
rect 800 8950 970 8990
rect 800 8920 810 8950
rect 840 8920 970 8950
rect 800 8900 970 8920
rect 1000 9020 1170 9040
rect 1000 8990 1010 9020
rect 1040 8990 1170 9020
rect 1000 8950 1170 8990
rect 1000 8920 1010 8950
rect 1040 8920 1170 8950
rect 1000 8900 1170 8920
rect 1200 9020 1370 9040
rect 1200 8990 1210 9020
rect 1240 8990 1370 9020
rect 1200 8950 1370 8990
rect 1200 8920 1210 8950
rect 1240 8920 1370 8950
rect 1200 8900 1370 8920
rect 1400 9020 1570 9040
rect 1400 8990 1410 9020
rect 1440 8990 1570 9020
rect 1400 8950 1570 8990
rect 1400 8920 1410 8950
rect 1440 8920 1570 8950
rect 1400 8900 1570 8920
rect 1600 9020 1770 9040
rect 1600 8990 1610 9020
rect 1640 8990 1770 9020
rect 1600 8950 1770 8990
rect 1600 8920 1610 8950
rect 1640 8920 1770 8950
rect 1600 8900 1770 8920
rect 1800 9020 1970 9040
rect 1800 8990 1810 9020
rect 1840 8990 1970 9020
rect 1800 8950 1970 8990
rect 1800 8920 1810 8950
rect 1840 8920 1970 8950
rect 1800 8900 1970 8920
rect 2000 9020 2170 9040
rect 2000 8990 2010 9020
rect 2040 8990 2170 9020
rect 2000 8950 2170 8990
rect 2000 8920 2010 8950
rect 2040 8920 2170 8950
rect 2000 8900 2170 8920
rect 2200 9020 2370 9040
rect 2200 8990 2210 9020
rect 2240 8990 2370 9020
rect 2200 8950 2370 8990
rect 2200 8920 2210 8950
rect 2240 8920 2370 8950
rect 2200 8900 2370 8920
rect 2400 9020 2570 9040
rect 2400 8990 2410 9020
rect 2440 8990 2570 9020
rect 2400 8950 2570 8990
rect 2400 8920 2410 8950
rect 2440 8920 2570 8950
rect 2400 8900 2570 8920
rect 2600 9020 2770 9040
rect 2600 8990 2610 9020
rect 2640 8990 2770 9020
rect 2600 8950 2770 8990
rect 2600 8920 2610 8950
rect 2640 8920 2770 8950
rect 2600 8900 2770 8920
rect 2800 9020 2970 9040
rect 2800 8990 2810 9020
rect 2840 8990 2970 9020
rect 2800 8950 2970 8990
rect 2800 8920 2810 8950
rect 2840 8920 2970 8950
rect 2800 8900 2970 8920
rect 3000 9020 3170 9040
rect 3000 8990 3010 9020
rect 3040 8990 3170 9020
rect 3000 8950 3170 8990
rect 3000 8920 3010 8950
rect 3040 8920 3170 8950
rect 3000 8900 3170 8920
rect 3200 9020 3370 9040
rect 3200 8990 3210 9020
rect 3240 8990 3370 9020
rect 3200 8950 3370 8990
rect 3200 8920 3210 8950
rect 3240 8920 3370 8950
rect 3200 8900 3370 8920
rect 3400 9020 3570 9040
rect 3400 8990 3410 9020
rect 3440 8990 3570 9020
rect 3400 8950 3570 8990
rect 3400 8920 3410 8950
rect 3440 8920 3570 8950
rect 3400 8900 3570 8920
rect 3600 9020 3770 9040
rect 3600 8990 3610 9020
rect 3640 8990 3770 9020
rect 3600 8950 3770 8990
rect 3600 8920 3610 8950
rect 3640 8920 3770 8950
rect 3600 8900 3770 8920
rect 3800 9020 3970 9040
rect 3800 8990 3810 9020
rect 3840 8990 3970 9020
rect 3800 8950 3970 8990
rect 3800 8920 3810 8950
rect 3840 8920 3970 8950
rect 3800 8900 3970 8920
rect 4000 9020 4170 9040
rect 4000 8990 4010 9020
rect 4040 8990 4170 9020
rect 4000 8950 4170 8990
rect 4000 8920 4010 8950
rect 4040 8920 4170 8950
rect 4000 8900 4170 8920
rect 4200 9020 4370 9040
rect 4200 8990 4210 9020
rect 4240 8990 4370 9020
rect 4200 8950 4370 8990
rect 4200 8920 4210 8950
rect 4240 8920 4370 8950
rect 4200 8900 4370 8920
rect 4400 9020 4570 9040
rect 4400 8990 4410 9020
rect 4440 8990 4570 9020
rect 4400 8950 4570 8990
rect 4400 8920 4410 8950
rect 4440 8920 4570 8950
rect 4400 8900 4570 8920
rect 4600 9020 4770 9040
rect 4600 8990 4610 9020
rect 4640 8990 4770 9020
rect 4600 8950 4770 8990
rect 4600 8920 4610 8950
rect 4640 8920 4770 8950
rect 4600 8900 4770 8920
rect 4800 9020 4970 9040
rect 4800 8990 4810 9020
rect 4840 8990 4970 9020
rect 4800 8950 4970 8990
rect 4800 8920 4810 8950
rect 4840 8920 4970 8950
rect 4800 8900 4970 8920
rect 5000 9020 5170 9040
rect 5000 8990 5010 9020
rect 5040 8990 5170 9020
rect 5000 8950 5170 8990
rect 5000 8920 5010 8950
rect 5040 8920 5170 8950
rect 5000 8900 5170 8920
rect 5200 9020 5370 9040
rect 5200 8990 5210 9020
rect 5240 8990 5370 9020
rect 5200 8950 5370 8990
rect 5200 8920 5210 8950
rect 5240 8920 5370 8950
rect 5200 8900 5370 8920
rect 5400 9020 5570 9040
rect 5400 8990 5410 9020
rect 5440 8990 5570 9020
rect 5400 8950 5570 8990
rect 5400 8920 5410 8950
rect 5440 8920 5570 8950
rect 5400 8900 5570 8920
rect 5600 9020 5770 9040
rect 5600 8990 5610 9020
rect 5640 8990 5770 9020
rect 5600 8950 5770 8990
rect 5600 8920 5610 8950
rect 5640 8920 5770 8950
rect 5600 8900 5770 8920
rect 5800 9020 5970 9040
rect 5800 8990 5810 9020
rect 5840 8990 5970 9020
rect 5800 8950 5970 8990
rect 5800 8920 5810 8950
rect 5840 8920 5970 8950
rect 5800 8900 5970 8920
rect 6000 9020 6170 9040
rect 6000 8990 6010 9020
rect 6040 8990 6170 9020
rect 6000 8950 6170 8990
rect 6000 8920 6010 8950
rect 6040 8920 6170 8950
rect 6000 8900 6170 8920
rect 6200 9020 6370 9040
rect 6200 8990 6210 9020
rect 6240 8990 6370 9020
rect 6200 8950 6370 8990
rect 6200 8920 6210 8950
rect 6240 8920 6370 8950
rect 6200 8900 6370 8920
rect 6400 9020 6570 9040
rect 6400 8990 6410 9020
rect 6440 8990 6570 9020
rect 6400 8950 6570 8990
rect 6400 8920 6410 8950
rect 6440 8920 6570 8950
rect 6400 8900 6570 8920
rect -200 8835 -30 8855
rect -200 8805 -190 8835
rect -160 8805 -30 8835
rect -200 8765 -30 8805
rect -200 8735 -190 8765
rect -160 8735 -30 8765
rect -200 8715 -30 8735
rect 0 8835 170 8855
rect 0 8805 10 8835
rect 40 8805 170 8835
rect 0 8765 170 8805
rect 0 8735 10 8765
rect 40 8735 170 8765
rect 0 8715 170 8735
rect 200 8835 370 8855
rect 200 8805 210 8835
rect 240 8805 370 8835
rect 200 8765 370 8805
rect 200 8735 210 8765
rect 240 8735 370 8765
rect 200 8715 370 8735
rect 400 8835 570 8855
rect 400 8805 410 8835
rect 440 8805 570 8835
rect 400 8765 570 8805
rect 400 8735 410 8765
rect 440 8735 570 8765
rect 400 8715 570 8735
rect 600 8835 770 8855
rect 600 8805 610 8835
rect 640 8805 770 8835
rect 600 8765 770 8805
rect 600 8735 610 8765
rect 640 8735 770 8765
rect 600 8715 770 8735
rect 800 8835 970 8855
rect 800 8805 810 8835
rect 840 8805 970 8835
rect 800 8765 970 8805
rect 800 8735 810 8765
rect 840 8735 970 8765
rect 800 8715 970 8735
rect 1000 8835 1170 8855
rect 1000 8805 1010 8835
rect 1040 8805 1170 8835
rect 1000 8765 1170 8805
rect 1000 8735 1010 8765
rect 1040 8735 1170 8765
rect 1000 8715 1170 8735
rect 1200 8835 1370 8855
rect 1200 8805 1210 8835
rect 1240 8805 1370 8835
rect 1200 8765 1370 8805
rect 1200 8735 1210 8765
rect 1240 8735 1370 8765
rect 1200 8715 1370 8735
rect 1400 8835 1570 8855
rect 1400 8805 1410 8835
rect 1440 8805 1570 8835
rect 1400 8765 1570 8805
rect 1400 8735 1410 8765
rect 1440 8735 1570 8765
rect 1400 8715 1570 8735
rect 1600 8835 1770 8855
rect 1600 8805 1610 8835
rect 1640 8805 1770 8835
rect 1600 8765 1770 8805
rect 1600 8735 1610 8765
rect 1640 8735 1770 8765
rect 1600 8715 1770 8735
rect 1800 8835 1970 8855
rect 1800 8805 1810 8835
rect 1840 8805 1970 8835
rect 1800 8765 1970 8805
rect 1800 8735 1810 8765
rect 1840 8735 1970 8765
rect 1800 8715 1970 8735
rect 2000 8835 2170 8855
rect 2000 8805 2010 8835
rect 2040 8805 2170 8835
rect 2000 8765 2170 8805
rect 2000 8735 2010 8765
rect 2040 8735 2170 8765
rect 2000 8715 2170 8735
rect 2200 8835 2370 8855
rect 2200 8805 2210 8835
rect 2240 8805 2370 8835
rect 2200 8765 2370 8805
rect 2200 8735 2210 8765
rect 2240 8735 2370 8765
rect 2200 8715 2370 8735
rect 2400 8835 2570 8855
rect 2400 8805 2410 8835
rect 2440 8805 2570 8835
rect 2400 8765 2570 8805
rect 2400 8735 2410 8765
rect 2440 8735 2570 8765
rect 2400 8715 2570 8735
rect 2600 8835 2770 8855
rect 2600 8805 2610 8835
rect 2640 8805 2770 8835
rect 2600 8765 2770 8805
rect 2600 8735 2610 8765
rect 2640 8735 2770 8765
rect 2600 8715 2770 8735
rect 2800 8835 2970 8855
rect 2800 8805 2810 8835
rect 2840 8805 2970 8835
rect 2800 8765 2970 8805
rect 2800 8735 2810 8765
rect 2840 8735 2970 8765
rect 2800 8715 2970 8735
rect 3000 8835 3170 8855
rect 3000 8805 3010 8835
rect 3040 8805 3170 8835
rect 3000 8765 3170 8805
rect 3000 8735 3010 8765
rect 3040 8735 3170 8765
rect 3000 8715 3170 8735
rect 3200 8835 3370 8855
rect 3200 8805 3210 8835
rect 3240 8805 3370 8835
rect 3200 8765 3370 8805
rect 3200 8735 3210 8765
rect 3240 8735 3370 8765
rect 3200 8715 3370 8735
rect 3400 8835 3570 8855
rect 3400 8805 3410 8835
rect 3440 8805 3570 8835
rect 3400 8765 3570 8805
rect 3400 8735 3410 8765
rect 3440 8735 3570 8765
rect 3400 8715 3570 8735
rect 3600 8835 3770 8855
rect 3600 8805 3610 8835
rect 3640 8805 3770 8835
rect 3600 8765 3770 8805
rect 3600 8735 3610 8765
rect 3640 8735 3770 8765
rect 3600 8715 3770 8735
rect 3800 8835 3970 8855
rect 3800 8805 3810 8835
rect 3840 8805 3970 8835
rect 3800 8765 3970 8805
rect 3800 8735 3810 8765
rect 3840 8735 3970 8765
rect 3800 8715 3970 8735
rect 4000 8835 4170 8855
rect 4000 8805 4010 8835
rect 4040 8805 4170 8835
rect 4000 8765 4170 8805
rect 4000 8735 4010 8765
rect 4040 8735 4170 8765
rect 4000 8715 4170 8735
rect 4200 8835 4370 8855
rect 4200 8805 4210 8835
rect 4240 8805 4370 8835
rect 4200 8765 4370 8805
rect 4200 8735 4210 8765
rect 4240 8735 4370 8765
rect 4200 8715 4370 8735
rect 4400 8835 4570 8855
rect 4400 8805 4410 8835
rect 4440 8805 4570 8835
rect 4400 8765 4570 8805
rect 4400 8735 4410 8765
rect 4440 8735 4570 8765
rect 4400 8715 4570 8735
rect 4600 8835 4770 8855
rect 4600 8805 4610 8835
rect 4640 8805 4770 8835
rect 4600 8765 4770 8805
rect 4600 8735 4610 8765
rect 4640 8735 4770 8765
rect 4600 8715 4770 8735
rect 4800 8835 4970 8855
rect 4800 8805 4810 8835
rect 4840 8805 4970 8835
rect 4800 8765 4970 8805
rect 4800 8735 4810 8765
rect 4840 8735 4970 8765
rect 4800 8715 4970 8735
rect 5000 8835 5170 8855
rect 5000 8805 5010 8835
rect 5040 8805 5170 8835
rect 5000 8765 5170 8805
rect 5000 8735 5010 8765
rect 5040 8735 5170 8765
rect 5000 8715 5170 8735
rect 5200 8835 5370 8855
rect 5200 8805 5210 8835
rect 5240 8805 5370 8835
rect 5200 8765 5370 8805
rect 5200 8735 5210 8765
rect 5240 8735 5370 8765
rect 5200 8715 5370 8735
rect 5400 8835 5570 8855
rect 5400 8805 5410 8835
rect 5440 8805 5570 8835
rect 5400 8765 5570 8805
rect 5400 8735 5410 8765
rect 5440 8735 5570 8765
rect 5400 8715 5570 8735
rect 5600 8835 5770 8855
rect 5600 8805 5610 8835
rect 5640 8805 5770 8835
rect 5600 8765 5770 8805
rect 5600 8735 5610 8765
rect 5640 8735 5770 8765
rect 5600 8715 5770 8735
rect 5800 8835 5970 8855
rect 5800 8805 5810 8835
rect 5840 8805 5970 8835
rect 5800 8765 5970 8805
rect 5800 8735 5810 8765
rect 5840 8735 5970 8765
rect 5800 8715 5970 8735
rect 6000 8835 6170 8855
rect 6000 8805 6010 8835
rect 6040 8805 6170 8835
rect 6000 8765 6170 8805
rect 6000 8735 6010 8765
rect 6040 8735 6170 8765
rect 6000 8715 6170 8735
rect 6200 8835 6370 8855
rect 6200 8805 6210 8835
rect 6240 8805 6370 8835
rect 6200 8765 6370 8805
rect 6200 8735 6210 8765
rect 6240 8735 6370 8765
rect 6200 8715 6370 8735
rect 6400 8835 6570 8855
rect 6400 8805 6410 8835
rect 6440 8805 6570 8835
rect 6400 8765 6570 8805
rect 6400 8735 6410 8765
rect 6440 8735 6570 8765
rect 6400 8715 6570 8735
rect -200 8650 -30 8670
rect -200 8620 -190 8650
rect -160 8620 -30 8650
rect -200 8580 -30 8620
rect -200 8550 -190 8580
rect -160 8550 -30 8580
rect -200 8530 -30 8550
rect 0 8650 170 8670
rect 0 8620 10 8650
rect 40 8620 170 8650
rect 0 8580 170 8620
rect 0 8550 10 8580
rect 40 8550 170 8580
rect 0 8530 170 8550
rect 200 8650 370 8670
rect 200 8620 210 8650
rect 240 8620 370 8650
rect 200 8580 370 8620
rect 200 8550 210 8580
rect 240 8550 370 8580
rect 200 8530 370 8550
rect 400 8650 570 8670
rect 400 8620 410 8650
rect 440 8620 570 8650
rect 400 8580 570 8620
rect 400 8550 410 8580
rect 440 8550 570 8580
rect 400 8530 570 8550
rect 600 8650 770 8670
rect 600 8620 610 8650
rect 640 8620 770 8650
rect 600 8580 770 8620
rect 600 8550 610 8580
rect 640 8550 770 8580
rect 600 8530 770 8550
rect 800 8650 970 8670
rect 800 8620 810 8650
rect 840 8620 970 8650
rect 800 8580 970 8620
rect 800 8550 810 8580
rect 840 8550 970 8580
rect 800 8530 970 8550
rect 1000 8650 1170 8670
rect 1000 8620 1010 8650
rect 1040 8620 1170 8650
rect 1000 8580 1170 8620
rect 1000 8550 1010 8580
rect 1040 8550 1170 8580
rect 1000 8530 1170 8550
rect 1200 8650 1370 8670
rect 1200 8620 1210 8650
rect 1240 8620 1370 8650
rect 1200 8580 1370 8620
rect 1200 8550 1210 8580
rect 1240 8550 1370 8580
rect 1200 8530 1370 8550
rect 1400 8650 1570 8670
rect 1400 8620 1410 8650
rect 1440 8620 1570 8650
rect 1400 8580 1570 8620
rect 1400 8550 1410 8580
rect 1440 8550 1570 8580
rect 1400 8530 1570 8550
rect 1600 8650 1770 8670
rect 1600 8620 1610 8650
rect 1640 8620 1770 8650
rect 1600 8580 1770 8620
rect 1600 8550 1610 8580
rect 1640 8550 1770 8580
rect 1600 8530 1770 8550
rect 1800 8650 1970 8670
rect 1800 8620 1810 8650
rect 1840 8620 1970 8650
rect 1800 8580 1970 8620
rect 1800 8550 1810 8580
rect 1840 8550 1970 8580
rect 1800 8530 1970 8550
rect 2000 8650 2170 8670
rect 2000 8620 2010 8650
rect 2040 8620 2170 8650
rect 2000 8580 2170 8620
rect 2000 8550 2010 8580
rect 2040 8550 2170 8580
rect 2000 8530 2170 8550
rect 2200 8650 2370 8670
rect 2200 8620 2210 8650
rect 2240 8620 2370 8650
rect 2200 8580 2370 8620
rect 2200 8550 2210 8580
rect 2240 8550 2370 8580
rect 2200 8530 2370 8550
rect 2400 8650 2570 8670
rect 2400 8620 2410 8650
rect 2440 8620 2570 8650
rect 2400 8580 2570 8620
rect 2400 8550 2410 8580
rect 2440 8550 2570 8580
rect 2400 8530 2570 8550
rect 2600 8650 2770 8670
rect 2600 8620 2610 8650
rect 2640 8620 2770 8650
rect 2600 8580 2770 8620
rect 2600 8550 2610 8580
rect 2640 8550 2770 8580
rect 2600 8530 2770 8550
rect 2800 8650 2970 8670
rect 2800 8620 2810 8650
rect 2840 8620 2970 8650
rect 2800 8580 2970 8620
rect 2800 8550 2810 8580
rect 2840 8550 2970 8580
rect 2800 8530 2970 8550
rect 3000 8650 3170 8670
rect 3000 8620 3010 8650
rect 3040 8620 3170 8650
rect 3000 8580 3170 8620
rect 3000 8550 3010 8580
rect 3040 8550 3170 8580
rect 3000 8530 3170 8550
rect 3200 8650 3370 8670
rect 3200 8620 3210 8650
rect 3240 8620 3370 8650
rect 3200 8580 3370 8620
rect 3200 8550 3210 8580
rect 3240 8550 3370 8580
rect 3200 8530 3370 8550
rect 3400 8650 3570 8670
rect 3400 8620 3410 8650
rect 3440 8620 3570 8650
rect 3400 8580 3570 8620
rect 3400 8550 3410 8580
rect 3440 8550 3570 8580
rect 3400 8530 3570 8550
rect 3600 8650 3770 8670
rect 3600 8620 3610 8650
rect 3640 8620 3770 8650
rect 3600 8580 3770 8620
rect 3600 8550 3610 8580
rect 3640 8550 3770 8580
rect 3600 8530 3770 8550
rect 3800 8650 3970 8670
rect 3800 8620 3810 8650
rect 3840 8620 3970 8650
rect 3800 8580 3970 8620
rect 3800 8550 3810 8580
rect 3840 8550 3970 8580
rect 3800 8530 3970 8550
rect 4000 8650 4170 8670
rect 4000 8620 4010 8650
rect 4040 8620 4170 8650
rect 4000 8580 4170 8620
rect 4000 8550 4010 8580
rect 4040 8550 4170 8580
rect 4000 8530 4170 8550
rect 4200 8650 4370 8670
rect 4200 8620 4210 8650
rect 4240 8620 4370 8650
rect 4200 8580 4370 8620
rect 4200 8550 4210 8580
rect 4240 8550 4370 8580
rect 4200 8530 4370 8550
rect 4400 8650 4570 8670
rect 4400 8620 4410 8650
rect 4440 8620 4570 8650
rect 4400 8580 4570 8620
rect 4400 8550 4410 8580
rect 4440 8550 4570 8580
rect 4400 8530 4570 8550
rect 4600 8650 4770 8670
rect 4600 8620 4610 8650
rect 4640 8620 4770 8650
rect 4600 8580 4770 8620
rect 4600 8550 4610 8580
rect 4640 8550 4770 8580
rect 4600 8530 4770 8550
rect 4800 8650 4970 8670
rect 4800 8620 4810 8650
rect 4840 8620 4970 8650
rect 4800 8580 4970 8620
rect 4800 8550 4810 8580
rect 4840 8550 4970 8580
rect 4800 8530 4970 8550
rect 5000 8650 5170 8670
rect 5000 8620 5010 8650
rect 5040 8620 5170 8650
rect 5000 8580 5170 8620
rect 5000 8550 5010 8580
rect 5040 8550 5170 8580
rect 5000 8530 5170 8550
rect 5200 8650 5370 8670
rect 5200 8620 5210 8650
rect 5240 8620 5370 8650
rect 5200 8580 5370 8620
rect 5200 8550 5210 8580
rect 5240 8550 5370 8580
rect 5200 8530 5370 8550
rect 5400 8650 5570 8670
rect 5400 8620 5410 8650
rect 5440 8620 5570 8650
rect 5400 8580 5570 8620
rect 5400 8550 5410 8580
rect 5440 8550 5570 8580
rect 5400 8530 5570 8550
rect 5600 8650 5770 8670
rect 5600 8620 5610 8650
rect 5640 8620 5770 8650
rect 5600 8580 5770 8620
rect 5600 8550 5610 8580
rect 5640 8550 5770 8580
rect 5600 8530 5770 8550
rect 5800 8650 5970 8670
rect 5800 8620 5810 8650
rect 5840 8620 5970 8650
rect 5800 8580 5970 8620
rect 5800 8550 5810 8580
rect 5840 8550 5970 8580
rect 5800 8530 5970 8550
rect 6000 8650 6170 8670
rect 6000 8620 6010 8650
rect 6040 8620 6170 8650
rect 6000 8580 6170 8620
rect 6000 8550 6010 8580
rect 6040 8550 6170 8580
rect 6000 8530 6170 8550
rect 6200 8650 6370 8670
rect 6200 8620 6210 8650
rect 6240 8620 6370 8650
rect 6200 8580 6370 8620
rect 6200 8550 6210 8580
rect 6240 8550 6370 8580
rect 6200 8530 6370 8550
rect 6400 8650 6570 8670
rect 6400 8620 6410 8650
rect 6440 8620 6570 8650
rect 6400 8580 6570 8620
rect 6400 8550 6410 8580
rect 6440 8550 6570 8580
rect 6400 8530 6570 8550
rect -200 8465 -30 8485
rect -200 8435 -190 8465
rect -160 8435 -30 8465
rect -200 8395 -30 8435
rect -200 8365 -190 8395
rect -160 8365 -30 8395
rect -200 8345 -30 8365
rect 0 8465 170 8485
rect 0 8435 10 8465
rect 40 8435 170 8465
rect 0 8395 170 8435
rect 0 8365 10 8395
rect 40 8365 170 8395
rect 0 8345 170 8365
rect 200 8465 370 8485
rect 200 8435 210 8465
rect 240 8435 370 8465
rect 200 8395 370 8435
rect 200 8365 210 8395
rect 240 8365 370 8395
rect 200 8345 370 8365
rect 400 8465 570 8485
rect 400 8435 410 8465
rect 440 8435 570 8465
rect 400 8395 570 8435
rect 400 8365 410 8395
rect 440 8365 570 8395
rect 400 8345 570 8365
rect 600 8465 770 8485
rect 600 8435 610 8465
rect 640 8435 770 8465
rect 600 8395 770 8435
rect 600 8365 610 8395
rect 640 8365 770 8395
rect 600 8345 770 8365
rect 800 8465 970 8485
rect 800 8435 810 8465
rect 840 8435 970 8465
rect 800 8395 970 8435
rect 800 8365 810 8395
rect 840 8365 970 8395
rect 800 8345 970 8365
rect 1000 8465 1170 8485
rect 1000 8435 1010 8465
rect 1040 8435 1170 8465
rect 1000 8395 1170 8435
rect 1000 8365 1010 8395
rect 1040 8365 1170 8395
rect 1000 8345 1170 8365
rect 1200 8465 1370 8485
rect 1200 8435 1210 8465
rect 1240 8435 1370 8465
rect 1200 8395 1370 8435
rect 1200 8365 1210 8395
rect 1240 8365 1370 8395
rect 1200 8345 1370 8365
rect 1400 8465 1570 8485
rect 1400 8435 1410 8465
rect 1440 8435 1570 8465
rect 1400 8395 1570 8435
rect 1400 8365 1410 8395
rect 1440 8365 1570 8395
rect 1400 8345 1570 8365
rect 1600 8465 1770 8485
rect 1600 8435 1610 8465
rect 1640 8435 1770 8465
rect 1600 8395 1770 8435
rect 1600 8365 1610 8395
rect 1640 8365 1770 8395
rect 1600 8345 1770 8365
rect 1800 8465 1970 8485
rect 1800 8435 1810 8465
rect 1840 8435 1970 8465
rect 1800 8395 1970 8435
rect 1800 8365 1810 8395
rect 1840 8365 1970 8395
rect 1800 8345 1970 8365
rect 2000 8465 2170 8485
rect 2000 8435 2010 8465
rect 2040 8435 2170 8465
rect 2000 8395 2170 8435
rect 2000 8365 2010 8395
rect 2040 8365 2170 8395
rect 2000 8345 2170 8365
rect 2200 8465 2370 8485
rect 2200 8435 2210 8465
rect 2240 8435 2370 8465
rect 2200 8395 2370 8435
rect 2200 8365 2210 8395
rect 2240 8365 2370 8395
rect 2200 8345 2370 8365
rect 2400 8465 2570 8485
rect 2400 8435 2410 8465
rect 2440 8435 2570 8465
rect 2400 8395 2570 8435
rect 2400 8365 2410 8395
rect 2440 8365 2570 8395
rect 2400 8345 2570 8365
rect 2600 8465 2770 8485
rect 2600 8435 2610 8465
rect 2640 8435 2770 8465
rect 2600 8395 2770 8435
rect 2600 8365 2610 8395
rect 2640 8365 2770 8395
rect 2600 8345 2770 8365
rect 2800 8465 2970 8485
rect 2800 8435 2810 8465
rect 2840 8435 2970 8465
rect 2800 8395 2970 8435
rect 2800 8365 2810 8395
rect 2840 8365 2970 8395
rect 2800 8345 2970 8365
rect 3000 8465 3170 8485
rect 3000 8435 3010 8465
rect 3040 8435 3170 8465
rect 3000 8395 3170 8435
rect 3000 8365 3010 8395
rect 3040 8365 3170 8395
rect 3000 8345 3170 8365
rect 3200 8465 3370 8485
rect 3200 8435 3210 8465
rect 3240 8435 3370 8465
rect 3200 8395 3370 8435
rect 3200 8365 3210 8395
rect 3240 8365 3370 8395
rect 3200 8345 3370 8365
rect 3400 8465 3570 8485
rect 3400 8435 3410 8465
rect 3440 8435 3570 8465
rect 3400 8395 3570 8435
rect 3400 8365 3410 8395
rect 3440 8365 3570 8395
rect 3400 8345 3570 8365
rect 3600 8465 3770 8485
rect 3600 8435 3610 8465
rect 3640 8435 3770 8465
rect 3600 8395 3770 8435
rect 3600 8365 3610 8395
rect 3640 8365 3770 8395
rect 3600 8345 3770 8365
rect 3800 8465 3970 8485
rect 3800 8435 3810 8465
rect 3840 8435 3970 8465
rect 3800 8395 3970 8435
rect 3800 8365 3810 8395
rect 3840 8365 3970 8395
rect 3800 8345 3970 8365
rect 4000 8465 4170 8485
rect 4000 8435 4010 8465
rect 4040 8435 4170 8465
rect 4000 8395 4170 8435
rect 4000 8365 4010 8395
rect 4040 8365 4170 8395
rect 4000 8345 4170 8365
rect 4200 8465 4370 8485
rect 4200 8435 4210 8465
rect 4240 8435 4370 8465
rect 4200 8395 4370 8435
rect 4200 8365 4210 8395
rect 4240 8365 4370 8395
rect 4200 8345 4370 8365
rect 4400 8465 4570 8485
rect 4400 8435 4410 8465
rect 4440 8435 4570 8465
rect 4400 8395 4570 8435
rect 4400 8365 4410 8395
rect 4440 8365 4570 8395
rect 4400 8345 4570 8365
rect 4600 8465 4770 8485
rect 4600 8435 4610 8465
rect 4640 8435 4770 8465
rect 4600 8395 4770 8435
rect 4600 8365 4610 8395
rect 4640 8365 4770 8395
rect 4600 8345 4770 8365
rect 4800 8465 4970 8485
rect 4800 8435 4810 8465
rect 4840 8435 4970 8465
rect 4800 8395 4970 8435
rect 4800 8365 4810 8395
rect 4840 8365 4970 8395
rect 4800 8345 4970 8365
rect 5000 8465 5170 8485
rect 5000 8435 5010 8465
rect 5040 8435 5170 8465
rect 5000 8395 5170 8435
rect 5000 8365 5010 8395
rect 5040 8365 5170 8395
rect 5000 8345 5170 8365
rect 5200 8465 5370 8485
rect 5200 8435 5210 8465
rect 5240 8435 5370 8465
rect 5200 8395 5370 8435
rect 5200 8365 5210 8395
rect 5240 8365 5370 8395
rect 5200 8345 5370 8365
rect 5400 8465 5570 8485
rect 5400 8435 5410 8465
rect 5440 8435 5570 8465
rect 5400 8395 5570 8435
rect 5400 8365 5410 8395
rect 5440 8365 5570 8395
rect 5400 8345 5570 8365
rect 5600 8465 5770 8485
rect 5600 8435 5610 8465
rect 5640 8435 5770 8465
rect 5600 8395 5770 8435
rect 5600 8365 5610 8395
rect 5640 8365 5770 8395
rect 5600 8345 5770 8365
rect 5800 8465 5970 8485
rect 5800 8435 5810 8465
rect 5840 8435 5970 8465
rect 5800 8395 5970 8435
rect 5800 8365 5810 8395
rect 5840 8365 5970 8395
rect 5800 8345 5970 8365
rect 6000 8465 6170 8485
rect 6000 8435 6010 8465
rect 6040 8435 6170 8465
rect 6000 8395 6170 8435
rect 6000 8365 6010 8395
rect 6040 8365 6170 8395
rect 6000 8345 6170 8365
rect 6200 8465 6370 8485
rect 6200 8435 6210 8465
rect 6240 8435 6370 8465
rect 6200 8395 6370 8435
rect 6200 8365 6210 8395
rect 6240 8365 6370 8395
rect 6200 8345 6370 8365
rect 6400 8465 6570 8485
rect 6400 8435 6410 8465
rect 6440 8435 6570 8465
rect 6400 8395 6570 8435
rect 6400 8365 6410 8395
rect 6440 8365 6570 8395
rect 6400 8345 6570 8365
rect -200 8280 -30 8300
rect -200 8250 -190 8280
rect -160 8250 -30 8280
rect -200 8210 -30 8250
rect -200 8180 -190 8210
rect -160 8180 -30 8210
rect -200 8160 -30 8180
rect 0 8280 170 8300
rect 0 8250 10 8280
rect 40 8250 170 8280
rect 0 8210 170 8250
rect 0 8180 10 8210
rect 40 8180 170 8210
rect 0 8160 170 8180
rect 200 8280 370 8300
rect 200 8250 210 8280
rect 240 8250 370 8280
rect 200 8210 370 8250
rect 200 8180 210 8210
rect 240 8180 370 8210
rect 200 8160 370 8180
rect 400 8280 570 8300
rect 400 8250 410 8280
rect 440 8250 570 8280
rect 400 8210 570 8250
rect 400 8180 410 8210
rect 440 8180 570 8210
rect 400 8160 570 8180
rect 600 8280 770 8300
rect 600 8250 610 8280
rect 640 8250 770 8280
rect 600 8210 770 8250
rect 600 8180 610 8210
rect 640 8180 770 8210
rect 600 8160 770 8180
rect 800 8280 970 8300
rect 800 8250 810 8280
rect 840 8250 970 8280
rect 800 8210 970 8250
rect 800 8180 810 8210
rect 840 8180 970 8210
rect 800 8160 970 8180
rect 1000 8280 1170 8300
rect 1000 8250 1010 8280
rect 1040 8250 1170 8280
rect 1000 8210 1170 8250
rect 1000 8180 1010 8210
rect 1040 8180 1170 8210
rect 1000 8160 1170 8180
rect 1200 8280 1370 8300
rect 1200 8250 1210 8280
rect 1240 8250 1370 8280
rect 1200 8210 1370 8250
rect 1200 8180 1210 8210
rect 1240 8180 1370 8210
rect 1200 8160 1370 8180
rect 1400 8280 1570 8300
rect 1400 8250 1410 8280
rect 1440 8250 1570 8280
rect 1400 8210 1570 8250
rect 1400 8180 1410 8210
rect 1440 8180 1570 8210
rect 1400 8160 1570 8180
rect 1600 8280 1770 8300
rect 1600 8250 1610 8280
rect 1640 8250 1770 8280
rect 1600 8210 1770 8250
rect 1600 8180 1610 8210
rect 1640 8180 1770 8210
rect 1600 8160 1770 8180
rect 1800 8280 1970 8300
rect 1800 8250 1810 8280
rect 1840 8250 1970 8280
rect 1800 8210 1970 8250
rect 1800 8180 1810 8210
rect 1840 8180 1970 8210
rect 1800 8160 1970 8180
rect 2000 8280 2170 8300
rect 2000 8250 2010 8280
rect 2040 8250 2170 8280
rect 2000 8210 2170 8250
rect 2000 8180 2010 8210
rect 2040 8180 2170 8210
rect 2000 8160 2170 8180
rect 2200 8280 2370 8300
rect 2200 8250 2210 8280
rect 2240 8250 2370 8280
rect 2200 8210 2370 8250
rect 2200 8180 2210 8210
rect 2240 8180 2370 8210
rect 2200 8160 2370 8180
rect 2400 8280 2570 8300
rect 2400 8250 2410 8280
rect 2440 8250 2570 8280
rect 2400 8210 2570 8250
rect 2400 8180 2410 8210
rect 2440 8180 2570 8210
rect 2400 8160 2570 8180
rect 2600 8280 2770 8300
rect 2600 8250 2610 8280
rect 2640 8250 2770 8280
rect 2600 8210 2770 8250
rect 2600 8180 2610 8210
rect 2640 8180 2770 8210
rect 2600 8160 2770 8180
rect 2800 8280 2970 8300
rect 2800 8250 2810 8280
rect 2840 8250 2970 8280
rect 2800 8210 2970 8250
rect 2800 8180 2810 8210
rect 2840 8180 2970 8210
rect 2800 8160 2970 8180
rect 3000 8280 3170 8300
rect 3000 8250 3010 8280
rect 3040 8250 3170 8280
rect 3000 8210 3170 8250
rect 3000 8180 3010 8210
rect 3040 8180 3170 8210
rect 3000 8160 3170 8180
rect 3200 8280 3370 8300
rect 3200 8250 3210 8280
rect 3240 8250 3370 8280
rect 3200 8210 3370 8250
rect 3200 8180 3210 8210
rect 3240 8180 3370 8210
rect 3200 8160 3370 8180
rect 3400 8280 3570 8300
rect 3400 8250 3410 8280
rect 3440 8250 3570 8280
rect 3400 8210 3570 8250
rect 3400 8180 3410 8210
rect 3440 8180 3570 8210
rect 3400 8160 3570 8180
rect 3600 8280 3770 8300
rect 3600 8250 3610 8280
rect 3640 8250 3770 8280
rect 3600 8210 3770 8250
rect 3600 8180 3610 8210
rect 3640 8180 3770 8210
rect 3600 8160 3770 8180
rect 3800 8280 3970 8300
rect 3800 8250 3810 8280
rect 3840 8250 3970 8280
rect 3800 8210 3970 8250
rect 3800 8180 3810 8210
rect 3840 8180 3970 8210
rect 3800 8160 3970 8180
rect 4000 8280 4170 8300
rect 4000 8250 4010 8280
rect 4040 8250 4170 8280
rect 4000 8210 4170 8250
rect 4000 8180 4010 8210
rect 4040 8180 4170 8210
rect 4000 8160 4170 8180
rect 4200 8280 4370 8300
rect 4200 8250 4210 8280
rect 4240 8250 4370 8280
rect 4200 8210 4370 8250
rect 4200 8180 4210 8210
rect 4240 8180 4370 8210
rect 4200 8160 4370 8180
rect 4400 8280 4570 8300
rect 4400 8250 4410 8280
rect 4440 8250 4570 8280
rect 4400 8210 4570 8250
rect 4400 8180 4410 8210
rect 4440 8180 4570 8210
rect 4400 8160 4570 8180
rect 4600 8280 4770 8300
rect 4600 8250 4610 8280
rect 4640 8250 4770 8280
rect 4600 8210 4770 8250
rect 4600 8180 4610 8210
rect 4640 8180 4770 8210
rect 4600 8160 4770 8180
rect 4800 8280 4970 8300
rect 4800 8250 4810 8280
rect 4840 8250 4970 8280
rect 4800 8210 4970 8250
rect 4800 8180 4810 8210
rect 4840 8180 4970 8210
rect 4800 8160 4970 8180
rect 5000 8280 5170 8300
rect 5000 8250 5010 8280
rect 5040 8250 5170 8280
rect 5000 8210 5170 8250
rect 5000 8180 5010 8210
rect 5040 8180 5170 8210
rect 5000 8160 5170 8180
rect 5200 8280 5370 8300
rect 5200 8250 5210 8280
rect 5240 8250 5370 8280
rect 5200 8210 5370 8250
rect 5200 8180 5210 8210
rect 5240 8180 5370 8210
rect 5200 8160 5370 8180
rect 5400 8280 5570 8300
rect 5400 8250 5410 8280
rect 5440 8250 5570 8280
rect 5400 8210 5570 8250
rect 5400 8180 5410 8210
rect 5440 8180 5570 8210
rect 5400 8160 5570 8180
rect 5600 8280 5770 8300
rect 5600 8250 5610 8280
rect 5640 8250 5770 8280
rect 5600 8210 5770 8250
rect 5600 8180 5610 8210
rect 5640 8180 5770 8210
rect 5600 8160 5770 8180
rect 5800 8280 5970 8300
rect 5800 8250 5810 8280
rect 5840 8250 5970 8280
rect 5800 8210 5970 8250
rect 5800 8180 5810 8210
rect 5840 8180 5970 8210
rect 5800 8160 5970 8180
rect 6000 8280 6170 8300
rect 6000 8250 6010 8280
rect 6040 8250 6170 8280
rect 6000 8210 6170 8250
rect 6000 8180 6010 8210
rect 6040 8180 6170 8210
rect 6000 8160 6170 8180
rect 6200 8280 6370 8300
rect 6200 8250 6210 8280
rect 6240 8250 6370 8280
rect 6200 8210 6370 8250
rect 6200 8180 6210 8210
rect 6240 8180 6370 8210
rect 6200 8160 6370 8180
rect 6400 8280 6570 8300
rect 6400 8250 6410 8280
rect 6440 8250 6570 8280
rect 6400 8210 6570 8250
rect 6400 8180 6410 8210
rect 6440 8180 6570 8210
rect 6400 8160 6570 8180
rect -200 8095 -30 8115
rect -200 8065 -190 8095
rect -160 8065 -30 8095
rect -200 8025 -30 8065
rect -200 7995 -190 8025
rect -160 7995 -30 8025
rect -200 7975 -30 7995
rect 0 8095 170 8115
rect 0 8065 10 8095
rect 40 8065 170 8095
rect 0 8025 170 8065
rect 0 7995 10 8025
rect 40 7995 170 8025
rect 0 7975 170 7995
rect 200 8095 370 8115
rect 200 8065 210 8095
rect 240 8065 370 8095
rect 200 8025 370 8065
rect 200 7995 210 8025
rect 240 7995 370 8025
rect 200 7975 370 7995
rect 400 8095 570 8115
rect 400 8065 410 8095
rect 440 8065 570 8095
rect 400 8025 570 8065
rect 400 7995 410 8025
rect 440 7995 570 8025
rect 400 7975 570 7995
rect 600 8095 770 8115
rect 600 8065 610 8095
rect 640 8065 770 8095
rect 600 8025 770 8065
rect 600 7995 610 8025
rect 640 7995 770 8025
rect 600 7975 770 7995
rect 800 8095 970 8115
rect 800 8065 810 8095
rect 840 8065 970 8095
rect 800 8025 970 8065
rect 800 7995 810 8025
rect 840 7995 970 8025
rect 800 7975 970 7995
rect 1000 8095 1170 8115
rect 1000 8065 1010 8095
rect 1040 8065 1170 8095
rect 1000 8025 1170 8065
rect 1000 7995 1010 8025
rect 1040 7995 1170 8025
rect 1000 7975 1170 7995
rect 1200 8095 1370 8115
rect 1200 8065 1210 8095
rect 1240 8065 1370 8095
rect 1200 8025 1370 8065
rect 1200 7995 1210 8025
rect 1240 7995 1370 8025
rect 1200 7975 1370 7995
rect 1400 8095 1570 8115
rect 1400 8065 1410 8095
rect 1440 8065 1570 8095
rect 1400 8025 1570 8065
rect 1400 7995 1410 8025
rect 1440 7995 1570 8025
rect 1400 7975 1570 7995
rect 1600 8095 1770 8115
rect 1600 8065 1610 8095
rect 1640 8065 1770 8095
rect 1600 8025 1770 8065
rect 1600 7995 1610 8025
rect 1640 7995 1770 8025
rect 1600 7975 1770 7995
rect 1800 8095 1970 8115
rect 1800 8065 1810 8095
rect 1840 8065 1970 8095
rect 1800 8025 1970 8065
rect 1800 7995 1810 8025
rect 1840 7995 1970 8025
rect 1800 7975 1970 7995
rect 2000 8095 2170 8115
rect 2000 8065 2010 8095
rect 2040 8065 2170 8095
rect 2000 8025 2170 8065
rect 2000 7995 2010 8025
rect 2040 7995 2170 8025
rect 2000 7975 2170 7995
rect 2200 8095 2370 8115
rect 2200 8065 2210 8095
rect 2240 8065 2370 8095
rect 2200 8025 2370 8065
rect 2200 7995 2210 8025
rect 2240 7995 2370 8025
rect 2200 7975 2370 7995
rect 2400 8095 2570 8115
rect 2400 8065 2410 8095
rect 2440 8065 2570 8095
rect 2400 8025 2570 8065
rect 2400 7995 2410 8025
rect 2440 7995 2570 8025
rect 2400 7975 2570 7995
rect 2600 8095 2770 8115
rect 2600 8065 2610 8095
rect 2640 8065 2770 8095
rect 2600 8025 2770 8065
rect 2600 7995 2610 8025
rect 2640 7995 2770 8025
rect 2600 7975 2770 7995
rect 2800 8095 2970 8115
rect 2800 8065 2810 8095
rect 2840 8065 2970 8095
rect 2800 8025 2970 8065
rect 2800 7995 2810 8025
rect 2840 7995 2970 8025
rect 2800 7975 2970 7995
rect 3000 8095 3170 8115
rect 3000 8065 3010 8095
rect 3040 8065 3170 8095
rect 3000 8025 3170 8065
rect 3000 7995 3010 8025
rect 3040 7995 3170 8025
rect 3000 7975 3170 7995
rect 3200 8095 3370 8115
rect 3200 8065 3210 8095
rect 3240 8065 3370 8095
rect 3200 8025 3370 8065
rect 3200 7995 3210 8025
rect 3240 7995 3370 8025
rect 3200 7975 3370 7995
rect 3400 8095 3570 8115
rect 3400 8065 3410 8095
rect 3440 8065 3570 8095
rect 3400 8025 3570 8065
rect 3400 7995 3410 8025
rect 3440 7995 3570 8025
rect 3400 7975 3570 7995
rect 3600 8095 3770 8115
rect 3600 8065 3610 8095
rect 3640 8065 3770 8095
rect 3600 8025 3770 8065
rect 3600 7995 3610 8025
rect 3640 7995 3770 8025
rect 3600 7975 3770 7995
rect 3800 8095 3970 8115
rect 3800 8065 3810 8095
rect 3840 8065 3970 8095
rect 3800 8025 3970 8065
rect 3800 7995 3810 8025
rect 3840 7995 3970 8025
rect 3800 7975 3970 7995
rect 4000 8095 4170 8115
rect 4000 8065 4010 8095
rect 4040 8065 4170 8095
rect 4000 8025 4170 8065
rect 4000 7995 4010 8025
rect 4040 7995 4170 8025
rect 4000 7975 4170 7995
rect 4200 8095 4370 8115
rect 4200 8065 4210 8095
rect 4240 8065 4370 8095
rect 4200 8025 4370 8065
rect 4200 7995 4210 8025
rect 4240 7995 4370 8025
rect 4200 7975 4370 7995
rect 4400 8095 4570 8115
rect 4400 8065 4410 8095
rect 4440 8065 4570 8095
rect 4400 8025 4570 8065
rect 4400 7995 4410 8025
rect 4440 7995 4570 8025
rect 4400 7975 4570 7995
rect 4600 8095 4770 8115
rect 4600 8065 4610 8095
rect 4640 8065 4770 8095
rect 4600 8025 4770 8065
rect 4600 7995 4610 8025
rect 4640 7995 4770 8025
rect 4600 7975 4770 7995
rect 4800 8095 4970 8115
rect 4800 8065 4810 8095
rect 4840 8065 4970 8095
rect 4800 8025 4970 8065
rect 4800 7995 4810 8025
rect 4840 7995 4970 8025
rect 4800 7975 4970 7995
rect 5000 8095 5170 8115
rect 5000 8065 5010 8095
rect 5040 8065 5170 8095
rect 5000 8025 5170 8065
rect 5000 7995 5010 8025
rect 5040 7995 5170 8025
rect 5000 7975 5170 7995
rect 5200 8095 5370 8115
rect 5200 8065 5210 8095
rect 5240 8065 5370 8095
rect 5200 8025 5370 8065
rect 5200 7995 5210 8025
rect 5240 7995 5370 8025
rect 5200 7975 5370 7995
rect 5400 8095 5570 8115
rect 5400 8065 5410 8095
rect 5440 8065 5570 8095
rect 5400 8025 5570 8065
rect 5400 7995 5410 8025
rect 5440 7995 5570 8025
rect 5400 7975 5570 7995
rect 5600 8095 5770 8115
rect 5600 8065 5610 8095
rect 5640 8065 5770 8095
rect 5600 8025 5770 8065
rect 5600 7995 5610 8025
rect 5640 7995 5770 8025
rect 5600 7975 5770 7995
rect 5800 8095 5970 8115
rect 5800 8065 5810 8095
rect 5840 8065 5970 8095
rect 5800 8025 5970 8065
rect 5800 7995 5810 8025
rect 5840 7995 5970 8025
rect 5800 7975 5970 7995
rect 6000 8095 6170 8115
rect 6000 8065 6010 8095
rect 6040 8065 6170 8095
rect 6000 8025 6170 8065
rect 6000 7995 6010 8025
rect 6040 7995 6170 8025
rect 6000 7975 6170 7995
rect 6200 8095 6370 8115
rect 6200 8065 6210 8095
rect 6240 8065 6370 8095
rect 6200 8025 6370 8065
rect 6200 7995 6210 8025
rect 6240 7995 6370 8025
rect 6200 7975 6370 7995
rect 6400 8095 6570 8115
rect 6400 8065 6410 8095
rect 6440 8065 6570 8095
rect 6400 8025 6570 8065
rect 6400 7995 6410 8025
rect 6440 7995 6570 8025
rect 6400 7975 6570 7995
rect -200 7910 -30 7930
rect -200 7880 -190 7910
rect -160 7880 -30 7910
rect -200 7840 -30 7880
rect -200 7810 -190 7840
rect -160 7810 -30 7840
rect -200 7790 -30 7810
rect 0 7910 170 7930
rect 0 7880 10 7910
rect 40 7880 170 7910
rect 0 7840 170 7880
rect 0 7810 10 7840
rect 40 7810 170 7840
rect 0 7790 170 7810
rect 200 7910 370 7930
rect 200 7880 210 7910
rect 240 7880 370 7910
rect 200 7840 370 7880
rect 200 7810 210 7840
rect 240 7810 370 7840
rect 200 7790 370 7810
rect 400 7910 570 7930
rect 400 7880 410 7910
rect 440 7880 570 7910
rect 400 7840 570 7880
rect 400 7810 410 7840
rect 440 7810 570 7840
rect 400 7790 570 7810
rect 600 7910 770 7930
rect 600 7880 610 7910
rect 640 7880 770 7910
rect 600 7840 770 7880
rect 600 7810 610 7840
rect 640 7810 770 7840
rect 600 7790 770 7810
rect 800 7910 970 7930
rect 800 7880 810 7910
rect 840 7880 970 7910
rect 800 7840 970 7880
rect 800 7810 810 7840
rect 840 7810 970 7840
rect 800 7790 970 7810
rect 1000 7910 1170 7930
rect 1000 7880 1010 7910
rect 1040 7880 1170 7910
rect 1000 7840 1170 7880
rect 1000 7810 1010 7840
rect 1040 7810 1170 7840
rect 1000 7790 1170 7810
rect 1200 7910 1370 7930
rect 1200 7880 1210 7910
rect 1240 7880 1370 7910
rect 1200 7840 1370 7880
rect 1200 7810 1210 7840
rect 1240 7810 1370 7840
rect 1200 7790 1370 7810
rect 1400 7910 1570 7930
rect 1400 7880 1410 7910
rect 1440 7880 1570 7910
rect 1400 7840 1570 7880
rect 1400 7810 1410 7840
rect 1440 7810 1570 7840
rect 1400 7790 1570 7810
rect 1600 7910 1770 7930
rect 1600 7880 1610 7910
rect 1640 7880 1770 7910
rect 1600 7840 1770 7880
rect 1600 7810 1610 7840
rect 1640 7810 1770 7840
rect 1600 7790 1770 7810
rect 1800 7910 1970 7930
rect 1800 7880 1810 7910
rect 1840 7880 1970 7910
rect 1800 7840 1970 7880
rect 1800 7810 1810 7840
rect 1840 7810 1970 7840
rect 1800 7790 1970 7810
rect 2000 7910 2170 7930
rect 2000 7880 2010 7910
rect 2040 7880 2170 7910
rect 2000 7840 2170 7880
rect 2000 7810 2010 7840
rect 2040 7810 2170 7840
rect 2000 7790 2170 7810
rect 2200 7910 2370 7930
rect 2200 7880 2210 7910
rect 2240 7880 2370 7910
rect 2200 7840 2370 7880
rect 2200 7810 2210 7840
rect 2240 7810 2370 7840
rect 2200 7790 2370 7810
rect 2400 7910 2570 7930
rect 2400 7880 2410 7910
rect 2440 7880 2570 7910
rect 2400 7840 2570 7880
rect 2400 7810 2410 7840
rect 2440 7810 2570 7840
rect 2400 7790 2570 7810
rect 2600 7910 2770 7930
rect 2600 7880 2610 7910
rect 2640 7880 2770 7910
rect 2600 7840 2770 7880
rect 2600 7810 2610 7840
rect 2640 7810 2770 7840
rect 2600 7790 2770 7810
rect 2800 7910 2970 7930
rect 2800 7880 2810 7910
rect 2840 7880 2970 7910
rect 2800 7840 2970 7880
rect 2800 7810 2810 7840
rect 2840 7810 2970 7840
rect 2800 7790 2970 7810
rect 3000 7910 3170 7930
rect 3000 7880 3010 7910
rect 3040 7880 3170 7910
rect 3000 7840 3170 7880
rect 3000 7810 3010 7840
rect 3040 7810 3170 7840
rect 3000 7790 3170 7810
rect 3200 7910 3370 7930
rect 3200 7880 3210 7910
rect 3240 7880 3370 7910
rect 3200 7840 3370 7880
rect 3200 7810 3210 7840
rect 3240 7810 3370 7840
rect 3200 7790 3370 7810
rect 3400 7910 3570 7930
rect 3400 7880 3410 7910
rect 3440 7880 3570 7910
rect 3400 7840 3570 7880
rect 3400 7810 3410 7840
rect 3440 7810 3570 7840
rect 3400 7790 3570 7810
rect 3600 7910 3770 7930
rect 3600 7880 3610 7910
rect 3640 7880 3770 7910
rect 3600 7840 3770 7880
rect 3600 7810 3610 7840
rect 3640 7810 3770 7840
rect 3600 7790 3770 7810
rect 3800 7910 3970 7930
rect 3800 7880 3810 7910
rect 3840 7880 3970 7910
rect 3800 7840 3970 7880
rect 3800 7810 3810 7840
rect 3840 7810 3970 7840
rect 3800 7790 3970 7810
rect 4000 7910 4170 7930
rect 4000 7880 4010 7910
rect 4040 7880 4170 7910
rect 4000 7840 4170 7880
rect 4000 7810 4010 7840
rect 4040 7810 4170 7840
rect 4000 7790 4170 7810
rect 4200 7910 4370 7930
rect 4200 7880 4210 7910
rect 4240 7880 4370 7910
rect 4200 7840 4370 7880
rect 4200 7810 4210 7840
rect 4240 7810 4370 7840
rect 4200 7790 4370 7810
rect 4400 7910 4570 7930
rect 4400 7880 4410 7910
rect 4440 7880 4570 7910
rect 4400 7840 4570 7880
rect 4400 7810 4410 7840
rect 4440 7810 4570 7840
rect 4400 7790 4570 7810
rect 4600 7910 4770 7930
rect 4600 7880 4610 7910
rect 4640 7880 4770 7910
rect 4600 7840 4770 7880
rect 4600 7810 4610 7840
rect 4640 7810 4770 7840
rect 4600 7790 4770 7810
rect 4800 7910 4970 7930
rect 4800 7880 4810 7910
rect 4840 7880 4970 7910
rect 4800 7840 4970 7880
rect 4800 7810 4810 7840
rect 4840 7810 4970 7840
rect 4800 7790 4970 7810
rect 5000 7910 5170 7930
rect 5000 7880 5010 7910
rect 5040 7880 5170 7910
rect 5000 7840 5170 7880
rect 5000 7810 5010 7840
rect 5040 7810 5170 7840
rect 5000 7790 5170 7810
rect 5200 7910 5370 7930
rect 5200 7880 5210 7910
rect 5240 7880 5370 7910
rect 5200 7840 5370 7880
rect 5200 7810 5210 7840
rect 5240 7810 5370 7840
rect 5200 7790 5370 7810
rect 5400 7910 5570 7930
rect 5400 7880 5410 7910
rect 5440 7880 5570 7910
rect 5400 7840 5570 7880
rect 5400 7810 5410 7840
rect 5440 7810 5570 7840
rect 5400 7790 5570 7810
rect 5600 7910 5770 7930
rect 5600 7880 5610 7910
rect 5640 7880 5770 7910
rect 5600 7840 5770 7880
rect 5600 7810 5610 7840
rect 5640 7810 5770 7840
rect 5600 7790 5770 7810
rect 5800 7910 5970 7930
rect 5800 7880 5810 7910
rect 5840 7880 5970 7910
rect 5800 7840 5970 7880
rect 5800 7810 5810 7840
rect 5840 7810 5970 7840
rect 5800 7790 5970 7810
rect 6000 7910 6170 7930
rect 6000 7880 6010 7910
rect 6040 7880 6170 7910
rect 6000 7840 6170 7880
rect 6000 7810 6010 7840
rect 6040 7810 6170 7840
rect 6000 7790 6170 7810
rect 6200 7910 6370 7930
rect 6200 7880 6210 7910
rect 6240 7880 6370 7910
rect 6200 7840 6370 7880
rect 6200 7810 6210 7840
rect 6240 7810 6370 7840
rect 6200 7790 6370 7810
rect 6400 7910 6570 7930
rect 6400 7880 6410 7910
rect 6440 7880 6570 7910
rect 6400 7840 6570 7880
rect 6400 7810 6410 7840
rect 6440 7810 6570 7840
rect 6400 7790 6570 7810
rect -200 7725 -30 7745
rect -200 7695 -190 7725
rect -160 7695 -30 7725
rect -200 7655 -30 7695
rect -200 7625 -190 7655
rect -160 7625 -30 7655
rect -200 7605 -30 7625
rect 0 7725 170 7745
rect 0 7695 10 7725
rect 40 7695 170 7725
rect 0 7655 170 7695
rect 0 7625 10 7655
rect 40 7625 170 7655
rect 0 7605 170 7625
rect 200 7725 370 7745
rect 200 7695 210 7725
rect 240 7695 370 7725
rect 200 7655 370 7695
rect 200 7625 210 7655
rect 240 7625 370 7655
rect 200 7605 370 7625
rect 400 7725 570 7745
rect 400 7695 410 7725
rect 440 7695 570 7725
rect 400 7655 570 7695
rect 400 7625 410 7655
rect 440 7625 570 7655
rect 400 7605 570 7625
rect 600 7725 770 7745
rect 600 7695 610 7725
rect 640 7695 770 7725
rect 600 7655 770 7695
rect 600 7625 610 7655
rect 640 7625 770 7655
rect 600 7605 770 7625
rect 800 7725 970 7745
rect 800 7695 810 7725
rect 840 7695 970 7725
rect 800 7655 970 7695
rect 800 7625 810 7655
rect 840 7625 970 7655
rect 800 7605 970 7625
rect 1000 7725 1170 7745
rect 1000 7695 1010 7725
rect 1040 7695 1170 7725
rect 1000 7655 1170 7695
rect 1000 7625 1010 7655
rect 1040 7625 1170 7655
rect 1000 7605 1170 7625
rect 1200 7725 1370 7745
rect 1200 7695 1210 7725
rect 1240 7695 1370 7725
rect 1200 7655 1370 7695
rect 1200 7625 1210 7655
rect 1240 7625 1370 7655
rect 1200 7605 1370 7625
rect 1400 7725 1570 7745
rect 1400 7695 1410 7725
rect 1440 7695 1570 7725
rect 1400 7655 1570 7695
rect 1400 7625 1410 7655
rect 1440 7625 1570 7655
rect 1400 7605 1570 7625
rect 1600 7725 1770 7745
rect 1600 7695 1610 7725
rect 1640 7695 1770 7725
rect 1600 7655 1770 7695
rect 1600 7625 1610 7655
rect 1640 7625 1770 7655
rect 1600 7605 1770 7625
rect 1800 7725 1970 7745
rect 1800 7695 1810 7725
rect 1840 7695 1970 7725
rect 1800 7655 1970 7695
rect 1800 7625 1810 7655
rect 1840 7625 1970 7655
rect 1800 7605 1970 7625
rect 2000 7725 2170 7745
rect 2000 7695 2010 7725
rect 2040 7695 2170 7725
rect 2000 7655 2170 7695
rect 2000 7625 2010 7655
rect 2040 7625 2170 7655
rect 2000 7605 2170 7625
rect 2200 7725 2370 7745
rect 2200 7695 2210 7725
rect 2240 7695 2370 7725
rect 2200 7655 2370 7695
rect 2200 7625 2210 7655
rect 2240 7625 2370 7655
rect 2200 7605 2370 7625
rect 2400 7725 2570 7745
rect 2400 7695 2410 7725
rect 2440 7695 2570 7725
rect 2400 7655 2570 7695
rect 2400 7625 2410 7655
rect 2440 7625 2570 7655
rect 2400 7605 2570 7625
rect 2600 7725 2770 7745
rect 2600 7695 2610 7725
rect 2640 7695 2770 7725
rect 2600 7655 2770 7695
rect 2600 7625 2610 7655
rect 2640 7625 2770 7655
rect 2600 7605 2770 7625
rect 2800 7725 2970 7745
rect 2800 7695 2810 7725
rect 2840 7695 2970 7725
rect 2800 7655 2970 7695
rect 2800 7625 2810 7655
rect 2840 7625 2970 7655
rect 2800 7605 2970 7625
rect 3000 7725 3170 7745
rect 3000 7695 3010 7725
rect 3040 7695 3170 7725
rect 3000 7655 3170 7695
rect 3000 7625 3010 7655
rect 3040 7625 3170 7655
rect 3000 7605 3170 7625
rect 3200 7725 3370 7745
rect 3200 7695 3210 7725
rect 3240 7695 3370 7725
rect 3200 7655 3370 7695
rect 3200 7625 3210 7655
rect 3240 7625 3370 7655
rect 3200 7605 3370 7625
rect 3400 7725 3570 7745
rect 3400 7695 3410 7725
rect 3440 7695 3570 7725
rect 3400 7655 3570 7695
rect 3400 7625 3410 7655
rect 3440 7625 3570 7655
rect 3400 7605 3570 7625
rect 3600 7725 3770 7745
rect 3600 7695 3610 7725
rect 3640 7695 3770 7725
rect 3600 7655 3770 7695
rect 3600 7625 3610 7655
rect 3640 7625 3770 7655
rect 3600 7605 3770 7625
rect 3800 7725 3970 7745
rect 3800 7695 3810 7725
rect 3840 7695 3970 7725
rect 3800 7655 3970 7695
rect 3800 7625 3810 7655
rect 3840 7625 3970 7655
rect 3800 7605 3970 7625
rect 4000 7725 4170 7745
rect 4000 7695 4010 7725
rect 4040 7695 4170 7725
rect 4000 7655 4170 7695
rect 4000 7625 4010 7655
rect 4040 7625 4170 7655
rect 4000 7605 4170 7625
rect 4200 7725 4370 7745
rect 4200 7695 4210 7725
rect 4240 7695 4370 7725
rect 4200 7655 4370 7695
rect 4200 7625 4210 7655
rect 4240 7625 4370 7655
rect 4200 7605 4370 7625
rect 4400 7725 4570 7745
rect 4400 7695 4410 7725
rect 4440 7695 4570 7725
rect 4400 7655 4570 7695
rect 4400 7625 4410 7655
rect 4440 7625 4570 7655
rect 4400 7605 4570 7625
rect 4600 7725 4770 7745
rect 4600 7695 4610 7725
rect 4640 7695 4770 7725
rect 4600 7655 4770 7695
rect 4600 7625 4610 7655
rect 4640 7625 4770 7655
rect 4600 7605 4770 7625
rect 4800 7725 4970 7745
rect 4800 7695 4810 7725
rect 4840 7695 4970 7725
rect 4800 7655 4970 7695
rect 4800 7625 4810 7655
rect 4840 7625 4970 7655
rect 4800 7605 4970 7625
rect 5000 7725 5170 7745
rect 5000 7695 5010 7725
rect 5040 7695 5170 7725
rect 5000 7655 5170 7695
rect 5000 7625 5010 7655
rect 5040 7625 5170 7655
rect 5000 7605 5170 7625
rect 5200 7725 5370 7745
rect 5200 7695 5210 7725
rect 5240 7695 5370 7725
rect 5200 7655 5370 7695
rect 5200 7625 5210 7655
rect 5240 7625 5370 7655
rect 5200 7605 5370 7625
rect 5400 7725 5570 7745
rect 5400 7695 5410 7725
rect 5440 7695 5570 7725
rect 5400 7655 5570 7695
rect 5400 7625 5410 7655
rect 5440 7625 5570 7655
rect 5400 7605 5570 7625
rect 5600 7725 5770 7745
rect 5600 7695 5610 7725
rect 5640 7695 5770 7725
rect 5600 7655 5770 7695
rect 5600 7625 5610 7655
rect 5640 7625 5770 7655
rect 5600 7605 5770 7625
rect 5800 7725 5970 7745
rect 5800 7695 5810 7725
rect 5840 7695 5970 7725
rect 5800 7655 5970 7695
rect 5800 7625 5810 7655
rect 5840 7625 5970 7655
rect 5800 7605 5970 7625
rect 6000 7725 6170 7745
rect 6000 7695 6010 7725
rect 6040 7695 6170 7725
rect 6000 7655 6170 7695
rect 6000 7625 6010 7655
rect 6040 7625 6170 7655
rect 6000 7605 6170 7625
rect 6200 7725 6370 7745
rect 6200 7695 6210 7725
rect 6240 7695 6370 7725
rect 6200 7655 6370 7695
rect 6200 7625 6210 7655
rect 6240 7625 6370 7655
rect 6200 7605 6370 7625
rect 6400 7725 6570 7745
rect 6400 7695 6410 7725
rect 6440 7695 6570 7725
rect 6400 7655 6570 7695
rect 6400 7625 6410 7655
rect 6440 7625 6570 7655
rect 6400 7605 6570 7625
rect -200 7540 -30 7560
rect -200 7510 -190 7540
rect -160 7510 -30 7540
rect -200 7470 -30 7510
rect -200 7440 -190 7470
rect -160 7440 -30 7470
rect -200 7420 -30 7440
rect 0 7540 170 7560
rect 0 7510 10 7540
rect 40 7510 170 7540
rect 0 7470 170 7510
rect 0 7440 10 7470
rect 40 7440 170 7470
rect 0 7420 170 7440
rect 200 7540 370 7560
rect 200 7510 210 7540
rect 240 7510 370 7540
rect 200 7470 370 7510
rect 200 7440 210 7470
rect 240 7440 370 7470
rect 200 7420 370 7440
rect 400 7540 570 7560
rect 400 7510 410 7540
rect 440 7510 570 7540
rect 400 7470 570 7510
rect 400 7440 410 7470
rect 440 7440 570 7470
rect 400 7420 570 7440
rect 600 7540 770 7560
rect 600 7510 610 7540
rect 640 7510 770 7540
rect 600 7470 770 7510
rect 600 7440 610 7470
rect 640 7440 770 7470
rect 600 7420 770 7440
rect 800 7540 970 7560
rect 800 7510 810 7540
rect 840 7510 970 7540
rect 800 7470 970 7510
rect 800 7440 810 7470
rect 840 7440 970 7470
rect 800 7420 970 7440
rect 1000 7540 1170 7560
rect 1000 7510 1010 7540
rect 1040 7510 1170 7540
rect 1000 7470 1170 7510
rect 1000 7440 1010 7470
rect 1040 7440 1170 7470
rect 1000 7420 1170 7440
rect 1200 7540 1370 7560
rect 1200 7510 1210 7540
rect 1240 7510 1370 7540
rect 1200 7470 1370 7510
rect 1200 7440 1210 7470
rect 1240 7440 1370 7470
rect 1200 7420 1370 7440
rect 1400 7540 1570 7560
rect 1400 7510 1410 7540
rect 1440 7510 1570 7540
rect 1400 7470 1570 7510
rect 1400 7440 1410 7470
rect 1440 7440 1570 7470
rect 1400 7420 1570 7440
rect 1600 7540 1770 7560
rect 1600 7510 1610 7540
rect 1640 7510 1770 7540
rect 1600 7470 1770 7510
rect 1600 7440 1610 7470
rect 1640 7440 1770 7470
rect 1600 7420 1770 7440
rect 1800 7540 1970 7560
rect 1800 7510 1810 7540
rect 1840 7510 1970 7540
rect 1800 7470 1970 7510
rect 1800 7440 1810 7470
rect 1840 7440 1970 7470
rect 1800 7420 1970 7440
rect 2000 7540 2170 7560
rect 2000 7510 2010 7540
rect 2040 7510 2170 7540
rect 2000 7470 2170 7510
rect 2000 7440 2010 7470
rect 2040 7440 2170 7470
rect 2000 7420 2170 7440
rect 2200 7540 2370 7560
rect 2200 7510 2210 7540
rect 2240 7510 2370 7540
rect 2200 7470 2370 7510
rect 2200 7440 2210 7470
rect 2240 7440 2370 7470
rect 2200 7420 2370 7440
rect 2400 7540 2570 7560
rect 2400 7510 2410 7540
rect 2440 7510 2570 7540
rect 2400 7470 2570 7510
rect 2400 7440 2410 7470
rect 2440 7440 2570 7470
rect 2400 7420 2570 7440
rect 2600 7540 2770 7560
rect 2600 7510 2610 7540
rect 2640 7510 2770 7540
rect 2600 7470 2770 7510
rect 2600 7440 2610 7470
rect 2640 7440 2770 7470
rect 2600 7420 2770 7440
rect 2800 7540 2970 7560
rect 2800 7510 2810 7540
rect 2840 7510 2970 7540
rect 2800 7470 2970 7510
rect 2800 7440 2810 7470
rect 2840 7440 2970 7470
rect 2800 7420 2970 7440
rect 3000 7540 3170 7560
rect 3000 7510 3010 7540
rect 3040 7510 3170 7540
rect 3000 7470 3170 7510
rect 3000 7440 3010 7470
rect 3040 7440 3170 7470
rect 3000 7420 3170 7440
rect 3200 7540 3370 7560
rect 3200 7510 3210 7540
rect 3240 7510 3370 7540
rect 3200 7470 3370 7510
rect 3200 7440 3210 7470
rect 3240 7440 3370 7470
rect 3200 7420 3370 7440
rect 3400 7540 3570 7560
rect 3400 7510 3410 7540
rect 3440 7510 3570 7540
rect 3400 7470 3570 7510
rect 3400 7440 3410 7470
rect 3440 7440 3570 7470
rect 3400 7420 3570 7440
rect 3600 7540 3770 7560
rect 3600 7510 3610 7540
rect 3640 7510 3770 7540
rect 3600 7470 3770 7510
rect 3600 7440 3610 7470
rect 3640 7440 3770 7470
rect 3600 7420 3770 7440
rect 3800 7540 3970 7560
rect 3800 7510 3810 7540
rect 3840 7510 3970 7540
rect 3800 7470 3970 7510
rect 3800 7440 3810 7470
rect 3840 7440 3970 7470
rect 3800 7420 3970 7440
rect 4000 7540 4170 7560
rect 4000 7510 4010 7540
rect 4040 7510 4170 7540
rect 4000 7470 4170 7510
rect 4000 7440 4010 7470
rect 4040 7440 4170 7470
rect 4000 7420 4170 7440
rect 4200 7540 4370 7560
rect 4200 7510 4210 7540
rect 4240 7510 4370 7540
rect 4200 7470 4370 7510
rect 4200 7440 4210 7470
rect 4240 7440 4370 7470
rect 4200 7420 4370 7440
rect 4400 7540 4570 7560
rect 4400 7510 4410 7540
rect 4440 7510 4570 7540
rect 4400 7470 4570 7510
rect 4400 7440 4410 7470
rect 4440 7440 4570 7470
rect 4400 7420 4570 7440
rect 4600 7540 4770 7560
rect 4600 7510 4610 7540
rect 4640 7510 4770 7540
rect 4600 7470 4770 7510
rect 4600 7440 4610 7470
rect 4640 7440 4770 7470
rect 4600 7420 4770 7440
rect 4800 7540 4970 7560
rect 4800 7510 4810 7540
rect 4840 7510 4970 7540
rect 4800 7470 4970 7510
rect 4800 7440 4810 7470
rect 4840 7440 4970 7470
rect 4800 7420 4970 7440
rect 5000 7540 5170 7560
rect 5000 7510 5010 7540
rect 5040 7510 5170 7540
rect 5000 7470 5170 7510
rect 5000 7440 5010 7470
rect 5040 7440 5170 7470
rect 5000 7420 5170 7440
rect 5200 7540 5370 7560
rect 5200 7510 5210 7540
rect 5240 7510 5370 7540
rect 5200 7470 5370 7510
rect 5200 7440 5210 7470
rect 5240 7440 5370 7470
rect 5200 7420 5370 7440
rect 5400 7540 5570 7560
rect 5400 7510 5410 7540
rect 5440 7510 5570 7540
rect 5400 7470 5570 7510
rect 5400 7440 5410 7470
rect 5440 7440 5570 7470
rect 5400 7420 5570 7440
rect 5600 7540 5770 7560
rect 5600 7510 5610 7540
rect 5640 7510 5770 7540
rect 5600 7470 5770 7510
rect 5600 7440 5610 7470
rect 5640 7440 5770 7470
rect 5600 7420 5770 7440
rect 5800 7540 5970 7560
rect 5800 7510 5810 7540
rect 5840 7510 5970 7540
rect 5800 7470 5970 7510
rect 5800 7440 5810 7470
rect 5840 7440 5970 7470
rect 5800 7420 5970 7440
rect 6000 7540 6170 7560
rect 6000 7510 6010 7540
rect 6040 7510 6170 7540
rect 6000 7470 6170 7510
rect 6000 7440 6010 7470
rect 6040 7440 6170 7470
rect 6000 7420 6170 7440
rect 6200 7540 6370 7560
rect 6200 7510 6210 7540
rect 6240 7510 6370 7540
rect 6200 7470 6370 7510
rect 6200 7440 6210 7470
rect 6240 7440 6370 7470
rect 6200 7420 6370 7440
rect 6400 7540 6570 7560
rect 6400 7510 6410 7540
rect 6440 7510 6570 7540
rect 6400 7470 6570 7510
rect 6400 7440 6410 7470
rect 6440 7440 6570 7470
rect 6400 7420 6570 7440
rect -200 7355 -30 7375
rect -200 7325 -190 7355
rect -160 7325 -30 7355
rect -200 7285 -30 7325
rect -200 7255 -190 7285
rect -160 7255 -30 7285
rect -200 7235 -30 7255
rect 0 7355 170 7375
rect 0 7325 10 7355
rect 40 7325 170 7355
rect 0 7285 170 7325
rect 0 7255 10 7285
rect 40 7255 170 7285
rect 0 7235 170 7255
rect 200 7355 370 7375
rect 200 7325 210 7355
rect 240 7325 370 7355
rect 200 7285 370 7325
rect 200 7255 210 7285
rect 240 7255 370 7285
rect 200 7235 370 7255
rect 400 7355 570 7375
rect 400 7325 410 7355
rect 440 7325 570 7355
rect 400 7285 570 7325
rect 400 7255 410 7285
rect 440 7255 570 7285
rect 400 7235 570 7255
rect 600 7355 770 7375
rect 600 7325 610 7355
rect 640 7325 770 7355
rect 600 7285 770 7325
rect 600 7255 610 7285
rect 640 7255 770 7285
rect 600 7235 770 7255
rect 800 7355 970 7375
rect 800 7325 810 7355
rect 840 7325 970 7355
rect 800 7285 970 7325
rect 800 7255 810 7285
rect 840 7255 970 7285
rect 800 7235 970 7255
rect 1000 7355 1170 7375
rect 1000 7325 1010 7355
rect 1040 7325 1170 7355
rect 1000 7285 1170 7325
rect 1000 7255 1010 7285
rect 1040 7255 1170 7285
rect 1000 7235 1170 7255
rect 1200 7355 1370 7375
rect 1200 7325 1210 7355
rect 1240 7325 1370 7355
rect 1200 7285 1370 7325
rect 1200 7255 1210 7285
rect 1240 7255 1370 7285
rect 1200 7235 1370 7255
rect 1400 7355 1570 7375
rect 1400 7325 1410 7355
rect 1440 7325 1570 7355
rect 1400 7285 1570 7325
rect 1400 7255 1410 7285
rect 1440 7255 1570 7285
rect 1400 7235 1570 7255
rect 1600 7355 1770 7375
rect 1600 7325 1610 7355
rect 1640 7325 1770 7355
rect 1600 7285 1770 7325
rect 1600 7255 1610 7285
rect 1640 7255 1770 7285
rect 1600 7235 1770 7255
rect 1800 7355 1970 7375
rect 1800 7325 1810 7355
rect 1840 7325 1970 7355
rect 1800 7285 1970 7325
rect 1800 7255 1810 7285
rect 1840 7255 1970 7285
rect 1800 7235 1970 7255
rect 2000 7355 2170 7375
rect 2000 7325 2010 7355
rect 2040 7325 2170 7355
rect 2000 7285 2170 7325
rect 2000 7255 2010 7285
rect 2040 7255 2170 7285
rect 2000 7235 2170 7255
rect 2200 7355 2370 7375
rect 2200 7325 2210 7355
rect 2240 7325 2370 7355
rect 2200 7285 2370 7325
rect 2200 7255 2210 7285
rect 2240 7255 2370 7285
rect 2200 7235 2370 7255
rect 2400 7355 2570 7375
rect 2400 7325 2410 7355
rect 2440 7325 2570 7355
rect 2400 7285 2570 7325
rect 2400 7255 2410 7285
rect 2440 7255 2570 7285
rect 2400 7235 2570 7255
rect 2600 7355 2770 7375
rect 2600 7325 2610 7355
rect 2640 7325 2770 7355
rect 2600 7285 2770 7325
rect 2600 7255 2610 7285
rect 2640 7255 2770 7285
rect 2600 7235 2770 7255
rect 2800 7355 2970 7375
rect 2800 7325 2810 7355
rect 2840 7325 2970 7355
rect 2800 7285 2970 7325
rect 2800 7255 2810 7285
rect 2840 7255 2970 7285
rect 2800 7235 2970 7255
rect 3000 7355 3170 7375
rect 3000 7325 3010 7355
rect 3040 7325 3170 7355
rect 3000 7285 3170 7325
rect 3000 7255 3010 7285
rect 3040 7255 3170 7285
rect 3000 7235 3170 7255
rect 3200 7355 3370 7375
rect 3200 7325 3210 7355
rect 3240 7325 3370 7355
rect 3200 7285 3370 7325
rect 3200 7255 3210 7285
rect 3240 7255 3370 7285
rect 3200 7235 3370 7255
rect 3400 7355 3570 7375
rect 3400 7325 3410 7355
rect 3440 7325 3570 7355
rect 3400 7285 3570 7325
rect 3400 7255 3410 7285
rect 3440 7255 3570 7285
rect 3400 7235 3570 7255
rect 3600 7355 3770 7375
rect 3600 7325 3610 7355
rect 3640 7325 3770 7355
rect 3600 7285 3770 7325
rect 3600 7255 3610 7285
rect 3640 7255 3770 7285
rect 3600 7235 3770 7255
rect 3800 7355 3970 7375
rect 3800 7325 3810 7355
rect 3840 7325 3970 7355
rect 3800 7285 3970 7325
rect 3800 7255 3810 7285
rect 3840 7255 3970 7285
rect 3800 7235 3970 7255
rect 4000 7355 4170 7375
rect 4000 7325 4010 7355
rect 4040 7325 4170 7355
rect 4000 7285 4170 7325
rect 4000 7255 4010 7285
rect 4040 7255 4170 7285
rect 4000 7235 4170 7255
rect 4200 7355 4370 7375
rect 4200 7325 4210 7355
rect 4240 7325 4370 7355
rect 4200 7285 4370 7325
rect 4200 7255 4210 7285
rect 4240 7255 4370 7285
rect 4200 7235 4370 7255
rect 4400 7355 4570 7375
rect 4400 7325 4410 7355
rect 4440 7325 4570 7355
rect 4400 7285 4570 7325
rect 4400 7255 4410 7285
rect 4440 7255 4570 7285
rect 4400 7235 4570 7255
rect 4600 7355 4770 7375
rect 4600 7325 4610 7355
rect 4640 7325 4770 7355
rect 4600 7285 4770 7325
rect 4600 7255 4610 7285
rect 4640 7255 4770 7285
rect 4600 7235 4770 7255
rect 4800 7355 4970 7375
rect 4800 7325 4810 7355
rect 4840 7325 4970 7355
rect 4800 7285 4970 7325
rect 4800 7255 4810 7285
rect 4840 7255 4970 7285
rect 4800 7235 4970 7255
rect 5000 7355 5170 7375
rect 5000 7325 5010 7355
rect 5040 7325 5170 7355
rect 5000 7285 5170 7325
rect 5000 7255 5010 7285
rect 5040 7255 5170 7285
rect 5000 7235 5170 7255
rect 5200 7355 5370 7375
rect 5200 7325 5210 7355
rect 5240 7325 5370 7355
rect 5200 7285 5370 7325
rect 5200 7255 5210 7285
rect 5240 7255 5370 7285
rect 5200 7235 5370 7255
rect 5400 7355 5570 7375
rect 5400 7325 5410 7355
rect 5440 7325 5570 7355
rect 5400 7285 5570 7325
rect 5400 7255 5410 7285
rect 5440 7255 5570 7285
rect 5400 7235 5570 7255
rect 5600 7355 5770 7375
rect 5600 7325 5610 7355
rect 5640 7325 5770 7355
rect 5600 7285 5770 7325
rect 5600 7255 5610 7285
rect 5640 7255 5770 7285
rect 5600 7235 5770 7255
rect 5800 7355 5970 7375
rect 5800 7325 5810 7355
rect 5840 7325 5970 7355
rect 5800 7285 5970 7325
rect 5800 7255 5810 7285
rect 5840 7255 5970 7285
rect 5800 7235 5970 7255
rect 6000 7355 6170 7375
rect 6000 7325 6010 7355
rect 6040 7325 6170 7355
rect 6000 7285 6170 7325
rect 6000 7255 6010 7285
rect 6040 7255 6170 7285
rect 6000 7235 6170 7255
rect 6200 7355 6370 7375
rect 6200 7325 6210 7355
rect 6240 7325 6370 7355
rect 6200 7285 6370 7325
rect 6200 7255 6210 7285
rect 6240 7255 6370 7285
rect 6200 7235 6370 7255
rect 6400 7355 6570 7375
rect 6400 7325 6410 7355
rect 6440 7325 6570 7355
rect 6400 7285 6570 7325
rect 6400 7255 6410 7285
rect 6440 7255 6570 7285
rect 6400 7235 6570 7255
rect -200 7170 -30 7190
rect -200 7140 -190 7170
rect -160 7140 -30 7170
rect -200 7100 -30 7140
rect -200 7070 -190 7100
rect -160 7070 -30 7100
rect -200 7050 -30 7070
rect 0 7170 170 7190
rect 0 7140 10 7170
rect 40 7140 170 7170
rect 0 7100 170 7140
rect 0 7070 10 7100
rect 40 7070 170 7100
rect 0 7050 170 7070
rect 200 7170 370 7190
rect 200 7140 210 7170
rect 240 7140 370 7170
rect 200 7100 370 7140
rect 200 7070 210 7100
rect 240 7070 370 7100
rect 200 7050 370 7070
rect 400 7170 570 7190
rect 400 7140 410 7170
rect 440 7140 570 7170
rect 400 7100 570 7140
rect 400 7070 410 7100
rect 440 7070 570 7100
rect 400 7050 570 7070
rect 600 7170 770 7190
rect 600 7140 610 7170
rect 640 7140 770 7170
rect 600 7100 770 7140
rect 600 7070 610 7100
rect 640 7070 770 7100
rect 600 7050 770 7070
rect 800 7170 970 7190
rect 800 7140 810 7170
rect 840 7140 970 7170
rect 800 7100 970 7140
rect 800 7070 810 7100
rect 840 7070 970 7100
rect 800 7050 970 7070
rect 1000 7170 1170 7190
rect 1000 7140 1010 7170
rect 1040 7140 1170 7170
rect 1000 7100 1170 7140
rect 1000 7070 1010 7100
rect 1040 7070 1170 7100
rect 1000 7050 1170 7070
rect 1200 7170 1370 7190
rect 1200 7140 1210 7170
rect 1240 7140 1370 7170
rect 1200 7100 1370 7140
rect 1200 7070 1210 7100
rect 1240 7070 1370 7100
rect 1200 7050 1370 7070
rect 1400 7170 1570 7190
rect 1400 7140 1410 7170
rect 1440 7140 1570 7170
rect 1400 7100 1570 7140
rect 1400 7070 1410 7100
rect 1440 7070 1570 7100
rect 1400 7050 1570 7070
rect 1600 7170 1770 7190
rect 1600 7140 1610 7170
rect 1640 7140 1770 7170
rect 1600 7100 1770 7140
rect 1600 7070 1610 7100
rect 1640 7070 1770 7100
rect 1600 7050 1770 7070
rect 1800 7170 1970 7190
rect 1800 7140 1810 7170
rect 1840 7140 1970 7170
rect 1800 7100 1970 7140
rect 1800 7070 1810 7100
rect 1840 7070 1970 7100
rect 1800 7050 1970 7070
rect 2000 7170 2170 7190
rect 2000 7140 2010 7170
rect 2040 7140 2170 7170
rect 2000 7100 2170 7140
rect 2000 7070 2010 7100
rect 2040 7070 2170 7100
rect 2000 7050 2170 7070
rect 2200 7170 2370 7190
rect 2200 7140 2210 7170
rect 2240 7140 2370 7170
rect 2200 7100 2370 7140
rect 2200 7070 2210 7100
rect 2240 7070 2370 7100
rect 2200 7050 2370 7070
rect 2400 7170 2570 7190
rect 2400 7140 2410 7170
rect 2440 7140 2570 7170
rect 2400 7100 2570 7140
rect 2400 7070 2410 7100
rect 2440 7070 2570 7100
rect 2400 7050 2570 7070
rect 2600 7170 2770 7190
rect 2600 7140 2610 7170
rect 2640 7140 2770 7170
rect 2600 7100 2770 7140
rect 2600 7070 2610 7100
rect 2640 7070 2770 7100
rect 2600 7050 2770 7070
rect 2800 7170 2970 7190
rect 2800 7140 2810 7170
rect 2840 7140 2970 7170
rect 2800 7100 2970 7140
rect 2800 7070 2810 7100
rect 2840 7070 2970 7100
rect 2800 7050 2970 7070
rect 3000 7170 3170 7190
rect 3000 7140 3010 7170
rect 3040 7140 3170 7170
rect 3000 7100 3170 7140
rect 3000 7070 3010 7100
rect 3040 7070 3170 7100
rect 3000 7050 3170 7070
rect 3200 7170 3370 7190
rect 3200 7140 3210 7170
rect 3240 7140 3370 7170
rect 3200 7100 3370 7140
rect 3200 7070 3210 7100
rect 3240 7070 3370 7100
rect 3200 7050 3370 7070
rect 3400 7170 3570 7190
rect 3400 7140 3410 7170
rect 3440 7140 3570 7170
rect 3400 7100 3570 7140
rect 3400 7070 3410 7100
rect 3440 7070 3570 7100
rect 3400 7050 3570 7070
rect 3600 7170 3770 7190
rect 3600 7140 3610 7170
rect 3640 7140 3770 7170
rect 3600 7100 3770 7140
rect 3600 7070 3610 7100
rect 3640 7070 3770 7100
rect 3600 7050 3770 7070
rect 3800 7170 3970 7190
rect 3800 7140 3810 7170
rect 3840 7140 3970 7170
rect 3800 7100 3970 7140
rect 3800 7070 3810 7100
rect 3840 7070 3970 7100
rect 3800 7050 3970 7070
rect 4000 7170 4170 7190
rect 4000 7140 4010 7170
rect 4040 7140 4170 7170
rect 4000 7100 4170 7140
rect 4000 7070 4010 7100
rect 4040 7070 4170 7100
rect 4000 7050 4170 7070
rect 4200 7170 4370 7190
rect 4200 7140 4210 7170
rect 4240 7140 4370 7170
rect 4200 7100 4370 7140
rect 4200 7070 4210 7100
rect 4240 7070 4370 7100
rect 4200 7050 4370 7070
rect 4400 7170 4570 7190
rect 4400 7140 4410 7170
rect 4440 7140 4570 7170
rect 4400 7100 4570 7140
rect 4400 7070 4410 7100
rect 4440 7070 4570 7100
rect 4400 7050 4570 7070
rect 4600 7170 4770 7190
rect 4600 7140 4610 7170
rect 4640 7140 4770 7170
rect 4600 7100 4770 7140
rect 4600 7070 4610 7100
rect 4640 7070 4770 7100
rect 4600 7050 4770 7070
rect 4800 7170 4970 7190
rect 4800 7140 4810 7170
rect 4840 7140 4970 7170
rect 4800 7100 4970 7140
rect 4800 7070 4810 7100
rect 4840 7070 4970 7100
rect 4800 7050 4970 7070
rect 5000 7170 5170 7190
rect 5000 7140 5010 7170
rect 5040 7140 5170 7170
rect 5000 7100 5170 7140
rect 5000 7070 5010 7100
rect 5040 7070 5170 7100
rect 5000 7050 5170 7070
rect 5200 7170 5370 7190
rect 5200 7140 5210 7170
rect 5240 7140 5370 7170
rect 5200 7100 5370 7140
rect 5200 7070 5210 7100
rect 5240 7070 5370 7100
rect 5200 7050 5370 7070
rect 5400 7170 5570 7190
rect 5400 7140 5410 7170
rect 5440 7140 5570 7170
rect 5400 7100 5570 7140
rect 5400 7070 5410 7100
rect 5440 7070 5570 7100
rect 5400 7050 5570 7070
rect 5600 7170 5770 7190
rect 5600 7140 5610 7170
rect 5640 7140 5770 7170
rect 5600 7100 5770 7140
rect 5600 7070 5610 7100
rect 5640 7070 5770 7100
rect 5600 7050 5770 7070
rect 5800 7170 5970 7190
rect 5800 7140 5810 7170
rect 5840 7140 5970 7170
rect 5800 7100 5970 7140
rect 5800 7070 5810 7100
rect 5840 7070 5970 7100
rect 5800 7050 5970 7070
rect 6000 7170 6170 7190
rect 6000 7140 6010 7170
rect 6040 7140 6170 7170
rect 6000 7100 6170 7140
rect 6000 7070 6010 7100
rect 6040 7070 6170 7100
rect 6000 7050 6170 7070
rect 6200 7170 6370 7190
rect 6200 7140 6210 7170
rect 6240 7140 6370 7170
rect 6200 7100 6370 7140
rect 6200 7070 6210 7100
rect 6240 7070 6370 7100
rect 6200 7050 6370 7070
rect 6400 7170 6570 7190
rect 6400 7140 6410 7170
rect 6440 7140 6570 7170
rect 6400 7100 6570 7140
rect 6400 7070 6410 7100
rect 6440 7070 6570 7100
rect 6400 7050 6570 7070
rect -200 6985 -30 7005
rect -200 6955 -190 6985
rect -160 6955 -30 6985
rect -200 6915 -30 6955
rect -200 6885 -190 6915
rect -160 6885 -30 6915
rect -200 6865 -30 6885
rect 0 6985 170 7005
rect 0 6955 10 6985
rect 40 6955 170 6985
rect 0 6915 170 6955
rect 0 6885 10 6915
rect 40 6885 170 6915
rect 0 6865 170 6885
rect 200 6985 370 7005
rect 200 6955 210 6985
rect 240 6955 370 6985
rect 200 6915 370 6955
rect 200 6885 210 6915
rect 240 6885 370 6915
rect 200 6865 370 6885
rect 400 6985 570 7005
rect 400 6955 410 6985
rect 440 6955 570 6985
rect 400 6915 570 6955
rect 400 6885 410 6915
rect 440 6885 570 6915
rect 400 6865 570 6885
rect 600 6985 770 7005
rect 600 6955 610 6985
rect 640 6955 770 6985
rect 600 6915 770 6955
rect 600 6885 610 6915
rect 640 6885 770 6915
rect 600 6865 770 6885
rect 800 6985 970 7005
rect 800 6955 810 6985
rect 840 6955 970 6985
rect 800 6915 970 6955
rect 800 6885 810 6915
rect 840 6885 970 6915
rect 800 6865 970 6885
rect 1000 6985 1170 7005
rect 1000 6955 1010 6985
rect 1040 6955 1170 6985
rect 1000 6915 1170 6955
rect 1000 6885 1010 6915
rect 1040 6885 1170 6915
rect 1000 6865 1170 6885
rect 1200 6985 1370 7005
rect 1200 6955 1210 6985
rect 1240 6955 1370 6985
rect 1200 6915 1370 6955
rect 1200 6885 1210 6915
rect 1240 6885 1370 6915
rect 1200 6865 1370 6885
rect 1400 6985 1570 7005
rect 1400 6955 1410 6985
rect 1440 6955 1570 6985
rect 1400 6915 1570 6955
rect 1400 6885 1410 6915
rect 1440 6885 1570 6915
rect 1400 6865 1570 6885
rect 1600 6985 1770 7005
rect 1600 6955 1610 6985
rect 1640 6955 1770 6985
rect 1600 6915 1770 6955
rect 1600 6885 1610 6915
rect 1640 6885 1770 6915
rect 1600 6865 1770 6885
rect 1800 6985 1970 7005
rect 1800 6955 1810 6985
rect 1840 6955 1970 6985
rect 1800 6915 1970 6955
rect 1800 6885 1810 6915
rect 1840 6885 1970 6915
rect 1800 6865 1970 6885
rect 2000 6985 2170 7005
rect 2000 6955 2010 6985
rect 2040 6955 2170 6985
rect 2000 6915 2170 6955
rect 2000 6885 2010 6915
rect 2040 6885 2170 6915
rect 2000 6865 2170 6885
rect 2200 6985 2370 7005
rect 2200 6955 2210 6985
rect 2240 6955 2370 6985
rect 2200 6915 2370 6955
rect 2200 6885 2210 6915
rect 2240 6885 2370 6915
rect 2200 6865 2370 6885
rect 2400 6985 2570 7005
rect 2400 6955 2410 6985
rect 2440 6955 2570 6985
rect 2400 6915 2570 6955
rect 2400 6885 2410 6915
rect 2440 6885 2570 6915
rect 2400 6865 2570 6885
rect 2600 6985 2770 7005
rect 2600 6955 2610 6985
rect 2640 6955 2770 6985
rect 2600 6915 2770 6955
rect 2600 6885 2610 6915
rect 2640 6885 2770 6915
rect 2600 6865 2770 6885
rect 2800 6985 2970 7005
rect 2800 6955 2810 6985
rect 2840 6955 2970 6985
rect 2800 6915 2970 6955
rect 2800 6885 2810 6915
rect 2840 6885 2970 6915
rect 2800 6865 2970 6885
rect 3000 6985 3170 7005
rect 3000 6955 3010 6985
rect 3040 6955 3170 6985
rect 3000 6915 3170 6955
rect 3000 6885 3010 6915
rect 3040 6885 3170 6915
rect 3000 6865 3170 6885
rect 3200 6985 3370 7005
rect 3200 6955 3210 6985
rect 3240 6955 3370 6985
rect 3200 6915 3370 6955
rect 3200 6885 3210 6915
rect 3240 6885 3370 6915
rect 3200 6865 3370 6885
rect 3400 6985 3570 7005
rect 3400 6955 3410 6985
rect 3440 6955 3570 6985
rect 3400 6915 3570 6955
rect 3400 6885 3410 6915
rect 3440 6885 3570 6915
rect 3400 6865 3570 6885
rect 3600 6985 3770 7005
rect 3600 6955 3610 6985
rect 3640 6955 3770 6985
rect 3600 6915 3770 6955
rect 3600 6885 3610 6915
rect 3640 6885 3770 6915
rect 3600 6865 3770 6885
rect 3800 6985 3970 7005
rect 3800 6955 3810 6985
rect 3840 6955 3970 6985
rect 3800 6915 3970 6955
rect 3800 6885 3810 6915
rect 3840 6885 3970 6915
rect 3800 6865 3970 6885
rect 4000 6985 4170 7005
rect 4000 6955 4010 6985
rect 4040 6955 4170 6985
rect 4000 6915 4170 6955
rect 4000 6885 4010 6915
rect 4040 6885 4170 6915
rect 4000 6865 4170 6885
rect 4200 6985 4370 7005
rect 4200 6955 4210 6985
rect 4240 6955 4370 6985
rect 4200 6915 4370 6955
rect 4200 6885 4210 6915
rect 4240 6885 4370 6915
rect 4200 6865 4370 6885
rect 4400 6985 4570 7005
rect 4400 6955 4410 6985
rect 4440 6955 4570 6985
rect 4400 6915 4570 6955
rect 4400 6885 4410 6915
rect 4440 6885 4570 6915
rect 4400 6865 4570 6885
rect 4600 6985 4770 7005
rect 4600 6955 4610 6985
rect 4640 6955 4770 6985
rect 4600 6915 4770 6955
rect 4600 6885 4610 6915
rect 4640 6885 4770 6915
rect 4600 6865 4770 6885
rect 4800 6985 4970 7005
rect 4800 6955 4810 6985
rect 4840 6955 4970 6985
rect 4800 6915 4970 6955
rect 4800 6885 4810 6915
rect 4840 6885 4970 6915
rect 4800 6865 4970 6885
rect 5000 6985 5170 7005
rect 5000 6955 5010 6985
rect 5040 6955 5170 6985
rect 5000 6915 5170 6955
rect 5000 6885 5010 6915
rect 5040 6885 5170 6915
rect 5000 6865 5170 6885
rect 5200 6985 5370 7005
rect 5200 6955 5210 6985
rect 5240 6955 5370 6985
rect 5200 6915 5370 6955
rect 5200 6885 5210 6915
rect 5240 6885 5370 6915
rect 5200 6865 5370 6885
rect 5400 6985 5570 7005
rect 5400 6955 5410 6985
rect 5440 6955 5570 6985
rect 5400 6915 5570 6955
rect 5400 6885 5410 6915
rect 5440 6885 5570 6915
rect 5400 6865 5570 6885
rect 5600 6985 5770 7005
rect 5600 6955 5610 6985
rect 5640 6955 5770 6985
rect 5600 6915 5770 6955
rect 5600 6885 5610 6915
rect 5640 6885 5770 6915
rect 5600 6865 5770 6885
rect 5800 6985 5970 7005
rect 5800 6955 5810 6985
rect 5840 6955 5970 6985
rect 5800 6915 5970 6955
rect 5800 6885 5810 6915
rect 5840 6885 5970 6915
rect 5800 6865 5970 6885
rect 6000 6985 6170 7005
rect 6000 6955 6010 6985
rect 6040 6955 6170 6985
rect 6000 6915 6170 6955
rect 6000 6885 6010 6915
rect 6040 6885 6170 6915
rect 6000 6865 6170 6885
rect 6200 6985 6370 7005
rect 6200 6955 6210 6985
rect 6240 6955 6370 6985
rect 6200 6915 6370 6955
rect 6200 6885 6210 6915
rect 6240 6885 6370 6915
rect 6200 6865 6370 6885
rect 6400 6985 6570 7005
rect 6400 6955 6410 6985
rect 6440 6955 6570 6985
rect 6400 6915 6570 6955
rect 6400 6885 6410 6915
rect 6440 6885 6570 6915
rect 6400 6865 6570 6885
rect -200 6800 -30 6820
rect -200 6770 -190 6800
rect -160 6770 -30 6800
rect -200 6730 -30 6770
rect -200 6700 -190 6730
rect -160 6700 -30 6730
rect -200 6680 -30 6700
rect 0 6800 170 6820
rect 0 6770 10 6800
rect 40 6770 170 6800
rect 0 6730 170 6770
rect 0 6700 10 6730
rect 40 6700 170 6730
rect 0 6680 170 6700
rect 200 6800 370 6820
rect 200 6770 210 6800
rect 240 6770 370 6800
rect 200 6730 370 6770
rect 200 6700 210 6730
rect 240 6700 370 6730
rect 200 6680 370 6700
rect 400 6800 570 6820
rect 400 6770 410 6800
rect 440 6770 570 6800
rect 400 6730 570 6770
rect 400 6700 410 6730
rect 440 6700 570 6730
rect 400 6680 570 6700
rect 600 6800 770 6820
rect 600 6770 610 6800
rect 640 6770 770 6800
rect 600 6730 770 6770
rect 600 6700 610 6730
rect 640 6700 770 6730
rect 600 6680 770 6700
rect 800 6800 970 6820
rect 800 6770 810 6800
rect 840 6770 970 6800
rect 800 6730 970 6770
rect 800 6700 810 6730
rect 840 6700 970 6730
rect 800 6680 970 6700
rect 1000 6800 1170 6820
rect 1000 6770 1010 6800
rect 1040 6770 1170 6800
rect 1000 6730 1170 6770
rect 1000 6700 1010 6730
rect 1040 6700 1170 6730
rect 1000 6680 1170 6700
rect 1200 6800 1370 6820
rect 1200 6770 1210 6800
rect 1240 6770 1370 6800
rect 1200 6730 1370 6770
rect 1200 6700 1210 6730
rect 1240 6700 1370 6730
rect 1200 6680 1370 6700
rect 1400 6800 1570 6820
rect 1400 6770 1410 6800
rect 1440 6770 1570 6800
rect 1400 6730 1570 6770
rect 1400 6700 1410 6730
rect 1440 6700 1570 6730
rect 1400 6680 1570 6700
rect 1600 6800 1770 6820
rect 1600 6770 1610 6800
rect 1640 6770 1770 6800
rect 1600 6730 1770 6770
rect 1600 6700 1610 6730
rect 1640 6700 1770 6730
rect 1600 6680 1770 6700
rect 1800 6800 1970 6820
rect 1800 6770 1810 6800
rect 1840 6770 1970 6800
rect 1800 6730 1970 6770
rect 1800 6700 1810 6730
rect 1840 6700 1970 6730
rect 1800 6680 1970 6700
rect 2000 6800 2170 6820
rect 2000 6770 2010 6800
rect 2040 6770 2170 6800
rect 2000 6730 2170 6770
rect 2000 6700 2010 6730
rect 2040 6700 2170 6730
rect 2000 6680 2170 6700
rect 2200 6800 2370 6820
rect 2200 6770 2210 6800
rect 2240 6770 2370 6800
rect 2200 6730 2370 6770
rect 2200 6700 2210 6730
rect 2240 6700 2370 6730
rect 2200 6680 2370 6700
rect 2400 6800 2570 6820
rect 2400 6770 2410 6800
rect 2440 6770 2570 6800
rect 2400 6730 2570 6770
rect 2400 6700 2410 6730
rect 2440 6700 2570 6730
rect 2400 6680 2570 6700
rect 2600 6800 2770 6820
rect 2600 6770 2610 6800
rect 2640 6770 2770 6800
rect 2600 6730 2770 6770
rect 2600 6700 2610 6730
rect 2640 6700 2770 6730
rect 2600 6680 2770 6700
rect 2800 6800 2970 6820
rect 2800 6770 2810 6800
rect 2840 6770 2970 6800
rect 2800 6730 2970 6770
rect 2800 6700 2810 6730
rect 2840 6700 2970 6730
rect 2800 6680 2970 6700
rect 3000 6800 3170 6820
rect 3000 6770 3010 6800
rect 3040 6770 3170 6800
rect 3000 6730 3170 6770
rect 3000 6700 3010 6730
rect 3040 6700 3170 6730
rect 3000 6680 3170 6700
rect 3200 6800 3370 6820
rect 3200 6770 3210 6800
rect 3240 6770 3370 6800
rect 3200 6730 3370 6770
rect 3200 6700 3210 6730
rect 3240 6700 3370 6730
rect 3200 6680 3370 6700
rect 3400 6800 3570 6820
rect 3400 6770 3410 6800
rect 3440 6770 3570 6800
rect 3400 6730 3570 6770
rect 3400 6700 3410 6730
rect 3440 6700 3570 6730
rect 3400 6680 3570 6700
rect 3600 6800 3770 6820
rect 3600 6770 3610 6800
rect 3640 6770 3770 6800
rect 3600 6730 3770 6770
rect 3600 6700 3610 6730
rect 3640 6700 3770 6730
rect 3600 6680 3770 6700
rect 3800 6800 3970 6820
rect 3800 6770 3810 6800
rect 3840 6770 3970 6800
rect 3800 6730 3970 6770
rect 3800 6700 3810 6730
rect 3840 6700 3970 6730
rect 3800 6680 3970 6700
rect 4000 6800 4170 6820
rect 4000 6770 4010 6800
rect 4040 6770 4170 6800
rect 4000 6730 4170 6770
rect 4000 6700 4010 6730
rect 4040 6700 4170 6730
rect 4000 6680 4170 6700
rect 4200 6800 4370 6820
rect 4200 6770 4210 6800
rect 4240 6770 4370 6800
rect 4200 6730 4370 6770
rect 4200 6700 4210 6730
rect 4240 6700 4370 6730
rect 4200 6680 4370 6700
rect 4400 6800 4570 6820
rect 4400 6770 4410 6800
rect 4440 6770 4570 6800
rect 4400 6730 4570 6770
rect 4400 6700 4410 6730
rect 4440 6700 4570 6730
rect 4400 6680 4570 6700
rect 4600 6800 4770 6820
rect 4600 6770 4610 6800
rect 4640 6770 4770 6800
rect 4600 6730 4770 6770
rect 4600 6700 4610 6730
rect 4640 6700 4770 6730
rect 4600 6680 4770 6700
rect 4800 6800 4970 6820
rect 4800 6770 4810 6800
rect 4840 6770 4970 6800
rect 4800 6730 4970 6770
rect 4800 6700 4810 6730
rect 4840 6700 4970 6730
rect 4800 6680 4970 6700
rect 5000 6800 5170 6820
rect 5000 6770 5010 6800
rect 5040 6770 5170 6800
rect 5000 6730 5170 6770
rect 5000 6700 5010 6730
rect 5040 6700 5170 6730
rect 5000 6680 5170 6700
rect 5200 6800 5370 6820
rect 5200 6770 5210 6800
rect 5240 6770 5370 6800
rect 5200 6730 5370 6770
rect 5200 6700 5210 6730
rect 5240 6700 5370 6730
rect 5200 6680 5370 6700
rect 5400 6800 5570 6820
rect 5400 6770 5410 6800
rect 5440 6770 5570 6800
rect 5400 6730 5570 6770
rect 5400 6700 5410 6730
rect 5440 6700 5570 6730
rect 5400 6680 5570 6700
rect 5600 6800 5770 6820
rect 5600 6770 5610 6800
rect 5640 6770 5770 6800
rect 5600 6730 5770 6770
rect 5600 6700 5610 6730
rect 5640 6700 5770 6730
rect 5600 6680 5770 6700
rect 5800 6800 5970 6820
rect 5800 6770 5810 6800
rect 5840 6770 5970 6800
rect 5800 6730 5970 6770
rect 5800 6700 5810 6730
rect 5840 6700 5970 6730
rect 5800 6680 5970 6700
rect 6000 6800 6170 6820
rect 6000 6770 6010 6800
rect 6040 6770 6170 6800
rect 6000 6730 6170 6770
rect 6000 6700 6010 6730
rect 6040 6700 6170 6730
rect 6000 6680 6170 6700
rect 6200 6800 6370 6820
rect 6200 6770 6210 6800
rect 6240 6770 6370 6800
rect 6200 6730 6370 6770
rect 6200 6700 6210 6730
rect 6240 6700 6370 6730
rect 6200 6680 6370 6700
rect 6400 6800 6570 6820
rect 6400 6770 6410 6800
rect 6440 6770 6570 6800
rect 6400 6730 6570 6770
rect 6400 6700 6410 6730
rect 6440 6700 6570 6730
rect 6400 6680 6570 6700
rect -200 6615 -30 6635
rect -200 6585 -190 6615
rect -160 6585 -30 6615
rect -200 6545 -30 6585
rect -200 6515 -190 6545
rect -160 6515 -30 6545
rect -200 6495 -30 6515
rect 0 6615 170 6635
rect 0 6585 10 6615
rect 40 6585 170 6615
rect 0 6545 170 6585
rect 0 6515 10 6545
rect 40 6515 170 6545
rect 0 6495 170 6515
rect 200 6615 370 6635
rect 200 6585 210 6615
rect 240 6585 370 6615
rect 200 6545 370 6585
rect 200 6515 210 6545
rect 240 6515 370 6545
rect 200 6495 370 6515
rect 400 6615 570 6635
rect 400 6585 410 6615
rect 440 6585 570 6615
rect 400 6545 570 6585
rect 400 6515 410 6545
rect 440 6515 570 6545
rect 400 6495 570 6515
rect 600 6615 770 6635
rect 600 6585 610 6615
rect 640 6585 770 6615
rect 600 6545 770 6585
rect 600 6515 610 6545
rect 640 6515 770 6545
rect 600 6495 770 6515
rect 800 6615 970 6635
rect 800 6585 810 6615
rect 840 6585 970 6615
rect 800 6545 970 6585
rect 800 6515 810 6545
rect 840 6515 970 6545
rect 800 6495 970 6515
rect 1000 6615 1170 6635
rect 1000 6585 1010 6615
rect 1040 6585 1170 6615
rect 1000 6545 1170 6585
rect 1000 6515 1010 6545
rect 1040 6515 1170 6545
rect 1000 6495 1170 6515
rect 1200 6615 1370 6635
rect 1200 6585 1210 6615
rect 1240 6585 1370 6615
rect 1200 6545 1370 6585
rect 1200 6515 1210 6545
rect 1240 6515 1370 6545
rect 1200 6495 1370 6515
rect 1400 6615 1570 6635
rect 1400 6585 1410 6615
rect 1440 6585 1570 6615
rect 1400 6545 1570 6585
rect 1400 6515 1410 6545
rect 1440 6515 1570 6545
rect 1400 6495 1570 6515
rect 1600 6615 1770 6635
rect 1600 6585 1610 6615
rect 1640 6585 1770 6615
rect 1600 6545 1770 6585
rect 1600 6515 1610 6545
rect 1640 6515 1770 6545
rect 1600 6495 1770 6515
rect 1800 6615 1970 6635
rect 1800 6585 1810 6615
rect 1840 6585 1970 6615
rect 1800 6545 1970 6585
rect 1800 6515 1810 6545
rect 1840 6515 1970 6545
rect 1800 6495 1970 6515
rect 2000 6615 2170 6635
rect 2000 6585 2010 6615
rect 2040 6585 2170 6615
rect 2000 6545 2170 6585
rect 2000 6515 2010 6545
rect 2040 6515 2170 6545
rect 2000 6495 2170 6515
rect 2200 6615 2370 6635
rect 2200 6585 2210 6615
rect 2240 6585 2370 6615
rect 2200 6545 2370 6585
rect 2200 6515 2210 6545
rect 2240 6515 2370 6545
rect 2200 6495 2370 6515
rect 2400 6615 2570 6635
rect 2400 6585 2410 6615
rect 2440 6585 2570 6615
rect 2400 6545 2570 6585
rect 2400 6515 2410 6545
rect 2440 6515 2570 6545
rect 2400 6495 2570 6515
rect 2600 6615 2770 6635
rect 2600 6585 2610 6615
rect 2640 6585 2770 6615
rect 2600 6545 2770 6585
rect 2600 6515 2610 6545
rect 2640 6515 2770 6545
rect 2600 6495 2770 6515
rect 2800 6615 2970 6635
rect 2800 6585 2810 6615
rect 2840 6585 2970 6615
rect 2800 6545 2970 6585
rect 2800 6515 2810 6545
rect 2840 6515 2970 6545
rect 2800 6495 2970 6515
rect 3000 6615 3170 6635
rect 3000 6585 3010 6615
rect 3040 6585 3170 6615
rect 3000 6545 3170 6585
rect 3000 6515 3010 6545
rect 3040 6515 3170 6545
rect 3000 6495 3170 6515
rect 3200 6615 3370 6635
rect 3200 6585 3210 6615
rect 3240 6585 3370 6615
rect 3200 6545 3370 6585
rect 3200 6515 3210 6545
rect 3240 6515 3370 6545
rect 3200 6495 3370 6515
rect 3400 6615 3570 6635
rect 3400 6585 3410 6615
rect 3440 6585 3570 6615
rect 3400 6545 3570 6585
rect 3400 6515 3410 6545
rect 3440 6515 3570 6545
rect 3400 6495 3570 6515
rect 3600 6615 3770 6635
rect 3600 6585 3610 6615
rect 3640 6585 3770 6615
rect 3600 6545 3770 6585
rect 3600 6515 3610 6545
rect 3640 6515 3770 6545
rect 3600 6495 3770 6515
rect 3800 6615 3970 6635
rect 3800 6585 3810 6615
rect 3840 6585 3970 6615
rect 3800 6545 3970 6585
rect 3800 6515 3810 6545
rect 3840 6515 3970 6545
rect 3800 6495 3970 6515
rect 4000 6615 4170 6635
rect 4000 6585 4010 6615
rect 4040 6585 4170 6615
rect 4000 6545 4170 6585
rect 4000 6515 4010 6545
rect 4040 6515 4170 6545
rect 4000 6495 4170 6515
rect 4200 6615 4370 6635
rect 4200 6585 4210 6615
rect 4240 6585 4370 6615
rect 4200 6545 4370 6585
rect 4200 6515 4210 6545
rect 4240 6515 4370 6545
rect 4200 6495 4370 6515
rect 4400 6615 4570 6635
rect 4400 6585 4410 6615
rect 4440 6585 4570 6615
rect 4400 6545 4570 6585
rect 4400 6515 4410 6545
rect 4440 6515 4570 6545
rect 4400 6495 4570 6515
rect 4600 6615 4770 6635
rect 4600 6585 4610 6615
rect 4640 6585 4770 6615
rect 4600 6545 4770 6585
rect 4600 6515 4610 6545
rect 4640 6515 4770 6545
rect 4600 6495 4770 6515
rect 4800 6615 4970 6635
rect 4800 6585 4810 6615
rect 4840 6585 4970 6615
rect 4800 6545 4970 6585
rect 4800 6515 4810 6545
rect 4840 6515 4970 6545
rect 4800 6495 4970 6515
rect 5000 6615 5170 6635
rect 5000 6585 5010 6615
rect 5040 6585 5170 6615
rect 5000 6545 5170 6585
rect 5000 6515 5010 6545
rect 5040 6515 5170 6545
rect 5000 6495 5170 6515
rect 5200 6615 5370 6635
rect 5200 6585 5210 6615
rect 5240 6585 5370 6615
rect 5200 6545 5370 6585
rect 5200 6515 5210 6545
rect 5240 6515 5370 6545
rect 5200 6495 5370 6515
rect 5400 6615 5570 6635
rect 5400 6585 5410 6615
rect 5440 6585 5570 6615
rect 5400 6545 5570 6585
rect 5400 6515 5410 6545
rect 5440 6515 5570 6545
rect 5400 6495 5570 6515
rect 5600 6615 5770 6635
rect 5600 6585 5610 6615
rect 5640 6585 5770 6615
rect 5600 6545 5770 6585
rect 5600 6515 5610 6545
rect 5640 6515 5770 6545
rect 5600 6495 5770 6515
rect 5800 6615 5970 6635
rect 5800 6585 5810 6615
rect 5840 6585 5970 6615
rect 5800 6545 5970 6585
rect 5800 6515 5810 6545
rect 5840 6515 5970 6545
rect 5800 6495 5970 6515
rect 6000 6615 6170 6635
rect 6000 6585 6010 6615
rect 6040 6585 6170 6615
rect 6000 6545 6170 6585
rect 6000 6515 6010 6545
rect 6040 6515 6170 6545
rect 6000 6495 6170 6515
rect 6200 6615 6370 6635
rect 6200 6585 6210 6615
rect 6240 6585 6370 6615
rect 6200 6545 6370 6585
rect 6200 6515 6210 6545
rect 6240 6515 6370 6545
rect 6200 6495 6370 6515
rect 6400 6615 6570 6635
rect 6400 6585 6410 6615
rect 6440 6585 6570 6615
rect 6400 6545 6570 6585
rect 6400 6515 6410 6545
rect 6440 6515 6570 6545
rect 6400 6495 6570 6515
rect -200 6430 -30 6450
rect -200 6400 -190 6430
rect -160 6400 -30 6430
rect -200 6360 -30 6400
rect -200 6330 -190 6360
rect -160 6330 -30 6360
rect -200 6310 -30 6330
rect 0 6430 170 6450
rect 0 6400 10 6430
rect 40 6400 170 6430
rect 0 6360 170 6400
rect 0 6330 10 6360
rect 40 6330 170 6360
rect 0 6310 170 6330
rect 200 6430 370 6450
rect 200 6400 210 6430
rect 240 6400 370 6430
rect 200 6360 370 6400
rect 200 6330 210 6360
rect 240 6330 370 6360
rect 200 6310 370 6330
rect 400 6430 570 6450
rect 400 6400 410 6430
rect 440 6400 570 6430
rect 400 6360 570 6400
rect 400 6330 410 6360
rect 440 6330 570 6360
rect 400 6310 570 6330
rect 600 6430 770 6450
rect 600 6400 610 6430
rect 640 6400 770 6430
rect 600 6360 770 6400
rect 600 6330 610 6360
rect 640 6330 770 6360
rect 600 6310 770 6330
rect 800 6430 970 6450
rect 800 6400 810 6430
rect 840 6400 970 6430
rect 800 6360 970 6400
rect 800 6330 810 6360
rect 840 6330 970 6360
rect 800 6310 970 6330
rect 1000 6430 1170 6450
rect 1000 6400 1010 6430
rect 1040 6400 1170 6430
rect 1000 6360 1170 6400
rect 1000 6330 1010 6360
rect 1040 6330 1170 6360
rect 1000 6310 1170 6330
rect 1200 6430 1370 6450
rect 1200 6400 1210 6430
rect 1240 6400 1370 6430
rect 1200 6360 1370 6400
rect 1200 6330 1210 6360
rect 1240 6330 1370 6360
rect 1200 6310 1370 6330
rect 1400 6430 1570 6450
rect 1400 6400 1410 6430
rect 1440 6400 1570 6430
rect 1400 6360 1570 6400
rect 1400 6330 1410 6360
rect 1440 6330 1570 6360
rect 1400 6310 1570 6330
rect 1600 6430 1770 6450
rect 1600 6400 1610 6430
rect 1640 6400 1770 6430
rect 1600 6360 1770 6400
rect 1600 6330 1610 6360
rect 1640 6330 1770 6360
rect 1600 6310 1770 6330
rect 1800 6430 1970 6450
rect 1800 6400 1810 6430
rect 1840 6400 1970 6430
rect 1800 6360 1970 6400
rect 1800 6330 1810 6360
rect 1840 6330 1970 6360
rect 1800 6310 1970 6330
rect 2000 6430 2170 6450
rect 2000 6400 2010 6430
rect 2040 6400 2170 6430
rect 2000 6360 2170 6400
rect 2000 6330 2010 6360
rect 2040 6330 2170 6360
rect 2000 6310 2170 6330
rect 2200 6430 2370 6450
rect 2200 6400 2210 6430
rect 2240 6400 2370 6430
rect 2200 6360 2370 6400
rect 2200 6330 2210 6360
rect 2240 6330 2370 6360
rect 2200 6310 2370 6330
rect 2400 6430 2570 6450
rect 2400 6400 2410 6430
rect 2440 6400 2570 6430
rect 2400 6360 2570 6400
rect 2400 6330 2410 6360
rect 2440 6330 2570 6360
rect 2400 6310 2570 6330
rect 2600 6430 2770 6450
rect 2600 6400 2610 6430
rect 2640 6400 2770 6430
rect 2600 6360 2770 6400
rect 2600 6330 2610 6360
rect 2640 6330 2770 6360
rect 2600 6310 2770 6330
rect 2800 6430 2970 6450
rect 2800 6400 2810 6430
rect 2840 6400 2970 6430
rect 2800 6360 2970 6400
rect 2800 6330 2810 6360
rect 2840 6330 2970 6360
rect 2800 6310 2970 6330
rect 3000 6430 3170 6450
rect 3000 6400 3010 6430
rect 3040 6400 3170 6430
rect 3000 6360 3170 6400
rect 3000 6330 3010 6360
rect 3040 6330 3170 6360
rect 3000 6310 3170 6330
rect 3200 6430 3370 6450
rect 3200 6400 3210 6430
rect 3240 6400 3370 6430
rect 3200 6360 3370 6400
rect 3200 6330 3210 6360
rect 3240 6330 3370 6360
rect 3200 6310 3370 6330
rect 3400 6430 3570 6450
rect 3400 6400 3410 6430
rect 3440 6400 3570 6430
rect 3400 6360 3570 6400
rect 3400 6330 3410 6360
rect 3440 6330 3570 6360
rect 3400 6310 3570 6330
rect 3600 6430 3770 6450
rect 3600 6400 3610 6430
rect 3640 6400 3770 6430
rect 3600 6360 3770 6400
rect 3600 6330 3610 6360
rect 3640 6330 3770 6360
rect 3600 6310 3770 6330
rect 3800 6430 3970 6450
rect 3800 6400 3810 6430
rect 3840 6400 3970 6430
rect 3800 6360 3970 6400
rect 3800 6330 3810 6360
rect 3840 6330 3970 6360
rect 3800 6310 3970 6330
rect 4000 6430 4170 6450
rect 4000 6400 4010 6430
rect 4040 6400 4170 6430
rect 4000 6360 4170 6400
rect 4000 6330 4010 6360
rect 4040 6330 4170 6360
rect 4000 6310 4170 6330
rect 4200 6430 4370 6450
rect 4200 6400 4210 6430
rect 4240 6400 4370 6430
rect 4200 6360 4370 6400
rect 4200 6330 4210 6360
rect 4240 6330 4370 6360
rect 4200 6310 4370 6330
rect 4400 6430 4570 6450
rect 4400 6400 4410 6430
rect 4440 6400 4570 6430
rect 4400 6360 4570 6400
rect 4400 6330 4410 6360
rect 4440 6330 4570 6360
rect 4400 6310 4570 6330
rect 4600 6430 4770 6450
rect 4600 6400 4610 6430
rect 4640 6400 4770 6430
rect 4600 6360 4770 6400
rect 4600 6330 4610 6360
rect 4640 6330 4770 6360
rect 4600 6310 4770 6330
rect 4800 6430 4970 6450
rect 4800 6400 4810 6430
rect 4840 6400 4970 6430
rect 4800 6360 4970 6400
rect 4800 6330 4810 6360
rect 4840 6330 4970 6360
rect 4800 6310 4970 6330
rect 5000 6430 5170 6450
rect 5000 6400 5010 6430
rect 5040 6400 5170 6430
rect 5000 6360 5170 6400
rect 5000 6330 5010 6360
rect 5040 6330 5170 6360
rect 5000 6310 5170 6330
rect 5200 6430 5370 6450
rect 5200 6400 5210 6430
rect 5240 6400 5370 6430
rect 5200 6360 5370 6400
rect 5200 6330 5210 6360
rect 5240 6330 5370 6360
rect 5200 6310 5370 6330
rect 5400 6430 5570 6450
rect 5400 6400 5410 6430
rect 5440 6400 5570 6430
rect 5400 6360 5570 6400
rect 5400 6330 5410 6360
rect 5440 6330 5570 6360
rect 5400 6310 5570 6330
rect 5600 6430 5770 6450
rect 5600 6400 5610 6430
rect 5640 6400 5770 6430
rect 5600 6360 5770 6400
rect 5600 6330 5610 6360
rect 5640 6330 5770 6360
rect 5600 6310 5770 6330
rect 5800 6430 5970 6450
rect 5800 6400 5810 6430
rect 5840 6400 5970 6430
rect 5800 6360 5970 6400
rect 5800 6330 5810 6360
rect 5840 6330 5970 6360
rect 5800 6310 5970 6330
rect 6000 6430 6170 6450
rect 6000 6400 6010 6430
rect 6040 6400 6170 6430
rect 6000 6360 6170 6400
rect 6000 6330 6010 6360
rect 6040 6330 6170 6360
rect 6000 6310 6170 6330
rect 6200 6430 6370 6450
rect 6200 6400 6210 6430
rect 6240 6400 6370 6430
rect 6200 6360 6370 6400
rect 6200 6330 6210 6360
rect 6240 6330 6370 6360
rect 6200 6310 6370 6330
rect 6400 6430 6570 6450
rect 6400 6400 6410 6430
rect 6440 6400 6570 6430
rect 6400 6360 6570 6400
rect 6400 6330 6410 6360
rect 6440 6330 6570 6360
rect 6400 6310 6570 6330
rect -200 6245 -30 6265
rect -200 6215 -190 6245
rect -160 6215 -30 6245
rect -200 6175 -30 6215
rect -200 6145 -190 6175
rect -160 6145 -30 6175
rect -200 6125 -30 6145
rect 0 6245 170 6265
rect 0 6215 10 6245
rect 40 6215 170 6245
rect 0 6175 170 6215
rect 0 6145 10 6175
rect 40 6145 170 6175
rect 0 6125 170 6145
rect 200 6245 370 6265
rect 200 6215 210 6245
rect 240 6215 370 6245
rect 200 6175 370 6215
rect 200 6145 210 6175
rect 240 6145 370 6175
rect 200 6125 370 6145
rect 400 6245 570 6265
rect 400 6215 410 6245
rect 440 6215 570 6245
rect 400 6175 570 6215
rect 400 6145 410 6175
rect 440 6145 570 6175
rect 400 6125 570 6145
rect 600 6245 770 6265
rect 600 6215 610 6245
rect 640 6215 770 6245
rect 600 6175 770 6215
rect 600 6145 610 6175
rect 640 6145 770 6175
rect 600 6125 770 6145
rect 800 6245 970 6265
rect 800 6215 810 6245
rect 840 6215 970 6245
rect 800 6175 970 6215
rect 800 6145 810 6175
rect 840 6145 970 6175
rect 800 6125 970 6145
rect 1000 6245 1170 6265
rect 1000 6215 1010 6245
rect 1040 6215 1170 6245
rect 1000 6175 1170 6215
rect 1000 6145 1010 6175
rect 1040 6145 1170 6175
rect 1000 6125 1170 6145
rect 1200 6245 1370 6265
rect 1200 6215 1210 6245
rect 1240 6215 1370 6245
rect 1200 6175 1370 6215
rect 1200 6145 1210 6175
rect 1240 6145 1370 6175
rect 1200 6125 1370 6145
rect 1400 6245 1570 6265
rect 1400 6215 1410 6245
rect 1440 6215 1570 6245
rect 1400 6175 1570 6215
rect 1400 6145 1410 6175
rect 1440 6145 1570 6175
rect 1400 6125 1570 6145
rect 1600 6245 1770 6265
rect 1600 6215 1610 6245
rect 1640 6215 1770 6245
rect 1600 6175 1770 6215
rect 1600 6145 1610 6175
rect 1640 6145 1770 6175
rect 1600 6125 1770 6145
rect 1800 6245 1970 6265
rect 1800 6215 1810 6245
rect 1840 6215 1970 6245
rect 1800 6175 1970 6215
rect 1800 6145 1810 6175
rect 1840 6145 1970 6175
rect 1800 6125 1970 6145
rect 2000 6245 2170 6265
rect 2000 6215 2010 6245
rect 2040 6215 2170 6245
rect 2000 6175 2170 6215
rect 2000 6145 2010 6175
rect 2040 6145 2170 6175
rect 2000 6125 2170 6145
rect 2200 6245 2370 6265
rect 2200 6215 2210 6245
rect 2240 6215 2370 6245
rect 2200 6175 2370 6215
rect 2200 6145 2210 6175
rect 2240 6145 2370 6175
rect 2200 6125 2370 6145
rect 2400 6245 2570 6265
rect 2400 6215 2410 6245
rect 2440 6215 2570 6245
rect 2400 6175 2570 6215
rect 2400 6145 2410 6175
rect 2440 6145 2570 6175
rect 2400 6125 2570 6145
rect 2600 6245 2770 6265
rect 2600 6215 2610 6245
rect 2640 6215 2770 6245
rect 2600 6175 2770 6215
rect 2600 6145 2610 6175
rect 2640 6145 2770 6175
rect 2600 6125 2770 6145
rect 2800 6245 2970 6265
rect 2800 6215 2810 6245
rect 2840 6215 2970 6245
rect 2800 6175 2970 6215
rect 2800 6145 2810 6175
rect 2840 6145 2970 6175
rect 2800 6125 2970 6145
rect 3000 6245 3170 6265
rect 3000 6215 3010 6245
rect 3040 6215 3170 6245
rect 3000 6175 3170 6215
rect 3000 6145 3010 6175
rect 3040 6145 3170 6175
rect 3000 6125 3170 6145
rect 3200 6245 3370 6265
rect 3200 6215 3210 6245
rect 3240 6215 3370 6245
rect 3200 6175 3370 6215
rect 3200 6145 3210 6175
rect 3240 6145 3370 6175
rect 3200 6125 3370 6145
rect 3400 6245 3570 6265
rect 3400 6215 3410 6245
rect 3440 6215 3570 6245
rect 3400 6175 3570 6215
rect 3400 6145 3410 6175
rect 3440 6145 3570 6175
rect 3400 6125 3570 6145
rect 3600 6245 3770 6265
rect 3600 6215 3610 6245
rect 3640 6215 3770 6245
rect 3600 6175 3770 6215
rect 3600 6145 3610 6175
rect 3640 6145 3770 6175
rect 3600 6125 3770 6145
rect 3800 6245 3970 6265
rect 3800 6215 3810 6245
rect 3840 6215 3970 6245
rect 3800 6175 3970 6215
rect 3800 6145 3810 6175
rect 3840 6145 3970 6175
rect 3800 6125 3970 6145
rect 4000 6245 4170 6265
rect 4000 6215 4010 6245
rect 4040 6215 4170 6245
rect 4000 6175 4170 6215
rect 4000 6145 4010 6175
rect 4040 6145 4170 6175
rect 4000 6125 4170 6145
rect 4200 6245 4370 6265
rect 4200 6215 4210 6245
rect 4240 6215 4370 6245
rect 4200 6175 4370 6215
rect 4200 6145 4210 6175
rect 4240 6145 4370 6175
rect 4200 6125 4370 6145
rect 4400 6245 4570 6265
rect 4400 6215 4410 6245
rect 4440 6215 4570 6245
rect 4400 6175 4570 6215
rect 4400 6145 4410 6175
rect 4440 6145 4570 6175
rect 4400 6125 4570 6145
rect 4600 6245 4770 6265
rect 4600 6215 4610 6245
rect 4640 6215 4770 6245
rect 4600 6175 4770 6215
rect 4600 6145 4610 6175
rect 4640 6145 4770 6175
rect 4600 6125 4770 6145
rect 4800 6245 4970 6265
rect 4800 6215 4810 6245
rect 4840 6215 4970 6245
rect 4800 6175 4970 6215
rect 4800 6145 4810 6175
rect 4840 6145 4970 6175
rect 4800 6125 4970 6145
rect 5000 6245 5170 6265
rect 5000 6215 5010 6245
rect 5040 6215 5170 6245
rect 5000 6175 5170 6215
rect 5000 6145 5010 6175
rect 5040 6145 5170 6175
rect 5000 6125 5170 6145
rect 5200 6245 5370 6265
rect 5200 6215 5210 6245
rect 5240 6215 5370 6245
rect 5200 6175 5370 6215
rect 5200 6145 5210 6175
rect 5240 6145 5370 6175
rect 5200 6125 5370 6145
rect 5400 6245 5570 6265
rect 5400 6215 5410 6245
rect 5440 6215 5570 6245
rect 5400 6175 5570 6215
rect 5400 6145 5410 6175
rect 5440 6145 5570 6175
rect 5400 6125 5570 6145
rect 5600 6245 5770 6265
rect 5600 6215 5610 6245
rect 5640 6215 5770 6245
rect 5600 6175 5770 6215
rect 5600 6145 5610 6175
rect 5640 6145 5770 6175
rect 5600 6125 5770 6145
rect 5800 6245 5970 6265
rect 5800 6215 5810 6245
rect 5840 6215 5970 6245
rect 5800 6175 5970 6215
rect 5800 6145 5810 6175
rect 5840 6145 5970 6175
rect 5800 6125 5970 6145
rect 6000 6245 6170 6265
rect 6000 6215 6010 6245
rect 6040 6215 6170 6245
rect 6000 6175 6170 6215
rect 6000 6145 6010 6175
rect 6040 6145 6170 6175
rect 6000 6125 6170 6145
rect 6200 6245 6370 6265
rect 6200 6215 6210 6245
rect 6240 6215 6370 6245
rect 6200 6175 6370 6215
rect 6200 6145 6210 6175
rect 6240 6145 6370 6175
rect 6200 6125 6370 6145
rect 6400 6245 6570 6265
rect 6400 6215 6410 6245
rect 6440 6215 6570 6245
rect 6400 6175 6570 6215
rect 6400 6145 6410 6175
rect 6440 6145 6570 6175
rect 6400 6125 6570 6145
rect -200 6060 -30 6080
rect -200 6030 -190 6060
rect -160 6030 -30 6060
rect -200 5990 -30 6030
rect -200 5960 -190 5990
rect -160 5960 -30 5990
rect -200 5940 -30 5960
rect 0 6060 170 6080
rect 0 6030 10 6060
rect 40 6030 170 6060
rect 0 5990 170 6030
rect 0 5960 10 5990
rect 40 5960 170 5990
rect 0 5940 170 5960
rect 200 6060 370 6080
rect 200 6030 210 6060
rect 240 6030 370 6060
rect 200 5990 370 6030
rect 200 5960 210 5990
rect 240 5960 370 5990
rect 200 5940 370 5960
rect 400 6060 570 6080
rect 400 6030 410 6060
rect 440 6030 570 6060
rect 400 5990 570 6030
rect 400 5960 410 5990
rect 440 5960 570 5990
rect 400 5940 570 5960
rect 600 6060 770 6080
rect 600 6030 610 6060
rect 640 6030 770 6060
rect 600 5990 770 6030
rect 600 5960 610 5990
rect 640 5960 770 5990
rect 600 5940 770 5960
rect 800 6060 970 6080
rect 800 6030 810 6060
rect 840 6030 970 6060
rect 800 5990 970 6030
rect 800 5960 810 5990
rect 840 5960 970 5990
rect 800 5940 970 5960
rect 1000 6060 1170 6080
rect 1000 6030 1010 6060
rect 1040 6030 1170 6060
rect 1000 5990 1170 6030
rect 1000 5960 1010 5990
rect 1040 5960 1170 5990
rect 1000 5940 1170 5960
rect 1200 6060 1370 6080
rect 1200 6030 1210 6060
rect 1240 6030 1370 6060
rect 1200 5990 1370 6030
rect 1200 5960 1210 5990
rect 1240 5960 1370 5990
rect 1200 5940 1370 5960
rect 1400 6060 1570 6080
rect 1400 6030 1410 6060
rect 1440 6030 1570 6060
rect 1400 5990 1570 6030
rect 1400 5960 1410 5990
rect 1440 5960 1570 5990
rect 1400 5940 1570 5960
rect 1600 6060 1770 6080
rect 1600 6030 1610 6060
rect 1640 6030 1770 6060
rect 1600 5990 1770 6030
rect 1600 5960 1610 5990
rect 1640 5960 1770 5990
rect 1600 5940 1770 5960
rect 1800 6060 1970 6080
rect 1800 6030 1810 6060
rect 1840 6030 1970 6060
rect 1800 5990 1970 6030
rect 1800 5960 1810 5990
rect 1840 5960 1970 5990
rect 1800 5940 1970 5960
rect 2000 6060 2170 6080
rect 2000 6030 2010 6060
rect 2040 6030 2170 6060
rect 2000 5990 2170 6030
rect 2000 5960 2010 5990
rect 2040 5960 2170 5990
rect 2000 5940 2170 5960
rect 2200 6060 2370 6080
rect 2200 6030 2210 6060
rect 2240 6030 2370 6060
rect 2200 5990 2370 6030
rect 2200 5960 2210 5990
rect 2240 5960 2370 5990
rect 2200 5940 2370 5960
rect 2400 6060 2570 6080
rect 2400 6030 2410 6060
rect 2440 6030 2570 6060
rect 2400 5990 2570 6030
rect 2400 5960 2410 5990
rect 2440 5960 2570 5990
rect 2400 5940 2570 5960
rect 2600 6060 2770 6080
rect 2600 6030 2610 6060
rect 2640 6030 2770 6060
rect 2600 5990 2770 6030
rect 2600 5960 2610 5990
rect 2640 5960 2770 5990
rect 2600 5940 2770 5960
rect 2800 6060 2970 6080
rect 2800 6030 2810 6060
rect 2840 6030 2970 6060
rect 2800 5990 2970 6030
rect 2800 5960 2810 5990
rect 2840 5960 2970 5990
rect 2800 5940 2970 5960
rect 3000 6060 3170 6080
rect 3000 6030 3010 6060
rect 3040 6030 3170 6060
rect 3000 5990 3170 6030
rect 3000 5960 3010 5990
rect 3040 5960 3170 5990
rect 3000 5940 3170 5960
rect 3200 6060 3370 6080
rect 3200 6030 3210 6060
rect 3240 6030 3370 6060
rect 3200 5990 3370 6030
rect 3200 5960 3210 5990
rect 3240 5960 3370 5990
rect 3200 5940 3370 5960
rect 3400 6060 3570 6080
rect 3400 6030 3410 6060
rect 3440 6030 3570 6060
rect 3400 5990 3570 6030
rect 3400 5960 3410 5990
rect 3440 5960 3570 5990
rect 3400 5940 3570 5960
rect 3600 6060 3770 6080
rect 3600 6030 3610 6060
rect 3640 6030 3770 6060
rect 3600 5990 3770 6030
rect 3600 5960 3610 5990
rect 3640 5960 3770 5990
rect 3600 5940 3770 5960
rect 3800 6060 3970 6080
rect 3800 6030 3810 6060
rect 3840 6030 3970 6060
rect 3800 5990 3970 6030
rect 3800 5960 3810 5990
rect 3840 5960 3970 5990
rect 3800 5940 3970 5960
rect 4000 6060 4170 6080
rect 4000 6030 4010 6060
rect 4040 6030 4170 6060
rect 4000 5990 4170 6030
rect 4000 5960 4010 5990
rect 4040 5960 4170 5990
rect 4000 5940 4170 5960
rect 4200 6060 4370 6080
rect 4200 6030 4210 6060
rect 4240 6030 4370 6060
rect 4200 5990 4370 6030
rect 4200 5960 4210 5990
rect 4240 5960 4370 5990
rect 4200 5940 4370 5960
rect 4400 6060 4570 6080
rect 4400 6030 4410 6060
rect 4440 6030 4570 6060
rect 4400 5990 4570 6030
rect 4400 5960 4410 5990
rect 4440 5960 4570 5990
rect 4400 5940 4570 5960
rect 4600 6060 4770 6080
rect 4600 6030 4610 6060
rect 4640 6030 4770 6060
rect 4600 5990 4770 6030
rect 4600 5960 4610 5990
rect 4640 5960 4770 5990
rect 4600 5940 4770 5960
rect 4800 6060 4970 6080
rect 4800 6030 4810 6060
rect 4840 6030 4970 6060
rect 4800 5990 4970 6030
rect 4800 5960 4810 5990
rect 4840 5960 4970 5990
rect 4800 5940 4970 5960
rect 5000 6060 5170 6080
rect 5000 6030 5010 6060
rect 5040 6030 5170 6060
rect 5000 5990 5170 6030
rect 5000 5960 5010 5990
rect 5040 5960 5170 5990
rect 5000 5940 5170 5960
rect 5200 6060 5370 6080
rect 5200 6030 5210 6060
rect 5240 6030 5370 6060
rect 5200 5990 5370 6030
rect 5200 5960 5210 5990
rect 5240 5960 5370 5990
rect 5200 5940 5370 5960
rect 5400 6060 5570 6080
rect 5400 6030 5410 6060
rect 5440 6030 5570 6060
rect 5400 5990 5570 6030
rect 5400 5960 5410 5990
rect 5440 5960 5570 5990
rect 5400 5940 5570 5960
rect 5600 6060 5770 6080
rect 5600 6030 5610 6060
rect 5640 6030 5770 6060
rect 5600 5990 5770 6030
rect 5600 5960 5610 5990
rect 5640 5960 5770 5990
rect 5600 5940 5770 5960
rect 5800 6060 5970 6080
rect 5800 6030 5810 6060
rect 5840 6030 5970 6060
rect 5800 5990 5970 6030
rect 5800 5960 5810 5990
rect 5840 5960 5970 5990
rect 5800 5940 5970 5960
rect 6000 6060 6170 6080
rect 6000 6030 6010 6060
rect 6040 6030 6170 6060
rect 6000 5990 6170 6030
rect 6000 5960 6010 5990
rect 6040 5960 6170 5990
rect 6000 5940 6170 5960
rect 6200 6060 6370 6080
rect 6200 6030 6210 6060
rect 6240 6030 6370 6060
rect 6200 5990 6370 6030
rect 6200 5960 6210 5990
rect 6240 5960 6370 5990
rect 6200 5940 6370 5960
rect 6400 6060 6570 6080
rect 6400 6030 6410 6060
rect 6440 6030 6570 6060
rect 6400 5990 6570 6030
rect 6400 5960 6410 5990
rect 6440 5960 6570 5990
rect 6400 5940 6570 5960
rect -200 5875 -30 5895
rect -200 5845 -190 5875
rect -160 5845 -30 5875
rect -200 5805 -30 5845
rect -200 5775 -190 5805
rect -160 5775 -30 5805
rect -200 5755 -30 5775
rect 0 5875 170 5895
rect 0 5845 10 5875
rect 40 5845 170 5875
rect 0 5805 170 5845
rect 0 5775 10 5805
rect 40 5775 170 5805
rect 0 5755 170 5775
rect 200 5875 370 5895
rect 200 5845 210 5875
rect 240 5845 370 5875
rect 200 5805 370 5845
rect 200 5775 210 5805
rect 240 5775 370 5805
rect 200 5755 370 5775
rect 400 5875 570 5895
rect 400 5845 410 5875
rect 440 5845 570 5875
rect 400 5805 570 5845
rect 400 5775 410 5805
rect 440 5775 570 5805
rect 400 5755 570 5775
rect 600 5875 770 5895
rect 600 5845 610 5875
rect 640 5845 770 5875
rect 600 5805 770 5845
rect 600 5775 610 5805
rect 640 5775 770 5805
rect 600 5755 770 5775
rect 800 5875 970 5895
rect 800 5845 810 5875
rect 840 5845 970 5875
rect 800 5805 970 5845
rect 800 5775 810 5805
rect 840 5775 970 5805
rect 800 5755 970 5775
rect 1000 5875 1170 5895
rect 1000 5845 1010 5875
rect 1040 5845 1170 5875
rect 1000 5805 1170 5845
rect 1000 5775 1010 5805
rect 1040 5775 1170 5805
rect 1000 5755 1170 5775
rect 1200 5875 1370 5895
rect 1200 5845 1210 5875
rect 1240 5845 1370 5875
rect 1200 5805 1370 5845
rect 1200 5775 1210 5805
rect 1240 5775 1370 5805
rect 1200 5755 1370 5775
rect 1400 5875 1570 5895
rect 1400 5845 1410 5875
rect 1440 5845 1570 5875
rect 1400 5805 1570 5845
rect 1400 5775 1410 5805
rect 1440 5775 1570 5805
rect 1400 5755 1570 5775
rect 1600 5875 1770 5895
rect 1600 5845 1610 5875
rect 1640 5845 1770 5875
rect 1600 5805 1770 5845
rect 1600 5775 1610 5805
rect 1640 5775 1770 5805
rect 1600 5755 1770 5775
rect 1800 5875 1970 5895
rect 1800 5845 1810 5875
rect 1840 5845 1970 5875
rect 1800 5805 1970 5845
rect 1800 5775 1810 5805
rect 1840 5775 1970 5805
rect 1800 5755 1970 5775
rect 2000 5875 2170 5895
rect 2000 5845 2010 5875
rect 2040 5845 2170 5875
rect 2000 5805 2170 5845
rect 2000 5775 2010 5805
rect 2040 5775 2170 5805
rect 2000 5755 2170 5775
rect 2200 5875 2370 5895
rect 2200 5845 2210 5875
rect 2240 5845 2370 5875
rect 2200 5805 2370 5845
rect 2200 5775 2210 5805
rect 2240 5775 2370 5805
rect 2200 5755 2370 5775
rect 2400 5875 2570 5895
rect 2400 5845 2410 5875
rect 2440 5845 2570 5875
rect 2400 5805 2570 5845
rect 2400 5775 2410 5805
rect 2440 5775 2570 5805
rect 2400 5755 2570 5775
rect 2600 5875 2770 5895
rect 2600 5845 2610 5875
rect 2640 5845 2770 5875
rect 2600 5805 2770 5845
rect 2600 5775 2610 5805
rect 2640 5775 2770 5805
rect 2600 5755 2770 5775
rect 2800 5875 2970 5895
rect 2800 5845 2810 5875
rect 2840 5845 2970 5875
rect 2800 5805 2970 5845
rect 2800 5775 2810 5805
rect 2840 5775 2970 5805
rect 2800 5755 2970 5775
rect 3000 5875 3170 5895
rect 3000 5845 3010 5875
rect 3040 5845 3170 5875
rect 3000 5805 3170 5845
rect 3000 5775 3010 5805
rect 3040 5775 3170 5805
rect 3000 5755 3170 5775
rect 3200 5875 3370 5895
rect 3200 5845 3210 5875
rect 3240 5845 3370 5875
rect 3200 5805 3370 5845
rect 3200 5775 3210 5805
rect 3240 5775 3370 5805
rect 3200 5755 3370 5775
rect 3400 5875 3570 5895
rect 3400 5845 3410 5875
rect 3440 5845 3570 5875
rect 3400 5805 3570 5845
rect 3400 5775 3410 5805
rect 3440 5775 3570 5805
rect 3400 5755 3570 5775
rect 3600 5875 3770 5895
rect 3600 5845 3610 5875
rect 3640 5845 3770 5875
rect 3600 5805 3770 5845
rect 3600 5775 3610 5805
rect 3640 5775 3770 5805
rect 3600 5755 3770 5775
rect 3800 5875 3970 5895
rect 3800 5845 3810 5875
rect 3840 5845 3970 5875
rect 3800 5805 3970 5845
rect 3800 5775 3810 5805
rect 3840 5775 3970 5805
rect 3800 5755 3970 5775
rect 4000 5875 4170 5895
rect 4000 5845 4010 5875
rect 4040 5845 4170 5875
rect 4000 5805 4170 5845
rect 4000 5775 4010 5805
rect 4040 5775 4170 5805
rect 4000 5755 4170 5775
rect 4200 5875 4370 5895
rect 4200 5845 4210 5875
rect 4240 5845 4370 5875
rect 4200 5805 4370 5845
rect 4200 5775 4210 5805
rect 4240 5775 4370 5805
rect 4200 5755 4370 5775
rect 4400 5875 4570 5895
rect 4400 5845 4410 5875
rect 4440 5845 4570 5875
rect 4400 5805 4570 5845
rect 4400 5775 4410 5805
rect 4440 5775 4570 5805
rect 4400 5755 4570 5775
rect 4600 5875 4770 5895
rect 4600 5845 4610 5875
rect 4640 5845 4770 5875
rect 4600 5805 4770 5845
rect 4600 5775 4610 5805
rect 4640 5775 4770 5805
rect 4600 5755 4770 5775
rect 4800 5875 4970 5895
rect 4800 5845 4810 5875
rect 4840 5845 4970 5875
rect 4800 5805 4970 5845
rect 4800 5775 4810 5805
rect 4840 5775 4970 5805
rect 4800 5755 4970 5775
rect 5000 5875 5170 5895
rect 5000 5845 5010 5875
rect 5040 5845 5170 5875
rect 5000 5805 5170 5845
rect 5000 5775 5010 5805
rect 5040 5775 5170 5805
rect 5000 5755 5170 5775
rect 5200 5875 5370 5895
rect 5200 5845 5210 5875
rect 5240 5845 5370 5875
rect 5200 5805 5370 5845
rect 5200 5775 5210 5805
rect 5240 5775 5370 5805
rect 5200 5755 5370 5775
rect 5400 5875 5570 5895
rect 5400 5845 5410 5875
rect 5440 5845 5570 5875
rect 5400 5805 5570 5845
rect 5400 5775 5410 5805
rect 5440 5775 5570 5805
rect 5400 5755 5570 5775
rect 5600 5875 5770 5895
rect 5600 5845 5610 5875
rect 5640 5845 5770 5875
rect 5600 5805 5770 5845
rect 5600 5775 5610 5805
rect 5640 5775 5770 5805
rect 5600 5755 5770 5775
rect 5800 5875 5970 5895
rect 5800 5845 5810 5875
rect 5840 5845 5970 5875
rect 5800 5805 5970 5845
rect 5800 5775 5810 5805
rect 5840 5775 5970 5805
rect 5800 5755 5970 5775
rect 6000 5875 6170 5895
rect 6000 5845 6010 5875
rect 6040 5845 6170 5875
rect 6000 5805 6170 5845
rect 6000 5775 6010 5805
rect 6040 5775 6170 5805
rect 6000 5755 6170 5775
rect 6200 5875 6370 5895
rect 6200 5845 6210 5875
rect 6240 5845 6370 5875
rect 6200 5805 6370 5845
rect 6200 5775 6210 5805
rect 6240 5775 6370 5805
rect 6200 5755 6370 5775
rect 6400 5875 6570 5895
rect 6400 5845 6410 5875
rect 6440 5845 6570 5875
rect 6400 5805 6570 5845
rect 6400 5775 6410 5805
rect 6440 5775 6570 5805
rect 6400 5755 6570 5775
rect -200 5690 -30 5710
rect -200 5660 -190 5690
rect -160 5660 -30 5690
rect -200 5620 -30 5660
rect -200 5590 -190 5620
rect -160 5590 -30 5620
rect -200 5570 -30 5590
rect 0 5690 170 5710
rect 0 5660 10 5690
rect 40 5660 170 5690
rect 0 5620 170 5660
rect 0 5590 10 5620
rect 40 5590 170 5620
rect 0 5570 170 5590
rect 200 5690 370 5710
rect 200 5660 210 5690
rect 240 5660 370 5690
rect 200 5620 370 5660
rect 200 5590 210 5620
rect 240 5590 370 5620
rect 200 5570 370 5590
rect 400 5690 570 5710
rect 400 5660 410 5690
rect 440 5660 570 5690
rect 400 5620 570 5660
rect 400 5590 410 5620
rect 440 5590 570 5620
rect 400 5570 570 5590
rect 600 5690 770 5710
rect 600 5660 610 5690
rect 640 5660 770 5690
rect 600 5620 770 5660
rect 600 5590 610 5620
rect 640 5590 770 5620
rect 600 5570 770 5590
rect 800 5690 970 5710
rect 800 5660 810 5690
rect 840 5660 970 5690
rect 800 5620 970 5660
rect 800 5590 810 5620
rect 840 5590 970 5620
rect 800 5570 970 5590
rect 1000 5690 1170 5710
rect 1000 5660 1010 5690
rect 1040 5660 1170 5690
rect 1000 5620 1170 5660
rect 1000 5590 1010 5620
rect 1040 5590 1170 5620
rect 1000 5570 1170 5590
rect 1200 5690 1370 5710
rect 1200 5660 1210 5690
rect 1240 5660 1370 5690
rect 1200 5620 1370 5660
rect 1200 5590 1210 5620
rect 1240 5590 1370 5620
rect 1200 5570 1370 5590
rect 1400 5690 1570 5710
rect 1400 5660 1410 5690
rect 1440 5660 1570 5690
rect 1400 5620 1570 5660
rect 1400 5590 1410 5620
rect 1440 5590 1570 5620
rect 1400 5570 1570 5590
rect 1600 5690 1770 5710
rect 1600 5660 1610 5690
rect 1640 5660 1770 5690
rect 1600 5620 1770 5660
rect 1600 5590 1610 5620
rect 1640 5590 1770 5620
rect 1600 5570 1770 5590
rect 1800 5690 1970 5710
rect 1800 5660 1810 5690
rect 1840 5660 1970 5690
rect 1800 5620 1970 5660
rect 1800 5590 1810 5620
rect 1840 5590 1970 5620
rect 1800 5570 1970 5590
rect 2000 5690 2170 5710
rect 2000 5660 2010 5690
rect 2040 5660 2170 5690
rect 2000 5620 2170 5660
rect 2000 5590 2010 5620
rect 2040 5590 2170 5620
rect 2000 5570 2170 5590
rect 2200 5690 2370 5710
rect 2200 5660 2210 5690
rect 2240 5660 2370 5690
rect 2200 5620 2370 5660
rect 2200 5590 2210 5620
rect 2240 5590 2370 5620
rect 2200 5570 2370 5590
rect 2400 5690 2570 5710
rect 2400 5660 2410 5690
rect 2440 5660 2570 5690
rect 2400 5620 2570 5660
rect 2400 5590 2410 5620
rect 2440 5590 2570 5620
rect 2400 5570 2570 5590
rect 2600 5690 2770 5710
rect 2600 5660 2610 5690
rect 2640 5660 2770 5690
rect 2600 5620 2770 5660
rect 2600 5590 2610 5620
rect 2640 5590 2770 5620
rect 2600 5570 2770 5590
rect 2800 5690 2970 5710
rect 2800 5660 2810 5690
rect 2840 5660 2970 5690
rect 2800 5620 2970 5660
rect 2800 5590 2810 5620
rect 2840 5590 2970 5620
rect 2800 5570 2970 5590
rect 3000 5690 3170 5710
rect 3000 5660 3010 5690
rect 3040 5660 3170 5690
rect 3000 5620 3170 5660
rect 3000 5590 3010 5620
rect 3040 5590 3170 5620
rect 3000 5570 3170 5590
rect 3200 5690 3370 5710
rect 3200 5660 3210 5690
rect 3240 5660 3370 5690
rect 3200 5620 3370 5660
rect 3200 5590 3210 5620
rect 3240 5590 3370 5620
rect 3200 5570 3370 5590
rect 3400 5690 3570 5710
rect 3400 5660 3410 5690
rect 3440 5660 3570 5690
rect 3400 5620 3570 5660
rect 3400 5590 3410 5620
rect 3440 5590 3570 5620
rect 3400 5570 3570 5590
rect 3600 5690 3770 5710
rect 3600 5660 3610 5690
rect 3640 5660 3770 5690
rect 3600 5620 3770 5660
rect 3600 5590 3610 5620
rect 3640 5590 3770 5620
rect 3600 5570 3770 5590
rect 3800 5690 3970 5710
rect 3800 5660 3810 5690
rect 3840 5660 3970 5690
rect 3800 5620 3970 5660
rect 3800 5590 3810 5620
rect 3840 5590 3970 5620
rect 3800 5570 3970 5590
rect 4000 5690 4170 5710
rect 4000 5660 4010 5690
rect 4040 5660 4170 5690
rect 4000 5620 4170 5660
rect 4000 5590 4010 5620
rect 4040 5590 4170 5620
rect 4000 5570 4170 5590
rect 4200 5690 4370 5710
rect 4200 5660 4210 5690
rect 4240 5660 4370 5690
rect 4200 5620 4370 5660
rect 4200 5590 4210 5620
rect 4240 5590 4370 5620
rect 4200 5570 4370 5590
rect 4400 5690 4570 5710
rect 4400 5660 4410 5690
rect 4440 5660 4570 5690
rect 4400 5620 4570 5660
rect 4400 5590 4410 5620
rect 4440 5590 4570 5620
rect 4400 5570 4570 5590
rect 4600 5690 4770 5710
rect 4600 5660 4610 5690
rect 4640 5660 4770 5690
rect 4600 5620 4770 5660
rect 4600 5590 4610 5620
rect 4640 5590 4770 5620
rect 4600 5570 4770 5590
rect 4800 5690 4970 5710
rect 4800 5660 4810 5690
rect 4840 5660 4970 5690
rect 4800 5620 4970 5660
rect 4800 5590 4810 5620
rect 4840 5590 4970 5620
rect 4800 5570 4970 5590
rect 5000 5690 5170 5710
rect 5000 5660 5010 5690
rect 5040 5660 5170 5690
rect 5000 5620 5170 5660
rect 5000 5590 5010 5620
rect 5040 5590 5170 5620
rect 5000 5570 5170 5590
rect 5200 5690 5370 5710
rect 5200 5660 5210 5690
rect 5240 5660 5370 5690
rect 5200 5620 5370 5660
rect 5200 5590 5210 5620
rect 5240 5590 5370 5620
rect 5200 5570 5370 5590
rect 5400 5690 5570 5710
rect 5400 5660 5410 5690
rect 5440 5660 5570 5690
rect 5400 5620 5570 5660
rect 5400 5590 5410 5620
rect 5440 5590 5570 5620
rect 5400 5570 5570 5590
rect 5600 5690 5770 5710
rect 5600 5660 5610 5690
rect 5640 5660 5770 5690
rect 5600 5620 5770 5660
rect 5600 5590 5610 5620
rect 5640 5590 5770 5620
rect 5600 5570 5770 5590
rect 5800 5690 5970 5710
rect 5800 5660 5810 5690
rect 5840 5660 5970 5690
rect 5800 5620 5970 5660
rect 5800 5590 5810 5620
rect 5840 5590 5970 5620
rect 5800 5570 5970 5590
rect 6000 5690 6170 5710
rect 6000 5660 6010 5690
rect 6040 5660 6170 5690
rect 6000 5620 6170 5660
rect 6000 5590 6010 5620
rect 6040 5590 6170 5620
rect 6000 5570 6170 5590
rect 6200 5690 6370 5710
rect 6200 5660 6210 5690
rect 6240 5660 6370 5690
rect 6200 5620 6370 5660
rect 6200 5590 6210 5620
rect 6240 5590 6370 5620
rect 6200 5570 6370 5590
rect 6400 5690 6570 5710
rect 6400 5660 6410 5690
rect 6440 5660 6570 5690
rect 6400 5620 6570 5660
rect 6400 5590 6410 5620
rect 6440 5590 6570 5620
rect 6400 5570 6570 5590
rect -200 5505 -30 5525
rect -200 5475 -190 5505
rect -160 5475 -30 5505
rect -200 5435 -30 5475
rect -200 5405 -190 5435
rect -160 5405 -30 5435
rect -200 5385 -30 5405
rect 0 5505 170 5525
rect 0 5475 10 5505
rect 40 5475 170 5505
rect 0 5435 170 5475
rect 0 5405 10 5435
rect 40 5405 170 5435
rect 0 5385 170 5405
rect 200 5505 370 5525
rect 200 5475 210 5505
rect 240 5475 370 5505
rect 200 5435 370 5475
rect 200 5405 210 5435
rect 240 5405 370 5435
rect 200 5385 370 5405
rect 400 5505 570 5525
rect 400 5475 410 5505
rect 440 5475 570 5505
rect 400 5435 570 5475
rect 400 5405 410 5435
rect 440 5405 570 5435
rect 400 5385 570 5405
rect 600 5505 770 5525
rect 600 5475 610 5505
rect 640 5475 770 5505
rect 600 5435 770 5475
rect 600 5405 610 5435
rect 640 5405 770 5435
rect 600 5385 770 5405
rect 800 5505 970 5525
rect 800 5475 810 5505
rect 840 5475 970 5505
rect 800 5435 970 5475
rect 800 5405 810 5435
rect 840 5405 970 5435
rect 800 5385 970 5405
rect 1000 5505 1170 5525
rect 1000 5475 1010 5505
rect 1040 5475 1170 5505
rect 1000 5435 1170 5475
rect 1000 5405 1010 5435
rect 1040 5405 1170 5435
rect 1000 5385 1170 5405
rect 1200 5505 1370 5525
rect 1200 5475 1210 5505
rect 1240 5475 1370 5505
rect 1200 5435 1370 5475
rect 1200 5405 1210 5435
rect 1240 5405 1370 5435
rect 1200 5385 1370 5405
rect 1400 5505 1570 5525
rect 1400 5475 1410 5505
rect 1440 5475 1570 5505
rect 1400 5435 1570 5475
rect 1400 5405 1410 5435
rect 1440 5405 1570 5435
rect 1400 5385 1570 5405
rect 1600 5505 1770 5525
rect 1600 5475 1610 5505
rect 1640 5475 1770 5505
rect 1600 5435 1770 5475
rect 1600 5405 1610 5435
rect 1640 5405 1770 5435
rect 1600 5385 1770 5405
rect 1800 5505 1970 5525
rect 1800 5475 1810 5505
rect 1840 5475 1970 5505
rect 1800 5435 1970 5475
rect 1800 5405 1810 5435
rect 1840 5405 1970 5435
rect 1800 5385 1970 5405
rect 2000 5505 2170 5525
rect 2000 5475 2010 5505
rect 2040 5475 2170 5505
rect 2000 5435 2170 5475
rect 2000 5405 2010 5435
rect 2040 5405 2170 5435
rect 2000 5385 2170 5405
rect 2200 5505 2370 5525
rect 2200 5475 2210 5505
rect 2240 5475 2370 5505
rect 2200 5435 2370 5475
rect 2200 5405 2210 5435
rect 2240 5405 2370 5435
rect 2200 5385 2370 5405
rect 2400 5505 2570 5525
rect 2400 5475 2410 5505
rect 2440 5475 2570 5505
rect 2400 5435 2570 5475
rect 2400 5405 2410 5435
rect 2440 5405 2570 5435
rect 2400 5385 2570 5405
rect 2600 5505 2770 5525
rect 2600 5475 2610 5505
rect 2640 5475 2770 5505
rect 2600 5435 2770 5475
rect 2600 5405 2610 5435
rect 2640 5405 2770 5435
rect 2600 5385 2770 5405
rect 2800 5505 2970 5525
rect 2800 5475 2810 5505
rect 2840 5475 2970 5505
rect 2800 5435 2970 5475
rect 2800 5405 2810 5435
rect 2840 5405 2970 5435
rect 2800 5385 2970 5405
rect 3000 5505 3170 5525
rect 3000 5475 3010 5505
rect 3040 5475 3170 5505
rect 3000 5435 3170 5475
rect 3000 5405 3010 5435
rect 3040 5405 3170 5435
rect 3000 5385 3170 5405
rect 3200 5505 3370 5525
rect 3200 5475 3210 5505
rect 3240 5475 3370 5505
rect 3200 5435 3370 5475
rect 3200 5405 3210 5435
rect 3240 5405 3370 5435
rect 3200 5385 3370 5405
rect 3400 5505 3570 5525
rect 3400 5475 3410 5505
rect 3440 5475 3570 5505
rect 3400 5435 3570 5475
rect 3400 5405 3410 5435
rect 3440 5405 3570 5435
rect 3400 5385 3570 5405
rect 3600 5505 3770 5525
rect 3600 5475 3610 5505
rect 3640 5475 3770 5505
rect 3600 5435 3770 5475
rect 3600 5405 3610 5435
rect 3640 5405 3770 5435
rect 3600 5385 3770 5405
rect 3800 5505 3970 5525
rect 3800 5475 3810 5505
rect 3840 5475 3970 5505
rect 3800 5435 3970 5475
rect 3800 5405 3810 5435
rect 3840 5405 3970 5435
rect 3800 5385 3970 5405
rect 4000 5505 4170 5525
rect 4000 5475 4010 5505
rect 4040 5475 4170 5505
rect 4000 5435 4170 5475
rect 4000 5405 4010 5435
rect 4040 5405 4170 5435
rect 4000 5385 4170 5405
rect 4200 5505 4370 5525
rect 4200 5475 4210 5505
rect 4240 5475 4370 5505
rect 4200 5435 4370 5475
rect 4200 5405 4210 5435
rect 4240 5405 4370 5435
rect 4200 5385 4370 5405
rect 4400 5505 4570 5525
rect 4400 5475 4410 5505
rect 4440 5475 4570 5505
rect 4400 5435 4570 5475
rect 4400 5405 4410 5435
rect 4440 5405 4570 5435
rect 4400 5385 4570 5405
rect 4600 5505 4770 5525
rect 4600 5475 4610 5505
rect 4640 5475 4770 5505
rect 4600 5435 4770 5475
rect 4600 5405 4610 5435
rect 4640 5405 4770 5435
rect 4600 5385 4770 5405
rect 4800 5505 4970 5525
rect 4800 5475 4810 5505
rect 4840 5475 4970 5505
rect 4800 5435 4970 5475
rect 4800 5405 4810 5435
rect 4840 5405 4970 5435
rect 4800 5385 4970 5405
rect 5000 5505 5170 5525
rect 5000 5475 5010 5505
rect 5040 5475 5170 5505
rect 5000 5435 5170 5475
rect 5000 5405 5010 5435
rect 5040 5405 5170 5435
rect 5000 5385 5170 5405
rect 5200 5505 5370 5525
rect 5200 5475 5210 5505
rect 5240 5475 5370 5505
rect 5200 5435 5370 5475
rect 5200 5405 5210 5435
rect 5240 5405 5370 5435
rect 5200 5385 5370 5405
rect 5400 5505 5570 5525
rect 5400 5475 5410 5505
rect 5440 5475 5570 5505
rect 5400 5435 5570 5475
rect 5400 5405 5410 5435
rect 5440 5405 5570 5435
rect 5400 5385 5570 5405
rect 5600 5505 5770 5525
rect 5600 5475 5610 5505
rect 5640 5475 5770 5505
rect 5600 5435 5770 5475
rect 5600 5405 5610 5435
rect 5640 5405 5770 5435
rect 5600 5385 5770 5405
rect 5800 5505 5970 5525
rect 5800 5475 5810 5505
rect 5840 5475 5970 5505
rect 5800 5435 5970 5475
rect 5800 5405 5810 5435
rect 5840 5405 5970 5435
rect 5800 5385 5970 5405
rect 6000 5505 6170 5525
rect 6000 5475 6010 5505
rect 6040 5475 6170 5505
rect 6000 5435 6170 5475
rect 6000 5405 6010 5435
rect 6040 5405 6170 5435
rect 6000 5385 6170 5405
rect 6200 5505 6370 5525
rect 6200 5475 6210 5505
rect 6240 5475 6370 5505
rect 6200 5435 6370 5475
rect 6200 5405 6210 5435
rect 6240 5405 6370 5435
rect 6200 5385 6370 5405
rect 6400 5505 6570 5525
rect 6400 5475 6410 5505
rect 6440 5475 6570 5505
rect 6400 5435 6570 5475
rect 6400 5405 6410 5435
rect 6440 5405 6570 5435
rect 6400 5385 6570 5405
rect -200 5320 -30 5340
rect -200 5290 -190 5320
rect -160 5290 -30 5320
rect -200 5250 -30 5290
rect -200 5220 -190 5250
rect -160 5220 -30 5250
rect -200 5200 -30 5220
rect 0 5320 170 5340
rect 0 5290 10 5320
rect 40 5290 170 5320
rect 0 5250 170 5290
rect 0 5220 10 5250
rect 40 5220 170 5250
rect 0 5200 170 5220
rect 200 5320 370 5340
rect 200 5290 210 5320
rect 240 5290 370 5320
rect 200 5250 370 5290
rect 200 5220 210 5250
rect 240 5220 370 5250
rect 200 5200 370 5220
rect 400 5320 570 5340
rect 400 5290 410 5320
rect 440 5290 570 5320
rect 400 5250 570 5290
rect 400 5220 410 5250
rect 440 5220 570 5250
rect 400 5200 570 5220
rect 600 5320 770 5340
rect 600 5290 610 5320
rect 640 5290 770 5320
rect 600 5250 770 5290
rect 600 5220 610 5250
rect 640 5220 770 5250
rect 600 5200 770 5220
rect 800 5320 970 5340
rect 800 5290 810 5320
rect 840 5290 970 5320
rect 800 5250 970 5290
rect 800 5220 810 5250
rect 840 5220 970 5250
rect 800 5200 970 5220
rect 1000 5320 1170 5340
rect 1000 5290 1010 5320
rect 1040 5290 1170 5320
rect 1000 5250 1170 5290
rect 1000 5220 1010 5250
rect 1040 5220 1170 5250
rect 1000 5200 1170 5220
rect 1200 5320 1370 5340
rect 1200 5290 1210 5320
rect 1240 5290 1370 5320
rect 1200 5250 1370 5290
rect 1200 5220 1210 5250
rect 1240 5220 1370 5250
rect 1200 5200 1370 5220
rect 1400 5320 1570 5340
rect 1400 5290 1410 5320
rect 1440 5290 1570 5320
rect 1400 5250 1570 5290
rect 1400 5220 1410 5250
rect 1440 5220 1570 5250
rect 1400 5200 1570 5220
rect 1600 5320 1770 5340
rect 1600 5290 1610 5320
rect 1640 5290 1770 5320
rect 1600 5250 1770 5290
rect 1600 5220 1610 5250
rect 1640 5220 1770 5250
rect 1600 5200 1770 5220
rect 1800 5320 1970 5340
rect 1800 5290 1810 5320
rect 1840 5290 1970 5320
rect 1800 5250 1970 5290
rect 1800 5220 1810 5250
rect 1840 5220 1970 5250
rect 1800 5200 1970 5220
rect 2000 5320 2170 5340
rect 2000 5290 2010 5320
rect 2040 5290 2170 5320
rect 2000 5250 2170 5290
rect 2000 5220 2010 5250
rect 2040 5220 2170 5250
rect 2000 5200 2170 5220
rect 2200 5320 2370 5340
rect 2200 5290 2210 5320
rect 2240 5290 2370 5320
rect 2200 5250 2370 5290
rect 2200 5220 2210 5250
rect 2240 5220 2370 5250
rect 2200 5200 2370 5220
rect 2400 5320 2570 5340
rect 2400 5290 2410 5320
rect 2440 5290 2570 5320
rect 2400 5250 2570 5290
rect 2400 5220 2410 5250
rect 2440 5220 2570 5250
rect 2400 5200 2570 5220
rect 2600 5320 2770 5340
rect 2600 5290 2610 5320
rect 2640 5290 2770 5320
rect 2600 5250 2770 5290
rect 2600 5220 2610 5250
rect 2640 5220 2770 5250
rect 2600 5200 2770 5220
rect 2800 5320 2970 5340
rect 2800 5290 2810 5320
rect 2840 5290 2970 5320
rect 2800 5250 2970 5290
rect 2800 5220 2810 5250
rect 2840 5220 2970 5250
rect 2800 5200 2970 5220
rect 3000 5320 3170 5340
rect 3000 5290 3010 5320
rect 3040 5290 3170 5320
rect 3000 5250 3170 5290
rect 3000 5220 3010 5250
rect 3040 5220 3170 5250
rect 3000 5200 3170 5220
rect 3200 5320 3370 5340
rect 3200 5290 3210 5320
rect 3240 5290 3370 5320
rect 3200 5250 3370 5290
rect 3200 5220 3210 5250
rect 3240 5220 3370 5250
rect 3200 5200 3370 5220
rect 3400 5320 3570 5340
rect 3400 5290 3410 5320
rect 3440 5290 3570 5320
rect 3400 5250 3570 5290
rect 3400 5220 3410 5250
rect 3440 5220 3570 5250
rect 3400 5200 3570 5220
rect 3600 5320 3770 5340
rect 3600 5290 3610 5320
rect 3640 5290 3770 5320
rect 3600 5250 3770 5290
rect 3600 5220 3610 5250
rect 3640 5220 3770 5250
rect 3600 5200 3770 5220
rect 3800 5320 3970 5340
rect 3800 5290 3810 5320
rect 3840 5290 3970 5320
rect 3800 5250 3970 5290
rect 3800 5220 3810 5250
rect 3840 5220 3970 5250
rect 3800 5200 3970 5220
rect 4000 5320 4170 5340
rect 4000 5290 4010 5320
rect 4040 5290 4170 5320
rect 4000 5250 4170 5290
rect 4000 5220 4010 5250
rect 4040 5220 4170 5250
rect 4000 5200 4170 5220
rect 4200 5320 4370 5340
rect 4200 5290 4210 5320
rect 4240 5290 4370 5320
rect 4200 5250 4370 5290
rect 4200 5220 4210 5250
rect 4240 5220 4370 5250
rect 4200 5200 4370 5220
rect 4400 5320 4570 5340
rect 4400 5290 4410 5320
rect 4440 5290 4570 5320
rect 4400 5250 4570 5290
rect 4400 5220 4410 5250
rect 4440 5220 4570 5250
rect 4400 5200 4570 5220
rect 4600 5320 4770 5340
rect 4600 5290 4610 5320
rect 4640 5290 4770 5320
rect 4600 5250 4770 5290
rect 4600 5220 4610 5250
rect 4640 5220 4770 5250
rect 4600 5200 4770 5220
rect 4800 5320 4970 5340
rect 4800 5290 4810 5320
rect 4840 5290 4970 5320
rect 4800 5250 4970 5290
rect 4800 5220 4810 5250
rect 4840 5220 4970 5250
rect 4800 5200 4970 5220
rect 5000 5320 5170 5340
rect 5000 5290 5010 5320
rect 5040 5290 5170 5320
rect 5000 5250 5170 5290
rect 5000 5220 5010 5250
rect 5040 5220 5170 5250
rect 5000 5200 5170 5220
rect 5200 5320 5370 5340
rect 5200 5290 5210 5320
rect 5240 5290 5370 5320
rect 5200 5250 5370 5290
rect 5200 5220 5210 5250
rect 5240 5220 5370 5250
rect 5200 5200 5370 5220
rect 5400 5320 5570 5340
rect 5400 5290 5410 5320
rect 5440 5290 5570 5320
rect 5400 5250 5570 5290
rect 5400 5220 5410 5250
rect 5440 5220 5570 5250
rect 5400 5200 5570 5220
rect 5600 5320 5770 5340
rect 5600 5290 5610 5320
rect 5640 5290 5770 5320
rect 5600 5250 5770 5290
rect 5600 5220 5610 5250
rect 5640 5220 5770 5250
rect 5600 5200 5770 5220
rect 5800 5320 5970 5340
rect 5800 5290 5810 5320
rect 5840 5290 5970 5320
rect 5800 5250 5970 5290
rect 5800 5220 5810 5250
rect 5840 5220 5970 5250
rect 5800 5200 5970 5220
rect 6000 5320 6170 5340
rect 6000 5290 6010 5320
rect 6040 5290 6170 5320
rect 6000 5250 6170 5290
rect 6000 5220 6010 5250
rect 6040 5220 6170 5250
rect 6000 5200 6170 5220
rect 6200 5320 6370 5340
rect 6200 5290 6210 5320
rect 6240 5290 6370 5320
rect 6200 5250 6370 5290
rect 6200 5220 6210 5250
rect 6240 5220 6370 5250
rect 6200 5200 6370 5220
rect 6400 5320 6570 5340
rect 6400 5290 6410 5320
rect 6440 5290 6570 5320
rect 6400 5250 6570 5290
rect 6400 5220 6410 5250
rect 6440 5220 6570 5250
rect 6400 5200 6570 5220
rect -200 5135 -30 5155
rect -200 5105 -190 5135
rect -160 5105 -30 5135
rect -200 5065 -30 5105
rect -200 5035 -190 5065
rect -160 5035 -30 5065
rect -200 5015 -30 5035
rect 0 5135 170 5155
rect 0 5105 10 5135
rect 40 5105 170 5135
rect 0 5065 170 5105
rect 0 5035 10 5065
rect 40 5035 170 5065
rect 0 5015 170 5035
rect 200 5135 370 5155
rect 200 5105 210 5135
rect 240 5105 370 5135
rect 200 5065 370 5105
rect 200 5035 210 5065
rect 240 5035 370 5065
rect 200 5015 370 5035
rect 400 5135 570 5155
rect 400 5105 410 5135
rect 440 5105 570 5135
rect 400 5065 570 5105
rect 400 5035 410 5065
rect 440 5035 570 5065
rect 400 5015 570 5035
rect 600 5135 770 5155
rect 600 5105 610 5135
rect 640 5105 770 5135
rect 600 5065 770 5105
rect 600 5035 610 5065
rect 640 5035 770 5065
rect 600 5015 770 5035
rect 800 5135 970 5155
rect 800 5105 810 5135
rect 840 5105 970 5135
rect 800 5065 970 5105
rect 800 5035 810 5065
rect 840 5035 970 5065
rect 800 5015 970 5035
rect 1000 5135 1170 5155
rect 1000 5105 1010 5135
rect 1040 5105 1170 5135
rect 1000 5065 1170 5105
rect 1000 5035 1010 5065
rect 1040 5035 1170 5065
rect 1000 5015 1170 5035
rect 1200 5135 1370 5155
rect 1200 5105 1210 5135
rect 1240 5105 1370 5135
rect 1200 5065 1370 5105
rect 1200 5035 1210 5065
rect 1240 5035 1370 5065
rect 1200 5015 1370 5035
rect 1400 5135 1570 5155
rect 1400 5105 1410 5135
rect 1440 5105 1570 5135
rect 1400 5065 1570 5105
rect 1400 5035 1410 5065
rect 1440 5035 1570 5065
rect 1400 5015 1570 5035
rect 1600 5135 1770 5155
rect 1600 5105 1610 5135
rect 1640 5105 1770 5135
rect 1600 5065 1770 5105
rect 1600 5035 1610 5065
rect 1640 5035 1770 5065
rect 1600 5015 1770 5035
rect 1800 5135 1970 5155
rect 1800 5105 1810 5135
rect 1840 5105 1970 5135
rect 1800 5065 1970 5105
rect 1800 5035 1810 5065
rect 1840 5035 1970 5065
rect 1800 5015 1970 5035
rect 2000 5135 2170 5155
rect 2000 5105 2010 5135
rect 2040 5105 2170 5135
rect 2000 5065 2170 5105
rect 2000 5035 2010 5065
rect 2040 5035 2170 5065
rect 2000 5015 2170 5035
rect 2200 5135 2370 5155
rect 2200 5105 2210 5135
rect 2240 5105 2370 5135
rect 2200 5065 2370 5105
rect 2200 5035 2210 5065
rect 2240 5035 2370 5065
rect 2200 5015 2370 5035
rect 2400 5135 2570 5155
rect 2400 5105 2410 5135
rect 2440 5105 2570 5135
rect 2400 5065 2570 5105
rect 2400 5035 2410 5065
rect 2440 5035 2570 5065
rect 2400 5015 2570 5035
rect 2600 5135 2770 5155
rect 2600 5105 2610 5135
rect 2640 5105 2770 5135
rect 2600 5065 2770 5105
rect 2600 5035 2610 5065
rect 2640 5035 2770 5065
rect 2600 5015 2770 5035
rect 2800 5135 2970 5155
rect 2800 5105 2810 5135
rect 2840 5105 2970 5135
rect 2800 5065 2970 5105
rect 2800 5035 2810 5065
rect 2840 5035 2970 5065
rect 2800 5015 2970 5035
rect 3000 5135 3170 5155
rect 3000 5105 3010 5135
rect 3040 5105 3170 5135
rect 3000 5065 3170 5105
rect 3000 5035 3010 5065
rect 3040 5035 3170 5065
rect 3000 5015 3170 5035
rect 3200 5135 3370 5155
rect 3200 5105 3210 5135
rect 3240 5105 3370 5135
rect 3200 5065 3370 5105
rect 3200 5035 3210 5065
rect 3240 5035 3370 5065
rect 3200 5015 3370 5035
rect 3400 5135 3570 5155
rect 3400 5105 3410 5135
rect 3440 5105 3570 5135
rect 3400 5065 3570 5105
rect 3400 5035 3410 5065
rect 3440 5035 3570 5065
rect 3400 5015 3570 5035
rect 3600 5135 3770 5155
rect 3600 5105 3610 5135
rect 3640 5105 3770 5135
rect 3600 5065 3770 5105
rect 3600 5035 3610 5065
rect 3640 5035 3770 5065
rect 3600 5015 3770 5035
rect 3800 5135 3970 5155
rect 3800 5105 3810 5135
rect 3840 5105 3970 5135
rect 3800 5065 3970 5105
rect 3800 5035 3810 5065
rect 3840 5035 3970 5065
rect 3800 5015 3970 5035
rect 4000 5135 4170 5155
rect 4000 5105 4010 5135
rect 4040 5105 4170 5135
rect 4000 5065 4170 5105
rect 4000 5035 4010 5065
rect 4040 5035 4170 5065
rect 4000 5015 4170 5035
rect 4200 5135 4370 5155
rect 4200 5105 4210 5135
rect 4240 5105 4370 5135
rect 4200 5065 4370 5105
rect 4200 5035 4210 5065
rect 4240 5035 4370 5065
rect 4200 5015 4370 5035
rect 4400 5135 4570 5155
rect 4400 5105 4410 5135
rect 4440 5105 4570 5135
rect 4400 5065 4570 5105
rect 4400 5035 4410 5065
rect 4440 5035 4570 5065
rect 4400 5015 4570 5035
rect 4600 5135 4770 5155
rect 4600 5105 4610 5135
rect 4640 5105 4770 5135
rect 4600 5065 4770 5105
rect 4600 5035 4610 5065
rect 4640 5035 4770 5065
rect 4600 5015 4770 5035
rect 4800 5135 4970 5155
rect 4800 5105 4810 5135
rect 4840 5105 4970 5135
rect 4800 5065 4970 5105
rect 4800 5035 4810 5065
rect 4840 5035 4970 5065
rect 4800 5015 4970 5035
rect 5000 5135 5170 5155
rect 5000 5105 5010 5135
rect 5040 5105 5170 5135
rect 5000 5065 5170 5105
rect 5000 5035 5010 5065
rect 5040 5035 5170 5065
rect 5000 5015 5170 5035
rect 5200 5135 5370 5155
rect 5200 5105 5210 5135
rect 5240 5105 5370 5135
rect 5200 5065 5370 5105
rect 5200 5035 5210 5065
rect 5240 5035 5370 5065
rect 5200 5015 5370 5035
rect 5400 5135 5570 5155
rect 5400 5105 5410 5135
rect 5440 5105 5570 5135
rect 5400 5065 5570 5105
rect 5400 5035 5410 5065
rect 5440 5035 5570 5065
rect 5400 5015 5570 5035
rect 5600 5135 5770 5155
rect 5600 5105 5610 5135
rect 5640 5105 5770 5135
rect 5600 5065 5770 5105
rect 5600 5035 5610 5065
rect 5640 5035 5770 5065
rect 5600 5015 5770 5035
rect 5800 5135 5970 5155
rect 5800 5105 5810 5135
rect 5840 5105 5970 5135
rect 5800 5065 5970 5105
rect 5800 5035 5810 5065
rect 5840 5035 5970 5065
rect 5800 5015 5970 5035
rect 6000 5135 6170 5155
rect 6000 5105 6010 5135
rect 6040 5105 6170 5135
rect 6000 5065 6170 5105
rect 6000 5035 6010 5065
rect 6040 5035 6170 5065
rect 6000 5015 6170 5035
rect 6200 5135 6370 5155
rect 6200 5105 6210 5135
rect 6240 5105 6370 5135
rect 6200 5065 6370 5105
rect 6200 5035 6210 5065
rect 6240 5035 6370 5065
rect 6200 5015 6370 5035
rect 6400 5135 6570 5155
rect 6400 5105 6410 5135
rect 6440 5105 6570 5135
rect 6400 5065 6570 5105
rect 6400 5035 6410 5065
rect 6440 5035 6570 5065
rect 6400 5015 6570 5035
rect -200 4950 -30 4970
rect -200 4920 -190 4950
rect -160 4920 -30 4950
rect -200 4880 -30 4920
rect -200 4850 -190 4880
rect -160 4850 -30 4880
rect -200 4830 -30 4850
rect 0 4950 170 4970
rect 0 4920 10 4950
rect 40 4920 170 4950
rect 0 4880 170 4920
rect 0 4850 10 4880
rect 40 4850 170 4880
rect 0 4830 170 4850
rect 200 4950 370 4970
rect 200 4920 210 4950
rect 240 4920 370 4950
rect 200 4880 370 4920
rect 200 4850 210 4880
rect 240 4850 370 4880
rect 200 4830 370 4850
rect 400 4950 570 4970
rect 400 4920 410 4950
rect 440 4920 570 4950
rect 400 4880 570 4920
rect 400 4850 410 4880
rect 440 4850 570 4880
rect 400 4830 570 4850
rect 600 4950 770 4970
rect 600 4920 610 4950
rect 640 4920 770 4950
rect 600 4880 770 4920
rect 600 4850 610 4880
rect 640 4850 770 4880
rect 600 4830 770 4850
rect 800 4950 970 4970
rect 800 4920 810 4950
rect 840 4920 970 4950
rect 800 4880 970 4920
rect 800 4850 810 4880
rect 840 4850 970 4880
rect 800 4830 970 4850
rect 1000 4950 1170 4970
rect 1000 4920 1010 4950
rect 1040 4920 1170 4950
rect 1000 4880 1170 4920
rect 1000 4850 1010 4880
rect 1040 4850 1170 4880
rect 1000 4830 1170 4850
rect 1200 4950 1370 4970
rect 1200 4920 1210 4950
rect 1240 4920 1370 4950
rect 1200 4880 1370 4920
rect 1200 4850 1210 4880
rect 1240 4850 1370 4880
rect 1200 4830 1370 4850
rect 1400 4950 1570 4970
rect 1400 4920 1410 4950
rect 1440 4920 1570 4950
rect 1400 4880 1570 4920
rect 1400 4850 1410 4880
rect 1440 4850 1570 4880
rect 1400 4830 1570 4850
rect 1600 4950 1770 4970
rect 1600 4920 1610 4950
rect 1640 4920 1770 4950
rect 1600 4880 1770 4920
rect 1600 4850 1610 4880
rect 1640 4850 1770 4880
rect 1600 4830 1770 4850
rect 1800 4950 1970 4970
rect 1800 4920 1810 4950
rect 1840 4920 1970 4950
rect 1800 4880 1970 4920
rect 1800 4850 1810 4880
rect 1840 4850 1970 4880
rect 1800 4830 1970 4850
rect 2000 4950 2170 4970
rect 2000 4920 2010 4950
rect 2040 4920 2170 4950
rect 2000 4880 2170 4920
rect 2000 4850 2010 4880
rect 2040 4850 2170 4880
rect 2000 4830 2170 4850
rect 2200 4950 2370 4970
rect 2200 4920 2210 4950
rect 2240 4920 2370 4950
rect 2200 4880 2370 4920
rect 2200 4850 2210 4880
rect 2240 4850 2370 4880
rect 2200 4830 2370 4850
rect 2400 4950 2570 4970
rect 2400 4920 2410 4950
rect 2440 4920 2570 4950
rect 2400 4880 2570 4920
rect 2400 4850 2410 4880
rect 2440 4850 2570 4880
rect 2400 4830 2570 4850
rect 2600 4950 2770 4970
rect 2600 4920 2610 4950
rect 2640 4920 2770 4950
rect 2600 4880 2770 4920
rect 2600 4850 2610 4880
rect 2640 4850 2770 4880
rect 2600 4830 2770 4850
rect 2800 4950 2970 4970
rect 2800 4920 2810 4950
rect 2840 4920 2970 4950
rect 2800 4880 2970 4920
rect 2800 4850 2810 4880
rect 2840 4850 2970 4880
rect 2800 4830 2970 4850
rect 3000 4950 3170 4970
rect 3000 4920 3010 4950
rect 3040 4920 3170 4950
rect 3000 4880 3170 4920
rect 3000 4850 3010 4880
rect 3040 4850 3170 4880
rect 3000 4830 3170 4850
rect 3200 4950 3370 4970
rect 3200 4920 3210 4950
rect 3240 4920 3370 4950
rect 3200 4880 3370 4920
rect 3200 4850 3210 4880
rect 3240 4850 3370 4880
rect 3200 4830 3370 4850
rect 3400 4950 3570 4970
rect 3400 4920 3410 4950
rect 3440 4920 3570 4950
rect 3400 4880 3570 4920
rect 3400 4850 3410 4880
rect 3440 4850 3570 4880
rect 3400 4830 3570 4850
rect 3600 4950 3770 4970
rect 3600 4920 3610 4950
rect 3640 4920 3770 4950
rect 3600 4880 3770 4920
rect 3600 4850 3610 4880
rect 3640 4850 3770 4880
rect 3600 4830 3770 4850
rect 3800 4950 3970 4970
rect 3800 4920 3810 4950
rect 3840 4920 3970 4950
rect 3800 4880 3970 4920
rect 3800 4850 3810 4880
rect 3840 4850 3970 4880
rect 3800 4830 3970 4850
rect 4000 4950 4170 4970
rect 4000 4920 4010 4950
rect 4040 4920 4170 4950
rect 4000 4880 4170 4920
rect 4000 4850 4010 4880
rect 4040 4850 4170 4880
rect 4000 4830 4170 4850
rect 4200 4950 4370 4970
rect 4200 4920 4210 4950
rect 4240 4920 4370 4950
rect 4200 4880 4370 4920
rect 4200 4850 4210 4880
rect 4240 4850 4370 4880
rect 4200 4830 4370 4850
rect 4400 4950 4570 4970
rect 4400 4920 4410 4950
rect 4440 4920 4570 4950
rect 4400 4880 4570 4920
rect 4400 4850 4410 4880
rect 4440 4850 4570 4880
rect 4400 4830 4570 4850
rect 4600 4950 4770 4970
rect 4600 4920 4610 4950
rect 4640 4920 4770 4950
rect 4600 4880 4770 4920
rect 4600 4850 4610 4880
rect 4640 4850 4770 4880
rect 4600 4830 4770 4850
rect 4800 4950 4970 4970
rect 4800 4920 4810 4950
rect 4840 4920 4970 4950
rect 4800 4880 4970 4920
rect 4800 4850 4810 4880
rect 4840 4850 4970 4880
rect 4800 4830 4970 4850
rect 5000 4950 5170 4970
rect 5000 4920 5010 4950
rect 5040 4920 5170 4950
rect 5000 4880 5170 4920
rect 5000 4850 5010 4880
rect 5040 4850 5170 4880
rect 5000 4830 5170 4850
rect 5200 4950 5370 4970
rect 5200 4920 5210 4950
rect 5240 4920 5370 4950
rect 5200 4880 5370 4920
rect 5200 4850 5210 4880
rect 5240 4850 5370 4880
rect 5200 4830 5370 4850
rect 5400 4950 5570 4970
rect 5400 4920 5410 4950
rect 5440 4920 5570 4950
rect 5400 4880 5570 4920
rect 5400 4850 5410 4880
rect 5440 4850 5570 4880
rect 5400 4830 5570 4850
rect 5600 4950 5770 4970
rect 5600 4920 5610 4950
rect 5640 4920 5770 4950
rect 5600 4880 5770 4920
rect 5600 4850 5610 4880
rect 5640 4850 5770 4880
rect 5600 4830 5770 4850
rect 5800 4950 5970 4970
rect 5800 4920 5810 4950
rect 5840 4920 5970 4950
rect 5800 4880 5970 4920
rect 5800 4850 5810 4880
rect 5840 4850 5970 4880
rect 5800 4830 5970 4850
rect 6000 4950 6170 4970
rect 6000 4920 6010 4950
rect 6040 4920 6170 4950
rect 6000 4880 6170 4920
rect 6000 4850 6010 4880
rect 6040 4850 6170 4880
rect 6000 4830 6170 4850
rect 6200 4950 6370 4970
rect 6200 4920 6210 4950
rect 6240 4920 6370 4950
rect 6200 4880 6370 4920
rect 6200 4850 6210 4880
rect 6240 4850 6370 4880
rect 6200 4830 6370 4850
rect 6400 4950 6570 4970
rect 6400 4920 6410 4950
rect 6440 4920 6570 4950
rect 6400 4880 6570 4920
rect 6400 4850 6410 4880
rect 6440 4850 6570 4880
rect 6400 4830 6570 4850
rect -200 4765 -30 4785
rect -200 4735 -190 4765
rect -160 4735 -30 4765
rect -200 4695 -30 4735
rect -200 4665 -190 4695
rect -160 4665 -30 4695
rect -200 4645 -30 4665
rect 0 4765 170 4785
rect 0 4735 10 4765
rect 40 4735 170 4765
rect 0 4695 170 4735
rect 0 4665 10 4695
rect 40 4665 170 4695
rect 0 4645 170 4665
rect 200 4765 370 4785
rect 200 4735 210 4765
rect 240 4735 370 4765
rect 200 4695 370 4735
rect 200 4665 210 4695
rect 240 4665 370 4695
rect 200 4645 370 4665
rect 400 4765 570 4785
rect 400 4735 410 4765
rect 440 4735 570 4765
rect 400 4695 570 4735
rect 400 4665 410 4695
rect 440 4665 570 4695
rect 400 4645 570 4665
rect 600 4765 770 4785
rect 600 4735 610 4765
rect 640 4735 770 4765
rect 600 4695 770 4735
rect 600 4665 610 4695
rect 640 4665 770 4695
rect 600 4645 770 4665
rect 800 4765 970 4785
rect 800 4735 810 4765
rect 840 4735 970 4765
rect 800 4695 970 4735
rect 800 4665 810 4695
rect 840 4665 970 4695
rect 800 4645 970 4665
rect 1000 4765 1170 4785
rect 1000 4735 1010 4765
rect 1040 4735 1170 4765
rect 1000 4695 1170 4735
rect 1000 4665 1010 4695
rect 1040 4665 1170 4695
rect 1000 4645 1170 4665
rect 1200 4765 1370 4785
rect 1200 4735 1210 4765
rect 1240 4735 1370 4765
rect 1200 4695 1370 4735
rect 1200 4665 1210 4695
rect 1240 4665 1370 4695
rect 1200 4645 1370 4665
rect 1400 4765 1570 4785
rect 1400 4735 1410 4765
rect 1440 4735 1570 4765
rect 1400 4695 1570 4735
rect 1400 4665 1410 4695
rect 1440 4665 1570 4695
rect 1400 4645 1570 4665
rect 1600 4765 1770 4785
rect 1600 4735 1610 4765
rect 1640 4735 1770 4765
rect 1600 4695 1770 4735
rect 1600 4665 1610 4695
rect 1640 4665 1770 4695
rect 1600 4645 1770 4665
rect 1800 4765 1970 4785
rect 1800 4735 1810 4765
rect 1840 4735 1970 4765
rect 1800 4695 1970 4735
rect 1800 4665 1810 4695
rect 1840 4665 1970 4695
rect 1800 4645 1970 4665
rect 2000 4765 2170 4785
rect 2000 4735 2010 4765
rect 2040 4735 2170 4765
rect 2000 4695 2170 4735
rect 2000 4665 2010 4695
rect 2040 4665 2170 4695
rect 2000 4645 2170 4665
rect 2200 4765 2370 4785
rect 2200 4735 2210 4765
rect 2240 4735 2370 4765
rect 2200 4695 2370 4735
rect 2200 4665 2210 4695
rect 2240 4665 2370 4695
rect 2200 4645 2370 4665
rect 2400 4765 2570 4785
rect 2400 4735 2410 4765
rect 2440 4735 2570 4765
rect 2400 4695 2570 4735
rect 2400 4665 2410 4695
rect 2440 4665 2570 4695
rect 2400 4645 2570 4665
rect 2600 4765 2770 4785
rect 2600 4735 2610 4765
rect 2640 4735 2770 4765
rect 2600 4695 2770 4735
rect 2600 4665 2610 4695
rect 2640 4665 2770 4695
rect 2600 4645 2770 4665
rect 2800 4765 2970 4785
rect 2800 4735 2810 4765
rect 2840 4735 2970 4765
rect 2800 4695 2970 4735
rect 2800 4665 2810 4695
rect 2840 4665 2970 4695
rect 2800 4645 2970 4665
rect 3000 4765 3170 4785
rect 3000 4735 3010 4765
rect 3040 4735 3170 4765
rect 3000 4695 3170 4735
rect 3000 4665 3010 4695
rect 3040 4665 3170 4695
rect 3000 4645 3170 4665
rect 3200 4765 3370 4785
rect 3200 4735 3210 4765
rect 3240 4735 3370 4765
rect 3200 4695 3370 4735
rect 3200 4665 3210 4695
rect 3240 4665 3370 4695
rect 3200 4645 3370 4665
rect 3400 4765 3570 4785
rect 3400 4735 3410 4765
rect 3440 4735 3570 4765
rect 3400 4695 3570 4735
rect 3400 4665 3410 4695
rect 3440 4665 3570 4695
rect 3400 4645 3570 4665
rect 3600 4765 3770 4785
rect 3600 4735 3610 4765
rect 3640 4735 3770 4765
rect 3600 4695 3770 4735
rect 3600 4665 3610 4695
rect 3640 4665 3770 4695
rect 3600 4645 3770 4665
rect 3800 4765 3970 4785
rect 3800 4735 3810 4765
rect 3840 4735 3970 4765
rect 3800 4695 3970 4735
rect 3800 4665 3810 4695
rect 3840 4665 3970 4695
rect 3800 4645 3970 4665
rect 4000 4765 4170 4785
rect 4000 4735 4010 4765
rect 4040 4735 4170 4765
rect 4000 4695 4170 4735
rect 4000 4665 4010 4695
rect 4040 4665 4170 4695
rect 4000 4645 4170 4665
rect 4200 4765 4370 4785
rect 4200 4735 4210 4765
rect 4240 4735 4370 4765
rect 4200 4695 4370 4735
rect 4200 4665 4210 4695
rect 4240 4665 4370 4695
rect 4200 4645 4370 4665
rect 4400 4765 4570 4785
rect 4400 4735 4410 4765
rect 4440 4735 4570 4765
rect 4400 4695 4570 4735
rect 4400 4665 4410 4695
rect 4440 4665 4570 4695
rect 4400 4645 4570 4665
rect 4600 4765 4770 4785
rect 4600 4735 4610 4765
rect 4640 4735 4770 4765
rect 4600 4695 4770 4735
rect 4600 4665 4610 4695
rect 4640 4665 4770 4695
rect 4600 4645 4770 4665
rect 4800 4765 4970 4785
rect 4800 4735 4810 4765
rect 4840 4735 4970 4765
rect 4800 4695 4970 4735
rect 4800 4665 4810 4695
rect 4840 4665 4970 4695
rect 4800 4645 4970 4665
rect 5000 4765 5170 4785
rect 5000 4735 5010 4765
rect 5040 4735 5170 4765
rect 5000 4695 5170 4735
rect 5000 4665 5010 4695
rect 5040 4665 5170 4695
rect 5000 4645 5170 4665
rect 5200 4765 5370 4785
rect 5200 4735 5210 4765
rect 5240 4735 5370 4765
rect 5200 4695 5370 4735
rect 5200 4665 5210 4695
rect 5240 4665 5370 4695
rect 5200 4645 5370 4665
rect 5400 4765 5570 4785
rect 5400 4735 5410 4765
rect 5440 4735 5570 4765
rect 5400 4695 5570 4735
rect 5400 4665 5410 4695
rect 5440 4665 5570 4695
rect 5400 4645 5570 4665
rect 5600 4765 5770 4785
rect 5600 4735 5610 4765
rect 5640 4735 5770 4765
rect 5600 4695 5770 4735
rect 5600 4665 5610 4695
rect 5640 4665 5770 4695
rect 5600 4645 5770 4665
rect 5800 4765 5970 4785
rect 5800 4735 5810 4765
rect 5840 4735 5970 4765
rect 5800 4695 5970 4735
rect 5800 4665 5810 4695
rect 5840 4665 5970 4695
rect 5800 4645 5970 4665
rect 6000 4765 6170 4785
rect 6000 4735 6010 4765
rect 6040 4735 6170 4765
rect 6000 4695 6170 4735
rect 6000 4665 6010 4695
rect 6040 4665 6170 4695
rect 6000 4645 6170 4665
rect 6200 4765 6370 4785
rect 6200 4735 6210 4765
rect 6240 4735 6370 4765
rect 6200 4695 6370 4735
rect 6200 4665 6210 4695
rect 6240 4665 6370 4695
rect 6200 4645 6370 4665
rect 6400 4765 6570 4785
rect 6400 4735 6410 4765
rect 6440 4735 6570 4765
rect 6400 4695 6570 4735
rect 6400 4665 6410 4695
rect 6440 4665 6570 4695
rect 6400 4645 6570 4665
rect -200 4580 -30 4600
rect -200 4550 -190 4580
rect -160 4550 -30 4580
rect -200 4510 -30 4550
rect -200 4480 -190 4510
rect -160 4480 -30 4510
rect -200 4460 -30 4480
rect 0 4580 170 4600
rect 0 4550 10 4580
rect 40 4550 170 4580
rect 0 4510 170 4550
rect 0 4480 10 4510
rect 40 4480 170 4510
rect 0 4460 170 4480
rect 200 4580 370 4600
rect 200 4550 210 4580
rect 240 4550 370 4580
rect 200 4510 370 4550
rect 200 4480 210 4510
rect 240 4480 370 4510
rect 200 4460 370 4480
rect 400 4580 570 4600
rect 400 4550 410 4580
rect 440 4550 570 4580
rect 400 4510 570 4550
rect 400 4480 410 4510
rect 440 4480 570 4510
rect 400 4460 570 4480
rect 600 4580 770 4600
rect 600 4550 610 4580
rect 640 4550 770 4580
rect 600 4510 770 4550
rect 600 4480 610 4510
rect 640 4480 770 4510
rect 600 4460 770 4480
rect 800 4580 970 4600
rect 800 4550 810 4580
rect 840 4550 970 4580
rect 800 4510 970 4550
rect 800 4480 810 4510
rect 840 4480 970 4510
rect 800 4460 970 4480
rect 1000 4580 1170 4600
rect 1000 4550 1010 4580
rect 1040 4550 1170 4580
rect 1000 4510 1170 4550
rect 1000 4480 1010 4510
rect 1040 4480 1170 4510
rect 1000 4460 1170 4480
rect 1200 4580 1370 4600
rect 1200 4550 1210 4580
rect 1240 4550 1370 4580
rect 1200 4510 1370 4550
rect 1200 4480 1210 4510
rect 1240 4480 1370 4510
rect 1200 4460 1370 4480
rect 1400 4580 1570 4600
rect 1400 4550 1410 4580
rect 1440 4550 1570 4580
rect 1400 4510 1570 4550
rect 1400 4480 1410 4510
rect 1440 4480 1570 4510
rect 1400 4460 1570 4480
rect 1600 4580 1770 4600
rect 1600 4550 1610 4580
rect 1640 4550 1770 4580
rect 1600 4510 1770 4550
rect 1600 4480 1610 4510
rect 1640 4480 1770 4510
rect 1600 4460 1770 4480
rect 1800 4580 1970 4600
rect 1800 4550 1810 4580
rect 1840 4550 1970 4580
rect 1800 4510 1970 4550
rect 1800 4480 1810 4510
rect 1840 4480 1970 4510
rect 1800 4460 1970 4480
rect 2000 4580 2170 4600
rect 2000 4550 2010 4580
rect 2040 4550 2170 4580
rect 2000 4510 2170 4550
rect 2000 4480 2010 4510
rect 2040 4480 2170 4510
rect 2000 4460 2170 4480
rect 2200 4580 2370 4600
rect 2200 4550 2210 4580
rect 2240 4550 2370 4580
rect 2200 4510 2370 4550
rect 2200 4480 2210 4510
rect 2240 4480 2370 4510
rect 2200 4460 2370 4480
rect 2400 4580 2570 4600
rect 2400 4550 2410 4580
rect 2440 4550 2570 4580
rect 2400 4510 2570 4550
rect 2400 4480 2410 4510
rect 2440 4480 2570 4510
rect 2400 4460 2570 4480
rect 2600 4580 2770 4600
rect 2600 4550 2610 4580
rect 2640 4550 2770 4580
rect 2600 4510 2770 4550
rect 2600 4480 2610 4510
rect 2640 4480 2770 4510
rect 2600 4460 2770 4480
rect 2800 4580 2970 4600
rect 2800 4550 2810 4580
rect 2840 4550 2970 4580
rect 2800 4510 2970 4550
rect 2800 4480 2810 4510
rect 2840 4480 2970 4510
rect 2800 4460 2970 4480
rect 3000 4580 3170 4600
rect 3000 4550 3010 4580
rect 3040 4550 3170 4580
rect 3000 4510 3170 4550
rect 3000 4480 3010 4510
rect 3040 4480 3170 4510
rect 3000 4460 3170 4480
rect 3200 4580 3370 4600
rect 3200 4550 3210 4580
rect 3240 4550 3370 4580
rect 3200 4510 3370 4550
rect 3200 4480 3210 4510
rect 3240 4480 3370 4510
rect 3200 4460 3370 4480
rect 3400 4580 3570 4600
rect 3400 4550 3410 4580
rect 3440 4550 3570 4580
rect 3400 4510 3570 4550
rect 3400 4480 3410 4510
rect 3440 4480 3570 4510
rect 3400 4460 3570 4480
rect 3600 4580 3770 4600
rect 3600 4550 3610 4580
rect 3640 4550 3770 4580
rect 3600 4510 3770 4550
rect 3600 4480 3610 4510
rect 3640 4480 3770 4510
rect 3600 4460 3770 4480
rect 3800 4580 3970 4600
rect 3800 4550 3810 4580
rect 3840 4550 3970 4580
rect 3800 4510 3970 4550
rect 3800 4480 3810 4510
rect 3840 4480 3970 4510
rect 3800 4460 3970 4480
rect 4000 4580 4170 4600
rect 4000 4550 4010 4580
rect 4040 4550 4170 4580
rect 4000 4510 4170 4550
rect 4000 4480 4010 4510
rect 4040 4480 4170 4510
rect 4000 4460 4170 4480
rect 4200 4580 4370 4600
rect 4200 4550 4210 4580
rect 4240 4550 4370 4580
rect 4200 4510 4370 4550
rect 4200 4480 4210 4510
rect 4240 4480 4370 4510
rect 4200 4460 4370 4480
rect 4400 4580 4570 4600
rect 4400 4550 4410 4580
rect 4440 4550 4570 4580
rect 4400 4510 4570 4550
rect 4400 4480 4410 4510
rect 4440 4480 4570 4510
rect 4400 4460 4570 4480
rect 4600 4580 4770 4600
rect 4600 4550 4610 4580
rect 4640 4550 4770 4580
rect 4600 4510 4770 4550
rect 4600 4480 4610 4510
rect 4640 4480 4770 4510
rect 4600 4460 4770 4480
rect 4800 4580 4970 4600
rect 4800 4550 4810 4580
rect 4840 4550 4970 4580
rect 4800 4510 4970 4550
rect 4800 4480 4810 4510
rect 4840 4480 4970 4510
rect 4800 4460 4970 4480
rect 5000 4580 5170 4600
rect 5000 4550 5010 4580
rect 5040 4550 5170 4580
rect 5000 4510 5170 4550
rect 5000 4480 5010 4510
rect 5040 4480 5170 4510
rect 5000 4460 5170 4480
rect 5200 4580 5370 4600
rect 5200 4550 5210 4580
rect 5240 4550 5370 4580
rect 5200 4510 5370 4550
rect 5200 4480 5210 4510
rect 5240 4480 5370 4510
rect 5200 4460 5370 4480
rect 5400 4580 5570 4600
rect 5400 4550 5410 4580
rect 5440 4550 5570 4580
rect 5400 4510 5570 4550
rect 5400 4480 5410 4510
rect 5440 4480 5570 4510
rect 5400 4460 5570 4480
rect 5600 4580 5770 4600
rect 5600 4550 5610 4580
rect 5640 4550 5770 4580
rect 5600 4510 5770 4550
rect 5600 4480 5610 4510
rect 5640 4480 5770 4510
rect 5600 4460 5770 4480
rect 5800 4580 5970 4600
rect 5800 4550 5810 4580
rect 5840 4550 5970 4580
rect 5800 4510 5970 4550
rect 5800 4480 5810 4510
rect 5840 4480 5970 4510
rect 5800 4460 5970 4480
rect 6000 4580 6170 4600
rect 6000 4550 6010 4580
rect 6040 4550 6170 4580
rect 6000 4510 6170 4550
rect 6000 4480 6010 4510
rect 6040 4480 6170 4510
rect 6000 4460 6170 4480
rect 6200 4580 6370 4600
rect 6200 4550 6210 4580
rect 6240 4550 6370 4580
rect 6200 4510 6370 4550
rect 6200 4480 6210 4510
rect 6240 4480 6370 4510
rect 6200 4460 6370 4480
rect 6400 4580 6570 4600
rect 6400 4550 6410 4580
rect 6440 4550 6570 4580
rect 6400 4510 6570 4550
rect 6400 4480 6410 4510
rect 6440 4480 6570 4510
rect 6400 4460 6570 4480
rect -200 4395 -30 4415
rect -200 4365 -190 4395
rect -160 4365 -30 4395
rect -200 4325 -30 4365
rect -200 4295 -190 4325
rect -160 4295 -30 4325
rect -200 4275 -30 4295
rect 0 4395 170 4415
rect 0 4365 10 4395
rect 40 4365 170 4395
rect 0 4325 170 4365
rect 0 4295 10 4325
rect 40 4295 170 4325
rect 0 4275 170 4295
rect 200 4395 370 4415
rect 200 4365 210 4395
rect 240 4365 370 4395
rect 200 4325 370 4365
rect 200 4295 210 4325
rect 240 4295 370 4325
rect 200 4275 370 4295
rect 400 4395 570 4415
rect 400 4365 410 4395
rect 440 4365 570 4395
rect 400 4325 570 4365
rect 400 4295 410 4325
rect 440 4295 570 4325
rect 400 4275 570 4295
rect 600 4395 770 4415
rect 600 4365 610 4395
rect 640 4365 770 4395
rect 600 4325 770 4365
rect 600 4295 610 4325
rect 640 4295 770 4325
rect 600 4275 770 4295
rect 800 4395 970 4415
rect 800 4365 810 4395
rect 840 4365 970 4395
rect 800 4325 970 4365
rect 800 4295 810 4325
rect 840 4295 970 4325
rect 800 4275 970 4295
rect 1000 4395 1170 4415
rect 1000 4365 1010 4395
rect 1040 4365 1170 4395
rect 1000 4325 1170 4365
rect 1000 4295 1010 4325
rect 1040 4295 1170 4325
rect 1000 4275 1170 4295
rect 1200 4395 1370 4415
rect 1200 4365 1210 4395
rect 1240 4365 1370 4395
rect 1200 4325 1370 4365
rect 1200 4295 1210 4325
rect 1240 4295 1370 4325
rect 1200 4275 1370 4295
rect 1400 4395 1570 4415
rect 1400 4365 1410 4395
rect 1440 4365 1570 4395
rect 1400 4325 1570 4365
rect 1400 4295 1410 4325
rect 1440 4295 1570 4325
rect 1400 4275 1570 4295
rect 1600 4395 1770 4415
rect 1600 4365 1610 4395
rect 1640 4365 1770 4395
rect 1600 4325 1770 4365
rect 1600 4295 1610 4325
rect 1640 4295 1770 4325
rect 1600 4275 1770 4295
rect 1800 4395 1970 4415
rect 1800 4365 1810 4395
rect 1840 4365 1970 4395
rect 1800 4325 1970 4365
rect 1800 4295 1810 4325
rect 1840 4295 1970 4325
rect 1800 4275 1970 4295
rect 2000 4395 2170 4415
rect 2000 4365 2010 4395
rect 2040 4365 2170 4395
rect 2000 4325 2170 4365
rect 2000 4295 2010 4325
rect 2040 4295 2170 4325
rect 2000 4275 2170 4295
rect 2200 4395 2370 4415
rect 2200 4365 2210 4395
rect 2240 4365 2370 4395
rect 2200 4325 2370 4365
rect 2200 4295 2210 4325
rect 2240 4295 2370 4325
rect 2200 4275 2370 4295
rect 2400 4395 2570 4415
rect 2400 4365 2410 4395
rect 2440 4365 2570 4395
rect 2400 4325 2570 4365
rect 2400 4295 2410 4325
rect 2440 4295 2570 4325
rect 2400 4275 2570 4295
rect 2600 4395 2770 4415
rect 2600 4365 2610 4395
rect 2640 4365 2770 4395
rect 2600 4325 2770 4365
rect 2600 4295 2610 4325
rect 2640 4295 2770 4325
rect 2600 4275 2770 4295
rect 2800 4395 2970 4415
rect 2800 4365 2810 4395
rect 2840 4365 2970 4395
rect 2800 4325 2970 4365
rect 2800 4295 2810 4325
rect 2840 4295 2970 4325
rect 2800 4275 2970 4295
rect 3000 4395 3170 4415
rect 3000 4365 3010 4395
rect 3040 4365 3170 4395
rect 3000 4325 3170 4365
rect 3000 4295 3010 4325
rect 3040 4295 3170 4325
rect 3000 4275 3170 4295
rect 3200 4395 3370 4415
rect 3200 4365 3210 4395
rect 3240 4365 3370 4395
rect 3200 4325 3370 4365
rect 3200 4295 3210 4325
rect 3240 4295 3370 4325
rect 3200 4275 3370 4295
rect 3400 4395 3570 4415
rect 3400 4365 3410 4395
rect 3440 4365 3570 4395
rect 3400 4325 3570 4365
rect 3400 4295 3410 4325
rect 3440 4295 3570 4325
rect 3400 4275 3570 4295
rect 3600 4395 3770 4415
rect 3600 4365 3610 4395
rect 3640 4365 3770 4395
rect 3600 4325 3770 4365
rect 3600 4295 3610 4325
rect 3640 4295 3770 4325
rect 3600 4275 3770 4295
rect 3800 4395 3970 4415
rect 3800 4365 3810 4395
rect 3840 4365 3970 4395
rect 3800 4325 3970 4365
rect 3800 4295 3810 4325
rect 3840 4295 3970 4325
rect 3800 4275 3970 4295
rect 4000 4395 4170 4415
rect 4000 4365 4010 4395
rect 4040 4365 4170 4395
rect 4000 4325 4170 4365
rect 4000 4295 4010 4325
rect 4040 4295 4170 4325
rect 4000 4275 4170 4295
rect 4200 4395 4370 4415
rect 4200 4365 4210 4395
rect 4240 4365 4370 4395
rect 4200 4325 4370 4365
rect 4200 4295 4210 4325
rect 4240 4295 4370 4325
rect 4200 4275 4370 4295
rect 4400 4395 4570 4415
rect 4400 4365 4410 4395
rect 4440 4365 4570 4395
rect 4400 4325 4570 4365
rect 4400 4295 4410 4325
rect 4440 4295 4570 4325
rect 4400 4275 4570 4295
rect 4600 4395 4770 4415
rect 4600 4365 4610 4395
rect 4640 4365 4770 4395
rect 4600 4325 4770 4365
rect 4600 4295 4610 4325
rect 4640 4295 4770 4325
rect 4600 4275 4770 4295
rect 4800 4395 4970 4415
rect 4800 4365 4810 4395
rect 4840 4365 4970 4395
rect 4800 4325 4970 4365
rect 4800 4295 4810 4325
rect 4840 4295 4970 4325
rect 4800 4275 4970 4295
rect 5000 4395 5170 4415
rect 5000 4365 5010 4395
rect 5040 4365 5170 4395
rect 5000 4325 5170 4365
rect 5000 4295 5010 4325
rect 5040 4295 5170 4325
rect 5000 4275 5170 4295
rect 5200 4395 5370 4415
rect 5200 4365 5210 4395
rect 5240 4365 5370 4395
rect 5200 4325 5370 4365
rect 5200 4295 5210 4325
rect 5240 4295 5370 4325
rect 5200 4275 5370 4295
rect 5400 4395 5570 4415
rect 5400 4365 5410 4395
rect 5440 4365 5570 4395
rect 5400 4325 5570 4365
rect 5400 4295 5410 4325
rect 5440 4295 5570 4325
rect 5400 4275 5570 4295
rect 5600 4395 5770 4415
rect 5600 4365 5610 4395
rect 5640 4365 5770 4395
rect 5600 4325 5770 4365
rect 5600 4295 5610 4325
rect 5640 4295 5770 4325
rect 5600 4275 5770 4295
rect 5800 4395 5970 4415
rect 5800 4365 5810 4395
rect 5840 4365 5970 4395
rect 5800 4325 5970 4365
rect 5800 4295 5810 4325
rect 5840 4295 5970 4325
rect 5800 4275 5970 4295
rect 6000 4395 6170 4415
rect 6000 4365 6010 4395
rect 6040 4365 6170 4395
rect 6000 4325 6170 4365
rect 6000 4295 6010 4325
rect 6040 4295 6170 4325
rect 6000 4275 6170 4295
rect 6200 4395 6370 4415
rect 6200 4365 6210 4395
rect 6240 4365 6370 4395
rect 6200 4325 6370 4365
rect 6200 4295 6210 4325
rect 6240 4295 6370 4325
rect 6200 4275 6370 4295
rect 6400 4395 6570 4415
rect 6400 4365 6410 4395
rect 6440 4365 6570 4395
rect 6400 4325 6570 4365
rect 6400 4295 6410 4325
rect 6440 4295 6570 4325
rect 6400 4275 6570 4295
rect -200 4210 -30 4230
rect -200 4180 -190 4210
rect -160 4180 -30 4210
rect -200 4140 -30 4180
rect -200 4110 -190 4140
rect -160 4110 -30 4140
rect -200 4090 -30 4110
rect 0 4210 170 4230
rect 0 4180 10 4210
rect 40 4180 170 4210
rect 0 4140 170 4180
rect 0 4110 10 4140
rect 40 4110 170 4140
rect 0 4090 170 4110
rect 200 4210 370 4230
rect 200 4180 210 4210
rect 240 4180 370 4210
rect 200 4140 370 4180
rect 200 4110 210 4140
rect 240 4110 370 4140
rect 200 4090 370 4110
rect 400 4210 570 4230
rect 400 4180 410 4210
rect 440 4180 570 4210
rect 400 4140 570 4180
rect 400 4110 410 4140
rect 440 4110 570 4140
rect 400 4090 570 4110
rect 600 4210 770 4230
rect 600 4180 610 4210
rect 640 4180 770 4210
rect 600 4140 770 4180
rect 600 4110 610 4140
rect 640 4110 770 4140
rect 600 4090 770 4110
rect 800 4210 970 4230
rect 800 4180 810 4210
rect 840 4180 970 4210
rect 800 4140 970 4180
rect 800 4110 810 4140
rect 840 4110 970 4140
rect 800 4090 970 4110
rect 1000 4210 1170 4230
rect 1000 4180 1010 4210
rect 1040 4180 1170 4210
rect 1000 4140 1170 4180
rect 1000 4110 1010 4140
rect 1040 4110 1170 4140
rect 1000 4090 1170 4110
rect 1200 4210 1370 4230
rect 1200 4180 1210 4210
rect 1240 4180 1370 4210
rect 1200 4140 1370 4180
rect 1200 4110 1210 4140
rect 1240 4110 1370 4140
rect 1200 4090 1370 4110
rect 1400 4210 1570 4230
rect 1400 4180 1410 4210
rect 1440 4180 1570 4210
rect 1400 4140 1570 4180
rect 1400 4110 1410 4140
rect 1440 4110 1570 4140
rect 1400 4090 1570 4110
rect 1600 4210 1770 4230
rect 1600 4180 1610 4210
rect 1640 4180 1770 4210
rect 1600 4140 1770 4180
rect 1600 4110 1610 4140
rect 1640 4110 1770 4140
rect 1600 4090 1770 4110
rect 1800 4210 1970 4230
rect 1800 4180 1810 4210
rect 1840 4180 1970 4210
rect 1800 4140 1970 4180
rect 1800 4110 1810 4140
rect 1840 4110 1970 4140
rect 1800 4090 1970 4110
rect 2000 4210 2170 4230
rect 2000 4180 2010 4210
rect 2040 4180 2170 4210
rect 2000 4140 2170 4180
rect 2000 4110 2010 4140
rect 2040 4110 2170 4140
rect 2000 4090 2170 4110
rect 2200 4210 2370 4230
rect 2200 4180 2210 4210
rect 2240 4180 2370 4210
rect 2200 4140 2370 4180
rect 2200 4110 2210 4140
rect 2240 4110 2370 4140
rect 2200 4090 2370 4110
rect 2400 4210 2570 4230
rect 2400 4180 2410 4210
rect 2440 4180 2570 4210
rect 2400 4140 2570 4180
rect 2400 4110 2410 4140
rect 2440 4110 2570 4140
rect 2400 4090 2570 4110
rect 2600 4210 2770 4230
rect 2600 4180 2610 4210
rect 2640 4180 2770 4210
rect 2600 4140 2770 4180
rect 2600 4110 2610 4140
rect 2640 4110 2770 4140
rect 2600 4090 2770 4110
rect 2800 4210 2970 4230
rect 2800 4180 2810 4210
rect 2840 4180 2970 4210
rect 2800 4140 2970 4180
rect 2800 4110 2810 4140
rect 2840 4110 2970 4140
rect 2800 4090 2970 4110
rect 3000 4210 3170 4230
rect 3000 4180 3010 4210
rect 3040 4180 3170 4210
rect 3000 4140 3170 4180
rect 3000 4110 3010 4140
rect 3040 4110 3170 4140
rect 3000 4090 3170 4110
rect 3200 4210 3370 4230
rect 3200 4180 3210 4210
rect 3240 4180 3370 4210
rect 3200 4140 3370 4180
rect 3200 4110 3210 4140
rect 3240 4110 3370 4140
rect 3200 4090 3370 4110
rect 3400 4210 3570 4230
rect 3400 4180 3410 4210
rect 3440 4180 3570 4210
rect 3400 4140 3570 4180
rect 3400 4110 3410 4140
rect 3440 4110 3570 4140
rect 3400 4090 3570 4110
rect 3600 4210 3770 4230
rect 3600 4180 3610 4210
rect 3640 4180 3770 4210
rect 3600 4140 3770 4180
rect 3600 4110 3610 4140
rect 3640 4110 3770 4140
rect 3600 4090 3770 4110
rect 3800 4210 3970 4230
rect 3800 4180 3810 4210
rect 3840 4180 3970 4210
rect 3800 4140 3970 4180
rect 3800 4110 3810 4140
rect 3840 4110 3970 4140
rect 3800 4090 3970 4110
rect 4000 4210 4170 4230
rect 4000 4180 4010 4210
rect 4040 4180 4170 4210
rect 4000 4140 4170 4180
rect 4000 4110 4010 4140
rect 4040 4110 4170 4140
rect 4000 4090 4170 4110
rect 4200 4210 4370 4230
rect 4200 4180 4210 4210
rect 4240 4180 4370 4210
rect 4200 4140 4370 4180
rect 4200 4110 4210 4140
rect 4240 4110 4370 4140
rect 4200 4090 4370 4110
rect 4400 4210 4570 4230
rect 4400 4180 4410 4210
rect 4440 4180 4570 4210
rect 4400 4140 4570 4180
rect 4400 4110 4410 4140
rect 4440 4110 4570 4140
rect 4400 4090 4570 4110
rect 4600 4210 4770 4230
rect 4600 4180 4610 4210
rect 4640 4180 4770 4210
rect 4600 4140 4770 4180
rect 4600 4110 4610 4140
rect 4640 4110 4770 4140
rect 4600 4090 4770 4110
rect 4800 4210 4970 4230
rect 4800 4180 4810 4210
rect 4840 4180 4970 4210
rect 4800 4140 4970 4180
rect 4800 4110 4810 4140
rect 4840 4110 4970 4140
rect 4800 4090 4970 4110
rect 5000 4210 5170 4230
rect 5000 4180 5010 4210
rect 5040 4180 5170 4210
rect 5000 4140 5170 4180
rect 5000 4110 5010 4140
rect 5040 4110 5170 4140
rect 5000 4090 5170 4110
rect 5200 4210 5370 4230
rect 5200 4180 5210 4210
rect 5240 4180 5370 4210
rect 5200 4140 5370 4180
rect 5200 4110 5210 4140
rect 5240 4110 5370 4140
rect 5200 4090 5370 4110
rect 5400 4210 5570 4230
rect 5400 4180 5410 4210
rect 5440 4180 5570 4210
rect 5400 4140 5570 4180
rect 5400 4110 5410 4140
rect 5440 4110 5570 4140
rect 5400 4090 5570 4110
rect 5600 4210 5770 4230
rect 5600 4180 5610 4210
rect 5640 4180 5770 4210
rect 5600 4140 5770 4180
rect 5600 4110 5610 4140
rect 5640 4110 5770 4140
rect 5600 4090 5770 4110
rect 5800 4210 5970 4230
rect 5800 4180 5810 4210
rect 5840 4180 5970 4210
rect 5800 4140 5970 4180
rect 5800 4110 5810 4140
rect 5840 4110 5970 4140
rect 5800 4090 5970 4110
rect 6000 4210 6170 4230
rect 6000 4180 6010 4210
rect 6040 4180 6170 4210
rect 6000 4140 6170 4180
rect 6000 4110 6010 4140
rect 6040 4110 6170 4140
rect 6000 4090 6170 4110
rect 6200 4210 6370 4230
rect 6200 4180 6210 4210
rect 6240 4180 6370 4210
rect 6200 4140 6370 4180
rect 6200 4110 6210 4140
rect 6240 4110 6370 4140
rect 6200 4090 6370 4110
rect 6400 4210 6570 4230
rect 6400 4180 6410 4210
rect 6440 4180 6570 4210
rect 6400 4140 6570 4180
rect 6400 4110 6410 4140
rect 6440 4110 6570 4140
rect 6400 4090 6570 4110
rect -200 4025 -30 4045
rect -200 3995 -190 4025
rect -160 3995 -30 4025
rect -200 3955 -30 3995
rect -200 3925 -190 3955
rect -160 3925 -30 3955
rect -200 3905 -30 3925
rect 0 4025 170 4045
rect 0 3995 10 4025
rect 40 3995 170 4025
rect 0 3955 170 3995
rect 0 3925 10 3955
rect 40 3925 170 3955
rect 0 3905 170 3925
rect 200 4025 370 4045
rect 200 3995 210 4025
rect 240 3995 370 4025
rect 200 3955 370 3995
rect 200 3925 210 3955
rect 240 3925 370 3955
rect 200 3905 370 3925
rect 400 4025 570 4045
rect 400 3995 410 4025
rect 440 3995 570 4025
rect 400 3955 570 3995
rect 400 3925 410 3955
rect 440 3925 570 3955
rect 400 3905 570 3925
rect 600 4025 770 4045
rect 600 3995 610 4025
rect 640 3995 770 4025
rect 600 3955 770 3995
rect 600 3925 610 3955
rect 640 3925 770 3955
rect 600 3905 770 3925
rect 800 4025 970 4045
rect 800 3995 810 4025
rect 840 3995 970 4025
rect 800 3955 970 3995
rect 800 3925 810 3955
rect 840 3925 970 3955
rect 800 3905 970 3925
rect 1000 4025 1170 4045
rect 1000 3995 1010 4025
rect 1040 3995 1170 4025
rect 1000 3955 1170 3995
rect 1000 3925 1010 3955
rect 1040 3925 1170 3955
rect 1000 3905 1170 3925
rect 1200 4025 1370 4045
rect 1200 3995 1210 4025
rect 1240 3995 1370 4025
rect 1200 3955 1370 3995
rect 1200 3925 1210 3955
rect 1240 3925 1370 3955
rect 1200 3905 1370 3925
rect 1400 4025 1570 4045
rect 1400 3995 1410 4025
rect 1440 3995 1570 4025
rect 1400 3955 1570 3995
rect 1400 3925 1410 3955
rect 1440 3925 1570 3955
rect 1400 3905 1570 3925
rect 1600 4025 1770 4045
rect 1600 3995 1610 4025
rect 1640 3995 1770 4025
rect 1600 3955 1770 3995
rect 1600 3925 1610 3955
rect 1640 3925 1770 3955
rect 1600 3905 1770 3925
rect 1800 4025 1970 4045
rect 1800 3995 1810 4025
rect 1840 3995 1970 4025
rect 1800 3955 1970 3995
rect 1800 3925 1810 3955
rect 1840 3925 1970 3955
rect 1800 3905 1970 3925
rect 2000 4025 2170 4045
rect 2000 3995 2010 4025
rect 2040 3995 2170 4025
rect 2000 3955 2170 3995
rect 2000 3925 2010 3955
rect 2040 3925 2170 3955
rect 2000 3905 2170 3925
rect 2200 4025 2370 4045
rect 2200 3995 2210 4025
rect 2240 3995 2370 4025
rect 2200 3955 2370 3995
rect 2200 3925 2210 3955
rect 2240 3925 2370 3955
rect 2200 3905 2370 3925
rect 2400 4025 2570 4045
rect 2400 3995 2410 4025
rect 2440 3995 2570 4025
rect 2400 3955 2570 3995
rect 2400 3925 2410 3955
rect 2440 3925 2570 3955
rect 2400 3905 2570 3925
rect 2600 4025 2770 4045
rect 2600 3995 2610 4025
rect 2640 3995 2770 4025
rect 2600 3955 2770 3995
rect 2600 3925 2610 3955
rect 2640 3925 2770 3955
rect 2600 3905 2770 3925
rect 2800 4025 2970 4045
rect 2800 3995 2810 4025
rect 2840 3995 2970 4025
rect 2800 3955 2970 3995
rect 2800 3925 2810 3955
rect 2840 3925 2970 3955
rect 2800 3905 2970 3925
rect 3000 4025 3170 4045
rect 3000 3995 3010 4025
rect 3040 3995 3170 4025
rect 3000 3955 3170 3995
rect 3000 3925 3010 3955
rect 3040 3925 3170 3955
rect 3000 3905 3170 3925
rect 3200 4025 3370 4045
rect 3200 3995 3210 4025
rect 3240 3995 3370 4025
rect 3200 3955 3370 3995
rect 3200 3925 3210 3955
rect 3240 3925 3370 3955
rect 3200 3905 3370 3925
rect 3400 4025 3570 4045
rect 3400 3995 3410 4025
rect 3440 3995 3570 4025
rect 3400 3955 3570 3995
rect 3400 3925 3410 3955
rect 3440 3925 3570 3955
rect 3400 3905 3570 3925
rect 3600 4025 3770 4045
rect 3600 3995 3610 4025
rect 3640 3995 3770 4025
rect 3600 3955 3770 3995
rect 3600 3925 3610 3955
rect 3640 3925 3770 3955
rect 3600 3905 3770 3925
rect 3800 4025 3970 4045
rect 3800 3995 3810 4025
rect 3840 3995 3970 4025
rect 3800 3955 3970 3995
rect 3800 3925 3810 3955
rect 3840 3925 3970 3955
rect 3800 3905 3970 3925
rect 4000 4025 4170 4045
rect 4000 3995 4010 4025
rect 4040 3995 4170 4025
rect 4000 3955 4170 3995
rect 4000 3925 4010 3955
rect 4040 3925 4170 3955
rect 4000 3905 4170 3925
rect 4200 4025 4370 4045
rect 4200 3995 4210 4025
rect 4240 3995 4370 4025
rect 4200 3955 4370 3995
rect 4200 3925 4210 3955
rect 4240 3925 4370 3955
rect 4200 3905 4370 3925
rect 4400 4025 4570 4045
rect 4400 3995 4410 4025
rect 4440 3995 4570 4025
rect 4400 3955 4570 3995
rect 4400 3925 4410 3955
rect 4440 3925 4570 3955
rect 4400 3905 4570 3925
rect 4600 4025 4770 4045
rect 4600 3995 4610 4025
rect 4640 3995 4770 4025
rect 4600 3955 4770 3995
rect 4600 3925 4610 3955
rect 4640 3925 4770 3955
rect 4600 3905 4770 3925
rect 4800 4025 4970 4045
rect 4800 3995 4810 4025
rect 4840 3995 4970 4025
rect 4800 3955 4970 3995
rect 4800 3925 4810 3955
rect 4840 3925 4970 3955
rect 4800 3905 4970 3925
rect 5000 4025 5170 4045
rect 5000 3995 5010 4025
rect 5040 3995 5170 4025
rect 5000 3955 5170 3995
rect 5000 3925 5010 3955
rect 5040 3925 5170 3955
rect 5000 3905 5170 3925
rect 5200 4025 5370 4045
rect 5200 3995 5210 4025
rect 5240 3995 5370 4025
rect 5200 3955 5370 3995
rect 5200 3925 5210 3955
rect 5240 3925 5370 3955
rect 5200 3905 5370 3925
rect 5400 4025 5570 4045
rect 5400 3995 5410 4025
rect 5440 3995 5570 4025
rect 5400 3955 5570 3995
rect 5400 3925 5410 3955
rect 5440 3925 5570 3955
rect 5400 3905 5570 3925
rect 5600 4025 5770 4045
rect 5600 3995 5610 4025
rect 5640 3995 5770 4025
rect 5600 3955 5770 3995
rect 5600 3925 5610 3955
rect 5640 3925 5770 3955
rect 5600 3905 5770 3925
rect 5800 4025 5970 4045
rect 5800 3995 5810 4025
rect 5840 3995 5970 4025
rect 5800 3955 5970 3995
rect 5800 3925 5810 3955
rect 5840 3925 5970 3955
rect 5800 3905 5970 3925
rect 6000 4025 6170 4045
rect 6000 3995 6010 4025
rect 6040 3995 6170 4025
rect 6000 3955 6170 3995
rect 6000 3925 6010 3955
rect 6040 3925 6170 3955
rect 6000 3905 6170 3925
rect 6200 4025 6370 4045
rect 6200 3995 6210 4025
rect 6240 3995 6370 4025
rect 6200 3955 6370 3995
rect 6200 3925 6210 3955
rect 6240 3925 6370 3955
rect 6200 3905 6370 3925
rect 6400 4025 6570 4045
rect 6400 3995 6410 4025
rect 6440 3995 6570 4025
rect 6400 3955 6570 3995
rect 6400 3925 6410 3955
rect 6440 3925 6570 3955
rect 6400 3905 6570 3925
rect -200 3840 -30 3860
rect -200 3810 -190 3840
rect -160 3810 -30 3840
rect -200 3770 -30 3810
rect -200 3740 -190 3770
rect -160 3740 -30 3770
rect -200 3720 -30 3740
rect 0 3840 170 3860
rect 0 3810 10 3840
rect 40 3810 170 3840
rect 0 3770 170 3810
rect 0 3740 10 3770
rect 40 3740 170 3770
rect 0 3720 170 3740
rect 200 3840 370 3860
rect 200 3810 210 3840
rect 240 3810 370 3840
rect 200 3770 370 3810
rect 200 3740 210 3770
rect 240 3740 370 3770
rect 200 3720 370 3740
rect 400 3840 570 3860
rect 400 3810 410 3840
rect 440 3810 570 3840
rect 400 3770 570 3810
rect 400 3740 410 3770
rect 440 3740 570 3770
rect 400 3720 570 3740
rect 600 3840 770 3860
rect 600 3810 610 3840
rect 640 3810 770 3840
rect 600 3770 770 3810
rect 600 3740 610 3770
rect 640 3740 770 3770
rect 600 3720 770 3740
rect 800 3840 970 3860
rect 800 3810 810 3840
rect 840 3810 970 3840
rect 800 3770 970 3810
rect 800 3740 810 3770
rect 840 3740 970 3770
rect 800 3720 970 3740
rect 1000 3840 1170 3860
rect 1000 3810 1010 3840
rect 1040 3810 1170 3840
rect 1000 3770 1170 3810
rect 1000 3740 1010 3770
rect 1040 3740 1170 3770
rect 1000 3720 1170 3740
rect 1200 3840 1370 3860
rect 1200 3810 1210 3840
rect 1240 3810 1370 3840
rect 1200 3770 1370 3810
rect 1200 3740 1210 3770
rect 1240 3740 1370 3770
rect 1200 3720 1370 3740
rect 1400 3840 1570 3860
rect 1400 3810 1410 3840
rect 1440 3810 1570 3840
rect 1400 3770 1570 3810
rect 1400 3740 1410 3770
rect 1440 3740 1570 3770
rect 1400 3720 1570 3740
rect 1600 3840 1770 3860
rect 1600 3810 1610 3840
rect 1640 3810 1770 3840
rect 1600 3770 1770 3810
rect 1600 3740 1610 3770
rect 1640 3740 1770 3770
rect 1600 3720 1770 3740
rect 1800 3840 1970 3860
rect 1800 3810 1810 3840
rect 1840 3810 1970 3840
rect 1800 3770 1970 3810
rect 1800 3740 1810 3770
rect 1840 3740 1970 3770
rect 1800 3720 1970 3740
rect 2000 3840 2170 3860
rect 2000 3810 2010 3840
rect 2040 3810 2170 3840
rect 2000 3770 2170 3810
rect 2000 3740 2010 3770
rect 2040 3740 2170 3770
rect 2000 3720 2170 3740
rect 2200 3840 2370 3860
rect 2200 3810 2210 3840
rect 2240 3810 2370 3840
rect 2200 3770 2370 3810
rect 2200 3740 2210 3770
rect 2240 3740 2370 3770
rect 2200 3720 2370 3740
rect 2400 3840 2570 3860
rect 2400 3810 2410 3840
rect 2440 3810 2570 3840
rect 2400 3770 2570 3810
rect 2400 3740 2410 3770
rect 2440 3740 2570 3770
rect 2400 3720 2570 3740
rect 2600 3840 2770 3860
rect 2600 3810 2610 3840
rect 2640 3810 2770 3840
rect 2600 3770 2770 3810
rect 2600 3740 2610 3770
rect 2640 3740 2770 3770
rect 2600 3720 2770 3740
rect 2800 3840 2970 3860
rect 2800 3810 2810 3840
rect 2840 3810 2970 3840
rect 2800 3770 2970 3810
rect 2800 3740 2810 3770
rect 2840 3740 2970 3770
rect 2800 3720 2970 3740
rect 3000 3840 3170 3860
rect 3000 3810 3010 3840
rect 3040 3810 3170 3840
rect 3000 3770 3170 3810
rect 3000 3740 3010 3770
rect 3040 3740 3170 3770
rect 3000 3720 3170 3740
rect 3200 3840 3370 3860
rect 3200 3810 3210 3840
rect 3240 3810 3370 3840
rect 3200 3770 3370 3810
rect 3200 3740 3210 3770
rect 3240 3740 3370 3770
rect 3200 3720 3370 3740
rect 3400 3840 3570 3860
rect 3400 3810 3410 3840
rect 3440 3810 3570 3840
rect 3400 3770 3570 3810
rect 3400 3740 3410 3770
rect 3440 3740 3570 3770
rect 3400 3720 3570 3740
rect 3600 3840 3770 3860
rect 3600 3810 3610 3840
rect 3640 3810 3770 3840
rect 3600 3770 3770 3810
rect 3600 3740 3610 3770
rect 3640 3740 3770 3770
rect 3600 3720 3770 3740
rect 3800 3840 3970 3860
rect 3800 3810 3810 3840
rect 3840 3810 3970 3840
rect 3800 3770 3970 3810
rect 3800 3740 3810 3770
rect 3840 3740 3970 3770
rect 3800 3720 3970 3740
rect 4000 3840 4170 3860
rect 4000 3810 4010 3840
rect 4040 3810 4170 3840
rect 4000 3770 4170 3810
rect 4000 3740 4010 3770
rect 4040 3740 4170 3770
rect 4000 3720 4170 3740
rect 4200 3840 4370 3860
rect 4200 3810 4210 3840
rect 4240 3810 4370 3840
rect 4200 3770 4370 3810
rect 4200 3740 4210 3770
rect 4240 3740 4370 3770
rect 4200 3720 4370 3740
rect 4400 3840 4570 3860
rect 4400 3810 4410 3840
rect 4440 3810 4570 3840
rect 4400 3770 4570 3810
rect 4400 3740 4410 3770
rect 4440 3740 4570 3770
rect 4400 3720 4570 3740
rect 4600 3840 4770 3860
rect 4600 3810 4610 3840
rect 4640 3810 4770 3840
rect 4600 3770 4770 3810
rect 4600 3740 4610 3770
rect 4640 3740 4770 3770
rect 4600 3720 4770 3740
rect 4800 3840 4970 3860
rect 4800 3810 4810 3840
rect 4840 3810 4970 3840
rect 4800 3770 4970 3810
rect 4800 3740 4810 3770
rect 4840 3740 4970 3770
rect 4800 3720 4970 3740
rect 5000 3840 5170 3860
rect 5000 3810 5010 3840
rect 5040 3810 5170 3840
rect 5000 3770 5170 3810
rect 5000 3740 5010 3770
rect 5040 3740 5170 3770
rect 5000 3720 5170 3740
rect 5200 3840 5370 3860
rect 5200 3810 5210 3840
rect 5240 3810 5370 3840
rect 5200 3770 5370 3810
rect 5200 3740 5210 3770
rect 5240 3740 5370 3770
rect 5200 3720 5370 3740
rect 5400 3840 5570 3860
rect 5400 3810 5410 3840
rect 5440 3810 5570 3840
rect 5400 3770 5570 3810
rect 5400 3740 5410 3770
rect 5440 3740 5570 3770
rect 5400 3720 5570 3740
rect 5600 3840 5770 3860
rect 5600 3810 5610 3840
rect 5640 3810 5770 3840
rect 5600 3770 5770 3810
rect 5600 3740 5610 3770
rect 5640 3740 5770 3770
rect 5600 3720 5770 3740
rect 5800 3840 5970 3860
rect 5800 3810 5810 3840
rect 5840 3810 5970 3840
rect 5800 3770 5970 3810
rect 5800 3740 5810 3770
rect 5840 3740 5970 3770
rect 5800 3720 5970 3740
rect 6000 3840 6170 3860
rect 6000 3810 6010 3840
rect 6040 3810 6170 3840
rect 6000 3770 6170 3810
rect 6000 3740 6010 3770
rect 6040 3740 6170 3770
rect 6000 3720 6170 3740
rect 6200 3840 6370 3860
rect 6200 3810 6210 3840
rect 6240 3810 6370 3840
rect 6200 3770 6370 3810
rect 6200 3740 6210 3770
rect 6240 3740 6370 3770
rect 6200 3720 6370 3740
rect 6400 3840 6570 3860
rect 6400 3810 6410 3840
rect 6440 3810 6570 3840
rect 6400 3770 6570 3810
rect 6400 3740 6410 3770
rect 6440 3740 6570 3770
rect 6400 3720 6570 3740
rect -200 3655 -30 3675
rect -200 3625 -190 3655
rect -160 3625 -30 3655
rect -200 3585 -30 3625
rect -200 3555 -190 3585
rect -160 3555 -30 3585
rect -200 3535 -30 3555
rect 0 3655 170 3675
rect 0 3625 10 3655
rect 40 3625 170 3655
rect 0 3585 170 3625
rect 0 3555 10 3585
rect 40 3555 170 3585
rect 0 3535 170 3555
rect 200 3655 370 3675
rect 200 3625 210 3655
rect 240 3625 370 3655
rect 200 3585 370 3625
rect 200 3555 210 3585
rect 240 3555 370 3585
rect 200 3535 370 3555
rect 400 3655 570 3675
rect 400 3625 410 3655
rect 440 3625 570 3655
rect 400 3585 570 3625
rect 400 3555 410 3585
rect 440 3555 570 3585
rect 400 3535 570 3555
rect 600 3655 770 3675
rect 600 3625 610 3655
rect 640 3625 770 3655
rect 600 3585 770 3625
rect 600 3555 610 3585
rect 640 3555 770 3585
rect 600 3535 770 3555
rect 800 3655 970 3675
rect 800 3625 810 3655
rect 840 3625 970 3655
rect 800 3585 970 3625
rect 800 3555 810 3585
rect 840 3555 970 3585
rect 800 3535 970 3555
rect 1000 3655 1170 3675
rect 1000 3625 1010 3655
rect 1040 3625 1170 3655
rect 1000 3585 1170 3625
rect 1000 3555 1010 3585
rect 1040 3555 1170 3585
rect 1000 3535 1170 3555
rect 1200 3655 1370 3675
rect 1200 3625 1210 3655
rect 1240 3625 1370 3655
rect 1200 3585 1370 3625
rect 1200 3555 1210 3585
rect 1240 3555 1370 3585
rect 1200 3535 1370 3555
rect 1400 3655 1570 3675
rect 1400 3625 1410 3655
rect 1440 3625 1570 3655
rect 1400 3585 1570 3625
rect 1400 3555 1410 3585
rect 1440 3555 1570 3585
rect 1400 3535 1570 3555
rect 1600 3655 1770 3675
rect 1600 3625 1610 3655
rect 1640 3625 1770 3655
rect 1600 3585 1770 3625
rect 1600 3555 1610 3585
rect 1640 3555 1770 3585
rect 1600 3535 1770 3555
rect 1800 3655 1970 3675
rect 1800 3625 1810 3655
rect 1840 3625 1970 3655
rect 1800 3585 1970 3625
rect 1800 3555 1810 3585
rect 1840 3555 1970 3585
rect 1800 3535 1970 3555
rect 2000 3655 2170 3675
rect 2000 3625 2010 3655
rect 2040 3625 2170 3655
rect 2000 3585 2170 3625
rect 2000 3555 2010 3585
rect 2040 3555 2170 3585
rect 2000 3535 2170 3555
rect 2200 3655 2370 3675
rect 2200 3625 2210 3655
rect 2240 3625 2370 3655
rect 2200 3585 2370 3625
rect 2200 3555 2210 3585
rect 2240 3555 2370 3585
rect 2200 3535 2370 3555
rect 2400 3655 2570 3675
rect 2400 3625 2410 3655
rect 2440 3625 2570 3655
rect 2400 3585 2570 3625
rect 2400 3555 2410 3585
rect 2440 3555 2570 3585
rect 2400 3535 2570 3555
rect 2600 3655 2770 3675
rect 2600 3625 2610 3655
rect 2640 3625 2770 3655
rect 2600 3585 2770 3625
rect 2600 3555 2610 3585
rect 2640 3555 2770 3585
rect 2600 3535 2770 3555
rect 2800 3655 2970 3675
rect 2800 3625 2810 3655
rect 2840 3625 2970 3655
rect 2800 3585 2970 3625
rect 2800 3555 2810 3585
rect 2840 3555 2970 3585
rect 2800 3535 2970 3555
rect 3000 3655 3170 3675
rect 3000 3625 3010 3655
rect 3040 3625 3170 3655
rect 3000 3585 3170 3625
rect 3000 3555 3010 3585
rect 3040 3555 3170 3585
rect 3000 3535 3170 3555
rect 3200 3655 3370 3675
rect 3200 3625 3210 3655
rect 3240 3625 3370 3655
rect 3200 3585 3370 3625
rect 3200 3555 3210 3585
rect 3240 3555 3370 3585
rect 3200 3535 3370 3555
rect 3400 3655 3570 3675
rect 3400 3625 3410 3655
rect 3440 3625 3570 3655
rect 3400 3585 3570 3625
rect 3400 3555 3410 3585
rect 3440 3555 3570 3585
rect 3400 3535 3570 3555
rect 3600 3655 3770 3675
rect 3600 3625 3610 3655
rect 3640 3625 3770 3655
rect 3600 3585 3770 3625
rect 3600 3555 3610 3585
rect 3640 3555 3770 3585
rect 3600 3535 3770 3555
rect 3800 3655 3970 3675
rect 3800 3625 3810 3655
rect 3840 3625 3970 3655
rect 3800 3585 3970 3625
rect 3800 3555 3810 3585
rect 3840 3555 3970 3585
rect 3800 3535 3970 3555
rect 4000 3655 4170 3675
rect 4000 3625 4010 3655
rect 4040 3625 4170 3655
rect 4000 3585 4170 3625
rect 4000 3555 4010 3585
rect 4040 3555 4170 3585
rect 4000 3535 4170 3555
rect 4200 3655 4370 3675
rect 4200 3625 4210 3655
rect 4240 3625 4370 3655
rect 4200 3585 4370 3625
rect 4200 3555 4210 3585
rect 4240 3555 4370 3585
rect 4200 3535 4370 3555
rect 4400 3655 4570 3675
rect 4400 3625 4410 3655
rect 4440 3625 4570 3655
rect 4400 3585 4570 3625
rect 4400 3555 4410 3585
rect 4440 3555 4570 3585
rect 4400 3535 4570 3555
rect 4600 3655 4770 3675
rect 4600 3625 4610 3655
rect 4640 3625 4770 3655
rect 4600 3585 4770 3625
rect 4600 3555 4610 3585
rect 4640 3555 4770 3585
rect 4600 3535 4770 3555
rect 4800 3655 4970 3675
rect 4800 3625 4810 3655
rect 4840 3625 4970 3655
rect 4800 3585 4970 3625
rect 4800 3555 4810 3585
rect 4840 3555 4970 3585
rect 4800 3535 4970 3555
rect 5000 3655 5170 3675
rect 5000 3625 5010 3655
rect 5040 3625 5170 3655
rect 5000 3585 5170 3625
rect 5000 3555 5010 3585
rect 5040 3555 5170 3585
rect 5000 3535 5170 3555
rect 5200 3655 5370 3675
rect 5200 3625 5210 3655
rect 5240 3625 5370 3655
rect 5200 3585 5370 3625
rect 5200 3555 5210 3585
rect 5240 3555 5370 3585
rect 5200 3535 5370 3555
rect 5400 3655 5570 3675
rect 5400 3625 5410 3655
rect 5440 3625 5570 3655
rect 5400 3585 5570 3625
rect 5400 3555 5410 3585
rect 5440 3555 5570 3585
rect 5400 3535 5570 3555
rect 5600 3655 5770 3675
rect 5600 3625 5610 3655
rect 5640 3625 5770 3655
rect 5600 3585 5770 3625
rect 5600 3555 5610 3585
rect 5640 3555 5770 3585
rect 5600 3535 5770 3555
rect 5800 3655 5970 3675
rect 5800 3625 5810 3655
rect 5840 3625 5970 3655
rect 5800 3585 5970 3625
rect 5800 3555 5810 3585
rect 5840 3555 5970 3585
rect 5800 3535 5970 3555
rect 6000 3655 6170 3675
rect 6000 3625 6010 3655
rect 6040 3625 6170 3655
rect 6000 3585 6170 3625
rect 6000 3555 6010 3585
rect 6040 3555 6170 3585
rect 6000 3535 6170 3555
rect 6200 3655 6370 3675
rect 6200 3625 6210 3655
rect 6240 3625 6370 3655
rect 6200 3585 6370 3625
rect 6200 3555 6210 3585
rect 6240 3555 6370 3585
rect 6200 3535 6370 3555
rect 6400 3655 6570 3675
rect 6400 3625 6410 3655
rect 6440 3625 6570 3655
rect 6400 3585 6570 3625
rect 6400 3555 6410 3585
rect 6440 3555 6570 3585
rect 6400 3535 6570 3555
rect -200 3470 -30 3490
rect -200 3440 -190 3470
rect -160 3440 -30 3470
rect -200 3400 -30 3440
rect -200 3370 -190 3400
rect -160 3370 -30 3400
rect -200 3350 -30 3370
rect 0 3470 170 3490
rect 0 3440 10 3470
rect 40 3440 170 3470
rect 0 3400 170 3440
rect 0 3370 10 3400
rect 40 3370 170 3400
rect 0 3350 170 3370
rect 200 3470 370 3490
rect 200 3440 210 3470
rect 240 3440 370 3470
rect 200 3400 370 3440
rect 200 3370 210 3400
rect 240 3370 370 3400
rect 200 3350 370 3370
rect 400 3470 570 3490
rect 400 3440 410 3470
rect 440 3440 570 3470
rect 400 3400 570 3440
rect 400 3370 410 3400
rect 440 3370 570 3400
rect 400 3350 570 3370
rect 600 3470 770 3490
rect 600 3440 610 3470
rect 640 3440 770 3470
rect 600 3400 770 3440
rect 600 3370 610 3400
rect 640 3370 770 3400
rect 600 3350 770 3370
rect 800 3470 970 3490
rect 800 3440 810 3470
rect 840 3440 970 3470
rect 800 3400 970 3440
rect 800 3370 810 3400
rect 840 3370 970 3400
rect 800 3350 970 3370
rect 1000 3470 1170 3490
rect 1000 3440 1010 3470
rect 1040 3440 1170 3470
rect 1000 3400 1170 3440
rect 1000 3370 1010 3400
rect 1040 3370 1170 3400
rect 1000 3350 1170 3370
rect 1200 3470 1370 3490
rect 1200 3440 1210 3470
rect 1240 3440 1370 3470
rect 1200 3400 1370 3440
rect 1200 3370 1210 3400
rect 1240 3370 1370 3400
rect 1200 3350 1370 3370
rect 1400 3470 1570 3490
rect 1400 3440 1410 3470
rect 1440 3440 1570 3470
rect 1400 3400 1570 3440
rect 1400 3370 1410 3400
rect 1440 3370 1570 3400
rect 1400 3350 1570 3370
rect 1600 3470 1770 3490
rect 1600 3440 1610 3470
rect 1640 3440 1770 3470
rect 1600 3400 1770 3440
rect 1600 3370 1610 3400
rect 1640 3370 1770 3400
rect 1600 3350 1770 3370
rect 1800 3470 1970 3490
rect 1800 3440 1810 3470
rect 1840 3440 1970 3470
rect 1800 3400 1970 3440
rect 1800 3370 1810 3400
rect 1840 3370 1970 3400
rect 1800 3350 1970 3370
rect 2000 3470 2170 3490
rect 2000 3440 2010 3470
rect 2040 3440 2170 3470
rect 2000 3400 2170 3440
rect 2000 3370 2010 3400
rect 2040 3370 2170 3400
rect 2000 3350 2170 3370
rect 2200 3470 2370 3490
rect 2200 3440 2210 3470
rect 2240 3440 2370 3470
rect 2200 3400 2370 3440
rect 2200 3370 2210 3400
rect 2240 3370 2370 3400
rect 2200 3350 2370 3370
rect 2400 3470 2570 3490
rect 2400 3440 2410 3470
rect 2440 3440 2570 3470
rect 2400 3400 2570 3440
rect 2400 3370 2410 3400
rect 2440 3370 2570 3400
rect 2400 3350 2570 3370
rect 2600 3470 2770 3490
rect 2600 3440 2610 3470
rect 2640 3440 2770 3470
rect 2600 3400 2770 3440
rect 2600 3370 2610 3400
rect 2640 3370 2770 3400
rect 2600 3350 2770 3370
rect 2800 3470 2970 3490
rect 2800 3440 2810 3470
rect 2840 3440 2970 3470
rect 2800 3400 2970 3440
rect 2800 3370 2810 3400
rect 2840 3370 2970 3400
rect 2800 3350 2970 3370
rect 3000 3470 3170 3490
rect 3000 3440 3010 3470
rect 3040 3440 3170 3470
rect 3000 3400 3170 3440
rect 3000 3370 3010 3400
rect 3040 3370 3170 3400
rect 3000 3350 3170 3370
rect 3200 3470 3370 3490
rect 3200 3440 3210 3470
rect 3240 3440 3370 3470
rect 3200 3400 3370 3440
rect 3200 3370 3210 3400
rect 3240 3370 3370 3400
rect 3200 3350 3370 3370
rect 3400 3470 3570 3490
rect 3400 3440 3410 3470
rect 3440 3440 3570 3470
rect 3400 3400 3570 3440
rect 3400 3370 3410 3400
rect 3440 3370 3570 3400
rect 3400 3350 3570 3370
rect 3600 3470 3770 3490
rect 3600 3440 3610 3470
rect 3640 3440 3770 3470
rect 3600 3400 3770 3440
rect 3600 3370 3610 3400
rect 3640 3370 3770 3400
rect 3600 3350 3770 3370
rect 3800 3470 3970 3490
rect 3800 3440 3810 3470
rect 3840 3440 3970 3470
rect 3800 3400 3970 3440
rect 3800 3370 3810 3400
rect 3840 3370 3970 3400
rect 3800 3350 3970 3370
rect 4000 3470 4170 3490
rect 4000 3440 4010 3470
rect 4040 3440 4170 3470
rect 4000 3400 4170 3440
rect 4000 3370 4010 3400
rect 4040 3370 4170 3400
rect 4000 3350 4170 3370
rect 4200 3470 4370 3490
rect 4200 3440 4210 3470
rect 4240 3440 4370 3470
rect 4200 3400 4370 3440
rect 4200 3370 4210 3400
rect 4240 3370 4370 3400
rect 4200 3350 4370 3370
rect 4400 3470 4570 3490
rect 4400 3440 4410 3470
rect 4440 3440 4570 3470
rect 4400 3400 4570 3440
rect 4400 3370 4410 3400
rect 4440 3370 4570 3400
rect 4400 3350 4570 3370
rect 4600 3470 4770 3490
rect 4600 3440 4610 3470
rect 4640 3440 4770 3470
rect 4600 3400 4770 3440
rect 4600 3370 4610 3400
rect 4640 3370 4770 3400
rect 4600 3350 4770 3370
rect 4800 3470 4970 3490
rect 4800 3440 4810 3470
rect 4840 3440 4970 3470
rect 4800 3400 4970 3440
rect 4800 3370 4810 3400
rect 4840 3370 4970 3400
rect 4800 3350 4970 3370
rect 5000 3470 5170 3490
rect 5000 3440 5010 3470
rect 5040 3440 5170 3470
rect 5000 3400 5170 3440
rect 5000 3370 5010 3400
rect 5040 3370 5170 3400
rect 5000 3350 5170 3370
rect 5200 3470 5370 3490
rect 5200 3440 5210 3470
rect 5240 3440 5370 3470
rect 5200 3400 5370 3440
rect 5200 3370 5210 3400
rect 5240 3370 5370 3400
rect 5200 3350 5370 3370
rect 5400 3470 5570 3490
rect 5400 3440 5410 3470
rect 5440 3440 5570 3470
rect 5400 3400 5570 3440
rect 5400 3370 5410 3400
rect 5440 3370 5570 3400
rect 5400 3350 5570 3370
rect 5600 3470 5770 3490
rect 5600 3440 5610 3470
rect 5640 3440 5770 3470
rect 5600 3400 5770 3440
rect 5600 3370 5610 3400
rect 5640 3370 5770 3400
rect 5600 3350 5770 3370
rect 5800 3470 5970 3490
rect 5800 3440 5810 3470
rect 5840 3440 5970 3470
rect 5800 3400 5970 3440
rect 5800 3370 5810 3400
rect 5840 3370 5970 3400
rect 5800 3350 5970 3370
rect 6000 3470 6170 3490
rect 6000 3440 6010 3470
rect 6040 3440 6170 3470
rect 6000 3400 6170 3440
rect 6000 3370 6010 3400
rect 6040 3370 6170 3400
rect 6000 3350 6170 3370
rect 6200 3470 6370 3490
rect 6200 3440 6210 3470
rect 6240 3440 6370 3470
rect 6200 3400 6370 3440
rect 6200 3370 6210 3400
rect 6240 3370 6370 3400
rect 6200 3350 6370 3370
rect 6400 3470 6570 3490
rect 6400 3440 6410 3470
rect 6440 3440 6570 3470
rect 6400 3400 6570 3440
rect 6400 3370 6410 3400
rect 6440 3370 6570 3400
rect 6400 3350 6570 3370
rect -200 3285 -30 3305
rect -200 3255 -190 3285
rect -160 3255 -30 3285
rect -200 3215 -30 3255
rect -200 3185 -190 3215
rect -160 3185 -30 3215
rect -200 3165 -30 3185
rect 0 3285 170 3305
rect 0 3255 10 3285
rect 40 3255 170 3285
rect 0 3215 170 3255
rect 0 3185 10 3215
rect 40 3185 170 3215
rect 0 3165 170 3185
rect 200 3285 370 3305
rect 200 3255 210 3285
rect 240 3255 370 3285
rect 200 3215 370 3255
rect 200 3185 210 3215
rect 240 3185 370 3215
rect 200 3165 370 3185
rect 400 3285 570 3305
rect 400 3255 410 3285
rect 440 3255 570 3285
rect 400 3215 570 3255
rect 400 3185 410 3215
rect 440 3185 570 3215
rect 400 3165 570 3185
rect 600 3285 770 3305
rect 600 3255 610 3285
rect 640 3255 770 3285
rect 600 3215 770 3255
rect 600 3185 610 3215
rect 640 3185 770 3215
rect 600 3165 770 3185
rect 800 3285 970 3305
rect 800 3255 810 3285
rect 840 3255 970 3285
rect 800 3215 970 3255
rect 800 3185 810 3215
rect 840 3185 970 3215
rect 800 3165 970 3185
rect 1000 3285 1170 3305
rect 1000 3255 1010 3285
rect 1040 3255 1170 3285
rect 1000 3215 1170 3255
rect 1000 3185 1010 3215
rect 1040 3185 1170 3215
rect 1000 3165 1170 3185
rect 1200 3285 1370 3305
rect 1200 3255 1210 3285
rect 1240 3255 1370 3285
rect 1200 3215 1370 3255
rect 1200 3185 1210 3215
rect 1240 3185 1370 3215
rect 1200 3165 1370 3185
rect 1400 3285 1570 3305
rect 1400 3255 1410 3285
rect 1440 3255 1570 3285
rect 1400 3215 1570 3255
rect 1400 3185 1410 3215
rect 1440 3185 1570 3215
rect 1400 3165 1570 3185
rect 1600 3285 1770 3305
rect 1600 3255 1610 3285
rect 1640 3255 1770 3285
rect 1600 3215 1770 3255
rect 1600 3185 1610 3215
rect 1640 3185 1770 3215
rect 1600 3165 1770 3185
rect 1800 3285 1970 3305
rect 1800 3255 1810 3285
rect 1840 3255 1970 3285
rect 1800 3215 1970 3255
rect 1800 3185 1810 3215
rect 1840 3185 1970 3215
rect 1800 3165 1970 3185
rect 2000 3285 2170 3305
rect 2000 3255 2010 3285
rect 2040 3255 2170 3285
rect 2000 3215 2170 3255
rect 2000 3185 2010 3215
rect 2040 3185 2170 3215
rect 2000 3165 2170 3185
rect 2200 3285 2370 3305
rect 2200 3255 2210 3285
rect 2240 3255 2370 3285
rect 2200 3215 2370 3255
rect 2200 3185 2210 3215
rect 2240 3185 2370 3215
rect 2200 3165 2370 3185
rect 2400 3285 2570 3305
rect 2400 3255 2410 3285
rect 2440 3255 2570 3285
rect 2400 3215 2570 3255
rect 2400 3185 2410 3215
rect 2440 3185 2570 3215
rect 2400 3165 2570 3185
rect 2600 3285 2770 3305
rect 2600 3255 2610 3285
rect 2640 3255 2770 3285
rect 2600 3215 2770 3255
rect 2600 3185 2610 3215
rect 2640 3185 2770 3215
rect 2600 3165 2770 3185
rect 2800 3285 2970 3305
rect 2800 3255 2810 3285
rect 2840 3255 2970 3285
rect 2800 3215 2970 3255
rect 2800 3185 2810 3215
rect 2840 3185 2970 3215
rect 2800 3165 2970 3185
rect 3000 3285 3170 3305
rect 3000 3255 3010 3285
rect 3040 3255 3170 3285
rect 3000 3215 3170 3255
rect 3000 3185 3010 3215
rect 3040 3185 3170 3215
rect 3000 3165 3170 3185
rect 3200 3285 3370 3305
rect 3200 3255 3210 3285
rect 3240 3255 3370 3285
rect 3200 3215 3370 3255
rect 3200 3185 3210 3215
rect 3240 3185 3370 3215
rect 3200 3165 3370 3185
rect 3400 3285 3570 3305
rect 3400 3255 3410 3285
rect 3440 3255 3570 3285
rect 3400 3215 3570 3255
rect 3400 3185 3410 3215
rect 3440 3185 3570 3215
rect 3400 3165 3570 3185
rect 3600 3285 3770 3305
rect 3600 3255 3610 3285
rect 3640 3255 3770 3285
rect 3600 3215 3770 3255
rect 3600 3185 3610 3215
rect 3640 3185 3770 3215
rect 3600 3165 3770 3185
rect 3800 3285 3970 3305
rect 3800 3255 3810 3285
rect 3840 3255 3970 3285
rect 3800 3215 3970 3255
rect 3800 3185 3810 3215
rect 3840 3185 3970 3215
rect 3800 3165 3970 3185
rect 4000 3285 4170 3305
rect 4000 3255 4010 3285
rect 4040 3255 4170 3285
rect 4000 3215 4170 3255
rect 4000 3185 4010 3215
rect 4040 3185 4170 3215
rect 4000 3165 4170 3185
rect 4200 3285 4370 3305
rect 4200 3255 4210 3285
rect 4240 3255 4370 3285
rect 4200 3215 4370 3255
rect 4200 3185 4210 3215
rect 4240 3185 4370 3215
rect 4200 3165 4370 3185
rect 4400 3285 4570 3305
rect 4400 3255 4410 3285
rect 4440 3255 4570 3285
rect 4400 3215 4570 3255
rect 4400 3185 4410 3215
rect 4440 3185 4570 3215
rect 4400 3165 4570 3185
rect 4600 3285 4770 3305
rect 4600 3255 4610 3285
rect 4640 3255 4770 3285
rect 4600 3215 4770 3255
rect 4600 3185 4610 3215
rect 4640 3185 4770 3215
rect 4600 3165 4770 3185
rect 4800 3285 4970 3305
rect 4800 3255 4810 3285
rect 4840 3255 4970 3285
rect 4800 3215 4970 3255
rect 4800 3185 4810 3215
rect 4840 3185 4970 3215
rect 4800 3165 4970 3185
rect 5000 3285 5170 3305
rect 5000 3255 5010 3285
rect 5040 3255 5170 3285
rect 5000 3215 5170 3255
rect 5000 3185 5010 3215
rect 5040 3185 5170 3215
rect 5000 3165 5170 3185
rect 5200 3285 5370 3305
rect 5200 3255 5210 3285
rect 5240 3255 5370 3285
rect 5200 3215 5370 3255
rect 5200 3185 5210 3215
rect 5240 3185 5370 3215
rect 5200 3165 5370 3185
rect 5400 3285 5570 3305
rect 5400 3255 5410 3285
rect 5440 3255 5570 3285
rect 5400 3215 5570 3255
rect 5400 3185 5410 3215
rect 5440 3185 5570 3215
rect 5400 3165 5570 3185
rect 5600 3285 5770 3305
rect 5600 3255 5610 3285
rect 5640 3255 5770 3285
rect 5600 3215 5770 3255
rect 5600 3185 5610 3215
rect 5640 3185 5770 3215
rect 5600 3165 5770 3185
rect 5800 3285 5970 3305
rect 5800 3255 5810 3285
rect 5840 3255 5970 3285
rect 5800 3215 5970 3255
rect 5800 3185 5810 3215
rect 5840 3185 5970 3215
rect 5800 3165 5970 3185
rect 6000 3285 6170 3305
rect 6000 3255 6010 3285
rect 6040 3255 6170 3285
rect 6000 3215 6170 3255
rect 6000 3185 6010 3215
rect 6040 3185 6170 3215
rect 6000 3165 6170 3185
rect 6200 3285 6370 3305
rect 6200 3255 6210 3285
rect 6240 3255 6370 3285
rect 6200 3215 6370 3255
rect 6200 3185 6210 3215
rect 6240 3185 6370 3215
rect 6200 3165 6370 3185
rect 6400 3285 6570 3305
rect 6400 3255 6410 3285
rect 6440 3255 6570 3285
rect 6400 3215 6570 3255
rect 6400 3185 6410 3215
rect 6440 3185 6570 3215
rect 6400 3165 6570 3185
rect -200 3100 -30 3120
rect -200 3070 -190 3100
rect -160 3070 -30 3100
rect -200 3030 -30 3070
rect -200 3000 -190 3030
rect -160 3000 -30 3030
rect -200 2980 -30 3000
rect 0 3100 170 3120
rect 0 3070 10 3100
rect 40 3070 170 3100
rect 0 3030 170 3070
rect 0 3000 10 3030
rect 40 3000 170 3030
rect 0 2980 170 3000
rect 200 3100 370 3120
rect 200 3070 210 3100
rect 240 3070 370 3100
rect 200 3030 370 3070
rect 200 3000 210 3030
rect 240 3000 370 3030
rect 200 2980 370 3000
rect 400 3100 570 3120
rect 400 3070 410 3100
rect 440 3070 570 3100
rect 400 3030 570 3070
rect 400 3000 410 3030
rect 440 3000 570 3030
rect 400 2980 570 3000
rect 600 3100 770 3120
rect 600 3070 610 3100
rect 640 3070 770 3100
rect 600 3030 770 3070
rect 600 3000 610 3030
rect 640 3000 770 3030
rect 600 2980 770 3000
rect 800 3100 970 3120
rect 800 3070 810 3100
rect 840 3070 970 3100
rect 800 3030 970 3070
rect 800 3000 810 3030
rect 840 3000 970 3030
rect 800 2980 970 3000
rect 1000 3100 1170 3120
rect 1000 3070 1010 3100
rect 1040 3070 1170 3100
rect 1000 3030 1170 3070
rect 1000 3000 1010 3030
rect 1040 3000 1170 3030
rect 1000 2980 1170 3000
rect 1200 3100 1370 3120
rect 1200 3070 1210 3100
rect 1240 3070 1370 3100
rect 1200 3030 1370 3070
rect 1200 3000 1210 3030
rect 1240 3000 1370 3030
rect 1200 2980 1370 3000
rect 1400 3100 1570 3120
rect 1400 3070 1410 3100
rect 1440 3070 1570 3100
rect 1400 3030 1570 3070
rect 1400 3000 1410 3030
rect 1440 3000 1570 3030
rect 1400 2980 1570 3000
rect 1600 3100 1770 3120
rect 1600 3070 1610 3100
rect 1640 3070 1770 3100
rect 1600 3030 1770 3070
rect 1600 3000 1610 3030
rect 1640 3000 1770 3030
rect 1600 2980 1770 3000
rect 1800 3100 1970 3120
rect 1800 3070 1810 3100
rect 1840 3070 1970 3100
rect 1800 3030 1970 3070
rect 1800 3000 1810 3030
rect 1840 3000 1970 3030
rect 1800 2980 1970 3000
rect 2000 3100 2170 3120
rect 2000 3070 2010 3100
rect 2040 3070 2170 3100
rect 2000 3030 2170 3070
rect 2000 3000 2010 3030
rect 2040 3000 2170 3030
rect 2000 2980 2170 3000
rect 2200 3100 2370 3120
rect 2200 3070 2210 3100
rect 2240 3070 2370 3100
rect 2200 3030 2370 3070
rect 2200 3000 2210 3030
rect 2240 3000 2370 3030
rect 2200 2980 2370 3000
rect 2400 3100 2570 3120
rect 2400 3070 2410 3100
rect 2440 3070 2570 3100
rect 2400 3030 2570 3070
rect 2400 3000 2410 3030
rect 2440 3000 2570 3030
rect 2400 2980 2570 3000
rect 2600 3100 2770 3120
rect 2600 3070 2610 3100
rect 2640 3070 2770 3100
rect 2600 3030 2770 3070
rect 2600 3000 2610 3030
rect 2640 3000 2770 3030
rect 2600 2980 2770 3000
rect 2800 3100 2970 3120
rect 2800 3070 2810 3100
rect 2840 3070 2970 3100
rect 2800 3030 2970 3070
rect 2800 3000 2810 3030
rect 2840 3000 2970 3030
rect 2800 2980 2970 3000
rect 3000 3100 3170 3120
rect 3000 3070 3010 3100
rect 3040 3070 3170 3100
rect 3000 3030 3170 3070
rect 3000 3000 3010 3030
rect 3040 3000 3170 3030
rect 3000 2980 3170 3000
rect 3200 3100 3370 3120
rect 3200 3070 3210 3100
rect 3240 3070 3370 3100
rect 3200 3030 3370 3070
rect 3200 3000 3210 3030
rect 3240 3000 3370 3030
rect 3200 2980 3370 3000
rect 3400 3100 3570 3120
rect 3400 3070 3410 3100
rect 3440 3070 3570 3100
rect 3400 3030 3570 3070
rect 3400 3000 3410 3030
rect 3440 3000 3570 3030
rect 3400 2980 3570 3000
rect 3600 3100 3770 3120
rect 3600 3070 3610 3100
rect 3640 3070 3770 3100
rect 3600 3030 3770 3070
rect 3600 3000 3610 3030
rect 3640 3000 3770 3030
rect 3600 2980 3770 3000
rect 3800 3100 3970 3120
rect 3800 3070 3810 3100
rect 3840 3070 3970 3100
rect 3800 3030 3970 3070
rect 3800 3000 3810 3030
rect 3840 3000 3970 3030
rect 3800 2980 3970 3000
rect 4000 3100 4170 3120
rect 4000 3070 4010 3100
rect 4040 3070 4170 3100
rect 4000 3030 4170 3070
rect 4000 3000 4010 3030
rect 4040 3000 4170 3030
rect 4000 2980 4170 3000
rect 4200 3100 4370 3120
rect 4200 3070 4210 3100
rect 4240 3070 4370 3100
rect 4200 3030 4370 3070
rect 4200 3000 4210 3030
rect 4240 3000 4370 3030
rect 4200 2980 4370 3000
rect 4400 3100 4570 3120
rect 4400 3070 4410 3100
rect 4440 3070 4570 3100
rect 4400 3030 4570 3070
rect 4400 3000 4410 3030
rect 4440 3000 4570 3030
rect 4400 2980 4570 3000
rect 4600 3100 4770 3120
rect 4600 3070 4610 3100
rect 4640 3070 4770 3100
rect 4600 3030 4770 3070
rect 4600 3000 4610 3030
rect 4640 3000 4770 3030
rect 4600 2980 4770 3000
rect 4800 3100 4970 3120
rect 4800 3070 4810 3100
rect 4840 3070 4970 3100
rect 4800 3030 4970 3070
rect 4800 3000 4810 3030
rect 4840 3000 4970 3030
rect 4800 2980 4970 3000
rect 5000 3100 5170 3120
rect 5000 3070 5010 3100
rect 5040 3070 5170 3100
rect 5000 3030 5170 3070
rect 5000 3000 5010 3030
rect 5040 3000 5170 3030
rect 5000 2980 5170 3000
rect 5200 3100 5370 3120
rect 5200 3070 5210 3100
rect 5240 3070 5370 3100
rect 5200 3030 5370 3070
rect 5200 3000 5210 3030
rect 5240 3000 5370 3030
rect 5200 2980 5370 3000
rect 5400 3100 5570 3120
rect 5400 3070 5410 3100
rect 5440 3070 5570 3100
rect 5400 3030 5570 3070
rect 5400 3000 5410 3030
rect 5440 3000 5570 3030
rect 5400 2980 5570 3000
rect 5600 3100 5770 3120
rect 5600 3070 5610 3100
rect 5640 3070 5770 3100
rect 5600 3030 5770 3070
rect 5600 3000 5610 3030
rect 5640 3000 5770 3030
rect 5600 2980 5770 3000
rect 5800 3100 5970 3120
rect 5800 3070 5810 3100
rect 5840 3070 5970 3100
rect 5800 3030 5970 3070
rect 5800 3000 5810 3030
rect 5840 3000 5970 3030
rect 5800 2980 5970 3000
rect 6000 3100 6170 3120
rect 6000 3070 6010 3100
rect 6040 3070 6170 3100
rect 6000 3030 6170 3070
rect 6000 3000 6010 3030
rect 6040 3000 6170 3030
rect 6000 2980 6170 3000
rect 6200 3100 6370 3120
rect 6200 3070 6210 3100
rect 6240 3070 6370 3100
rect 6200 3030 6370 3070
rect 6200 3000 6210 3030
rect 6240 3000 6370 3030
rect 6200 2980 6370 3000
rect 6400 3100 6570 3120
rect 6400 3070 6410 3100
rect 6440 3070 6570 3100
rect 6400 3030 6570 3070
rect 6400 3000 6410 3030
rect 6440 3000 6570 3030
rect 6400 2980 6570 3000
rect -200 2915 -30 2935
rect -200 2885 -190 2915
rect -160 2885 -30 2915
rect -200 2845 -30 2885
rect -200 2815 -190 2845
rect -160 2815 -30 2845
rect -200 2795 -30 2815
rect 0 2915 170 2935
rect 0 2885 10 2915
rect 40 2885 170 2915
rect 0 2845 170 2885
rect 0 2815 10 2845
rect 40 2815 170 2845
rect 0 2795 170 2815
rect 200 2915 370 2935
rect 200 2885 210 2915
rect 240 2885 370 2915
rect 200 2845 370 2885
rect 200 2815 210 2845
rect 240 2815 370 2845
rect 200 2795 370 2815
rect 400 2915 570 2935
rect 400 2885 410 2915
rect 440 2885 570 2915
rect 400 2845 570 2885
rect 400 2815 410 2845
rect 440 2815 570 2845
rect 400 2795 570 2815
rect 600 2915 770 2935
rect 600 2885 610 2915
rect 640 2885 770 2915
rect 600 2845 770 2885
rect 600 2815 610 2845
rect 640 2815 770 2845
rect 600 2795 770 2815
rect 800 2915 970 2935
rect 800 2885 810 2915
rect 840 2885 970 2915
rect 800 2845 970 2885
rect 800 2815 810 2845
rect 840 2815 970 2845
rect 800 2795 970 2815
rect 1000 2915 1170 2935
rect 1000 2885 1010 2915
rect 1040 2885 1170 2915
rect 1000 2845 1170 2885
rect 1000 2815 1010 2845
rect 1040 2815 1170 2845
rect 1000 2795 1170 2815
rect 1200 2915 1370 2935
rect 1200 2885 1210 2915
rect 1240 2885 1370 2915
rect 1200 2845 1370 2885
rect 1200 2815 1210 2845
rect 1240 2815 1370 2845
rect 1200 2795 1370 2815
rect 1400 2915 1570 2935
rect 1400 2885 1410 2915
rect 1440 2885 1570 2915
rect 1400 2845 1570 2885
rect 1400 2815 1410 2845
rect 1440 2815 1570 2845
rect 1400 2795 1570 2815
rect 1600 2915 1770 2935
rect 1600 2885 1610 2915
rect 1640 2885 1770 2915
rect 1600 2845 1770 2885
rect 1600 2815 1610 2845
rect 1640 2815 1770 2845
rect 1600 2795 1770 2815
rect 1800 2915 1970 2935
rect 1800 2885 1810 2915
rect 1840 2885 1970 2915
rect 1800 2845 1970 2885
rect 1800 2815 1810 2845
rect 1840 2815 1970 2845
rect 1800 2795 1970 2815
rect 2000 2915 2170 2935
rect 2000 2885 2010 2915
rect 2040 2885 2170 2915
rect 2000 2845 2170 2885
rect 2000 2815 2010 2845
rect 2040 2815 2170 2845
rect 2000 2795 2170 2815
rect 2200 2915 2370 2935
rect 2200 2885 2210 2915
rect 2240 2885 2370 2915
rect 2200 2845 2370 2885
rect 2200 2815 2210 2845
rect 2240 2815 2370 2845
rect 2200 2795 2370 2815
rect 2400 2915 2570 2935
rect 2400 2885 2410 2915
rect 2440 2885 2570 2915
rect 2400 2845 2570 2885
rect 2400 2815 2410 2845
rect 2440 2815 2570 2845
rect 2400 2795 2570 2815
rect 2600 2915 2770 2935
rect 2600 2885 2610 2915
rect 2640 2885 2770 2915
rect 2600 2845 2770 2885
rect 2600 2815 2610 2845
rect 2640 2815 2770 2845
rect 2600 2795 2770 2815
rect 2800 2915 2970 2935
rect 2800 2885 2810 2915
rect 2840 2885 2970 2915
rect 2800 2845 2970 2885
rect 2800 2815 2810 2845
rect 2840 2815 2970 2845
rect 2800 2795 2970 2815
rect 3000 2915 3170 2935
rect 3000 2885 3010 2915
rect 3040 2885 3170 2915
rect 3000 2845 3170 2885
rect 3000 2815 3010 2845
rect 3040 2815 3170 2845
rect 3000 2795 3170 2815
rect 3200 2915 3370 2935
rect 3200 2885 3210 2915
rect 3240 2885 3370 2915
rect 3200 2845 3370 2885
rect 3200 2815 3210 2845
rect 3240 2815 3370 2845
rect 3200 2795 3370 2815
rect 3400 2915 3570 2935
rect 3400 2885 3410 2915
rect 3440 2885 3570 2915
rect 3400 2845 3570 2885
rect 3400 2815 3410 2845
rect 3440 2815 3570 2845
rect 3400 2795 3570 2815
rect 3600 2915 3770 2935
rect 3600 2885 3610 2915
rect 3640 2885 3770 2915
rect 3600 2845 3770 2885
rect 3600 2815 3610 2845
rect 3640 2815 3770 2845
rect 3600 2795 3770 2815
rect 3800 2915 3970 2935
rect 3800 2885 3810 2915
rect 3840 2885 3970 2915
rect 3800 2845 3970 2885
rect 3800 2815 3810 2845
rect 3840 2815 3970 2845
rect 3800 2795 3970 2815
rect 4000 2915 4170 2935
rect 4000 2885 4010 2915
rect 4040 2885 4170 2915
rect 4000 2845 4170 2885
rect 4000 2815 4010 2845
rect 4040 2815 4170 2845
rect 4000 2795 4170 2815
rect 4200 2915 4370 2935
rect 4200 2885 4210 2915
rect 4240 2885 4370 2915
rect 4200 2845 4370 2885
rect 4200 2815 4210 2845
rect 4240 2815 4370 2845
rect 4200 2795 4370 2815
rect 4400 2915 4570 2935
rect 4400 2885 4410 2915
rect 4440 2885 4570 2915
rect 4400 2845 4570 2885
rect 4400 2815 4410 2845
rect 4440 2815 4570 2845
rect 4400 2795 4570 2815
rect 4600 2915 4770 2935
rect 4600 2885 4610 2915
rect 4640 2885 4770 2915
rect 4600 2845 4770 2885
rect 4600 2815 4610 2845
rect 4640 2815 4770 2845
rect 4600 2795 4770 2815
rect 4800 2915 4970 2935
rect 4800 2885 4810 2915
rect 4840 2885 4970 2915
rect 4800 2845 4970 2885
rect 4800 2815 4810 2845
rect 4840 2815 4970 2845
rect 4800 2795 4970 2815
rect 5000 2915 5170 2935
rect 5000 2885 5010 2915
rect 5040 2885 5170 2915
rect 5000 2845 5170 2885
rect 5000 2815 5010 2845
rect 5040 2815 5170 2845
rect 5000 2795 5170 2815
rect 5200 2915 5370 2935
rect 5200 2885 5210 2915
rect 5240 2885 5370 2915
rect 5200 2845 5370 2885
rect 5200 2815 5210 2845
rect 5240 2815 5370 2845
rect 5200 2795 5370 2815
rect 5400 2915 5570 2935
rect 5400 2885 5410 2915
rect 5440 2885 5570 2915
rect 5400 2845 5570 2885
rect 5400 2815 5410 2845
rect 5440 2815 5570 2845
rect 5400 2795 5570 2815
rect 5600 2915 5770 2935
rect 5600 2885 5610 2915
rect 5640 2885 5770 2915
rect 5600 2845 5770 2885
rect 5600 2815 5610 2845
rect 5640 2815 5770 2845
rect 5600 2795 5770 2815
rect 5800 2915 5970 2935
rect 5800 2885 5810 2915
rect 5840 2885 5970 2915
rect 5800 2845 5970 2885
rect 5800 2815 5810 2845
rect 5840 2815 5970 2845
rect 5800 2795 5970 2815
rect 6000 2915 6170 2935
rect 6000 2885 6010 2915
rect 6040 2885 6170 2915
rect 6000 2845 6170 2885
rect 6000 2815 6010 2845
rect 6040 2815 6170 2845
rect 6000 2795 6170 2815
rect 6200 2915 6370 2935
rect 6200 2885 6210 2915
rect 6240 2885 6370 2915
rect 6200 2845 6370 2885
rect 6200 2815 6210 2845
rect 6240 2815 6370 2845
rect 6200 2795 6370 2815
rect 6400 2915 6570 2935
rect 6400 2885 6410 2915
rect 6440 2885 6570 2915
rect 6400 2845 6570 2885
rect 6400 2815 6410 2845
rect 6440 2815 6570 2845
rect 6400 2795 6570 2815
rect -200 2730 -30 2750
rect -200 2700 -190 2730
rect -160 2700 -30 2730
rect -200 2660 -30 2700
rect -200 2630 -190 2660
rect -160 2630 -30 2660
rect -200 2610 -30 2630
rect 0 2730 170 2750
rect 0 2700 10 2730
rect 40 2700 170 2730
rect 0 2660 170 2700
rect 0 2630 10 2660
rect 40 2630 170 2660
rect 0 2610 170 2630
rect 200 2730 370 2750
rect 200 2700 210 2730
rect 240 2700 370 2730
rect 200 2660 370 2700
rect 200 2630 210 2660
rect 240 2630 370 2660
rect 200 2610 370 2630
rect 400 2730 570 2750
rect 400 2700 410 2730
rect 440 2700 570 2730
rect 400 2660 570 2700
rect 400 2630 410 2660
rect 440 2630 570 2660
rect 400 2610 570 2630
rect 600 2730 770 2750
rect 600 2700 610 2730
rect 640 2700 770 2730
rect 600 2660 770 2700
rect 600 2630 610 2660
rect 640 2630 770 2660
rect 600 2610 770 2630
rect 800 2730 970 2750
rect 800 2700 810 2730
rect 840 2700 970 2730
rect 800 2660 970 2700
rect 800 2630 810 2660
rect 840 2630 970 2660
rect 800 2610 970 2630
rect 1000 2730 1170 2750
rect 1000 2700 1010 2730
rect 1040 2700 1170 2730
rect 1000 2660 1170 2700
rect 1000 2630 1010 2660
rect 1040 2630 1170 2660
rect 1000 2610 1170 2630
rect 1200 2730 1370 2750
rect 1200 2700 1210 2730
rect 1240 2700 1370 2730
rect 1200 2660 1370 2700
rect 1200 2630 1210 2660
rect 1240 2630 1370 2660
rect 1200 2610 1370 2630
rect 1400 2730 1570 2750
rect 1400 2700 1410 2730
rect 1440 2700 1570 2730
rect 1400 2660 1570 2700
rect 1400 2630 1410 2660
rect 1440 2630 1570 2660
rect 1400 2610 1570 2630
rect 1600 2730 1770 2750
rect 1600 2700 1610 2730
rect 1640 2700 1770 2730
rect 1600 2660 1770 2700
rect 1600 2630 1610 2660
rect 1640 2630 1770 2660
rect 1600 2610 1770 2630
rect 1800 2730 1970 2750
rect 1800 2700 1810 2730
rect 1840 2700 1970 2730
rect 1800 2660 1970 2700
rect 1800 2630 1810 2660
rect 1840 2630 1970 2660
rect 1800 2610 1970 2630
rect 2000 2730 2170 2750
rect 2000 2700 2010 2730
rect 2040 2700 2170 2730
rect 2000 2660 2170 2700
rect 2000 2630 2010 2660
rect 2040 2630 2170 2660
rect 2000 2610 2170 2630
rect 2200 2730 2370 2750
rect 2200 2700 2210 2730
rect 2240 2700 2370 2730
rect 2200 2660 2370 2700
rect 2200 2630 2210 2660
rect 2240 2630 2370 2660
rect 2200 2610 2370 2630
rect 2400 2730 2570 2750
rect 2400 2700 2410 2730
rect 2440 2700 2570 2730
rect 2400 2660 2570 2700
rect 2400 2630 2410 2660
rect 2440 2630 2570 2660
rect 2400 2610 2570 2630
rect 2600 2730 2770 2750
rect 2600 2700 2610 2730
rect 2640 2700 2770 2730
rect 2600 2660 2770 2700
rect 2600 2630 2610 2660
rect 2640 2630 2770 2660
rect 2600 2610 2770 2630
rect 2800 2730 2970 2750
rect 2800 2700 2810 2730
rect 2840 2700 2970 2730
rect 2800 2660 2970 2700
rect 2800 2630 2810 2660
rect 2840 2630 2970 2660
rect 2800 2610 2970 2630
rect 3000 2730 3170 2750
rect 3000 2700 3010 2730
rect 3040 2700 3170 2730
rect 3000 2660 3170 2700
rect 3000 2630 3010 2660
rect 3040 2630 3170 2660
rect 3000 2610 3170 2630
rect 3200 2730 3370 2750
rect 3200 2700 3210 2730
rect 3240 2700 3370 2730
rect 3200 2660 3370 2700
rect 3200 2630 3210 2660
rect 3240 2630 3370 2660
rect 3200 2610 3370 2630
rect 3400 2730 3570 2750
rect 3400 2700 3410 2730
rect 3440 2700 3570 2730
rect 3400 2660 3570 2700
rect 3400 2630 3410 2660
rect 3440 2630 3570 2660
rect 3400 2610 3570 2630
rect 3600 2730 3770 2750
rect 3600 2700 3610 2730
rect 3640 2700 3770 2730
rect 3600 2660 3770 2700
rect 3600 2630 3610 2660
rect 3640 2630 3770 2660
rect 3600 2610 3770 2630
rect 3800 2730 3970 2750
rect 3800 2700 3810 2730
rect 3840 2700 3970 2730
rect 3800 2660 3970 2700
rect 3800 2630 3810 2660
rect 3840 2630 3970 2660
rect 3800 2610 3970 2630
rect 4000 2730 4170 2750
rect 4000 2700 4010 2730
rect 4040 2700 4170 2730
rect 4000 2660 4170 2700
rect 4000 2630 4010 2660
rect 4040 2630 4170 2660
rect 4000 2610 4170 2630
rect 4200 2730 4370 2750
rect 4200 2700 4210 2730
rect 4240 2700 4370 2730
rect 4200 2660 4370 2700
rect 4200 2630 4210 2660
rect 4240 2630 4370 2660
rect 4200 2610 4370 2630
rect 4400 2730 4570 2750
rect 4400 2700 4410 2730
rect 4440 2700 4570 2730
rect 4400 2660 4570 2700
rect 4400 2630 4410 2660
rect 4440 2630 4570 2660
rect 4400 2610 4570 2630
rect 4600 2730 4770 2750
rect 4600 2700 4610 2730
rect 4640 2700 4770 2730
rect 4600 2660 4770 2700
rect 4600 2630 4610 2660
rect 4640 2630 4770 2660
rect 4600 2610 4770 2630
rect 4800 2730 4970 2750
rect 4800 2700 4810 2730
rect 4840 2700 4970 2730
rect 4800 2660 4970 2700
rect 4800 2630 4810 2660
rect 4840 2630 4970 2660
rect 4800 2610 4970 2630
rect 5000 2730 5170 2750
rect 5000 2700 5010 2730
rect 5040 2700 5170 2730
rect 5000 2660 5170 2700
rect 5000 2630 5010 2660
rect 5040 2630 5170 2660
rect 5000 2610 5170 2630
rect 5200 2730 5370 2750
rect 5200 2700 5210 2730
rect 5240 2700 5370 2730
rect 5200 2660 5370 2700
rect 5200 2630 5210 2660
rect 5240 2630 5370 2660
rect 5200 2610 5370 2630
rect 5400 2730 5570 2750
rect 5400 2700 5410 2730
rect 5440 2700 5570 2730
rect 5400 2660 5570 2700
rect 5400 2630 5410 2660
rect 5440 2630 5570 2660
rect 5400 2610 5570 2630
rect 5600 2730 5770 2750
rect 5600 2700 5610 2730
rect 5640 2700 5770 2730
rect 5600 2660 5770 2700
rect 5600 2630 5610 2660
rect 5640 2630 5770 2660
rect 5600 2610 5770 2630
rect 5800 2730 5970 2750
rect 5800 2700 5810 2730
rect 5840 2700 5970 2730
rect 5800 2660 5970 2700
rect 5800 2630 5810 2660
rect 5840 2630 5970 2660
rect 5800 2610 5970 2630
rect 6000 2730 6170 2750
rect 6000 2700 6010 2730
rect 6040 2700 6170 2730
rect 6000 2660 6170 2700
rect 6000 2630 6010 2660
rect 6040 2630 6170 2660
rect 6000 2610 6170 2630
rect 6200 2730 6370 2750
rect 6200 2700 6210 2730
rect 6240 2700 6370 2730
rect 6200 2660 6370 2700
rect 6200 2630 6210 2660
rect 6240 2630 6370 2660
rect 6200 2610 6370 2630
rect 6400 2730 6570 2750
rect 6400 2700 6410 2730
rect 6440 2700 6570 2730
rect 6400 2660 6570 2700
rect 6400 2630 6410 2660
rect 6440 2630 6570 2660
rect 6400 2610 6570 2630
rect -200 2545 -30 2565
rect -200 2515 -190 2545
rect -160 2515 -30 2545
rect -200 2475 -30 2515
rect -200 2445 -190 2475
rect -160 2445 -30 2475
rect -200 2425 -30 2445
rect 0 2545 170 2565
rect 0 2515 10 2545
rect 40 2515 170 2545
rect 0 2475 170 2515
rect 0 2445 10 2475
rect 40 2445 170 2475
rect 0 2425 170 2445
rect 200 2545 370 2565
rect 200 2515 210 2545
rect 240 2515 370 2545
rect 200 2475 370 2515
rect 200 2445 210 2475
rect 240 2445 370 2475
rect 200 2425 370 2445
rect 400 2545 570 2565
rect 400 2515 410 2545
rect 440 2515 570 2545
rect 400 2475 570 2515
rect 400 2445 410 2475
rect 440 2445 570 2475
rect 400 2425 570 2445
rect 600 2545 770 2565
rect 600 2515 610 2545
rect 640 2515 770 2545
rect 600 2475 770 2515
rect 600 2445 610 2475
rect 640 2445 770 2475
rect 600 2425 770 2445
rect 800 2545 970 2565
rect 800 2515 810 2545
rect 840 2515 970 2545
rect 800 2475 970 2515
rect 800 2445 810 2475
rect 840 2445 970 2475
rect 800 2425 970 2445
rect 1000 2545 1170 2565
rect 1000 2515 1010 2545
rect 1040 2515 1170 2545
rect 1000 2475 1170 2515
rect 1000 2445 1010 2475
rect 1040 2445 1170 2475
rect 1000 2425 1170 2445
rect 1200 2545 1370 2565
rect 1200 2515 1210 2545
rect 1240 2515 1370 2545
rect 1200 2475 1370 2515
rect 1200 2445 1210 2475
rect 1240 2445 1370 2475
rect 1200 2425 1370 2445
rect 1400 2545 1570 2565
rect 1400 2515 1410 2545
rect 1440 2515 1570 2545
rect 1400 2475 1570 2515
rect 1400 2445 1410 2475
rect 1440 2445 1570 2475
rect 1400 2425 1570 2445
rect 1600 2545 1770 2565
rect 1600 2515 1610 2545
rect 1640 2515 1770 2545
rect 1600 2475 1770 2515
rect 1600 2445 1610 2475
rect 1640 2445 1770 2475
rect 1600 2425 1770 2445
rect 1800 2545 1970 2565
rect 1800 2515 1810 2545
rect 1840 2515 1970 2545
rect 1800 2475 1970 2515
rect 1800 2445 1810 2475
rect 1840 2445 1970 2475
rect 1800 2425 1970 2445
rect 2000 2545 2170 2565
rect 2000 2515 2010 2545
rect 2040 2515 2170 2545
rect 2000 2475 2170 2515
rect 2000 2445 2010 2475
rect 2040 2445 2170 2475
rect 2000 2425 2170 2445
rect 2200 2545 2370 2565
rect 2200 2515 2210 2545
rect 2240 2515 2370 2545
rect 2200 2475 2370 2515
rect 2200 2445 2210 2475
rect 2240 2445 2370 2475
rect 2200 2425 2370 2445
rect 2400 2545 2570 2565
rect 2400 2515 2410 2545
rect 2440 2515 2570 2545
rect 2400 2475 2570 2515
rect 2400 2445 2410 2475
rect 2440 2445 2570 2475
rect 2400 2425 2570 2445
rect 2600 2545 2770 2565
rect 2600 2515 2610 2545
rect 2640 2515 2770 2545
rect 2600 2475 2770 2515
rect 2600 2445 2610 2475
rect 2640 2445 2770 2475
rect 2600 2425 2770 2445
rect 2800 2545 2970 2565
rect 2800 2515 2810 2545
rect 2840 2515 2970 2545
rect 2800 2475 2970 2515
rect 2800 2445 2810 2475
rect 2840 2445 2970 2475
rect 2800 2425 2970 2445
rect 3000 2545 3170 2565
rect 3000 2515 3010 2545
rect 3040 2515 3170 2545
rect 3000 2475 3170 2515
rect 3000 2445 3010 2475
rect 3040 2445 3170 2475
rect 3000 2425 3170 2445
rect 3200 2545 3370 2565
rect 3200 2515 3210 2545
rect 3240 2515 3370 2545
rect 3200 2475 3370 2515
rect 3200 2445 3210 2475
rect 3240 2445 3370 2475
rect 3200 2425 3370 2445
rect 3400 2545 3570 2565
rect 3400 2515 3410 2545
rect 3440 2515 3570 2545
rect 3400 2475 3570 2515
rect 3400 2445 3410 2475
rect 3440 2445 3570 2475
rect 3400 2425 3570 2445
rect 3600 2545 3770 2565
rect 3600 2515 3610 2545
rect 3640 2515 3770 2545
rect 3600 2475 3770 2515
rect 3600 2445 3610 2475
rect 3640 2445 3770 2475
rect 3600 2425 3770 2445
rect 3800 2545 3970 2565
rect 3800 2515 3810 2545
rect 3840 2515 3970 2545
rect 3800 2475 3970 2515
rect 3800 2445 3810 2475
rect 3840 2445 3970 2475
rect 3800 2425 3970 2445
rect 4000 2545 4170 2565
rect 4000 2515 4010 2545
rect 4040 2515 4170 2545
rect 4000 2475 4170 2515
rect 4000 2445 4010 2475
rect 4040 2445 4170 2475
rect 4000 2425 4170 2445
rect 4200 2545 4370 2565
rect 4200 2515 4210 2545
rect 4240 2515 4370 2545
rect 4200 2475 4370 2515
rect 4200 2445 4210 2475
rect 4240 2445 4370 2475
rect 4200 2425 4370 2445
rect 4400 2545 4570 2565
rect 4400 2515 4410 2545
rect 4440 2515 4570 2545
rect 4400 2475 4570 2515
rect 4400 2445 4410 2475
rect 4440 2445 4570 2475
rect 4400 2425 4570 2445
rect 4600 2545 4770 2565
rect 4600 2515 4610 2545
rect 4640 2515 4770 2545
rect 4600 2475 4770 2515
rect 4600 2445 4610 2475
rect 4640 2445 4770 2475
rect 4600 2425 4770 2445
rect 4800 2545 4970 2565
rect 4800 2515 4810 2545
rect 4840 2515 4970 2545
rect 4800 2475 4970 2515
rect 4800 2445 4810 2475
rect 4840 2445 4970 2475
rect 4800 2425 4970 2445
rect 5000 2545 5170 2565
rect 5000 2515 5010 2545
rect 5040 2515 5170 2545
rect 5000 2475 5170 2515
rect 5000 2445 5010 2475
rect 5040 2445 5170 2475
rect 5000 2425 5170 2445
rect 5200 2545 5370 2565
rect 5200 2515 5210 2545
rect 5240 2515 5370 2545
rect 5200 2475 5370 2515
rect 5200 2445 5210 2475
rect 5240 2445 5370 2475
rect 5200 2425 5370 2445
rect 5400 2545 5570 2565
rect 5400 2515 5410 2545
rect 5440 2515 5570 2545
rect 5400 2475 5570 2515
rect 5400 2445 5410 2475
rect 5440 2445 5570 2475
rect 5400 2425 5570 2445
rect 5600 2545 5770 2565
rect 5600 2515 5610 2545
rect 5640 2515 5770 2545
rect 5600 2475 5770 2515
rect 5600 2445 5610 2475
rect 5640 2445 5770 2475
rect 5600 2425 5770 2445
rect 5800 2545 5970 2565
rect 5800 2515 5810 2545
rect 5840 2515 5970 2545
rect 5800 2475 5970 2515
rect 5800 2445 5810 2475
rect 5840 2445 5970 2475
rect 5800 2425 5970 2445
rect 6000 2545 6170 2565
rect 6000 2515 6010 2545
rect 6040 2515 6170 2545
rect 6000 2475 6170 2515
rect 6000 2445 6010 2475
rect 6040 2445 6170 2475
rect 6000 2425 6170 2445
rect 6200 2545 6370 2565
rect 6200 2515 6210 2545
rect 6240 2515 6370 2545
rect 6200 2475 6370 2515
rect 6200 2445 6210 2475
rect 6240 2445 6370 2475
rect 6200 2425 6370 2445
rect 6400 2545 6570 2565
rect 6400 2515 6410 2545
rect 6440 2515 6570 2545
rect 6400 2475 6570 2515
rect 6400 2445 6410 2475
rect 6440 2445 6570 2475
rect 6400 2425 6570 2445
rect -200 2360 -30 2380
rect -200 2330 -190 2360
rect -160 2330 -30 2360
rect -200 2290 -30 2330
rect -200 2260 -190 2290
rect -160 2260 -30 2290
rect -200 2240 -30 2260
rect 0 2360 170 2380
rect 0 2330 10 2360
rect 40 2330 170 2360
rect 0 2290 170 2330
rect 0 2260 10 2290
rect 40 2260 170 2290
rect 0 2240 170 2260
rect 200 2360 370 2380
rect 200 2330 210 2360
rect 240 2330 370 2360
rect 200 2290 370 2330
rect 200 2260 210 2290
rect 240 2260 370 2290
rect 200 2240 370 2260
rect 400 2360 570 2380
rect 400 2330 410 2360
rect 440 2330 570 2360
rect 400 2290 570 2330
rect 400 2260 410 2290
rect 440 2260 570 2290
rect 400 2240 570 2260
rect 600 2360 770 2380
rect 600 2330 610 2360
rect 640 2330 770 2360
rect 600 2290 770 2330
rect 600 2260 610 2290
rect 640 2260 770 2290
rect 600 2240 770 2260
rect 800 2360 970 2380
rect 800 2330 810 2360
rect 840 2330 970 2360
rect 800 2290 970 2330
rect 800 2260 810 2290
rect 840 2260 970 2290
rect 800 2240 970 2260
rect 1000 2360 1170 2380
rect 1000 2330 1010 2360
rect 1040 2330 1170 2360
rect 1000 2290 1170 2330
rect 1000 2260 1010 2290
rect 1040 2260 1170 2290
rect 1000 2240 1170 2260
rect 1200 2360 1370 2380
rect 1200 2330 1210 2360
rect 1240 2330 1370 2360
rect 1200 2290 1370 2330
rect 1200 2260 1210 2290
rect 1240 2260 1370 2290
rect 1200 2240 1370 2260
rect 1400 2360 1570 2380
rect 1400 2330 1410 2360
rect 1440 2330 1570 2360
rect 1400 2290 1570 2330
rect 1400 2260 1410 2290
rect 1440 2260 1570 2290
rect 1400 2240 1570 2260
rect 1600 2360 1770 2380
rect 1600 2330 1610 2360
rect 1640 2330 1770 2360
rect 1600 2290 1770 2330
rect 1600 2260 1610 2290
rect 1640 2260 1770 2290
rect 1600 2240 1770 2260
rect 1800 2360 1970 2380
rect 1800 2330 1810 2360
rect 1840 2330 1970 2360
rect 1800 2290 1970 2330
rect 1800 2260 1810 2290
rect 1840 2260 1970 2290
rect 1800 2240 1970 2260
rect 2000 2360 2170 2380
rect 2000 2330 2010 2360
rect 2040 2330 2170 2360
rect 2000 2290 2170 2330
rect 2000 2260 2010 2290
rect 2040 2260 2170 2290
rect 2000 2240 2170 2260
rect 2200 2360 2370 2380
rect 2200 2330 2210 2360
rect 2240 2330 2370 2360
rect 2200 2290 2370 2330
rect 2200 2260 2210 2290
rect 2240 2260 2370 2290
rect 2200 2240 2370 2260
rect 2400 2360 2570 2380
rect 2400 2330 2410 2360
rect 2440 2330 2570 2360
rect 2400 2290 2570 2330
rect 2400 2260 2410 2290
rect 2440 2260 2570 2290
rect 2400 2240 2570 2260
rect 2600 2360 2770 2380
rect 2600 2330 2610 2360
rect 2640 2330 2770 2360
rect 2600 2290 2770 2330
rect 2600 2260 2610 2290
rect 2640 2260 2770 2290
rect 2600 2240 2770 2260
rect 2800 2360 2970 2380
rect 2800 2330 2810 2360
rect 2840 2330 2970 2360
rect 2800 2290 2970 2330
rect 2800 2260 2810 2290
rect 2840 2260 2970 2290
rect 2800 2240 2970 2260
rect 3000 2360 3170 2380
rect 3000 2330 3010 2360
rect 3040 2330 3170 2360
rect 3000 2290 3170 2330
rect 3000 2260 3010 2290
rect 3040 2260 3170 2290
rect 3000 2240 3170 2260
rect 3200 2360 3370 2380
rect 3200 2330 3210 2360
rect 3240 2330 3370 2360
rect 3200 2290 3370 2330
rect 3200 2260 3210 2290
rect 3240 2260 3370 2290
rect 3200 2240 3370 2260
rect 3400 2360 3570 2380
rect 3400 2330 3410 2360
rect 3440 2330 3570 2360
rect 3400 2290 3570 2330
rect 3400 2260 3410 2290
rect 3440 2260 3570 2290
rect 3400 2240 3570 2260
rect 3600 2360 3770 2380
rect 3600 2330 3610 2360
rect 3640 2330 3770 2360
rect 3600 2290 3770 2330
rect 3600 2260 3610 2290
rect 3640 2260 3770 2290
rect 3600 2240 3770 2260
rect 3800 2360 3970 2380
rect 3800 2330 3810 2360
rect 3840 2330 3970 2360
rect 3800 2290 3970 2330
rect 3800 2260 3810 2290
rect 3840 2260 3970 2290
rect 3800 2240 3970 2260
rect 4000 2360 4170 2380
rect 4000 2330 4010 2360
rect 4040 2330 4170 2360
rect 4000 2290 4170 2330
rect 4000 2260 4010 2290
rect 4040 2260 4170 2290
rect 4000 2240 4170 2260
rect 4200 2360 4370 2380
rect 4200 2330 4210 2360
rect 4240 2330 4370 2360
rect 4200 2290 4370 2330
rect 4200 2260 4210 2290
rect 4240 2260 4370 2290
rect 4200 2240 4370 2260
rect 4400 2360 4570 2380
rect 4400 2330 4410 2360
rect 4440 2330 4570 2360
rect 4400 2290 4570 2330
rect 4400 2260 4410 2290
rect 4440 2260 4570 2290
rect 4400 2240 4570 2260
rect 4600 2360 4770 2380
rect 4600 2330 4610 2360
rect 4640 2330 4770 2360
rect 4600 2290 4770 2330
rect 4600 2260 4610 2290
rect 4640 2260 4770 2290
rect 4600 2240 4770 2260
rect 4800 2360 4970 2380
rect 4800 2330 4810 2360
rect 4840 2330 4970 2360
rect 4800 2290 4970 2330
rect 4800 2260 4810 2290
rect 4840 2260 4970 2290
rect 4800 2240 4970 2260
rect 5000 2360 5170 2380
rect 5000 2330 5010 2360
rect 5040 2330 5170 2360
rect 5000 2290 5170 2330
rect 5000 2260 5010 2290
rect 5040 2260 5170 2290
rect 5000 2240 5170 2260
rect 5200 2360 5370 2380
rect 5200 2330 5210 2360
rect 5240 2330 5370 2360
rect 5200 2290 5370 2330
rect 5200 2260 5210 2290
rect 5240 2260 5370 2290
rect 5200 2240 5370 2260
rect 5400 2360 5570 2380
rect 5400 2330 5410 2360
rect 5440 2330 5570 2360
rect 5400 2290 5570 2330
rect 5400 2260 5410 2290
rect 5440 2260 5570 2290
rect 5400 2240 5570 2260
rect 5600 2360 5770 2380
rect 5600 2330 5610 2360
rect 5640 2330 5770 2360
rect 5600 2290 5770 2330
rect 5600 2260 5610 2290
rect 5640 2260 5770 2290
rect 5600 2240 5770 2260
rect 5800 2360 5970 2380
rect 5800 2330 5810 2360
rect 5840 2330 5970 2360
rect 5800 2290 5970 2330
rect 5800 2260 5810 2290
rect 5840 2260 5970 2290
rect 5800 2240 5970 2260
rect 6000 2360 6170 2380
rect 6000 2330 6010 2360
rect 6040 2330 6170 2360
rect 6000 2290 6170 2330
rect 6000 2260 6010 2290
rect 6040 2260 6170 2290
rect 6000 2240 6170 2260
rect 6200 2360 6370 2380
rect 6200 2330 6210 2360
rect 6240 2330 6370 2360
rect 6200 2290 6370 2330
rect 6200 2260 6210 2290
rect 6240 2260 6370 2290
rect 6200 2240 6370 2260
rect 6400 2360 6570 2380
rect 6400 2330 6410 2360
rect 6440 2330 6570 2360
rect 6400 2290 6570 2330
rect 6400 2260 6410 2290
rect 6440 2260 6570 2290
rect 6400 2240 6570 2260
rect -200 2175 -30 2195
rect -200 2145 -190 2175
rect -160 2145 -30 2175
rect -200 2105 -30 2145
rect -200 2075 -190 2105
rect -160 2075 -30 2105
rect -200 2055 -30 2075
rect 0 2175 170 2195
rect 0 2145 10 2175
rect 40 2145 170 2175
rect 0 2105 170 2145
rect 0 2075 10 2105
rect 40 2075 170 2105
rect 0 2055 170 2075
rect 200 2175 370 2195
rect 200 2145 210 2175
rect 240 2145 370 2175
rect 200 2105 370 2145
rect 200 2075 210 2105
rect 240 2075 370 2105
rect 200 2055 370 2075
rect 400 2175 570 2195
rect 400 2145 410 2175
rect 440 2145 570 2175
rect 400 2105 570 2145
rect 400 2075 410 2105
rect 440 2075 570 2105
rect 400 2055 570 2075
rect 600 2175 770 2195
rect 600 2145 610 2175
rect 640 2145 770 2175
rect 600 2105 770 2145
rect 600 2075 610 2105
rect 640 2075 770 2105
rect 600 2055 770 2075
rect 800 2175 970 2195
rect 800 2145 810 2175
rect 840 2145 970 2175
rect 800 2105 970 2145
rect 800 2075 810 2105
rect 840 2075 970 2105
rect 800 2055 970 2075
rect 1000 2175 1170 2195
rect 1000 2145 1010 2175
rect 1040 2145 1170 2175
rect 1000 2105 1170 2145
rect 1000 2075 1010 2105
rect 1040 2075 1170 2105
rect 1000 2055 1170 2075
rect 1200 2175 1370 2195
rect 1200 2145 1210 2175
rect 1240 2145 1370 2175
rect 1200 2105 1370 2145
rect 1200 2075 1210 2105
rect 1240 2075 1370 2105
rect 1200 2055 1370 2075
rect 1400 2175 1570 2195
rect 1400 2145 1410 2175
rect 1440 2145 1570 2175
rect 1400 2105 1570 2145
rect 1400 2075 1410 2105
rect 1440 2075 1570 2105
rect 1400 2055 1570 2075
rect 1600 2175 1770 2195
rect 1600 2145 1610 2175
rect 1640 2145 1770 2175
rect 1600 2105 1770 2145
rect 1600 2075 1610 2105
rect 1640 2075 1770 2105
rect 1600 2055 1770 2075
rect 1800 2175 1970 2195
rect 1800 2145 1810 2175
rect 1840 2145 1970 2175
rect 1800 2105 1970 2145
rect 1800 2075 1810 2105
rect 1840 2075 1970 2105
rect 1800 2055 1970 2075
rect 2000 2175 2170 2195
rect 2000 2145 2010 2175
rect 2040 2145 2170 2175
rect 2000 2105 2170 2145
rect 2000 2075 2010 2105
rect 2040 2075 2170 2105
rect 2000 2055 2170 2075
rect 2200 2175 2370 2195
rect 2200 2145 2210 2175
rect 2240 2145 2370 2175
rect 2200 2105 2370 2145
rect 2200 2075 2210 2105
rect 2240 2075 2370 2105
rect 2200 2055 2370 2075
rect 2400 2175 2570 2195
rect 2400 2145 2410 2175
rect 2440 2145 2570 2175
rect 2400 2105 2570 2145
rect 2400 2075 2410 2105
rect 2440 2075 2570 2105
rect 2400 2055 2570 2075
rect 2600 2175 2770 2195
rect 2600 2145 2610 2175
rect 2640 2145 2770 2175
rect 2600 2105 2770 2145
rect 2600 2075 2610 2105
rect 2640 2075 2770 2105
rect 2600 2055 2770 2075
rect 2800 2175 2970 2195
rect 2800 2145 2810 2175
rect 2840 2145 2970 2175
rect 2800 2105 2970 2145
rect 2800 2075 2810 2105
rect 2840 2075 2970 2105
rect 2800 2055 2970 2075
rect 3000 2175 3170 2195
rect 3000 2145 3010 2175
rect 3040 2145 3170 2175
rect 3000 2105 3170 2145
rect 3000 2075 3010 2105
rect 3040 2075 3170 2105
rect 3000 2055 3170 2075
rect 3200 2175 3370 2195
rect 3200 2145 3210 2175
rect 3240 2145 3370 2175
rect 3200 2105 3370 2145
rect 3200 2075 3210 2105
rect 3240 2075 3370 2105
rect 3200 2055 3370 2075
rect 3400 2175 3570 2195
rect 3400 2145 3410 2175
rect 3440 2145 3570 2175
rect 3400 2105 3570 2145
rect 3400 2075 3410 2105
rect 3440 2075 3570 2105
rect 3400 2055 3570 2075
rect 3600 2175 3770 2195
rect 3600 2145 3610 2175
rect 3640 2145 3770 2175
rect 3600 2105 3770 2145
rect 3600 2075 3610 2105
rect 3640 2075 3770 2105
rect 3600 2055 3770 2075
rect 3800 2175 3970 2195
rect 3800 2145 3810 2175
rect 3840 2145 3970 2175
rect 3800 2105 3970 2145
rect 3800 2075 3810 2105
rect 3840 2075 3970 2105
rect 3800 2055 3970 2075
rect 4000 2175 4170 2195
rect 4000 2145 4010 2175
rect 4040 2145 4170 2175
rect 4000 2105 4170 2145
rect 4000 2075 4010 2105
rect 4040 2075 4170 2105
rect 4000 2055 4170 2075
rect 4200 2175 4370 2195
rect 4200 2145 4210 2175
rect 4240 2145 4370 2175
rect 4200 2105 4370 2145
rect 4200 2075 4210 2105
rect 4240 2075 4370 2105
rect 4200 2055 4370 2075
rect 4400 2175 4570 2195
rect 4400 2145 4410 2175
rect 4440 2145 4570 2175
rect 4400 2105 4570 2145
rect 4400 2075 4410 2105
rect 4440 2075 4570 2105
rect 4400 2055 4570 2075
rect 4600 2175 4770 2195
rect 4600 2145 4610 2175
rect 4640 2145 4770 2175
rect 4600 2105 4770 2145
rect 4600 2075 4610 2105
rect 4640 2075 4770 2105
rect 4600 2055 4770 2075
rect 4800 2175 4970 2195
rect 4800 2145 4810 2175
rect 4840 2145 4970 2175
rect 4800 2105 4970 2145
rect 4800 2075 4810 2105
rect 4840 2075 4970 2105
rect 4800 2055 4970 2075
rect 5000 2175 5170 2195
rect 5000 2145 5010 2175
rect 5040 2145 5170 2175
rect 5000 2105 5170 2145
rect 5000 2075 5010 2105
rect 5040 2075 5170 2105
rect 5000 2055 5170 2075
rect 5200 2175 5370 2195
rect 5200 2145 5210 2175
rect 5240 2145 5370 2175
rect 5200 2105 5370 2145
rect 5200 2075 5210 2105
rect 5240 2075 5370 2105
rect 5200 2055 5370 2075
rect 5400 2175 5570 2195
rect 5400 2145 5410 2175
rect 5440 2145 5570 2175
rect 5400 2105 5570 2145
rect 5400 2075 5410 2105
rect 5440 2075 5570 2105
rect 5400 2055 5570 2075
rect 5600 2175 5770 2195
rect 5600 2145 5610 2175
rect 5640 2145 5770 2175
rect 5600 2105 5770 2145
rect 5600 2075 5610 2105
rect 5640 2075 5770 2105
rect 5600 2055 5770 2075
rect 5800 2175 5970 2195
rect 5800 2145 5810 2175
rect 5840 2145 5970 2175
rect 5800 2105 5970 2145
rect 5800 2075 5810 2105
rect 5840 2075 5970 2105
rect 5800 2055 5970 2075
rect 6000 2175 6170 2195
rect 6000 2145 6010 2175
rect 6040 2145 6170 2175
rect 6000 2105 6170 2145
rect 6000 2075 6010 2105
rect 6040 2075 6170 2105
rect 6000 2055 6170 2075
rect 6200 2175 6370 2195
rect 6200 2145 6210 2175
rect 6240 2145 6370 2175
rect 6200 2105 6370 2145
rect 6200 2075 6210 2105
rect 6240 2075 6370 2105
rect 6200 2055 6370 2075
rect 6400 2175 6570 2195
rect 6400 2145 6410 2175
rect 6440 2145 6570 2175
rect 6400 2105 6570 2145
rect 6400 2075 6410 2105
rect 6440 2075 6570 2105
rect 6400 2055 6570 2075
rect -200 1990 -30 2010
rect -200 1960 -190 1990
rect -160 1960 -30 1990
rect -200 1920 -30 1960
rect -200 1890 -190 1920
rect -160 1890 -30 1920
rect -200 1870 -30 1890
rect 0 1990 170 2010
rect 0 1960 10 1990
rect 40 1960 170 1990
rect 0 1920 170 1960
rect 0 1890 10 1920
rect 40 1890 170 1920
rect 0 1870 170 1890
rect 200 1990 370 2010
rect 200 1960 210 1990
rect 240 1960 370 1990
rect 200 1920 370 1960
rect 200 1890 210 1920
rect 240 1890 370 1920
rect 200 1870 370 1890
rect 400 1990 570 2010
rect 400 1960 410 1990
rect 440 1960 570 1990
rect 400 1920 570 1960
rect 400 1890 410 1920
rect 440 1890 570 1920
rect 400 1870 570 1890
rect 600 1990 770 2010
rect 600 1960 610 1990
rect 640 1960 770 1990
rect 600 1920 770 1960
rect 600 1890 610 1920
rect 640 1890 770 1920
rect 600 1870 770 1890
rect 800 1990 970 2010
rect 800 1960 810 1990
rect 840 1960 970 1990
rect 800 1920 970 1960
rect 800 1890 810 1920
rect 840 1890 970 1920
rect 800 1870 970 1890
rect 1000 1990 1170 2010
rect 1000 1960 1010 1990
rect 1040 1960 1170 1990
rect 1000 1920 1170 1960
rect 1000 1890 1010 1920
rect 1040 1890 1170 1920
rect 1000 1870 1170 1890
rect 1200 1990 1370 2010
rect 1200 1960 1210 1990
rect 1240 1960 1370 1990
rect 1200 1920 1370 1960
rect 1200 1890 1210 1920
rect 1240 1890 1370 1920
rect 1200 1870 1370 1890
rect 1400 1990 1570 2010
rect 1400 1960 1410 1990
rect 1440 1960 1570 1990
rect 1400 1920 1570 1960
rect 1400 1890 1410 1920
rect 1440 1890 1570 1920
rect 1400 1870 1570 1890
rect 1600 1990 1770 2010
rect 1600 1960 1610 1990
rect 1640 1960 1770 1990
rect 1600 1920 1770 1960
rect 1600 1890 1610 1920
rect 1640 1890 1770 1920
rect 1600 1870 1770 1890
rect 1800 1990 1970 2010
rect 1800 1960 1810 1990
rect 1840 1960 1970 1990
rect 1800 1920 1970 1960
rect 1800 1890 1810 1920
rect 1840 1890 1970 1920
rect 1800 1870 1970 1890
rect 2000 1990 2170 2010
rect 2000 1960 2010 1990
rect 2040 1960 2170 1990
rect 2000 1920 2170 1960
rect 2000 1890 2010 1920
rect 2040 1890 2170 1920
rect 2000 1870 2170 1890
rect 2200 1990 2370 2010
rect 2200 1960 2210 1990
rect 2240 1960 2370 1990
rect 2200 1920 2370 1960
rect 2200 1890 2210 1920
rect 2240 1890 2370 1920
rect 2200 1870 2370 1890
rect 2400 1990 2570 2010
rect 2400 1960 2410 1990
rect 2440 1960 2570 1990
rect 2400 1920 2570 1960
rect 2400 1890 2410 1920
rect 2440 1890 2570 1920
rect 2400 1870 2570 1890
rect 2600 1990 2770 2010
rect 2600 1960 2610 1990
rect 2640 1960 2770 1990
rect 2600 1920 2770 1960
rect 2600 1890 2610 1920
rect 2640 1890 2770 1920
rect 2600 1870 2770 1890
rect 2800 1990 2970 2010
rect 2800 1960 2810 1990
rect 2840 1960 2970 1990
rect 2800 1920 2970 1960
rect 2800 1890 2810 1920
rect 2840 1890 2970 1920
rect 2800 1870 2970 1890
rect 3000 1990 3170 2010
rect 3000 1960 3010 1990
rect 3040 1960 3170 1990
rect 3000 1920 3170 1960
rect 3000 1890 3010 1920
rect 3040 1890 3170 1920
rect 3000 1870 3170 1890
rect 3200 1990 3370 2010
rect 3200 1960 3210 1990
rect 3240 1960 3370 1990
rect 3200 1920 3370 1960
rect 3200 1890 3210 1920
rect 3240 1890 3370 1920
rect 3200 1870 3370 1890
rect 3400 1990 3570 2010
rect 3400 1960 3410 1990
rect 3440 1960 3570 1990
rect 3400 1920 3570 1960
rect 3400 1890 3410 1920
rect 3440 1890 3570 1920
rect 3400 1870 3570 1890
rect 3600 1990 3770 2010
rect 3600 1960 3610 1990
rect 3640 1960 3770 1990
rect 3600 1920 3770 1960
rect 3600 1890 3610 1920
rect 3640 1890 3770 1920
rect 3600 1870 3770 1890
rect 3800 1990 3970 2010
rect 3800 1960 3810 1990
rect 3840 1960 3970 1990
rect 3800 1920 3970 1960
rect 3800 1890 3810 1920
rect 3840 1890 3970 1920
rect 3800 1870 3970 1890
rect 4000 1990 4170 2010
rect 4000 1960 4010 1990
rect 4040 1960 4170 1990
rect 4000 1920 4170 1960
rect 4000 1890 4010 1920
rect 4040 1890 4170 1920
rect 4000 1870 4170 1890
rect 4200 1990 4370 2010
rect 4200 1960 4210 1990
rect 4240 1960 4370 1990
rect 4200 1920 4370 1960
rect 4200 1890 4210 1920
rect 4240 1890 4370 1920
rect 4200 1870 4370 1890
rect 4400 1990 4570 2010
rect 4400 1960 4410 1990
rect 4440 1960 4570 1990
rect 4400 1920 4570 1960
rect 4400 1890 4410 1920
rect 4440 1890 4570 1920
rect 4400 1870 4570 1890
rect 4600 1990 4770 2010
rect 4600 1960 4610 1990
rect 4640 1960 4770 1990
rect 4600 1920 4770 1960
rect 4600 1890 4610 1920
rect 4640 1890 4770 1920
rect 4600 1870 4770 1890
rect 4800 1990 4970 2010
rect 4800 1960 4810 1990
rect 4840 1960 4970 1990
rect 4800 1920 4970 1960
rect 4800 1890 4810 1920
rect 4840 1890 4970 1920
rect 4800 1870 4970 1890
rect 5000 1990 5170 2010
rect 5000 1960 5010 1990
rect 5040 1960 5170 1990
rect 5000 1920 5170 1960
rect 5000 1890 5010 1920
rect 5040 1890 5170 1920
rect 5000 1870 5170 1890
rect 5200 1990 5370 2010
rect 5200 1960 5210 1990
rect 5240 1960 5370 1990
rect 5200 1920 5370 1960
rect 5200 1890 5210 1920
rect 5240 1890 5370 1920
rect 5200 1870 5370 1890
rect 5400 1990 5570 2010
rect 5400 1960 5410 1990
rect 5440 1960 5570 1990
rect 5400 1920 5570 1960
rect 5400 1890 5410 1920
rect 5440 1890 5570 1920
rect 5400 1870 5570 1890
rect 5600 1990 5770 2010
rect 5600 1960 5610 1990
rect 5640 1960 5770 1990
rect 5600 1920 5770 1960
rect 5600 1890 5610 1920
rect 5640 1890 5770 1920
rect 5600 1870 5770 1890
rect 5800 1990 5970 2010
rect 5800 1960 5810 1990
rect 5840 1960 5970 1990
rect 5800 1920 5970 1960
rect 5800 1890 5810 1920
rect 5840 1890 5970 1920
rect 5800 1870 5970 1890
rect 6000 1990 6170 2010
rect 6000 1960 6010 1990
rect 6040 1960 6170 1990
rect 6000 1920 6170 1960
rect 6000 1890 6010 1920
rect 6040 1890 6170 1920
rect 6000 1870 6170 1890
rect 6200 1990 6370 2010
rect 6200 1960 6210 1990
rect 6240 1960 6370 1990
rect 6200 1920 6370 1960
rect 6200 1890 6210 1920
rect 6240 1890 6370 1920
rect 6200 1870 6370 1890
rect 6400 1990 6570 2010
rect 6400 1960 6410 1990
rect 6440 1960 6570 1990
rect 6400 1920 6570 1960
rect 6400 1890 6410 1920
rect 6440 1890 6570 1920
rect 6400 1870 6570 1890
rect -200 1805 -30 1825
rect -200 1775 -190 1805
rect -160 1775 -30 1805
rect -200 1735 -30 1775
rect -200 1705 -190 1735
rect -160 1705 -30 1735
rect -200 1685 -30 1705
rect 0 1805 170 1825
rect 0 1775 10 1805
rect 40 1775 170 1805
rect 0 1735 170 1775
rect 0 1705 10 1735
rect 40 1705 170 1735
rect 0 1685 170 1705
rect 200 1805 370 1825
rect 200 1775 210 1805
rect 240 1775 370 1805
rect 200 1735 370 1775
rect 200 1705 210 1735
rect 240 1705 370 1735
rect 200 1685 370 1705
rect 400 1805 570 1825
rect 400 1775 410 1805
rect 440 1775 570 1805
rect 400 1735 570 1775
rect 400 1705 410 1735
rect 440 1705 570 1735
rect 400 1685 570 1705
rect 600 1805 770 1825
rect 600 1775 610 1805
rect 640 1775 770 1805
rect 600 1735 770 1775
rect 600 1705 610 1735
rect 640 1705 770 1735
rect 600 1685 770 1705
rect 800 1805 970 1825
rect 800 1775 810 1805
rect 840 1775 970 1805
rect 800 1735 970 1775
rect 800 1705 810 1735
rect 840 1705 970 1735
rect 800 1685 970 1705
rect 1000 1805 1170 1825
rect 1000 1775 1010 1805
rect 1040 1775 1170 1805
rect 1000 1735 1170 1775
rect 1000 1705 1010 1735
rect 1040 1705 1170 1735
rect 1000 1685 1170 1705
rect 1200 1805 1370 1825
rect 1200 1775 1210 1805
rect 1240 1775 1370 1805
rect 1200 1735 1370 1775
rect 1200 1705 1210 1735
rect 1240 1705 1370 1735
rect 1200 1685 1370 1705
rect 1400 1805 1570 1825
rect 1400 1775 1410 1805
rect 1440 1775 1570 1805
rect 1400 1735 1570 1775
rect 1400 1705 1410 1735
rect 1440 1705 1570 1735
rect 1400 1685 1570 1705
rect 1600 1805 1770 1825
rect 1600 1775 1610 1805
rect 1640 1775 1770 1805
rect 1600 1735 1770 1775
rect 1600 1705 1610 1735
rect 1640 1705 1770 1735
rect 1600 1685 1770 1705
rect 1800 1805 1970 1825
rect 1800 1775 1810 1805
rect 1840 1775 1970 1805
rect 1800 1735 1970 1775
rect 1800 1705 1810 1735
rect 1840 1705 1970 1735
rect 1800 1685 1970 1705
rect 2000 1805 2170 1825
rect 2000 1775 2010 1805
rect 2040 1775 2170 1805
rect 2000 1735 2170 1775
rect 2000 1705 2010 1735
rect 2040 1705 2170 1735
rect 2000 1685 2170 1705
rect 2200 1805 2370 1825
rect 2200 1775 2210 1805
rect 2240 1775 2370 1805
rect 2200 1735 2370 1775
rect 2200 1705 2210 1735
rect 2240 1705 2370 1735
rect 2200 1685 2370 1705
rect 2400 1805 2570 1825
rect 2400 1775 2410 1805
rect 2440 1775 2570 1805
rect 2400 1735 2570 1775
rect 2400 1705 2410 1735
rect 2440 1705 2570 1735
rect 2400 1685 2570 1705
rect 2600 1805 2770 1825
rect 2600 1775 2610 1805
rect 2640 1775 2770 1805
rect 2600 1735 2770 1775
rect 2600 1705 2610 1735
rect 2640 1705 2770 1735
rect 2600 1685 2770 1705
rect 2800 1805 2970 1825
rect 2800 1775 2810 1805
rect 2840 1775 2970 1805
rect 2800 1735 2970 1775
rect 2800 1705 2810 1735
rect 2840 1705 2970 1735
rect 2800 1685 2970 1705
rect 3000 1805 3170 1825
rect 3000 1775 3010 1805
rect 3040 1775 3170 1805
rect 3000 1735 3170 1775
rect 3000 1705 3010 1735
rect 3040 1705 3170 1735
rect 3000 1685 3170 1705
rect 3200 1805 3370 1825
rect 3200 1775 3210 1805
rect 3240 1775 3370 1805
rect 3200 1735 3370 1775
rect 3200 1705 3210 1735
rect 3240 1705 3370 1735
rect 3200 1685 3370 1705
rect 3400 1805 3570 1825
rect 3400 1775 3410 1805
rect 3440 1775 3570 1805
rect 3400 1735 3570 1775
rect 3400 1705 3410 1735
rect 3440 1705 3570 1735
rect 3400 1685 3570 1705
rect 3600 1805 3770 1825
rect 3600 1775 3610 1805
rect 3640 1775 3770 1805
rect 3600 1735 3770 1775
rect 3600 1705 3610 1735
rect 3640 1705 3770 1735
rect 3600 1685 3770 1705
rect 3800 1805 3970 1825
rect 3800 1775 3810 1805
rect 3840 1775 3970 1805
rect 3800 1735 3970 1775
rect 3800 1705 3810 1735
rect 3840 1705 3970 1735
rect 3800 1685 3970 1705
rect 4000 1805 4170 1825
rect 4000 1775 4010 1805
rect 4040 1775 4170 1805
rect 4000 1735 4170 1775
rect 4000 1705 4010 1735
rect 4040 1705 4170 1735
rect 4000 1685 4170 1705
rect 4200 1805 4370 1825
rect 4200 1775 4210 1805
rect 4240 1775 4370 1805
rect 4200 1735 4370 1775
rect 4200 1705 4210 1735
rect 4240 1705 4370 1735
rect 4200 1685 4370 1705
rect 4400 1805 4570 1825
rect 4400 1775 4410 1805
rect 4440 1775 4570 1805
rect 4400 1735 4570 1775
rect 4400 1705 4410 1735
rect 4440 1705 4570 1735
rect 4400 1685 4570 1705
rect 4600 1805 4770 1825
rect 4600 1775 4610 1805
rect 4640 1775 4770 1805
rect 4600 1735 4770 1775
rect 4600 1705 4610 1735
rect 4640 1705 4770 1735
rect 4600 1685 4770 1705
rect 4800 1805 4970 1825
rect 4800 1775 4810 1805
rect 4840 1775 4970 1805
rect 4800 1735 4970 1775
rect 4800 1705 4810 1735
rect 4840 1705 4970 1735
rect 4800 1685 4970 1705
rect 5000 1805 5170 1825
rect 5000 1775 5010 1805
rect 5040 1775 5170 1805
rect 5000 1735 5170 1775
rect 5000 1705 5010 1735
rect 5040 1705 5170 1735
rect 5000 1685 5170 1705
rect 5200 1805 5370 1825
rect 5200 1775 5210 1805
rect 5240 1775 5370 1805
rect 5200 1735 5370 1775
rect 5200 1705 5210 1735
rect 5240 1705 5370 1735
rect 5200 1685 5370 1705
rect 5400 1805 5570 1825
rect 5400 1775 5410 1805
rect 5440 1775 5570 1805
rect 5400 1735 5570 1775
rect 5400 1705 5410 1735
rect 5440 1705 5570 1735
rect 5400 1685 5570 1705
rect 5600 1805 5770 1825
rect 5600 1775 5610 1805
rect 5640 1775 5770 1805
rect 5600 1735 5770 1775
rect 5600 1705 5610 1735
rect 5640 1705 5770 1735
rect 5600 1685 5770 1705
rect 5800 1805 5970 1825
rect 5800 1775 5810 1805
rect 5840 1775 5970 1805
rect 5800 1735 5970 1775
rect 5800 1705 5810 1735
rect 5840 1705 5970 1735
rect 5800 1685 5970 1705
rect 6000 1805 6170 1825
rect 6000 1775 6010 1805
rect 6040 1775 6170 1805
rect 6000 1735 6170 1775
rect 6000 1705 6010 1735
rect 6040 1705 6170 1735
rect 6000 1685 6170 1705
rect 6200 1805 6370 1825
rect 6200 1775 6210 1805
rect 6240 1775 6370 1805
rect 6200 1735 6370 1775
rect 6200 1705 6210 1735
rect 6240 1705 6370 1735
rect 6200 1685 6370 1705
rect 6400 1805 6570 1825
rect 6400 1775 6410 1805
rect 6440 1775 6570 1805
rect 6400 1735 6570 1775
rect 6400 1705 6410 1735
rect 6440 1705 6570 1735
rect 6400 1685 6570 1705
rect -200 1620 -30 1640
rect -200 1590 -190 1620
rect -160 1590 -30 1620
rect -200 1550 -30 1590
rect -200 1520 -190 1550
rect -160 1520 -30 1550
rect -200 1500 -30 1520
rect 0 1620 170 1640
rect 0 1590 10 1620
rect 40 1590 170 1620
rect 0 1550 170 1590
rect 0 1520 10 1550
rect 40 1520 170 1550
rect 0 1500 170 1520
rect 200 1620 370 1640
rect 200 1590 210 1620
rect 240 1590 370 1620
rect 200 1550 370 1590
rect 200 1520 210 1550
rect 240 1520 370 1550
rect 200 1500 370 1520
rect 400 1620 570 1640
rect 400 1590 410 1620
rect 440 1590 570 1620
rect 400 1550 570 1590
rect 400 1520 410 1550
rect 440 1520 570 1550
rect 400 1500 570 1520
rect 600 1620 770 1640
rect 600 1590 610 1620
rect 640 1590 770 1620
rect 600 1550 770 1590
rect 600 1520 610 1550
rect 640 1520 770 1550
rect 600 1500 770 1520
rect 800 1620 970 1640
rect 800 1590 810 1620
rect 840 1590 970 1620
rect 800 1550 970 1590
rect 800 1520 810 1550
rect 840 1520 970 1550
rect 800 1500 970 1520
rect 1000 1620 1170 1640
rect 1000 1590 1010 1620
rect 1040 1590 1170 1620
rect 1000 1550 1170 1590
rect 1000 1520 1010 1550
rect 1040 1520 1170 1550
rect 1000 1500 1170 1520
rect 1200 1620 1370 1640
rect 1200 1590 1210 1620
rect 1240 1590 1370 1620
rect 1200 1550 1370 1590
rect 1200 1520 1210 1550
rect 1240 1520 1370 1550
rect 1200 1500 1370 1520
rect 1400 1620 1570 1640
rect 1400 1590 1410 1620
rect 1440 1590 1570 1620
rect 1400 1550 1570 1590
rect 1400 1520 1410 1550
rect 1440 1520 1570 1550
rect 1400 1500 1570 1520
rect 1600 1620 1770 1640
rect 1600 1590 1610 1620
rect 1640 1590 1770 1620
rect 1600 1550 1770 1590
rect 1600 1520 1610 1550
rect 1640 1520 1770 1550
rect 1600 1500 1770 1520
rect 1800 1620 1970 1640
rect 1800 1590 1810 1620
rect 1840 1590 1970 1620
rect 1800 1550 1970 1590
rect 1800 1520 1810 1550
rect 1840 1520 1970 1550
rect 1800 1500 1970 1520
rect 2000 1620 2170 1640
rect 2000 1590 2010 1620
rect 2040 1590 2170 1620
rect 2000 1550 2170 1590
rect 2000 1520 2010 1550
rect 2040 1520 2170 1550
rect 2000 1500 2170 1520
rect 2200 1620 2370 1640
rect 2200 1590 2210 1620
rect 2240 1590 2370 1620
rect 2200 1550 2370 1590
rect 2200 1520 2210 1550
rect 2240 1520 2370 1550
rect 2200 1500 2370 1520
rect 2400 1620 2570 1640
rect 2400 1590 2410 1620
rect 2440 1590 2570 1620
rect 2400 1550 2570 1590
rect 2400 1520 2410 1550
rect 2440 1520 2570 1550
rect 2400 1500 2570 1520
rect 2600 1620 2770 1640
rect 2600 1590 2610 1620
rect 2640 1590 2770 1620
rect 2600 1550 2770 1590
rect 2600 1520 2610 1550
rect 2640 1520 2770 1550
rect 2600 1500 2770 1520
rect 2800 1620 2970 1640
rect 2800 1590 2810 1620
rect 2840 1590 2970 1620
rect 2800 1550 2970 1590
rect 2800 1520 2810 1550
rect 2840 1520 2970 1550
rect 2800 1500 2970 1520
rect 3000 1620 3170 1640
rect 3000 1590 3010 1620
rect 3040 1590 3170 1620
rect 3000 1550 3170 1590
rect 3000 1520 3010 1550
rect 3040 1520 3170 1550
rect 3000 1500 3170 1520
rect 3200 1620 3370 1640
rect 3200 1590 3210 1620
rect 3240 1590 3370 1620
rect 3200 1550 3370 1590
rect 3200 1520 3210 1550
rect 3240 1520 3370 1550
rect 3200 1500 3370 1520
rect 3400 1620 3570 1640
rect 3400 1590 3410 1620
rect 3440 1590 3570 1620
rect 3400 1550 3570 1590
rect 3400 1520 3410 1550
rect 3440 1520 3570 1550
rect 3400 1500 3570 1520
rect 3600 1620 3770 1640
rect 3600 1590 3610 1620
rect 3640 1590 3770 1620
rect 3600 1550 3770 1590
rect 3600 1520 3610 1550
rect 3640 1520 3770 1550
rect 3600 1500 3770 1520
rect 3800 1620 3970 1640
rect 3800 1590 3810 1620
rect 3840 1590 3970 1620
rect 3800 1550 3970 1590
rect 3800 1520 3810 1550
rect 3840 1520 3970 1550
rect 3800 1500 3970 1520
rect 4000 1620 4170 1640
rect 4000 1590 4010 1620
rect 4040 1590 4170 1620
rect 4000 1550 4170 1590
rect 4000 1520 4010 1550
rect 4040 1520 4170 1550
rect 4000 1500 4170 1520
rect 4200 1620 4370 1640
rect 4200 1590 4210 1620
rect 4240 1590 4370 1620
rect 4200 1550 4370 1590
rect 4200 1520 4210 1550
rect 4240 1520 4370 1550
rect 4200 1500 4370 1520
rect 4400 1620 4570 1640
rect 4400 1590 4410 1620
rect 4440 1590 4570 1620
rect 4400 1550 4570 1590
rect 4400 1520 4410 1550
rect 4440 1520 4570 1550
rect 4400 1500 4570 1520
rect 4600 1620 4770 1640
rect 4600 1590 4610 1620
rect 4640 1590 4770 1620
rect 4600 1550 4770 1590
rect 4600 1520 4610 1550
rect 4640 1520 4770 1550
rect 4600 1500 4770 1520
rect 4800 1620 4970 1640
rect 4800 1590 4810 1620
rect 4840 1590 4970 1620
rect 4800 1550 4970 1590
rect 4800 1520 4810 1550
rect 4840 1520 4970 1550
rect 4800 1500 4970 1520
rect 5000 1620 5170 1640
rect 5000 1590 5010 1620
rect 5040 1590 5170 1620
rect 5000 1550 5170 1590
rect 5000 1520 5010 1550
rect 5040 1520 5170 1550
rect 5000 1500 5170 1520
rect 5200 1620 5370 1640
rect 5200 1590 5210 1620
rect 5240 1590 5370 1620
rect 5200 1550 5370 1590
rect 5200 1520 5210 1550
rect 5240 1520 5370 1550
rect 5200 1500 5370 1520
rect 5400 1620 5570 1640
rect 5400 1590 5410 1620
rect 5440 1590 5570 1620
rect 5400 1550 5570 1590
rect 5400 1520 5410 1550
rect 5440 1520 5570 1550
rect 5400 1500 5570 1520
rect 5600 1620 5770 1640
rect 5600 1590 5610 1620
rect 5640 1590 5770 1620
rect 5600 1550 5770 1590
rect 5600 1520 5610 1550
rect 5640 1520 5770 1550
rect 5600 1500 5770 1520
rect 5800 1620 5970 1640
rect 5800 1590 5810 1620
rect 5840 1590 5970 1620
rect 5800 1550 5970 1590
rect 5800 1520 5810 1550
rect 5840 1520 5970 1550
rect 5800 1500 5970 1520
rect 6000 1620 6170 1640
rect 6000 1590 6010 1620
rect 6040 1590 6170 1620
rect 6000 1550 6170 1590
rect 6000 1520 6010 1550
rect 6040 1520 6170 1550
rect 6000 1500 6170 1520
rect 6200 1620 6370 1640
rect 6200 1590 6210 1620
rect 6240 1590 6370 1620
rect 6200 1550 6370 1590
rect 6200 1520 6210 1550
rect 6240 1520 6370 1550
rect 6200 1500 6370 1520
rect 6400 1620 6570 1640
rect 6400 1590 6410 1620
rect 6440 1590 6570 1620
rect 6400 1550 6570 1590
rect 6400 1520 6410 1550
rect 6440 1520 6570 1550
rect 6400 1500 6570 1520
rect -200 1435 -30 1455
rect -200 1405 -190 1435
rect -160 1405 -30 1435
rect -200 1365 -30 1405
rect -200 1335 -190 1365
rect -160 1335 -30 1365
rect -200 1315 -30 1335
rect 0 1435 170 1455
rect 0 1405 10 1435
rect 40 1405 170 1435
rect 0 1365 170 1405
rect 0 1335 10 1365
rect 40 1335 170 1365
rect 0 1315 170 1335
rect 200 1435 370 1455
rect 200 1405 210 1435
rect 240 1405 370 1435
rect 200 1365 370 1405
rect 200 1335 210 1365
rect 240 1335 370 1365
rect 200 1315 370 1335
rect 400 1435 570 1455
rect 400 1405 410 1435
rect 440 1405 570 1435
rect 400 1365 570 1405
rect 400 1335 410 1365
rect 440 1335 570 1365
rect 400 1315 570 1335
rect 600 1435 770 1455
rect 600 1405 610 1435
rect 640 1405 770 1435
rect 600 1365 770 1405
rect 600 1335 610 1365
rect 640 1335 770 1365
rect 600 1315 770 1335
rect 800 1435 970 1455
rect 800 1405 810 1435
rect 840 1405 970 1435
rect 800 1365 970 1405
rect 800 1335 810 1365
rect 840 1335 970 1365
rect 800 1315 970 1335
rect 1000 1435 1170 1455
rect 1000 1405 1010 1435
rect 1040 1405 1170 1435
rect 1000 1365 1170 1405
rect 1000 1335 1010 1365
rect 1040 1335 1170 1365
rect 1000 1315 1170 1335
rect 1200 1435 1370 1455
rect 1200 1405 1210 1435
rect 1240 1405 1370 1435
rect 1200 1365 1370 1405
rect 1200 1335 1210 1365
rect 1240 1335 1370 1365
rect 1200 1315 1370 1335
rect 1400 1435 1570 1455
rect 1400 1405 1410 1435
rect 1440 1405 1570 1435
rect 1400 1365 1570 1405
rect 1400 1335 1410 1365
rect 1440 1335 1570 1365
rect 1400 1315 1570 1335
rect 1600 1435 1770 1455
rect 1600 1405 1610 1435
rect 1640 1405 1770 1435
rect 1600 1365 1770 1405
rect 1600 1335 1610 1365
rect 1640 1335 1770 1365
rect 1600 1315 1770 1335
rect 1800 1435 1970 1455
rect 1800 1405 1810 1435
rect 1840 1405 1970 1435
rect 1800 1365 1970 1405
rect 1800 1335 1810 1365
rect 1840 1335 1970 1365
rect 1800 1315 1970 1335
rect 2000 1435 2170 1455
rect 2000 1405 2010 1435
rect 2040 1405 2170 1435
rect 2000 1365 2170 1405
rect 2000 1335 2010 1365
rect 2040 1335 2170 1365
rect 2000 1315 2170 1335
rect 2200 1435 2370 1455
rect 2200 1405 2210 1435
rect 2240 1405 2370 1435
rect 2200 1365 2370 1405
rect 2200 1335 2210 1365
rect 2240 1335 2370 1365
rect 2200 1315 2370 1335
rect 2400 1435 2570 1455
rect 2400 1405 2410 1435
rect 2440 1405 2570 1435
rect 2400 1365 2570 1405
rect 2400 1335 2410 1365
rect 2440 1335 2570 1365
rect 2400 1315 2570 1335
rect 2600 1435 2770 1455
rect 2600 1405 2610 1435
rect 2640 1405 2770 1435
rect 2600 1365 2770 1405
rect 2600 1335 2610 1365
rect 2640 1335 2770 1365
rect 2600 1315 2770 1335
rect 2800 1435 2970 1455
rect 2800 1405 2810 1435
rect 2840 1405 2970 1435
rect 2800 1365 2970 1405
rect 2800 1335 2810 1365
rect 2840 1335 2970 1365
rect 2800 1315 2970 1335
rect 3000 1435 3170 1455
rect 3000 1405 3010 1435
rect 3040 1405 3170 1435
rect 3000 1365 3170 1405
rect 3000 1335 3010 1365
rect 3040 1335 3170 1365
rect 3000 1315 3170 1335
rect 3200 1435 3370 1455
rect 3200 1405 3210 1435
rect 3240 1405 3370 1435
rect 3200 1365 3370 1405
rect 3200 1335 3210 1365
rect 3240 1335 3370 1365
rect 3200 1315 3370 1335
rect 3400 1435 3570 1455
rect 3400 1405 3410 1435
rect 3440 1405 3570 1435
rect 3400 1365 3570 1405
rect 3400 1335 3410 1365
rect 3440 1335 3570 1365
rect 3400 1315 3570 1335
rect 3600 1435 3770 1455
rect 3600 1405 3610 1435
rect 3640 1405 3770 1435
rect 3600 1365 3770 1405
rect 3600 1335 3610 1365
rect 3640 1335 3770 1365
rect 3600 1315 3770 1335
rect 3800 1435 3970 1455
rect 3800 1405 3810 1435
rect 3840 1405 3970 1435
rect 3800 1365 3970 1405
rect 3800 1335 3810 1365
rect 3840 1335 3970 1365
rect 3800 1315 3970 1335
rect 4000 1435 4170 1455
rect 4000 1405 4010 1435
rect 4040 1405 4170 1435
rect 4000 1365 4170 1405
rect 4000 1335 4010 1365
rect 4040 1335 4170 1365
rect 4000 1315 4170 1335
rect 4200 1435 4370 1455
rect 4200 1405 4210 1435
rect 4240 1405 4370 1435
rect 4200 1365 4370 1405
rect 4200 1335 4210 1365
rect 4240 1335 4370 1365
rect 4200 1315 4370 1335
rect 4400 1435 4570 1455
rect 4400 1405 4410 1435
rect 4440 1405 4570 1435
rect 4400 1365 4570 1405
rect 4400 1335 4410 1365
rect 4440 1335 4570 1365
rect 4400 1315 4570 1335
rect 4600 1435 4770 1455
rect 4600 1405 4610 1435
rect 4640 1405 4770 1435
rect 4600 1365 4770 1405
rect 4600 1335 4610 1365
rect 4640 1335 4770 1365
rect 4600 1315 4770 1335
rect 4800 1435 4970 1455
rect 4800 1405 4810 1435
rect 4840 1405 4970 1435
rect 4800 1365 4970 1405
rect 4800 1335 4810 1365
rect 4840 1335 4970 1365
rect 4800 1315 4970 1335
rect 5000 1435 5170 1455
rect 5000 1405 5010 1435
rect 5040 1405 5170 1435
rect 5000 1365 5170 1405
rect 5000 1335 5010 1365
rect 5040 1335 5170 1365
rect 5000 1315 5170 1335
rect 5200 1435 5370 1455
rect 5200 1405 5210 1435
rect 5240 1405 5370 1435
rect 5200 1365 5370 1405
rect 5200 1335 5210 1365
rect 5240 1335 5370 1365
rect 5200 1315 5370 1335
rect 5400 1435 5570 1455
rect 5400 1405 5410 1435
rect 5440 1405 5570 1435
rect 5400 1365 5570 1405
rect 5400 1335 5410 1365
rect 5440 1335 5570 1365
rect 5400 1315 5570 1335
rect 5600 1435 5770 1455
rect 5600 1405 5610 1435
rect 5640 1405 5770 1435
rect 5600 1365 5770 1405
rect 5600 1335 5610 1365
rect 5640 1335 5770 1365
rect 5600 1315 5770 1335
rect 5800 1435 5970 1455
rect 5800 1405 5810 1435
rect 5840 1405 5970 1435
rect 5800 1365 5970 1405
rect 5800 1335 5810 1365
rect 5840 1335 5970 1365
rect 5800 1315 5970 1335
rect 6000 1435 6170 1455
rect 6000 1405 6010 1435
rect 6040 1405 6170 1435
rect 6000 1365 6170 1405
rect 6000 1335 6010 1365
rect 6040 1335 6170 1365
rect 6000 1315 6170 1335
rect 6200 1435 6370 1455
rect 6200 1405 6210 1435
rect 6240 1405 6370 1435
rect 6200 1365 6370 1405
rect 6200 1335 6210 1365
rect 6240 1335 6370 1365
rect 6200 1315 6370 1335
rect 6400 1435 6570 1455
rect 6400 1405 6410 1435
rect 6440 1405 6570 1435
rect 6400 1365 6570 1405
rect 6400 1335 6410 1365
rect 6440 1335 6570 1365
rect 6400 1315 6570 1335
rect -200 1250 -30 1270
rect -200 1220 -190 1250
rect -160 1220 -30 1250
rect -200 1180 -30 1220
rect -200 1150 -190 1180
rect -160 1150 -30 1180
rect -200 1130 -30 1150
rect 0 1250 170 1270
rect 0 1220 10 1250
rect 40 1220 170 1250
rect 0 1180 170 1220
rect 0 1150 10 1180
rect 40 1150 170 1180
rect 0 1130 170 1150
rect 200 1250 370 1270
rect 200 1220 210 1250
rect 240 1220 370 1250
rect 200 1180 370 1220
rect 200 1150 210 1180
rect 240 1150 370 1180
rect 200 1130 370 1150
rect 400 1250 570 1270
rect 400 1220 410 1250
rect 440 1220 570 1250
rect 400 1180 570 1220
rect 400 1150 410 1180
rect 440 1150 570 1180
rect 400 1130 570 1150
rect 600 1250 770 1270
rect 600 1220 610 1250
rect 640 1220 770 1250
rect 600 1180 770 1220
rect 600 1150 610 1180
rect 640 1150 770 1180
rect 600 1130 770 1150
rect 800 1250 970 1270
rect 800 1220 810 1250
rect 840 1220 970 1250
rect 800 1180 970 1220
rect 800 1150 810 1180
rect 840 1150 970 1180
rect 800 1130 970 1150
rect 1000 1250 1170 1270
rect 1000 1220 1010 1250
rect 1040 1220 1170 1250
rect 1000 1180 1170 1220
rect 1000 1150 1010 1180
rect 1040 1150 1170 1180
rect 1000 1130 1170 1150
rect 1200 1250 1370 1270
rect 1200 1220 1210 1250
rect 1240 1220 1370 1250
rect 1200 1180 1370 1220
rect 1200 1150 1210 1180
rect 1240 1150 1370 1180
rect 1200 1130 1370 1150
rect 1400 1250 1570 1270
rect 1400 1220 1410 1250
rect 1440 1220 1570 1250
rect 1400 1180 1570 1220
rect 1400 1150 1410 1180
rect 1440 1150 1570 1180
rect 1400 1130 1570 1150
rect 1600 1250 1770 1270
rect 1600 1220 1610 1250
rect 1640 1220 1770 1250
rect 1600 1180 1770 1220
rect 1600 1150 1610 1180
rect 1640 1150 1770 1180
rect 1600 1130 1770 1150
rect 1800 1250 1970 1270
rect 1800 1220 1810 1250
rect 1840 1220 1970 1250
rect 1800 1180 1970 1220
rect 1800 1150 1810 1180
rect 1840 1150 1970 1180
rect 1800 1130 1970 1150
rect 2000 1250 2170 1270
rect 2000 1220 2010 1250
rect 2040 1220 2170 1250
rect 2000 1180 2170 1220
rect 2000 1150 2010 1180
rect 2040 1150 2170 1180
rect 2000 1130 2170 1150
rect 2200 1250 2370 1270
rect 2200 1220 2210 1250
rect 2240 1220 2370 1250
rect 2200 1180 2370 1220
rect 2200 1150 2210 1180
rect 2240 1150 2370 1180
rect 2200 1130 2370 1150
rect 2400 1250 2570 1270
rect 2400 1220 2410 1250
rect 2440 1220 2570 1250
rect 2400 1180 2570 1220
rect 2400 1150 2410 1180
rect 2440 1150 2570 1180
rect 2400 1130 2570 1150
rect 2600 1250 2770 1270
rect 2600 1220 2610 1250
rect 2640 1220 2770 1250
rect 2600 1180 2770 1220
rect 2600 1150 2610 1180
rect 2640 1150 2770 1180
rect 2600 1130 2770 1150
rect 2800 1250 2970 1270
rect 2800 1220 2810 1250
rect 2840 1220 2970 1250
rect 2800 1180 2970 1220
rect 2800 1150 2810 1180
rect 2840 1150 2970 1180
rect 2800 1130 2970 1150
rect 3000 1250 3170 1270
rect 3000 1220 3010 1250
rect 3040 1220 3170 1250
rect 3000 1180 3170 1220
rect 3000 1150 3010 1180
rect 3040 1150 3170 1180
rect 3000 1130 3170 1150
rect 3200 1250 3370 1270
rect 3200 1220 3210 1250
rect 3240 1220 3370 1250
rect 3200 1180 3370 1220
rect 3200 1150 3210 1180
rect 3240 1150 3370 1180
rect 3200 1130 3370 1150
rect 3400 1250 3570 1270
rect 3400 1220 3410 1250
rect 3440 1220 3570 1250
rect 3400 1180 3570 1220
rect 3400 1150 3410 1180
rect 3440 1150 3570 1180
rect 3400 1130 3570 1150
rect 3600 1250 3770 1270
rect 3600 1220 3610 1250
rect 3640 1220 3770 1250
rect 3600 1180 3770 1220
rect 3600 1150 3610 1180
rect 3640 1150 3770 1180
rect 3600 1130 3770 1150
rect 3800 1250 3970 1270
rect 3800 1220 3810 1250
rect 3840 1220 3970 1250
rect 3800 1180 3970 1220
rect 3800 1150 3810 1180
rect 3840 1150 3970 1180
rect 3800 1130 3970 1150
rect 4000 1250 4170 1270
rect 4000 1220 4010 1250
rect 4040 1220 4170 1250
rect 4000 1180 4170 1220
rect 4000 1150 4010 1180
rect 4040 1150 4170 1180
rect 4000 1130 4170 1150
rect 4200 1250 4370 1270
rect 4200 1220 4210 1250
rect 4240 1220 4370 1250
rect 4200 1180 4370 1220
rect 4200 1150 4210 1180
rect 4240 1150 4370 1180
rect 4200 1130 4370 1150
rect 4400 1250 4570 1270
rect 4400 1220 4410 1250
rect 4440 1220 4570 1250
rect 4400 1180 4570 1220
rect 4400 1150 4410 1180
rect 4440 1150 4570 1180
rect 4400 1130 4570 1150
rect 4600 1250 4770 1270
rect 4600 1220 4610 1250
rect 4640 1220 4770 1250
rect 4600 1180 4770 1220
rect 4600 1150 4610 1180
rect 4640 1150 4770 1180
rect 4600 1130 4770 1150
rect 4800 1250 4970 1270
rect 4800 1220 4810 1250
rect 4840 1220 4970 1250
rect 4800 1180 4970 1220
rect 4800 1150 4810 1180
rect 4840 1150 4970 1180
rect 4800 1130 4970 1150
rect 5000 1250 5170 1270
rect 5000 1220 5010 1250
rect 5040 1220 5170 1250
rect 5000 1180 5170 1220
rect 5000 1150 5010 1180
rect 5040 1150 5170 1180
rect 5000 1130 5170 1150
rect 5200 1250 5370 1270
rect 5200 1220 5210 1250
rect 5240 1220 5370 1250
rect 5200 1180 5370 1220
rect 5200 1150 5210 1180
rect 5240 1150 5370 1180
rect 5200 1130 5370 1150
rect 5400 1250 5570 1270
rect 5400 1220 5410 1250
rect 5440 1220 5570 1250
rect 5400 1180 5570 1220
rect 5400 1150 5410 1180
rect 5440 1150 5570 1180
rect 5400 1130 5570 1150
rect 5600 1250 5770 1270
rect 5600 1220 5610 1250
rect 5640 1220 5770 1250
rect 5600 1180 5770 1220
rect 5600 1150 5610 1180
rect 5640 1150 5770 1180
rect 5600 1130 5770 1150
rect 5800 1250 5970 1270
rect 5800 1220 5810 1250
rect 5840 1220 5970 1250
rect 5800 1180 5970 1220
rect 5800 1150 5810 1180
rect 5840 1150 5970 1180
rect 5800 1130 5970 1150
rect 6000 1250 6170 1270
rect 6000 1220 6010 1250
rect 6040 1220 6170 1250
rect 6000 1180 6170 1220
rect 6000 1150 6010 1180
rect 6040 1150 6170 1180
rect 6000 1130 6170 1150
rect 6200 1250 6370 1270
rect 6200 1220 6210 1250
rect 6240 1220 6370 1250
rect 6200 1180 6370 1220
rect 6200 1150 6210 1180
rect 6240 1150 6370 1180
rect 6200 1130 6370 1150
rect 6400 1250 6570 1270
rect 6400 1220 6410 1250
rect 6440 1220 6570 1250
rect 6400 1180 6570 1220
rect 6400 1150 6410 1180
rect 6440 1150 6570 1180
rect 6400 1130 6570 1150
rect -200 1065 -30 1085
rect -200 1035 -190 1065
rect -160 1035 -30 1065
rect -200 995 -30 1035
rect -200 965 -190 995
rect -160 965 -30 995
rect -200 945 -30 965
rect 0 1065 170 1085
rect 0 1035 10 1065
rect 40 1035 170 1065
rect 0 995 170 1035
rect 0 965 10 995
rect 40 965 170 995
rect 0 945 170 965
rect 200 1065 370 1085
rect 200 1035 210 1065
rect 240 1035 370 1065
rect 200 995 370 1035
rect 200 965 210 995
rect 240 965 370 995
rect 200 945 370 965
rect 400 1065 570 1085
rect 400 1035 410 1065
rect 440 1035 570 1065
rect 400 995 570 1035
rect 400 965 410 995
rect 440 965 570 995
rect 400 945 570 965
rect 600 1065 770 1085
rect 600 1035 610 1065
rect 640 1035 770 1065
rect 600 995 770 1035
rect 600 965 610 995
rect 640 965 770 995
rect 600 945 770 965
rect 800 1065 970 1085
rect 800 1035 810 1065
rect 840 1035 970 1065
rect 800 995 970 1035
rect 800 965 810 995
rect 840 965 970 995
rect 800 945 970 965
rect 1000 1065 1170 1085
rect 1000 1035 1010 1065
rect 1040 1035 1170 1065
rect 1000 995 1170 1035
rect 1000 965 1010 995
rect 1040 965 1170 995
rect 1000 945 1170 965
rect 1200 1065 1370 1085
rect 1200 1035 1210 1065
rect 1240 1035 1370 1065
rect 1200 995 1370 1035
rect 1200 965 1210 995
rect 1240 965 1370 995
rect 1200 945 1370 965
rect 1400 1065 1570 1085
rect 1400 1035 1410 1065
rect 1440 1035 1570 1065
rect 1400 995 1570 1035
rect 1400 965 1410 995
rect 1440 965 1570 995
rect 1400 945 1570 965
rect 1600 1065 1770 1085
rect 1600 1035 1610 1065
rect 1640 1035 1770 1065
rect 1600 995 1770 1035
rect 1600 965 1610 995
rect 1640 965 1770 995
rect 1600 945 1770 965
rect 1800 1065 1970 1085
rect 1800 1035 1810 1065
rect 1840 1035 1970 1065
rect 1800 995 1970 1035
rect 1800 965 1810 995
rect 1840 965 1970 995
rect 1800 945 1970 965
rect 2000 1065 2170 1085
rect 2000 1035 2010 1065
rect 2040 1035 2170 1065
rect 2000 995 2170 1035
rect 2000 965 2010 995
rect 2040 965 2170 995
rect 2000 945 2170 965
rect 2200 1065 2370 1085
rect 2200 1035 2210 1065
rect 2240 1035 2370 1065
rect 2200 995 2370 1035
rect 2200 965 2210 995
rect 2240 965 2370 995
rect 2200 945 2370 965
rect 2400 1065 2570 1085
rect 2400 1035 2410 1065
rect 2440 1035 2570 1065
rect 2400 995 2570 1035
rect 2400 965 2410 995
rect 2440 965 2570 995
rect 2400 945 2570 965
rect 2600 1065 2770 1085
rect 2600 1035 2610 1065
rect 2640 1035 2770 1065
rect 2600 995 2770 1035
rect 2600 965 2610 995
rect 2640 965 2770 995
rect 2600 945 2770 965
rect 2800 1065 2970 1085
rect 2800 1035 2810 1065
rect 2840 1035 2970 1065
rect 2800 995 2970 1035
rect 2800 965 2810 995
rect 2840 965 2970 995
rect 2800 945 2970 965
rect 3000 1065 3170 1085
rect 3000 1035 3010 1065
rect 3040 1035 3170 1065
rect 3000 995 3170 1035
rect 3000 965 3010 995
rect 3040 965 3170 995
rect 3000 945 3170 965
rect 3200 1065 3370 1085
rect 3200 1035 3210 1065
rect 3240 1035 3370 1065
rect 3200 995 3370 1035
rect 3200 965 3210 995
rect 3240 965 3370 995
rect 3200 945 3370 965
rect 3400 1065 3570 1085
rect 3400 1035 3410 1065
rect 3440 1035 3570 1065
rect 3400 995 3570 1035
rect 3400 965 3410 995
rect 3440 965 3570 995
rect 3400 945 3570 965
rect 3600 1065 3770 1085
rect 3600 1035 3610 1065
rect 3640 1035 3770 1065
rect 3600 995 3770 1035
rect 3600 965 3610 995
rect 3640 965 3770 995
rect 3600 945 3770 965
rect 3800 1065 3970 1085
rect 3800 1035 3810 1065
rect 3840 1035 3970 1065
rect 3800 995 3970 1035
rect 3800 965 3810 995
rect 3840 965 3970 995
rect 3800 945 3970 965
rect 4000 1065 4170 1085
rect 4000 1035 4010 1065
rect 4040 1035 4170 1065
rect 4000 995 4170 1035
rect 4000 965 4010 995
rect 4040 965 4170 995
rect 4000 945 4170 965
rect 4200 1065 4370 1085
rect 4200 1035 4210 1065
rect 4240 1035 4370 1065
rect 4200 995 4370 1035
rect 4200 965 4210 995
rect 4240 965 4370 995
rect 4200 945 4370 965
rect 4400 1065 4570 1085
rect 4400 1035 4410 1065
rect 4440 1035 4570 1065
rect 4400 995 4570 1035
rect 4400 965 4410 995
rect 4440 965 4570 995
rect 4400 945 4570 965
rect 4600 1065 4770 1085
rect 4600 1035 4610 1065
rect 4640 1035 4770 1065
rect 4600 995 4770 1035
rect 4600 965 4610 995
rect 4640 965 4770 995
rect 4600 945 4770 965
rect 4800 1065 4970 1085
rect 4800 1035 4810 1065
rect 4840 1035 4970 1065
rect 4800 995 4970 1035
rect 4800 965 4810 995
rect 4840 965 4970 995
rect 4800 945 4970 965
rect 5000 1065 5170 1085
rect 5000 1035 5010 1065
rect 5040 1035 5170 1065
rect 5000 995 5170 1035
rect 5000 965 5010 995
rect 5040 965 5170 995
rect 5000 945 5170 965
rect 5200 1065 5370 1085
rect 5200 1035 5210 1065
rect 5240 1035 5370 1065
rect 5200 995 5370 1035
rect 5200 965 5210 995
rect 5240 965 5370 995
rect 5200 945 5370 965
rect 5400 1065 5570 1085
rect 5400 1035 5410 1065
rect 5440 1035 5570 1065
rect 5400 995 5570 1035
rect 5400 965 5410 995
rect 5440 965 5570 995
rect 5400 945 5570 965
rect 5600 1065 5770 1085
rect 5600 1035 5610 1065
rect 5640 1035 5770 1065
rect 5600 995 5770 1035
rect 5600 965 5610 995
rect 5640 965 5770 995
rect 5600 945 5770 965
rect 5800 1065 5970 1085
rect 5800 1035 5810 1065
rect 5840 1035 5970 1065
rect 5800 995 5970 1035
rect 5800 965 5810 995
rect 5840 965 5970 995
rect 5800 945 5970 965
rect 6000 1065 6170 1085
rect 6000 1035 6010 1065
rect 6040 1035 6170 1065
rect 6000 995 6170 1035
rect 6000 965 6010 995
rect 6040 965 6170 995
rect 6000 945 6170 965
rect 6200 1065 6370 1085
rect 6200 1035 6210 1065
rect 6240 1035 6370 1065
rect 6200 995 6370 1035
rect 6200 965 6210 995
rect 6240 965 6370 995
rect 6200 945 6370 965
rect 6400 1065 6570 1085
rect 6400 1035 6410 1065
rect 6440 1035 6570 1065
rect 6400 995 6570 1035
rect 6400 965 6410 995
rect 6440 965 6570 995
rect 6400 945 6570 965
rect -200 880 -30 900
rect -200 850 -190 880
rect -160 850 -30 880
rect -200 810 -30 850
rect -200 780 -190 810
rect -160 780 -30 810
rect -200 760 -30 780
rect 0 880 170 900
rect 0 850 10 880
rect 40 850 170 880
rect 0 810 170 850
rect 0 780 10 810
rect 40 780 170 810
rect 0 760 170 780
rect 200 880 370 900
rect 200 850 210 880
rect 240 850 370 880
rect 200 810 370 850
rect 200 780 210 810
rect 240 780 370 810
rect 200 760 370 780
rect 400 880 570 900
rect 400 850 410 880
rect 440 850 570 880
rect 400 810 570 850
rect 400 780 410 810
rect 440 780 570 810
rect 400 760 570 780
rect 600 880 770 900
rect 600 850 610 880
rect 640 850 770 880
rect 600 810 770 850
rect 600 780 610 810
rect 640 780 770 810
rect 600 760 770 780
rect 800 880 970 900
rect 800 850 810 880
rect 840 850 970 880
rect 800 810 970 850
rect 800 780 810 810
rect 840 780 970 810
rect 800 760 970 780
rect 1000 880 1170 900
rect 1000 850 1010 880
rect 1040 850 1170 880
rect 1000 810 1170 850
rect 1000 780 1010 810
rect 1040 780 1170 810
rect 1000 760 1170 780
rect 1200 880 1370 900
rect 1200 850 1210 880
rect 1240 850 1370 880
rect 1200 810 1370 850
rect 1200 780 1210 810
rect 1240 780 1370 810
rect 1200 760 1370 780
rect 1400 880 1570 900
rect 1400 850 1410 880
rect 1440 850 1570 880
rect 1400 810 1570 850
rect 1400 780 1410 810
rect 1440 780 1570 810
rect 1400 760 1570 780
rect 1600 880 1770 900
rect 1600 850 1610 880
rect 1640 850 1770 880
rect 1600 810 1770 850
rect 1600 780 1610 810
rect 1640 780 1770 810
rect 1600 760 1770 780
rect 1800 880 1970 900
rect 1800 850 1810 880
rect 1840 850 1970 880
rect 1800 810 1970 850
rect 1800 780 1810 810
rect 1840 780 1970 810
rect 1800 760 1970 780
rect 2000 880 2170 900
rect 2000 850 2010 880
rect 2040 850 2170 880
rect 2000 810 2170 850
rect 2000 780 2010 810
rect 2040 780 2170 810
rect 2000 760 2170 780
rect 2200 880 2370 900
rect 2200 850 2210 880
rect 2240 850 2370 880
rect 2200 810 2370 850
rect 2200 780 2210 810
rect 2240 780 2370 810
rect 2200 760 2370 780
rect 2400 880 2570 900
rect 2400 850 2410 880
rect 2440 850 2570 880
rect 2400 810 2570 850
rect 2400 780 2410 810
rect 2440 780 2570 810
rect 2400 760 2570 780
rect 2600 880 2770 900
rect 2600 850 2610 880
rect 2640 850 2770 880
rect 2600 810 2770 850
rect 2600 780 2610 810
rect 2640 780 2770 810
rect 2600 760 2770 780
rect 2800 880 2970 900
rect 2800 850 2810 880
rect 2840 850 2970 880
rect 2800 810 2970 850
rect 2800 780 2810 810
rect 2840 780 2970 810
rect 2800 760 2970 780
rect 3000 880 3170 900
rect 3000 850 3010 880
rect 3040 850 3170 880
rect 3000 810 3170 850
rect 3000 780 3010 810
rect 3040 780 3170 810
rect 3000 760 3170 780
rect 3200 880 3370 900
rect 3200 850 3210 880
rect 3240 850 3370 880
rect 3200 810 3370 850
rect 3200 780 3210 810
rect 3240 780 3370 810
rect 3200 760 3370 780
rect 3400 880 3570 900
rect 3400 850 3410 880
rect 3440 850 3570 880
rect 3400 810 3570 850
rect 3400 780 3410 810
rect 3440 780 3570 810
rect 3400 760 3570 780
rect 3600 880 3770 900
rect 3600 850 3610 880
rect 3640 850 3770 880
rect 3600 810 3770 850
rect 3600 780 3610 810
rect 3640 780 3770 810
rect 3600 760 3770 780
rect 3800 880 3970 900
rect 3800 850 3810 880
rect 3840 850 3970 880
rect 3800 810 3970 850
rect 3800 780 3810 810
rect 3840 780 3970 810
rect 3800 760 3970 780
rect 4000 880 4170 900
rect 4000 850 4010 880
rect 4040 850 4170 880
rect 4000 810 4170 850
rect 4000 780 4010 810
rect 4040 780 4170 810
rect 4000 760 4170 780
rect 4200 880 4370 900
rect 4200 850 4210 880
rect 4240 850 4370 880
rect 4200 810 4370 850
rect 4200 780 4210 810
rect 4240 780 4370 810
rect 4200 760 4370 780
rect 4400 880 4570 900
rect 4400 850 4410 880
rect 4440 850 4570 880
rect 4400 810 4570 850
rect 4400 780 4410 810
rect 4440 780 4570 810
rect 4400 760 4570 780
rect 4600 880 4770 900
rect 4600 850 4610 880
rect 4640 850 4770 880
rect 4600 810 4770 850
rect 4600 780 4610 810
rect 4640 780 4770 810
rect 4600 760 4770 780
rect 4800 880 4970 900
rect 4800 850 4810 880
rect 4840 850 4970 880
rect 4800 810 4970 850
rect 4800 780 4810 810
rect 4840 780 4970 810
rect 4800 760 4970 780
rect 5000 880 5170 900
rect 5000 850 5010 880
rect 5040 850 5170 880
rect 5000 810 5170 850
rect 5000 780 5010 810
rect 5040 780 5170 810
rect 5000 760 5170 780
rect 5200 880 5370 900
rect 5200 850 5210 880
rect 5240 850 5370 880
rect 5200 810 5370 850
rect 5200 780 5210 810
rect 5240 780 5370 810
rect 5200 760 5370 780
rect 5400 880 5570 900
rect 5400 850 5410 880
rect 5440 850 5570 880
rect 5400 810 5570 850
rect 5400 780 5410 810
rect 5440 780 5570 810
rect 5400 760 5570 780
rect 5600 880 5770 900
rect 5600 850 5610 880
rect 5640 850 5770 880
rect 5600 810 5770 850
rect 5600 780 5610 810
rect 5640 780 5770 810
rect 5600 760 5770 780
rect 5800 880 5970 900
rect 5800 850 5810 880
rect 5840 850 5970 880
rect 5800 810 5970 850
rect 5800 780 5810 810
rect 5840 780 5970 810
rect 5800 760 5970 780
rect 6000 880 6170 900
rect 6000 850 6010 880
rect 6040 850 6170 880
rect 6000 810 6170 850
rect 6000 780 6010 810
rect 6040 780 6170 810
rect 6000 760 6170 780
rect 6200 880 6370 900
rect 6200 850 6210 880
rect 6240 850 6370 880
rect 6200 810 6370 850
rect 6200 780 6210 810
rect 6240 780 6370 810
rect 6200 760 6370 780
rect 6400 880 6570 900
rect 6400 850 6410 880
rect 6440 850 6570 880
rect 6400 810 6570 850
rect 6400 780 6410 810
rect 6440 780 6570 810
rect 6400 760 6570 780
rect -200 695 -30 715
rect -200 665 -190 695
rect -160 665 -30 695
rect -200 625 -30 665
rect -200 595 -190 625
rect -160 595 -30 625
rect -200 575 -30 595
rect 0 695 170 715
rect 0 665 10 695
rect 40 665 170 695
rect 0 625 170 665
rect 0 595 10 625
rect 40 595 170 625
rect 0 575 170 595
rect 200 695 370 715
rect 200 665 210 695
rect 240 665 370 695
rect 200 625 370 665
rect 200 595 210 625
rect 240 595 370 625
rect 200 575 370 595
rect 400 695 570 715
rect 400 665 410 695
rect 440 665 570 695
rect 400 625 570 665
rect 400 595 410 625
rect 440 595 570 625
rect 400 575 570 595
rect 600 695 770 715
rect 600 665 610 695
rect 640 665 770 695
rect 600 625 770 665
rect 600 595 610 625
rect 640 595 770 625
rect 600 575 770 595
rect 800 695 970 715
rect 800 665 810 695
rect 840 665 970 695
rect 800 625 970 665
rect 800 595 810 625
rect 840 595 970 625
rect 800 575 970 595
rect 1000 695 1170 715
rect 1000 665 1010 695
rect 1040 665 1170 695
rect 1000 625 1170 665
rect 1000 595 1010 625
rect 1040 595 1170 625
rect 1000 575 1170 595
rect 1200 695 1370 715
rect 1200 665 1210 695
rect 1240 665 1370 695
rect 1200 625 1370 665
rect 1200 595 1210 625
rect 1240 595 1370 625
rect 1200 575 1370 595
rect 1400 695 1570 715
rect 1400 665 1410 695
rect 1440 665 1570 695
rect 1400 625 1570 665
rect 1400 595 1410 625
rect 1440 595 1570 625
rect 1400 575 1570 595
rect 1600 695 1770 715
rect 1600 665 1610 695
rect 1640 665 1770 695
rect 1600 625 1770 665
rect 1600 595 1610 625
rect 1640 595 1770 625
rect 1600 575 1770 595
rect 1800 695 1970 715
rect 1800 665 1810 695
rect 1840 665 1970 695
rect 1800 625 1970 665
rect 1800 595 1810 625
rect 1840 595 1970 625
rect 1800 575 1970 595
rect 2000 695 2170 715
rect 2000 665 2010 695
rect 2040 665 2170 695
rect 2000 625 2170 665
rect 2000 595 2010 625
rect 2040 595 2170 625
rect 2000 575 2170 595
rect 2200 695 2370 715
rect 2200 665 2210 695
rect 2240 665 2370 695
rect 2200 625 2370 665
rect 2200 595 2210 625
rect 2240 595 2370 625
rect 2200 575 2370 595
rect 2400 695 2570 715
rect 2400 665 2410 695
rect 2440 665 2570 695
rect 2400 625 2570 665
rect 2400 595 2410 625
rect 2440 595 2570 625
rect 2400 575 2570 595
rect 2600 695 2770 715
rect 2600 665 2610 695
rect 2640 665 2770 695
rect 2600 625 2770 665
rect 2600 595 2610 625
rect 2640 595 2770 625
rect 2600 575 2770 595
rect 2800 695 2970 715
rect 2800 665 2810 695
rect 2840 665 2970 695
rect 2800 625 2970 665
rect 2800 595 2810 625
rect 2840 595 2970 625
rect 2800 575 2970 595
rect 3000 695 3170 715
rect 3000 665 3010 695
rect 3040 665 3170 695
rect 3000 625 3170 665
rect 3000 595 3010 625
rect 3040 595 3170 625
rect 3000 575 3170 595
rect 3200 695 3370 715
rect 3200 665 3210 695
rect 3240 665 3370 695
rect 3200 625 3370 665
rect 3200 595 3210 625
rect 3240 595 3370 625
rect 3200 575 3370 595
rect 3400 695 3570 715
rect 3400 665 3410 695
rect 3440 665 3570 695
rect 3400 625 3570 665
rect 3400 595 3410 625
rect 3440 595 3570 625
rect 3400 575 3570 595
rect 3600 695 3770 715
rect 3600 665 3610 695
rect 3640 665 3770 695
rect 3600 625 3770 665
rect 3600 595 3610 625
rect 3640 595 3770 625
rect 3600 575 3770 595
rect 3800 695 3970 715
rect 3800 665 3810 695
rect 3840 665 3970 695
rect 3800 625 3970 665
rect 3800 595 3810 625
rect 3840 595 3970 625
rect 3800 575 3970 595
rect 4000 695 4170 715
rect 4000 665 4010 695
rect 4040 665 4170 695
rect 4000 625 4170 665
rect 4000 595 4010 625
rect 4040 595 4170 625
rect 4000 575 4170 595
rect 4200 695 4370 715
rect 4200 665 4210 695
rect 4240 665 4370 695
rect 4200 625 4370 665
rect 4200 595 4210 625
rect 4240 595 4370 625
rect 4200 575 4370 595
rect 4400 695 4570 715
rect 4400 665 4410 695
rect 4440 665 4570 695
rect 4400 625 4570 665
rect 4400 595 4410 625
rect 4440 595 4570 625
rect 4400 575 4570 595
rect 4600 695 4770 715
rect 4600 665 4610 695
rect 4640 665 4770 695
rect 4600 625 4770 665
rect 4600 595 4610 625
rect 4640 595 4770 625
rect 4600 575 4770 595
rect 4800 695 4970 715
rect 4800 665 4810 695
rect 4840 665 4970 695
rect 4800 625 4970 665
rect 4800 595 4810 625
rect 4840 595 4970 625
rect 4800 575 4970 595
rect 5000 695 5170 715
rect 5000 665 5010 695
rect 5040 665 5170 695
rect 5000 625 5170 665
rect 5000 595 5010 625
rect 5040 595 5170 625
rect 5000 575 5170 595
rect 5200 695 5370 715
rect 5200 665 5210 695
rect 5240 665 5370 695
rect 5200 625 5370 665
rect 5200 595 5210 625
rect 5240 595 5370 625
rect 5200 575 5370 595
rect 5400 695 5570 715
rect 5400 665 5410 695
rect 5440 665 5570 695
rect 5400 625 5570 665
rect 5400 595 5410 625
rect 5440 595 5570 625
rect 5400 575 5570 595
rect 5600 695 5770 715
rect 5600 665 5610 695
rect 5640 665 5770 695
rect 5600 625 5770 665
rect 5600 595 5610 625
rect 5640 595 5770 625
rect 5600 575 5770 595
rect 5800 695 5970 715
rect 5800 665 5810 695
rect 5840 665 5970 695
rect 5800 625 5970 665
rect 5800 595 5810 625
rect 5840 595 5970 625
rect 5800 575 5970 595
rect 6000 695 6170 715
rect 6000 665 6010 695
rect 6040 665 6170 695
rect 6000 625 6170 665
rect 6000 595 6010 625
rect 6040 595 6170 625
rect 6000 575 6170 595
rect 6200 695 6370 715
rect 6200 665 6210 695
rect 6240 665 6370 695
rect 6200 625 6370 665
rect 6200 595 6210 625
rect 6240 595 6370 625
rect 6200 575 6370 595
rect 6400 695 6570 715
rect 6400 665 6410 695
rect 6440 665 6570 695
rect 6400 625 6570 665
rect 6400 595 6410 625
rect 6440 595 6570 625
rect 6400 575 6570 595
rect -200 510 -30 530
rect -200 480 -190 510
rect -160 480 -30 510
rect -200 440 -30 480
rect -200 410 -190 440
rect -160 410 -30 440
rect -200 390 -30 410
rect 0 510 170 530
rect 0 480 10 510
rect 40 480 170 510
rect 0 440 170 480
rect 0 410 10 440
rect 40 410 170 440
rect 0 390 170 410
rect 200 510 370 530
rect 200 480 210 510
rect 240 480 370 510
rect 200 440 370 480
rect 200 410 210 440
rect 240 410 370 440
rect 200 390 370 410
rect 400 510 570 530
rect 400 480 410 510
rect 440 480 570 510
rect 400 440 570 480
rect 400 410 410 440
rect 440 410 570 440
rect 400 390 570 410
rect 600 510 770 530
rect 600 480 610 510
rect 640 480 770 510
rect 600 440 770 480
rect 600 410 610 440
rect 640 410 770 440
rect 600 390 770 410
rect 800 510 970 530
rect 800 480 810 510
rect 840 480 970 510
rect 800 440 970 480
rect 800 410 810 440
rect 840 410 970 440
rect 800 390 970 410
rect 1000 510 1170 530
rect 1000 480 1010 510
rect 1040 480 1170 510
rect 1000 440 1170 480
rect 1000 410 1010 440
rect 1040 410 1170 440
rect 1000 390 1170 410
rect 1200 510 1370 530
rect 1200 480 1210 510
rect 1240 480 1370 510
rect 1200 440 1370 480
rect 1200 410 1210 440
rect 1240 410 1370 440
rect 1200 390 1370 410
rect 1400 510 1570 530
rect 1400 480 1410 510
rect 1440 480 1570 510
rect 1400 440 1570 480
rect 1400 410 1410 440
rect 1440 410 1570 440
rect 1400 390 1570 410
rect 1600 510 1770 530
rect 1600 480 1610 510
rect 1640 480 1770 510
rect 1600 440 1770 480
rect 1600 410 1610 440
rect 1640 410 1770 440
rect 1600 390 1770 410
rect 1800 510 1970 530
rect 1800 480 1810 510
rect 1840 480 1970 510
rect 1800 440 1970 480
rect 1800 410 1810 440
rect 1840 410 1970 440
rect 1800 390 1970 410
rect 2000 510 2170 530
rect 2000 480 2010 510
rect 2040 480 2170 510
rect 2000 440 2170 480
rect 2000 410 2010 440
rect 2040 410 2170 440
rect 2000 390 2170 410
rect 2200 510 2370 530
rect 2200 480 2210 510
rect 2240 480 2370 510
rect 2200 440 2370 480
rect 2200 410 2210 440
rect 2240 410 2370 440
rect 2200 390 2370 410
rect 2400 510 2570 530
rect 2400 480 2410 510
rect 2440 480 2570 510
rect 2400 440 2570 480
rect 2400 410 2410 440
rect 2440 410 2570 440
rect 2400 390 2570 410
rect 2600 510 2770 530
rect 2600 480 2610 510
rect 2640 480 2770 510
rect 2600 440 2770 480
rect 2600 410 2610 440
rect 2640 410 2770 440
rect 2600 390 2770 410
rect 2800 510 2970 530
rect 2800 480 2810 510
rect 2840 480 2970 510
rect 2800 440 2970 480
rect 2800 410 2810 440
rect 2840 410 2970 440
rect 2800 390 2970 410
rect 3000 510 3170 530
rect 3000 480 3010 510
rect 3040 480 3170 510
rect 3000 440 3170 480
rect 3000 410 3010 440
rect 3040 410 3170 440
rect 3000 390 3170 410
rect 3200 510 3370 530
rect 3200 480 3210 510
rect 3240 480 3370 510
rect 3200 440 3370 480
rect 3200 410 3210 440
rect 3240 410 3370 440
rect 3200 390 3370 410
rect 3400 510 3570 530
rect 3400 480 3410 510
rect 3440 480 3570 510
rect 3400 440 3570 480
rect 3400 410 3410 440
rect 3440 410 3570 440
rect 3400 390 3570 410
rect 3600 510 3770 530
rect 3600 480 3610 510
rect 3640 480 3770 510
rect 3600 440 3770 480
rect 3600 410 3610 440
rect 3640 410 3770 440
rect 3600 390 3770 410
rect 3800 510 3970 530
rect 3800 480 3810 510
rect 3840 480 3970 510
rect 3800 440 3970 480
rect 3800 410 3810 440
rect 3840 410 3970 440
rect 3800 390 3970 410
rect 4000 510 4170 530
rect 4000 480 4010 510
rect 4040 480 4170 510
rect 4000 440 4170 480
rect 4000 410 4010 440
rect 4040 410 4170 440
rect 4000 390 4170 410
rect 4200 510 4370 530
rect 4200 480 4210 510
rect 4240 480 4370 510
rect 4200 440 4370 480
rect 4200 410 4210 440
rect 4240 410 4370 440
rect 4200 390 4370 410
rect 4400 510 4570 530
rect 4400 480 4410 510
rect 4440 480 4570 510
rect 4400 440 4570 480
rect 4400 410 4410 440
rect 4440 410 4570 440
rect 4400 390 4570 410
rect 4600 510 4770 530
rect 4600 480 4610 510
rect 4640 480 4770 510
rect 4600 440 4770 480
rect 4600 410 4610 440
rect 4640 410 4770 440
rect 4600 390 4770 410
rect 4800 510 4970 530
rect 4800 480 4810 510
rect 4840 480 4970 510
rect 4800 440 4970 480
rect 4800 410 4810 440
rect 4840 410 4970 440
rect 4800 390 4970 410
rect 5000 510 5170 530
rect 5000 480 5010 510
rect 5040 480 5170 510
rect 5000 440 5170 480
rect 5000 410 5010 440
rect 5040 410 5170 440
rect 5000 390 5170 410
rect 5200 510 5370 530
rect 5200 480 5210 510
rect 5240 480 5370 510
rect 5200 440 5370 480
rect 5200 410 5210 440
rect 5240 410 5370 440
rect 5200 390 5370 410
rect 5400 510 5570 530
rect 5400 480 5410 510
rect 5440 480 5570 510
rect 5400 440 5570 480
rect 5400 410 5410 440
rect 5440 410 5570 440
rect 5400 390 5570 410
rect 5600 510 5770 530
rect 5600 480 5610 510
rect 5640 480 5770 510
rect 5600 440 5770 480
rect 5600 410 5610 440
rect 5640 410 5770 440
rect 5600 390 5770 410
rect 5800 510 5970 530
rect 5800 480 5810 510
rect 5840 480 5970 510
rect 5800 440 5970 480
rect 5800 410 5810 440
rect 5840 410 5970 440
rect 5800 390 5970 410
rect 6000 510 6170 530
rect 6000 480 6010 510
rect 6040 480 6170 510
rect 6000 440 6170 480
rect 6000 410 6010 440
rect 6040 410 6170 440
rect 6000 390 6170 410
rect 6200 510 6370 530
rect 6200 480 6210 510
rect 6240 480 6370 510
rect 6200 440 6370 480
rect 6200 410 6210 440
rect 6240 410 6370 440
rect 6200 390 6370 410
rect 6400 510 6570 530
rect 6400 480 6410 510
rect 6440 480 6570 510
rect 6400 440 6570 480
rect 6400 410 6410 440
rect 6440 410 6570 440
rect 6400 390 6570 410
rect -200 325 -30 345
rect -200 295 -190 325
rect -160 295 -30 325
rect -200 255 -30 295
rect -200 225 -190 255
rect -160 225 -30 255
rect -200 205 -30 225
rect 0 325 170 345
rect 0 295 10 325
rect 40 295 170 325
rect 0 255 170 295
rect 0 225 10 255
rect 40 225 170 255
rect 0 205 170 225
rect 200 325 370 345
rect 200 295 210 325
rect 240 295 370 325
rect 200 255 370 295
rect 200 225 210 255
rect 240 225 370 255
rect 200 205 370 225
rect 400 325 570 345
rect 400 295 410 325
rect 440 295 570 325
rect 400 255 570 295
rect 400 225 410 255
rect 440 225 570 255
rect 400 205 570 225
rect 600 325 770 345
rect 600 295 610 325
rect 640 295 770 325
rect 600 255 770 295
rect 600 225 610 255
rect 640 225 770 255
rect 600 205 770 225
rect 800 325 970 345
rect 800 295 810 325
rect 840 295 970 325
rect 800 255 970 295
rect 800 225 810 255
rect 840 225 970 255
rect 800 205 970 225
rect 1000 325 1170 345
rect 1000 295 1010 325
rect 1040 295 1170 325
rect 1000 255 1170 295
rect 1000 225 1010 255
rect 1040 225 1170 255
rect 1000 205 1170 225
rect 1200 325 1370 345
rect 1200 295 1210 325
rect 1240 295 1370 325
rect 1200 255 1370 295
rect 1200 225 1210 255
rect 1240 225 1370 255
rect 1200 205 1370 225
rect 1400 325 1570 345
rect 1400 295 1410 325
rect 1440 295 1570 325
rect 1400 255 1570 295
rect 1400 225 1410 255
rect 1440 225 1570 255
rect 1400 205 1570 225
rect 1600 325 1770 345
rect 1600 295 1610 325
rect 1640 295 1770 325
rect 1600 255 1770 295
rect 1600 225 1610 255
rect 1640 225 1770 255
rect 1600 205 1770 225
rect 1800 325 1970 345
rect 1800 295 1810 325
rect 1840 295 1970 325
rect 1800 255 1970 295
rect 1800 225 1810 255
rect 1840 225 1970 255
rect 1800 205 1970 225
rect 2000 325 2170 345
rect 2000 295 2010 325
rect 2040 295 2170 325
rect 2000 255 2170 295
rect 2000 225 2010 255
rect 2040 225 2170 255
rect 2000 205 2170 225
rect 2200 325 2370 345
rect 2200 295 2210 325
rect 2240 295 2370 325
rect 2200 255 2370 295
rect 2200 225 2210 255
rect 2240 225 2370 255
rect 2200 205 2370 225
rect 2400 325 2570 345
rect 2400 295 2410 325
rect 2440 295 2570 325
rect 2400 255 2570 295
rect 2400 225 2410 255
rect 2440 225 2570 255
rect 2400 205 2570 225
rect 2600 325 2770 345
rect 2600 295 2610 325
rect 2640 295 2770 325
rect 2600 255 2770 295
rect 2600 225 2610 255
rect 2640 225 2770 255
rect 2600 205 2770 225
rect 2800 325 2970 345
rect 2800 295 2810 325
rect 2840 295 2970 325
rect 2800 255 2970 295
rect 2800 225 2810 255
rect 2840 225 2970 255
rect 2800 205 2970 225
rect 3000 325 3170 345
rect 3000 295 3010 325
rect 3040 295 3170 325
rect 3000 255 3170 295
rect 3000 225 3010 255
rect 3040 225 3170 255
rect 3000 205 3170 225
rect 3200 325 3370 345
rect 3200 295 3210 325
rect 3240 295 3370 325
rect 3200 255 3370 295
rect 3200 225 3210 255
rect 3240 225 3370 255
rect 3200 205 3370 225
rect 3400 325 3570 345
rect 3400 295 3410 325
rect 3440 295 3570 325
rect 3400 255 3570 295
rect 3400 225 3410 255
rect 3440 225 3570 255
rect 3400 205 3570 225
rect 3600 325 3770 345
rect 3600 295 3610 325
rect 3640 295 3770 325
rect 3600 255 3770 295
rect 3600 225 3610 255
rect 3640 225 3770 255
rect 3600 205 3770 225
rect 3800 325 3970 345
rect 3800 295 3810 325
rect 3840 295 3970 325
rect 3800 255 3970 295
rect 3800 225 3810 255
rect 3840 225 3970 255
rect 3800 205 3970 225
rect 4000 325 4170 345
rect 4000 295 4010 325
rect 4040 295 4170 325
rect 4000 255 4170 295
rect 4000 225 4010 255
rect 4040 225 4170 255
rect 4000 205 4170 225
rect 4200 325 4370 345
rect 4200 295 4210 325
rect 4240 295 4370 325
rect 4200 255 4370 295
rect 4200 225 4210 255
rect 4240 225 4370 255
rect 4200 205 4370 225
rect 4400 325 4570 345
rect 4400 295 4410 325
rect 4440 295 4570 325
rect 4400 255 4570 295
rect 4400 225 4410 255
rect 4440 225 4570 255
rect 4400 205 4570 225
rect 4600 325 4770 345
rect 4600 295 4610 325
rect 4640 295 4770 325
rect 4600 255 4770 295
rect 4600 225 4610 255
rect 4640 225 4770 255
rect 4600 205 4770 225
rect 4800 325 4970 345
rect 4800 295 4810 325
rect 4840 295 4970 325
rect 4800 255 4970 295
rect 4800 225 4810 255
rect 4840 225 4970 255
rect 4800 205 4970 225
rect 5000 325 5170 345
rect 5000 295 5010 325
rect 5040 295 5170 325
rect 5000 255 5170 295
rect 5000 225 5010 255
rect 5040 225 5170 255
rect 5000 205 5170 225
rect 5200 325 5370 345
rect 5200 295 5210 325
rect 5240 295 5370 325
rect 5200 255 5370 295
rect 5200 225 5210 255
rect 5240 225 5370 255
rect 5200 205 5370 225
rect 5400 325 5570 345
rect 5400 295 5410 325
rect 5440 295 5570 325
rect 5400 255 5570 295
rect 5400 225 5410 255
rect 5440 225 5570 255
rect 5400 205 5570 225
rect 5600 325 5770 345
rect 5600 295 5610 325
rect 5640 295 5770 325
rect 5600 255 5770 295
rect 5600 225 5610 255
rect 5640 225 5770 255
rect 5600 205 5770 225
rect 5800 325 5970 345
rect 5800 295 5810 325
rect 5840 295 5970 325
rect 5800 255 5970 295
rect 5800 225 5810 255
rect 5840 225 5970 255
rect 5800 205 5970 225
rect 6000 325 6170 345
rect 6000 295 6010 325
rect 6040 295 6170 325
rect 6000 255 6170 295
rect 6000 225 6010 255
rect 6040 225 6170 255
rect 6000 205 6170 225
rect 6200 325 6370 345
rect 6200 295 6210 325
rect 6240 295 6370 325
rect 6200 255 6370 295
rect 6200 225 6210 255
rect 6240 225 6370 255
rect 6200 205 6370 225
rect 6400 325 6570 345
rect 6400 295 6410 325
rect 6440 295 6570 325
rect 6400 255 6570 295
rect 6400 225 6410 255
rect 6440 225 6570 255
rect 6400 205 6570 225
rect -200 140 -30 160
rect -200 110 -190 140
rect -160 110 -30 140
rect -200 70 -30 110
rect -200 40 -190 70
rect -160 40 -30 70
rect -200 20 -30 40
rect 0 140 170 160
rect 0 110 10 140
rect 40 110 170 140
rect 0 70 170 110
rect 0 40 10 70
rect 40 40 170 70
rect 0 20 170 40
rect 200 140 370 160
rect 200 110 210 140
rect 240 110 370 140
rect 200 70 370 110
rect 200 40 210 70
rect 240 40 370 70
rect 200 20 370 40
rect 400 140 570 160
rect 400 110 410 140
rect 440 110 570 140
rect 400 70 570 110
rect 400 40 410 70
rect 440 40 570 70
rect 400 20 570 40
rect 600 140 770 160
rect 600 110 610 140
rect 640 110 770 140
rect 600 70 770 110
rect 600 40 610 70
rect 640 40 770 70
rect 600 20 770 40
rect 800 140 970 160
rect 800 110 810 140
rect 840 110 970 140
rect 800 70 970 110
rect 800 40 810 70
rect 840 40 970 70
rect 800 20 970 40
rect 1000 140 1170 160
rect 1000 110 1010 140
rect 1040 110 1170 140
rect 1000 70 1170 110
rect 1000 40 1010 70
rect 1040 40 1170 70
rect 1000 20 1170 40
rect 1200 140 1370 160
rect 1200 110 1210 140
rect 1240 110 1370 140
rect 1200 70 1370 110
rect 1200 40 1210 70
rect 1240 40 1370 70
rect 1200 20 1370 40
rect 1400 140 1570 160
rect 1400 110 1410 140
rect 1440 110 1570 140
rect 1400 70 1570 110
rect 1400 40 1410 70
rect 1440 40 1570 70
rect 1400 20 1570 40
rect 1600 140 1770 160
rect 1600 110 1610 140
rect 1640 110 1770 140
rect 1600 70 1770 110
rect 1600 40 1610 70
rect 1640 40 1770 70
rect 1600 20 1770 40
rect 1800 140 1970 160
rect 1800 110 1810 140
rect 1840 110 1970 140
rect 1800 70 1970 110
rect 1800 40 1810 70
rect 1840 40 1970 70
rect 1800 20 1970 40
rect 2000 140 2170 160
rect 2000 110 2010 140
rect 2040 110 2170 140
rect 2000 70 2170 110
rect 2000 40 2010 70
rect 2040 40 2170 70
rect 2000 20 2170 40
rect 2200 140 2370 160
rect 2200 110 2210 140
rect 2240 110 2370 140
rect 2200 70 2370 110
rect 2200 40 2210 70
rect 2240 40 2370 70
rect 2200 20 2370 40
rect 2400 140 2570 160
rect 2400 110 2410 140
rect 2440 110 2570 140
rect 2400 70 2570 110
rect 2400 40 2410 70
rect 2440 40 2570 70
rect 2400 20 2570 40
rect 2600 140 2770 160
rect 2600 110 2610 140
rect 2640 110 2770 140
rect 2600 70 2770 110
rect 2600 40 2610 70
rect 2640 40 2770 70
rect 2600 20 2770 40
rect 2800 140 2970 160
rect 2800 110 2810 140
rect 2840 110 2970 140
rect 2800 70 2970 110
rect 2800 40 2810 70
rect 2840 40 2970 70
rect 2800 20 2970 40
rect 3000 140 3170 160
rect 3000 110 3010 140
rect 3040 110 3170 140
rect 3000 70 3170 110
rect 3000 40 3010 70
rect 3040 40 3170 70
rect 3000 20 3170 40
rect 3200 140 3370 160
rect 3200 110 3210 140
rect 3240 110 3370 140
rect 3200 70 3370 110
rect 3200 40 3210 70
rect 3240 40 3370 70
rect 3200 20 3370 40
rect 3400 140 3570 160
rect 3400 110 3410 140
rect 3440 110 3570 140
rect 3400 70 3570 110
rect 3400 40 3410 70
rect 3440 40 3570 70
rect 3400 20 3570 40
rect 3600 140 3770 160
rect 3600 110 3610 140
rect 3640 110 3770 140
rect 3600 70 3770 110
rect 3600 40 3610 70
rect 3640 40 3770 70
rect 3600 20 3770 40
rect 3800 140 3970 160
rect 3800 110 3810 140
rect 3840 110 3970 140
rect 3800 70 3970 110
rect 3800 40 3810 70
rect 3840 40 3970 70
rect 3800 20 3970 40
rect 4000 140 4170 160
rect 4000 110 4010 140
rect 4040 110 4170 140
rect 4000 70 4170 110
rect 4000 40 4010 70
rect 4040 40 4170 70
rect 4000 20 4170 40
rect 4200 140 4370 160
rect 4200 110 4210 140
rect 4240 110 4370 140
rect 4200 70 4370 110
rect 4200 40 4210 70
rect 4240 40 4370 70
rect 4200 20 4370 40
rect 4400 140 4570 160
rect 4400 110 4410 140
rect 4440 110 4570 140
rect 4400 70 4570 110
rect 4400 40 4410 70
rect 4440 40 4570 70
rect 4400 20 4570 40
rect 4600 140 4770 160
rect 4600 110 4610 140
rect 4640 110 4770 140
rect 4600 70 4770 110
rect 4600 40 4610 70
rect 4640 40 4770 70
rect 4600 20 4770 40
rect 4800 140 4970 160
rect 4800 110 4810 140
rect 4840 110 4970 140
rect 4800 70 4970 110
rect 4800 40 4810 70
rect 4840 40 4970 70
rect 4800 20 4970 40
rect 5000 140 5170 160
rect 5000 110 5010 140
rect 5040 110 5170 140
rect 5000 70 5170 110
rect 5000 40 5010 70
rect 5040 40 5170 70
rect 5000 20 5170 40
rect 5200 140 5370 160
rect 5200 110 5210 140
rect 5240 110 5370 140
rect 5200 70 5370 110
rect 5200 40 5210 70
rect 5240 40 5370 70
rect 5200 20 5370 40
rect 5400 140 5570 160
rect 5400 110 5410 140
rect 5440 110 5570 140
rect 5400 70 5570 110
rect 5400 40 5410 70
rect 5440 40 5570 70
rect 5400 20 5570 40
rect 5600 140 5770 160
rect 5600 110 5610 140
rect 5640 110 5770 140
rect 5600 70 5770 110
rect 5600 40 5610 70
rect 5640 40 5770 70
rect 5600 20 5770 40
rect 5800 140 5970 160
rect 5800 110 5810 140
rect 5840 110 5970 140
rect 5800 70 5970 110
rect 5800 40 5810 70
rect 5840 40 5970 70
rect 5800 20 5970 40
rect 6000 140 6170 160
rect 6000 110 6010 140
rect 6040 110 6170 140
rect 6000 70 6170 110
rect 6000 40 6010 70
rect 6040 40 6170 70
rect 6000 20 6170 40
rect 6200 140 6370 160
rect 6200 110 6210 140
rect 6240 110 6370 140
rect 6200 70 6370 110
rect 6200 40 6210 70
rect 6240 40 6370 70
rect 6200 20 6370 40
rect 6400 140 6570 160
rect 6400 110 6410 140
rect 6440 110 6570 140
rect 6400 70 6570 110
rect 6400 40 6410 70
rect 6440 40 6570 70
rect 6400 20 6570 40
rect -200 -45 -30 -25
rect -200 -75 -190 -45
rect -160 -75 -30 -45
rect -200 -115 -30 -75
rect -200 -145 -190 -115
rect -160 -145 -30 -115
rect -200 -165 -30 -145
rect 0 -45 170 -25
rect 0 -75 10 -45
rect 40 -75 170 -45
rect 0 -115 170 -75
rect 0 -145 10 -115
rect 40 -145 170 -115
rect 0 -165 170 -145
rect 200 -45 370 -25
rect 200 -75 210 -45
rect 240 -75 370 -45
rect 200 -115 370 -75
rect 200 -145 210 -115
rect 240 -145 370 -115
rect 200 -165 370 -145
rect 400 -45 570 -25
rect 400 -75 410 -45
rect 440 -75 570 -45
rect 400 -115 570 -75
rect 400 -145 410 -115
rect 440 -145 570 -115
rect 400 -165 570 -145
rect 600 -45 770 -25
rect 600 -75 610 -45
rect 640 -75 770 -45
rect 600 -115 770 -75
rect 600 -145 610 -115
rect 640 -145 770 -115
rect 600 -165 770 -145
rect 800 -45 970 -25
rect 800 -75 810 -45
rect 840 -75 970 -45
rect 800 -115 970 -75
rect 800 -145 810 -115
rect 840 -145 970 -115
rect 800 -165 970 -145
rect 1000 -45 1170 -25
rect 1000 -75 1010 -45
rect 1040 -75 1170 -45
rect 1000 -115 1170 -75
rect 1000 -145 1010 -115
rect 1040 -145 1170 -115
rect 1000 -165 1170 -145
rect 1200 -45 1370 -25
rect 1200 -75 1210 -45
rect 1240 -75 1370 -45
rect 1200 -115 1370 -75
rect 1200 -145 1210 -115
rect 1240 -145 1370 -115
rect 1200 -165 1370 -145
rect 1400 -45 1570 -25
rect 1400 -75 1410 -45
rect 1440 -75 1570 -45
rect 1400 -115 1570 -75
rect 1400 -145 1410 -115
rect 1440 -145 1570 -115
rect 1400 -165 1570 -145
rect 1600 -45 1770 -25
rect 1600 -75 1610 -45
rect 1640 -75 1770 -45
rect 1600 -115 1770 -75
rect 1600 -145 1610 -115
rect 1640 -145 1770 -115
rect 1600 -165 1770 -145
rect 1800 -45 1970 -25
rect 1800 -75 1810 -45
rect 1840 -75 1970 -45
rect 1800 -115 1970 -75
rect 1800 -145 1810 -115
rect 1840 -145 1970 -115
rect 1800 -165 1970 -145
rect 2000 -45 2170 -25
rect 2000 -75 2010 -45
rect 2040 -75 2170 -45
rect 2000 -115 2170 -75
rect 2000 -145 2010 -115
rect 2040 -145 2170 -115
rect 2000 -165 2170 -145
rect 2200 -45 2370 -25
rect 2200 -75 2210 -45
rect 2240 -75 2370 -45
rect 2200 -115 2370 -75
rect 2200 -145 2210 -115
rect 2240 -145 2370 -115
rect 2200 -165 2370 -145
rect 2400 -45 2570 -25
rect 2400 -75 2410 -45
rect 2440 -75 2570 -45
rect 2400 -115 2570 -75
rect 2400 -145 2410 -115
rect 2440 -145 2570 -115
rect 2400 -165 2570 -145
rect 2600 -45 2770 -25
rect 2600 -75 2610 -45
rect 2640 -75 2770 -45
rect 2600 -115 2770 -75
rect 2600 -145 2610 -115
rect 2640 -145 2770 -115
rect 2600 -165 2770 -145
rect 2800 -45 2970 -25
rect 2800 -75 2810 -45
rect 2840 -75 2970 -45
rect 2800 -115 2970 -75
rect 2800 -145 2810 -115
rect 2840 -145 2970 -115
rect 2800 -165 2970 -145
rect 3000 -45 3170 -25
rect 3000 -75 3010 -45
rect 3040 -75 3170 -45
rect 3000 -115 3170 -75
rect 3000 -145 3010 -115
rect 3040 -145 3170 -115
rect 3000 -165 3170 -145
rect 3200 -45 3370 -25
rect 3200 -75 3210 -45
rect 3240 -75 3370 -45
rect 3200 -115 3370 -75
rect 3200 -145 3210 -115
rect 3240 -145 3370 -115
rect 3200 -165 3370 -145
rect 3400 -45 3570 -25
rect 3400 -75 3410 -45
rect 3440 -75 3570 -45
rect 3400 -115 3570 -75
rect 3400 -145 3410 -115
rect 3440 -145 3570 -115
rect 3400 -165 3570 -145
rect 3600 -45 3770 -25
rect 3600 -75 3610 -45
rect 3640 -75 3770 -45
rect 3600 -115 3770 -75
rect 3600 -145 3610 -115
rect 3640 -145 3770 -115
rect 3600 -165 3770 -145
rect 3800 -45 3970 -25
rect 3800 -75 3810 -45
rect 3840 -75 3970 -45
rect 3800 -115 3970 -75
rect 3800 -145 3810 -115
rect 3840 -145 3970 -115
rect 3800 -165 3970 -145
rect 4000 -45 4170 -25
rect 4000 -75 4010 -45
rect 4040 -75 4170 -45
rect 4000 -115 4170 -75
rect 4000 -145 4010 -115
rect 4040 -145 4170 -115
rect 4000 -165 4170 -145
rect 4200 -45 4370 -25
rect 4200 -75 4210 -45
rect 4240 -75 4370 -45
rect 4200 -115 4370 -75
rect 4200 -145 4210 -115
rect 4240 -145 4370 -115
rect 4200 -165 4370 -145
rect 4400 -45 4570 -25
rect 4400 -75 4410 -45
rect 4440 -75 4570 -45
rect 4400 -115 4570 -75
rect 4400 -145 4410 -115
rect 4440 -145 4570 -115
rect 4400 -165 4570 -145
rect 4600 -45 4770 -25
rect 4600 -75 4610 -45
rect 4640 -75 4770 -45
rect 4600 -115 4770 -75
rect 4600 -145 4610 -115
rect 4640 -145 4770 -115
rect 4600 -165 4770 -145
rect 4800 -45 4970 -25
rect 4800 -75 4810 -45
rect 4840 -75 4970 -45
rect 4800 -115 4970 -75
rect 4800 -145 4810 -115
rect 4840 -145 4970 -115
rect 4800 -165 4970 -145
rect 5000 -45 5170 -25
rect 5000 -75 5010 -45
rect 5040 -75 5170 -45
rect 5000 -115 5170 -75
rect 5000 -145 5010 -115
rect 5040 -145 5170 -115
rect 5000 -165 5170 -145
rect 5200 -45 5370 -25
rect 5200 -75 5210 -45
rect 5240 -75 5370 -45
rect 5200 -115 5370 -75
rect 5200 -145 5210 -115
rect 5240 -145 5370 -115
rect 5200 -165 5370 -145
rect 5400 -45 5570 -25
rect 5400 -75 5410 -45
rect 5440 -75 5570 -45
rect 5400 -115 5570 -75
rect 5400 -145 5410 -115
rect 5440 -145 5570 -115
rect 5400 -165 5570 -145
rect 5600 -45 5770 -25
rect 5600 -75 5610 -45
rect 5640 -75 5770 -45
rect 5600 -115 5770 -75
rect 5600 -145 5610 -115
rect 5640 -145 5770 -115
rect 5600 -165 5770 -145
rect 5800 -45 5970 -25
rect 5800 -75 5810 -45
rect 5840 -75 5970 -45
rect 5800 -115 5970 -75
rect 5800 -145 5810 -115
rect 5840 -145 5970 -115
rect 5800 -165 5970 -145
rect 6000 -45 6170 -25
rect 6000 -75 6010 -45
rect 6040 -75 6170 -45
rect 6000 -115 6170 -75
rect 6000 -145 6010 -115
rect 6040 -145 6170 -115
rect 6000 -165 6170 -145
rect 6200 -45 6370 -25
rect 6200 -75 6210 -45
rect 6240 -75 6370 -45
rect 6200 -115 6370 -75
rect 6200 -145 6210 -115
rect 6240 -145 6370 -115
rect 6200 -165 6370 -145
rect 6400 -45 6570 -25
rect 6400 -75 6410 -45
rect 6440 -75 6570 -45
rect 6400 -115 6570 -75
rect 6400 -145 6410 -115
rect 6440 -145 6570 -115
rect 6400 -165 6570 -145
<< via3 >>
rect -145 12090 -105 12095
rect -145 12060 -140 12090
rect -140 12060 -110 12090
rect -110 12060 -105 12090
rect -145 12055 -105 12060
rect -95 12090 -55 12095
rect -95 12060 -90 12090
rect -90 12060 -60 12090
rect -60 12060 -55 12090
rect -95 12055 -55 12060
rect 6455 12065 6495 12070
rect 6455 12035 6460 12065
rect 6460 12035 6490 12065
rect 6490 12035 6495 12065
rect 6455 12030 6495 12035
rect 6505 12065 6545 12070
rect 6505 12035 6510 12065
rect 6510 12035 6540 12065
rect 6540 12035 6545 12065
rect 6505 12030 6545 12035
<< mimcap >>
rect -150 11970 -50 11980
rect -150 11890 -140 11970
rect -60 11890 -50 11970
rect -150 11880 -50 11890
rect 50 11970 150 11980
rect 50 11890 60 11970
rect 140 11890 150 11970
rect 50 11880 150 11890
rect 250 11970 350 11980
rect 250 11890 260 11970
rect 340 11890 350 11970
rect 250 11880 350 11890
rect 450 11970 550 11980
rect 450 11890 460 11970
rect 540 11890 550 11970
rect 450 11880 550 11890
rect 650 11970 750 11980
rect 650 11890 660 11970
rect 740 11890 750 11970
rect 650 11880 750 11890
rect 850 11970 950 11980
rect 850 11890 860 11970
rect 940 11890 950 11970
rect 850 11880 950 11890
rect 1050 11970 1150 11980
rect 1050 11890 1060 11970
rect 1140 11890 1150 11970
rect 1050 11880 1150 11890
rect 1250 11970 1350 11980
rect 1250 11890 1260 11970
rect 1340 11890 1350 11970
rect 1250 11880 1350 11890
rect 1450 11970 1550 11980
rect 1450 11890 1460 11970
rect 1540 11890 1550 11970
rect 1450 11880 1550 11890
rect 1650 11970 1750 11980
rect 1650 11890 1660 11970
rect 1740 11890 1750 11970
rect 1650 11880 1750 11890
rect 1850 11970 1950 11980
rect 1850 11890 1860 11970
rect 1940 11890 1950 11970
rect 1850 11880 1950 11890
rect 2050 11970 2150 11980
rect 2050 11890 2060 11970
rect 2140 11890 2150 11970
rect 2050 11880 2150 11890
rect 2250 11970 2350 11980
rect 2250 11890 2260 11970
rect 2340 11890 2350 11970
rect 2250 11880 2350 11890
rect 2450 11970 2550 11980
rect 2450 11890 2460 11970
rect 2540 11890 2550 11970
rect 2450 11880 2550 11890
rect 2650 11970 2750 11980
rect 2650 11890 2660 11970
rect 2740 11890 2750 11970
rect 2650 11880 2750 11890
rect 2850 11970 2950 11980
rect 2850 11890 2860 11970
rect 2940 11890 2950 11970
rect 2850 11880 2950 11890
rect 3050 11970 3150 11980
rect 3050 11890 3060 11970
rect 3140 11890 3150 11970
rect 3050 11880 3150 11890
rect 3250 11970 3350 11980
rect 3250 11890 3260 11970
rect 3340 11890 3350 11970
rect 3250 11880 3350 11890
rect 3450 11970 3550 11980
rect 3450 11890 3460 11970
rect 3540 11890 3550 11970
rect 3450 11880 3550 11890
rect 3650 11970 3750 11980
rect 3650 11890 3660 11970
rect 3740 11890 3750 11970
rect 3650 11880 3750 11890
rect 3850 11970 3950 11980
rect 3850 11890 3860 11970
rect 3940 11890 3950 11970
rect 3850 11880 3950 11890
rect 4050 11970 4150 11980
rect 4050 11890 4060 11970
rect 4140 11890 4150 11970
rect 4050 11880 4150 11890
rect 4250 11970 4350 11980
rect 4250 11890 4260 11970
rect 4340 11890 4350 11970
rect 4250 11880 4350 11890
rect 4450 11970 4550 11980
rect 4450 11890 4460 11970
rect 4540 11890 4550 11970
rect 4450 11880 4550 11890
rect 4650 11970 4750 11980
rect 4650 11890 4660 11970
rect 4740 11890 4750 11970
rect 4650 11880 4750 11890
rect 4850 11970 4950 11980
rect 4850 11890 4860 11970
rect 4940 11890 4950 11970
rect 4850 11880 4950 11890
rect 5050 11970 5150 11980
rect 5050 11890 5060 11970
rect 5140 11890 5150 11970
rect 5050 11880 5150 11890
rect 5250 11970 5350 11980
rect 5250 11890 5260 11970
rect 5340 11890 5350 11970
rect 5250 11880 5350 11890
rect 5450 11970 5550 11980
rect 5450 11890 5460 11970
rect 5540 11890 5550 11970
rect 5450 11880 5550 11890
rect 5650 11970 5750 11980
rect 5650 11890 5660 11970
rect 5740 11890 5750 11970
rect 5650 11880 5750 11890
rect 5850 11970 5950 11980
rect 5850 11890 5860 11970
rect 5940 11890 5950 11970
rect 5850 11880 5950 11890
rect 6050 11970 6150 11980
rect 6050 11890 6060 11970
rect 6140 11890 6150 11970
rect 6050 11880 6150 11890
rect 6250 11970 6350 11980
rect 6250 11890 6260 11970
rect 6340 11890 6350 11970
rect 6250 11880 6350 11890
rect 6450 11970 6550 11980
rect 6450 11890 6460 11970
rect 6540 11890 6550 11970
rect 6450 11880 6550 11890
rect -150 11785 -50 11795
rect -150 11705 -140 11785
rect -60 11705 -50 11785
rect -150 11695 -50 11705
rect 50 11785 150 11795
rect 50 11705 60 11785
rect 140 11705 150 11785
rect 50 11695 150 11705
rect 250 11785 350 11795
rect 250 11705 260 11785
rect 340 11705 350 11785
rect 250 11695 350 11705
rect 450 11785 550 11795
rect 450 11705 460 11785
rect 540 11705 550 11785
rect 450 11695 550 11705
rect 650 11785 750 11795
rect 650 11705 660 11785
rect 740 11705 750 11785
rect 650 11695 750 11705
rect 850 11785 950 11795
rect 850 11705 860 11785
rect 940 11705 950 11785
rect 850 11695 950 11705
rect 1050 11785 1150 11795
rect 1050 11705 1060 11785
rect 1140 11705 1150 11785
rect 1050 11695 1150 11705
rect 1250 11785 1350 11795
rect 1250 11705 1260 11785
rect 1340 11705 1350 11785
rect 1250 11695 1350 11705
rect 1450 11785 1550 11795
rect 1450 11705 1460 11785
rect 1540 11705 1550 11785
rect 1450 11695 1550 11705
rect 1650 11785 1750 11795
rect 1650 11705 1660 11785
rect 1740 11705 1750 11785
rect 1650 11695 1750 11705
rect 1850 11785 1950 11795
rect 1850 11705 1860 11785
rect 1940 11705 1950 11785
rect 1850 11695 1950 11705
rect 2050 11785 2150 11795
rect 2050 11705 2060 11785
rect 2140 11705 2150 11785
rect 2050 11695 2150 11705
rect 2250 11785 2350 11795
rect 2250 11705 2260 11785
rect 2340 11705 2350 11785
rect 2250 11695 2350 11705
rect 2450 11785 2550 11795
rect 2450 11705 2460 11785
rect 2540 11705 2550 11785
rect 2450 11695 2550 11705
rect 2650 11785 2750 11795
rect 2650 11705 2660 11785
rect 2740 11705 2750 11785
rect 2650 11695 2750 11705
rect 2850 11785 2950 11795
rect 2850 11705 2860 11785
rect 2940 11705 2950 11785
rect 2850 11695 2950 11705
rect 3050 11785 3150 11795
rect 3050 11705 3060 11785
rect 3140 11705 3150 11785
rect 3050 11695 3150 11705
rect 3250 11785 3350 11795
rect 3250 11705 3260 11785
rect 3340 11705 3350 11785
rect 3250 11695 3350 11705
rect 3450 11785 3550 11795
rect 3450 11705 3460 11785
rect 3540 11705 3550 11785
rect 3450 11695 3550 11705
rect 3650 11785 3750 11795
rect 3650 11705 3660 11785
rect 3740 11705 3750 11785
rect 3650 11695 3750 11705
rect 3850 11785 3950 11795
rect 3850 11705 3860 11785
rect 3940 11705 3950 11785
rect 3850 11695 3950 11705
rect 4050 11785 4150 11795
rect 4050 11705 4060 11785
rect 4140 11705 4150 11785
rect 4050 11695 4150 11705
rect 4250 11785 4350 11795
rect 4250 11705 4260 11785
rect 4340 11705 4350 11785
rect 4250 11695 4350 11705
rect 4450 11785 4550 11795
rect 4450 11705 4460 11785
rect 4540 11705 4550 11785
rect 4450 11695 4550 11705
rect 4650 11785 4750 11795
rect 4650 11705 4660 11785
rect 4740 11705 4750 11785
rect 4650 11695 4750 11705
rect 4850 11785 4950 11795
rect 4850 11705 4860 11785
rect 4940 11705 4950 11785
rect 4850 11695 4950 11705
rect 5050 11785 5150 11795
rect 5050 11705 5060 11785
rect 5140 11705 5150 11785
rect 5050 11695 5150 11705
rect 5250 11785 5350 11795
rect 5250 11705 5260 11785
rect 5340 11705 5350 11785
rect 5250 11695 5350 11705
rect 5450 11785 5550 11795
rect 5450 11705 5460 11785
rect 5540 11705 5550 11785
rect 5450 11695 5550 11705
rect 5650 11785 5750 11795
rect 5650 11705 5660 11785
rect 5740 11705 5750 11785
rect 5650 11695 5750 11705
rect 5850 11785 5950 11795
rect 5850 11705 5860 11785
rect 5940 11705 5950 11785
rect 5850 11695 5950 11705
rect 6050 11785 6150 11795
rect 6050 11705 6060 11785
rect 6140 11705 6150 11785
rect 6050 11695 6150 11705
rect 6250 11785 6350 11795
rect 6250 11705 6260 11785
rect 6340 11705 6350 11785
rect 6250 11695 6350 11705
rect 6450 11785 6550 11795
rect 6450 11705 6460 11785
rect 6540 11705 6550 11785
rect 6450 11695 6550 11705
rect -150 11600 -50 11610
rect -150 11520 -140 11600
rect -60 11520 -50 11600
rect -150 11510 -50 11520
rect 50 11600 150 11610
rect 50 11520 60 11600
rect 140 11520 150 11600
rect 50 11510 150 11520
rect 250 11600 350 11610
rect 250 11520 260 11600
rect 340 11520 350 11600
rect 250 11510 350 11520
rect 450 11600 550 11610
rect 450 11520 460 11600
rect 540 11520 550 11600
rect 450 11510 550 11520
rect 650 11600 750 11610
rect 650 11520 660 11600
rect 740 11520 750 11600
rect 650 11510 750 11520
rect 850 11600 950 11610
rect 850 11520 860 11600
rect 940 11520 950 11600
rect 850 11510 950 11520
rect 1050 11600 1150 11610
rect 1050 11520 1060 11600
rect 1140 11520 1150 11600
rect 1050 11510 1150 11520
rect 1250 11600 1350 11610
rect 1250 11520 1260 11600
rect 1340 11520 1350 11600
rect 1250 11510 1350 11520
rect 1450 11600 1550 11610
rect 1450 11520 1460 11600
rect 1540 11520 1550 11600
rect 1450 11510 1550 11520
rect 1650 11600 1750 11610
rect 1650 11520 1660 11600
rect 1740 11520 1750 11600
rect 1650 11510 1750 11520
rect 1850 11600 1950 11610
rect 1850 11520 1860 11600
rect 1940 11520 1950 11600
rect 1850 11510 1950 11520
rect 2050 11600 2150 11610
rect 2050 11520 2060 11600
rect 2140 11520 2150 11600
rect 2050 11510 2150 11520
rect 2250 11600 2350 11610
rect 2250 11520 2260 11600
rect 2340 11520 2350 11600
rect 2250 11510 2350 11520
rect 2450 11600 2550 11610
rect 2450 11520 2460 11600
rect 2540 11520 2550 11600
rect 2450 11510 2550 11520
rect 2650 11600 2750 11610
rect 2650 11520 2660 11600
rect 2740 11520 2750 11600
rect 2650 11510 2750 11520
rect 2850 11600 2950 11610
rect 2850 11520 2860 11600
rect 2940 11520 2950 11600
rect 2850 11510 2950 11520
rect 3050 11600 3150 11610
rect 3050 11520 3060 11600
rect 3140 11520 3150 11600
rect 3050 11510 3150 11520
rect 3250 11600 3350 11610
rect 3250 11520 3260 11600
rect 3340 11520 3350 11600
rect 3250 11510 3350 11520
rect 3450 11600 3550 11610
rect 3450 11520 3460 11600
rect 3540 11520 3550 11600
rect 3450 11510 3550 11520
rect 3650 11600 3750 11610
rect 3650 11520 3660 11600
rect 3740 11520 3750 11600
rect 3650 11510 3750 11520
rect 3850 11600 3950 11610
rect 3850 11520 3860 11600
rect 3940 11520 3950 11600
rect 3850 11510 3950 11520
rect 4050 11600 4150 11610
rect 4050 11520 4060 11600
rect 4140 11520 4150 11600
rect 4050 11510 4150 11520
rect 4250 11600 4350 11610
rect 4250 11520 4260 11600
rect 4340 11520 4350 11600
rect 4250 11510 4350 11520
rect 4450 11600 4550 11610
rect 4450 11520 4460 11600
rect 4540 11520 4550 11600
rect 4450 11510 4550 11520
rect 4650 11600 4750 11610
rect 4650 11520 4660 11600
rect 4740 11520 4750 11600
rect 4650 11510 4750 11520
rect 4850 11600 4950 11610
rect 4850 11520 4860 11600
rect 4940 11520 4950 11600
rect 4850 11510 4950 11520
rect 5050 11600 5150 11610
rect 5050 11520 5060 11600
rect 5140 11520 5150 11600
rect 5050 11510 5150 11520
rect 5250 11600 5350 11610
rect 5250 11520 5260 11600
rect 5340 11520 5350 11600
rect 5250 11510 5350 11520
rect 5450 11600 5550 11610
rect 5450 11520 5460 11600
rect 5540 11520 5550 11600
rect 5450 11510 5550 11520
rect 5650 11600 5750 11610
rect 5650 11520 5660 11600
rect 5740 11520 5750 11600
rect 5650 11510 5750 11520
rect 5850 11600 5950 11610
rect 5850 11520 5860 11600
rect 5940 11520 5950 11600
rect 5850 11510 5950 11520
rect 6050 11600 6150 11610
rect 6050 11520 6060 11600
rect 6140 11520 6150 11600
rect 6050 11510 6150 11520
rect 6250 11600 6350 11610
rect 6250 11520 6260 11600
rect 6340 11520 6350 11600
rect 6250 11510 6350 11520
rect 6450 11600 6550 11610
rect 6450 11520 6460 11600
rect 6540 11520 6550 11600
rect 6450 11510 6550 11520
rect -150 11415 -50 11425
rect -150 11335 -140 11415
rect -60 11335 -50 11415
rect -150 11325 -50 11335
rect 50 11415 150 11425
rect 50 11335 60 11415
rect 140 11335 150 11415
rect 50 11325 150 11335
rect 250 11415 350 11425
rect 250 11335 260 11415
rect 340 11335 350 11415
rect 250 11325 350 11335
rect 450 11415 550 11425
rect 450 11335 460 11415
rect 540 11335 550 11415
rect 450 11325 550 11335
rect 650 11415 750 11425
rect 650 11335 660 11415
rect 740 11335 750 11415
rect 650 11325 750 11335
rect 850 11415 950 11425
rect 850 11335 860 11415
rect 940 11335 950 11415
rect 850 11325 950 11335
rect 1050 11415 1150 11425
rect 1050 11335 1060 11415
rect 1140 11335 1150 11415
rect 1050 11325 1150 11335
rect 1250 11415 1350 11425
rect 1250 11335 1260 11415
rect 1340 11335 1350 11415
rect 1250 11325 1350 11335
rect 1450 11415 1550 11425
rect 1450 11335 1460 11415
rect 1540 11335 1550 11415
rect 1450 11325 1550 11335
rect 1650 11415 1750 11425
rect 1650 11335 1660 11415
rect 1740 11335 1750 11415
rect 1650 11325 1750 11335
rect 1850 11415 1950 11425
rect 1850 11335 1860 11415
rect 1940 11335 1950 11415
rect 1850 11325 1950 11335
rect 2050 11415 2150 11425
rect 2050 11335 2060 11415
rect 2140 11335 2150 11415
rect 2050 11325 2150 11335
rect 2250 11415 2350 11425
rect 2250 11335 2260 11415
rect 2340 11335 2350 11415
rect 2250 11325 2350 11335
rect 2450 11415 2550 11425
rect 2450 11335 2460 11415
rect 2540 11335 2550 11415
rect 2450 11325 2550 11335
rect 2650 11415 2750 11425
rect 2650 11335 2660 11415
rect 2740 11335 2750 11415
rect 2650 11325 2750 11335
rect 2850 11415 2950 11425
rect 2850 11335 2860 11415
rect 2940 11335 2950 11415
rect 2850 11325 2950 11335
rect 3050 11415 3150 11425
rect 3050 11335 3060 11415
rect 3140 11335 3150 11415
rect 3050 11325 3150 11335
rect 3250 11415 3350 11425
rect 3250 11335 3260 11415
rect 3340 11335 3350 11415
rect 3250 11325 3350 11335
rect 3450 11415 3550 11425
rect 3450 11335 3460 11415
rect 3540 11335 3550 11415
rect 3450 11325 3550 11335
rect 3650 11415 3750 11425
rect 3650 11335 3660 11415
rect 3740 11335 3750 11415
rect 3650 11325 3750 11335
rect 3850 11415 3950 11425
rect 3850 11335 3860 11415
rect 3940 11335 3950 11415
rect 3850 11325 3950 11335
rect 4050 11415 4150 11425
rect 4050 11335 4060 11415
rect 4140 11335 4150 11415
rect 4050 11325 4150 11335
rect 4250 11415 4350 11425
rect 4250 11335 4260 11415
rect 4340 11335 4350 11415
rect 4250 11325 4350 11335
rect 4450 11415 4550 11425
rect 4450 11335 4460 11415
rect 4540 11335 4550 11415
rect 4450 11325 4550 11335
rect 4650 11415 4750 11425
rect 4650 11335 4660 11415
rect 4740 11335 4750 11415
rect 4650 11325 4750 11335
rect 4850 11415 4950 11425
rect 4850 11335 4860 11415
rect 4940 11335 4950 11415
rect 4850 11325 4950 11335
rect 5050 11415 5150 11425
rect 5050 11335 5060 11415
rect 5140 11335 5150 11415
rect 5050 11325 5150 11335
rect 5250 11415 5350 11425
rect 5250 11335 5260 11415
rect 5340 11335 5350 11415
rect 5250 11325 5350 11335
rect 5450 11415 5550 11425
rect 5450 11335 5460 11415
rect 5540 11335 5550 11415
rect 5450 11325 5550 11335
rect 5650 11415 5750 11425
rect 5650 11335 5660 11415
rect 5740 11335 5750 11415
rect 5650 11325 5750 11335
rect 5850 11415 5950 11425
rect 5850 11335 5860 11415
rect 5940 11335 5950 11415
rect 5850 11325 5950 11335
rect 6050 11415 6150 11425
rect 6050 11335 6060 11415
rect 6140 11335 6150 11415
rect 6050 11325 6150 11335
rect 6250 11415 6350 11425
rect 6250 11335 6260 11415
rect 6340 11335 6350 11415
rect 6250 11325 6350 11335
rect 6450 11415 6550 11425
rect 6450 11335 6460 11415
rect 6540 11335 6550 11415
rect 6450 11325 6550 11335
rect -150 11230 -50 11240
rect -150 11150 -140 11230
rect -60 11150 -50 11230
rect -150 11140 -50 11150
rect 50 11230 150 11240
rect 50 11150 60 11230
rect 140 11150 150 11230
rect 50 11140 150 11150
rect 250 11230 350 11240
rect 250 11150 260 11230
rect 340 11150 350 11230
rect 250 11140 350 11150
rect 450 11230 550 11240
rect 450 11150 460 11230
rect 540 11150 550 11230
rect 450 11140 550 11150
rect 650 11230 750 11240
rect 650 11150 660 11230
rect 740 11150 750 11230
rect 650 11140 750 11150
rect 850 11230 950 11240
rect 850 11150 860 11230
rect 940 11150 950 11230
rect 850 11140 950 11150
rect 1050 11230 1150 11240
rect 1050 11150 1060 11230
rect 1140 11150 1150 11230
rect 1050 11140 1150 11150
rect 1250 11230 1350 11240
rect 1250 11150 1260 11230
rect 1340 11150 1350 11230
rect 1250 11140 1350 11150
rect 1450 11230 1550 11240
rect 1450 11150 1460 11230
rect 1540 11150 1550 11230
rect 1450 11140 1550 11150
rect 1650 11230 1750 11240
rect 1650 11150 1660 11230
rect 1740 11150 1750 11230
rect 1650 11140 1750 11150
rect 1850 11230 1950 11240
rect 1850 11150 1860 11230
rect 1940 11150 1950 11230
rect 1850 11140 1950 11150
rect 2050 11230 2150 11240
rect 2050 11150 2060 11230
rect 2140 11150 2150 11230
rect 2050 11140 2150 11150
rect 2250 11230 2350 11240
rect 2250 11150 2260 11230
rect 2340 11150 2350 11230
rect 2250 11140 2350 11150
rect 2450 11230 2550 11240
rect 2450 11150 2460 11230
rect 2540 11150 2550 11230
rect 2450 11140 2550 11150
rect 2650 11230 2750 11240
rect 2650 11150 2660 11230
rect 2740 11150 2750 11230
rect 2650 11140 2750 11150
rect 2850 11230 2950 11240
rect 2850 11150 2860 11230
rect 2940 11150 2950 11230
rect 2850 11140 2950 11150
rect 3050 11230 3150 11240
rect 3050 11150 3060 11230
rect 3140 11150 3150 11230
rect 3050 11140 3150 11150
rect 3250 11230 3350 11240
rect 3250 11150 3260 11230
rect 3340 11150 3350 11230
rect 3250 11140 3350 11150
rect 3450 11230 3550 11240
rect 3450 11150 3460 11230
rect 3540 11150 3550 11230
rect 3450 11140 3550 11150
rect 3650 11230 3750 11240
rect 3650 11150 3660 11230
rect 3740 11150 3750 11230
rect 3650 11140 3750 11150
rect 3850 11230 3950 11240
rect 3850 11150 3860 11230
rect 3940 11150 3950 11230
rect 3850 11140 3950 11150
rect 4050 11230 4150 11240
rect 4050 11150 4060 11230
rect 4140 11150 4150 11230
rect 4050 11140 4150 11150
rect 4250 11230 4350 11240
rect 4250 11150 4260 11230
rect 4340 11150 4350 11230
rect 4250 11140 4350 11150
rect 4450 11230 4550 11240
rect 4450 11150 4460 11230
rect 4540 11150 4550 11230
rect 4450 11140 4550 11150
rect 4650 11230 4750 11240
rect 4650 11150 4660 11230
rect 4740 11150 4750 11230
rect 4650 11140 4750 11150
rect 4850 11230 4950 11240
rect 4850 11150 4860 11230
rect 4940 11150 4950 11230
rect 4850 11140 4950 11150
rect 5050 11230 5150 11240
rect 5050 11150 5060 11230
rect 5140 11150 5150 11230
rect 5050 11140 5150 11150
rect 5250 11230 5350 11240
rect 5250 11150 5260 11230
rect 5340 11150 5350 11230
rect 5250 11140 5350 11150
rect 5450 11230 5550 11240
rect 5450 11150 5460 11230
rect 5540 11150 5550 11230
rect 5450 11140 5550 11150
rect 5650 11230 5750 11240
rect 5650 11150 5660 11230
rect 5740 11150 5750 11230
rect 5650 11140 5750 11150
rect 5850 11230 5950 11240
rect 5850 11150 5860 11230
rect 5940 11150 5950 11230
rect 5850 11140 5950 11150
rect 6050 11230 6150 11240
rect 6050 11150 6060 11230
rect 6140 11150 6150 11230
rect 6050 11140 6150 11150
rect 6250 11230 6350 11240
rect 6250 11150 6260 11230
rect 6340 11150 6350 11230
rect 6250 11140 6350 11150
rect 6450 11230 6550 11240
rect 6450 11150 6460 11230
rect 6540 11150 6550 11230
rect 6450 11140 6550 11150
rect -150 11045 -50 11055
rect -150 10965 -140 11045
rect -60 10965 -50 11045
rect -150 10955 -50 10965
rect 50 11045 150 11055
rect 50 10965 60 11045
rect 140 10965 150 11045
rect 50 10955 150 10965
rect 250 11045 350 11055
rect 250 10965 260 11045
rect 340 10965 350 11045
rect 250 10955 350 10965
rect 450 11045 550 11055
rect 450 10965 460 11045
rect 540 10965 550 11045
rect 450 10955 550 10965
rect 650 11045 750 11055
rect 650 10965 660 11045
rect 740 10965 750 11045
rect 650 10955 750 10965
rect 850 11045 950 11055
rect 850 10965 860 11045
rect 940 10965 950 11045
rect 850 10955 950 10965
rect 1050 11045 1150 11055
rect 1050 10965 1060 11045
rect 1140 10965 1150 11045
rect 1050 10955 1150 10965
rect 1250 11045 1350 11055
rect 1250 10965 1260 11045
rect 1340 10965 1350 11045
rect 1250 10955 1350 10965
rect 1450 11045 1550 11055
rect 1450 10965 1460 11045
rect 1540 10965 1550 11045
rect 1450 10955 1550 10965
rect 1650 11045 1750 11055
rect 1650 10965 1660 11045
rect 1740 10965 1750 11045
rect 1650 10955 1750 10965
rect 1850 11045 1950 11055
rect 1850 10965 1860 11045
rect 1940 10965 1950 11045
rect 1850 10955 1950 10965
rect 2050 11045 2150 11055
rect 2050 10965 2060 11045
rect 2140 10965 2150 11045
rect 2050 10955 2150 10965
rect 2250 11045 2350 11055
rect 2250 10965 2260 11045
rect 2340 10965 2350 11045
rect 2250 10955 2350 10965
rect 2450 11045 2550 11055
rect 2450 10965 2460 11045
rect 2540 10965 2550 11045
rect 2450 10955 2550 10965
rect 2650 11045 2750 11055
rect 2650 10965 2660 11045
rect 2740 10965 2750 11045
rect 2650 10955 2750 10965
rect 2850 11045 2950 11055
rect 2850 10965 2860 11045
rect 2940 10965 2950 11045
rect 2850 10955 2950 10965
rect 3050 11045 3150 11055
rect 3050 10965 3060 11045
rect 3140 10965 3150 11045
rect 3050 10955 3150 10965
rect 3250 11045 3350 11055
rect 3250 10965 3260 11045
rect 3340 10965 3350 11045
rect 3250 10955 3350 10965
rect 3450 11045 3550 11055
rect 3450 10965 3460 11045
rect 3540 10965 3550 11045
rect 3450 10955 3550 10965
rect 3650 11045 3750 11055
rect 3650 10965 3660 11045
rect 3740 10965 3750 11045
rect 3650 10955 3750 10965
rect 3850 11045 3950 11055
rect 3850 10965 3860 11045
rect 3940 10965 3950 11045
rect 3850 10955 3950 10965
rect 4050 11045 4150 11055
rect 4050 10965 4060 11045
rect 4140 10965 4150 11045
rect 4050 10955 4150 10965
rect 4250 11045 4350 11055
rect 4250 10965 4260 11045
rect 4340 10965 4350 11045
rect 4250 10955 4350 10965
rect 4450 11045 4550 11055
rect 4450 10965 4460 11045
rect 4540 10965 4550 11045
rect 4450 10955 4550 10965
rect 4650 11045 4750 11055
rect 4650 10965 4660 11045
rect 4740 10965 4750 11045
rect 4650 10955 4750 10965
rect 4850 11045 4950 11055
rect 4850 10965 4860 11045
rect 4940 10965 4950 11045
rect 4850 10955 4950 10965
rect 5050 11045 5150 11055
rect 5050 10965 5060 11045
rect 5140 10965 5150 11045
rect 5050 10955 5150 10965
rect 5250 11045 5350 11055
rect 5250 10965 5260 11045
rect 5340 10965 5350 11045
rect 5250 10955 5350 10965
rect 5450 11045 5550 11055
rect 5450 10965 5460 11045
rect 5540 10965 5550 11045
rect 5450 10955 5550 10965
rect 5650 11045 5750 11055
rect 5650 10965 5660 11045
rect 5740 10965 5750 11045
rect 5650 10955 5750 10965
rect 5850 11045 5950 11055
rect 5850 10965 5860 11045
rect 5940 10965 5950 11045
rect 5850 10955 5950 10965
rect 6050 11045 6150 11055
rect 6050 10965 6060 11045
rect 6140 10965 6150 11045
rect 6050 10955 6150 10965
rect 6250 11045 6350 11055
rect 6250 10965 6260 11045
rect 6340 10965 6350 11045
rect 6250 10955 6350 10965
rect 6450 11045 6550 11055
rect 6450 10965 6460 11045
rect 6540 10965 6550 11045
rect 6450 10955 6550 10965
rect -150 10860 -50 10870
rect -150 10780 -140 10860
rect -60 10780 -50 10860
rect -150 10770 -50 10780
rect 50 10860 150 10870
rect 50 10780 60 10860
rect 140 10780 150 10860
rect 50 10770 150 10780
rect 250 10860 350 10870
rect 250 10780 260 10860
rect 340 10780 350 10860
rect 250 10770 350 10780
rect 450 10860 550 10870
rect 450 10780 460 10860
rect 540 10780 550 10860
rect 450 10770 550 10780
rect 650 10860 750 10870
rect 650 10780 660 10860
rect 740 10780 750 10860
rect 650 10770 750 10780
rect 850 10860 950 10870
rect 850 10780 860 10860
rect 940 10780 950 10860
rect 850 10770 950 10780
rect 1050 10860 1150 10870
rect 1050 10780 1060 10860
rect 1140 10780 1150 10860
rect 1050 10770 1150 10780
rect 1250 10860 1350 10870
rect 1250 10780 1260 10860
rect 1340 10780 1350 10860
rect 1250 10770 1350 10780
rect 1450 10860 1550 10870
rect 1450 10780 1460 10860
rect 1540 10780 1550 10860
rect 1450 10770 1550 10780
rect 1650 10860 1750 10870
rect 1650 10780 1660 10860
rect 1740 10780 1750 10860
rect 1650 10770 1750 10780
rect 1850 10860 1950 10870
rect 1850 10780 1860 10860
rect 1940 10780 1950 10860
rect 1850 10770 1950 10780
rect 2050 10860 2150 10870
rect 2050 10780 2060 10860
rect 2140 10780 2150 10860
rect 2050 10770 2150 10780
rect 2250 10860 2350 10870
rect 2250 10780 2260 10860
rect 2340 10780 2350 10860
rect 2250 10770 2350 10780
rect 2450 10860 2550 10870
rect 2450 10780 2460 10860
rect 2540 10780 2550 10860
rect 2450 10770 2550 10780
rect 2650 10860 2750 10870
rect 2650 10780 2660 10860
rect 2740 10780 2750 10860
rect 2650 10770 2750 10780
rect 2850 10860 2950 10870
rect 2850 10780 2860 10860
rect 2940 10780 2950 10860
rect 2850 10770 2950 10780
rect 3050 10860 3150 10870
rect 3050 10780 3060 10860
rect 3140 10780 3150 10860
rect 3050 10770 3150 10780
rect 3250 10860 3350 10870
rect 3250 10780 3260 10860
rect 3340 10780 3350 10860
rect 3250 10770 3350 10780
rect 3450 10860 3550 10870
rect 3450 10780 3460 10860
rect 3540 10780 3550 10860
rect 3450 10770 3550 10780
rect 3650 10860 3750 10870
rect 3650 10780 3660 10860
rect 3740 10780 3750 10860
rect 3650 10770 3750 10780
rect 3850 10860 3950 10870
rect 3850 10780 3860 10860
rect 3940 10780 3950 10860
rect 3850 10770 3950 10780
rect 4050 10860 4150 10870
rect 4050 10780 4060 10860
rect 4140 10780 4150 10860
rect 4050 10770 4150 10780
rect 4250 10860 4350 10870
rect 4250 10780 4260 10860
rect 4340 10780 4350 10860
rect 4250 10770 4350 10780
rect 4450 10860 4550 10870
rect 4450 10780 4460 10860
rect 4540 10780 4550 10860
rect 4450 10770 4550 10780
rect 4650 10860 4750 10870
rect 4650 10780 4660 10860
rect 4740 10780 4750 10860
rect 4650 10770 4750 10780
rect 4850 10860 4950 10870
rect 4850 10780 4860 10860
rect 4940 10780 4950 10860
rect 4850 10770 4950 10780
rect 5050 10860 5150 10870
rect 5050 10780 5060 10860
rect 5140 10780 5150 10860
rect 5050 10770 5150 10780
rect 5250 10860 5350 10870
rect 5250 10780 5260 10860
rect 5340 10780 5350 10860
rect 5250 10770 5350 10780
rect 5450 10860 5550 10870
rect 5450 10780 5460 10860
rect 5540 10780 5550 10860
rect 5450 10770 5550 10780
rect 5650 10860 5750 10870
rect 5650 10780 5660 10860
rect 5740 10780 5750 10860
rect 5650 10770 5750 10780
rect 5850 10860 5950 10870
rect 5850 10780 5860 10860
rect 5940 10780 5950 10860
rect 5850 10770 5950 10780
rect 6050 10860 6150 10870
rect 6050 10780 6060 10860
rect 6140 10780 6150 10860
rect 6050 10770 6150 10780
rect 6250 10860 6350 10870
rect 6250 10780 6260 10860
rect 6340 10780 6350 10860
rect 6250 10770 6350 10780
rect 6450 10860 6550 10870
rect 6450 10780 6460 10860
rect 6540 10780 6550 10860
rect 6450 10770 6550 10780
rect -150 10675 -50 10685
rect -150 10595 -140 10675
rect -60 10595 -50 10675
rect -150 10585 -50 10595
rect 50 10675 150 10685
rect 50 10595 60 10675
rect 140 10595 150 10675
rect 50 10585 150 10595
rect 250 10675 350 10685
rect 250 10595 260 10675
rect 340 10595 350 10675
rect 250 10585 350 10595
rect 450 10675 550 10685
rect 450 10595 460 10675
rect 540 10595 550 10675
rect 450 10585 550 10595
rect 650 10675 750 10685
rect 650 10595 660 10675
rect 740 10595 750 10675
rect 650 10585 750 10595
rect 850 10675 950 10685
rect 850 10595 860 10675
rect 940 10595 950 10675
rect 850 10585 950 10595
rect 1050 10675 1150 10685
rect 1050 10595 1060 10675
rect 1140 10595 1150 10675
rect 1050 10585 1150 10595
rect 1250 10675 1350 10685
rect 1250 10595 1260 10675
rect 1340 10595 1350 10675
rect 1250 10585 1350 10595
rect 1450 10675 1550 10685
rect 1450 10595 1460 10675
rect 1540 10595 1550 10675
rect 1450 10585 1550 10595
rect 1650 10675 1750 10685
rect 1650 10595 1660 10675
rect 1740 10595 1750 10675
rect 1650 10585 1750 10595
rect 1850 10675 1950 10685
rect 1850 10595 1860 10675
rect 1940 10595 1950 10675
rect 1850 10585 1950 10595
rect 2050 10675 2150 10685
rect 2050 10595 2060 10675
rect 2140 10595 2150 10675
rect 2050 10585 2150 10595
rect 2250 10675 2350 10685
rect 2250 10595 2260 10675
rect 2340 10595 2350 10675
rect 2250 10585 2350 10595
rect 2450 10675 2550 10685
rect 2450 10595 2460 10675
rect 2540 10595 2550 10675
rect 2450 10585 2550 10595
rect 2650 10675 2750 10685
rect 2650 10595 2660 10675
rect 2740 10595 2750 10675
rect 2650 10585 2750 10595
rect 2850 10675 2950 10685
rect 2850 10595 2860 10675
rect 2940 10595 2950 10675
rect 2850 10585 2950 10595
rect 3050 10675 3150 10685
rect 3050 10595 3060 10675
rect 3140 10595 3150 10675
rect 3050 10585 3150 10595
rect 3250 10675 3350 10685
rect 3250 10595 3260 10675
rect 3340 10595 3350 10675
rect 3250 10585 3350 10595
rect 3450 10675 3550 10685
rect 3450 10595 3460 10675
rect 3540 10595 3550 10675
rect 3450 10585 3550 10595
rect 3650 10675 3750 10685
rect 3650 10595 3660 10675
rect 3740 10595 3750 10675
rect 3650 10585 3750 10595
rect 3850 10675 3950 10685
rect 3850 10595 3860 10675
rect 3940 10595 3950 10675
rect 3850 10585 3950 10595
rect 4050 10675 4150 10685
rect 4050 10595 4060 10675
rect 4140 10595 4150 10675
rect 4050 10585 4150 10595
rect 4250 10675 4350 10685
rect 4250 10595 4260 10675
rect 4340 10595 4350 10675
rect 4250 10585 4350 10595
rect 4450 10675 4550 10685
rect 4450 10595 4460 10675
rect 4540 10595 4550 10675
rect 4450 10585 4550 10595
rect 4650 10675 4750 10685
rect 4650 10595 4660 10675
rect 4740 10595 4750 10675
rect 4650 10585 4750 10595
rect 4850 10675 4950 10685
rect 4850 10595 4860 10675
rect 4940 10595 4950 10675
rect 4850 10585 4950 10595
rect 5050 10675 5150 10685
rect 5050 10595 5060 10675
rect 5140 10595 5150 10675
rect 5050 10585 5150 10595
rect 5250 10675 5350 10685
rect 5250 10595 5260 10675
rect 5340 10595 5350 10675
rect 5250 10585 5350 10595
rect 5450 10675 5550 10685
rect 5450 10595 5460 10675
rect 5540 10595 5550 10675
rect 5450 10585 5550 10595
rect 5650 10675 5750 10685
rect 5650 10595 5660 10675
rect 5740 10595 5750 10675
rect 5650 10585 5750 10595
rect 5850 10675 5950 10685
rect 5850 10595 5860 10675
rect 5940 10595 5950 10675
rect 5850 10585 5950 10595
rect 6050 10675 6150 10685
rect 6050 10595 6060 10675
rect 6140 10595 6150 10675
rect 6050 10585 6150 10595
rect 6250 10675 6350 10685
rect 6250 10595 6260 10675
rect 6340 10595 6350 10675
rect 6250 10585 6350 10595
rect 6450 10675 6550 10685
rect 6450 10595 6460 10675
rect 6540 10595 6550 10675
rect 6450 10585 6550 10595
rect -150 10490 -50 10500
rect -150 10410 -140 10490
rect -60 10410 -50 10490
rect -150 10400 -50 10410
rect 50 10490 150 10500
rect 50 10410 60 10490
rect 140 10410 150 10490
rect 50 10400 150 10410
rect 250 10490 350 10500
rect 250 10410 260 10490
rect 340 10410 350 10490
rect 250 10400 350 10410
rect 450 10490 550 10500
rect 450 10410 460 10490
rect 540 10410 550 10490
rect 450 10400 550 10410
rect 650 10490 750 10500
rect 650 10410 660 10490
rect 740 10410 750 10490
rect 650 10400 750 10410
rect 850 10490 950 10500
rect 850 10410 860 10490
rect 940 10410 950 10490
rect 850 10400 950 10410
rect 1050 10490 1150 10500
rect 1050 10410 1060 10490
rect 1140 10410 1150 10490
rect 1050 10400 1150 10410
rect 1250 10490 1350 10500
rect 1250 10410 1260 10490
rect 1340 10410 1350 10490
rect 1250 10400 1350 10410
rect 1450 10490 1550 10500
rect 1450 10410 1460 10490
rect 1540 10410 1550 10490
rect 1450 10400 1550 10410
rect 1650 10490 1750 10500
rect 1650 10410 1660 10490
rect 1740 10410 1750 10490
rect 1650 10400 1750 10410
rect 1850 10490 1950 10500
rect 1850 10410 1860 10490
rect 1940 10410 1950 10490
rect 1850 10400 1950 10410
rect 2050 10490 2150 10500
rect 2050 10410 2060 10490
rect 2140 10410 2150 10490
rect 2050 10400 2150 10410
rect 2250 10490 2350 10500
rect 2250 10410 2260 10490
rect 2340 10410 2350 10490
rect 2250 10400 2350 10410
rect 2450 10490 2550 10500
rect 2450 10410 2460 10490
rect 2540 10410 2550 10490
rect 2450 10400 2550 10410
rect 2650 10490 2750 10500
rect 2650 10410 2660 10490
rect 2740 10410 2750 10490
rect 2650 10400 2750 10410
rect 2850 10490 2950 10500
rect 2850 10410 2860 10490
rect 2940 10410 2950 10490
rect 2850 10400 2950 10410
rect 3050 10490 3150 10500
rect 3050 10410 3060 10490
rect 3140 10410 3150 10490
rect 3050 10400 3150 10410
rect 3250 10490 3350 10500
rect 3250 10410 3260 10490
rect 3340 10410 3350 10490
rect 3250 10400 3350 10410
rect 3450 10490 3550 10500
rect 3450 10410 3460 10490
rect 3540 10410 3550 10490
rect 3450 10400 3550 10410
rect 3650 10490 3750 10500
rect 3650 10410 3660 10490
rect 3740 10410 3750 10490
rect 3650 10400 3750 10410
rect 3850 10490 3950 10500
rect 3850 10410 3860 10490
rect 3940 10410 3950 10490
rect 3850 10400 3950 10410
rect 4050 10490 4150 10500
rect 4050 10410 4060 10490
rect 4140 10410 4150 10490
rect 4050 10400 4150 10410
rect 4250 10490 4350 10500
rect 4250 10410 4260 10490
rect 4340 10410 4350 10490
rect 4250 10400 4350 10410
rect 4450 10490 4550 10500
rect 4450 10410 4460 10490
rect 4540 10410 4550 10490
rect 4450 10400 4550 10410
rect 4650 10490 4750 10500
rect 4650 10410 4660 10490
rect 4740 10410 4750 10490
rect 4650 10400 4750 10410
rect 4850 10490 4950 10500
rect 4850 10410 4860 10490
rect 4940 10410 4950 10490
rect 4850 10400 4950 10410
rect 5050 10490 5150 10500
rect 5050 10410 5060 10490
rect 5140 10410 5150 10490
rect 5050 10400 5150 10410
rect 5250 10490 5350 10500
rect 5250 10410 5260 10490
rect 5340 10410 5350 10490
rect 5250 10400 5350 10410
rect 5450 10490 5550 10500
rect 5450 10410 5460 10490
rect 5540 10410 5550 10490
rect 5450 10400 5550 10410
rect 5650 10490 5750 10500
rect 5650 10410 5660 10490
rect 5740 10410 5750 10490
rect 5650 10400 5750 10410
rect 5850 10490 5950 10500
rect 5850 10410 5860 10490
rect 5940 10410 5950 10490
rect 5850 10400 5950 10410
rect 6050 10490 6150 10500
rect 6050 10410 6060 10490
rect 6140 10410 6150 10490
rect 6050 10400 6150 10410
rect 6250 10490 6350 10500
rect 6250 10410 6260 10490
rect 6340 10410 6350 10490
rect 6250 10400 6350 10410
rect 6450 10490 6550 10500
rect 6450 10410 6460 10490
rect 6540 10410 6550 10490
rect 6450 10400 6550 10410
rect -150 10305 -50 10315
rect -150 10225 -140 10305
rect -60 10225 -50 10305
rect -150 10215 -50 10225
rect 50 10305 150 10315
rect 50 10225 60 10305
rect 140 10225 150 10305
rect 50 10215 150 10225
rect 250 10305 350 10315
rect 250 10225 260 10305
rect 340 10225 350 10305
rect 250 10215 350 10225
rect 450 10305 550 10315
rect 450 10225 460 10305
rect 540 10225 550 10305
rect 450 10215 550 10225
rect 650 10305 750 10315
rect 650 10225 660 10305
rect 740 10225 750 10305
rect 650 10215 750 10225
rect 850 10305 950 10315
rect 850 10225 860 10305
rect 940 10225 950 10305
rect 850 10215 950 10225
rect 1050 10305 1150 10315
rect 1050 10225 1060 10305
rect 1140 10225 1150 10305
rect 1050 10215 1150 10225
rect 1250 10305 1350 10315
rect 1250 10225 1260 10305
rect 1340 10225 1350 10305
rect 1250 10215 1350 10225
rect 1450 10305 1550 10315
rect 1450 10225 1460 10305
rect 1540 10225 1550 10305
rect 1450 10215 1550 10225
rect 1650 10305 1750 10315
rect 1650 10225 1660 10305
rect 1740 10225 1750 10305
rect 1650 10215 1750 10225
rect 1850 10305 1950 10315
rect 1850 10225 1860 10305
rect 1940 10225 1950 10305
rect 1850 10215 1950 10225
rect 2050 10305 2150 10315
rect 2050 10225 2060 10305
rect 2140 10225 2150 10305
rect 2050 10215 2150 10225
rect 2250 10305 2350 10315
rect 2250 10225 2260 10305
rect 2340 10225 2350 10305
rect 2250 10215 2350 10225
rect 2450 10305 2550 10315
rect 2450 10225 2460 10305
rect 2540 10225 2550 10305
rect 2450 10215 2550 10225
rect 2650 10305 2750 10315
rect 2650 10225 2660 10305
rect 2740 10225 2750 10305
rect 2650 10215 2750 10225
rect 2850 10305 2950 10315
rect 2850 10225 2860 10305
rect 2940 10225 2950 10305
rect 2850 10215 2950 10225
rect 3050 10305 3150 10315
rect 3050 10225 3060 10305
rect 3140 10225 3150 10305
rect 3050 10215 3150 10225
rect 3250 10305 3350 10315
rect 3250 10225 3260 10305
rect 3340 10225 3350 10305
rect 3250 10215 3350 10225
rect 3450 10305 3550 10315
rect 3450 10225 3460 10305
rect 3540 10225 3550 10305
rect 3450 10215 3550 10225
rect 3650 10305 3750 10315
rect 3650 10225 3660 10305
rect 3740 10225 3750 10305
rect 3650 10215 3750 10225
rect 3850 10305 3950 10315
rect 3850 10225 3860 10305
rect 3940 10225 3950 10305
rect 3850 10215 3950 10225
rect 4050 10305 4150 10315
rect 4050 10225 4060 10305
rect 4140 10225 4150 10305
rect 4050 10215 4150 10225
rect 4250 10305 4350 10315
rect 4250 10225 4260 10305
rect 4340 10225 4350 10305
rect 4250 10215 4350 10225
rect 4450 10305 4550 10315
rect 4450 10225 4460 10305
rect 4540 10225 4550 10305
rect 4450 10215 4550 10225
rect 4650 10305 4750 10315
rect 4650 10225 4660 10305
rect 4740 10225 4750 10305
rect 4650 10215 4750 10225
rect 4850 10305 4950 10315
rect 4850 10225 4860 10305
rect 4940 10225 4950 10305
rect 4850 10215 4950 10225
rect 5050 10305 5150 10315
rect 5050 10225 5060 10305
rect 5140 10225 5150 10305
rect 5050 10215 5150 10225
rect 5250 10305 5350 10315
rect 5250 10225 5260 10305
rect 5340 10225 5350 10305
rect 5250 10215 5350 10225
rect 5450 10305 5550 10315
rect 5450 10225 5460 10305
rect 5540 10225 5550 10305
rect 5450 10215 5550 10225
rect 5650 10305 5750 10315
rect 5650 10225 5660 10305
rect 5740 10225 5750 10305
rect 5650 10215 5750 10225
rect 5850 10305 5950 10315
rect 5850 10225 5860 10305
rect 5940 10225 5950 10305
rect 5850 10215 5950 10225
rect 6050 10305 6150 10315
rect 6050 10225 6060 10305
rect 6140 10225 6150 10305
rect 6050 10215 6150 10225
rect 6250 10305 6350 10315
rect 6250 10225 6260 10305
rect 6340 10225 6350 10305
rect 6250 10215 6350 10225
rect 6450 10305 6550 10315
rect 6450 10225 6460 10305
rect 6540 10225 6550 10305
rect 6450 10215 6550 10225
rect -150 10120 -50 10130
rect -150 10040 -140 10120
rect -60 10040 -50 10120
rect -150 10030 -50 10040
rect 50 10120 150 10130
rect 50 10040 60 10120
rect 140 10040 150 10120
rect 50 10030 150 10040
rect 250 10120 350 10130
rect 250 10040 260 10120
rect 340 10040 350 10120
rect 250 10030 350 10040
rect 450 10120 550 10130
rect 450 10040 460 10120
rect 540 10040 550 10120
rect 450 10030 550 10040
rect 650 10120 750 10130
rect 650 10040 660 10120
rect 740 10040 750 10120
rect 650 10030 750 10040
rect 850 10120 950 10130
rect 850 10040 860 10120
rect 940 10040 950 10120
rect 850 10030 950 10040
rect 1050 10120 1150 10130
rect 1050 10040 1060 10120
rect 1140 10040 1150 10120
rect 1050 10030 1150 10040
rect 1250 10120 1350 10130
rect 1250 10040 1260 10120
rect 1340 10040 1350 10120
rect 1250 10030 1350 10040
rect 1450 10120 1550 10130
rect 1450 10040 1460 10120
rect 1540 10040 1550 10120
rect 1450 10030 1550 10040
rect 1650 10120 1750 10130
rect 1650 10040 1660 10120
rect 1740 10040 1750 10120
rect 1650 10030 1750 10040
rect 1850 10120 1950 10130
rect 1850 10040 1860 10120
rect 1940 10040 1950 10120
rect 1850 10030 1950 10040
rect 2050 10120 2150 10130
rect 2050 10040 2060 10120
rect 2140 10040 2150 10120
rect 2050 10030 2150 10040
rect 2250 10120 2350 10130
rect 2250 10040 2260 10120
rect 2340 10040 2350 10120
rect 2250 10030 2350 10040
rect 2450 10120 2550 10130
rect 2450 10040 2460 10120
rect 2540 10040 2550 10120
rect 2450 10030 2550 10040
rect 2650 10120 2750 10130
rect 2650 10040 2660 10120
rect 2740 10040 2750 10120
rect 2650 10030 2750 10040
rect 2850 10120 2950 10130
rect 2850 10040 2860 10120
rect 2940 10040 2950 10120
rect 2850 10030 2950 10040
rect 3050 10120 3150 10130
rect 3050 10040 3060 10120
rect 3140 10040 3150 10120
rect 3050 10030 3150 10040
rect 3250 10120 3350 10130
rect 3250 10040 3260 10120
rect 3340 10040 3350 10120
rect 3250 10030 3350 10040
rect 3450 10120 3550 10130
rect 3450 10040 3460 10120
rect 3540 10040 3550 10120
rect 3450 10030 3550 10040
rect 3650 10120 3750 10130
rect 3650 10040 3660 10120
rect 3740 10040 3750 10120
rect 3650 10030 3750 10040
rect 3850 10120 3950 10130
rect 3850 10040 3860 10120
rect 3940 10040 3950 10120
rect 3850 10030 3950 10040
rect 4050 10120 4150 10130
rect 4050 10040 4060 10120
rect 4140 10040 4150 10120
rect 4050 10030 4150 10040
rect 4250 10120 4350 10130
rect 4250 10040 4260 10120
rect 4340 10040 4350 10120
rect 4250 10030 4350 10040
rect 4450 10120 4550 10130
rect 4450 10040 4460 10120
rect 4540 10040 4550 10120
rect 4450 10030 4550 10040
rect 4650 10120 4750 10130
rect 4650 10040 4660 10120
rect 4740 10040 4750 10120
rect 4650 10030 4750 10040
rect 4850 10120 4950 10130
rect 4850 10040 4860 10120
rect 4940 10040 4950 10120
rect 4850 10030 4950 10040
rect 5050 10120 5150 10130
rect 5050 10040 5060 10120
rect 5140 10040 5150 10120
rect 5050 10030 5150 10040
rect 5250 10120 5350 10130
rect 5250 10040 5260 10120
rect 5340 10040 5350 10120
rect 5250 10030 5350 10040
rect 5450 10120 5550 10130
rect 5450 10040 5460 10120
rect 5540 10040 5550 10120
rect 5450 10030 5550 10040
rect 5650 10120 5750 10130
rect 5650 10040 5660 10120
rect 5740 10040 5750 10120
rect 5650 10030 5750 10040
rect 5850 10120 5950 10130
rect 5850 10040 5860 10120
rect 5940 10040 5950 10120
rect 5850 10030 5950 10040
rect 6050 10120 6150 10130
rect 6050 10040 6060 10120
rect 6140 10040 6150 10120
rect 6050 10030 6150 10040
rect 6250 10120 6350 10130
rect 6250 10040 6260 10120
rect 6340 10040 6350 10120
rect 6250 10030 6350 10040
rect 6450 10120 6550 10130
rect 6450 10040 6460 10120
rect 6540 10040 6550 10120
rect 6450 10030 6550 10040
rect -150 9935 -50 9945
rect -150 9855 -140 9935
rect -60 9855 -50 9935
rect -150 9845 -50 9855
rect 50 9935 150 9945
rect 50 9855 60 9935
rect 140 9855 150 9935
rect 50 9845 150 9855
rect 250 9935 350 9945
rect 250 9855 260 9935
rect 340 9855 350 9935
rect 250 9845 350 9855
rect 450 9935 550 9945
rect 450 9855 460 9935
rect 540 9855 550 9935
rect 450 9845 550 9855
rect 650 9935 750 9945
rect 650 9855 660 9935
rect 740 9855 750 9935
rect 650 9845 750 9855
rect 850 9935 950 9945
rect 850 9855 860 9935
rect 940 9855 950 9935
rect 850 9845 950 9855
rect 1050 9935 1150 9945
rect 1050 9855 1060 9935
rect 1140 9855 1150 9935
rect 1050 9845 1150 9855
rect 1250 9935 1350 9945
rect 1250 9855 1260 9935
rect 1340 9855 1350 9935
rect 1250 9845 1350 9855
rect 1450 9935 1550 9945
rect 1450 9855 1460 9935
rect 1540 9855 1550 9935
rect 1450 9845 1550 9855
rect 1650 9935 1750 9945
rect 1650 9855 1660 9935
rect 1740 9855 1750 9935
rect 1650 9845 1750 9855
rect 1850 9935 1950 9945
rect 1850 9855 1860 9935
rect 1940 9855 1950 9935
rect 1850 9845 1950 9855
rect 2050 9935 2150 9945
rect 2050 9855 2060 9935
rect 2140 9855 2150 9935
rect 2050 9845 2150 9855
rect 2250 9935 2350 9945
rect 2250 9855 2260 9935
rect 2340 9855 2350 9935
rect 2250 9845 2350 9855
rect 2450 9935 2550 9945
rect 2450 9855 2460 9935
rect 2540 9855 2550 9935
rect 2450 9845 2550 9855
rect 2650 9935 2750 9945
rect 2650 9855 2660 9935
rect 2740 9855 2750 9935
rect 2650 9845 2750 9855
rect 2850 9935 2950 9945
rect 2850 9855 2860 9935
rect 2940 9855 2950 9935
rect 2850 9845 2950 9855
rect 3050 9935 3150 9945
rect 3050 9855 3060 9935
rect 3140 9855 3150 9935
rect 3050 9845 3150 9855
rect 3250 9935 3350 9945
rect 3250 9855 3260 9935
rect 3340 9855 3350 9935
rect 3250 9845 3350 9855
rect 3450 9935 3550 9945
rect 3450 9855 3460 9935
rect 3540 9855 3550 9935
rect 3450 9845 3550 9855
rect 3650 9935 3750 9945
rect 3650 9855 3660 9935
rect 3740 9855 3750 9935
rect 3650 9845 3750 9855
rect 3850 9935 3950 9945
rect 3850 9855 3860 9935
rect 3940 9855 3950 9935
rect 3850 9845 3950 9855
rect 4050 9935 4150 9945
rect 4050 9855 4060 9935
rect 4140 9855 4150 9935
rect 4050 9845 4150 9855
rect 4250 9935 4350 9945
rect 4250 9855 4260 9935
rect 4340 9855 4350 9935
rect 4250 9845 4350 9855
rect 4450 9935 4550 9945
rect 4450 9855 4460 9935
rect 4540 9855 4550 9935
rect 4450 9845 4550 9855
rect 4650 9935 4750 9945
rect 4650 9855 4660 9935
rect 4740 9855 4750 9935
rect 4650 9845 4750 9855
rect 4850 9935 4950 9945
rect 4850 9855 4860 9935
rect 4940 9855 4950 9935
rect 4850 9845 4950 9855
rect 5050 9935 5150 9945
rect 5050 9855 5060 9935
rect 5140 9855 5150 9935
rect 5050 9845 5150 9855
rect 5250 9935 5350 9945
rect 5250 9855 5260 9935
rect 5340 9855 5350 9935
rect 5250 9845 5350 9855
rect 5450 9935 5550 9945
rect 5450 9855 5460 9935
rect 5540 9855 5550 9935
rect 5450 9845 5550 9855
rect 5650 9935 5750 9945
rect 5650 9855 5660 9935
rect 5740 9855 5750 9935
rect 5650 9845 5750 9855
rect 5850 9935 5950 9945
rect 5850 9855 5860 9935
rect 5940 9855 5950 9935
rect 5850 9845 5950 9855
rect 6050 9935 6150 9945
rect 6050 9855 6060 9935
rect 6140 9855 6150 9935
rect 6050 9845 6150 9855
rect 6250 9935 6350 9945
rect 6250 9855 6260 9935
rect 6340 9855 6350 9935
rect 6250 9845 6350 9855
rect 6450 9935 6550 9945
rect 6450 9855 6460 9935
rect 6540 9855 6550 9935
rect 6450 9845 6550 9855
rect -150 9750 -50 9760
rect -150 9670 -140 9750
rect -60 9670 -50 9750
rect -150 9660 -50 9670
rect 50 9750 150 9760
rect 50 9670 60 9750
rect 140 9670 150 9750
rect 50 9660 150 9670
rect 250 9750 350 9760
rect 250 9670 260 9750
rect 340 9670 350 9750
rect 250 9660 350 9670
rect 450 9750 550 9760
rect 450 9670 460 9750
rect 540 9670 550 9750
rect 450 9660 550 9670
rect 650 9750 750 9760
rect 650 9670 660 9750
rect 740 9670 750 9750
rect 650 9660 750 9670
rect 850 9750 950 9760
rect 850 9670 860 9750
rect 940 9670 950 9750
rect 850 9660 950 9670
rect 1050 9750 1150 9760
rect 1050 9670 1060 9750
rect 1140 9670 1150 9750
rect 1050 9660 1150 9670
rect 1250 9750 1350 9760
rect 1250 9670 1260 9750
rect 1340 9670 1350 9750
rect 1250 9660 1350 9670
rect 1450 9750 1550 9760
rect 1450 9670 1460 9750
rect 1540 9670 1550 9750
rect 1450 9660 1550 9670
rect 1650 9750 1750 9760
rect 1650 9670 1660 9750
rect 1740 9670 1750 9750
rect 1650 9660 1750 9670
rect 1850 9750 1950 9760
rect 1850 9670 1860 9750
rect 1940 9670 1950 9750
rect 1850 9660 1950 9670
rect 2050 9750 2150 9760
rect 2050 9670 2060 9750
rect 2140 9670 2150 9750
rect 2050 9660 2150 9670
rect 2250 9750 2350 9760
rect 2250 9670 2260 9750
rect 2340 9670 2350 9750
rect 2250 9660 2350 9670
rect 2450 9750 2550 9760
rect 2450 9670 2460 9750
rect 2540 9670 2550 9750
rect 2450 9660 2550 9670
rect 2650 9750 2750 9760
rect 2650 9670 2660 9750
rect 2740 9670 2750 9750
rect 2650 9660 2750 9670
rect 2850 9750 2950 9760
rect 2850 9670 2860 9750
rect 2940 9670 2950 9750
rect 2850 9660 2950 9670
rect 3050 9750 3150 9760
rect 3050 9670 3060 9750
rect 3140 9670 3150 9750
rect 3050 9660 3150 9670
rect 3250 9750 3350 9760
rect 3250 9670 3260 9750
rect 3340 9670 3350 9750
rect 3250 9660 3350 9670
rect 3450 9750 3550 9760
rect 3450 9670 3460 9750
rect 3540 9670 3550 9750
rect 3450 9660 3550 9670
rect 3650 9750 3750 9760
rect 3650 9670 3660 9750
rect 3740 9670 3750 9750
rect 3650 9660 3750 9670
rect 3850 9750 3950 9760
rect 3850 9670 3860 9750
rect 3940 9670 3950 9750
rect 3850 9660 3950 9670
rect 4050 9750 4150 9760
rect 4050 9670 4060 9750
rect 4140 9670 4150 9750
rect 4050 9660 4150 9670
rect 4250 9750 4350 9760
rect 4250 9670 4260 9750
rect 4340 9670 4350 9750
rect 4250 9660 4350 9670
rect 4450 9750 4550 9760
rect 4450 9670 4460 9750
rect 4540 9670 4550 9750
rect 4450 9660 4550 9670
rect 4650 9750 4750 9760
rect 4650 9670 4660 9750
rect 4740 9670 4750 9750
rect 4650 9660 4750 9670
rect 4850 9750 4950 9760
rect 4850 9670 4860 9750
rect 4940 9670 4950 9750
rect 4850 9660 4950 9670
rect 5050 9750 5150 9760
rect 5050 9670 5060 9750
rect 5140 9670 5150 9750
rect 5050 9660 5150 9670
rect 5250 9750 5350 9760
rect 5250 9670 5260 9750
rect 5340 9670 5350 9750
rect 5250 9660 5350 9670
rect 5450 9750 5550 9760
rect 5450 9670 5460 9750
rect 5540 9670 5550 9750
rect 5450 9660 5550 9670
rect 5650 9750 5750 9760
rect 5650 9670 5660 9750
rect 5740 9670 5750 9750
rect 5650 9660 5750 9670
rect 5850 9750 5950 9760
rect 5850 9670 5860 9750
rect 5940 9670 5950 9750
rect 5850 9660 5950 9670
rect 6050 9750 6150 9760
rect 6050 9670 6060 9750
rect 6140 9670 6150 9750
rect 6050 9660 6150 9670
rect 6250 9750 6350 9760
rect 6250 9670 6260 9750
rect 6340 9670 6350 9750
rect 6250 9660 6350 9670
rect 6450 9750 6550 9760
rect 6450 9670 6460 9750
rect 6540 9670 6550 9750
rect 6450 9660 6550 9670
rect -150 9565 -50 9575
rect -150 9485 -140 9565
rect -60 9485 -50 9565
rect -150 9475 -50 9485
rect 50 9565 150 9575
rect 50 9485 60 9565
rect 140 9485 150 9565
rect 50 9475 150 9485
rect 250 9565 350 9575
rect 250 9485 260 9565
rect 340 9485 350 9565
rect 250 9475 350 9485
rect 450 9565 550 9575
rect 450 9485 460 9565
rect 540 9485 550 9565
rect 450 9475 550 9485
rect 650 9565 750 9575
rect 650 9485 660 9565
rect 740 9485 750 9565
rect 650 9475 750 9485
rect 850 9565 950 9575
rect 850 9485 860 9565
rect 940 9485 950 9565
rect 850 9475 950 9485
rect 1050 9565 1150 9575
rect 1050 9485 1060 9565
rect 1140 9485 1150 9565
rect 1050 9475 1150 9485
rect 1250 9565 1350 9575
rect 1250 9485 1260 9565
rect 1340 9485 1350 9565
rect 1250 9475 1350 9485
rect 1450 9565 1550 9575
rect 1450 9485 1460 9565
rect 1540 9485 1550 9565
rect 1450 9475 1550 9485
rect 1650 9565 1750 9575
rect 1650 9485 1660 9565
rect 1740 9485 1750 9565
rect 1650 9475 1750 9485
rect 1850 9565 1950 9575
rect 1850 9485 1860 9565
rect 1940 9485 1950 9565
rect 1850 9475 1950 9485
rect 2050 9565 2150 9575
rect 2050 9485 2060 9565
rect 2140 9485 2150 9565
rect 2050 9475 2150 9485
rect 2250 9565 2350 9575
rect 2250 9485 2260 9565
rect 2340 9485 2350 9565
rect 2250 9475 2350 9485
rect 2450 9565 2550 9575
rect 2450 9485 2460 9565
rect 2540 9485 2550 9565
rect 2450 9475 2550 9485
rect 2650 9565 2750 9575
rect 2650 9485 2660 9565
rect 2740 9485 2750 9565
rect 2650 9475 2750 9485
rect 2850 9565 2950 9575
rect 2850 9485 2860 9565
rect 2940 9485 2950 9565
rect 2850 9475 2950 9485
rect 3050 9565 3150 9575
rect 3050 9485 3060 9565
rect 3140 9485 3150 9565
rect 3050 9475 3150 9485
rect 3250 9565 3350 9575
rect 3250 9485 3260 9565
rect 3340 9485 3350 9565
rect 3250 9475 3350 9485
rect 3450 9565 3550 9575
rect 3450 9485 3460 9565
rect 3540 9485 3550 9565
rect 3450 9475 3550 9485
rect 3650 9565 3750 9575
rect 3650 9485 3660 9565
rect 3740 9485 3750 9565
rect 3650 9475 3750 9485
rect 3850 9565 3950 9575
rect 3850 9485 3860 9565
rect 3940 9485 3950 9565
rect 3850 9475 3950 9485
rect 4050 9565 4150 9575
rect 4050 9485 4060 9565
rect 4140 9485 4150 9565
rect 4050 9475 4150 9485
rect 4250 9565 4350 9575
rect 4250 9485 4260 9565
rect 4340 9485 4350 9565
rect 4250 9475 4350 9485
rect 4450 9565 4550 9575
rect 4450 9485 4460 9565
rect 4540 9485 4550 9565
rect 4450 9475 4550 9485
rect 4650 9565 4750 9575
rect 4650 9485 4660 9565
rect 4740 9485 4750 9565
rect 4650 9475 4750 9485
rect 4850 9565 4950 9575
rect 4850 9485 4860 9565
rect 4940 9485 4950 9565
rect 4850 9475 4950 9485
rect 5050 9565 5150 9575
rect 5050 9485 5060 9565
rect 5140 9485 5150 9565
rect 5050 9475 5150 9485
rect 5250 9565 5350 9575
rect 5250 9485 5260 9565
rect 5340 9485 5350 9565
rect 5250 9475 5350 9485
rect 5450 9565 5550 9575
rect 5450 9485 5460 9565
rect 5540 9485 5550 9565
rect 5450 9475 5550 9485
rect 5650 9565 5750 9575
rect 5650 9485 5660 9565
rect 5740 9485 5750 9565
rect 5650 9475 5750 9485
rect 5850 9565 5950 9575
rect 5850 9485 5860 9565
rect 5940 9485 5950 9565
rect 5850 9475 5950 9485
rect 6050 9565 6150 9575
rect 6050 9485 6060 9565
rect 6140 9485 6150 9565
rect 6050 9475 6150 9485
rect 6250 9565 6350 9575
rect 6250 9485 6260 9565
rect 6340 9485 6350 9565
rect 6250 9475 6350 9485
rect 6450 9565 6550 9575
rect 6450 9485 6460 9565
rect 6540 9485 6550 9565
rect 6450 9475 6550 9485
rect -150 9380 -50 9390
rect -150 9300 -140 9380
rect -60 9300 -50 9380
rect -150 9290 -50 9300
rect 50 9380 150 9390
rect 50 9300 60 9380
rect 140 9300 150 9380
rect 50 9290 150 9300
rect 250 9380 350 9390
rect 250 9300 260 9380
rect 340 9300 350 9380
rect 250 9290 350 9300
rect 450 9380 550 9390
rect 450 9300 460 9380
rect 540 9300 550 9380
rect 450 9290 550 9300
rect 650 9380 750 9390
rect 650 9300 660 9380
rect 740 9300 750 9380
rect 650 9290 750 9300
rect 850 9380 950 9390
rect 850 9300 860 9380
rect 940 9300 950 9380
rect 850 9290 950 9300
rect 1050 9380 1150 9390
rect 1050 9300 1060 9380
rect 1140 9300 1150 9380
rect 1050 9290 1150 9300
rect 1250 9380 1350 9390
rect 1250 9300 1260 9380
rect 1340 9300 1350 9380
rect 1250 9290 1350 9300
rect 1450 9380 1550 9390
rect 1450 9300 1460 9380
rect 1540 9300 1550 9380
rect 1450 9290 1550 9300
rect 1650 9380 1750 9390
rect 1650 9300 1660 9380
rect 1740 9300 1750 9380
rect 1650 9290 1750 9300
rect 1850 9380 1950 9390
rect 1850 9300 1860 9380
rect 1940 9300 1950 9380
rect 1850 9290 1950 9300
rect 2050 9380 2150 9390
rect 2050 9300 2060 9380
rect 2140 9300 2150 9380
rect 2050 9290 2150 9300
rect 2250 9380 2350 9390
rect 2250 9300 2260 9380
rect 2340 9300 2350 9380
rect 2250 9290 2350 9300
rect 2450 9380 2550 9390
rect 2450 9300 2460 9380
rect 2540 9300 2550 9380
rect 2450 9290 2550 9300
rect 2650 9380 2750 9390
rect 2650 9300 2660 9380
rect 2740 9300 2750 9380
rect 2650 9290 2750 9300
rect 2850 9380 2950 9390
rect 2850 9300 2860 9380
rect 2940 9300 2950 9380
rect 2850 9290 2950 9300
rect 3050 9380 3150 9390
rect 3050 9300 3060 9380
rect 3140 9300 3150 9380
rect 3050 9290 3150 9300
rect 3250 9380 3350 9390
rect 3250 9300 3260 9380
rect 3340 9300 3350 9380
rect 3250 9290 3350 9300
rect 3450 9380 3550 9390
rect 3450 9300 3460 9380
rect 3540 9300 3550 9380
rect 3450 9290 3550 9300
rect 3650 9380 3750 9390
rect 3650 9300 3660 9380
rect 3740 9300 3750 9380
rect 3650 9290 3750 9300
rect 3850 9380 3950 9390
rect 3850 9300 3860 9380
rect 3940 9300 3950 9380
rect 3850 9290 3950 9300
rect 4050 9380 4150 9390
rect 4050 9300 4060 9380
rect 4140 9300 4150 9380
rect 4050 9290 4150 9300
rect 4250 9380 4350 9390
rect 4250 9300 4260 9380
rect 4340 9300 4350 9380
rect 4250 9290 4350 9300
rect 4450 9380 4550 9390
rect 4450 9300 4460 9380
rect 4540 9300 4550 9380
rect 4450 9290 4550 9300
rect 4650 9380 4750 9390
rect 4650 9300 4660 9380
rect 4740 9300 4750 9380
rect 4650 9290 4750 9300
rect 4850 9380 4950 9390
rect 4850 9300 4860 9380
rect 4940 9300 4950 9380
rect 4850 9290 4950 9300
rect 5050 9380 5150 9390
rect 5050 9300 5060 9380
rect 5140 9300 5150 9380
rect 5050 9290 5150 9300
rect 5250 9380 5350 9390
rect 5250 9300 5260 9380
rect 5340 9300 5350 9380
rect 5250 9290 5350 9300
rect 5450 9380 5550 9390
rect 5450 9300 5460 9380
rect 5540 9300 5550 9380
rect 5450 9290 5550 9300
rect 5650 9380 5750 9390
rect 5650 9300 5660 9380
rect 5740 9300 5750 9380
rect 5650 9290 5750 9300
rect 5850 9380 5950 9390
rect 5850 9300 5860 9380
rect 5940 9300 5950 9380
rect 5850 9290 5950 9300
rect 6050 9380 6150 9390
rect 6050 9300 6060 9380
rect 6140 9300 6150 9380
rect 6050 9290 6150 9300
rect 6250 9380 6350 9390
rect 6250 9300 6260 9380
rect 6340 9300 6350 9380
rect 6250 9290 6350 9300
rect 6450 9380 6550 9390
rect 6450 9300 6460 9380
rect 6540 9300 6550 9380
rect 6450 9290 6550 9300
rect -150 9195 -50 9205
rect -150 9115 -140 9195
rect -60 9115 -50 9195
rect -150 9105 -50 9115
rect 50 9195 150 9205
rect 50 9115 60 9195
rect 140 9115 150 9195
rect 50 9105 150 9115
rect 250 9195 350 9205
rect 250 9115 260 9195
rect 340 9115 350 9195
rect 250 9105 350 9115
rect 450 9195 550 9205
rect 450 9115 460 9195
rect 540 9115 550 9195
rect 450 9105 550 9115
rect 650 9195 750 9205
rect 650 9115 660 9195
rect 740 9115 750 9195
rect 650 9105 750 9115
rect 850 9195 950 9205
rect 850 9115 860 9195
rect 940 9115 950 9195
rect 850 9105 950 9115
rect 1050 9195 1150 9205
rect 1050 9115 1060 9195
rect 1140 9115 1150 9195
rect 1050 9105 1150 9115
rect 1250 9195 1350 9205
rect 1250 9115 1260 9195
rect 1340 9115 1350 9195
rect 1250 9105 1350 9115
rect 1450 9195 1550 9205
rect 1450 9115 1460 9195
rect 1540 9115 1550 9195
rect 1450 9105 1550 9115
rect 1650 9195 1750 9205
rect 1650 9115 1660 9195
rect 1740 9115 1750 9195
rect 1650 9105 1750 9115
rect 1850 9195 1950 9205
rect 1850 9115 1860 9195
rect 1940 9115 1950 9195
rect 1850 9105 1950 9115
rect 2050 9195 2150 9205
rect 2050 9115 2060 9195
rect 2140 9115 2150 9195
rect 2050 9105 2150 9115
rect 2250 9195 2350 9205
rect 2250 9115 2260 9195
rect 2340 9115 2350 9195
rect 2250 9105 2350 9115
rect 2450 9195 2550 9205
rect 2450 9115 2460 9195
rect 2540 9115 2550 9195
rect 2450 9105 2550 9115
rect 2650 9195 2750 9205
rect 2650 9115 2660 9195
rect 2740 9115 2750 9195
rect 2650 9105 2750 9115
rect 2850 9195 2950 9205
rect 2850 9115 2860 9195
rect 2940 9115 2950 9195
rect 2850 9105 2950 9115
rect 3050 9195 3150 9205
rect 3050 9115 3060 9195
rect 3140 9115 3150 9195
rect 3050 9105 3150 9115
rect 3250 9195 3350 9205
rect 3250 9115 3260 9195
rect 3340 9115 3350 9195
rect 3250 9105 3350 9115
rect 3450 9195 3550 9205
rect 3450 9115 3460 9195
rect 3540 9115 3550 9195
rect 3450 9105 3550 9115
rect 3650 9195 3750 9205
rect 3650 9115 3660 9195
rect 3740 9115 3750 9195
rect 3650 9105 3750 9115
rect 3850 9195 3950 9205
rect 3850 9115 3860 9195
rect 3940 9115 3950 9195
rect 3850 9105 3950 9115
rect 4050 9195 4150 9205
rect 4050 9115 4060 9195
rect 4140 9115 4150 9195
rect 4050 9105 4150 9115
rect 4250 9195 4350 9205
rect 4250 9115 4260 9195
rect 4340 9115 4350 9195
rect 4250 9105 4350 9115
rect 4450 9195 4550 9205
rect 4450 9115 4460 9195
rect 4540 9115 4550 9195
rect 4450 9105 4550 9115
rect 4650 9195 4750 9205
rect 4650 9115 4660 9195
rect 4740 9115 4750 9195
rect 4650 9105 4750 9115
rect 4850 9195 4950 9205
rect 4850 9115 4860 9195
rect 4940 9115 4950 9195
rect 4850 9105 4950 9115
rect 5050 9195 5150 9205
rect 5050 9115 5060 9195
rect 5140 9115 5150 9195
rect 5050 9105 5150 9115
rect 5250 9195 5350 9205
rect 5250 9115 5260 9195
rect 5340 9115 5350 9195
rect 5250 9105 5350 9115
rect 5450 9195 5550 9205
rect 5450 9115 5460 9195
rect 5540 9115 5550 9195
rect 5450 9105 5550 9115
rect 5650 9195 5750 9205
rect 5650 9115 5660 9195
rect 5740 9115 5750 9195
rect 5650 9105 5750 9115
rect 5850 9195 5950 9205
rect 5850 9115 5860 9195
rect 5940 9115 5950 9195
rect 5850 9105 5950 9115
rect 6050 9195 6150 9205
rect 6050 9115 6060 9195
rect 6140 9115 6150 9195
rect 6050 9105 6150 9115
rect 6250 9195 6350 9205
rect 6250 9115 6260 9195
rect 6340 9115 6350 9195
rect 6250 9105 6350 9115
rect 6450 9195 6550 9205
rect 6450 9115 6460 9195
rect 6540 9115 6550 9195
rect 6450 9105 6550 9115
rect -150 9010 -50 9020
rect -150 8930 -140 9010
rect -60 8930 -50 9010
rect -150 8920 -50 8930
rect 50 9010 150 9020
rect 50 8930 60 9010
rect 140 8930 150 9010
rect 50 8920 150 8930
rect 250 9010 350 9020
rect 250 8930 260 9010
rect 340 8930 350 9010
rect 250 8920 350 8930
rect 450 9010 550 9020
rect 450 8930 460 9010
rect 540 8930 550 9010
rect 450 8920 550 8930
rect 650 9010 750 9020
rect 650 8930 660 9010
rect 740 8930 750 9010
rect 650 8920 750 8930
rect 850 9010 950 9020
rect 850 8930 860 9010
rect 940 8930 950 9010
rect 850 8920 950 8930
rect 1050 9010 1150 9020
rect 1050 8930 1060 9010
rect 1140 8930 1150 9010
rect 1050 8920 1150 8930
rect 1250 9010 1350 9020
rect 1250 8930 1260 9010
rect 1340 8930 1350 9010
rect 1250 8920 1350 8930
rect 1450 9010 1550 9020
rect 1450 8930 1460 9010
rect 1540 8930 1550 9010
rect 1450 8920 1550 8930
rect 1650 9010 1750 9020
rect 1650 8930 1660 9010
rect 1740 8930 1750 9010
rect 1650 8920 1750 8930
rect 1850 9010 1950 9020
rect 1850 8930 1860 9010
rect 1940 8930 1950 9010
rect 1850 8920 1950 8930
rect 2050 9010 2150 9020
rect 2050 8930 2060 9010
rect 2140 8930 2150 9010
rect 2050 8920 2150 8930
rect 2250 9010 2350 9020
rect 2250 8930 2260 9010
rect 2340 8930 2350 9010
rect 2250 8920 2350 8930
rect 2450 9010 2550 9020
rect 2450 8930 2460 9010
rect 2540 8930 2550 9010
rect 2450 8920 2550 8930
rect 2650 9010 2750 9020
rect 2650 8930 2660 9010
rect 2740 8930 2750 9010
rect 2650 8920 2750 8930
rect 2850 9010 2950 9020
rect 2850 8930 2860 9010
rect 2940 8930 2950 9010
rect 2850 8920 2950 8930
rect 3050 9010 3150 9020
rect 3050 8930 3060 9010
rect 3140 8930 3150 9010
rect 3050 8920 3150 8930
rect 3250 9010 3350 9020
rect 3250 8930 3260 9010
rect 3340 8930 3350 9010
rect 3250 8920 3350 8930
rect 3450 9010 3550 9020
rect 3450 8930 3460 9010
rect 3540 8930 3550 9010
rect 3450 8920 3550 8930
rect 3650 9010 3750 9020
rect 3650 8930 3660 9010
rect 3740 8930 3750 9010
rect 3650 8920 3750 8930
rect 3850 9010 3950 9020
rect 3850 8930 3860 9010
rect 3940 8930 3950 9010
rect 3850 8920 3950 8930
rect 4050 9010 4150 9020
rect 4050 8930 4060 9010
rect 4140 8930 4150 9010
rect 4050 8920 4150 8930
rect 4250 9010 4350 9020
rect 4250 8930 4260 9010
rect 4340 8930 4350 9010
rect 4250 8920 4350 8930
rect 4450 9010 4550 9020
rect 4450 8930 4460 9010
rect 4540 8930 4550 9010
rect 4450 8920 4550 8930
rect 4650 9010 4750 9020
rect 4650 8930 4660 9010
rect 4740 8930 4750 9010
rect 4650 8920 4750 8930
rect 4850 9010 4950 9020
rect 4850 8930 4860 9010
rect 4940 8930 4950 9010
rect 4850 8920 4950 8930
rect 5050 9010 5150 9020
rect 5050 8930 5060 9010
rect 5140 8930 5150 9010
rect 5050 8920 5150 8930
rect 5250 9010 5350 9020
rect 5250 8930 5260 9010
rect 5340 8930 5350 9010
rect 5250 8920 5350 8930
rect 5450 9010 5550 9020
rect 5450 8930 5460 9010
rect 5540 8930 5550 9010
rect 5450 8920 5550 8930
rect 5650 9010 5750 9020
rect 5650 8930 5660 9010
rect 5740 8930 5750 9010
rect 5650 8920 5750 8930
rect 5850 9010 5950 9020
rect 5850 8930 5860 9010
rect 5940 8930 5950 9010
rect 5850 8920 5950 8930
rect 6050 9010 6150 9020
rect 6050 8930 6060 9010
rect 6140 8930 6150 9010
rect 6050 8920 6150 8930
rect 6250 9010 6350 9020
rect 6250 8930 6260 9010
rect 6340 8930 6350 9010
rect 6250 8920 6350 8930
rect 6450 9010 6550 9020
rect 6450 8930 6460 9010
rect 6540 8930 6550 9010
rect 6450 8920 6550 8930
rect -150 8825 -50 8835
rect -150 8745 -140 8825
rect -60 8745 -50 8825
rect -150 8735 -50 8745
rect 50 8825 150 8835
rect 50 8745 60 8825
rect 140 8745 150 8825
rect 50 8735 150 8745
rect 250 8825 350 8835
rect 250 8745 260 8825
rect 340 8745 350 8825
rect 250 8735 350 8745
rect 450 8825 550 8835
rect 450 8745 460 8825
rect 540 8745 550 8825
rect 450 8735 550 8745
rect 650 8825 750 8835
rect 650 8745 660 8825
rect 740 8745 750 8825
rect 650 8735 750 8745
rect 850 8825 950 8835
rect 850 8745 860 8825
rect 940 8745 950 8825
rect 850 8735 950 8745
rect 1050 8825 1150 8835
rect 1050 8745 1060 8825
rect 1140 8745 1150 8825
rect 1050 8735 1150 8745
rect 1250 8825 1350 8835
rect 1250 8745 1260 8825
rect 1340 8745 1350 8825
rect 1250 8735 1350 8745
rect 1450 8825 1550 8835
rect 1450 8745 1460 8825
rect 1540 8745 1550 8825
rect 1450 8735 1550 8745
rect 1650 8825 1750 8835
rect 1650 8745 1660 8825
rect 1740 8745 1750 8825
rect 1650 8735 1750 8745
rect 1850 8825 1950 8835
rect 1850 8745 1860 8825
rect 1940 8745 1950 8825
rect 1850 8735 1950 8745
rect 2050 8825 2150 8835
rect 2050 8745 2060 8825
rect 2140 8745 2150 8825
rect 2050 8735 2150 8745
rect 2250 8825 2350 8835
rect 2250 8745 2260 8825
rect 2340 8745 2350 8825
rect 2250 8735 2350 8745
rect 2450 8825 2550 8835
rect 2450 8745 2460 8825
rect 2540 8745 2550 8825
rect 2450 8735 2550 8745
rect 2650 8825 2750 8835
rect 2650 8745 2660 8825
rect 2740 8745 2750 8825
rect 2650 8735 2750 8745
rect 2850 8825 2950 8835
rect 2850 8745 2860 8825
rect 2940 8745 2950 8825
rect 2850 8735 2950 8745
rect 3050 8825 3150 8835
rect 3050 8745 3060 8825
rect 3140 8745 3150 8825
rect 3050 8735 3150 8745
rect 3250 8825 3350 8835
rect 3250 8745 3260 8825
rect 3340 8745 3350 8825
rect 3250 8735 3350 8745
rect 3450 8825 3550 8835
rect 3450 8745 3460 8825
rect 3540 8745 3550 8825
rect 3450 8735 3550 8745
rect 3650 8825 3750 8835
rect 3650 8745 3660 8825
rect 3740 8745 3750 8825
rect 3650 8735 3750 8745
rect 3850 8825 3950 8835
rect 3850 8745 3860 8825
rect 3940 8745 3950 8825
rect 3850 8735 3950 8745
rect 4050 8825 4150 8835
rect 4050 8745 4060 8825
rect 4140 8745 4150 8825
rect 4050 8735 4150 8745
rect 4250 8825 4350 8835
rect 4250 8745 4260 8825
rect 4340 8745 4350 8825
rect 4250 8735 4350 8745
rect 4450 8825 4550 8835
rect 4450 8745 4460 8825
rect 4540 8745 4550 8825
rect 4450 8735 4550 8745
rect 4650 8825 4750 8835
rect 4650 8745 4660 8825
rect 4740 8745 4750 8825
rect 4650 8735 4750 8745
rect 4850 8825 4950 8835
rect 4850 8745 4860 8825
rect 4940 8745 4950 8825
rect 4850 8735 4950 8745
rect 5050 8825 5150 8835
rect 5050 8745 5060 8825
rect 5140 8745 5150 8825
rect 5050 8735 5150 8745
rect 5250 8825 5350 8835
rect 5250 8745 5260 8825
rect 5340 8745 5350 8825
rect 5250 8735 5350 8745
rect 5450 8825 5550 8835
rect 5450 8745 5460 8825
rect 5540 8745 5550 8825
rect 5450 8735 5550 8745
rect 5650 8825 5750 8835
rect 5650 8745 5660 8825
rect 5740 8745 5750 8825
rect 5650 8735 5750 8745
rect 5850 8825 5950 8835
rect 5850 8745 5860 8825
rect 5940 8745 5950 8825
rect 5850 8735 5950 8745
rect 6050 8825 6150 8835
rect 6050 8745 6060 8825
rect 6140 8745 6150 8825
rect 6050 8735 6150 8745
rect 6250 8825 6350 8835
rect 6250 8745 6260 8825
rect 6340 8745 6350 8825
rect 6250 8735 6350 8745
rect 6450 8825 6550 8835
rect 6450 8745 6460 8825
rect 6540 8745 6550 8825
rect 6450 8735 6550 8745
rect -150 8640 -50 8650
rect -150 8560 -140 8640
rect -60 8560 -50 8640
rect -150 8550 -50 8560
rect 50 8640 150 8650
rect 50 8560 60 8640
rect 140 8560 150 8640
rect 50 8550 150 8560
rect 250 8640 350 8650
rect 250 8560 260 8640
rect 340 8560 350 8640
rect 250 8550 350 8560
rect 450 8640 550 8650
rect 450 8560 460 8640
rect 540 8560 550 8640
rect 450 8550 550 8560
rect 650 8640 750 8650
rect 650 8560 660 8640
rect 740 8560 750 8640
rect 650 8550 750 8560
rect 850 8640 950 8650
rect 850 8560 860 8640
rect 940 8560 950 8640
rect 850 8550 950 8560
rect 1050 8640 1150 8650
rect 1050 8560 1060 8640
rect 1140 8560 1150 8640
rect 1050 8550 1150 8560
rect 1250 8640 1350 8650
rect 1250 8560 1260 8640
rect 1340 8560 1350 8640
rect 1250 8550 1350 8560
rect 1450 8640 1550 8650
rect 1450 8560 1460 8640
rect 1540 8560 1550 8640
rect 1450 8550 1550 8560
rect 1650 8640 1750 8650
rect 1650 8560 1660 8640
rect 1740 8560 1750 8640
rect 1650 8550 1750 8560
rect 1850 8640 1950 8650
rect 1850 8560 1860 8640
rect 1940 8560 1950 8640
rect 1850 8550 1950 8560
rect 2050 8640 2150 8650
rect 2050 8560 2060 8640
rect 2140 8560 2150 8640
rect 2050 8550 2150 8560
rect 2250 8640 2350 8650
rect 2250 8560 2260 8640
rect 2340 8560 2350 8640
rect 2250 8550 2350 8560
rect 2450 8640 2550 8650
rect 2450 8560 2460 8640
rect 2540 8560 2550 8640
rect 2450 8550 2550 8560
rect 2650 8640 2750 8650
rect 2650 8560 2660 8640
rect 2740 8560 2750 8640
rect 2650 8550 2750 8560
rect 2850 8640 2950 8650
rect 2850 8560 2860 8640
rect 2940 8560 2950 8640
rect 2850 8550 2950 8560
rect 3050 8640 3150 8650
rect 3050 8560 3060 8640
rect 3140 8560 3150 8640
rect 3050 8550 3150 8560
rect 3250 8640 3350 8650
rect 3250 8560 3260 8640
rect 3340 8560 3350 8640
rect 3250 8550 3350 8560
rect 3450 8640 3550 8650
rect 3450 8560 3460 8640
rect 3540 8560 3550 8640
rect 3450 8550 3550 8560
rect 3650 8640 3750 8650
rect 3650 8560 3660 8640
rect 3740 8560 3750 8640
rect 3650 8550 3750 8560
rect 3850 8640 3950 8650
rect 3850 8560 3860 8640
rect 3940 8560 3950 8640
rect 3850 8550 3950 8560
rect 4050 8640 4150 8650
rect 4050 8560 4060 8640
rect 4140 8560 4150 8640
rect 4050 8550 4150 8560
rect 4250 8640 4350 8650
rect 4250 8560 4260 8640
rect 4340 8560 4350 8640
rect 4250 8550 4350 8560
rect 4450 8640 4550 8650
rect 4450 8560 4460 8640
rect 4540 8560 4550 8640
rect 4450 8550 4550 8560
rect 4650 8640 4750 8650
rect 4650 8560 4660 8640
rect 4740 8560 4750 8640
rect 4650 8550 4750 8560
rect 4850 8640 4950 8650
rect 4850 8560 4860 8640
rect 4940 8560 4950 8640
rect 4850 8550 4950 8560
rect 5050 8640 5150 8650
rect 5050 8560 5060 8640
rect 5140 8560 5150 8640
rect 5050 8550 5150 8560
rect 5250 8640 5350 8650
rect 5250 8560 5260 8640
rect 5340 8560 5350 8640
rect 5250 8550 5350 8560
rect 5450 8640 5550 8650
rect 5450 8560 5460 8640
rect 5540 8560 5550 8640
rect 5450 8550 5550 8560
rect 5650 8640 5750 8650
rect 5650 8560 5660 8640
rect 5740 8560 5750 8640
rect 5650 8550 5750 8560
rect 5850 8640 5950 8650
rect 5850 8560 5860 8640
rect 5940 8560 5950 8640
rect 5850 8550 5950 8560
rect 6050 8640 6150 8650
rect 6050 8560 6060 8640
rect 6140 8560 6150 8640
rect 6050 8550 6150 8560
rect 6250 8640 6350 8650
rect 6250 8560 6260 8640
rect 6340 8560 6350 8640
rect 6250 8550 6350 8560
rect 6450 8640 6550 8650
rect 6450 8560 6460 8640
rect 6540 8560 6550 8640
rect 6450 8550 6550 8560
rect -150 8455 -50 8465
rect -150 8375 -140 8455
rect -60 8375 -50 8455
rect -150 8365 -50 8375
rect 50 8455 150 8465
rect 50 8375 60 8455
rect 140 8375 150 8455
rect 50 8365 150 8375
rect 250 8455 350 8465
rect 250 8375 260 8455
rect 340 8375 350 8455
rect 250 8365 350 8375
rect 450 8455 550 8465
rect 450 8375 460 8455
rect 540 8375 550 8455
rect 450 8365 550 8375
rect 650 8455 750 8465
rect 650 8375 660 8455
rect 740 8375 750 8455
rect 650 8365 750 8375
rect 850 8455 950 8465
rect 850 8375 860 8455
rect 940 8375 950 8455
rect 850 8365 950 8375
rect 1050 8455 1150 8465
rect 1050 8375 1060 8455
rect 1140 8375 1150 8455
rect 1050 8365 1150 8375
rect 1250 8455 1350 8465
rect 1250 8375 1260 8455
rect 1340 8375 1350 8455
rect 1250 8365 1350 8375
rect 1450 8455 1550 8465
rect 1450 8375 1460 8455
rect 1540 8375 1550 8455
rect 1450 8365 1550 8375
rect 1650 8455 1750 8465
rect 1650 8375 1660 8455
rect 1740 8375 1750 8455
rect 1650 8365 1750 8375
rect 1850 8455 1950 8465
rect 1850 8375 1860 8455
rect 1940 8375 1950 8455
rect 1850 8365 1950 8375
rect 2050 8455 2150 8465
rect 2050 8375 2060 8455
rect 2140 8375 2150 8455
rect 2050 8365 2150 8375
rect 2250 8455 2350 8465
rect 2250 8375 2260 8455
rect 2340 8375 2350 8455
rect 2250 8365 2350 8375
rect 2450 8455 2550 8465
rect 2450 8375 2460 8455
rect 2540 8375 2550 8455
rect 2450 8365 2550 8375
rect 2650 8455 2750 8465
rect 2650 8375 2660 8455
rect 2740 8375 2750 8455
rect 2650 8365 2750 8375
rect 2850 8455 2950 8465
rect 2850 8375 2860 8455
rect 2940 8375 2950 8455
rect 2850 8365 2950 8375
rect 3050 8455 3150 8465
rect 3050 8375 3060 8455
rect 3140 8375 3150 8455
rect 3050 8365 3150 8375
rect 3250 8455 3350 8465
rect 3250 8375 3260 8455
rect 3340 8375 3350 8455
rect 3250 8365 3350 8375
rect 3450 8455 3550 8465
rect 3450 8375 3460 8455
rect 3540 8375 3550 8455
rect 3450 8365 3550 8375
rect 3650 8455 3750 8465
rect 3650 8375 3660 8455
rect 3740 8375 3750 8455
rect 3650 8365 3750 8375
rect 3850 8455 3950 8465
rect 3850 8375 3860 8455
rect 3940 8375 3950 8455
rect 3850 8365 3950 8375
rect 4050 8455 4150 8465
rect 4050 8375 4060 8455
rect 4140 8375 4150 8455
rect 4050 8365 4150 8375
rect 4250 8455 4350 8465
rect 4250 8375 4260 8455
rect 4340 8375 4350 8455
rect 4250 8365 4350 8375
rect 4450 8455 4550 8465
rect 4450 8375 4460 8455
rect 4540 8375 4550 8455
rect 4450 8365 4550 8375
rect 4650 8455 4750 8465
rect 4650 8375 4660 8455
rect 4740 8375 4750 8455
rect 4650 8365 4750 8375
rect 4850 8455 4950 8465
rect 4850 8375 4860 8455
rect 4940 8375 4950 8455
rect 4850 8365 4950 8375
rect 5050 8455 5150 8465
rect 5050 8375 5060 8455
rect 5140 8375 5150 8455
rect 5050 8365 5150 8375
rect 5250 8455 5350 8465
rect 5250 8375 5260 8455
rect 5340 8375 5350 8455
rect 5250 8365 5350 8375
rect 5450 8455 5550 8465
rect 5450 8375 5460 8455
rect 5540 8375 5550 8455
rect 5450 8365 5550 8375
rect 5650 8455 5750 8465
rect 5650 8375 5660 8455
rect 5740 8375 5750 8455
rect 5650 8365 5750 8375
rect 5850 8455 5950 8465
rect 5850 8375 5860 8455
rect 5940 8375 5950 8455
rect 5850 8365 5950 8375
rect 6050 8455 6150 8465
rect 6050 8375 6060 8455
rect 6140 8375 6150 8455
rect 6050 8365 6150 8375
rect 6250 8455 6350 8465
rect 6250 8375 6260 8455
rect 6340 8375 6350 8455
rect 6250 8365 6350 8375
rect 6450 8455 6550 8465
rect 6450 8375 6460 8455
rect 6540 8375 6550 8455
rect 6450 8365 6550 8375
rect -150 8270 -50 8280
rect -150 8190 -140 8270
rect -60 8190 -50 8270
rect -150 8180 -50 8190
rect 50 8270 150 8280
rect 50 8190 60 8270
rect 140 8190 150 8270
rect 50 8180 150 8190
rect 250 8270 350 8280
rect 250 8190 260 8270
rect 340 8190 350 8270
rect 250 8180 350 8190
rect 450 8270 550 8280
rect 450 8190 460 8270
rect 540 8190 550 8270
rect 450 8180 550 8190
rect 650 8270 750 8280
rect 650 8190 660 8270
rect 740 8190 750 8270
rect 650 8180 750 8190
rect 850 8270 950 8280
rect 850 8190 860 8270
rect 940 8190 950 8270
rect 850 8180 950 8190
rect 1050 8270 1150 8280
rect 1050 8190 1060 8270
rect 1140 8190 1150 8270
rect 1050 8180 1150 8190
rect 1250 8270 1350 8280
rect 1250 8190 1260 8270
rect 1340 8190 1350 8270
rect 1250 8180 1350 8190
rect 1450 8270 1550 8280
rect 1450 8190 1460 8270
rect 1540 8190 1550 8270
rect 1450 8180 1550 8190
rect 1650 8270 1750 8280
rect 1650 8190 1660 8270
rect 1740 8190 1750 8270
rect 1650 8180 1750 8190
rect 1850 8270 1950 8280
rect 1850 8190 1860 8270
rect 1940 8190 1950 8270
rect 1850 8180 1950 8190
rect 2050 8270 2150 8280
rect 2050 8190 2060 8270
rect 2140 8190 2150 8270
rect 2050 8180 2150 8190
rect 2250 8270 2350 8280
rect 2250 8190 2260 8270
rect 2340 8190 2350 8270
rect 2250 8180 2350 8190
rect 2450 8270 2550 8280
rect 2450 8190 2460 8270
rect 2540 8190 2550 8270
rect 2450 8180 2550 8190
rect 2650 8270 2750 8280
rect 2650 8190 2660 8270
rect 2740 8190 2750 8270
rect 2650 8180 2750 8190
rect 2850 8270 2950 8280
rect 2850 8190 2860 8270
rect 2940 8190 2950 8270
rect 2850 8180 2950 8190
rect 3050 8270 3150 8280
rect 3050 8190 3060 8270
rect 3140 8190 3150 8270
rect 3050 8180 3150 8190
rect 3250 8270 3350 8280
rect 3250 8190 3260 8270
rect 3340 8190 3350 8270
rect 3250 8180 3350 8190
rect 3450 8270 3550 8280
rect 3450 8190 3460 8270
rect 3540 8190 3550 8270
rect 3450 8180 3550 8190
rect 3650 8270 3750 8280
rect 3650 8190 3660 8270
rect 3740 8190 3750 8270
rect 3650 8180 3750 8190
rect 3850 8270 3950 8280
rect 3850 8190 3860 8270
rect 3940 8190 3950 8270
rect 3850 8180 3950 8190
rect 4050 8270 4150 8280
rect 4050 8190 4060 8270
rect 4140 8190 4150 8270
rect 4050 8180 4150 8190
rect 4250 8270 4350 8280
rect 4250 8190 4260 8270
rect 4340 8190 4350 8270
rect 4250 8180 4350 8190
rect 4450 8270 4550 8280
rect 4450 8190 4460 8270
rect 4540 8190 4550 8270
rect 4450 8180 4550 8190
rect 4650 8270 4750 8280
rect 4650 8190 4660 8270
rect 4740 8190 4750 8270
rect 4650 8180 4750 8190
rect 4850 8270 4950 8280
rect 4850 8190 4860 8270
rect 4940 8190 4950 8270
rect 4850 8180 4950 8190
rect 5050 8270 5150 8280
rect 5050 8190 5060 8270
rect 5140 8190 5150 8270
rect 5050 8180 5150 8190
rect 5250 8270 5350 8280
rect 5250 8190 5260 8270
rect 5340 8190 5350 8270
rect 5250 8180 5350 8190
rect 5450 8270 5550 8280
rect 5450 8190 5460 8270
rect 5540 8190 5550 8270
rect 5450 8180 5550 8190
rect 5650 8270 5750 8280
rect 5650 8190 5660 8270
rect 5740 8190 5750 8270
rect 5650 8180 5750 8190
rect 5850 8270 5950 8280
rect 5850 8190 5860 8270
rect 5940 8190 5950 8270
rect 5850 8180 5950 8190
rect 6050 8270 6150 8280
rect 6050 8190 6060 8270
rect 6140 8190 6150 8270
rect 6050 8180 6150 8190
rect 6250 8270 6350 8280
rect 6250 8190 6260 8270
rect 6340 8190 6350 8270
rect 6250 8180 6350 8190
rect 6450 8270 6550 8280
rect 6450 8190 6460 8270
rect 6540 8190 6550 8270
rect 6450 8180 6550 8190
rect -150 8085 -50 8095
rect -150 8005 -140 8085
rect -60 8005 -50 8085
rect -150 7995 -50 8005
rect 50 8085 150 8095
rect 50 8005 60 8085
rect 140 8005 150 8085
rect 50 7995 150 8005
rect 250 8085 350 8095
rect 250 8005 260 8085
rect 340 8005 350 8085
rect 250 7995 350 8005
rect 450 8085 550 8095
rect 450 8005 460 8085
rect 540 8005 550 8085
rect 450 7995 550 8005
rect 650 8085 750 8095
rect 650 8005 660 8085
rect 740 8005 750 8085
rect 650 7995 750 8005
rect 850 8085 950 8095
rect 850 8005 860 8085
rect 940 8005 950 8085
rect 850 7995 950 8005
rect 1050 8085 1150 8095
rect 1050 8005 1060 8085
rect 1140 8005 1150 8085
rect 1050 7995 1150 8005
rect 1250 8085 1350 8095
rect 1250 8005 1260 8085
rect 1340 8005 1350 8085
rect 1250 7995 1350 8005
rect 1450 8085 1550 8095
rect 1450 8005 1460 8085
rect 1540 8005 1550 8085
rect 1450 7995 1550 8005
rect 1650 8085 1750 8095
rect 1650 8005 1660 8085
rect 1740 8005 1750 8085
rect 1650 7995 1750 8005
rect 1850 8085 1950 8095
rect 1850 8005 1860 8085
rect 1940 8005 1950 8085
rect 1850 7995 1950 8005
rect 2050 8085 2150 8095
rect 2050 8005 2060 8085
rect 2140 8005 2150 8085
rect 2050 7995 2150 8005
rect 2250 8085 2350 8095
rect 2250 8005 2260 8085
rect 2340 8005 2350 8085
rect 2250 7995 2350 8005
rect 2450 8085 2550 8095
rect 2450 8005 2460 8085
rect 2540 8005 2550 8085
rect 2450 7995 2550 8005
rect 2650 8085 2750 8095
rect 2650 8005 2660 8085
rect 2740 8005 2750 8085
rect 2650 7995 2750 8005
rect 2850 8085 2950 8095
rect 2850 8005 2860 8085
rect 2940 8005 2950 8085
rect 2850 7995 2950 8005
rect 3050 8085 3150 8095
rect 3050 8005 3060 8085
rect 3140 8005 3150 8085
rect 3050 7995 3150 8005
rect 3250 8085 3350 8095
rect 3250 8005 3260 8085
rect 3340 8005 3350 8085
rect 3250 7995 3350 8005
rect 3450 8085 3550 8095
rect 3450 8005 3460 8085
rect 3540 8005 3550 8085
rect 3450 7995 3550 8005
rect 3650 8085 3750 8095
rect 3650 8005 3660 8085
rect 3740 8005 3750 8085
rect 3650 7995 3750 8005
rect 3850 8085 3950 8095
rect 3850 8005 3860 8085
rect 3940 8005 3950 8085
rect 3850 7995 3950 8005
rect 4050 8085 4150 8095
rect 4050 8005 4060 8085
rect 4140 8005 4150 8085
rect 4050 7995 4150 8005
rect 4250 8085 4350 8095
rect 4250 8005 4260 8085
rect 4340 8005 4350 8085
rect 4250 7995 4350 8005
rect 4450 8085 4550 8095
rect 4450 8005 4460 8085
rect 4540 8005 4550 8085
rect 4450 7995 4550 8005
rect 4650 8085 4750 8095
rect 4650 8005 4660 8085
rect 4740 8005 4750 8085
rect 4650 7995 4750 8005
rect 4850 8085 4950 8095
rect 4850 8005 4860 8085
rect 4940 8005 4950 8085
rect 4850 7995 4950 8005
rect 5050 8085 5150 8095
rect 5050 8005 5060 8085
rect 5140 8005 5150 8085
rect 5050 7995 5150 8005
rect 5250 8085 5350 8095
rect 5250 8005 5260 8085
rect 5340 8005 5350 8085
rect 5250 7995 5350 8005
rect 5450 8085 5550 8095
rect 5450 8005 5460 8085
rect 5540 8005 5550 8085
rect 5450 7995 5550 8005
rect 5650 8085 5750 8095
rect 5650 8005 5660 8085
rect 5740 8005 5750 8085
rect 5650 7995 5750 8005
rect 5850 8085 5950 8095
rect 5850 8005 5860 8085
rect 5940 8005 5950 8085
rect 5850 7995 5950 8005
rect 6050 8085 6150 8095
rect 6050 8005 6060 8085
rect 6140 8005 6150 8085
rect 6050 7995 6150 8005
rect 6250 8085 6350 8095
rect 6250 8005 6260 8085
rect 6340 8005 6350 8085
rect 6250 7995 6350 8005
rect 6450 8085 6550 8095
rect 6450 8005 6460 8085
rect 6540 8005 6550 8085
rect 6450 7995 6550 8005
rect -150 7900 -50 7910
rect -150 7820 -140 7900
rect -60 7820 -50 7900
rect -150 7810 -50 7820
rect 50 7900 150 7910
rect 50 7820 60 7900
rect 140 7820 150 7900
rect 50 7810 150 7820
rect 250 7900 350 7910
rect 250 7820 260 7900
rect 340 7820 350 7900
rect 250 7810 350 7820
rect 450 7900 550 7910
rect 450 7820 460 7900
rect 540 7820 550 7900
rect 450 7810 550 7820
rect 650 7900 750 7910
rect 650 7820 660 7900
rect 740 7820 750 7900
rect 650 7810 750 7820
rect 850 7900 950 7910
rect 850 7820 860 7900
rect 940 7820 950 7900
rect 850 7810 950 7820
rect 1050 7900 1150 7910
rect 1050 7820 1060 7900
rect 1140 7820 1150 7900
rect 1050 7810 1150 7820
rect 1250 7900 1350 7910
rect 1250 7820 1260 7900
rect 1340 7820 1350 7900
rect 1250 7810 1350 7820
rect 1450 7900 1550 7910
rect 1450 7820 1460 7900
rect 1540 7820 1550 7900
rect 1450 7810 1550 7820
rect 1650 7900 1750 7910
rect 1650 7820 1660 7900
rect 1740 7820 1750 7900
rect 1650 7810 1750 7820
rect 1850 7900 1950 7910
rect 1850 7820 1860 7900
rect 1940 7820 1950 7900
rect 1850 7810 1950 7820
rect 2050 7900 2150 7910
rect 2050 7820 2060 7900
rect 2140 7820 2150 7900
rect 2050 7810 2150 7820
rect 2250 7900 2350 7910
rect 2250 7820 2260 7900
rect 2340 7820 2350 7900
rect 2250 7810 2350 7820
rect 2450 7900 2550 7910
rect 2450 7820 2460 7900
rect 2540 7820 2550 7900
rect 2450 7810 2550 7820
rect 2650 7900 2750 7910
rect 2650 7820 2660 7900
rect 2740 7820 2750 7900
rect 2650 7810 2750 7820
rect 2850 7900 2950 7910
rect 2850 7820 2860 7900
rect 2940 7820 2950 7900
rect 2850 7810 2950 7820
rect 3050 7900 3150 7910
rect 3050 7820 3060 7900
rect 3140 7820 3150 7900
rect 3050 7810 3150 7820
rect 3250 7900 3350 7910
rect 3250 7820 3260 7900
rect 3340 7820 3350 7900
rect 3250 7810 3350 7820
rect 3450 7900 3550 7910
rect 3450 7820 3460 7900
rect 3540 7820 3550 7900
rect 3450 7810 3550 7820
rect 3650 7900 3750 7910
rect 3650 7820 3660 7900
rect 3740 7820 3750 7900
rect 3650 7810 3750 7820
rect 3850 7900 3950 7910
rect 3850 7820 3860 7900
rect 3940 7820 3950 7900
rect 3850 7810 3950 7820
rect 4050 7900 4150 7910
rect 4050 7820 4060 7900
rect 4140 7820 4150 7900
rect 4050 7810 4150 7820
rect 4250 7900 4350 7910
rect 4250 7820 4260 7900
rect 4340 7820 4350 7900
rect 4250 7810 4350 7820
rect 4450 7900 4550 7910
rect 4450 7820 4460 7900
rect 4540 7820 4550 7900
rect 4450 7810 4550 7820
rect 4650 7900 4750 7910
rect 4650 7820 4660 7900
rect 4740 7820 4750 7900
rect 4650 7810 4750 7820
rect 4850 7900 4950 7910
rect 4850 7820 4860 7900
rect 4940 7820 4950 7900
rect 4850 7810 4950 7820
rect 5050 7900 5150 7910
rect 5050 7820 5060 7900
rect 5140 7820 5150 7900
rect 5050 7810 5150 7820
rect 5250 7900 5350 7910
rect 5250 7820 5260 7900
rect 5340 7820 5350 7900
rect 5250 7810 5350 7820
rect 5450 7900 5550 7910
rect 5450 7820 5460 7900
rect 5540 7820 5550 7900
rect 5450 7810 5550 7820
rect 5650 7900 5750 7910
rect 5650 7820 5660 7900
rect 5740 7820 5750 7900
rect 5650 7810 5750 7820
rect 5850 7900 5950 7910
rect 5850 7820 5860 7900
rect 5940 7820 5950 7900
rect 5850 7810 5950 7820
rect 6050 7900 6150 7910
rect 6050 7820 6060 7900
rect 6140 7820 6150 7900
rect 6050 7810 6150 7820
rect 6250 7900 6350 7910
rect 6250 7820 6260 7900
rect 6340 7820 6350 7900
rect 6250 7810 6350 7820
rect 6450 7900 6550 7910
rect 6450 7820 6460 7900
rect 6540 7820 6550 7900
rect 6450 7810 6550 7820
rect -150 7715 -50 7725
rect -150 7635 -140 7715
rect -60 7635 -50 7715
rect -150 7625 -50 7635
rect 50 7715 150 7725
rect 50 7635 60 7715
rect 140 7635 150 7715
rect 50 7625 150 7635
rect 250 7715 350 7725
rect 250 7635 260 7715
rect 340 7635 350 7715
rect 250 7625 350 7635
rect 450 7715 550 7725
rect 450 7635 460 7715
rect 540 7635 550 7715
rect 450 7625 550 7635
rect 650 7715 750 7725
rect 650 7635 660 7715
rect 740 7635 750 7715
rect 650 7625 750 7635
rect 850 7715 950 7725
rect 850 7635 860 7715
rect 940 7635 950 7715
rect 850 7625 950 7635
rect 1050 7715 1150 7725
rect 1050 7635 1060 7715
rect 1140 7635 1150 7715
rect 1050 7625 1150 7635
rect 1250 7715 1350 7725
rect 1250 7635 1260 7715
rect 1340 7635 1350 7715
rect 1250 7625 1350 7635
rect 1450 7715 1550 7725
rect 1450 7635 1460 7715
rect 1540 7635 1550 7715
rect 1450 7625 1550 7635
rect 1650 7715 1750 7725
rect 1650 7635 1660 7715
rect 1740 7635 1750 7715
rect 1650 7625 1750 7635
rect 1850 7715 1950 7725
rect 1850 7635 1860 7715
rect 1940 7635 1950 7715
rect 1850 7625 1950 7635
rect 2050 7715 2150 7725
rect 2050 7635 2060 7715
rect 2140 7635 2150 7715
rect 2050 7625 2150 7635
rect 2250 7715 2350 7725
rect 2250 7635 2260 7715
rect 2340 7635 2350 7715
rect 2250 7625 2350 7635
rect 2450 7715 2550 7725
rect 2450 7635 2460 7715
rect 2540 7635 2550 7715
rect 2450 7625 2550 7635
rect 2650 7715 2750 7725
rect 2650 7635 2660 7715
rect 2740 7635 2750 7715
rect 2650 7625 2750 7635
rect 2850 7715 2950 7725
rect 2850 7635 2860 7715
rect 2940 7635 2950 7715
rect 2850 7625 2950 7635
rect 3050 7715 3150 7725
rect 3050 7635 3060 7715
rect 3140 7635 3150 7715
rect 3050 7625 3150 7635
rect 3250 7715 3350 7725
rect 3250 7635 3260 7715
rect 3340 7635 3350 7715
rect 3250 7625 3350 7635
rect 3450 7715 3550 7725
rect 3450 7635 3460 7715
rect 3540 7635 3550 7715
rect 3450 7625 3550 7635
rect 3650 7715 3750 7725
rect 3650 7635 3660 7715
rect 3740 7635 3750 7715
rect 3650 7625 3750 7635
rect 3850 7715 3950 7725
rect 3850 7635 3860 7715
rect 3940 7635 3950 7715
rect 3850 7625 3950 7635
rect 4050 7715 4150 7725
rect 4050 7635 4060 7715
rect 4140 7635 4150 7715
rect 4050 7625 4150 7635
rect 4250 7715 4350 7725
rect 4250 7635 4260 7715
rect 4340 7635 4350 7715
rect 4250 7625 4350 7635
rect 4450 7715 4550 7725
rect 4450 7635 4460 7715
rect 4540 7635 4550 7715
rect 4450 7625 4550 7635
rect 4650 7715 4750 7725
rect 4650 7635 4660 7715
rect 4740 7635 4750 7715
rect 4650 7625 4750 7635
rect 4850 7715 4950 7725
rect 4850 7635 4860 7715
rect 4940 7635 4950 7715
rect 4850 7625 4950 7635
rect 5050 7715 5150 7725
rect 5050 7635 5060 7715
rect 5140 7635 5150 7715
rect 5050 7625 5150 7635
rect 5250 7715 5350 7725
rect 5250 7635 5260 7715
rect 5340 7635 5350 7715
rect 5250 7625 5350 7635
rect 5450 7715 5550 7725
rect 5450 7635 5460 7715
rect 5540 7635 5550 7715
rect 5450 7625 5550 7635
rect 5650 7715 5750 7725
rect 5650 7635 5660 7715
rect 5740 7635 5750 7715
rect 5650 7625 5750 7635
rect 5850 7715 5950 7725
rect 5850 7635 5860 7715
rect 5940 7635 5950 7715
rect 5850 7625 5950 7635
rect 6050 7715 6150 7725
rect 6050 7635 6060 7715
rect 6140 7635 6150 7715
rect 6050 7625 6150 7635
rect 6250 7715 6350 7725
rect 6250 7635 6260 7715
rect 6340 7635 6350 7715
rect 6250 7625 6350 7635
rect 6450 7715 6550 7725
rect 6450 7635 6460 7715
rect 6540 7635 6550 7715
rect 6450 7625 6550 7635
rect -150 7530 -50 7540
rect -150 7450 -140 7530
rect -60 7450 -50 7530
rect -150 7440 -50 7450
rect 50 7530 150 7540
rect 50 7450 60 7530
rect 140 7450 150 7530
rect 50 7440 150 7450
rect 250 7530 350 7540
rect 250 7450 260 7530
rect 340 7450 350 7530
rect 250 7440 350 7450
rect 450 7530 550 7540
rect 450 7450 460 7530
rect 540 7450 550 7530
rect 450 7440 550 7450
rect 650 7530 750 7540
rect 650 7450 660 7530
rect 740 7450 750 7530
rect 650 7440 750 7450
rect 850 7530 950 7540
rect 850 7450 860 7530
rect 940 7450 950 7530
rect 850 7440 950 7450
rect 1050 7530 1150 7540
rect 1050 7450 1060 7530
rect 1140 7450 1150 7530
rect 1050 7440 1150 7450
rect 1250 7530 1350 7540
rect 1250 7450 1260 7530
rect 1340 7450 1350 7530
rect 1250 7440 1350 7450
rect 1450 7530 1550 7540
rect 1450 7450 1460 7530
rect 1540 7450 1550 7530
rect 1450 7440 1550 7450
rect 1650 7530 1750 7540
rect 1650 7450 1660 7530
rect 1740 7450 1750 7530
rect 1650 7440 1750 7450
rect 1850 7530 1950 7540
rect 1850 7450 1860 7530
rect 1940 7450 1950 7530
rect 1850 7440 1950 7450
rect 2050 7530 2150 7540
rect 2050 7450 2060 7530
rect 2140 7450 2150 7530
rect 2050 7440 2150 7450
rect 2250 7530 2350 7540
rect 2250 7450 2260 7530
rect 2340 7450 2350 7530
rect 2250 7440 2350 7450
rect 2450 7530 2550 7540
rect 2450 7450 2460 7530
rect 2540 7450 2550 7530
rect 2450 7440 2550 7450
rect 2650 7530 2750 7540
rect 2650 7450 2660 7530
rect 2740 7450 2750 7530
rect 2650 7440 2750 7450
rect 2850 7530 2950 7540
rect 2850 7450 2860 7530
rect 2940 7450 2950 7530
rect 2850 7440 2950 7450
rect 3050 7530 3150 7540
rect 3050 7450 3060 7530
rect 3140 7450 3150 7530
rect 3050 7440 3150 7450
rect 3250 7530 3350 7540
rect 3250 7450 3260 7530
rect 3340 7450 3350 7530
rect 3250 7440 3350 7450
rect 3450 7530 3550 7540
rect 3450 7450 3460 7530
rect 3540 7450 3550 7530
rect 3450 7440 3550 7450
rect 3650 7530 3750 7540
rect 3650 7450 3660 7530
rect 3740 7450 3750 7530
rect 3650 7440 3750 7450
rect 3850 7530 3950 7540
rect 3850 7450 3860 7530
rect 3940 7450 3950 7530
rect 3850 7440 3950 7450
rect 4050 7530 4150 7540
rect 4050 7450 4060 7530
rect 4140 7450 4150 7530
rect 4050 7440 4150 7450
rect 4250 7530 4350 7540
rect 4250 7450 4260 7530
rect 4340 7450 4350 7530
rect 4250 7440 4350 7450
rect 4450 7530 4550 7540
rect 4450 7450 4460 7530
rect 4540 7450 4550 7530
rect 4450 7440 4550 7450
rect 4650 7530 4750 7540
rect 4650 7450 4660 7530
rect 4740 7450 4750 7530
rect 4650 7440 4750 7450
rect 4850 7530 4950 7540
rect 4850 7450 4860 7530
rect 4940 7450 4950 7530
rect 4850 7440 4950 7450
rect 5050 7530 5150 7540
rect 5050 7450 5060 7530
rect 5140 7450 5150 7530
rect 5050 7440 5150 7450
rect 5250 7530 5350 7540
rect 5250 7450 5260 7530
rect 5340 7450 5350 7530
rect 5250 7440 5350 7450
rect 5450 7530 5550 7540
rect 5450 7450 5460 7530
rect 5540 7450 5550 7530
rect 5450 7440 5550 7450
rect 5650 7530 5750 7540
rect 5650 7450 5660 7530
rect 5740 7450 5750 7530
rect 5650 7440 5750 7450
rect 5850 7530 5950 7540
rect 5850 7450 5860 7530
rect 5940 7450 5950 7530
rect 5850 7440 5950 7450
rect 6050 7530 6150 7540
rect 6050 7450 6060 7530
rect 6140 7450 6150 7530
rect 6050 7440 6150 7450
rect 6250 7530 6350 7540
rect 6250 7450 6260 7530
rect 6340 7450 6350 7530
rect 6250 7440 6350 7450
rect 6450 7530 6550 7540
rect 6450 7450 6460 7530
rect 6540 7450 6550 7530
rect 6450 7440 6550 7450
rect -150 7345 -50 7355
rect -150 7265 -140 7345
rect -60 7265 -50 7345
rect -150 7255 -50 7265
rect 50 7345 150 7355
rect 50 7265 60 7345
rect 140 7265 150 7345
rect 50 7255 150 7265
rect 250 7345 350 7355
rect 250 7265 260 7345
rect 340 7265 350 7345
rect 250 7255 350 7265
rect 450 7345 550 7355
rect 450 7265 460 7345
rect 540 7265 550 7345
rect 450 7255 550 7265
rect 650 7345 750 7355
rect 650 7265 660 7345
rect 740 7265 750 7345
rect 650 7255 750 7265
rect 850 7345 950 7355
rect 850 7265 860 7345
rect 940 7265 950 7345
rect 850 7255 950 7265
rect 1050 7345 1150 7355
rect 1050 7265 1060 7345
rect 1140 7265 1150 7345
rect 1050 7255 1150 7265
rect 1250 7345 1350 7355
rect 1250 7265 1260 7345
rect 1340 7265 1350 7345
rect 1250 7255 1350 7265
rect 1450 7345 1550 7355
rect 1450 7265 1460 7345
rect 1540 7265 1550 7345
rect 1450 7255 1550 7265
rect 1650 7345 1750 7355
rect 1650 7265 1660 7345
rect 1740 7265 1750 7345
rect 1650 7255 1750 7265
rect 1850 7345 1950 7355
rect 1850 7265 1860 7345
rect 1940 7265 1950 7345
rect 1850 7255 1950 7265
rect 2050 7345 2150 7355
rect 2050 7265 2060 7345
rect 2140 7265 2150 7345
rect 2050 7255 2150 7265
rect 2250 7345 2350 7355
rect 2250 7265 2260 7345
rect 2340 7265 2350 7345
rect 2250 7255 2350 7265
rect 2450 7345 2550 7355
rect 2450 7265 2460 7345
rect 2540 7265 2550 7345
rect 2450 7255 2550 7265
rect 2650 7345 2750 7355
rect 2650 7265 2660 7345
rect 2740 7265 2750 7345
rect 2650 7255 2750 7265
rect 2850 7345 2950 7355
rect 2850 7265 2860 7345
rect 2940 7265 2950 7345
rect 2850 7255 2950 7265
rect 3050 7345 3150 7355
rect 3050 7265 3060 7345
rect 3140 7265 3150 7345
rect 3050 7255 3150 7265
rect 3250 7345 3350 7355
rect 3250 7265 3260 7345
rect 3340 7265 3350 7345
rect 3250 7255 3350 7265
rect 3450 7345 3550 7355
rect 3450 7265 3460 7345
rect 3540 7265 3550 7345
rect 3450 7255 3550 7265
rect 3650 7345 3750 7355
rect 3650 7265 3660 7345
rect 3740 7265 3750 7345
rect 3650 7255 3750 7265
rect 3850 7345 3950 7355
rect 3850 7265 3860 7345
rect 3940 7265 3950 7345
rect 3850 7255 3950 7265
rect 4050 7345 4150 7355
rect 4050 7265 4060 7345
rect 4140 7265 4150 7345
rect 4050 7255 4150 7265
rect 4250 7345 4350 7355
rect 4250 7265 4260 7345
rect 4340 7265 4350 7345
rect 4250 7255 4350 7265
rect 4450 7345 4550 7355
rect 4450 7265 4460 7345
rect 4540 7265 4550 7345
rect 4450 7255 4550 7265
rect 4650 7345 4750 7355
rect 4650 7265 4660 7345
rect 4740 7265 4750 7345
rect 4650 7255 4750 7265
rect 4850 7345 4950 7355
rect 4850 7265 4860 7345
rect 4940 7265 4950 7345
rect 4850 7255 4950 7265
rect 5050 7345 5150 7355
rect 5050 7265 5060 7345
rect 5140 7265 5150 7345
rect 5050 7255 5150 7265
rect 5250 7345 5350 7355
rect 5250 7265 5260 7345
rect 5340 7265 5350 7345
rect 5250 7255 5350 7265
rect 5450 7345 5550 7355
rect 5450 7265 5460 7345
rect 5540 7265 5550 7345
rect 5450 7255 5550 7265
rect 5650 7345 5750 7355
rect 5650 7265 5660 7345
rect 5740 7265 5750 7345
rect 5650 7255 5750 7265
rect 5850 7345 5950 7355
rect 5850 7265 5860 7345
rect 5940 7265 5950 7345
rect 5850 7255 5950 7265
rect 6050 7345 6150 7355
rect 6050 7265 6060 7345
rect 6140 7265 6150 7345
rect 6050 7255 6150 7265
rect 6250 7345 6350 7355
rect 6250 7265 6260 7345
rect 6340 7265 6350 7345
rect 6250 7255 6350 7265
rect 6450 7345 6550 7355
rect 6450 7265 6460 7345
rect 6540 7265 6550 7345
rect 6450 7255 6550 7265
rect -150 7160 -50 7170
rect -150 7080 -140 7160
rect -60 7080 -50 7160
rect -150 7070 -50 7080
rect 50 7160 150 7170
rect 50 7080 60 7160
rect 140 7080 150 7160
rect 50 7070 150 7080
rect 250 7160 350 7170
rect 250 7080 260 7160
rect 340 7080 350 7160
rect 250 7070 350 7080
rect 450 7160 550 7170
rect 450 7080 460 7160
rect 540 7080 550 7160
rect 450 7070 550 7080
rect 650 7160 750 7170
rect 650 7080 660 7160
rect 740 7080 750 7160
rect 650 7070 750 7080
rect 850 7160 950 7170
rect 850 7080 860 7160
rect 940 7080 950 7160
rect 850 7070 950 7080
rect 1050 7160 1150 7170
rect 1050 7080 1060 7160
rect 1140 7080 1150 7160
rect 1050 7070 1150 7080
rect 1250 7160 1350 7170
rect 1250 7080 1260 7160
rect 1340 7080 1350 7160
rect 1250 7070 1350 7080
rect 1450 7160 1550 7170
rect 1450 7080 1460 7160
rect 1540 7080 1550 7160
rect 1450 7070 1550 7080
rect 1650 7160 1750 7170
rect 1650 7080 1660 7160
rect 1740 7080 1750 7160
rect 1650 7070 1750 7080
rect 1850 7160 1950 7170
rect 1850 7080 1860 7160
rect 1940 7080 1950 7160
rect 1850 7070 1950 7080
rect 2050 7160 2150 7170
rect 2050 7080 2060 7160
rect 2140 7080 2150 7160
rect 2050 7070 2150 7080
rect 2250 7160 2350 7170
rect 2250 7080 2260 7160
rect 2340 7080 2350 7160
rect 2250 7070 2350 7080
rect 2450 7160 2550 7170
rect 2450 7080 2460 7160
rect 2540 7080 2550 7160
rect 2450 7070 2550 7080
rect 2650 7160 2750 7170
rect 2650 7080 2660 7160
rect 2740 7080 2750 7160
rect 2650 7070 2750 7080
rect 2850 7160 2950 7170
rect 2850 7080 2860 7160
rect 2940 7080 2950 7160
rect 2850 7070 2950 7080
rect 3050 7160 3150 7170
rect 3050 7080 3060 7160
rect 3140 7080 3150 7160
rect 3050 7070 3150 7080
rect 3250 7160 3350 7170
rect 3250 7080 3260 7160
rect 3340 7080 3350 7160
rect 3250 7070 3350 7080
rect 3450 7160 3550 7170
rect 3450 7080 3460 7160
rect 3540 7080 3550 7160
rect 3450 7070 3550 7080
rect 3650 7160 3750 7170
rect 3650 7080 3660 7160
rect 3740 7080 3750 7160
rect 3650 7070 3750 7080
rect 3850 7160 3950 7170
rect 3850 7080 3860 7160
rect 3940 7080 3950 7160
rect 3850 7070 3950 7080
rect 4050 7160 4150 7170
rect 4050 7080 4060 7160
rect 4140 7080 4150 7160
rect 4050 7070 4150 7080
rect 4250 7160 4350 7170
rect 4250 7080 4260 7160
rect 4340 7080 4350 7160
rect 4250 7070 4350 7080
rect 4450 7160 4550 7170
rect 4450 7080 4460 7160
rect 4540 7080 4550 7160
rect 4450 7070 4550 7080
rect 4650 7160 4750 7170
rect 4650 7080 4660 7160
rect 4740 7080 4750 7160
rect 4650 7070 4750 7080
rect 4850 7160 4950 7170
rect 4850 7080 4860 7160
rect 4940 7080 4950 7160
rect 4850 7070 4950 7080
rect 5050 7160 5150 7170
rect 5050 7080 5060 7160
rect 5140 7080 5150 7160
rect 5050 7070 5150 7080
rect 5250 7160 5350 7170
rect 5250 7080 5260 7160
rect 5340 7080 5350 7160
rect 5250 7070 5350 7080
rect 5450 7160 5550 7170
rect 5450 7080 5460 7160
rect 5540 7080 5550 7160
rect 5450 7070 5550 7080
rect 5650 7160 5750 7170
rect 5650 7080 5660 7160
rect 5740 7080 5750 7160
rect 5650 7070 5750 7080
rect 5850 7160 5950 7170
rect 5850 7080 5860 7160
rect 5940 7080 5950 7160
rect 5850 7070 5950 7080
rect 6050 7160 6150 7170
rect 6050 7080 6060 7160
rect 6140 7080 6150 7160
rect 6050 7070 6150 7080
rect 6250 7160 6350 7170
rect 6250 7080 6260 7160
rect 6340 7080 6350 7160
rect 6250 7070 6350 7080
rect 6450 7160 6550 7170
rect 6450 7080 6460 7160
rect 6540 7080 6550 7160
rect 6450 7070 6550 7080
rect -150 6975 -50 6985
rect -150 6895 -140 6975
rect -60 6895 -50 6975
rect -150 6885 -50 6895
rect 50 6975 150 6985
rect 50 6895 60 6975
rect 140 6895 150 6975
rect 50 6885 150 6895
rect 250 6975 350 6985
rect 250 6895 260 6975
rect 340 6895 350 6975
rect 250 6885 350 6895
rect 450 6975 550 6985
rect 450 6895 460 6975
rect 540 6895 550 6975
rect 450 6885 550 6895
rect 650 6975 750 6985
rect 650 6895 660 6975
rect 740 6895 750 6975
rect 650 6885 750 6895
rect 850 6975 950 6985
rect 850 6895 860 6975
rect 940 6895 950 6975
rect 850 6885 950 6895
rect 1050 6975 1150 6985
rect 1050 6895 1060 6975
rect 1140 6895 1150 6975
rect 1050 6885 1150 6895
rect 1250 6975 1350 6985
rect 1250 6895 1260 6975
rect 1340 6895 1350 6975
rect 1250 6885 1350 6895
rect 1450 6975 1550 6985
rect 1450 6895 1460 6975
rect 1540 6895 1550 6975
rect 1450 6885 1550 6895
rect 1650 6975 1750 6985
rect 1650 6895 1660 6975
rect 1740 6895 1750 6975
rect 1650 6885 1750 6895
rect 1850 6975 1950 6985
rect 1850 6895 1860 6975
rect 1940 6895 1950 6975
rect 1850 6885 1950 6895
rect 2050 6975 2150 6985
rect 2050 6895 2060 6975
rect 2140 6895 2150 6975
rect 2050 6885 2150 6895
rect 2250 6975 2350 6985
rect 2250 6895 2260 6975
rect 2340 6895 2350 6975
rect 2250 6885 2350 6895
rect 2450 6975 2550 6985
rect 2450 6895 2460 6975
rect 2540 6895 2550 6975
rect 2450 6885 2550 6895
rect 2650 6975 2750 6985
rect 2650 6895 2660 6975
rect 2740 6895 2750 6975
rect 2650 6885 2750 6895
rect 2850 6975 2950 6985
rect 2850 6895 2860 6975
rect 2940 6895 2950 6975
rect 2850 6885 2950 6895
rect 3050 6975 3150 6985
rect 3050 6895 3060 6975
rect 3140 6895 3150 6975
rect 3050 6885 3150 6895
rect 3250 6975 3350 6985
rect 3250 6895 3260 6975
rect 3340 6895 3350 6975
rect 3250 6885 3350 6895
rect 3450 6975 3550 6985
rect 3450 6895 3460 6975
rect 3540 6895 3550 6975
rect 3450 6885 3550 6895
rect 3650 6975 3750 6985
rect 3650 6895 3660 6975
rect 3740 6895 3750 6975
rect 3650 6885 3750 6895
rect 3850 6975 3950 6985
rect 3850 6895 3860 6975
rect 3940 6895 3950 6975
rect 3850 6885 3950 6895
rect 4050 6975 4150 6985
rect 4050 6895 4060 6975
rect 4140 6895 4150 6975
rect 4050 6885 4150 6895
rect 4250 6975 4350 6985
rect 4250 6895 4260 6975
rect 4340 6895 4350 6975
rect 4250 6885 4350 6895
rect 4450 6975 4550 6985
rect 4450 6895 4460 6975
rect 4540 6895 4550 6975
rect 4450 6885 4550 6895
rect 4650 6975 4750 6985
rect 4650 6895 4660 6975
rect 4740 6895 4750 6975
rect 4650 6885 4750 6895
rect 4850 6975 4950 6985
rect 4850 6895 4860 6975
rect 4940 6895 4950 6975
rect 4850 6885 4950 6895
rect 5050 6975 5150 6985
rect 5050 6895 5060 6975
rect 5140 6895 5150 6975
rect 5050 6885 5150 6895
rect 5250 6975 5350 6985
rect 5250 6895 5260 6975
rect 5340 6895 5350 6975
rect 5250 6885 5350 6895
rect 5450 6975 5550 6985
rect 5450 6895 5460 6975
rect 5540 6895 5550 6975
rect 5450 6885 5550 6895
rect 5650 6975 5750 6985
rect 5650 6895 5660 6975
rect 5740 6895 5750 6975
rect 5650 6885 5750 6895
rect 5850 6975 5950 6985
rect 5850 6895 5860 6975
rect 5940 6895 5950 6975
rect 5850 6885 5950 6895
rect 6050 6975 6150 6985
rect 6050 6895 6060 6975
rect 6140 6895 6150 6975
rect 6050 6885 6150 6895
rect 6250 6975 6350 6985
rect 6250 6895 6260 6975
rect 6340 6895 6350 6975
rect 6250 6885 6350 6895
rect 6450 6975 6550 6985
rect 6450 6895 6460 6975
rect 6540 6895 6550 6975
rect 6450 6885 6550 6895
rect -150 6790 -50 6800
rect -150 6710 -140 6790
rect -60 6710 -50 6790
rect -150 6700 -50 6710
rect 50 6790 150 6800
rect 50 6710 60 6790
rect 140 6710 150 6790
rect 50 6700 150 6710
rect 250 6790 350 6800
rect 250 6710 260 6790
rect 340 6710 350 6790
rect 250 6700 350 6710
rect 450 6790 550 6800
rect 450 6710 460 6790
rect 540 6710 550 6790
rect 450 6700 550 6710
rect 650 6790 750 6800
rect 650 6710 660 6790
rect 740 6710 750 6790
rect 650 6700 750 6710
rect 850 6790 950 6800
rect 850 6710 860 6790
rect 940 6710 950 6790
rect 850 6700 950 6710
rect 1050 6790 1150 6800
rect 1050 6710 1060 6790
rect 1140 6710 1150 6790
rect 1050 6700 1150 6710
rect 1250 6790 1350 6800
rect 1250 6710 1260 6790
rect 1340 6710 1350 6790
rect 1250 6700 1350 6710
rect 1450 6790 1550 6800
rect 1450 6710 1460 6790
rect 1540 6710 1550 6790
rect 1450 6700 1550 6710
rect 1650 6790 1750 6800
rect 1650 6710 1660 6790
rect 1740 6710 1750 6790
rect 1650 6700 1750 6710
rect 1850 6790 1950 6800
rect 1850 6710 1860 6790
rect 1940 6710 1950 6790
rect 1850 6700 1950 6710
rect 2050 6790 2150 6800
rect 2050 6710 2060 6790
rect 2140 6710 2150 6790
rect 2050 6700 2150 6710
rect 2250 6790 2350 6800
rect 2250 6710 2260 6790
rect 2340 6710 2350 6790
rect 2250 6700 2350 6710
rect 2450 6790 2550 6800
rect 2450 6710 2460 6790
rect 2540 6710 2550 6790
rect 2450 6700 2550 6710
rect 2650 6790 2750 6800
rect 2650 6710 2660 6790
rect 2740 6710 2750 6790
rect 2650 6700 2750 6710
rect 2850 6790 2950 6800
rect 2850 6710 2860 6790
rect 2940 6710 2950 6790
rect 2850 6700 2950 6710
rect 3050 6790 3150 6800
rect 3050 6710 3060 6790
rect 3140 6710 3150 6790
rect 3050 6700 3150 6710
rect 3250 6790 3350 6800
rect 3250 6710 3260 6790
rect 3340 6710 3350 6790
rect 3250 6700 3350 6710
rect 3450 6790 3550 6800
rect 3450 6710 3460 6790
rect 3540 6710 3550 6790
rect 3450 6700 3550 6710
rect 3650 6790 3750 6800
rect 3650 6710 3660 6790
rect 3740 6710 3750 6790
rect 3650 6700 3750 6710
rect 3850 6790 3950 6800
rect 3850 6710 3860 6790
rect 3940 6710 3950 6790
rect 3850 6700 3950 6710
rect 4050 6790 4150 6800
rect 4050 6710 4060 6790
rect 4140 6710 4150 6790
rect 4050 6700 4150 6710
rect 4250 6790 4350 6800
rect 4250 6710 4260 6790
rect 4340 6710 4350 6790
rect 4250 6700 4350 6710
rect 4450 6790 4550 6800
rect 4450 6710 4460 6790
rect 4540 6710 4550 6790
rect 4450 6700 4550 6710
rect 4650 6790 4750 6800
rect 4650 6710 4660 6790
rect 4740 6710 4750 6790
rect 4650 6700 4750 6710
rect 4850 6790 4950 6800
rect 4850 6710 4860 6790
rect 4940 6710 4950 6790
rect 4850 6700 4950 6710
rect 5050 6790 5150 6800
rect 5050 6710 5060 6790
rect 5140 6710 5150 6790
rect 5050 6700 5150 6710
rect 5250 6790 5350 6800
rect 5250 6710 5260 6790
rect 5340 6710 5350 6790
rect 5250 6700 5350 6710
rect 5450 6790 5550 6800
rect 5450 6710 5460 6790
rect 5540 6710 5550 6790
rect 5450 6700 5550 6710
rect 5650 6790 5750 6800
rect 5650 6710 5660 6790
rect 5740 6710 5750 6790
rect 5650 6700 5750 6710
rect 5850 6790 5950 6800
rect 5850 6710 5860 6790
rect 5940 6710 5950 6790
rect 5850 6700 5950 6710
rect 6050 6790 6150 6800
rect 6050 6710 6060 6790
rect 6140 6710 6150 6790
rect 6050 6700 6150 6710
rect 6250 6790 6350 6800
rect 6250 6710 6260 6790
rect 6340 6710 6350 6790
rect 6250 6700 6350 6710
rect 6450 6790 6550 6800
rect 6450 6710 6460 6790
rect 6540 6710 6550 6790
rect 6450 6700 6550 6710
rect -150 6605 -50 6615
rect -150 6525 -140 6605
rect -60 6525 -50 6605
rect -150 6515 -50 6525
rect 50 6605 150 6615
rect 50 6525 60 6605
rect 140 6525 150 6605
rect 50 6515 150 6525
rect 250 6605 350 6615
rect 250 6525 260 6605
rect 340 6525 350 6605
rect 250 6515 350 6525
rect 450 6605 550 6615
rect 450 6525 460 6605
rect 540 6525 550 6605
rect 450 6515 550 6525
rect 650 6605 750 6615
rect 650 6525 660 6605
rect 740 6525 750 6605
rect 650 6515 750 6525
rect 850 6605 950 6615
rect 850 6525 860 6605
rect 940 6525 950 6605
rect 850 6515 950 6525
rect 1050 6605 1150 6615
rect 1050 6525 1060 6605
rect 1140 6525 1150 6605
rect 1050 6515 1150 6525
rect 1250 6605 1350 6615
rect 1250 6525 1260 6605
rect 1340 6525 1350 6605
rect 1250 6515 1350 6525
rect 1450 6605 1550 6615
rect 1450 6525 1460 6605
rect 1540 6525 1550 6605
rect 1450 6515 1550 6525
rect 1650 6605 1750 6615
rect 1650 6525 1660 6605
rect 1740 6525 1750 6605
rect 1650 6515 1750 6525
rect 1850 6605 1950 6615
rect 1850 6525 1860 6605
rect 1940 6525 1950 6605
rect 1850 6515 1950 6525
rect 2050 6605 2150 6615
rect 2050 6525 2060 6605
rect 2140 6525 2150 6605
rect 2050 6515 2150 6525
rect 2250 6605 2350 6615
rect 2250 6525 2260 6605
rect 2340 6525 2350 6605
rect 2250 6515 2350 6525
rect 2450 6605 2550 6615
rect 2450 6525 2460 6605
rect 2540 6525 2550 6605
rect 2450 6515 2550 6525
rect 2650 6605 2750 6615
rect 2650 6525 2660 6605
rect 2740 6525 2750 6605
rect 2650 6515 2750 6525
rect 2850 6605 2950 6615
rect 2850 6525 2860 6605
rect 2940 6525 2950 6605
rect 2850 6515 2950 6525
rect 3050 6605 3150 6615
rect 3050 6525 3060 6605
rect 3140 6525 3150 6605
rect 3050 6515 3150 6525
rect 3250 6605 3350 6615
rect 3250 6525 3260 6605
rect 3340 6525 3350 6605
rect 3250 6515 3350 6525
rect 3450 6605 3550 6615
rect 3450 6525 3460 6605
rect 3540 6525 3550 6605
rect 3450 6515 3550 6525
rect 3650 6605 3750 6615
rect 3650 6525 3660 6605
rect 3740 6525 3750 6605
rect 3650 6515 3750 6525
rect 3850 6605 3950 6615
rect 3850 6525 3860 6605
rect 3940 6525 3950 6605
rect 3850 6515 3950 6525
rect 4050 6605 4150 6615
rect 4050 6525 4060 6605
rect 4140 6525 4150 6605
rect 4050 6515 4150 6525
rect 4250 6605 4350 6615
rect 4250 6525 4260 6605
rect 4340 6525 4350 6605
rect 4250 6515 4350 6525
rect 4450 6605 4550 6615
rect 4450 6525 4460 6605
rect 4540 6525 4550 6605
rect 4450 6515 4550 6525
rect 4650 6605 4750 6615
rect 4650 6525 4660 6605
rect 4740 6525 4750 6605
rect 4650 6515 4750 6525
rect 4850 6605 4950 6615
rect 4850 6525 4860 6605
rect 4940 6525 4950 6605
rect 4850 6515 4950 6525
rect 5050 6605 5150 6615
rect 5050 6525 5060 6605
rect 5140 6525 5150 6605
rect 5050 6515 5150 6525
rect 5250 6605 5350 6615
rect 5250 6525 5260 6605
rect 5340 6525 5350 6605
rect 5250 6515 5350 6525
rect 5450 6605 5550 6615
rect 5450 6525 5460 6605
rect 5540 6525 5550 6605
rect 5450 6515 5550 6525
rect 5650 6605 5750 6615
rect 5650 6525 5660 6605
rect 5740 6525 5750 6605
rect 5650 6515 5750 6525
rect 5850 6605 5950 6615
rect 5850 6525 5860 6605
rect 5940 6525 5950 6605
rect 5850 6515 5950 6525
rect 6050 6605 6150 6615
rect 6050 6525 6060 6605
rect 6140 6525 6150 6605
rect 6050 6515 6150 6525
rect 6250 6605 6350 6615
rect 6250 6525 6260 6605
rect 6340 6525 6350 6605
rect 6250 6515 6350 6525
rect 6450 6605 6550 6615
rect 6450 6525 6460 6605
rect 6540 6525 6550 6605
rect 6450 6515 6550 6525
rect -150 6420 -50 6430
rect -150 6340 -140 6420
rect -60 6340 -50 6420
rect -150 6330 -50 6340
rect 50 6420 150 6430
rect 50 6340 60 6420
rect 140 6340 150 6420
rect 50 6330 150 6340
rect 250 6420 350 6430
rect 250 6340 260 6420
rect 340 6340 350 6420
rect 250 6330 350 6340
rect 450 6420 550 6430
rect 450 6340 460 6420
rect 540 6340 550 6420
rect 450 6330 550 6340
rect 650 6420 750 6430
rect 650 6340 660 6420
rect 740 6340 750 6420
rect 650 6330 750 6340
rect 850 6420 950 6430
rect 850 6340 860 6420
rect 940 6340 950 6420
rect 850 6330 950 6340
rect 1050 6420 1150 6430
rect 1050 6340 1060 6420
rect 1140 6340 1150 6420
rect 1050 6330 1150 6340
rect 1250 6420 1350 6430
rect 1250 6340 1260 6420
rect 1340 6340 1350 6420
rect 1250 6330 1350 6340
rect 1450 6420 1550 6430
rect 1450 6340 1460 6420
rect 1540 6340 1550 6420
rect 1450 6330 1550 6340
rect 1650 6420 1750 6430
rect 1650 6340 1660 6420
rect 1740 6340 1750 6420
rect 1650 6330 1750 6340
rect 1850 6420 1950 6430
rect 1850 6340 1860 6420
rect 1940 6340 1950 6420
rect 1850 6330 1950 6340
rect 2050 6420 2150 6430
rect 2050 6340 2060 6420
rect 2140 6340 2150 6420
rect 2050 6330 2150 6340
rect 2250 6420 2350 6430
rect 2250 6340 2260 6420
rect 2340 6340 2350 6420
rect 2250 6330 2350 6340
rect 2450 6420 2550 6430
rect 2450 6340 2460 6420
rect 2540 6340 2550 6420
rect 2450 6330 2550 6340
rect 2650 6420 2750 6430
rect 2650 6340 2660 6420
rect 2740 6340 2750 6420
rect 2650 6330 2750 6340
rect 2850 6420 2950 6430
rect 2850 6340 2860 6420
rect 2940 6340 2950 6420
rect 2850 6330 2950 6340
rect 3050 6420 3150 6430
rect 3050 6340 3060 6420
rect 3140 6340 3150 6420
rect 3050 6330 3150 6340
rect 3250 6420 3350 6430
rect 3250 6340 3260 6420
rect 3340 6340 3350 6420
rect 3250 6330 3350 6340
rect 3450 6420 3550 6430
rect 3450 6340 3460 6420
rect 3540 6340 3550 6420
rect 3450 6330 3550 6340
rect 3650 6420 3750 6430
rect 3650 6340 3660 6420
rect 3740 6340 3750 6420
rect 3650 6330 3750 6340
rect 3850 6420 3950 6430
rect 3850 6340 3860 6420
rect 3940 6340 3950 6420
rect 3850 6330 3950 6340
rect 4050 6420 4150 6430
rect 4050 6340 4060 6420
rect 4140 6340 4150 6420
rect 4050 6330 4150 6340
rect 4250 6420 4350 6430
rect 4250 6340 4260 6420
rect 4340 6340 4350 6420
rect 4250 6330 4350 6340
rect 4450 6420 4550 6430
rect 4450 6340 4460 6420
rect 4540 6340 4550 6420
rect 4450 6330 4550 6340
rect 4650 6420 4750 6430
rect 4650 6340 4660 6420
rect 4740 6340 4750 6420
rect 4650 6330 4750 6340
rect 4850 6420 4950 6430
rect 4850 6340 4860 6420
rect 4940 6340 4950 6420
rect 4850 6330 4950 6340
rect 5050 6420 5150 6430
rect 5050 6340 5060 6420
rect 5140 6340 5150 6420
rect 5050 6330 5150 6340
rect 5250 6420 5350 6430
rect 5250 6340 5260 6420
rect 5340 6340 5350 6420
rect 5250 6330 5350 6340
rect 5450 6420 5550 6430
rect 5450 6340 5460 6420
rect 5540 6340 5550 6420
rect 5450 6330 5550 6340
rect 5650 6420 5750 6430
rect 5650 6340 5660 6420
rect 5740 6340 5750 6420
rect 5650 6330 5750 6340
rect 5850 6420 5950 6430
rect 5850 6340 5860 6420
rect 5940 6340 5950 6420
rect 5850 6330 5950 6340
rect 6050 6420 6150 6430
rect 6050 6340 6060 6420
rect 6140 6340 6150 6420
rect 6050 6330 6150 6340
rect 6250 6420 6350 6430
rect 6250 6340 6260 6420
rect 6340 6340 6350 6420
rect 6250 6330 6350 6340
rect 6450 6420 6550 6430
rect 6450 6340 6460 6420
rect 6540 6340 6550 6420
rect 6450 6330 6550 6340
rect -150 6235 -50 6245
rect -150 6155 -140 6235
rect -60 6155 -50 6235
rect -150 6145 -50 6155
rect 50 6235 150 6245
rect 50 6155 60 6235
rect 140 6155 150 6235
rect 50 6145 150 6155
rect 250 6235 350 6245
rect 250 6155 260 6235
rect 340 6155 350 6235
rect 250 6145 350 6155
rect 450 6235 550 6245
rect 450 6155 460 6235
rect 540 6155 550 6235
rect 450 6145 550 6155
rect 650 6235 750 6245
rect 650 6155 660 6235
rect 740 6155 750 6235
rect 650 6145 750 6155
rect 850 6235 950 6245
rect 850 6155 860 6235
rect 940 6155 950 6235
rect 850 6145 950 6155
rect 1050 6235 1150 6245
rect 1050 6155 1060 6235
rect 1140 6155 1150 6235
rect 1050 6145 1150 6155
rect 1250 6235 1350 6245
rect 1250 6155 1260 6235
rect 1340 6155 1350 6235
rect 1250 6145 1350 6155
rect 1450 6235 1550 6245
rect 1450 6155 1460 6235
rect 1540 6155 1550 6235
rect 1450 6145 1550 6155
rect 1650 6235 1750 6245
rect 1650 6155 1660 6235
rect 1740 6155 1750 6235
rect 1650 6145 1750 6155
rect 1850 6235 1950 6245
rect 1850 6155 1860 6235
rect 1940 6155 1950 6235
rect 1850 6145 1950 6155
rect 2050 6235 2150 6245
rect 2050 6155 2060 6235
rect 2140 6155 2150 6235
rect 2050 6145 2150 6155
rect 2250 6235 2350 6245
rect 2250 6155 2260 6235
rect 2340 6155 2350 6235
rect 2250 6145 2350 6155
rect 2450 6235 2550 6245
rect 2450 6155 2460 6235
rect 2540 6155 2550 6235
rect 2450 6145 2550 6155
rect 2650 6235 2750 6245
rect 2650 6155 2660 6235
rect 2740 6155 2750 6235
rect 2650 6145 2750 6155
rect 2850 6235 2950 6245
rect 2850 6155 2860 6235
rect 2940 6155 2950 6235
rect 2850 6145 2950 6155
rect 3050 6235 3150 6245
rect 3050 6155 3060 6235
rect 3140 6155 3150 6235
rect 3050 6145 3150 6155
rect 3250 6235 3350 6245
rect 3250 6155 3260 6235
rect 3340 6155 3350 6235
rect 3250 6145 3350 6155
rect 3450 6235 3550 6245
rect 3450 6155 3460 6235
rect 3540 6155 3550 6235
rect 3450 6145 3550 6155
rect 3650 6235 3750 6245
rect 3650 6155 3660 6235
rect 3740 6155 3750 6235
rect 3650 6145 3750 6155
rect 3850 6235 3950 6245
rect 3850 6155 3860 6235
rect 3940 6155 3950 6235
rect 3850 6145 3950 6155
rect 4050 6235 4150 6245
rect 4050 6155 4060 6235
rect 4140 6155 4150 6235
rect 4050 6145 4150 6155
rect 4250 6235 4350 6245
rect 4250 6155 4260 6235
rect 4340 6155 4350 6235
rect 4250 6145 4350 6155
rect 4450 6235 4550 6245
rect 4450 6155 4460 6235
rect 4540 6155 4550 6235
rect 4450 6145 4550 6155
rect 4650 6235 4750 6245
rect 4650 6155 4660 6235
rect 4740 6155 4750 6235
rect 4650 6145 4750 6155
rect 4850 6235 4950 6245
rect 4850 6155 4860 6235
rect 4940 6155 4950 6235
rect 4850 6145 4950 6155
rect 5050 6235 5150 6245
rect 5050 6155 5060 6235
rect 5140 6155 5150 6235
rect 5050 6145 5150 6155
rect 5250 6235 5350 6245
rect 5250 6155 5260 6235
rect 5340 6155 5350 6235
rect 5250 6145 5350 6155
rect 5450 6235 5550 6245
rect 5450 6155 5460 6235
rect 5540 6155 5550 6235
rect 5450 6145 5550 6155
rect 5650 6235 5750 6245
rect 5650 6155 5660 6235
rect 5740 6155 5750 6235
rect 5650 6145 5750 6155
rect 5850 6235 5950 6245
rect 5850 6155 5860 6235
rect 5940 6155 5950 6235
rect 5850 6145 5950 6155
rect 6050 6235 6150 6245
rect 6050 6155 6060 6235
rect 6140 6155 6150 6235
rect 6050 6145 6150 6155
rect 6250 6235 6350 6245
rect 6250 6155 6260 6235
rect 6340 6155 6350 6235
rect 6250 6145 6350 6155
rect 6450 6235 6550 6245
rect 6450 6155 6460 6235
rect 6540 6155 6550 6235
rect 6450 6145 6550 6155
rect -150 6050 -50 6060
rect -150 5970 -140 6050
rect -60 5970 -50 6050
rect -150 5960 -50 5970
rect 50 6050 150 6060
rect 50 5970 60 6050
rect 140 5970 150 6050
rect 50 5960 150 5970
rect 250 6050 350 6060
rect 250 5970 260 6050
rect 340 5970 350 6050
rect 250 5960 350 5970
rect 450 6050 550 6060
rect 450 5970 460 6050
rect 540 5970 550 6050
rect 450 5960 550 5970
rect 650 6050 750 6060
rect 650 5970 660 6050
rect 740 5970 750 6050
rect 650 5960 750 5970
rect 850 6050 950 6060
rect 850 5970 860 6050
rect 940 5970 950 6050
rect 850 5960 950 5970
rect 1050 6050 1150 6060
rect 1050 5970 1060 6050
rect 1140 5970 1150 6050
rect 1050 5960 1150 5970
rect 1250 6050 1350 6060
rect 1250 5970 1260 6050
rect 1340 5970 1350 6050
rect 1250 5960 1350 5970
rect 1450 6050 1550 6060
rect 1450 5970 1460 6050
rect 1540 5970 1550 6050
rect 1450 5960 1550 5970
rect 1650 6050 1750 6060
rect 1650 5970 1660 6050
rect 1740 5970 1750 6050
rect 1650 5960 1750 5970
rect 1850 6050 1950 6060
rect 1850 5970 1860 6050
rect 1940 5970 1950 6050
rect 1850 5960 1950 5970
rect 2050 6050 2150 6060
rect 2050 5970 2060 6050
rect 2140 5970 2150 6050
rect 2050 5960 2150 5970
rect 2250 6050 2350 6060
rect 2250 5970 2260 6050
rect 2340 5970 2350 6050
rect 2250 5960 2350 5970
rect 2450 6050 2550 6060
rect 2450 5970 2460 6050
rect 2540 5970 2550 6050
rect 2450 5960 2550 5970
rect 2650 6050 2750 6060
rect 2650 5970 2660 6050
rect 2740 5970 2750 6050
rect 2650 5960 2750 5970
rect 2850 6050 2950 6060
rect 2850 5970 2860 6050
rect 2940 5970 2950 6050
rect 2850 5960 2950 5970
rect 3050 6050 3150 6060
rect 3050 5970 3060 6050
rect 3140 5970 3150 6050
rect 3050 5960 3150 5970
rect 3250 6050 3350 6060
rect 3250 5970 3260 6050
rect 3340 5970 3350 6050
rect 3250 5960 3350 5970
rect 3450 6050 3550 6060
rect 3450 5970 3460 6050
rect 3540 5970 3550 6050
rect 3450 5960 3550 5970
rect 3650 6050 3750 6060
rect 3650 5970 3660 6050
rect 3740 5970 3750 6050
rect 3650 5960 3750 5970
rect 3850 6050 3950 6060
rect 3850 5970 3860 6050
rect 3940 5970 3950 6050
rect 3850 5960 3950 5970
rect 4050 6050 4150 6060
rect 4050 5970 4060 6050
rect 4140 5970 4150 6050
rect 4050 5960 4150 5970
rect 4250 6050 4350 6060
rect 4250 5970 4260 6050
rect 4340 5970 4350 6050
rect 4250 5960 4350 5970
rect 4450 6050 4550 6060
rect 4450 5970 4460 6050
rect 4540 5970 4550 6050
rect 4450 5960 4550 5970
rect 4650 6050 4750 6060
rect 4650 5970 4660 6050
rect 4740 5970 4750 6050
rect 4650 5960 4750 5970
rect 4850 6050 4950 6060
rect 4850 5970 4860 6050
rect 4940 5970 4950 6050
rect 4850 5960 4950 5970
rect 5050 6050 5150 6060
rect 5050 5970 5060 6050
rect 5140 5970 5150 6050
rect 5050 5960 5150 5970
rect 5250 6050 5350 6060
rect 5250 5970 5260 6050
rect 5340 5970 5350 6050
rect 5250 5960 5350 5970
rect 5450 6050 5550 6060
rect 5450 5970 5460 6050
rect 5540 5970 5550 6050
rect 5450 5960 5550 5970
rect 5650 6050 5750 6060
rect 5650 5970 5660 6050
rect 5740 5970 5750 6050
rect 5650 5960 5750 5970
rect 5850 6050 5950 6060
rect 5850 5970 5860 6050
rect 5940 5970 5950 6050
rect 5850 5960 5950 5970
rect 6050 6050 6150 6060
rect 6050 5970 6060 6050
rect 6140 5970 6150 6050
rect 6050 5960 6150 5970
rect 6250 6050 6350 6060
rect 6250 5970 6260 6050
rect 6340 5970 6350 6050
rect 6250 5960 6350 5970
rect 6450 6050 6550 6060
rect 6450 5970 6460 6050
rect 6540 5970 6550 6050
rect 6450 5960 6550 5970
rect -150 5865 -50 5875
rect -150 5785 -140 5865
rect -60 5785 -50 5865
rect -150 5775 -50 5785
rect 50 5865 150 5875
rect 50 5785 60 5865
rect 140 5785 150 5865
rect 50 5775 150 5785
rect 250 5865 350 5875
rect 250 5785 260 5865
rect 340 5785 350 5865
rect 250 5775 350 5785
rect 450 5865 550 5875
rect 450 5785 460 5865
rect 540 5785 550 5865
rect 450 5775 550 5785
rect 650 5865 750 5875
rect 650 5785 660 5865
rect 740 5785 750 5865
rect 650 5775 750 5785
rect 850 5865 950 5875
rect 850 5785 860 5865
rect 940 5785 950 5865
rect 850 5775 950 5785
rect 1050 5865 1150 5875
rect 1050 5785 1060 5865
rect 1140 5785 1150 5865
rect 1050 5775 1150 5785
rect 1250 5865 1350 5875
rect 1250 5785 1260 5865
rect 1340 5785 1350 5865
rect 1250 5775 1350 5785
rect 1450 5865 1550 5875
rect 1450 5785 1460 5865
rect 1540 5785 1550 5865
rect 1450 5775 1550 5785
rect 1650 5865 1750 5875
rect 1650 5785 1660 5865
rect 1740 5785 1750 5865
rect 1650 5775 1750 5785
rect 1850 5865 1950 5875
rect 1850 5785 1860 5865
rect 1940 5785 1950 5865
rect 1850 5775 1950 5785
rect 2050 5865 2150 5875
rect 2050 5785 2060 5865
rect 2140 5785 2150 5865
rect 2050 5775 2150 5785
rect 2250 5865 2350 5875
rect 2250 5785 2260 5865
rect 2340 5785 2350 5865
rect 2250 5775 2350 5785
rect 2450 5865 2550 5875
rect 2450 5785 2460 5865
rect 2540 5785 2550 5865
rect 2450 5775 2550 5785
rect 2650 5865 2750 5875
rect 2650 5785 2660 5865
rect 2740 5785 2750 5865
rect 2650 5775 2750 5785
rect 2850 5865 2950 5875
rect 2850 5785 2860 5865
rect 2940 5785 2950 5865
rect 2850 5775 2950 5785
rect 3050 5865 3150 5875
rect 3050 5785 3060 5865
rect 3140 5785 3150 5865
rect 3050 5775 3150 5785
rect 3250 5865 3350 5875
rect 3250 5785 3260 5865
rect 3340 5785 3350 5865
rect 3250 5775 3350 5785
rect 3450 5865 3550 5875
rect 3450 5785 3460 5865
rect 3540 5785 3550 5865
rect 3450 5775 3550 5785
rect 3650 5865 3750 5875
rect 3650 5785 3660 5865
rect 3740 5785 3750 5865
rect 3650 5775 3750 5785
rect 3850 5865 3950 5875
rect 3850 5785 3860 5865
rect 3940 5785 3950 5865
rect 3850 5775 3950 5785
rect 4050 5865 4150 5875
rect 4050 5785 4060 5865
rect 4140 5785 4150 5865
rect 4050 5775 4150 5785
rect 4250 5865 4350 5875
rect 4250 5785 4260 5865
rect 4340 5785 4350 5865
rect 4250 5775 4350 5785
rect 4450 5865 4550 5875
rect 4450 5785 4460 5865
rect 4540 5785 4550 5865
rect 4450 5775 4550 5785
rect 4650 5865 4750 5875
rect 4650 5785 4660 5865
rect 4740 5785 4750 5865
rect 4650 5775 4750 5785
rect 4850 5865 4950 5875
rect 4850 5785 4860 5865
rect 4940 5785 4950 5865
rect 4850 5775 4950 5785
rect 5050 5865 5150 5875
rect 5050 5785 5060 5865
rect 5140 5785 5150 5865
rect 5050 5775 5150 5785
rect 5250 5865 5350 5875
rect 5250 5785 5260 5865
rect 5340 5785 5350 5865
rect 5250 5775 5350 5785
rect 5450 5865 5550 5875
rect 5450 5785 5460 5865
rect 5540 5785 5550 5865
rect 5450 5775 5550 5785
rect 5650 5865 5750 5875
rect 5650 5785 5660 5865
rect 5740 5785 5750 5865
rect 5650 5775 5750 5785
rect 5850 5865 5950 5875
rect 5850 5785 5860 5865
rect 5940 5785 5950 5865
rect 5850 5775 5950 5785
rect 6050 5865 6150 5875
rect 6050 5785 6060 5865
rect 6140 5785 6150 5865
rect 6050 5775 6150 5785
rect 6250 5865 6350 5875
rect 6250 5785 6260 5865
rect 6340 5785 6350 5865
rect 6250 5775 6350 5785
rect 6450 5865 6550 5875
rect 6450 5785 6460 5865
rect 6540 5785 6550 5865
rect 6450 5775 6550 5785
rect -150 5680 -50 5690
rect -150 5600 -140 5680
rect -60 5600 -50 5680
rect -150 5590 -50 5600
rect 50 5680 150 5690
rect 50 5600 60 5680
rect 140 5600 150 5680
rect 50 5590 150 5600
rect 250 5680 350 5690
rect 250 5600 260 5680
rect 340 5600 350 5680
rect 250 5590 350 5600
rect 450 5680 550 5690
rect 450 5600 460 5680
rect 540 5600 550 5680
rect 450 5590 550 5600
rect 650 5680 750 5690
rect 650 5600 660 5680
rect 740 5600 750 5680
rect 650 5590 750 5600
rect 850 5680 950 5690
rect 850 5600 860 5680
rect 940 5600 950 5680
rect 850 5590 950 5600
rect 1050 5680 1150 5690
rect 1050 5600 1060 5680
rect 1140 5600 1150 5680
rect 1050 5590 1150 5600
rect 1250 5680 1350 5690
rect 1250 5600 1260 5680
rect 1340 5600 1350 5680
rect 1250 5590 1350 5600
rect 1450 5680 1550 5690
rect 1450 5600 1460 5680
rect 1540 5600 1550 5680
rect 1450 5590 1550 5600
rect 1650 5680 1750 5690
rect 1650 5600 1660 5680
rect 1740 5600 1750 5680
rect 1650 5590 1750 5600
rect 1850 5680 1950 5690
rect 1850 5600 1860 5680
rect 1940 5600 1950 5680
rect 1850 5590 1950 5600
rect 2050 5680 2150 5690
rect 2050 5600 2060 5680
rect 2140 5600 2150 5680
rect 2050 5590 2150 5600
rect 2250 5680 2350 5690
rect 2250 5600 2260 5680
rect 2340 5600 2350 5680
rect 2250 5590 2350 5600
rect 2450 5680 2550 5690
rect 2450 5600 2460 5680
rect 2540 5600 2550 5680
rect 2450 5590 2550 5600
rect 2650 5680 2750 5690
rect 2650 5600 2660 5680
rect 2740 5600 2750 5680
rect 2650 5590 2750 5600
rect 2850 5680 2950 5690
rect 2850 5600 2860 5680
rect 2940 5600 2950 5680
rect 2850 5590 2950 5600
rect 3050 5680 3150 5690
rect 3050 5600 3060 5680
rect 3140 5600 3150 5680
rect 3050 5590 3150 5600
rect 3250 5680 3350 5690
rect 3250 5600 3260 5680
rect 3340 5600 3350 5680
rect 3250 5590 3350 5600
rect 3450 5680 3550 5690
rect 3450 5600 3460 5680
rect 3540 5600 3550 5680
rect 3450 5590 3550 5600
rect 3650 5680 3750 5690
rect 3650 5600 3660 5680
rect 3740 5600 3750 5680
rect 3650 5590 3750 5600
rect 3850 5680 3950 5690
rect 3850 5600 3860 5680
rect 3940 5600 3950 5680
rect 3850 5590 3950 5600
rect 4050 5680 4150 5690
rect 4050 5600 4060 5680
rect 4140 5600 4150 5680
rect 4050 5590 4150 5600
rect 4250 5680 4350 5690
rect 4250 5600 4260 5680
rect 4340 5600 4350 5680
rect 4250 5590 4350 5600
rect 4450 5680 4550 5690
rect 4450 5600 4460 5680
rect 4540 5600 4550 5680
rect 4450 5590 4550 5600
rect 4650 5680 4750 5690
rect 4650 5600 4660 5680
rect 4740 5600 4750 5680
rect 4650 5590 4750 5600
rect 4850 5680 4950 5690
rect 4850 5600 4860 5680
rect 4940 5600 4950 5680
rect 4850 5590 4950 5600
rect 5050 5680 5150 5690
rect 5050 5600 5060 5680
rect 5140 5600 5150 5680
rect 5050 5590 5150 5600
rect 5250 5680 5350 5690
rect 5250 5600 5260 5680
rect 5340 5600 5350 5680
rect 5250 5590 5350 5600
rect 5450 5680 5550 5690
rect 5450 5600 5460 5680
rect 5540 5600 5550 5680
rect 5450 5590 5550 5600
rect 5650 5680 5750 5690
rect 5650 5600 5660 5680
rect 5740 5600 5750 5680
rect 5650 5590 5750 5600
rect 5850 5680 5950 5690
rect 5850 5600 5860 5680
rect 5940 5600 5950 5680
rect 5850 5590 5950 5600
rect 6050 5680 6150 5690
rect 6050 5600 6060 5680
rect 6140 5600 6150 5680
rect 6050 5590 6150 5600
rect 6250 5680 6350 5690
rect 6250 5600 6260 5680
rect 6340 5600 6350 5680
rect 6250 5590 6350 5600
rect 6450 5680 6550 5690
rect 6450 5600 6460 5680
rect 6540 5600 6550 5680
rect 6450 5590 6550 5600
rect -150 5495 -50 5505
rect -150 5415 -140 5495
rect -60 5415 -50 5495
rect -150 5405 -50 5415
rect 50 5495 150 5505
rect 50 5415 60 5495
rect 140 5415 150 5495
rect 50 5405 150 5415
rect 250 5495 350 5505
rect 250 5415 260 5495
rect 340 5415 350 5495
rect 250 5405 350 5415
rect 450 5495 550 5505
rect 450 5415 460 5495
rect 540 5415 550 5495
rect 450 5405 550 5415
rect 650 5495 750 5505
rect 650 5415 660 5495
rect 740 5415 750 5495
rect 650 5405 750 5415
rect 850 5495 950 5505
rect 850 5415 860 5495
rect 940 5415 950 5495
rect 850 5405 950 5415
rect 1050 5495 1150 5505
rect 1050 5415 1060 5495
rect 1140 5415 1150 5495
rect 1050 5405 1150 5415
rect 1250 5495 1350 5505
rect 1250 5415 1260 5495
rect 1340 5415 1350 5495
rect 1250 5405 1350 5415
rect 1450 5495 1550 5505
rect 1450 5415 1460 5495
rect 1540 5415 1550 5495
rect 1450 5405 1550 5415
rect 1650 5495 1750 5505
rect 1650 5415 1660 5495
rect 1740 5415 1750 5495
rect 1650 5405 1750 5415
rect 1850 5495 1950 5505
rect 1850 5415 1860 5495
rect 1940 5415 1950 5495
rect 1850 5405 1950 5415
rect 2050 5495 2150 5505
rect 2050 5415 2060 5495
rect 2140 5415 2150 5495
rect 2050 5405 2150 5415
rect 2250 5495 2350 5505
rect 2250 5415 2260 5495
rect 2340 5415 2350 5495
rect 2250 5405 2350 5415
rect 2450 5495 2550 5505
rect 2450 5415 2460 5495
rect 2540 5415 2550 5495
rect 2450 5405 2550 5415
rect 2650 5495 2750 5505
rect 2650 5415 2660 5495
rect 2740 5415 2750 5495
rect 2650 5405 2750 5415
rect 2850 5495 2950 5505
rect 2850 5415 2860 5495
rect 2940 5415 2950 5495
rect 2850 5405 2950 5415
rect 3050 5495 3150 5505
rect 3050 5415 3060 5495
rect 3140 5415 3150 5495
rect 3050 5405 3150 5415
rect 3250 5495 3350 5505
rect 3250 5415 3260 5495
rect 3340 5415 3350 5495
rect 3250 5405 3350 5415
rect 3450 5495 3550 5505
rect 3450 5415 3460 5495
rect 3540 5415 3550 5495
rect 3450 5405 3550 5415
rect 3650 5495 3750 5505
rect 3650 5415 3660 5495
rect 3740 5415 3750 5495
rect 3650 5405 3750 5415
rect 3850 5495 3950 5505
rect 3850 5415 3860 5495
rect 3940 5415 3950 5495
rect 3850 5405 3950 5415
rect 4050 5495 4150 5505
rect 4050 5415 4060 5495
rect 4140 5415 4150 5495
rect 4050 5405 4150 5415
rect 4250 5495 4350 5505
rect 4250 5415 4260 5495
rect 4340 5415 4350 5495
rect 4250 5405 4350 5415
rect 4450 5495 4550 5505
rect 4450 5415 4460 5495
rect 4540 5415 4550 5495
rect 4450 5405 4550 5415
rect 4650 5495 4750 5505
rect 4650 5415 4660 5495
rect 4740 5415 4750 5495
rect 4650 5405 4750 5415
rect 4850 5495 4950 5505
rect 4850 5415 4860 5495
rect 4940 5415 4950 5495
rect 4850 5405 4950 5415
rect 5050 5495 5150 5505
rect 5050 5415 5060 5495
rect 5140 5415 5150 5495
rect 5050 5405 5150 5415
rect 5250 5495 5350 5505
rect 5250 5415 5260 5495
rect 5340 5415 5350 5495
rect 5250 5405 5350 5415
rect 5450 5495 5550 5505
rect 5450 5415 5460 5495
rect 5540 5415 5550 5495
rect 5450 5405 5550 5415
rect 5650 5495 5750 5505
rect 5650 5415 5660 5495
rect 5740 5415 5750 5495
rect 5650 5405 5750 5415
rect 5850 5495 5950 5505
rect 5850 5415 5860 5495
rect 5940 5415 5950 5495
rect 5850 5405 5950 5415
rect 6050 5495 6150 5505
rect 6050 5415 6060 5495
rect 6140 5415 6150 5495
rect 6050 5405 6150 5415
rect 6250 5495 6350 5505
rect 6250 5415 6260 5495
rect 6340 5415 6350 5495
rect 6250 5405 6350 5415
rect 6450 5495 6550 5505
rect 6450 5415 6460 5495
rect 6540 5415 6550 5495
rect 6450 5405 6550 5415
rect -150 5310 -50 5320
rect -150 5230 -140 5310
rect -60 5230 -50 5310
rect -150 5220 -50 5230
rect 50 5310 150 5320
rect 50 5230 60 5310
rect 140 5230 150 5310
rect 50 5220 150 5230
rect 250 5310 350 5320
rect 250 5230 260 5310
rect 340 5230 350 5310
rect 250 5220 350 5230
rect 450 5310 550 5320
rect 450 5230 460 5310
rect 540 5230 550 5310
rect 450 5220 550 5230
rect 650 5310 750 5320
rect 650 5230 660 5310
rect 740 5230 750 5310
rect 650 5220 750 5230
rect 850 5310 950 5320
rect 850 5230 860 5310
rect 940 5230 950 5310
rect 850 5220 950 5230
rect 1050 5310 1150 5320
rect 1050 5230 1060 5310
rect 1140 5230 1150 5310
rect 1050 5220 1150 5230
rect 1250 5310 1350 5320
rect 1250 5230 1260 5310
rect 1340 5230 1350 5310
rect 1250 5220 1350 5230
rect 1450 5310 1550 5320
rect 1450 5230 1460 5310
rect 1540 5230 1550 5310
rect 1450 5220 1550 5230
rect 1650 5310 1750 5320
rect 1650 5230 1660 5310
rect 1740 5230 1750 5310
rect 1650 5220 1750 5230
rect 1850 5310 1950 5320
rect 1850 5230 1860 5310
rect 1940 5230 1950 5310
rect 1850 5220 1950 5230
rect 2050 5310 2150 5320
rect 2050 5230 2060 5310
rect 2140 5230 2150 5310
rect 2050 5220 2150 5230
rect 2250 5310 2350 5320
rect 2250 5230 2260 5310
rect 2340 5230 2350 5310
rect 2250 5220 2350 5230
rect 2450 5310 2550 5320
rect 2450 5230 2460 5310
rect 2540 5230 2550 5310
rect 2450 5220 2550 5230
rect 2650 5310 2750 5320
rect 2650 5230 2660 5310
rect 2740 5230 2750 5310
rect 2650 5220 2750 5230
rect 2850 5310 2950 5320
rect 2850 5230 2860 5310
rect 2940 5230 2950 5310
rect 2850 5220 2950 5230
rect 3050 5310 3150 5320
rect 3050 5230 3060 5310
rect 3140 5230 3150 5310
rect 3050 5220 3150 5230
rect 3250 5310 3350 5320
rect 3250 5230 3260 5310
rect 3340 5230 3350 5310
rect 3250 5220 3350 5230
rect 3450 5310 3550 5320
rect 3450 5230 3460 5310
rect 3540 5230 3550 5310
rect 3450 5220 3550 5230
rect 3650 5310 3750 5320
rect 3650 5230 3660 5310
rect 3740 5230 3750 5310
rect 3650 5220 3750 5230
rect 3850 5310 3950 5320
rect 3850 5230 3860 5310
rect 3940 5230 3950 5310
rect 3850 5220 3950 5230
rect 4050 5310 4150 5320
rect 4050 5230 4060 5310
rect 4140 5230 4150 5310
rect 4050 5220 4150 5230
rect 4250 5310 4350 5320
rect 4250 5230 4260 5310
rect 4340 5230 4350 5310
rect 4250 5220 4350 5230
rect 4450 5310 4550 5320
rect 4450 5230 4460 5310
rect 4540 5230 4550 5310
rect 4450 5220 4550 5230
rect 4650 5310 4750 5320
rect 4650 5230 4660 5310
rect 4740 5230 4750 5310
rect 4650 5220 4750 5230
rect 4850 5310 4950 5320
rect 4850 5230 4860 5310
rect 4940 5230 4950 5310
rect 4850 5220 4950 5230
rect 5050 5310 5150 5320
rect 5050 5230 5060 5310
rect 5140 5230 5150 5310
rect 5050 5220 5150 5230
rect 5250 5310 5350 5320
rect 5250 5230 5260 5310
rect 5340 5230 5350 5310
rect 5250 5220 5350 5230
rect 5450 5310 5550 5320
rect 5450 5230 5460 5310
rect 5540 5230 5550 5310
rect 5450 5220 5550 5230
rect 5650 5310 5750 5320
rect 5650 5230 5660 5310
rect 5740 5230 5750 5310
rect 5650 5220 5750 5230
rect 5850 5310 5950 5320
rect 5850 5230 5860 5310
rect 5940 5230 5950 5310
rect 5850 5220 5950 5230
rect 6050 5310 6150 5320
rect 6050 5230 6060 5310
rect 6140 5230 6150 5310
rect 6050 5220 6150 5230
rect 6250 5310 6350 5320
rect 6250 5230 6260 5310
rect 6340 5230 6350 5310
rect 6250 5220 6350 5230
rect 6450 5310 6550 5320
rect 6450 5230 6460 5310
rect 6540 5230 6550 5310
rect 6450 5220 6550 5230
rect -150 5125 -50 5135
rect -150 5045 -140 5125
rect -60 5045 -50 5125
rect -150 5035 -50 5045
rect 50 5125 150 5135
rect 50 5045 60 5125
rect 140 5045 150 5125
rect 50 5035 150 5045
rect 250 5125 350 5135
rect 250 5045 260 5125
rect 340 5045 350 5125
rect 250 5035 350 5045
rect 450 5125 550 5135
rect 450 5045 460 5125
rect 540 5045 550 5125
rect 450 5035 550 5045
rect 650 5125 750 5135
rect 650 5045 660 5125
rect 740 5045 750 5125
rect 650 5035 750 5045
rect 850 5125 950 5135
rect 850 5045 860 5125
rect 940 5045 950 5125
rect 850 5035 950 5045
rect 1050 5125 1150 5135
rect 1050 5045 1060 5125
rect 1140 5045 1150 5125
rect 1050 5035 1150 5045
rect 1250 5125 1350 5135
rect 1250 5045 1260 5125
rect 1340 5045 1350 5125
rect 1250 5035 1350 5045
rect 1450 5125 1550 5135
rect 1450 5045 1460 5125
rect 1540 5045 1550 5125
rect 1450 5035 1550 5045
rect 1650 5125 1750 5135
rect 1650 5045 1660 5125
rect 1740 5045 1750 5125
rect 1650 5035 1750 5045
rect 1850 5125 1950 5135
rect 1850 5045 1860 5125
rect 1940 5045 1950 5125
rect 1850 5035 1950 5045
rect 2050 5125 2150 5135
rect 2050 5045 2060 5125
rect 2140 5045 2150 5125
rect 2050 5035 2150 5045
rect 2250 5125 2350 5135
rect 2250 5045 2260 5125
rect 2340 5045 2350 5125
rect 2250 5035 2350 5045
rect 2450 5125 2550 5135
rect 2450 5045 2460 5125
rect 2540 5045 2550 5125
rect 2450 5035 2550 5045
rect 2650 5125 2750 5135
rect 2650 5045 2660 5125
rect 2740 5045 2750 5125
rect 2650 5035 2750 5045
rect 2850 5125 2950 5135
rect 2850 5045 2860 5125
rect 2940 5045 2950 5125
rect 2850 5035 2950 5045
rect 3050 5125 3150 5135
rect 3050 5045 3060 5125
rect 3140 5045 3150 5125
rect 3050 5035 3150 5045
rect 3250 5125 3350 5135
rect 3250 5045 3260 5125
rect 3340 5045 3350 5125
rect 3250 5035 3350 5045
rect 3450 5125 3550 5135
rect 3450 5045 3460 5125
rect 3540 5045 3550 5125
rect 3450 5035 3550 5045
rect 3650 5125 3750 5135
rect 3650 5045 3660 5125
rect 3740 5045 3750 5125
rect 3650 5035 3750 5045
rect 3850 5125 3950 5135
rect 3850 5045 3860 5125
rect 3940 5045 3950 5125
rect 3850 5035 3950 5045
rect 4050 5125 4150 5135
rect 4050 5045 4060 5125
rect 4140 5045 4150 5125
rect 4050 5035 4150 5045
rect 4250 5125 4350 5135
rect 4250 5045 4260 5125
rect 4340 5045 4350 5125
rect 4250 5035 4350 5045
rect 4450 5125 4550 5135
rect 4450 5045 4460 5125
rect 4540 5045 4550 5125
rect 4450 5035 4550 5045
rect 4650 5125 4750 5135
rect 4650 5045 4660 5125
rect 4740 5045 4750 5125
rect 4650 5035 4750 5045
rect 4850 5125 4950 5135
rect 4850 5045 4860 5125
rect 4940 5045 4950 5125
rect 4850 5035 4950 5045
rect 5050 5125 5150 5135
rect 5050 5045 5060 5125
rect 5140 5045 5150 5125
rect 5050 5035 5150 5045
rect 5250 5125 5350 5135
rect 5250 5045 5260 5125
rect 5340 5045 5350 5125
rect 5250 5035 5350 5045
rect 5450 5125 5550 5135
rect 5450 5045 5460 5125
rect 5540 5045 5550 5125
rect 5450 5035 5550 5045
rect 5650 5125 5750 5135
rect 5650 5045 5660 5125
rect 5740 5045 5750 5125
rect 5650 5035 5750 5045
rect 5850 5125 5950 5135
rect 5850 5045 5860 5125
rect 5940 5045 5950 5125
rect 5850 5035 5950 5045
rect 6050 5125 6150 5135
rect 6050 5045 6060 5125
rect 6140 5045 6150 5125
rect 6050 5035 6150 5045
rect 6250 5125 6350 5135
rect 6250 5045 6260 5125
rect 6340 5045 6350 5125
rect 6250 5035 6350 5045
rect 6450 5125 6550 5135
rect 6450 5045 6460 5125
rect 6540 5045 6550 5125
rect 6450 5035 6550 5045
rect -150 4940 -50 4950
rect -150 4860 -140 4940
rect -60 4860 -50 4940
rect -150 4850 -50 4860
rect 50 4940 150 4950
rect 50 4860 60 4940
rect 140 4860 150 4940
rect 50 4850 150 4860
rect 250 4940 350 4950
rect 250 4860 260 4940
rect 340 4860 350 4940
rect 250 4850 350 4860
rect 450 4940 550 4950
rect 450 4860 460 4940
rect 540 4860 550 4940
rect 450 4850 550 4860
rect 650 4940 750 4950
rect 650 4860 660 4940
rect 740 4860 750 4940
rect 650 4850 750 4860
rect 850 4940 950 4950
rect 850 4860 860 4940
rect 940 4860 950 4940
rect 850 4850 950 4860
rect 1050 4940 1150 4950
rect 1050 4860 1060 4940
rect 1140 4860 1150 4940
rect 1050 4850 1150 4860
rect 1250 4940 1350 4950
rect 1250 4860 1260 4940
rect 1340 4860 1350 4940
rect 1250 4850 1350 4860
rect 1450 4940 1550 4950
rect 1450 4860 1460 4940
rect 1540 4860 1550 4940
rect 1450 4850 1550 4860
rect 1650 4940 1750 4950
rect 1650 4860 1660 4940
rect 1740 4860 1750 4940
rect 1650 4850 1750 4860
rect 1850 4940 1950 4950
rect 1850 4860 1860 4940
rect 1940 4860 1950 4940
rect 1850 4850 1950 4860
rect 2050 4940 2150 4950
rect 2050 4860 2060 4940
rect 2140 4860 2150 4940
rect 2050 4850 2150 4860
rect 2250 4940 2350 4950
rect 2250 4860 2260 4940
rect 2340 4860 2350 4940
rect 2250 4850 2350 4860
rect 2450 4940 2550 4950
rect 2450 4860 2460 4940
rect 2540 4860 2550 4940
rect 2450 4850 2550 4860
rect 2650 4940 2750 4950
rect 2650 4860 2660 4940
rect 2740 4860 2750 4940
rect 2650 4850 2750 4860
rect 2850 4940 2950 4950
rect 2850 4860 2860 4940
rect 2940 4860 2950 4940
rect 2850 4850 2950 4860
rect 3050 4940 3150 4950
rect 3050 4860 3060 4940
rect 3140 4860 3150 4940
rect 3050 4850 3150 4860
rect 3250 4940 3350 4950
rect 3250 4860 3260 4940
rect 3340 4860 3350 4940
rect 3250 4850 3350 4860
rect 3450 4940 3550 4950
rect 3450 4860 3460 4940
rect 3540 4860 3550 4940
rect 3450 4850 3550 4860
rect 3650 4940 3750 4950
rect 3650 4860 3660 4940
rect 3740 4860 3750 4940
rect 3650 4850 3750 4860
rect 3850 4940 3950 4950
rect 3850 4860 3860 4940
rect 3940 4860 3950 4940
rect 3850 4850 3950 4860
rect 4050 4940 4150 4950
rect 4050 4860 4060 4940
rect 4140 4860 4150 4940
rect 4050 4850 4150 4860
rect 4250 4940 4350 4950
rect 4250 4860 4260 4940
rect 4340 4860 4350 4940
rect 4250 4850 4350 4860
rect 4450 4940 4550 4950
rect 4450 4860 4460 4940
rect 4540 4860 4550 4940
rect 4450 4850 4550 4860
rect 4650 4940 4750 4950
rect 4650 4860 4660 4940
rect 4740 4860 4750 4940
rect 4650 4850 4750 4860
rect 4850 4940 4950 4950
rect 4850 4860 4860 4940
rect 4940 4860 4950 4940
rect 4850 4850 4950 4860
rect 5050 4940 5150 4950
rect 5050 4860 5060 4940
rect 5140 4860 5150 4940
rect 5050 4850 5150 4860
rect 5250 4940 5350 4950
rect 5250 4860 5260 4940
rect 5340 4860 5350 4940
rect 5250 4850 5350 4860
rect 5450 4940 5550 4950
rect 5450 4860 5460 4940
rect 5540 4860 5550 4940
rect 5450 4850 5550 4860
rect 5650 4940 5750 4950
rect 5650 4860 5660 4940
rect 5740 4860 5750 4940
rect 5650 4850 5750 4860
rect 5850 4940 5950 4950
rect 5850 4860 5860 4940
rect 5940 4860 5950 4940
rect 5850 4850 5950 4860
rect 6050 4940 6150 4950
rect 6050 4860 6060 4940
rect 6140 4860 6150 4940
rect 6050 4850 6150 4860
rect 6250 4940 6350 4950
rect 6250 4860 6260 4940
rect 6340 4860 6350 4940
rect 6250 4850 6350 4860
rect 6450 4940 6550 4950
rect 6450 4860 6460 4940
rect 6540 4860 6550 4940
rect 6450 4850 6550 4860
rect -150 4755 -50 4765
rect -150 4675 -140 4755
rect -60 4675 -50 4755
rect -150 4665 -50 4675
rect 50 4755 150 4765
rect 50 4675 60 4755
rect 140 4675 150 4755
rect 50 4665 150 4675
rect 250 4755 350 4765
rect 250 4675 260 4755
rect 340 4675 350 4755
rect 250 4665 350 4675
rect 450 4755 550 4765
rect 450 4675 460 4755
rect 540 4675 550 4755
rect 450 4665 550 4675
rect 650 4755 750 4765
rect 650 4675 660 4755
rect 740 4675 750 4755
rect 650 4665 750 4675
rect 850 4755 950 4765
rect 850 4675 860 4755
rect 940 4675 950 4755
rect 850 4665 950 4675
rect 1050 4755 1150 4765
rect 1050 4675 1060 4755
rect 1140 4675 1150 4755
rect 1050 4665 1150 4675
rect 1250 4755 1350 4765
rect 1250 4675 1260 4755
rect 1340 4675 1350 4755
rect 1250 4665 1350 4675
rect 1450 4755 1550 4765
rect 1450 4675 1460 4755
rect 1540 4675 1550 4755
rect 1450 4665 1550 4675
rect 1650 4755 1750 4765
rect 1650 4675 1660 4755
rect 1740 4675 1750 4755
rect 1650 4665 1750 4675
rect 1850 4755 1950 4765
rect 1850 4675 1860 4755
rect 1940 4675 1950 4755
rect 1850 4665 1950 4675
rect 2050 4755 2150 4765
rect 2050 4675 2060 4755
rect 2140 4675 2150 4755
rect 2050 4665 2150 4675
rect 2250 4755 2350 4765
rect 2250 4675 2260 4755
rect 2340 4675 2350 4755
rect 2250 4665 2350 4675
rect 2450 4755 2550 4765
rect 2450 4675 2460 4755
rect 2540 4675 2550 4755
rect 2450 4665 2550 4675
rect 2650 4755 2750 4765
rect 2650 4675 2660 4755
rect 2740 4675 2750 4755
rect 2650 4665 2750 4675
rect 2850 4755 2950 4765
rect 2850 4675 2860 4755
rect 2940 4675 2950 4755
rect 2850 4665 2950 4675
rect 3050 4755 3150 4765
rect 3050 4675 3060 4755
rect 3140 4675 3150 4755
rect 3050 4665 3150 4675
rect 3250 4755 3350 4765
rect 3250 4675 3260 4755
rect 3340 4675 3350 4755
rect 3250 4665 3350 4675
rect 3450 4755 3550 4765
rect 3450 4675 3460 4755
rect 3540 4675 3550 4755
rect 3450 4665 3550 4675
rect 3650 4755 3750 4765
rect 3650 4675 3660 4755
rect 3740 4675 3750 4755
rect 3650 4665 3750 4675
rect 3850 4755 3950 4765
rect 3850 4675 3860 4755
rect 3940 4675 3950 4755
rect 3850 4665 3950 4675
rect 4050 4755 4150 4765
rect 4050 4675 4060 4755
rect 4140 4675 4150 4755
rect 4050 4665 4150 4675
rect 4250 4755 4350 4765
rect 4250 4675 4260 4755
rect 4340 4675 4350 4755
rect 4250 4665 4350 4675
rect 4450 4755 4550 4765
rect 4450 4675 4460 4755
rect 4540 4675 4550 4755
rect 4450 4665 4550 4675
rect 4650 4755 4750 4765
rect 4650 4675 4660 4755
rect 4740 4675 4750 4755
rect 4650 4665 4750 4675
rect 4850 4755 4950 4765
rect 4850 4675 4860 4755
rect 4940 4675 4950 4755
rect 4850 4665 4950 4675
rect 5050 4755 5150 4765
rect 5050 4675 5060 4755
rect 5140 4675 5150 4755
rect 5050 4665 5150 4675
rect 5250 4755 5350 4765
rect 5250 4675 5260 4755
rect 5340 4675 5350 4755
rect 5250 4665 5350 4675
rect 5450 4755 5550 4765
rect 5450 4675 5460 4755
rect 5540 4675 5550 4755
rect 5450 4665 5550 4675
rect 5650 4755 5750 4765
rect 5650 4675 5660 4755
rect 5740 4675 5750 4755
rect 5650 4665 5750 4675
rect 5850 4755 5950 4765
rect 5850 4675 5860 4755
rect 5940 4675 5950 4755
rect 5850 4665 5950 4675
rect 6050 4755 6150 4765
rect 6050 4675 6060 4755
rect 6140 4675 6150 4755
rect 6050 4665 6150 4675
rect 6250 4755 6350 4765
rect 6250 4675 6260 4755
rect 6340 4675 6350 4755
rect 6250 4665 6350 4675
rect 6450 4755 6550 4765
rect 6450 4675 6460 4755
rect 6540 4675 6550 4755
rect 6450 4665 6550 4675
rect -150 4570 -50 4580
rect -150 4490 -140 4570
rect -60 4490 -50 4570
rect -150 4480 -50 4490
rect 50 4570 150 4580
rect 50 4490 60 4570
rect 140 4490 150 4570
rect 50 4480 150 4490
rect 250 4570 350 4580
rect 250 4490 260 4570
rect 340 4490 350 4570
rect 250 4480 350 4490
rect 450 4570 550 4580
rect 450 4490 460 4570
rect 540 4490 550 4570
rect 450 4480 550 4490
rect 650 4570 750 4580
rect 650 4490 660 4570
rect 740 4490 750 4570
rect 650 4480 750 4490
rect 850 4570 950 4580
rect 850 4490 860 4570
rect 940 4490 950 4570
rect 850 4480 950 4490
rect 1050 4570 1150 4580
rect 1050 4490 1060 4570
rect 1140 4490 1150 4570
rect 1050 4480 1150 4490
rect 1250 4570 1350 4580
rect 1250 4490 1260 4570
rect 1340 4490 1350 4570
rect 1250 4480 1350 4490
rect 1450 4570 1550 4580
rect 1450 4490 1460 4570
rect 1540 4490 1550 4570
rect 1450 4480 1550 4490
rect 1650 4570 1750 4580
rect 1650 4490 1660 4570
rect 1740 4490 1750 4570
rect 1650 4480 1750 4490
rect 1850 4570 1950 4580
rect 1850 4490 1860 4570
rect 1940 4490 1950 4570
rect 1850 4480 1950 4490
rect 2050 4570 2150 4580
rect 2050 4490 2060 4570
rect 2140 4490 2150 4570
rect 2050 4480 2150 4490
rect 2250 4570 2350 4580
rect 2250 4490 2260 4570
rect 2340 4490 2350 4570
rect 2250 4480 2350 4490
rect 2450 4570 2550 4580
rect 2450 4490 2460 4570
rect 2540 4490 2550 4570
rect 2450 4480 2550 4490
rect 2650 4570 2750 4580
rect 2650 4490 2660 4570
rect 2740 4490 2750 4570
rect 2650 4480 2750 4490
rect 2850 4570 2950 4580
rect 2850 4490 2860 4570
rect 2940 4490 2950 4570
rect 2850 4480 2950 4490
rect 3050 4570 3150 4580
rect 3050 4490 3060 4570
rect 3140 4490 3150 4570
rect 3050 4480 3150 4490
rect 3250 4570 3350 4580
rect 3250 4490 3260 4570
rect 3340 4490 3350 4570
rect 3250 4480 3350 4490
rect 3450 4570 3550 4580
rect 3450 4490 3460 4570
rect 3540 4490 3550 4570
rect 3450 4480 3550 4490
rect 3650 4570 3750 4580
rect 3650 4490 3660 4570
rect 3740 4490 3750 4570
rect 3650 4480 3750 4490
rect 3850 4570 3950 4580
rect 3850 4490 3860 4570
rect 3940 4490 3950 4570
rect 3850 4480 3950 4490
rect 4050 4570 4150 4580
rect 4050 4490 4060 4570
rect 4140 4490 4150 4570
rect 4050 4480 4150 4490
rect 4250 4570 4350 4580
rect 4250 4490 4260 4570
rect 4340 4490 4350 4570
rect 4250 4480 4350 4490
rect 4450 4570 4550 4580
rect 4450 4490 4460 4570
rect 4540 4490 4550 4570
rect 4450 4480 4550 4490
rect 4650 4570 4750 4580
rect 4650 4490 4660 4570
rect 4740 4490 4750 4570
rect 4650 4480 4750 4490
rect 4850 4570 4950 4580
rect 4850 4490 4860 4570
rect 4940 4490 4950 4570
rect 4850 4480 4950 4490
rect 5050 4570 5150 4580
rect 5050 4490 5060 4570
rect 5140 4490 5150 4570
rect 5050 4480 5150 4490
rect 5250 4570 5350 4580
rect 5250 4490 5260 4570
rect 5340 4490 5350 4570
rect 5250 4480 5350 4490
rect 5450 4570 5550 4580
rect 5450 4490 5460 4570
rect 5540 4490 5550 4570
rect 5450 4480 5550 4490
rect 5650 4570 5750 4580
rect 5650 4490 5660 4570
rect 5740 4490 5750 4570
rect 5650 4480 5750 4490
rect 5850 4570 5950 4580
rect 5850 4490 5860 4570
rect 5940 4490 5950 4570
rect 5850 4480 5950 4490
rect 6050 4570 6150 4580
rect 6050 4490 6060 4570
rect 6140 4490 6150 4570
rect 6050 4480 6150 4490
rect 6250 4570 6350 4580
rect 6250 4490 6260 4570
rect 6340 4490 6350 4570
rect 6250 4480 6350 4490
rect 6450 4570 6550 4580
rect 6450 4490 6460 4570
rect 6540 4490 6550 4570
rect 6450 4480 6550 4490
rect -150 4385 -50 4395
rect -150 4305 -140 4385
rect -60 4305 -50 4385
rect -150 4295 -50 4305
rect 50 4385 150 4395
rect 50 4305 60 4385
rect 140 4305 150 4385
rect 50 4295 150 4305
rect 250 4385 350 4395
rect 250 4305 260 4385
rect 340 4305 350 4385
rect 250 4295 350 4305
rect 450 4385 550 4395
rect 450 4305 460 4385
rect 540 4305 550 4385
rect 450 4295 550 4305
rect 650 4385 750 4395
rect 650 4305 660 4385
rect 740 4305 750 4385
rect 650 4295 750 4305
rect 850 4385 950 4395
rect 850 4305 860 4385
rect 940 4305 950 4385
rect 850 4295 950 4305
rect 1050 4385 1150 4395
rect 1050 4305 1060 4385
rect 1140 4305 1150 4385
rect 1050 4295 1150 4305
rect 1250 4385 1350 4395
rect 1250 4305 1260 4385
rect 1340 4305 1350 4385
rect 1250 4295 1350 4305
rect 1450 4385 1550 4395
rect 1450 4305 1460 4385
rect 1540 4305 1550 4385
rect 1450 4295 1550 4305
rect 1650 4385 1750 4395
rect 1650 4305 1660 4385
rect 1740 4305 1750 4385
rect 1650 4295 1750 4305
rect 1850 4385 1950 4395
rect 1850 4305 1860 4385
rect 1940 4305 1950 4385
rect 1850 4295 1950 4305
rect 2050 4385 2150 4395
rect 2050 4305 2060 4385
rect 2140 4305 2150 4385
rect 2050 4295 2150 4305
rect 2250 4385 2350 4395
rect 2250 4305 2260 4385
rect 2340 4305 2350 4385
rect 2250 4295 2350 4305
rect 2450 4385 2550 4395
rect 2450 4305 2460 4385
rect 2540 4305 2550 4385
rect 2450 4295 2550 4305
rect 2650 4385 2750 4395
rect 2650 4305 2660 4385
rect 2740 4305 2750 4385
rect 2650 4295 2750 4305
rect 2850 4385 2950 4395
rect 2850 4305 2860 4385
rect 2940 4305 2950 4385
rect 2850 4295 2950 4305
rect 3050 4385 3150 4395
rect 3050 4305 3060 4385
rect 3140 4305 3150 4385
rect 3050 4295 3150 4305
rect 3250 4385 3350 4395
rect 3250 4305 3260 4385
rect 3340 4305 3350 4385
rect 3250 4295 3350 4305
rect 3450 4385 3550 4395
rect 3450 4305 3460 4385
rect 3540 4305 3550 4385
rect 3450 4295 3550 4305
rect 3650 4385 3750 4395
rect 3650 4305 3660 4385
rect 3740 4305 3750 4385
rect 3650 4295 3750 4305
rect 3850 4385 3950 4395
rect 3850 4305 3860 4385
rect 3940 4305 3950 4385
rect 3850 4295 3950 4305
rect 4050 4385 4150 4395
rect 4050 4305 4060 4385
rect 4140 4305 4150 4385
rect 4050 4295 4150 4305
rect 4250 4385 4350 4395
rect 4250 4305 4260 4385
rect 4340 4305 4350 4385
rect 4250 4295 4350 4305
rect 4450 4385 4550 4395
rect 4450 4305 4460 4385
rect 4540 4305 4550 4385
rect 4450 4295 4550 4305
rect 4650 4385 4750 4395
rect 4650 4305 4660 4385
rect 4740 4305 4750 4385
rect 4650 4295 4750 4305
rect 4850 4385 4950 4395
rect 4850 4305 4860 4385
rect 4940 4305 4950 4385
rect 4850 4295 4950 4305
rect 5050 4385 5150 4395
rect 5050 4305 5060 4385
rect 5140 4305 5150 4385
rect 5050 4295 5150 4305
rect 5250 4385 5350 4395
rect 5250 4305 5260 4385
rect 5340 4305 5350 4385
rect 5250 4295 5350 4305
rect 5450 4385 5550 4395
rect 5450 4305 5460 4385
rect 5540 4305 5550 4385
rect 5450 4295 5550 4305
rect 5650 4385 5750 4395
rect 5650 4305 5660 4385
rect 5740 4305 5750 4385
rect 5650 4295 5750 4305
rect 5850 4385 5950 4395
rect 5850 4305 5860 4385
rect 5940 4305 5950 4385
rect 5850 4295 5950 4305
rect 6050 4385 6150 4395
rect 6050 4305 6060 4385
rect 6140 4305 6150 4385
rect 6050 4295 6150 4305
rect 6250 4385 6350 4395
rect 6250 4305 6260 4385
rect 6340 4305 6350 4385
rect 6250 4295 6350 4305
rect 6450 4385 6550 4395
rect 6450 4305 6460 4385
rect 6540 4305 6550 4385
rect 6450 4295 6550 4305
rect -150 4200 -50 4210
rect -150 4120 -140 4200
rect -60 4120 -50 4200
rect -150 4110 -50 4120
rect 50 4200 150 4210
rect 50 4120 60 4200
rect 140 4120 150 4200
rect 50 4110 150 4120
rect 250 4200 350 4210
rect 250 4120 260 4200
rect 340 4120 350 4200
rect 250 4110 350 4120
rect 450 4200 550 4210
rect 450 4120 460 4200
rect 540 4120 550 4200
rect 450 4110 550 4120
rect 650 4200 750 4210
rect 650 4120 660 4200
rect 740 4120 750 4200
rect 650 4110 750 4120
rect 850 4200 950 4210
rect 850 4120 860 4200
rect 940 4120 950 4200
rect 850 4110 950 4120
rect 1050 4200 1150 4210
rect 1050 4120 1060 4200
rect 1140 4120 1150 4200
rect 1050 4110 1150 4120
rect 1250 4200 1350 4210
rect 1250 4120 1260 4200
rect 1340 4120 1350 4200
rect 1250 4110 1350 4120
rect 1450 4200 1550 4210
rect 1450 4120 1460 4200
rect 1540 4120 1550 4200
rect 1450 4110 1550 4120
rect 1650 4200 1750 4210
rect 1650 4120 1660 4200
rect 1740 4120 1750 4200
rect 1650 4110 1750 4120
rect 1850 4200 1950 4210
rect 1850 4120 1860 4200
rect 1940 4120 1950 4200
rect 1850 4110 1950 4120
rect 2050 4200 2150 4210
rect 2050 4120 2060 4200
rect 2140 4120 2150 4200
rect 2050 4110 2150 4120
rect 2250 4200 2350 4210
rect 2250 4120 2260 4200
rect 2340 4120 2350 4200
rect 2250 4110 2350 4120
rect 2450 4200 2550 4210
rect 2450 4120 2460 4200
rect 2540 4120 2550 4200
rect 2450 4110 2550 4120
rect 2650 4200 2750 4210
rect 2650 4120 2660 4200
rect 2740 4120 2750 4200
rect 2650 4110 2750 4120
rect 2850 4200 2950 4210
rect 2850 4120 2860 4200
rect 2940 4120 2950 4200
rect 2850 4110 2950 4120
rect 3050 4200 3150 4210
rect 3050 4120 3060 4200
rect 3140 4120 3150 4200
rect 3050 4110 3150 4120
rect 3250 4200 3350 4210
rect 3250 4120 3260 4200
rect 3340 4120 3350 4200
rect 3250 4110 3350 4120
rect 3450 4200 3550 4210
rect 3450 4120 3460 4200
rect 3540 4120 3550 4200
rect 3450 4110 3550 4120
rect 3650 4200 3750 4210
rect 3650 4120 3660 4200
rect 3740 4120 3750 4200
rect 3650 4110 3750 4120
rect 3850 4200 3950 4210
rect 3850 4120 3860 4200
rect 3940 4120 3950 4200
rect 3850 4110 3950 4120
rect 4050 4200 4150 4210
rect 4050 4120 4060 4200
rect 4140 4120 4150 4200
rect 4050 4110 4150 4120
rect 4250 4200 4350 4210
rect 4250 4120 4260 4200
rect 4340 4120 4350 4200
rect 4250 4110 4350 4120
rect 4450 4200 4550 4210
rect 4450 4120 4460 4200
rect 4540 4120 4550 4200
rect 4450 4110 4550 4120
rect 4650 4200 4750 4210
rect 4650 4120 4660 4200
rect 4740 4120 4750 4200
rect 4650 4110 4750 4120
rect 4850 4200 4950 4210
rect 4850 4120 4860 4200
rect 4940 4120 4950 4200
rect 4850 4110 4950 4120
rect 5050 4200 5150 4210
rect 5050 4120 5060 4200
rect 5140 4120 5150 4200
rect 5050 4110 5150 4120
rect 5250 4200 5350 4210
rect 5250 4120 5260 4200
rect 5340 4120 5350 4200
rect 5250 4110 5350 4120
rect 5450 4200 5550 4210
rect 5450 4120 5460 4200
rect 5540 4120 5550 4200
rect 5450 4110 5550 4120
rect 5650 4200 5750 4210
rect 5650 4120 5660 4200
rect 5740 4120 5750 4200
rect 5650 4110 5750 4120
rect 5850 4200 5950 4210
rect 5850 4120 5860 4200
rect 5940 4120 5950 4200
rect 5850 4110 5950 4120
rect 6050 4200 6150 4210
rect 6050 4120 6060 4200
rect 6140 4120 6150 4200
rect 6050 4110 6150 4120
rect 6250 4200 6350 4210
rect 6250 4120 6260 4200
rect 6340 4120 6350 4200
rect 6250 4110 6350 4120
rect 6450 4200 6550 4210
rect 6450 4120 6460 4200
rect 6540 4120 6550 4200
rect 6450 4110 6550 4120
rect -150 4015 -50 4025
rect -150 3935 -140 4015
rect -60 3935 -50 4015
rect -150 3925 -50 3935
rect 50 4015 150 4025
rect 50 3935 60 4015
rect 140 3935 150 4015
rect 50 3925 150 3935
rect 250 4015 350 4025
rect 250 3935 260 4015
rect 340 3935 350 4015
rect 250 3925 350 3935
rect 450 4015 550 4025
rect 450 3935 460 4015
rect 540 3935 550 4015
rect 450 3925 550 3935
rect 650 4015 750 4025
rect 650 3935 660 4015
rect 740 3935 750 4015
rect 650 3925 750 3935
rect 850 4015 950 4025
rect 850 3935 860 4015
rect 940 3935 950 4015
rect 850 3925 950 3935
rect 1050 4015 1150 4025
rect 1050 3935 1060 4015
rect 1140 3935 1150 4015
rect 1050 3925 1150 3935
rect 1250 4015 1350 4025
rect 1250 3935 1260 4015
rect 1340 3935 1350 4015
rect 1250 3925 1350 3935
rect 1450 4015 1550 4025
rect 1450 3935 1460 4015
rect 1540 3935 1550 4015
rect 1450 3925 1550 3935
rect 1650 4015 1750 4025
rect 1650 3935 1660 4015
rect 1740 3935 1750 4015
rect 1650 3925 1750 3935
rect 1850 4015 1950 4025
rect 1850 3935 1860 4015
rect 1940 3935 1950 4015
rect 1850 3925 1950 3935
rect 2050 4015 2150 4025
rect 2050 3935 2060 4015
rect 2140 3935 2150 4015
rect 2050 3925 2150 3935
rect 2250 4015 2350 4025
rect 2250 3935 2260 4015
rect 2340 3935 2350 4015
rect 2250 3925 2350 3935
rect 2450 4015 2550 4025
rect 2450 3935 2460 4015
rect 2540 3935 2550 4015
rect 2450 3925 2550 3935
rect 2650 4015 2750 4025
rect 2650 3935 2660 4015
rect 2740 3935 2750 4015
rect 2650 3925 2750 3935
rect 2850 4015 2950 4025
rect 2850 3935 2860 4015
rect 2940 3935 2950 4015
rect 2850 3925 2950 3935
rect 3050 4015 3150 4025
rect 3050 3935 3060 4015
rect 3140 3935 3150 4015
rect 3050 3925 3150 3935
rect 3250 4015 3350 4025
rect 3250 3935 3260 4015
rect 3340 3935 3350 4015
rect 3250 3925 3350 3935
rect 3450 4015 3550 4025
rect 3450 3935 3460 4015
rect 3540 3935 3550 4015
rect 3450 3925 3550 3935
rect 3650 4015 3750 4025
rect 3650 3935 3660 4015
rect 3740 3935 3750 4015
rect 3650 3925 3750 3935
rect 3850 4015 3950 4025
rect 3850 3935 3860 4015
rect 3940 3935 3950 4015
rect 3850 3925 3950 3935
rect 4050 4015 4150 4025
rect 4050 3935 4060 4015
rect 4140 3935 4150 4015
rect 4050 3925 4150 3935
rect 4250 4015 4350 4025
rect 4250 3935 4260 4015
rect 4340 3935 4350 4015
rect 4250 3925 4350 3935
rect 4450 4015 4550 4025
rect 4450 3935 4460 4015
rect 4540 3935 4550 4015
rect 4450 3925 4550 3935
rect 4650 4015 4750 4025
rect 4650 3935 4660 4015
rect 4740 3935 4750 4015
rect 4650 3925 4750 3935
rect 4850 4015 4950 4025
rect 4850 3935 4860 4015
rect 4940 3935 4950 4015
rect 4850 3925 4950 3935
rect 5050 4015 5150 4025
rect 5050 3935 5060 4015
rect 5140 3935 5150 4015
rect 5050 3925 5150 3935
rect 5250 4015 5350 4025
rect 5250 3935 5260 4015
rect 5340 3935 5350 4015
rect 5250 3925 5350 3935
rect 5450 4015 5550 4025
rect 5450 3935 5460 4015
rect 5540 3935 5550 4015
rect 5450 3925 5550 3935
rect 5650 4015 5750 4025
rect 5650 3935 5660 4015
rect 5740 3935 5750 4015
rect 5650 3925 5750 3935
rect 5850 4015 5950 4025
rect 5850 3935 5860 4015
rect 5940 3935 5950 4015
rect 5850 3925 5950 3935
rect 6050 4015 6150 4025
rect 6050 3935 6060 4015
rect 6140 3935 6150 4015
rect 6050 3925 6150 3935
rect 6250 4015 6350 4025
rect 6250 3935 6260 4015
rect 6340 3935 6350 4015
rect 6250 3925 6350 3935
rect 6450 4015 6550 4025
rect 6450 3935 6460 4015
rect 6540 3935 6550 4015
rect 6450 3925 6550 3935
rect -150 3830 -50 3840
rect -150 3750 -140 3830
rect -60 3750 -50 3830
rect -150 3740 -50 3750
rect 50 3830 150 3840
rect 50 3750 60 3830
rect 140 3750 150 3830
rect 50 3740 150 3750
rect 250 3830 350 3840
rect 250 3750 260 3830
rect 340 3750 350 3830
rect 250 3740 350 3750
rect 450 3830 550 3840
rect 450 3750 460 3830
rect 540 3750 550 3830
rect 450 3740 550 3750
rect 650 3830 750 3840
rect 650 3750 660 3830
rect 740 3750 750 3830
rect 650 3740 750 3750
rect 850 3830 950 3840
rect 850 3750 860 3830
rect 940 3750 950 3830
rect 850 3740 950 3750
rect 1050 3830 1150 3840
rect 1050 3750 1060 3830
rect 1140 3750 1150 3830
rect 1050 3740 1150 3750
rect 1250 3830 1350 3840
rect 1250 3750 1260 3830
rect 1340 3750 1350 3830
rect 1250 3740 1350 3750
rect 1450 3830 1550 3840
rect 1450 3750 1460 3830
rect 1540 3750 1550 3830
rect 1450 3740 1550 3750
rect 1650 3830 1750 3840
rect 1650 3750 1660 3830
rect 1740 3750 1750 3830
rect 1650 3740 1750 3750
rect 1850 3830 1950 3840
rect 1850 3750 1860 3830
rect 1940 3750 1950 3830
rect 1850 3740 1950 3750
rect 2050 3830 2150 3840
rect 2050 3750 2060 3830
rect 2140 3750 2150 3830
rect 2050 3740 2150 3750
rect 2250 3830 2350 3840
rect 2250 3750 2260 3830
rect 2340 3750 2350 3830
rect 2250 3740 2350 3750
rect 2450 3830 2550 3840
rect 2450 3750 2460 3830
rect 2540 3750 2550 3830
rect 2450 3740 2550 3750
rect 2650 3830 2750 3840
rect 2650 3750 2660 3830
rect 2740 3750 2750 3830
rect 2650 3740 2750 3750
rect 2850 3830 2950 3840
rect 2850 3750 2860 3830
rect 2940 3750 2950 3830
rect 2850 3740 2950 3750
rect 3050 3830 3150 3840
rect 3050 3750 3060 3830
rect 3140 3750 3150 3830
rect 3050 3740 3150 3750
rect 3250 3830 3350 3840
rect 3250 3750 3260 3830
rect 3340 3750 3350 3830
rect 3250 3740 3350 3750
rect 3450 3830 3550 3840
rect 3450 3750 3460 3830
rect 3540 3750 3550 3830
rect 3450 3740 3550 3750
rect 3650 3830 3750 3840
rect 3650 3750 3660 3830
rect 3740 3750 3750 3830
rect 3650 3740 3750 3750
rect 3850 3830 3950 3840
rect 3850 3750 3860 3830
rect 3940 3750 3950 3830
rect 3850 3740 3950 3750
rect 4050 3830 4150 3840
rect 4050 3750 4060 3830
rect 4140 3750 4150 3830
rect 4050 3740 4150 3750
rect 4250 3830 4350 3840
rect 4250 3750 4260 3830
rect 4340 3750 4350 3830
rect 4250 3740 4350 3750
rect 4450 3830 4550 3840
rect 4450 3750 4460 3830
rect 4540 3750 4550 3830
rect 4450 3740 4550 3750
rect 4650 3830 4750 3840
rect 4650 3750 4660 3830
rect 4740 3750 4750 3830
rect 4650 3740 4750 3750
rect 4850 3830 4950 3840
rect 4850 3750 4860 3830
rect 4940 3750 4950 3830
rect 4850 3740 4950 3750
rect 5050 3830 5150 3840
rect 5050 3750 5060 3830
rect 5140 3750 5150 3830
rect 5050 3740 5150 3750
rect 5250 3830 5350 3840
rect 5250 3750 5260 3830
rect 5340 3750 5350 3830
rect 5250 3740 5350 3750
rect 5450 3830 5550 3840
rect 5450 3750 5460 3830
rect 5540 3750 5550 3830
rect 5450 3740 5550 3750
rect 5650 3830 5750 3840
rect 5650 3750 5660 3830
rect 5740 3750 5750 3830
rect 5650 3740 5750 3750
rect 5850 3830 5950 3840
rect 5850 3750 5860 3830
rect 5940 3750 5950 3830
rect 5850 3740 5950 3750
rect 6050 3830 6150 3840
rect 6050 3750 6060 3830
rect 6140 3750 6150 3830
rect 6050 3740 6150 3750
rect 6250 3830 6350 3840
rect 6250 3750 6260 3830
rect 6340 3750 6350 3830
rect 6250 3740 6350 3750
rect 6450 3830 6550 3840
rect 6450 3750 6460 3830
rect 6540 3750 6550 3830
rect 6450 3740 6550 3750
rect -150 3645 -50 3655
rect -150 3565 -140 3645
rect -60 3565 -50 3645
rect -150 3555 -50 3565
rect 50 3645 150 3655
rect 50 3565 60 3645
rect 140 3565 150 3645
rect 50 3555 150 3565
rect 250 3645 350 3655
rect 250 3565 260 3645
rect 340 3565 350 3645
rect 250 3555 350 3565
rect 450 3645 550 3655
rect 450 3565 460 3645
rect 540 3565 550 3645
rect 450 3555 550 3565
rect 650 3645 750 3655
rect 650 3565 660 3645
rect 740 3565 750 3645
rect 650 3555 750 3565
rect 850 3645 950 3655
rect 850 3565 860 3645
rect 940 3565 950 3645
rect 850 3555 950 3565
rect 1050 3645 1150 3655
rect 1050 3565 1060 3645
rect 1140 3565 1150 3645
rect 1050 3555 1150 3565
rect 1250 3645 1350 3655
rect 1250 3565 1260 3645
rect 1340 3565 1350 3645
rect 1250 3555 1350 3565
rect 1450 3645 1550 3655
rect 1450 3565 1460 3645
rect 1540 3565 1550 3645
rect 1450 3555 1550 3565
rect 1650 3645 1750 3655
rect 1650 3565 1660 3645
rect 1740 3565 1750 3645
rect 1650 3555 1750 3565
rect 1850 3645 1950 3655
rect 1850 3565 1860 3645
rect 1940 3565 1950 3645
rect 1850 3555 1950 3565
rect 2050 3645 2150 3655
rect 2050 3565 2060 3645
rect 2140 3565 2150 3645
rect 2050 3555 2150 3565
rect 2250 3645 2350 3655
rect 2250 3565 2260 3645
rect 2340 3565 2350 3645
rect 2250 3555 2350 3565
rect 2450 3645 2550 3655
rect 2450 3565 2460 3645
rect 2540 3565 2550 3645
rect 2450 3555 2550 3565
rect 2650 3645 2750 3655
rect 2650 3565 2660 3645
rect 2740 3565 2750 3645
rect 2650 3555 2750 3565
rect 2850 3645 2950 3655
rect 2850 3565 2860 3645
rect 2940 3565 2950 3645
rect 2850 3555 2950 3565
rect 3050 3645 3150 3655
rect 3050 3565 3060 3645
rect 3140 3565 3150 3645
rect 3050 3555 3150 3565
rect 3250 3645 3350 3655
rect 3250 3565 3260 3645
rect 3340 3565 3350 3645
rect 3250 3555 3350 3565
rect 3450 3645 3550 3655
rect 3450 3565 3460 3645
rect 3540 3565 3550 3645
rect 3450 3555 3550 3565
rect 3650 3645 3750 3655
rect 3650 3565 3660 3645
rect 3740 3565 3750 3645
rect 3650 3555 3750 3565
rect 3850 3645 3950 3655
rect 3850 3565 3860 3645
rect 3940 3565 3950 3645
rect 3850 3555 3950 3565
rect 4050 3645 4150 3655
rect 4050 3565 4060 3645
rect 4140 3565 4150 3645
rect 4050 3555 4150 3565
rect 4250 3645 4350 3655
rect 4250 3565 4260 3645
rect 4340 3565 4350 3645
rect 4250 3555 4350 3565
rect 4450 3645 4550 3655
rect 4450 3565 4460 3645
rect 4540 3565 4550 3645
rect 4450 3555 4550 3565
rect 4650 3645 4750 3655
rect 4650 3565 4660 3645
rect 4740 3565 4750 3645
rect 4650 3555 4750 3565
rect 4850 3645 4950 3655
rect 4850 3565 4860 3645
rect 4940 3565 4950 3645
rect 4850 3555 4950 3565
rect 5050 3645 5150 3655
rect 5050 3565 5060 3645
rect 5140 3565 5150 3645
rect 5050 3555 5150 3565
rect 5250 3645 5350 3655
rect 5250 3565 5260 3645
rect 5340 3565 5350 3645
rect 5250 3555 5350 3565
rect 5450 3645 5550 3655
rect 5450 3565 5460 3645
rect 5540 3565 5550 3645
rect 5450 3555 5550 3565
rect 5650 3645 5750 3655
rect 5650 3565 5660 3645
rect 5740 3565 5750 3645
rect 5650 3555 5750 3565
rect 5850 3645 5950 3655
rect 5850 3565 5860 3645
rect 5940 3565 5950 3645
rect 5850 3555 5950 3565
rect 6050 3645 6150 3655
rect 6050 3565 6060 3645
rect 6140 3565 6150 3645
rect 6050 3555 6150 3565
rect 6250 3645 6350 3655
rect 6250 3565 6260 3645
rect 6340 3565 6350 3645
rect 6250 3555 6350 3565
rect 6450 3645 6550 3655
rect 6450 3565 6460 3645
rect 6540 3565 6550 3645
rect 6450 3555 6550 3565
rect -150 3460 -50 3470
rect -150 3380 -140 3460
rect -60 3380 -50 3460
rect -150 3370 -50 3380
rect 50 3460 150 3470
rect 50 3380 60 3460
rect 140 3380 150 3460
rect 50 3370 150 3380
rect 250 3460 350 3470
rect 250 3380 260 3460
rect 340 3380 350 3460
rect 250 3370 350 3380
rect 450 3460 550 3470
rect 450 3380 460 3460
rect 540 3380 550 3460
rect 450 3370 550 3380
rect 650 3460 750 3470
rect 650 3380 660 3460
rect 740 3380 750 3460
rect 650 3370 750 3380
rect 850 3460 950 3470
rect 850 3380 860 3460
rect 940 3380 950 3460
rect 850 3370 950 3380
rect 1050 3460 1150 3470
rect 1050 3380 1060 3460
rect 1140 3380 1150 3460
rect 1050 3370 1150 3380
rect 1250 3460 1350 3470
rect 1250 3380 1260 3460
rect 1340 3380 1350 3460
rect 1250 3370 1350 3380
rect 1450 3460 1550 3470
rect 1450 3380 1460 3460
rect 1540 3380 1550 3460
rect 1450 3370 1550 3380
rect 1650 3460 1750 3470
rect 1650 3380 1660 3460
rect 1740 3380 1750 3460
rect 1650 3370 1750 3380
rect 1850 3460 1950 3470
rect 1850 3380 1860 3460
rect 1940 3380 1950 3460
rect 1850 3370 1950 3380
rect 2050 3460 2150 3470
rect 2050 3380 2060 3460
rect 2140 3380 2150 3460
rect 2050 3370 2150 3380
rect 2250 3460 2350 3470
rect 2250 3380 2260 3460
rect 2340 3380 2350 3460
rect 2250 3370 2350 3380
rect 2450 3460 2550 3470
rect 2450 3380 2460 3460
rect 2540 3380 2550 3460
rect 2450 3370 2550 3380
rect 2650 3460 2750 3470
rect 2650 3380 2660 3460
rect 2740 3380 2750 3460
rect 2650 3370 2750 3380
rect 2850 3460 2950 3470
rect 2850 3380 2860 3460
rect 2940 3380 2950 3460
rect 2850 3370 2950 3380
rect 3050 3460 3150 3470
rect 3050 3380 3060 3460
rect 3140 3380 3150 3460
rect 3050 3370 3150 3380
rect 3250 3460 3350 3470
rect 3250 3380 3260 3460
rect 3340 3380 3350 3460
rect 3250 3370 3350 3380
rect 3450 3460 3550 3470
rect 3450 3380 3460 3460
rect 3540 3380 3550 3460
rect 3450 3370 3550 3380
rect 3650 3460 3750 3470
rect 3650 3380 3660 3460
rect 3740 3380 3750 3460
rect 3650 3370 3750 3380
rect 3850 3460 3950 3470
rect 3850 3380 3860 3460
rect 3940 3380 3950 3460
rect 3850 3370 3950 3380
rect 4050 3460 4150 3470
rect 4050 3380 4060 3460
rect 4140 3380 4150 3460
rect 4050 3370 4150 3380
rect 4250 3460 4350 3470
rect 4250 3380 4260 3460
rect 4340 3380 4350 3460
rect 4250 3370 4350 3380
rect 4450 3460 4550 3470
rect 4450 3380 4460 3460
rect 4540 3380 4550 3460
rect 4450 3370 4550 3380
rect 4650 3460 4750 3470
rect 4650 3380 4660 3460
rect 4740 3380 4750 3460
rect 4650 3370 4750 3380
rect 4850 3460 4950 3470
rect 4850 3380 4860 3460
rect 4940 3380 4950 3460
rect 4850 3370 4950 3380
rect 5050 3460 5150 3470
rect 5050 3380 5060 3460
rect 5140 3380 5150 3460
rect 5050 3370 5150 3380
rect 5250 3460 5350 3470
rect 5250 3380 5260 3460
rect 5340 3380 5350 3460
rect 5250 3370 5350 3380
rect 5450 3460 5550 3470
rect 5450 3380 5460 3460
rect 5540 3380 5550 3460
rect 5450 3370 5550 3380
rect 5650 3460 5750 3470
rect 5650 3380 5660 3460
rect 5740 3380 5750 3460
rect 5650 3370 5750 3380
rect 5850 3460 5950 3470
rect 5850 3380 5860 3460
rect 5940 3380 5950 3460
rect 5850 3370 5950 3380
rect 6050 3460 6150 3470
rect 6050 3380 6060 3460
rect 6140 3380 6150 3460
rect 6050 3370 6150 3380
rect 6250 3460 6350 3470
rect 6250 3380 6260 3460
rect 6340 3380 6350 3460
rect 6250 3370 6350 3380
rect 6450 3460 6550 3470
rect 6450 3380 6460 3460
rect 6540 3380 6550 3460
rect 6450 3370 6550 3380
rect -150 3275 -50 3285
rect -150 3195 -140 3275
rect -60 3195 -50 3275
rect -150 3185 -50 3195
rect 50 3275 150 3285
rect 50 3195 60 3275
rect 140 3195 150 3275
rect 50 3185 150 3195
rect 250 3275 350 3285
rect 250 3195 260 3275
rect 340 3195 350 3275
rect 250 3185 350 3195
rect 450 3275 550 3285
rect 450 3195 460 3275
rect 540 3195 550 3275
rect 450 3185 550 3195
rect 650 3275 750 3285
rect 650 3195 660 3275
rect 740 3195 750 3275
rect 650 3185 750 3195
rect 850 3275 950 3285
rect 850 3195 860 3275
rect 940 3195 950 3275
rect 850 3185 950 3195
rect 1050 3275 1150 3285
rect 1050 3195 1060 3275
rect 1140 3195 1150 3275
rect 1050 3185 1150 3195
rect 1250 3275 1350 3285
rect 1250 3195 1260 3275
rect 1340 3195 1350 3275
rect 1250 3185 1350 3195
rect 1450 3275 1550 3285
rect 1450 3195 1460 3275
rect 1540 3195 1550 3275
rect 1450 3185 1550 3195
rect 1650 3275 1750 3285
rect 1650 3195 1660 3275
rect 1740 3195 1750 3275
rect 1650 3185 1750 3195
rect 1850 3275 1950 3285
rect 1850 3195 1860 3275
rect 1940 3195 1950 3275
rect 1850 3185 1950 3195
rect 2050 3275 2150 3285
rect 2050 3195 2060 3275
rect 2140 3195 2150 3275
rect 2050 3185 2150 3195
rect 2250 3275 2350 3285
rect 2250 3195 2260 3275
rect 2340 3195 2350 3275
rect 2250 3185 2350 3195
rect 2450 3275 2550 3285
rect 2450 3195 2460 3275
rect 2540 3195 2550 3275
rect 2450 3185 2550 3195
rect 2650 3275 2750 3285
rect 2650 3195 2660 3275
rect 2740 3195 2750 3275
rect 2650 3185 2750 3195
rect 2850 3275 2950 3285
rect 2850 3195 2860 3275
rect 2940 3195 2950 3275
rect 2850 3185 2950 3195
rect 3050 3275 3150 3285
rect 3050 3195 3060 3275
rect 3140 3195 3150 3275
rect 3050 3185 3150 3195
rect 3250 3275 3350 3285
rect 3250 3195 3260 3275
rect 3340 3195 3350 3275
rect 3250 3185 3350 3195
rect 3450 3275 3550 3285
rect 3450 3195 3460 3275
rect 3540 3195 3550 3275
rect 3450 3185 3550 3195
rect 3650 3275 3750 3285
rect 3650 3195 3660 3275
rect 3740 3195 3750 3275
rect 3650 3185 3750 3195
rect 3850 3275 3950 3285
rect 3850 3195 3860 3275
rect 3940 3195 3950 3275
rect 3850 3185 3950 3195
rect 4050 3275 4150 3285
rect 4050 3195 4060 3275
rect 4140 3195 4150 3275
rect 4050 3185 4150 3195
rect 4250 3275 4350 3285
rect 4250 3195 4260 3275
rect 4340 3195 4350 3275
rect 4250 3185 4350 3195
rect 4450 3275 4550 3285
rect 4450 3195 4460 3275
rect 4540 3195 4550 3275
rect 4450 3185 4550 3195
rect 4650 3275 4750 3285
rect 4650 3195 4660 3275
rect 4740 3195 4750 3275
rect 4650 3185 4750 3195
rect 4850 3275 4950 3285
rect 4850 3195 4860 3275
rect 4940 3195 4950 3275
rect 4850 3185 4950 3195
rect 5050 3275 5150 3285
rect 5050 3195 5060 3275
rect 5140 3195 5150 3275
rect 5050 3185 5150 3195
rect 5250 3275 5350 3285
rect 5250 3195 5260 3275
rect 5340 3195 5350 3275
rect 5250 3185 5350 3195
rect 5450 3275 5550 3285
rect 5450 3195 5460 3275
rect 5540 3195 5550 3275
rect 5450 3185 5550 3195
rect 5650 3275 5750 3285
rect 5650 3195 5660 3275
rect 5740 3195 5750 3275
rect 5650 3185 5750 3195
rect 5850 3275 5950 3285
rect 5850 3195 5860 3275
rect 5940 3195 5950 3275
rect 5850 3185 5950 3195
rect 6050 3275 6150 3285
rect 6050 3195 6060 3275
rect 6140 3195 6150 3275
rect 6050 3185 6150 3195
rect 6250 3275 6350 3285
rect 6250 3195 6260 3275
rect 6340 3195 6350 3275
rect 6250 3185 6350 3195
rect 6450 3275 6550 3285
rect 6450 3195 6460 3275
rect 6540 3195 6550 3275
rect 6450 3185 6550 3195
rect -150 3090 -50 3100
rect -150 3010 -140 3090
rect -60 3010 -50 3090
rect -150 3000 -50 3010
rect 50 3090 150 3100
rect 50 3010 60 3090
rect 140 3010 150 3090
rect 50 3000 150 3010
rect 250 3090 350 3100
rect 250 3010 260 3090
rect 340 3010 350 3090
rect 250 3000 350 3010
rect 450 3090 550 3100
rect 450 3010 460 3090
rect 540 3010 550 3090
rect 450 3000 550 3010
rect 650 3090 750 3100
rect 650 3010 660 3090
rect 740 3010 750 3090
rect 650 3000 750 3010
rect 850 3090 950 3100
rect 850 3010 860 3090
rect 940 3010 950 3090
rect 850 3000 950 3010
rect 1050 3090 1150 3100
rect 1050 3010 1060 3090
rect 1140 3010 1150 3090
rect 1050 3000 1150 3010
rect 1250 3090 1350 3100
rect 1250 3010 1260 3090
rect 1340 3010 1350 3090
rect 1250 3000 1350 3010
rect 1450 3090 1550 3100
rect 1450 3010 1460 3090
rect 1540 3010 1550 3090
rect 1450 3000 1550 3010
rect 1650 3090 1750 3100
rect 1650 3010 1660 3090
rect 1740 3010 1750 3090
rect 1650 3000 1750 3010
rect 1850 3090 1950 3100
rect 1850 3010 1860 3090
rect 1940 3010 1950 3090
rect 1850 3000 1950 3010
rect 2050 3090 2150 3100
rect 2050 3010 2060 3090
rect 2140 3010 2150 3090
rect 2050 3000 2150 3010
rect 2250 3090 2350 3100
rect 2250 3010 2260 3090
rect 2340 3010 2350 3090
rect 2250 3000 2350 3010
rect 2450 3090 2550 3100
rect 2450 3010 2460 3090
rect 2540 3010 2550 3090
rect 2450 3000 2550 3010
rect 2650 3090 2750 3100
rect 2650 3010 2660 3090
rect 2740 3010 2750 3090
rect 2650 3000 2750 3010
rect 2850 3090 2950 3100
rect 2850 3010 2860 3090
rect 2940 3010 2950 3090
rect 2850 3000 2950 3010
rect 3050 3090 3150 3100
rect 3050 3010 3060 3090
rect 3140 3010 3150 3090
rect 3050 3000 3150 3010
rect 3250 3090 3350 3100
rect 3250 3010 3260 3090
rect 3340 3010 3350 3090
rect 3250 3000 3350 3010
rect 3450 3090 3550 3100
rect 3450 3010 3460 3090
rect 3540 3010 3550 3090
rect 3450 3000 3550 3010
rect 3650 3090 3750 3100
rect 3650 3010 3660 3090
rect 3740 3010 3750 3090
rect 3650 3000 3750 3010
rect 3850 3090 3950 3100
rect 3850 3010 3860 3090
rect 3940 3010 3950 3090
rect 3850 3000 3950 3010
rect 4050 3090 4150 3100
rect 4050 3010 4060 3090
rect 4140 3010 4150 3090
rect 4050 3000 4150 3010
rect 4250 3090 4350 3100
rect 4250 3010 4260 3090
rect 4340 3010 4350 3090
rect 4250 3000 4350 3010
rect 4450 3090 4550 3100
rect 4450 3010 4460 3090
rect 4540 3010 4550 3090
rect 4450 3000 4550 3010
rect 4650 3090 4750 3100
rect 4650 3010 4660 3090
rect 4740 3010 4750 3090
rect 4650 3000 4750 3010
rect 4850 3090 4950 3100
rect 4850 3010 4860 3090
rect 4940 3010 4950 3090
rect 4850 3000 4950 3010
rect 5050 3090 5150 3100
rect 5050 3010 5060 3090
rect 5140 3010 5150 3090
rect 5050 3000 5150 3010
rect 5250 3090 5350 3100
rect 5250 3010 5260 3090
rect 5340 3010 5350 3090
rect 5250 3000 5350 3010
rect 5450 3090 5550 3100
rect 5450 3010 5460 3090
rect 5540 3010 5550 3090
rect 5450 3000 5550 3010
rect 5650 3090 5750 3100
rect 5650 3010 5660 3090
rect 5740 3010 5750 3090
rect 5650 3000 5750 3010
rect 5850 3090 5950 3100
rect 5850 3010 5860 3090
rect 5940 3010 5950 3090
rect 5850 3000 5950 3010
rect 6050 3090 6150 3100
rect 6050 3010 6060 3090
rect 6140 3010 6150 3090
rect 6050 3000 6150 3010
rect 6250 3090 6350 3100
rect 6250 3010 6260 3090
rect 6340 3010 6350 3090
rect 6250 3000 6350 3010
rect 6450 3090 6550 3100
rect 6450 3010 6460 3090
rect 6540 3010 6550 3090
rect 6450 3000 6550 3010
rect -150 2905 -50 2915
rect -150 2825 -140 2905
rect -60 2825 -50 2905
rect -150 2815 -50 2825
rect 50 2905 150 2915
rect 50 2825 60 2905
rect 140 2825 150 2905
rect 50 2815 150 2825
rect 250 2905 350 2915
rect 250 2825 260 2905
rect 340 2825 350 2905
rect 250 2815 350 2825
rect 450 2905 550 2915
rect 450 2825 460 2905
rect 540 2825 550 2905
rect 450 2815 550 2825
rect 650 2905 750 2915
rect 650 2825 660 2905
rect 740 2825 750 2905
rect 650 2815 750 2825
rect 850 2905 950 2915
rect 850 2825 860 2905
rect 940 2825 950 2905
rect 850 2815 950 2825
rect 1050 2905 1150 2915
rect 1050 2825 1060 2905
rect 1140 2825 1150 2905
rect 1050 2815 1150 2825
rect 1250 2905 1350 2915
rect 1250 2825 1260 2905
rect 1340 2825 1350 2905
rect 1250 2815 1350 2825
rect 1450 2905 1550 2915
rect 1450 2825 1460 2905
rect 1540 2825 1550 2905
rect 1450 2815 1550 2825
rect 1650 2905 1750 2915
rect 1650 2825 1660 2905
rect 1740 2825 1750 2905
rect 1650 2815 1750 2825
rect 1850 2905 1950 2915
rect 1850 2825 1860 2905
rect 1940 2825 1950 2905
rect 1850 2815 1950 2825
rect 2050 2905 2150 2915
rect 2050 2825 2060 2905
rect 2140 2825 2150 2905
rect 2050 2815 2150 2825
rect 2250 2905 2350 2915
rect 2250 2825 2260 2905
rect 2340 2825 2350 2905
rect 2250 2815 2350 2825
rect 2450 2905 2550 2915
rect 2450 2825 2460 2905
rect 2540 2825 2550 2905
rect 2450 2815 2550 2825
rect 2650 2905 2750 2915
rect 2650 2825 2660 2905
rect 2740 2825 2750 2905
rect 2650 2815 2750 2825
rect 2850 2905 2950 2915
rect 2850 2825 2860 2905
rect 2940 2825 2950 2905
rect 2850 2815 2950 2825
rect 3050 2905 3150 2915
rect 3050 2825 3060 2905
rect 3140 2825 3150 2905
rect 3050 2815 3150 2825
rect 3250 2905 3350 2915
rect 3250 2825 3260 2905
rect 3340 2825 3350 2905
rect 3250 2815 3350 2825
rect 3450 2905 3550 2915
rect 3450 2825 3460 2905
rect 3540 2825 3550 2905
rect 3450 2815 3550 2825
rect 3650 2905 3750 2915
rect 3650 2825 3660 2905
rect 3740 2825 3750 2905
rect 3650 2815 3750 2825
rect 3850 2905 3950 2915
rect 3850 2825 3860 2905
rect 3940 2825 3950 2905
rect 3850 2815 3950 2825
rect 4050 2905 4150 2915
rect 4050 2825 4060 2905
rect 4140 2825 4150 2905
rect 4050 2815 4150 2825
rect 4250 2905 4350 2915
rect 4250 2825 4260 2905
rect 4340 2825 4350 2905
rect 4250 2815 4350 2825
rect 4450 2905 4550 2915
rect 4450 2825 4460 2905
rect 4540 2825 4550 2905
rect 4450 2815 4550 2825
rect 4650 2905 4750 2915
rect 4650 2825 4660 2905
rect 4740 2825 4750 2905
rect 4650 2815 4750 2825
rect 4850 2905 4950 2915
rect 4850 2825 4860 2905
rect 4940 2825 4950 2905
rect 4850 2815 4950 2825
rect 5050 2905 5150 2915
rect 5050 2825 5060 2905
rect 5140 2825 5150 2905
rect 5050 2815 5150 2825
rect 5250 2905 5350 2915
rect 5250 2825 5260 2905
rect 5340 2825 5350 2905
rect 5250 2815 5350 2825
rect 5450 2905 5550 2915
rect 5450 2825 5460 2905
rect 5540 2825 5550 2905
rect 5450 2815 5550 2825
rect 5650 2905 5750 2915
rect 5650 2825 5660 2905
rect 5740 2825 5750 2905
rect 5650 2815 5750 2825
rect 5850 2905 5950 2915
rect 5850 2825 5860 2905
rect 5940 2825 5950 2905
rect 5850 2815 5950 2825
rect 6050 2905 6150 2915
rect 6050 2825 6060 2905
rect 6140 2825 6150 2905
rect 6050 2815 6150 2825
rect 6250 2905 6350 2915
rect 6250 2825 6260 2905
rect 6340 2825 6350 2905
rect 6250 2815 6350 2825
rect 6450 2905 6550 2915
rect 6450 2825 6460 2905
rect 6540 2825 6550 2905
rect 6450 2815 6550 2825
rect -150 2720 -50 2730
rect -150 2640 -140 2720
rect -60 2640 -50 2720
rect -150 2630 -50 2640
rect 50 2720 150 2730
rect 50 2640 60 2720
rect 140 2640 150 2720
rect 50 2630 150 2640
rect 250 2720 350 2730
rect 250 2640 260 2720
rect 340 2640 350 2720
rect 250 2630 350 2640
rect 450 2720 550 2730
rect 450 2640 460 2720
rect 540 2640 550 2720
rect 450 2630 550 2640
rect 650 2720 750 2730
rect 650 2640 660 2720
rect 740 2640 750 2720
rect 650 2630 750 2640
rect 850 2720 950 2730
rect 850 2640 860 2720
rect 940 2640 950 2720
rect 850 2630 950 2640
rect 1050 2720 1150 2730
rect 1050 2640 1060 2720
rect 1140 2640 1150 2720
rect 1050 2630 1150 2640
rect 1250 2720 1350 2730
rect 1250 2640 1260 2720
rect 1340 2640 1350 2720
rect 1250 2630 1350 2640
rect 1450 2720 1550 2730
rect 1450 2640 1460 2720
rect 1540 2640 1550 2720
rect 1450 2630 1550 2640
rect 1650 2720 1750 2730
rect 1650 2640 1660 2720
rect 1740 2640 1750 2720
rect 1650 2630 1750 2640
rect 1850 2720 1950 2730
rect 1850 2640 1860 2720
rect 1940 2640 1950 2720
rect 1850 2630 1950 2640
rect 2050 2720 2150 2730
rect 2050 2640 2060 2720
rect 2140 2640 2150 2720
rect 2050 2630 2150 2640
rect 2250 2720 2350 2730
rect 2250 2640 2260 2720
rect 2340 2640 2350 2720
rect 2250 2630 2350 2640
rect 2450 2720 2550 2730
rect 2450 2640 2460 2720
rect 2540 2640 2550 2720
rect 2450 2630 2550 2640
rect 2650 2720 2750 2730
rect 2650 2640 2660 2720
rect 2740 2640 2750 2720
rect 2650 2630 2750 2640
rect 2850 2720 2950 2730
rect 2850 2640 2860 2720
rect 2940 2640 2950 2720
rect 2850 2630 2950 2640
rect 3050 2720 3150 2730
rect 3050 2640 3060 2720
rect 3140 2640 3150 2720
rect 3050 2630 3150 2640
rect 3250 2720 3350 2730
rect 3250 2640 3260 2720
rect 3340 2640 3350 2720
rect 3250 2630 3350 2640
rect 3450 2720 3550 2730
rect 3450 2640 3460 2720
rect 3540 2640 3550 2720
rect 3450 2630 3550 2640
rect 3650 2720 3750 2730
rect 3650 2640 3660 2720
rect 3740 2640 3750 2720
rect 3650 2630 3750 2640
rect 3850 2720 3950 2730
rect 3850 2640 3860 2720
rect 3940 2640 3950 2720
rect 3850 2630 3950 2640
rect 4050 2720 4150 2730
rect 4050 2640 4060 2720
rect 4140 2640 4150 2720
rect 4050 2630 4150 2640
rect 4250 2720 4350 2730
rect 4250 2640 4260 2720
rect 4340 2640 4350 2720
rect 4250 2630 4350 2640
rect 4450 2720 4550 2730
rect 4450 2640 4460 2720
rect 4540 2640 4550 2720
rect 4450 2630 4550 2640
rect 4650 2720 4750 2730
rect 4650 2640 4660 2720
rect 4740 2640 4750 2720
rect 4650 2630 4750 2640
rect 4850 2720 4950 2730
rect 4850 2640 4860 2720
rect 4940 2640 4950 2720
rect 4850 2630 4950 2640
rect 5050 2720 5150 2730
rect 5050 2640 5060 2720
rect 5140 2640 5150 2720
rect 5050 2630 5150 2640
rect 5250 2720 5350 2730
rect 5250 2640 5260 2720
rect 5340 2640 5350 2720
rect 5250 2630 5350 2640
rect 5450 2720 5550 2730
rect 5450 2640 5460 2720
rect 5540 2640 5550 2720
rect 5450 2630 5550 2640
rect 5650 2720 5750 2730
rect 5650 2640 5660 2720
rect 5740 2640 5750 2720
rect 5650 2630 5750 2640
rect 5850 2720 5950 2730
rect 5850 2640 5860 2720
rect 5940 2640 5950 2720
rect 5850 2630 5950 2640
rect 6050 2720 6150 2730
rect 6050 2640 6060 2720
rect 6140 2640 6150 2720
rect 6050 2630 6150 2640
rect 6250 2720 6350 2730
rect 6250 2640 6260 2720
rect 6340 2640 6350 2720
rect 6250 2630 6350 2640
rect 6450 2720 6550 2730
rect 6450 2640 6460 2720
rect 6540 2640 6550 2720
rect 6450 2630 6550 2640
rect -150 2535 -50 2545
rect -150 2455 -140 2535
rect -60 2455 -50 2535
rect -150 2445 -50 2455
rect 50 2535 150 2545
rect 50 2455 60 2535
rect 140 2455 150 2535
rect 50 2445 150 2455
rect 250 2535 350 2545
rect 250 2455 260 2535
rect 340 2455 350 2535
rect 250 2445 350 2455
rect 450 2535 550 2545
rect 450 2455 460 2535
rect 540 2455 550 2535
rect 450 2445 550 2455
rect 650 2535 750 2545
rect 650 2455 660 2535
rect 740 2455 750 2535
rect 650 2445 750 2455
rect 850 2535 950 2545
rect 850 2455 860 2535
rect 940 2455 950 2535
rect 850 2445 950 2455
rect 1050 2535 1150 2545
rect 1050 2455 1060 2535
rect 1140 2455 1150 2535
rect 1050 2445 1150 2455
rect 1250 2535 1350 2545
rect 1250 2455 1260 2535
rect 1340 2455 1350 2535
rect 1250 2445 1350 2455
rect 1450 2535 1550 2545
rect 1450 2455 1460 2535
rect 1540 2455 1550 2535
rect 1450 2445 1550 2455
rect 1650 2535 1750 2545
rect 1650 2455 1660 2535
rect 1740 2455 1750 2535
rect 1650 2445 1750 2455
rect 1850 2535 1950 2545
rect 1850 2455 1860 2535
rect 1940 2455 1950 2535
rect 1850 2445 1950 2455
rect 2050 2535 2150 2545
rect 2050 2455 2060 2535
rect 2140 2455 2150 2535
rect 2050 2445 2150 2455
rect 2250 2535 2350 2545
rect 2250 2455 2260 2535
rect 2340 2455 2350 2535
rect 2250 2445 2350 2455
rect 2450 2535 2550 2545
rect 2450 2455 2460 2535
rect 2540 2455 2550 2535
rect 2450 2445 2550 2455
rect 2650 2535 2750 2545
rect 2650 2455 2660 2535
rect 2740 2455 2750 2535
rect 2650 2445 2750 2455
rect 2850 2535 2950 2545
rect 2850 2455 2860 2535
rect 2940 2455 2950 2535
rect 2850 2445 2950 2455
rect 3050 2535 3150 2545
rect 3050 2455 3060 2535
rect 3140 2455 3150 2535
rect 3050 2445 3150 2455
rect 3250 2535 3350 2545
rect 3250 2455 3260 2535
rect 3340 2455 3350 2535
rect 3250 2445 3350 2455
rect 3450 2535 3550 2545
rect 3450 2455 3460 2535
rect 3540 2455 3550 2535
rect 3450 2445 3550 2455
rect 3650 2535 3750 2545
rect 3650 2455 3660 2535
rect 3740 2455 3750 2535
rect 3650 2445 3750 2455
rect 3850 2535 3950 2545
rect 3850 2455 3860 2535
rect 3940 2455 3950 2535
rect 3850 2445 3950 2455
rect 4050 2535 4150 2545
rect 4050 2455 4060 2535
rect 4140 2455 4150 2535
rect 4050 2445 4150 2455
rect 4250 2535 4350 2545
rect 4250 2455 4260 2535
rect 4340 2455 4350 2535
rect 4250 2445 4350 2455
rect 4450 2535 4550 2545
rect 4450 2455 4460 2535
rect 4540 2455 4550 2535
rect 4450 2445 4550 2455
rect 4650 2535 4750 2545
rect 4650 2455 4660 2535
rect 4740 2455 4750 2535
rect 4650 2445 4750 2455
rect 4850 2535 4950 2545
rect 4850 2455 4860 2535
rect 4940 2455 4950 2535
rect 4850 2445 4950 2455
rect 5050 2535 5150 2545
rect 5050 2455 5060 2535
rect 5140 2455 5150 2535
rect 5050 2445 5150 2455
rect 5250 2535 5350 2545
rect 5250 2455 5260 2535
rect 5340 2455 5350 2535
rect 5250 2445 5350 2455
rect 5450 2535 5550 2545
rect 5450 2455 5460 2535
rect 5540 2455 5550 2535
rect 5450 2445 5550 2455
rect 5650 2535 5750 2545
rect 5650 2455 5660 2535
rect 5740 2455 5750 2535
rect 5650 2445 5750 2455
rect 5850 2535 5950 2545
rect 5850 2455 5860 2535
rect 5940 2455 5950 2535
rect 5850 2445 5950 2455
rect 6050 2535 6150 2545
rect 6050 2455 6060 2535
rect 6140 2455 6150 2535
rect 6050 2445 6150 2455
rect 6250 2535 6350 2545
rect 6250 2455 6260 2535
rect 6340 2455 6350 2535
rect 6250 2445 6350 2455
rect 6450 2535 6550 2545
rect 6450 2455 6460 2535
rect 6540 2455 6550 2535
rect 6450 2445 6550 2455
rect -150 2350 -50 2360
rect -150 2270 -140 2350
rect -60 2270 -50 2350
rect -150 2260 -50 2270
rect 50 2350 150 2360
rect 50 2270 60 2350
rect 140 2270 150 2350
rect 50 2260 150 2270
rect 250 2350 350 2360
rect 250 2270 260 2350
rect 340 2270 350 2350
rect 250 2260 350 2270
rect 450 2350 550 2360
rect 450 2270 460 2350
rect 540 2270 550 2350
rect 450 2260 550 2270
rect 650 2350 750 2360
rect 650 2270 660 2350
rect 740 2270 750 2350
rect 650 2260 750 2270
rect 850 2350 950 2360
rect 850 2270 860 2350
rect 940 2270 950 2350
rect 850 2260 950 2270
rect 1050 2350 1150 2360
rect 1050 2270 1060 2350
rect 1140 2270 1150 2350
rect 1050 2260 1150 2270
rect 1250 2350 1350 2360
rect 1250 2270 1260 2350
rect 1340 2270 1350 2350
rect 1250 2260 1350 2270
rect 1450 2350 1550 2360
rect 1450 2270 1460 2350
rect 1540 2270 1550 2350
rect 1450 2260 1550 2270
rect 1650 2350 1750 2360
rect 1650 2270 1660 2350
rect 1740 2270 1750 2350
rect 1650 2260 1750 2270
rect 1850 2350 1950 2360
rect 1850 2270 1860 2350
rect 1940 2270 1950 2350
rect 1850 2260 1950 2270
rect 2050 2350 2150 2360
rect 2050 2270 2060 2350
rect 2140 2270 2150 2350
rect 2050 2260 2150 2270
rect 2250 2350 2350 2360
rect 2250 2270 2260 2350
rect 2340 2270 2350 2350
rect 2250 2260 2350 2270
rect 2450 2350 2550 2360
rect 2450 2270 2460 2350
rect 2540 2270 2550 2350
rect 2450 2260 2550 2270
rect 2650 2350 2750 2360
rect 2650 2270 2660 2350
rect 2740 2270 2750 2350
rect 2650 2260 2750 2270
rect 2850 2350 2950 2360
rect 2850 2270 2860 2350
rect 2940 2270 2950 2350
rect 2850 2260 2950 2270
rect 3050 2350 3150 2360
rect 3050 2270 3060 2350
rect 3140 2270 3150 2350
rect 3050 2260 3150 2270
rect 3250 2350 3350 2360
rect 3250 2270 3260 2350
rect 3340 2270 3350 2350
rect 3250 2260 3350 2270
rect 3450 2350 3550 2360
rect 3450 2270 3460 2350
rect 3540 2270 3550 2350
rect 3450 2260 3550 2270
rect 3650 2350 3750 2360
rect 3650 2270 3660 2350
rect 3740 2270 3750 2350
rect 3650 2260 3750 2270
rect 3850 2350 3950 2360
rect 3850 2270 3860 2350
rect 3940 2270 3950 2350
rect 3850 2260 3950 2270
rect 4050 2350 4150 2360
rect 4050 2270 4060 2350
rect 4140 2270 4150 2350
rect 4050 2260 4150 2270
rect 4250 2350 4350 2360
rect 4250 2270 4260 2350
rect 4340 2270 4350 2350
rect 4250 2260 4350 2270
rect 4450 2350 4550 2360
rect 4450 2270 4460 2350
rect 4540 2270 4550 2350
rect 4450 2260 4550 2270
rect 4650 2350 4750 2360
rect 4650 2270 4660 2350
rect 4740 2270 4750 2350
rect 4650 2260 4750 2270
rect 4850 2350 4950 2360
rect 4850 2270 4860 2350
rect 4940 2270 4950 2350
rect 4850 2260 4950 2270
rect 5050 2350 5150 2360
rect 5050 2270 5060 2350
rect 5140 2270 5150 2350
rect 5050 2260 5150 2270
rect 5250 2350 5350 2360
rect 5250 2270 5260 2350
rect 5340 2270 5350 2350
rect 5250 2260 5350 2270
rect 5450 2350 5550 2360
rect 5450 2270 5460 2350
rect 5540 2270 5550 2350
rect 5450 2260 5550 2270
rect 5650 2350 5750 2360
rect 5650 2270 5660 2350
rect 5740 2270 5750 2350
rect 5650 2260 5750 2270
rect 5850 2350 5950 2360
rect 5850 2270 5860 2350
rect 5940 2270 5950 2350
rect 5850 2260 5950 2270
rect 6050 2350 6150 2360
rect 6050 2270 6060 2350
rect 6140 2270 6150 2350
rect 6050 2260 6150 2270
rect 6250 2350 6350 2360
rect 6250 2270 6260 2350
rect 6340 2270 6350 2350
rect 6250 2260 6350 2270
rect 6450 2350 6550 2360
rect 6450 2270 6460 2350
rect 6540 2270 6550 2350
rect 6450 2260 6550 2270
rect -150 2165 -50 2175
rect -150 2085 -140 2165
rect -60 2085 -50 2165
rect -150 2075 -50 2085
rect 50 2165 150 2175
rect 50 2085 60 2165
rect 140 2085 150 2165
rect 50 2075 150 2085
rect 250 2165 350 2175
rect 250 2085 260 2165
rect 340 2085 350 2165
rect 250 2075 350 2085
rect 450 2165 550 2175
rect 450 2085 460 2165
rect 540 2085 550 2165
rect 450 2075 550 2085
rect 650 2165 750 2175
rect 650 2085 660 2165
rect 740 2085 750 2165
rect 650 2075 750 2085
rect 850 2165 950 2175
rect 850 2085 860 2165
rect 940 2085 950 2165
rect 850 2075 950 2085
rect 1050 2165 1150 2175
rect 1050 2085 1060 2165
rect 1140 2085 1150 2165
rect 1050 2075 1150 2085
rect 1250 2165 1350 2175
rect 1250 2085 1260 2165
rect 1340 2085 1350 2165
rect 1250 2075 1350 2085
rect 1450 2165 1550 2175
rect 1450 2085 1460 2165
rect 1540 2085 1550 2165
rect 1450 2075 1550 2085
rect 1650 2165 1750 2175
rect 1650 2085 1660 2165
rect 1740 2085 1750 2165
rect 1650 2075 1750 2085
rect 1850 2165 1950 2175
rect 1850 2085 1860 2165
rect 1940 2085 1950 2165
rect 1850 2075 1950 2085
rect 2050 2165 2150 2175
rect 2050 2085 2060 2165
rect 2140 2085 2150 2165
rect 2050 2075 2150 2085
rect 2250 2165 2350 2175
rect 2250 2085 2260 2165
rect 2340 2085 2350 2165
rect 2250 2075 2350 2085
rect 2450 2165 2550 2175
rect 2450 2085 2460 2165
rect 2540 2085 2550 2165
rect 2450 2075 2550 2085
rect 2650 2165 2750 2175
rect 2650 2085 2660 2165
rect 2740 2085 2750 2165
rect 2650 2075 2750 2085
rect 2850 2165 2950 2175
rect 2850 2085 2860 2165
rect 2940 2085 2950 2165
rect 2850 2075 2950 2085
rect 3050 2165 3150 2175
rect 3050 2085 3060 2165
rect 3140 2085 3150 2165
rect 3050 2075 3150 2085
rect 3250 2165 3350 2175
rect 3250 2085 3260 2165
rect 3340 2085 3350 2165
rect 3250 2075 3350 2085
rect 3450 2165 3550 2175
rect 3450 2085 3460 2165
rect 3540 2085 3550 2165
rect 3450 2075 3550 2085
rect 3650 2165 3750 2175
rect 3650 2085 3660 2165
rect 3740 2085 3750 2165
rect 3650 2075 3750 2085
rect 3850 2165 3950 2175
rect 3850 2085 3860 2165
rect 3940 2085 3950 2165
rect 3850 2075 3950 2085
rect 4050 2165 4150 2175
rect 4050 2085 4060 2165
rect 4140 2085 4150 2165
rect 4050 2075 4150 2085
rect 4250 2165 4350 2175
rect 4250 2085 4260 2165
rect 4340 2085 4350 2165
rect 4250 2075 4350 2085
rect 4450 2165 4550 2175
rect 4450 2085 4460 2165
rect 4540 2085 4550 2165
rect 4450 2075 4550 2085
rect 4650 2165 4750 2175
rect 4650 2085 4660 2165
rect 4740 2085 4750 2165
rect 4650 2075 4750 2085
rect 4850 2165 4950 2175
rect 4850 2085 4860 2165
rect 4940 2085 4950 2165
rect 4850 2075 4950 2085
rect 5050 2165 5150 2175
rect 5050 2085 5060 2165
rect 5140 2085 5150 2165
rect 5050 2075 5150 2085
rect 5250 2165 5350 2175
rect 5250 2085 5260 2165
rect 5340 2085 5350 2165
rect 5250 2075 5350 2085
rect 5450 2165 5550 2175
rect 5450 2085 5460 2165
rect 5540 2085 5550 2165
rect 5450 2075 5550 2085
rect 5650 2165 5750 2175
rect 5650 2085 5660 2165
rect 5740 2085 5750 2165
rect 5650 2075 5750 2085
rect 5850 2165 5950 2175
rect 5850 2085 5860 2165
rect 5940 2085 5950 2165
rect 5850 2075 5950 2085
rect 6050 2165 6150 2175
rect 6050 2085 6060 2165
rect 6140 2085 6150 2165
rect 6050 2075 6150 2085
rect 6250 2165 6350 2175
rect 6250 2085 6260 2165
rect 6340 2085 6350 2165
rect 6250 2075 6350 2085
rect 6450 2165 6550 2175
rect 6450 2085 6460 2165
rect 6540 2085 6550 2165
rect 6450 2075 6550 2085
rect -150 1980 -50 1990
rect -150 1900 -140 1980
rect -60 1900 -50 1980
rect -150 1890 -50 1900
rect 50 1980 150 1990
rect 50 1900 60 1980
rect 140 1900 150 1980
rect 50 1890 150 1900
rect 250 1980 350 1990
rect 250 1900 260 1980
rect 340 1900 350 1980
rect 250 1890 350 1900
rect 450 1980 550 1990
rect 450 1900 460 1980
rect 540 1900 550 1980
rect 450 1890 550 1900
rect 650 1980 750 1990
rect 650 1900 660 1980
rect 740 1900 750 1980
rect 650 1890 750 1900
rect 850 1980 950 1990
rect 850 1900 860 1980
rect 940 1900 950 1980
rect 850 1890 950 1900
rect 1050 1980 1150 1990
rect 1050 1900 1060 1980
rect 1140 1900 1150 1980
rect 1050 1890 1150 1900
rect 1250 1980 1350 1990
rect 1250 1900 1260 1980
rect 1340 1900 1350 1980
rect 1250 1890 1350 1900
rect 1450 1980 1550 1990
rect 1450 1900 1460 1980
rect 1540 1900 1550 1980
rect 1450 1890 1550 1900
rect 1650 1980 1750 1990
rect 1650 1900 1660 1980
rect 1740 1900 1750 1980
rect 1650 1890 1750 1900
rect 1850 1980 1950 1990
rect 1850 1900 1860 1980
rect 1940 1900 1950 1980
rect 1850 1890 1950 1900
rect 2050 1980 2150 1990
rect 2050 1900 2060 1980
rect 2140 1900 2150 1980
rect 2050 1890 2150 1900
rect 2250 1980 2350 1990
rect 2250 1900 2260 1980
rect 2340 1900 2350 1980
rect 2250 1890 2350 1900
rect 2450 1980 2550 1990
rect 2450 1900 2460 1980
rect 2540 1900 2550 1980
rect 2450 1890 2550 1900
rect 2650 1980 2750 1990
rect 2650 1900 2660 1980
rect 2740 1900 2750 1980
rect 2650 1890 2750 1900
rect 2850 1980 2950 1990
rect 2850 1900 2860 1980
rect 2940 1900 2950 1980
rect 2850 1890 2950 1900
rect 3050 1980 3150 1990
rect 3050 1900 3060 1980
rect 3140 1900 3150 1980
rect 3050 1890 3150 1900
rect 3250 1980 3350 1990
rect 3250 1900 3260 1980
rect 3340 1900 3350 1980
rect 3250 1890 3350 1900
rect 3450 1980 3550 1990
rect 3450 1900 3460 1980
rect 3540 1900 3550 1980
rect 3450 1890 3550 1900
rect 3650 1980 3750 1990
rect 3650 1900 3660 1980
rect 3740 1900 3750 1980
rect 3650 1890 3750 1900
rect 3850 1980 3950 1990
rect 3850 1900 3860 1980
rect 3940 1900 3950 1980
rect 3850 1890 3950 1900
rect 4050 1980 4150 1990
rect 4050 1900 4060 1980
rect 4140 1900 4150 1980
rect 4050 1890 4150 1900
rect 4250 1980 4350 1990
rect 4250 1900 4260 1980
rect 4340 1900 4350 1980
rect 4250 1890 4350 1900
rect 4450 1980 4550 1990
rect 4450 1900 4460 1980
rect 4540 1900 4550 1980
rect 4450 1890 4550 1900
rect 4650 1980 4750 1990
rect 4650 1900 4660 1980
rect 4740 1900 4750 1980
rect 4650 1890 4750 1900
rect 4850 1980 4950 1990
rect 4850 1900 4860 1980
rect 4940 1900 4950 1980
rect 4850 1890 4950 1900
rect 5050 1980 5150 1990
rect 5050 1900 5060 1980
rect 5140 1900 5150 1980
rect 5050 1890 5150 1900
rect 5250 1980 5350 1990
rect 5250 1900 5260 1980
rect 5340 1900 5350 1980
rect 5250 1890 5350 1900
rect 5450 1980 5550 1990
rect 5450 1900 5460 1980
rect 5540 1900 5550 1980
rect 5450 1890 5550 1900
rect 5650 1980 5750 1990
rect 5650 1900 5660 1980
rect 5740 1900 5750 1980
rect 5650 1890 5750 1900
rect 5850 1980 5950 1990
rect 5850 1900 5860 1980
rect 5940 1900 5950 1980
rect 5850 1890 5950 1900
rect 6050 1980 6150 1990
rect 6050 1900 6060 1980
rect 6140 1900 6150 1980
rect 6050 1890 6150 1900
rect 6250 1980 6350 1990
rect 6250 1900 6260 1980
rect 6340 1900 6350 1980
rect 6250 1890 6350 1900
rect 6450 1980 6550 1990
rect 6450 1900 6460 1980
rect 6540 1900 6550 1980
rect 6450 1890 6550 1900
rect -150 1795 -50 1805
rect -150 1715 -140 1795
rect -60 1715 -50 1795
rect -150 1705 -50 1715
rect 50 1795 150 1805
rect 50 1715 60 1795
rect 140 1715 150 1795
rect 50 1705 150 1715
rect 250 1795 350 1805
rect 250 1715 260 1795
rect 340 1715 350 1795
rect 250 1705 350 1715
rect 450 1795 550 1805
rect 450 1715 460 1795
rect 540 1715 550 1795
rect 450 1705 550 1715
rect 650 1795 750 1805
rect 650 1715 660 1795
rect 740 1715 750 1795
rect 650 1705 750 1715
rect 850 1795 950 1805
rect 850 1715 860 1795
rect 940 1715 950 1795
rect 850 1705 950 1715
rect 1050 1795 1150 1805
rect 1050 1715 1060 1795
rect 1140 1715 1150 1795
rect 1050 1705 1150 1715
rect 1250 1795 1350 1805
rect 1250 1715 1260 1795
rect 1340 1715 1350 1795
rect 1250 1705 1350 1715
rect 1450 1795 1550 1805
rect 1450 1715 1460 1795
rect 1540 1715 1550 1795
rect 1450 1705 1550 1715
rect 1650 1795 1750 1805
rect 1650 1715 1660 1795
rect 1740 1715 1750 1795
rect 1650 1705 1750 1715
rect 1850 1795 1950 1805
rect 1850 1715 1860 1795
rect 1940 1715 1950 1795
rect 1850 1705 1950 1715
rect 2050 1795 2150 1805
rect 2050 1715 2060 1795
rect 2140 1715 2150 1795
rect 2050 1705 2150 1715
rect 2250 1795 2350 1805
rect 2250 1715 2260 1795
rect 2340 1715 2350 1795
rect 2250 1705 2350 1715
rect 2450 1795 2550 1805
rect 2450 1715 2460 1795
rect 2540 1715 2550 1795
rect 2450 1705 2550 1715
rect 2650 1795 2750 1805
rect 2650 1715 2660 1795
rect 2740 1715 2750 1795
rect 2650 1705 2750 1715
rect 2850 1795 2950 1805
rect 2850 1715 2860 1795
rect 2940 1715 2950 1795
rect 2850 1705 2950 1715
rect 3050 1795 3150 1805
rect 3050 1715 3060 1795
rect 3140 1715 3150 1795
rect 3050 1705 3150 1715
rect 3250 1795 3350 1805
rect 3250 1715 3260 1795
rect 3340 1715 3350 1795
rect 3250 1705 3350 1715
rect 3450 1795 3550 1805
rect 3450 1715 3460 1795
rect 3540 1715 3550 1795
rect 3450 1705 3550 1715
rect 3650 1795 3750 1805
rect 3650 1715 3660 1795
rect 3740 1715 3750 1795
rect 3650 1705 3750 1715
rect 3850 1795 3950 1805
rect 3850 1715 3860 1795
rect 3940 1715 3950 1795
rect 3850 1705 3950 1715
rect 4050 1795 4150 1805
rect 4050 1715 4060 1795
rect 4140 1715 4150 1795
rect 4050 1705 4150 1715
rect 4250 1795 4350 1805
rect 4250 1715 4260 1795
rect 4340 1715 4350 1795
rect 4250 1705 4350 1715
rect 4450 1795 4550 1805
rect 4450 1715 4460 1795
rect 4540 1715 4550 1795
rect 4450 1705 4550 1715
rect 4650 1795 4750 1805
rect 4650 1715 4660 1795
rect 4740 1715 4750 1795
rect 4650 1705 4750 1715
rect 4850 1795 4950 1805
rect 4850 1715 4860 1795
rect 4940 1715 4950 1795
rect 4850 1705 4950 1715
rect 5050 1795 5150 1805
rect 5050 1715 5060 1795
rect 5140 1715 5150 1795
rect 5050 1705 5150 1715
rect 5250 1795 5350 1805
rect 5250 1715 5260 1795
rect 5340 1715 5350 1795
rect 5250 1705 5350 1715
rect 5450 1795 5550 1805
rect 5450 1715 5460 1795
rect 5540 1715 5550 1795
rect 5450 1705 5550 1715
rect 5650 1795 5750 1805
rect 5650 1715 5660 1795
rect 5740 1715 5750 1795
rect 5650 1705 5750 1715
rect 5850 1795 5950 1805
rect 5850 1715 5860 1795
rect 5940 1715 5950 1795
rect 5850 1705 5950 1715
rect 6050 1795 6150 1805
rect 6050 1715 6060 1795
rect 6140 1715 6150 1795
rect 6050 1705 6150 1715
rect 6250 1795 6350 1805
rect 6250 1715 6260 1795
rect 6340 1715 6350 1795
rect 6250 1705 6350 1715
rect 6450 1795 6550 1805
rect 6450 1715 6460 1795
rect 6540 1715 6550 1795
rect 6450 1705 6550 1715
rect -150 1610 -50 1620
rect -150 1530 -140 1610
rect -60 1530 -50 1610
rect -150 1520 -50 1530
rect 50 1610 150 1620
rect 50 1530 60 1610
rect 140 1530 150 1610
rect 50 1520 150 1530
rect 250 1610 350 1620
rect 250 1530 260 1610
rect 340 1530 350 1610
rect 250 1520 350 1530
rect 450 1610 550 1620
rect 450 1530 460 1610
rect 540 1530 550 1610
rect 450 1520 550 1530
rect 650 1610 750 1620
rect 650 1530 660 1610
rect 740 1530 750 1610
rect 650 1520 750 1530
rect 850 1610 950 1620
rect 850 1530 860 1610
rect 940 1530 950 1610
rect 850 1520 950 1530
rect 1050 1610 1150 1620
rect 1050 1530 1060 1610
rect 1140 1530 1150 1610
rect 1050 1520 1150 1530
rect 1250 1610 1350 1620
rect 1250 1530 1260 1610
rect 1340 1530 1350 1610
rect 1250 1520 1350 1530
rect 1450 1610 1550 1620
rect 1450 1530 1460 1610
rect 1540 1530 1550 1610
rect 1450 1520 1550 1530
rect 1650 1610 1750 1620
rect 1650 1530 1660 1610
rect 1740 1530 1750 1610
rect 1650 1520 1750 1530
rect 1850 1610 1950 1620
rect 1850 1530 1860 1610
rect 1940 1530 1950 1610
rect 1850 1520 1950 1530
rect 2050 1610 2150 1620
rect 2050 1530 2060 1610
rect 2140 1530 2150 1610
rect 2050 1520 2150 1530
rect 2250 1610 2350 1620
rect 2250 1530 2260 1610
rect 2340 1530 2350 1610
rect 2250 1520 2350 1530
rect 2450 1610 2550 1620
rect 2450 1530 2460 1610
rect 2540 1530 2550 1610
rect 2450 1520 2550 1530
rect 2650 1610 2750 1620
rect 2650 1530 2660 1610
rect 2740 1530 2750 1610
rect 2650 1520 2750 1530
rect 2850 1610 2950 1620
rect 2850 1530 2860 1610
rect 2940 1530 2950 1610
rect 2850 1520 2950 1530
rect 3050 1610 3150 1620
rect 3050 1530 3060 1610
rect 3140 1530 3150 1610
rect 3050 1520 3150 1530
rect 3250 1610 3350 1620
rect 3250 1530 3260 1610
rect 3340 1530 3350 1610
rect 3250 1520 3350 1530
rect 3450 1610 3550 1620
rect 3450 1530 3460 1610
rect 3540 1530 3550 1610
rect 3450 1520 3550 1530
rect 3650 1610 3750 1620
rect 3650 1530 3660 1610
rect 3740 1530 3750 1610
rect 3650 1520 3750 1530
rect 3850 1610 3950 1620
rect 3850 1530 3860 1610
rect 3940 1530 3950 1610
rect 3850 1520 3950 1530
rect 4050 1610 4150 1620
rect 4050 1530 4060 1610
rect 4140 1530 4150 1610
rect 4050 1520 4150 1530
rect 4250 1610 4350 1620
rect 4250 1530 4260 1610
rect 4340 1530 4350 1610
rect 4250 1520 4350 1530
rect 4450 1610 4550 1620
rect 4450 1530 4460 1610
rect 4540 1530 4550 1610
rect 4450 1520 4550 1530
rect 4650 1610 4750 1620
rect 4650 1530 4660 1610
rect 4740 1530 4750 1610
rect 4650 1520 4750 1530
rect 4850 1610 4950 1620
rect 4850 1530 4860 1610
rect 4940 1530 4950 1610
rect 4850 1520 4950 1530
rect 5050 1610 5150 1620
rect 5050 1530 5060 1610
rect 5140 1530 5150 1610
rect 5050 1520 5150 1530
rect 5250 1610 5350 1620
rect 5250 1530 5260 1610
rect 5340 1530 5350 1610
rect 5250 1520 5350 1530
rect 5450 1610 5550 1620
rect 5450 1530 5460 1610
rect 5540 1530 5550 1610
rect 5450 1520 5550 1530
rect 5650 1610 5750 1620
rect 5650 1530 5660 1610
rect 5740 1530 5750 1610
rect 5650 1520 5750 1530
rect 5850 1610 5950 1620
rect 5850 1530 5860 1610
rect 5940 1530 5950 1610
rect 5850 1520 5950 1530
rect 6050 1610 6150 1620
rect 6050 1530 6060 1610
rect 6140 1530 6150 1610
rect 6050 1520 6150 1530
rect 6250 1610 6350 1620
rect 6250 1530 6260 1610
rect 6340 1530 6350 1610
rect 6250 1520 6350 1530
rect 6450 1610 6550 1620
rect 6450 1530 6460 1610
rect 6540 1530 6550 1610
rect 6450 1520 6550 1530
rect -150 1425 -50 1435
rect -150 1345 -140 1425
rect -60 1345 -50 1425
rect -150 1335 -50 1345
rect 50 1425 150 1435
rect 50 1345 60 1425
rect 140 1345 150 1425
rect 50 1335 150 1345
rect 250 1425 350 1435
rect 250 1345 260 1425
rect 340 1345 350 1425
rect 250 1335 350 1345
rect 450 1425 550 1435
rect 450 1345 460 1425
rect 540 1345 550 1425
rect 450 1335 550 1345
rect 650 1425 750 1435
rect 650 1345 660 1425
rect 740 1345 750 1425
rect 650 1335 750 1345
rect 850 1425 950 1435
rect 850 1345 860 1425
rect 940 1345 950 1425
rect 850 1335 950 1345
rect 1050 1425 1150 1435
rect 1050 1345 1060 1425
rect 1140 1345 1150 1425
rect 1050 1335 1150 1345
rect 1250 1425 1350 1435
rect 1250 1345 1260 1425
rect 1340 1345 1350 1425
rect 1250 1335 1350 1345
rect 1450 1425 1550 1435
rect 1450 1345 1460 1425
rect 1540 1345 1550 1425
rect 1450 1335 1550 1345
rect 1650 1425 1750 1435
rect 1650 1345 1660 1425
rect 1740 1345 1750 1425
rect 1650 1335 1750 1345
rect 1850 1425 1950 1435
rect 1850 1345 1860 1425
rect 1940 1345 1950 1425
rect 1850 1335 1950 1345
rect 2050 1425 2150 1435
rect 2050 1345 2060 1425
rect 2140 1345 2150 1425
rect 2050 1335 2150 1345
rect 2250 1425 2350 1435
rect 2250 1345 2260 1425
rect 2340 1345 2350 1425
rect 2250 1335 2350 1345
rect 2450 1425 2550 1435
rect 2450 1345 2460 1425
rect 2540 1345 2550 1425
rect 2450 1335 2550 1345
rect 2650 1425 2750 1435
rect 2650 1345 2660 1425
rect 2740 1345 2750 1425
rect 2650 1335 2750 1345
rect 2850 1425 2950 1435
rect 2850 1345 2860 1425
rect 2940 1345 2950 1425
rect 2850 1335 2950 1345
rect 3050 1425 3150 1435
rect 3050 1345 3060 1425
rect 3140 1345 3150 1425
rect 3050 1335 3150 1345
rect 3250 1425 3350 1435
rect 3250 1345 3260 1425
rect 3340 1345 3350 1425
rect 3250 1335 3350 1345
rect 3450 1425 3550 1435
rect 3450 1345 3460 1425
rect 3540 1345 3550 1425
rect 3450 1335 3550 1345
rect 3650 1425 3750 1435
rect 3650 1345 3660 1425
rect 3740 1345 3750 1425
rect 3650 1335 3750 1345
rect 3850 1425 3950 1435
rect 3850 1345 3860 1425
rect 3940 1345 3950 1425
rect 3850 1335 3950 1345
rect 4050 1425 4150 1435
rect 4050 1345 4060 1425
rect 4140 1345 4150 1425
rect 4050 1335 4150 1345
rect 4250 1425 4350 1435
rect 4250 1345 4260 1425
rect 4340 1345 4350 1425
rect 4250 1335 4350 1345
rect 4450 1425 4550 1435
rect 4450 1345 4460 1425
rect 4540 1345 4550 1425
rect 4450 1335 4550 1345
rect 4650 1425 4750 1435
rect 4650 1345 4660 1425
rect 4740 1345 4750 1425
rect 4650 1335 4750 1345
rect 4850 1425 4950 1435
rect 4850 1345 4860 1425
rect 4940 1345 4950 1425
rect 4850 1335 4950 1345
rect 5050 1425 5150 1435
rect 5050 1345 5060 1425
rect 5140 1345 5150 1425
rect 5050 1335 5150 1345
rect 5250 1425 5350 1435
rect 5250 1345 5260 1425
rect 5340 1345 5350 1425
rect 5250 1335 5350 1345
rect 5450 1425 5550 1435
rect 5450 1345 5460 1425
rect 5540 1345 5550 1425
rect 5450 1335 5550 1345
rect 5650 1425 5750 1435
rect 5650 1345 5660 1425
rect 5740 1345 5750 1425
rect 5650 1335 5750 1345
rect 5850 1425 5950 1435
rect 5850 1345 5860 1425
rect 5940 1345 5950 1425
rect 5850 1335 5950 1345
rect 6050 1425 6150 1435
rect 6050 1345 6060 1425
rect 6140 1345 6150 1425
rect 6050 1335 6150 1345
rect 6250 1425 6350 1435
rect 6250 1345 6260 1425
rect 6340 1345 6350 1425
rect 6250 1335 6350 1345
rect 6450 1425 6550 1435
rect 6450 1345 6460 1425
rect 6540 1345 6550 1425
rect 6450 1335 6550 1345
rect -150 1240 -50 1250
rect -150 1160 -140 1240
rect -60 1160 -50 1240
rect -150 1150 -50 1160
rect 50 1240 150 1250
rect 50 1160 60 1240
rect 140 1160 150 1240
rect 50 1150 150 1160
rect 250 1240 350 1250
rect 250 1160 260 1240
rect 340 1160 350 1240
rect 250 1150 350 1160
rect 450 1240 550 1250
rect 450 1160 460 1240
rect 540 1160 550 1240
rect 450 1150 550 1160
rect 650 1240 750 1250
rect 650 1160 660 1240
rect 740 1160 750 1240
rect 650 1150 750 1160
rect 850 1240 950 1250
rect 850 1160 860 1240
rect 940 1160 950 1240
rect 850 1150 950 1160
rect 1050 1240 1150 1250
rect 1050 1160 1060 1240
rect 1140 1160 1150 1240
rect 1050 1150 1150 1160
rect 1250 1240 1350 1250
rect 1250 1160 1260 1240
rect 1340 1160 1350 1240
rect 1250 1150 1350 1160
rect 1450 1240 1550 1250
rect 1450 1160 1460 1240
rect 1540 1160 1550 1240
rect 1450 1150 1550 1160
rect 1650 1240 1750 1250
rect 1650 1160 1660 1240
rect 1740 1160 1750 1240
rect 1650 1150 1750 1160
rect 1850 1240 1950 1250
rect 1850 1160 1860 1240
rect 1940 1160 1950 1240
rect 1850 1150 1950 1160
rect 2050 1240 2150 1250
rect 2050 1160 2060 1240
rect 2140 1160 2150 1240
rect 2050 1150 2150 1160
rect 2250 1240 2350 1250
rect 2250 1160 2260 1240
rect 2340 1160 2350 1240
rect 2250 1150 2350 1160
rect 2450 1240 2550 1250
rect 2450 1160 2460 1240
rect 2540 1160 2550 1240
rect 2450 1150 2550 1160
rect 2650 1240 2750 1250
rect 2650 1160 2660 1240
rect 2740 1160 2750 1240
rect 2650 1150 2750 1160
rect 2850 1240 2950 1250
rect 2850 1160 2860 1240
rect 2940 1160 2950 1240
rect 2850 1150 2950 1160
rect 3050 1240 3150 1250
rect 3050 1160 3060 1240
rect 3140 1160 3150 1240
rect 3050 1150 3150 1160
rect 3250 1240 3350 1250
rect 3250 1160 3260 1240
rect 3340 1160 3350 1240
rect 3250 1150 3350 1160
rect 3450 1240 3550 1250
rect 3450 1160 3460 1240
rect 3540 1160 3550 1240
rect 3450 1150 3550 1160
rect 3650 1240 3750 1250
rect 3650 1160 3660 1240
rect 3740 1160 3750 1240
rect 3650 1150 3750 1160
rect 3850 1240 3950 1250
rect 3850 1160 3860 1240
rect 3940 1160 3950 1240
rect 3850 1150 3950 1160
rect 4050 1240 4150 1250
rect 4050 1160 4060 1240
rect 4140 1160 4150 1240
rect 4050 1150 4150 1160
rect 4250 1240 4350 1250
rect 4250 1160 4260 1240
rect 4340 1160 4350 1240
rect 4250 1150 4350 1160
rect 4450 1240 4550 1250
rect 4450 1160 4460 1240
rect 4540 1160 4550 1240
rect 4450 1150 4550 1160
rect 4650 1240 4750 1250
rect 4650 1160 4660 1240
rect 4740 1160 4750 1240
rect 4650 1150 4750 1160
rect 4850 1240 4950 1250
rect 4850 1160 4860 1240
rect 4940 1160 4950 1240
rect 4850 1150 4950 1160
rect 5050 1240 5150 1250
rect 5050 1160 5060 1240
rect 5140 1160 5150 1240
rect 5050 1150 5150 1160
rect 5250 1240 5350 1250
rect 5250 1160 5260 1240
rect 5340 1160 5350 1240
rect 5250 1150 5350 1160
rect 5450 1240 5550 1250
rect 5450 1160 5460 1240
rect 5540 1160 5550 1240
rect 5450 1150 5550 1160
rect 5650 1240 5750 1250
rect 5650 1160 5660 1240
rect 5740 1160 5750 1240
rect 5650 1150 5750 1160
rect 5850 1240 5950 1250
rect 5850 1160 5860 1240
rect 5940 1160 5950 1240
rect 5850 1150 5950 1160
rect 6050 1240 6150 1250
rect 6050 1160 6060 1240
rect 6140 1160 6150 1240
rect 6050 1150 6150 1160
rect 6250 1240 6350 1250
rect 6250 1160 6260 1240
rect 6340 1160 6350 1240
rect 6250 1150 6350 1160
rect 6450 1240 6550 1250
rect 6450 1160 6460 1240
rect 6540 1160 6550 1240
rect 6450 1150 6550 1160
rect -150 1055 -50 1065
rect -150 975 -140 1055
rect -60 975 -50 1055
rect -150 965 -50 975
rect 50 1055 150 1065
rect 50 975 60 1055
rect 140 975 150 1055
rect 50 965 150 975
rect 250 1055 350 1065
rect 250 975 260 1055
rect 340 975 350 1055
rect 250 965 350 975
rect 450 1055 550 1065
rect 450 975 460 1055
rect 540 975 550 1055
rect 450 965 550 975
rect 650 1055 750 1065
rect 650 975 660 1055
rect 740 975 750 1055
rect 650 965 750 975
rect 850 1055 950 1065
rect 850 975 860 1055
rect 940 975 950 1055
rect 850 965 950 975
rect 1050 1055 1150 1065
rect 1050 975 1060 1055
rect 1140 975 1150 1055
rect 1050 965 1150 975
rect 1250 1055 1350 1065
rect 1250 975 1260 1055
rect 1340 975 1350 1055
rect 1250 965 1350 975
rect 1450 1055 1550 1065
rect 1450 975 1460 1055
rect 1540 975 1550 1055
rect 1450 965 1550 975
rect 1650 1055 1750 1065
rect 1650 975 1660 1055
rect 1740 975 1750 1055
rect 1650 965 1750 975
rect 1850 1055 1950 1065
rect 1850 975 1860 1055
rect 1940 975 1950 1055
rect 1850 965 1950 975
rect 2050 1055 2150 1065
rect 2050 975 2060 1055
rect 2140 975 2150 1055
rect 2050 965 2150 975
rect 2250 1055 2350 1065
rect 2250 975 2260 1055
rect 2340 975 2350 1055
rect 2250 965 2350 975
rect 2450 1055 2550 1065
rect 2450 975 2460 1055
rect 2540 975 2550 1055
rect 2450 965 2550 975
rect 2650 1055 2750 1065
rect 2650 975 2660 1055
rect 2740 975 2750 1055
rect 2650 965 2750 975
rect 2850 1055 2950 1065
rect 2850 975 2860 1055
rect 2940 975 2950 1055
rect 2850 965 2950 975
rect 3050 1055 3150 1065
rect 3050 975 3060 1055
rect 3140 975 3150 1055
rect 3050 965 3150 975
rect 3250 1055 3350 1065
rect 3250 975 3260 1055
rect 3340 975 3350 1055
rect 3250 965 3350 975
rect 3450 1055 3550 1065
rect 3450 975 3460 1055
rect 3540 975 3550 1055
rect 3450 965 3550 975
rect 3650 1055 3750 1065
rect 3650 975 3660 1055
rect 3740 975 3750 1055
rect 3650 965 3750 975
rect 3850 1055 3950 1065
rect 3850 975 3860 1055
rect 3940 975 3950 1055
rect 3850 965 3950 975
rect 4050 1055 4150 1065
rect 4050 975 4060 1055
rect 4140 975 4150 1055
rect 4050 965 4150 975
rect 4250 1055 4350 1065
rect 4250 975 4260 1055
rect 4340 975 4350 1055
rect 4250 965 4350 975
rect 4450 1055 4550 1065
rect 4450 975 4460 1055
rect 4540 975 4550 1055
rect 4450 965 4550 975
rect 4650 1055 4750 1065
rect 4650 975 4660 1055
rect 4740 975 4750 1055
rect 4650 965 4750 975
rect 4850 1055 4950 1065
rect 4850 975 4860 1055
rect 4940 975 4950 1055
rect 4850 965 4950 975
rect 5050 1055 5150 1065
rect 5050 975 5060 1055
rect 5140 975 5150 1055
rect 5050 965 5150 975
rect 5250 1055 5350 1065
rect 5250 975 5260 1055
rect 5340 975 5350 1055
rect 5250 965 5350 975
rect 5450 1055 5550 1065
rect 5450 975 5460 1055
rect 5540 975 5550 1055
rect 5450 965 5550 975
rect 5650 1055 5750 1065
rect 5650 975 5660 1055
rect 5740 975 5750 1055
rect 5650 965 5750 975
rect 5850 1055 5950 1065
rect 5850 975 5860 1055
rect 5940 975 5950 1055
rect 5850 965 5950 975
rect 6050 1055 6150 1065
rect 6050 975 6060 1055
rect 6140 975 6150 1055
rect 6050 965 6150 975
rect 6250 1055 6350 1065
rect 6250 975 6260 1055
rect 6340 975 6350 1055
rect 6250 965 6350 975
rect 6450 1055 6550 1065
rect 6450 975 6460 1055
rect 6540 975 6550 1055
rect 6450 965 6550 975
rect -150 870 -50 880
rect -150 790 -140 870
rect -60 790 -50 870
rect -150 780 -50 790
rect 50 870 150 880
rect 50 790 60 870
rect 140 790 150 870
rect 50 780 150 790
rect 250 870 350 880
rect 250 790 260 870
rect 340 790 350 870
rect 250 780 350 790
rect 450 870 550 880
rect 450 790 460 870
rect 540 790 550 870
rect 450 780 550 790
rect 650 870 750 880
rect 650 790 660 870
rect 740 790 750 870
rect 650 780 750 790
rect 850 870 950 880
rect 850 790 860 870
rect 940 790 950 870
rect 850 780 950 790
rect 1050 870 1150 880
rect 1050 790 1060 870
rect 1140 790 1150 870
rect 1050 780 1150 790
rect 1250 870 1350 880
rect 1250 790 1260 870
rect 1340 790 1350 870
rect 1250 780 1350 790
rect 1450 870 1550 880
rect 1450 790 1460 870
rect 1540 790 1550 870
rect 1450 780 1550 790
rect 1650 870 1750 880
rect 1650 790 1660 870
rect 1740 790 1750 870
rect 1650 780 1750 790
rect 1850 870 1950 880
rect 1850 790 1860 870
rect 1940 790 1950 870
rect 1850 780 1950 790
rect 2050 870 2150 880
rect 2050 790 2060 870
rect 2140 790 2150 870
rect 2050 780 2150 790
rect 2250 870 2350 880
rect 2250 790 2260 870
rect 2340 790 2350 870
rect 2250 780 2350 790
rect 2450 870 2550 880
rect 2450 790 2460 870
rect 2540 790 2550 870
rect 2450 780 2550 790
rect 2650 870 2750 880
rect 2650 790 2660 870
rect 2740 790 2750 870
rect 2650 780 2750 790
rect 2850 870 2950 880
rect 2850 790 2860 870
rect 2940 790 2950 870
rect 2850 780 2950 790
rect 3050 870 3150 880
rect 3050 790 3060 870
rect 3140 790 3150 870
rect 3050 780 3150 790
rect 3250 870 3350 880
rect 3250 790 3260 870
rect 3340 790 3350 870
rect 3250 780 3350 790
rect 3450 870 3550 880
rect 3450 790 3460 870
rect 3540 790 3550 870
rect 3450 780 3550 790
rect 3650 870 3750 880
rect 3650 790 3660 870
rect 3740 790 3750 870
rect 3650 780 3750 790
rect 3850 870 3950 880
rect 3850 790 3860 870
rect 3940 790 3950 870
rect 3850 780 3950 790
rect 4050 870 4150 880
rect 4050 790 4060 870
rect 4140 790 4150 870
rect 4050 780 4150 790
rect 4250 870 4350 880
rect 4250 790 4260 870
rect 4340 790 4350 870
rect 4250 780 4350 790
rect 4450 870 4550 880
rect 4450 790 4460 870
rect 4540 790 4550 870
rect 4450 780 4550 790
rect 4650 870 4750 880
rect 4650 790 4660 870
rect 4740 790 4750 870
rect 4650 780 4750 790
rect 4850 870 4950 880
rect 4850 790 4860 870
rect 4940 790 4950 870
rect 4850 780 4950 790
rect 5050 870 5150 880
rect 5050 790 5060 870
rect 5140 790 5150 870
rect 5050 780 5150 790
rect 5250 870 5350 880
rect 5250 790 5260 870
rect 5340 790 5350 870
rect 5250 780 5350 790
rect 5450 870 5550 880
rect 5450 790 5460 870
rect 5540 790 5550 870
rect 5450 780 5550 790
rect 5650 870 5750 880
rect 5650 790 5660 870
rect 5740 790 5750 870
rect 5650 780 5750 790
rect 5850 870 5950 880
rect 5850 790 5860 870
rect 5940 790 5950 870
rect 5850 780 5950 790
rect 6050 870 6150 880
rect 6050 790 6060 870
rect 6140 790 6150 870
rect 6050 780 6150 790
rect 6250 870 6350 880
rect 6250 790 6260 870
rect 6340 790 6350 870
rect 6250 780 6350 790
rect 6450 870 6550 880
rect 6450 790 6460 870
rect 6540 790 6550 870
rect 6450 780 6550 790
rect -150 685 -50 695
rect -150 605 -140 685
rect -60 605 -50 685
rect -150 595 -50 605
rect 50 685 150 695
rect 50 605 60 685
rect 140 605 150 685
rect 50 595 150 605
rect 250 685 350 695
rect 250 605 260 685
rect 340 605 350 685
rect 250 595 350 605
rect 450 685 550 695
rect 450 605 460 685
rect 540 605 550 685
rect 450 595 550 605
rect 650 685 750 695
rect 650 605 660 685
rect 740 605 750 685
rect 650 595 750 605
rect 850 685 950 695
rect 850 605 860 685
rect 940 605 950 685
rect 850 595 950 605
rect 1050 685 1150 695
rect 1050 605 1060 685
rect 1140 605 1150 685
rect 1050 595 1150 605
rect 1250 685 1350 695
rect 1250 605 1260 685
rect 1340 605 1350 685
rect 1250 595 1350 605
rect 1450 685 1550 695
rect 1450 605 1460 685
rect 1540 605 1550 685
rect 1450 595 1550 605
rect 1650 685 1750 695
rect 1650 605 1660 685
rect 1740 605 1750 685
rect 1650 595 1750 605
rect 1850 685 1950 695
rect 1850 605 1860 685
rect 1940 605 1950 685
rect 1850 595 1950 605
rect 2050 685 2150 695
rect 2050 605 2060 685
rect 2140 605 2150 685
rect 2050 595 2150 605
rect 2250 685 2350 695
rect 2250 605 2260 685
rect 2340 605 2350 685
rect 2250 595 2350 605
rect 2450 685 2550 695
rect 2450 605 2460 685
rect 2540 605 2550 685
rect 2450 595 2550 605
rect 2650 685 2750 695
rect 2650 605 2660 685
rect 2740 605 2750 685
rect 2650 595 2750 605
rect 2850 685 2950 695
rect 2850 605 2860 685
rect 2940 605 2950 685
rect 2850 595 2950 605
rect 3050 685 3150 695
rect 3050 605 3060 685
rect 3140 605 3150 685
rect 3050 595 3150 605
rect 3250 685 3350 695
rect 3250 605 3260 685
rect 3340 605 3350 685
rect 3250 595 3350 605
rect 3450 685 3550 695
rect 3450 605 3460 685
rect 3540 605 3550 685
rect 3450 595 3550 605
rect 3650 685 3750 695
rect 3650 605 3660 685
rect 3740 605 3750 685
rect 3650 595 3750 605
rect 3850 685 3950 695
rect 3850 605 3860 685
rect 3940 605 3950 685
rect 3850 595 3950 605
rect 4050 685 4150 695
rect 4050 605 4060 685
rect 4140 605 4150 685
rect 4050 595 4150 605
rect 4250 685 4350 695
rect 4250 605 4260 685
rect 4340 605 4350 685
rect 4250 595 4350 605
rect 4450 685 4550 695
rect 4450 605 4460 685
rect 4540 605 4550 685
rect 4450 595 4550 605
rect 4650 685 4750 695
rect 4650 605 4660 685
rect 4740 605 4750 685
rect 4650 595 4750 605
rect 4850 685 4950 695
rect 4850 605 4860 685
rect 4940 605 4950 685
rect 4850 595 4950 605
rect 5050 685 5150 695
rect 5050 605 5060 685
rect 5140 605 5150 685
rect 5050 595 5150 605
rect 5250 685 5350 695
rect 5250 605 5260 685
rect 5340 605 5350 685
rect 5250 595 5350 605
rect 5450 685 5550 695
rect 5450 605 5460 685
rect 5540 605 5550 685
rect 5450 595 5550 605
rect 5650 685 5750 695
rect 5650 605 5660 685
rect 5740 605 5750 685
rect 5650 595 5750 605
rect 5850 685 5950 695
rect 5850 605 5860 685
rect 5940 605 5950 685
rect 5850 595 5950 605
rect 6050 685 6150 695
rect 6050 605 6060 685
rect 6140 605 6150 685
rect 6050 595 6150 605
rect 6250 685 6350 695
rect 6250 605 6260 685
rect 6340 605 6350 685
rect 6250 595 6350 605
rect 6450 685 6550 695
rect 6450 605 6460 685
rect 6540 605 6550 685
rect 6450 595 6550 605
rect -150 500 -50 510
rect -150 420 -140 500
rect -60 420 -50 500
rect -150 410 -50 420
rect 50 500 150 510
rect 50 420 60 500
rect 140 420 150 500
rect 50 410 150 420
rect 250 500 350 510
rect 250 420 260 500
rect 340 420 350 500
rect 250 410 350 420
rect 450 500 550 510
rect 450 420 460 500
rect 540 420 550 500
rect 450 410 550 420
rect 650 500 750 510
rect 650 420 660 500
rect 740 420 750 500
rect 650 410 750 420
rect 850 500 950 510
rect 850 420 860 500
rect 940 420 950 500
rect 850 410 950 420
rect 1050 500 1150 510
rect 1050 420 1060 500
rect 1140 420 1150 500
rect 1050 410 1150 420
rect 1250 500 1350 510
rect 1250 420 1260 500
rect 1340 420 1350 500
rect 1250 410 1350 420
rect 1450 500 1550 510
rect 1450 420 1460 500
rect 1540 420 1550 500
rect 1450 410 1550 420
rect 1650 500 1750 510
rect 1650 420 1660 500
rect 1740 420 1750 500
rect 1650 410 1750 420
rect 1850 500 1950 510
rect 1850 420 1860 500
rect 1940 420 1950 500
rect 1850 410 1950 420
rect 2050 500 2150 510
rect 2050 420 2060 500
rect 2140 420 2150 500
rect 2050 410 2150 420
rect 2250 500 2350 510
rect 2250 420 2260 500
rect 2340 420 2350 500
rect 2250 410 2350 420
rect 2450 500 2550 510
rect 2450 420 2460 500
rect 2540 420 2550 500
rect 2450 410 2550 420
rect 2650 500 2750 510
rect 2650 420 2660 500
rect 2740 420 2750 500
rect 2650 410 2750 420
rect 2850 500 2950 510
rect 2850 420 2860 500
rect 2940 420 2950 500
rect 2850 410 2950 420
rect 3050 500 3150 510
rect 3050 420 3060 500
rect 3140 420 3150 500
rect 3050 410 3150 420
rect 3250 500 3350 510
rect 3250 420 3260 500
rect 3340 420 3350 500
rect 3250 410 3350 420
rect 3450 500 3550 510
rect 3450 420 3460 500
rect 3540 420 3550 500
rect 3450 410 3550 420
rect 3650 500 3750 510
rect 3650 420 3660 500
rect 3740 420 3750 500
rect 3650 410 3750 420
rect 3850 500 3950 510
rect 3850 420 3860 500
rect 3940 420 3950 500
rect 3850 410 3950 420
rect 4050 500 4150 510
rect 4050 420 4060 500
rect 4140 420 4150 500
rect 4050 410 4150 420
rect 4250 500 4350 510
rect 4250 420 4260 500
rect 4340 420 4350 500
rect 4250 410 4350 420
rect 4450 500 4550 510
rect 4450 420 4460 500
rect 4540 420 4550 500
rect 4450 410 4550 420
rect 4650 500 4750 510
rect 4650 420 4660 500
rect 4740 420 4750 500
rect 4650 410 4750 420
rect 4850 500 4950 510
rect 4850 420 4860 500
rect 4940 420 4950 500
rect 4850 410 4950 420
rect 5050 500 5150 510
rect 5050 420 5060 500
rect 5140 420 5150 500
rect 5050 410 5150 420
rect 5250 500 5350 510
rect 5250 420 5260 500
rect 5340 420 5350 500
rect 5250 410 5350 420
rect 5450 500 5550 510
rect 5450 420 5460 500
rect 5540 420 5550 500
rect 5450 410 5550 420
rect 5650 500 5750 510
rect 5650 420 5660 500
rect 5740 420 5750 500
rect 5650 410 5750 420
rect 5850 500 5950 510
rect 5850 420 5860 500
rect 5940 420 5950 500
rect 5850 410 5950 420
rect 6050 500 6150 510
rect 6050 420 6060 500
rect 6140 420 6150 500
rect 6050 410 6150 420
rect 6250 500 6350 510
rect 6250 420 6260 500
rect 6340 420 6350 500
rect 6250 410 6350 420
rect 6450 500 6550 510
rect 6450 420 6460 500
rect 6540 420 6550 500
rect 6450 410 6550 420
rect -150 315 -50 325
rect -150 235 -140 315
rect -60 235 -50 315
rect -150 225 -50 235
rect 50 315 150 325
rect 50 235 60 315
rect 140 235 150 315
rect 50 225 150 235
rect 250 315 350 325
rect 250 235 260 315
rect 340 235 350 315
rect 250 225 350 235
rect 450 315 550 325
rect 450 235 460 315
rect 540 235 550 315
rect 450 225 550 235
rect 650 315 750 325
rect 650 235 660 315
rect 740 235 750 315
rect 650 225 750 235
rect 850 315 950 325
rect 850 235 860 315
rect 940 235 950 315
rect 850 225 950 235
rect 1050 315 1150 325
rect 1050 235 1060 315
rect 1140 235 1150 315
rect 1050 225 1150 235
rect 1250 315 1350 325
rect 1250 235 1260 315
rect 1340 235 1350 315
rect 1250 225 1350 235
rect 1450 315 1550 325
rect 1450 235 1460 315
rect 1540 235 1550 315
rect 1450 225 1550 235
rect 1650 315 1750 325
rect 1650 235 1660 315
rect 1740 235 1750 315
rect 1650 225 1750 235
rect 1850 315 1950 325
rect 1850 235 1860 315
rect 1940 235 1950 315
rect 1850 225 1950 235
rect 2050 315 2150 325
rect 2050 235 2060 315
rect 2140 235 2150 315
rect 2050 225 2150 235
rect 2250 315 2350 325
rect 2250 235 2260 315
rect 2340 235 2350 315
rect 2250 225 2350 235
rect 2450 315 2550 325
rect 2450 235 2460 315
rect 2540 235 2550 315
rect 2450 225 2550 235
rect 2650 315 2750 325
rect 2650 235 2660 315
rect 2740 235 2750 315
rect 2650 225 2750 235
rect 2850 315 2950 325
rect 2850 235 2860 315
rect 2940 235 2950 315
rect 2850 225 2950 235
rect 3050 315 3150 325
rect 3050 235 3060 315
rect 3140 235 3150 315
rect 3050 225 3150 235
rect 3250 315 3350 325
rect 3250 235 3260 315
rect 3340 235 3350 315
rect 3250 225 3350 235
rect 3450 315 3550 325
rect 3450 235 3460 315
rect 3540 235 3550 315
rect 3450 225 3550 235
rect 3650 315 3750 325
rect 3650 235 3660 315
rect 3740 235 3750 315
rect 3650 225 3750 235
rect 3850 315 3950 325
rect 3850 235 3860 315
rect 3940 235 3950 315
rect 3850 225 3950 235
rect 4050 315 4150 325
rect 4050 235 4060 315
rect 4140 235 4150 315
rect 4050 225 4150 235
rect 4250 315 4350 325
rect 4250 235 4260 315
rect 4340 235 4350 315
rect 4250 225 4350 235
rect 4450 315 4550 325
rect 4450 235 4460 315
rect 4540 235 4550 315
rect 4450 225 4550 235
rect 4650 315 4750 325
rect 4650 235 4660 315
rect 4740 235 4750 315
rect 4650 225 4750 235
rect 4850 315 4950 325
rect 4850 235 4860 315
rect 4940 235 4950 315
rect 4850 225 4950 235
rect 5050 315 5150 325
rect 5050 235 5060 315
rect 5140 235 5150 315
rect 5050 225 5150 235
rect 5250 315 5350 325
rect 5250 235 5260 315
rect 5340 235 5350 315
rect 5250 225 5350 235
rect 5450 315 5550 325
rect 5450 235 5460 315
rect 5540 235 5550 315
rect 5450 225 5550 235
rect 5650 315 5750 325
rect 5650 235 5660 315
rect 5740 235 5750 315
rect 5650 225 5750 235
rect 5850 315 5950 325
rect 5850 235 5860 315
rect 5940 235 5950 315
rect 5850 225 5950 235
rect 6050 315 6150 325
rect 6050 235 6060 315
rect 6140 235 6150 315
rect 6050 225 6150 235
rect 6250 315 6350 325
rect 6250 235 6260 315
rect 6340 235 6350 315
rect 6250 225 6350 235
rect 6450 315 6550 325
rect 6450 235 6460 315
rect 6540 235 6550 315
rect 6450 225 6550 235
rect -150 130 -50 140
rect -150 50 -140 130
rect -60 50 -50 130
rect -150 40 -50 50
rect 50 130 150 140
rect 50 50 60 130
rect 140 50 150 130
rect 50 40 150 50
rect 250 130 350 140
rect 250 50 260 130
rect 340 50 350 130
rect 250 40 350 50
rect 450 130 550 140
rect 450 50 460 130
rect 540 50 550 130
rect 450 40 550 50
rect 650 130 750 140
rect 650 50 660 130
rect 740 50 750 130
rect 650 40 750 50
rect 850 130 950 140
rect 850 50 860 130
rect 940 50 950 130
rect 850 40 950 50
rect 1050 130 1150 140
rect 1050 50 1060 130
rect 1140 50 1150 130
rect 1050 40 1150 50
rect 1250 130 1350 140
rect 1250 50 1260 130
rect 1340 50 1350 130
rect 1250 40 1350 50
rect 1450 130 1550 140
rect 1450 50 1460 130
rect 1540 50 1550 130
rect 1450 40 1550 50
rect 1650 130 1750 140
rect 1650 50 1660 130
rect 1740 50 1750 130
rect 1650 40 1750 50
rect 1850 130 1950 140
rect 1850 50 1860 130
rect 1940 50 1950 130
rect 1850 40 1950 50
rect 2050 130 2150 140
rect 2050 50 2060 130
rect 2140 50 2150 130
rect 2050 40 2150 50
rect 2250 130 2350 140
rect 2250 50 2260 130
rect 2340 50 2350 130
rect 2250 40 2350 50
rect 2450 130 2550 140
rect 2450 50 2460 130
rect 2540 50 2550 130
rect 2450 40 2550 50
rect 2650 130 2750 140
rect 2650 50 2660 130
rect 2740 50 2750 130
rect 2650 40 2750 50
rect 2850 130 2950 140
rect 2850 50 2860 130
rect 2940 50 2950 130
rect 2850 40 2950 50
rect 3050 130 3150 140
rect 3050 50 3060 130
rect 3140 50 3150 130
rect 3050 40 3150 50
rect 3250 130 3350 140
rect 3250 50 3260 130
rect 3340 50 3350 130
rect 3250 40 3350 50
rect 3450 130 3550 140
rect 3450 50 3460 130
rect 3540 50 3550 130
rect 3450 40 3550 50
rect 3650 130 3750 140
rect 3650 50 3660 130
rect 3740 50 3750 130
rect 3650 40 3750 50
rect 3850 130 3950 140
rect 3850 50 3860 130
rect 3940 50 3950 130
rect 3850 40 3950 50
rect 4050 130 4150 140
rect 4050 50 4060 130
rect 4140 50 4150 130
rect 4050 40 4150 50
rect 4250 130 4350 140
rect 4250 50 4260 130
rect 4340 50 4350 130
rect 4250 40 4350 50
rect 4450 130 4550 140
rect 4450 50 4460 130
rect 4540 50 4550 130
rect 4450 40 4550 50
rect 4650 130 4750 140
rect 4650 50 4660 130
rect 4740 50 4750 130
rect 4650 40 4750 50
rect 4850 130 4950 140
rect 4850 50 4860 130
rect 4940 50 4950 130
rect 4850 40 4950 50
rect 5050 130 5150 140
rect 5050 50 5060 130
rect 5140 50 5150 130
rect 5050 40 5150 50
rect 5250 130 5350 140
rect 5250 50 5260 130
rect 5340 50 5350 130
rect 5250 40 5350 50
rect 5450 130 5550 140
rect 5450 50 5460 130
rect 5540 50 5550 130
rect 5450 40 5550 50
rect 5650 130 5750 140
rect 5650 50 5660 130
rect 5740 50 5750 130
rect 5650 40 5750 50
rect 5850 130 5950 140
rect 5850 50 5860 130
rect 5940 50 5950 130
rect 5850 40 5950 50
rect 6050 130 6150 140
rect 6050 50 6060 130
rect 6140 50 6150 130
rect 6050 40 6150 50
rect 6250 130 6350 140
rect 6250 50 6260 130
rect 6340 50 6350 130
rect 6250 40 6350 50
rect 6450 130 6550 140
rect 6450 50 6460 130
rect 6540 50 6550 130
rect 6450 40 6550 50
rect -150 -55 -50 -45
rect -150 -135 -140 -55
rect -60 -135 -50 -55
rect -150 -145 -50 -135
rect 50 -55 150 -45
rect 50 -135 60 -55
rect 140 -135 150 -55
rect 50 -145 150 -135
rect 250 -55 350 -45
rect 250 -135 260 -55
rect 340 -135 350 -55
rect 250 -145 350 -135
rect 450 -55 550 -45
rect 450 -135 460 -55
rect 540 -135 550 -55
rect 450 -145 550 -135
rect 650 -55 750 -45
rect 650 -135 660 -55
rect 740 -135 750 -55
rect 650 -145 750 -135
rect 850 -55 950 -45
rect 850 -135 860 -55
rect 940 -135 950 -55
rect 850 -145 950 -135
rect 1050 -55 1150 -45
rect 1050 -135 1060 -55
rect 1140 -135 1150 -55
rect 1050 -145 1150 -135
rect 1250 -55 1350 -45
rect 1250 -135 1260 -55
rect 1340 -135 1350 -55
rect 1250 -145 1350 -135
rect 1450 -55 1550 -45
rect 1450 -135 1460 -55
rect 1540 -135 1550 -55
rect 1450 -145 1550 -135
rect 1650 -55 1750 -45
rect 1650 -135 1660 -55
rect 1740 -135 1750 -55
rect 1650 -145 1750 -135
rect 1850 -55 1950 -45
rect 1850 -135 1860 -55
rect 1940 -135 1950 -55
rect 1850 -145 1950 -135
rect 2050 -55 2150 -45
rect 2050 -135 2060 -55
rect 2140 -135 2150 -55
rect 2050 -145 2150 -135
rect 2250 -55 2350 -45
rect 2250 -135 2260 -55
rect 2340 -135 2350 -55
rect 2250 -145 2350 -135
rect 2450 -55 2550 -45
rect 2450 -135 2460 -55
rect 2540 -135 2550 -55
rect 2450 -145 2550 -135
rect 2650 -55 2750 -45
rect 2650 -135 2660 -55
rect 2740 -135 2750 -55
rect 2650 -145 2750 -135
rect 2850 -55 2950 -45
rect 2850 -135 2860 -55
rect 2940 -135 2950 -55
rect 2850 -145 2950 -135
rect 3050 -55 3150 -45
rect 3050 -135 3060 -55
rect 3140 -135 3150 -55
rect 3050 -145 3150 -135
rect 3250 -55 3350 -45
rect 3250 -135 3260 -55
rect 3340 -135 3350 -55
rect 3250 -145 3350 -135
rect 3450 -55 3550 -45
rect 3450 -135 3460 -55
rect 3540 -135 3550 -55
rect 3450 -145 3550 -135
rect 3650 -55 3750 -45
rect 3650 -135 3660 -55
rect 3740 -135 3750 -55
rect 3650 -145 3750 -135
rect 3850 -55 3950 -45
rect 3850 -135 3860 -55
rect 3940 -135 3950 -55
rect 3850 -145 3950 -135
rect 4050 -55 4150 -45
rect 4050 -135 4060 -55
rect 4140 -135 4150 -55
rect 4050 -145 4150 -135
rect 4250 -55 4350 -45
rect 4250 -135 4260 -55
rect 4340 -135 4350 -55
rect 4250 -145 4350 -135
rect 4450 -55 4550 -45
rect 4450 -135 4460 -55
rect 4540 -135 4550 -55
rect 4450 -145 4550 -135
rect 4650 -55 4750 -45
rect 4650 -135 4660 -55
rect 4740 -135 4750 -55
rect 4650 -145 4750 -135
rect 4850 -55 4950 -45
rect 4850 -135 4860 -55
rect 4940 -135 4950 -55
rect 4850 -145 4950 -135
rect 5050 -55 5150 -45
rect 5050 -135 5060 -55
rect 5140 -135 5150 -55
rect 5050 -145 5150 -135
rect 5250 -55 5350 -45
rect 5250 -135 5260 -55
rect 5340 -135 5350 -55
rect 5250 -145 5350 -135
rect 5450 -55 5550 -45
rect 5450 -135 5460 -55
rect 5540 -135 5550 -55
rect 5450 -145 5550 -135
rect 5650 -55 5750 -45
rect 5650 -135 5660 -55
rect 5740 -135 5750 -55
rect 5650 -145 5750 -135
rect 5850 -55 5950 -45
rect 5850 -135 5860 -55
rect 5940 -135 5950 -55
rect 5850 -145 5950 -135
rect 6050 -55 6150 -45
rect 6050 -135 6060 -55
rect 6140 -135 6150 -55
rect 6050 -145 6150 -135
rect 6250 -55 6350 -45
rect 6250 -135 6260 -55
rect 6340 -135 6350 -55
rect 6250 -145 6350 -135
rect 6450 -55 6550 -45
rect 6450 -135 6460 -55
rect 6540 -135 6550 -55
rect 6450 -145 6550 -135
<< mimcapcontact >>
rect -140 11890 -60 11970
rect 60 11890 140 11970
rect 260 11890 340 11970
rect 460 11890 540 11970
rect 660 11890 740 11970
rect 860 11890 940 11970
rect 1060 11890 1140 11970
rect 1260 11890 1340 11970
rect 1460 11890 1540 11970
rect 1660 11890 1740 11970
rect 1860 11890 1940 11970
rect 2060 11890 2140 11970
rect 2260 11890 2340 11970
rect 2460 11890 2540 11970
rect 2660 11890 2740 11970
rect 2860 11890 2940 11970
rect 3060 11890 3140 11970
rect 3260 11890 3340 11970
rect 3460 11890 3540 11970
rect 3660 11890 3740 11970
rect 3860 11890 3940 11970
rect 4060 11890 4140 11970
rect 4260 11890 4340 11970
rect 4460 11890 4540 11970
rect 4660 11890 4740 11970
rect 4860 11890 4940 11970
rect 5060 11890 5140 11970
rect 5260 11890 5340 11970
rect 5460 11890 5540 11970
rect 5660 11890 5740 11970
rect 5860 11890 5940 11970
rect 6060 11890 6140 11970
rect 6260 11890 6340 11970
rect 6460 11890 6540 11970
rect -140 11705 -60 11785
rect 60 11705 140 11785
rect 260 11705 340 11785
rect 460 11705 540 11785
rect 660 11705 740 11785
rect 860 11705 940 11785
rect 1060 11705 1140 11785
rect 1260 11705 1340 11785
rect 1460 11705 1540 11785
rect 1660 11705 1740 11785
rect 1860 11705 1940 11785
rect 2060 11705 2140 11785
rect 2260 11705 2340 11785
rect 2460 11705 2540 11785
rect 2660 11705 2740 11785
rect 2860 11705 2940 11785
rect 3060 11705 3140 11785
rect 3260 11705 3340 11785
rect 3460 11705 3540 11785
rect 3660 11705 3740 11785
rect 3860 11705 3940 11785
rect 4060 11705 4140 11785
rect 4260 11705 4340 11785
rect 4460 11705 4540 11785
rect 4660 11705 4740 11785
rect 4860 11705 4940 11785
rect 5060 11705 5140 11785
rect 5260 11705 5340 11785
rect 5460 11705 5540 11785
rect 5660 11705 5740 11785
rect 5860 11705 5940 11785
rect 6060 11705 6140 11785
rect 6260 11705 6340 11785
rect 6460 11705 6540 11785
rect -140 11520 -60 11600
rect 60 11520 140 11600
rect 260 11520 340 11600
rect 460 11520 540 11600
rect 660 11520 740 11600
rect 860 11520 940 11600
rect 1060 11520 1140 11600
rect 1260 11520 1340 11600
rect 1460 11520 1540 11600
rect 1660 11520 1740 11600
rect 1860 11520 1940 11600
rect 2060 11520 2140 11600
rect 2260 11520 2340 11600
rect 2460 11520 2540 11600
rect 2660 11520 2740 11600
rect 2860 11520 2940 11600
rect 3060 11520 3140 11600
rect 3260 11520 3340 11600
rect 3460 11520 3540 11600
rect 3660 11520 3740 11600
rect 3860 11520 3940 11600
rect 4060 11520 4140 11600
rect 4260 11520 4340 11600
rect 4460 11520 4540 11600
rect 4660 11520 4740 11600
rect 4860 11520 4940 11600
rect 5060 11520 5140 11600
rect 5260 11520 5340 11600
rect 5460 11520 5540 11600
rect 5660 11520 5740 11600
rect 5860 11520 5940 11600
rect 6060 11520 6140 11600
rect 6260 11520 6340 11600
rect 6460 11520 6540 11600
rect -140 11335 -60 11415
rect 60 11335 140 11415
rect 260 11335 340 11415
rect 460 11335 540 11415
rect 660 11335 740 11415
rect 860 11335 940 11415
rect 1060 11335 1140 11415
rect 1260 11335 1340 11415
rect 1460 11335 1540 11415
rect 1660 11335 1740 11415
rect 1860 11335 1940 11415
rect 2060 11335 2140 11415
rect 2260 11335 2340 11415
rect 2460 11335 2540 11415
rect 2660 11335 2740 11415
rect 2860 11335 2940 11415
rect 3060 11335 3140 11415
rect 3260 11335 3340 11415
rect 3460 11335 3540 11415
rect 3660 11335 3740 11415
rect 3860 11335 3940 11415
rect 4060 11335 4140 11415
rect 4260 11335 4340 11415
rect 4460 11335 4540 11415
rect 4660 11335 4740 11415
rect 4860 11335 4940 11415
rect 5060 11335 5140 11415
rect 5260 11335 5340 11415
rect 5460 11335 5540 11415
rect 5660 11335 5740 11415
rect 5860 11335 5940 11415
rect 6060 11335 6140 11415
rect 6260 11335 6340 11415
rect 6460 11335 6540 11415
rect -140 11150 -60 11230
rect 60 11150 140 11230
rect 260 11150 340 11230
rect 460 11150 540 11230
rect 660 11150 740 11230
rect 860 11150 940 11230
rect 1060 11150 1140 11230
rect 1260 11150 1340 11230
rect 1460 11150 1540 11230
rect 1660 11150 1740 11230
rect 1860 11150 1940 11230
rect 2060 11150 2140 11230
rect 2260 11150 2340 11230
rect 2460 11150 2540 11230
rect 2660 11150 2740 11230
rect 2860 11150 2940 11230
rect 3060 11150 3140 11230
rect 3260 11150 3340 11230
rect 3460 11150 3540 11230
rect 3660 11150 3740 11230
rect 3860 11150 3940 11230
rect 4060 11150 4140 11230
rect 4260 11150 4340 11230
rect 4460 11150 4540 11230
rect 4660 11150 4740 11230
rect 4860 11150 4940 11230
rect 5060 11150 5140 11230
rect 5260 11150 5340 11230
rect 5460 11150 5540 11230
rect 5660 11150 5740 11230
rect 5860 11150 5940 11230
rect 6060 11150 6140 11230
rect 6260 11150 6340 11230
rect 6460 11150 6540 11230
rect -140 10965 -60 11045
rect 60 10965 140 11045
rect 260 10965 340 11045
rect 460 10965 540 11045
rect 660 10965 740 11045
rect 860 10965 940 11045
rect 1060 10965 1140 11045
rect 1260 10965 1340 11045
rect 1460 10965 1540 11045
rect 1660 10965 1740 11045
rect 1860 10965 1940 11045
rect 2060 10965 2140 11045
rect 2260 10965 2340 11045
rect 2460 10965 2540 11045
rect 2660 10965 2740 11045
rect 2860 10965 2940 11045
rect 3060 10965 3140 11045
rect 3260 10965 3340 11045
rect 3460 10965 3540 11045
rect 3660 10965 3740 11045
rect 3860 10965 3940 11045
rect 4060 10965 4140 11045
rect 4260 10965 4340 11045
rect 4460 10965 4540 11045
rect 4660 10965 4740 11045
rect 4860 10965 4940 11045
rect 5060 10965 5140 11045
rect 5260 10965 5340 11045
rect 5460 10965 5540 11045
rect 5660 10965 5740 11045
rect 5860 10965 5940 11045
rect 6060 10965 6140 11045
rect 6260 10965 6340 11045
rect 6460 10965 6540 11045
rect -140 10780 -60 10860
rect 60 10780 140 10860
rect 260 10780 340 10860
rect 460 10780 540 10860
rect 660 10780 740 10860
rect 860 10780 940 10860
rect 1060 10780 1140 10860
rect 1260 10780 1340 10860
rect 1460 10780 1540 10860
rect 1660 10780 1740 10860
rect 1860 10780 1940 10860
rect 2060 10780 2140 10860
rect 2260 10780 2340 10860
rect 2460 10780 2540 10860
rect 2660 10780 2740 10860
rect 2860 10780 2940 10860
rect 3060 10780 3140 10860
rect 3260 10780 3340 10860
rect 3460 10780 3540 10860
rect 3660 10780 3740 10860
rect 3860 10780 3940 10860
rect 4060 10780 4140 10860
rect 4260 10780 4340 10860
rect 4460 10780 4540 10860
rect 4660 10780 4740 10860
rect 4860 10780 4940 10860
rect 5060 10780 5140 10860
rect 5260 10780 5340 10860
rect 5460 10780 5540 10860
rect 5660 10780 5740 10860
rect 5860 10780 5940 10860
rect 6060 10780 6140 10860
rect 6260 10780 6340 10860
rect 6460 10780 6540 10860
rect -140 10595 -60 10675
rect 60 10595 140 10675
rect 260 10595 340 10675
rect 460 10595 540 10675
rect 660 10595 740 10675
rect 860 10595 940 10675
rect 1060 10595 1140 10675
rect 1260 10595 1340 10675
rect 1460 10595 1540 10675
rect 1660 10595 1740 10675
rect 1860 10595 1940 10675
rect 2060 10595 2140 10675
rect 2260 10595 2340 10675
rect 2460 10595 2540 10675
rect 2660 10595 2740 10675
rect 2860 10595 2940 10675
rect 3060 10595 3140 10675
rect 3260 10595 3340 10675
rect 3460 10595 3540 10675
rect 3660 10595 3740 10675
rect 3860 10595 3940 10675
rect 4060 10595 4140 10675
rect 4260 10595 4340 10675
rect 4460 10595 4540 10675
rect 4660 10595 4740 10675
rect 4860 10595 4940 10675
rect 5060 10595 5140 10675
rect 5260 10595 5340 10675
rect 5460 10595 5540 10675
rect 5660 10595 5740 10675
rect 5860 10595 5940 10675
rect 6060 10595 6140 10675
rect 6260 10595 6340 10675
rect 6460 10595 6540 10675
rect -140 10410 -60 10490
rect 60 10410 140 10490
rect 260 10410 340 10490
rect 460 10410 540 10490
rect 660 10410 740 10490
rect 860 10410 940 10490
rect 1060 10410 1140 10490
rect 1260 10410 1340 10490
rect 1460 10410 1540 10490
rect 1660 10410 1740 10490
rect 1860 10410 1940 10490
rect 2060 10410 2140 10490
rect 2260 10410 2340 10490
rect 2460 10410 2540 10490
rect 2660 10410 2740 10490
rect 2860 10410 2940 10490
rect 3060 10410 3140 10490
rect 3260 10410 3340 10490
rect 3460 10410 3540 10490
rect 3660 10410 3740 10490
rect 3860 10410 3940 10490
rect 4060 10410 4140 10490
rect 4260 10410 4340 10490
rect 4460 10410 4540 10490
rect 4660 10410 4740 10490
rect 4860 10410 4940 10490
rect 5060 10410 5140 10490
rect 5260 10410 5340 10490
rect 5460 10410 5540 10490
rect 5660 10410 5740 10490
rect 5860 10410 5940 10490
rect 6060 10410 6140 10490
rect 6260 10410 6340 10490
rect 6460 10410 6540 10490
rect -140 10225 -60 10305
rect 60 10225 140 10305
rect 260 10225 340 10305
rect 460 10225 540 10305
rect 660 10225 740 10305
rect 860 10225 940 10305
rect 1060 10225 1140 10305
rect 1260 10225 1340 10305
rect 1460 10225 1540 10305
rect 1660 10225 1740 10305
rect 1860 10225 1940 10305
rect 2060 10225 2140 10305
rect 2260 10225 2340 10305
rect 2460 10225 2540 10305
rect 2660 10225 2740 10305
rect 2860 10225 2940 10305
rect 3060 10225 3140 10305
rect 3260 10225 3340 10305
rect 3460 10225 3540 10305
rect 3660 10225 3740 10305
rect 3860 10225 3940 10305
rect 4060 10225 4140 10305
rect 4260 10225 4340 10305
rect 4460 10225 4540 10305
rect 4660 10225 4740 10305
rect 4860 10225 4940 10305
rect 5060 10225 5140 10305
rect 5260 10225 5340 10305
rect 5460 10225 5540 10305
rect 5660 10225 5740 10305
rect 5860 10225 5940 10305
rect 6060 10225 6140 10305
rect 6260 10225 6340 10305
rect 6460 10225 6540 10305
rect -140 10040 -60 10120
rect 60 10040 140 10120
rect 260 10040 340 10120
rect 460 10040 540 10120
rect 660 10040 740 10120
rect 860 10040 940 10120
rect 1060 10040 1140 10120
rect 1260 10040 1340 10120
rect 1460 10040 1540 10120
rect 1660 10040 1740 10120
rect 1860 10040 1940 10120
rect 2060 10040 2140 10120
rect 2260 10040 2340 10120
rect 2460 10040 2540 10120
rect 2660 10040 2740 10120
rect 2860 10040 2940 10120
rect 3060 10040 3140 10120
rect 3260 10040 3340 10120
rect 3460 10040 3540 10120
rect 3660 10040 3740 10120
rect 3860 10040 3940 10120
rect 4060 10040 4140 10120
rect 4260 10040 4340 10120
rect 4460 10040 4540 10120
rect 4660 10040 4740 10120
rect 4860 10040 4940 10120
rect 5060 10040 5140 10120
rect 5260 10040 5340 10120
rect 5460 10040 5540 10120
rect 5660 10040 5740 10120
rect 5860 10040 5940 10120
rect 6060 10040 6140 10120
rect 6260 10040 6340 10120
rect 6460 10040 6540 10120
rect -140 9855 -60 9935
rect 60 9855 140 9935
rect 260 9855 340 9935
rect 460 9855 540 9935
rect 660 9855 740 9935
rect 860 9855 940 9935
rect 1060 9855 1140 9935
rect 1260 9855 1340 9935
rect 1460 9855 1540 9935
rect 1660 9855 1740 9935
rect 1860 9855 1940 9935
rect 2060 9855 2140 9935
rect 2260 9855 2340 9935
rect 2460 9855 2540 9935
rect 2660 9855 2740 9935
rect 2860 9855 2940 9935
rect 3060 9855 3140 9935
rect 3260 9855 3340 9935
rect 3460 9855 3540 9935
rect 3660 9855 3740 9935
rect 3860 9855 3940 9935
rect 4060 9855 4140 9935
rect 4260 9855 4340 9935
rect 4460 9855 4540 9935
rect 4660 9855 4740 9935
rect 4860 9855 4940 9935
rect 5060 9855 5140 9935
rect 5260 9855 5340 9935
rect 5460 9855 5540 9935
rect 5660 9855 5740 9935
rect 5860 9855 5940 9935
rect 6060 9855 6140 9935
rect 6260 9855 6340 9935
rect 6460 9855 6540 9935
rect -140 9670 -60 9750
rect 60 9670 140 9750
rect 260 9670 340 9750
rect 460 9670 540 9750
rect 660 9670 740 9750
rect 860 9670 940 9750
rect 1060 9670 1140 9750
rect 1260 9670 1340 9750
rect 1460 9670 1540 9750
rect 1660 9670 1740 9750
rect 1860 9670 1940 9750
rect 2060 9670 2140 9750
rect 2260 9670 2340 9750
rect 2460 9670 2540 9750
rect 2660 9670 2740 9750
rect 2860 9670 2940 9750
rect 3060 9670 3140 9750
rect 3260 9670 3340 9750
rect 3460 9670 3540 9750
rect 3660 9670 3740 9750
rect 3860 9670 3940 9750
rect 4060 9670 4140 9750
rect 4260 9670 4340 9750
rect 4460 9670 4540 9750
rect 4660 9670 4740 9750
rect 4860 9670 4940 9750
rect 5060 9670 5140 9750
rect 5260 9670 5340 9750
rect 5460 9670 5540 9750
rect 5660 9670 5740 9750
rect 5860 9670 5940 9750
rect 6060 9670 6140 9750
rect 6260 9670 6340 9750
rect 6460 9670 6540 9750
rect -140 9485 -60 9565
rect 60 9485 140 9565
rect 260 9485 340 9565
rect 460 9485 540 9565
rect 660 9485 740 9565
rect 860 9485 940 9565
rect 1060 9485 1140 9565
rect 1260 9485 1340 9565
rect 1460 9485 1540 9565
rect 1660 9485 1740 9565
rect 1860 9485 1940 9565
rect 2060 9485 2140 9565
rect 2260 9485 2340 9565
rect 2460 9485 2540 9565
rect 2660 9485 2740 9565
rect 2860 9485 2940 9565
rect 3060 9485 3140 9565
rect 3260 9485 3340 9565
rect 3460 9485 3540 9565
rect 3660 9485 3740 9565
rect 3860 9485 3940 9565
rect 4060 9485 4140 9565
rect 4260 9485 4340 9565
rect 4460 9485 4540 9565
rect 4660 9485 4740 9565
rect 4860 9485 4940 9565
rect 5060 9485 5140 9565
rect 5260 9485 5340 9565
rect 5460 9485 5540 9565
rect 5660 9485 5740 9565
rect 5860 9485 5940 9565
rect 6060 9485 6140 9565
rect 6260 9485 6340 9565
rect 6460 9485 6540 9565
rect -140 9300 -60 9380
rect 60 9300 140 9380
rect 260 9300 340 9380
rect 460 9300 540 9380
rect 660 9300 740 9380
rect 860 9300 940 9380
rect 1060 9300 1140 9380
rect 1260 9300 1340 9380
rect 1460 9300 1540 9380
rect 1660 9300 1740 9380
rect 1860 9300 1940 9380
rect 2060 9300 2140 9380
rect 2260 9300 2340 9380
rect 2460 9300 2540 9380
rect 2660 9300 2740 9380
rect 2860 9300 2940 9380
rect 3060 9300 3140 9380
rect 3260 9300 3340 9380
rect 3460 9300 3540 9380
rect 3660 9300 3740 9380
rect 3860 9300 3940 9380
rect 4060 9300 4140 9380
rect 4260 9300 4340 9380
rect 4460 9300 4540 9380
rect 4660 9300 4740 9380
rect 4860 9300 4940 9380
rect 5060 9300 5140 9380
rect 5260 9300 5340 9380
rect 5460 9300 5540 9380
rect 5660 9300 5740 9380
rect 5860 9300 5940 9380
rect 6060 9300 6140 9380
rect 6260 9300 6340 9380
rect 6460 9300 6540 9380
rect -140 9115 -60 9195
rect 60 9115 140 9195
rect 260 9115 340 9195
rect 460 9115 540 9195
rect 660 9115 740 9195
rect 860 9115 940 9195
rect 1060 9115 1140 9195
rect 1260 9115 1340 9195
rect 1460 9115 1540 9195
rect 1660 9115 1740 9195
rect 1860 9115 1940 9195
rect 2060 9115 2140 9195
rect 2260 9115 2340 9195
rect 2460 9115 2540 9195
rect 2660 9115 2740 9195
rect 2860 9115 2940 9195
rect 3060 9115 3140 9195
rect 3260 9115 3340 9195
rect 3460 9115 3540 9195
rect 3660 9115 3740 9195
rect 3860 9115 3940 9195
rect 4060 9115 4140 9195
rect 4260 9115 4340 9195
rect 4460 9115 4540 9195
rect 4660 9115 4740 9195
rect 4860 9115 4940 9195
rect 5060 9115 5140 9195
rect 5260 9115 5340 9195
rect 5460 9115 5540 9195
rect 5660 9115 5740 9195
rect 5860 9115 5940 9195
rect 6060 9115 6140 9195
rect 6260 9115 6340 9195
rect 6460 9115 6540 9195
rect -140 8930 -60 9010
rect 60 8930 140 9010
rect 260 8930 340 9010
rect 460 8930 540 9010
rect 660 8930 740 9010
rect 860 8930 940 9010
rect 1060 8930 1140 9010
rect 1260 8930 1340 9010
rect 1460 8930 1540 9010
rect 1660 8930 1740 9010
rect 1860 8930 1940 9010
rect 2060 8930 2140 9010
rect 2260 8930 2340 9010
rect 2460 8930 2540 9010
rect 2660 8930 2740 9010
rect 2860 8930 2940 9010
rect 3060 8930 3140 9010
rect 3260 8930 3340 9010
rect 3460 8930 3540 9010
rect 3660 8930 3740 9010
rect 3860 8930 3940 9010
rect 4060 8930 4140 9010
rect 4260 8930 4340 9010
rect 4460 8930 4540 9010
rect 4660 8930 4740 9010
rect 4860 8930 4940 9010
rect 5060 8930 5140 9010
rect 5260 8930 5340 9010
rect 5460 8930 5540 9010
rect 5660 8930 5740 9010
rect 5860 8930 5940 9010
rect 6060 8930 6140 9010
rect 6260 8930 6340 9010
rect 6460 8930 6540 9010
rect -140 8745 -60 8825
rect 60 8745 140 8825
rect 260 8745 340 8825
rect 460 8745 540 8825
rect 660 8745 740 8825
rect 860 8745 940 8825
rect 1060 8745 1140 8825
rect 1260 8745 1340 8825
rect 1460 8745 1540 8825
rect 1660 8745 1740 8825
rect 1860 8745 1940 8825
rect 2060 8745 2140 8825
rect 2260 8745 2340 8825
rect 2460 8745 2540 8825
rect 2660 8745 2740 8825
rect 2860 8745 2940 8825
rect 3060 8745 3140 8825
rect 3260 8745 3340 8825
rect 3460 8745 3540 8825
rect 3660 8745 3740 8825
rect 3860 8745 3940 8825
rect 4060 8745 4140 8825
rect 4260 8745 4340 8825
rect 4460 8745 4540 8825
rect 4660 8745 4740 8825
rect 4860 8745 4940 8825
rect 5060 8745 5140 8825
rect 5260 8745 5340 8825
rect 5460 8745 5540 8825
rect 5660 8745 5740 8825
rect 5860 8745 5940 8825
rect 6060 8745 6140 8825
rect 6260 8745 6340 8825
rect 6460 8745 6540 8825
rect -140 8560 -60 8640
rect 60 8560 140 8640
rect 260 8560 340 8640
rect 460 8560 540 8640
rect 660 8560 740 8640
rect 860 8560 940 8640
rect 1060 8560 1140 8640
rect 1260 8560 1340 8640
rect 1460 8560 1540 8640
rect 1660 8560 1740 8640
rect 1860 8560 1940 8640
rect 2060 8560 2140 8640
rect 2260 8560 2340 8640
rect 2460 8560 2540 8640
rect 2660 8560 2740 8640
rect 2860 8560 2940 8640
rect 3060 8560 3140 8640
rect 3260 8560 3340 8640
rect 3460 8560 3540 8640
rect 3660 8560 3740 8640
rect 3860 8560 3940 8640
rect 4060 8560 4140 8640
rect 4260 8560 4340 8640
rect 4460 8560 4540 8640
rect 4660 8560 4740 8640
rect 4860 8560 4940 8640
rect 5060 8560 5140 8640
rect 5260 8560 5340 8640
rect 5460 8560 5540 8640
rect 5660 8560 5740 8640
rect 5860 8560 5940 8640
rect 6060 8560 6140 8640
rect 6260 8560 6340 8640
rect 6460 8560 6540 8640
rect -140 8375 -60 8455
rect 60 8375 140 8455
rect 260 8375 340 8455
rect 460 8375 540 8455
rect 660 8375 740 8455
rect 860 8375 940 8455
rect 1060 8375 1140 8455
rect 1260 8375 1340 8455
rect 1460 8375 1540 8455
rect 1660 8375 1740 8455
rect 1860 8375 1940 8455
rect 2060 8375 2140 8455
rect 2260 8375 2340 8455
rect 2460 8375 2540 8455
rect 2660 8375 2740 8455
rect 2860 8375 2940 8455
rect 3060 8375 3140 8455
rect 3260 8375 3340 8455
rect 3460 8375 3540 8455
rect 3660 8375 3740 8455
rect 3860 8375 3940 8455
rect 4060 8375 4140 8455
rect 4260 8375 4340 8455
rect 4460 8375 4540 8455
rect 4660 8375 4740 8455
rect 4860 8375 4940 8455
rect 5060 8375 5140 8455
rect 5260 8375 5340 8455
rect 5460 8375 5540 8455
rect 5660 8375 5740 8455
rect 5860 8375 5940 8455
rect 6060 8375 6140 8455
rect 6260 8375 6340 8455
rect 6460 8375 6540 8455
rect -140 8190 -60 8270
rect 60 8190 140 8270
rect 260 8190 340 8270
rect 460 8190 540 8270
rect 660 8190 740 8270
rect 860 8190 940 8270
rect 1060 8190 1140 8270
rect 1260 8190 1340 8270
rect 1460 8190 1540 8270
rect 1660 8190 1740 8270
rect 1860 8190 1940 8270
rect 2060 8190 2140 8270
rect 2260 8190 2340 8270
rect 2460 8190 2540 8270
rect 2660 8190 2740 8270
rect 2860 8190 2940 8270
rect 3060 8190 3140 8270
rect 3260 8190 3340 8270
rect 3460 8190 3540 8270
rect 3660 8190 3740 8270
rect 3860 8190 3940 8270
rect 4060 8190 4140 8270
rect 4260 8190 4340 8270
rect 4460 8190 4540 8270
rect 4660 8190 4740 8270
rect 4860 8190 4940 8270
rect 5060 8190 5140 8270
rect 5260 8190 5340 8270
rect 5460 8190 5540 8270
rect 5660 8190 5740 8270
rect 5860 8190 5940 8270
rect 6060 8190 6140 8270
rect 6260 8190 6340 8270
rect 6460 8190 6540 8270
rect -140 8005 -60 8085
rect 60 8005 140 8085
rect 260 8005 340 8085
rect 460 8005 540 8085
rect 660 8005 740 8085
rect 860 8005 940 8085
rect 1060 8005 1140 8085
rect 1260 8005 1340 8085
rect 1460 8005 1540 8085
rect 1660 8005 1740 8085
rect 1860 8005 1940 8085
rect 2060 8005 2140 8085
rect 2260 8005 2340 8085
rect 2460 8005 2540 8085
rect 2660 8005 2740 8085
rect 2860 8005 2940 8085
rect 3060 8005 3140 8085
rect 3260 8005 3340 8085
rect 3460 8005 3540 8085
rect 3660 8005 3740 8085
rect 3860 8005 3940 8085
rect 4060 8005 4140 8085
rect 4260 8005 4340 8085
rect 4460 8005 4540 8085
rect 4660 8005 4740 8085
rect 4860 8005 4940 8085
rect 5060 8005 5140 8085
rect 5260 8005 5340 8085
rect 5460 8005 5540 8085
rect 5660 8005 5740 8085
rect 5860 8005 5940 8085
rect 6060 8005 6140 8085
rect 6260 8005 6340 8085
rect 6460 8005 6540 8085
rect -140 7820 -60 7900
rect 60 7820 140 7900
rect 260 7820 340 7900
rect 460 7820 540 7900
rect 660 7820 740 7900
rect 860 7820 940 7900
rect 1060 7820 1140 7900
rect 1260 7820 1340 7900
rect 1460 7820 1540 7900
rect 1660 7820 1740 7900
rect 1860 7820 1940 7900
rect 2060 7820 2140 7900
rect 2260 7820 2340 7900
rect 2460 7820 2540 7900
rect 2660 7820 2740 7900
rect 2860 7820 2940 7900
rect 3060 7820 3140 7900
rect 3260 7820 3340 7900
rect 3460 7820 3540 7900
rect 3660 7820 3740 7900
rect 3860 7820 3940 7900
rect 4060 7820 4140 7900
rect 4260 7820 4340 7900
rect 4460 7820 4540 7900
rect 4660 7820 4740 7900
rect 4860 7820 4940 7900
rect 5060 7820 5140 7900
rect 5260 7820 5340 7900
rect 5460 7820 5540 7900
rect 5660 7820 5740 7900
rect 5860 7820 5940 7900
rect 6060 7820 6140 7900
rect 6260 7820 6340 7900
rect 6460 7820 6540 7900
rect -140 7635 -60 7715
rect 60 7635 140 7715
rect 260 7635 340 7715
rect 460 7635 540 7715
rect 660 7635 740 7715
rect 860 7635 940 7715
rect 1060 7635 1140 7715
rect 1260 7635 1340 7715
rect 1460 7635 1540 7715
rect 1660 7635 1740 7715
rect 1860 7635 1940 7715
rect 2060 7635 2140 7715
rect 2260 7635 2340 7715
rect 2460 7635 2540 7715
rect 2660 7635 2740 7715
rect 2860 7635 2940 7715
rect 3060 7635 3140 7715
rect 3260 7635 3340 7715
rect 3460 7635 3540 7715
rect 3660 7635 3740 7715
rect 3860 7635 3940 7715
rect 4060 7635 4140 7715
rect 4260 7635 4340 7715
rect 4460 7635 4540 7715
rect 4660 7635 4740 7715
rect 4860 7635 4940 7715
rect 5060 7635 5140 7715
rect 5260 7635 5340 7715
rect 5460 7635 5540 7715
rect 5660 7635 5740 7715
rect 5860 7635 5940 7715
rect 6060 7635 6140 7715
rect 6260 7635 6340 7715
rect 6460 7635 6540 7715
rect -140 7450 -60 7530
rect 60 7450 140 7530
rect 260 7450 340 7530
rect 460 7450 540 7530
rect 660 7450 740 7530
rect 860 7450 940 7530
rect 1060 7450 1140 7530
rect 1260 7450 1340 7530
rect 1460 7450 1540 7530
rect 1660 7450 1740 7530
rect 1860 7450 1940 7530
rect 2060 7450 2140 7530
rect 2260 7450 2340 7530
rect 2460 7450 2540 7530
rect 2660 7450 2740 7530
rect 2860 7450 2940 7530
rect 3060 7450 3140 7530
rect 3260 7450 3340 7530
rect 3460 7450 3540 7530
rect 3660 7450 3740 7530
rect 3860 7450 3940 7530
rect 4060 7450 4140 7530
rect 4260 7450 4340 7530
rect 4460 7450 4540 7530
rect 4660 7450 4740 7530
rect 4860 7450 4940 7530
rect 5060 7450 5140 7530
rect 5260 7450 5340 7530
rect 5460 7450 5540 7530
rect 5660 7450 5740 7530
rect 5860 7450 5940 7530
rect 6060 7450 6140 7530
rect 6260 7450 6340 7530
rect 6460 7450 6540 7530
rect -140 7265 -60 7345
rect 60 7265 140 7345
rect 260 7265 340 7345
rect 460 7265 540 7345
rect 660 7265 740 7345
rect 860 7265 940 7345
rect 1060 7265 1140 7345
rect 1260 7265 1340 7345
rect 1460 7265 1540 7345
rect 1660 7265 1740 7345
rect 1860 7265 1940 7345
rect 2060 7265 2140 7345
rect 2260 7265 2340 7345
rect 2460 7265 2540 7345
rect 2660 7265 2740 7345
rect 2860 7265 2940 7345
rect 3060 7265 3140 7345
rect 3260 7265 3340 7345
rect 3460 7265 3540 7345
rect 3660 7265 3740 7345
rect 3860 7265 3940 7345
rect 4060 7265 4140 7345
rect 4260 7265 4340 7345
rect 4460 7265 4540 7345
rect 4660 7265 4740 7345
rect 4860 7265 4940 7345
rect 5060 7265 5140 7345
rect 5260 7265 5340 7345
rect 5460 7265 5540 7345
rect 5660 7265 5740 7345
rect 5860 7265 5940 7345
rect 6060 7265 6140 7345
rect 6260 7265 6340 7345
rect 6460 7265 6540 7345
rect -140 7080 -60 7160
rect 60 7080 140 7160
rect 260 7080 340 7160
rect 460 7080 540 7160
rect 660 7080 740 7160
rect 860 7080 940 7160
rect 1060 7080 1140 7160
rect 1260 7080 1340 7160
rect 1460 7080 1540 7160
rect 1660 7080 1740 7160
rect 1860 7080 1940 7160
rect 2060 7080 2140 7160
rect 2260 7080 2340 7160
rect 2460 7080 2540 7160
rect 2660 7080 2740 7160
rect 2860 7080 2940 7160
rect 3060 7080 3140 7160
rect 3260 7080 3340 7160
rect 3460 7080 3540 7160
rect 3660 7080 3740 7160
rect 3860 7080 3940 7160
rect 4060 7080 4140 7160
rect 4260 7080 4340 7160
rect 4460 7080 4540 7160
rect 4660 7080 4740 7160
rect 4860 7080 4940 7160
rect 5060 7080 5140 7160
rect 5260 7080 5340 7160
rect 5460 7080 5540 7160
rect 5660 7080 5740 7160
rect 5860 7080 5940 7160
rect 6060 7080 6140 7160
rect 6260 7080 6340 7160
rect 6460 7080 6540 7160
rect -140 6895 -60 6975
rect 60 6895 140 6975
rect 260 6895 340 6975
rect 460 6895 540 6975
rect 660 6895 740 6975
rect 860 6895 940 6975
rect 1060 6895 1140 6975
rect 1260 6895 1340 6975
rect 1460 6895 1540 6975
rect 1660 6895 1740 6975
rect 1860 6895 1940 6975
rect 2060 6895 2140 6975
rect 2260 6895 2340 6975
rect 2460 6895 2540 6975
rect 2660 6895 2740 6975
rect 2860 6895 2940 6975
rect 3060 6895 3140 6975
rect 3260 6895 3340 6975
rect 3460 6895 3540 6975
rect 3660 6895 3740 6975
rect 3860 6895 3940 6975
rect 4060 6895 4140 6975
rect 4260 6895 4340 6975
rect 4460 6895 4540 6975
rect 4660 6895 4740 6975
rect 4860 6895 4940 6975
rect 5060 6895 5140 6975
rect 5260 6895 5340 6975
rect 5460 6895 5540 6975
rect 5660 6895 5740 6975
rect 5860 6895 5940 6975
rect 6060 6895 6140 6975
rect 6260 6895 6340 6975
rect 6460 6895 6540 6975
rect -140 6710 -60 6790
rect 60 6710 140 6790
rect 260 6710 340 6790
rect 460 6710 540 6790
rect 660 6710 740 6790
rect 860 6710 940 6790
rect 1060 6710 1140 6790
rect 1260 6710 1340 6790
rect 1460 6710 1540 6790
rect 1660 6710 1740 6790
rect 1860 6710 1940 6790
rect 2060 6710 2140 6790
rect 2260 6710 2340 6790
rect 2460 6710 2540 6790
rect 2660 6710 2740 6790
rect 2860 6710 2940 6790
rect 3060 6710 3140 6790
rect 3260 6710 3340 6790
rect 3460 6710 3540 6790
rect 3660 6710 3740 6790
rect 3860 6710 3940 6790
rect 4060 6710 4140 6790
rect 4260 6710 4340 6790
rect 4460 6710 4540 6790
rect 4660 6710 4740 6790
rect 4860 6710 4940 6790
rect 5060 6710 5140 6790
rect 5260 6710 5340 6790
rect 5460 6710 5540 6790
rect 5660 6710 5740 6790
rect 5860 6710 5940 6790
rect 6060 6710 6140 6790
rect 6260 6710 6340 6790
rect 6460 6710 6540 6790
rect -140 6525 -60 6605
rect 60 6525 140 6605
rect 260 6525 340 6605
rect 460 6525 540 6605
rect 660 6525 740 6605
rect 860 6525 940 6605
rect 1060 6525 1140 6605
rect 1260 6525 1340 6605
rect 1460 6525 1540 6605
rect 1660 6525 1740 6605
rect 1860 6525 1940 6605
rect 2060 6525 2140 6605
rect 2260 6525 2340 6605
rect 2460 6525 2540 6605
rect 2660 6525 2740 6605
rect 2860 6525 2940 6605
rect 3060 6525 3140 6605
rect 3260 6525 3340 6605
rect 3460 6525 3540 6605
rect 3660 6525 3740 6605
rect 3860 6525 3940 6605
rect 4060 6525 4140 6605
rect 4260 6525 4340 6605
rect 4460 6525 4540 6605
rect 4660 6525 4740 6605
rect 4860 6525 4940 6605
rect 5060 6525 5140 6605
rect 5260 6525 5340 6605
rect 5460 6525 5540 6605
rect 5660 6525 5740 6605
rect 5860 6525 5940 6605
rect 6060 6525 6140 6605
rect 6260 6525 6340 6605
rect 6460 6525 6540 6605
rect -140 6340 -60 6420
rect 60 6340 140 6420
rect 260 6340 340 6420
rect 460 6340 540 6420
rect 660 6340 740 6420
rect 860 6340 940 6420
rect 1060 6340 1140 6420
rect 1260 6340 1340 6420
rect 1460 6340 1540 6420
rect 1660 6340 1740 6420
rect 1860 6340 1940 6420
rect 2060 6340 2140 6420
rect 2260 6340 2340 6420
rect 2460 6340 2540 6420
rect 2660 6340 2740 6420
rect 2860 6340 2940 6420
rect 3060 6340 3140 6420
rect 3260 6340 3340 6420
rect 3460 6340 3540 6420
rect 3660 6340 3740 6420
rect 3860 6340 3940 6420
rect 4060 6340 4140 6420
rect 4260 6340 4340 6420
rect 4460 6340 4540 6420
rect 4660 6340 4740 6420
rect 4860 6340 4940 6420
rect 5060 6340 5140 6420
rect 5260 6340 5340 6420
rect 5460 6340 5540 6420
rect 5660 6340 5740 6420
rect 5860 6340 5940 6420
rect 6060 6340 6140 6420
rect 6260 6340 6340 6420
rect 6460 6340 6540 6420
rect -140 6155 -60 6235
rect 60 6155 140 6235
rect 260 6155 340 6235
rect 460 6155 540 6235
rect 660 6155 740 6235
rect 860 6155 940 6235
rect 1060 6155 1140 6235
rect 1260 6155 1340 6235
rect 1460 6155 1540 6235
rect 1660 6155 1740 6235
rect 1860 6155 1940 6235
rect 2060 6155 2140 6235
rect 2260 6155 2340 6235
rect 2460 6155 2540 6235
rect 2660 6155 2740 6235
rect 2860 6155 2940 6235
rect 3060 6155 3140 6235
rect 3260 6155 3340 6235
rect 3460 6155 3540 6235
rect 3660 6155 3740 6235
rect 3860 6155 3940 6235
rect 4060 6155 4140 6235
rect 4260 6155 4340 6235
rect 4460 6155 4540 6235
rect 4660 6155 4740 6235
rect 4860 6155 4940 6235
rect 5060 6155 5140 6235
rect 5260 6155 5340 6235
rect 5460 6155 5540 6235
rect 5660 6155 5740 6235
rect 5860 6155 5940 6235
rect 6060 6155 6140 6235
rect 6260 6155 6340 6235
rect 6460 6155 6540 6235
rect -140 5970 -60 6050
rect 60 5970 140 6050
rect 260 5970 340 6050
rect 460 5970 540 6050
rect 660 5970 740 6050
rect 860 5970 940 6050
rect 1060 5970 1140 6050
rect 1260 5970 1340 6050
rect 1460 5970 1540 6050
rect 1660 5970 1740 6050
rect 1860 5970 1940 6050
rect 2060 5970 2140 6050
rect 2260 5970 2340 6050
rect 2460 5970 2540 6050
rect 2660 5970 2740 6050
rect 2860 5970 2940 6050
rect 3060 5970 3140 6050
rect 3260 5970 3340 6050
rect 3460 5970 3540 6050
rect 3660 5970 3740 6050
rect 3860 5970 3940 6050
rect 4060 5970 4140 6050
rect 4260 5970 4340 6050
rect 4460 5970 4540 6050
rect 4660 5970 4740 6050
rect 4860 5970 4940 6050
rect 5060 5970 5140 6050
rect 5260 5970 5340 6050
rect 5460 5970 5540 6050
rect 5660 5970 5740 6050
rect 5860 5970 5940 6050
rect 6060 5970 6140 6050
rect 6260 5970 6340 6050
rect 6460 5970 6540 6050
rect -140 5785 -60 5865
rect 60 5785 140 5865
rect 260 5785 340 5865
rect 460 5785 540 5865
rect 660 5785 740 5865
rect 860 5785 940 5865
rect 1060 5785 1140 5865
rect 1260 5785 1340 5865
rect 1460 5785 1540 5865
rect 1660 5785 1740 5865
rect 1860 5785 1940 5865
rect 2060 5785 2140 5865
rect 2260 5785 2340 5865
rect 2460 5785 2540 5865
rect 2660 5785 2740 5865
rect 2860 5785 2940 5865
rect 3060 5785 3140 5865
rect 3260 5785 3340 5865
rect 3460 5785 3540 5865
rect 3660 5785 3740 5865
rect 3860 5785 3940 5865
rect 4060 5785 4140 5865
rect 4260 5785 4340 5865
rect 4460 5785 4540 5865
rect 4660 5785 4740 5865
rect 4860 5785 4940 5865
rect 5060 5785 5140 5865
rect 5260 5785 5340 5865
rect 5460 5785 5540 5865
rect 5660 5785 5740 5865
rect 5860 5785 5940 5865
rect 6060 5785 6140 5865
rect 6260 5785 6340 5865
rect 6460 5785 6540 5865
rect -140 5600 -60 5680
rect 60 5600 140 5680
rect 260 5600 340 5680
rect 460 5600 540 5680
rect 660 5600 740 5680
rect 860 5600 940 5680
rect 1060 5600 1140 5680
rect 1260 5600 1340 5680
rect 1460 5600 1540 5680
rect 1660 5600 1740 5680
rect 1860 5600 1940 5680
rect 2060 5600 2140 5680
rect 2260 5600 2340 5680
rect 2460 5600 2540 5680
rect 2660 5600 2740 5680
rect 2860 5600 2940 5680
rect 3060 5600 3140 5680
rect 3260 5600 3340 5680
rect 3460 5600 3540 5680
rect 3660 5600 3740 5680
rect 3860 5600 3940 5680
rect 4060 5600 4140 5680
rect 4260 5600 4340 5680
rect 4460 5600 4540 5680
rect 4660 5600 4740 5680
rect 4860 5600 4940 5680
rect 5060 5600 5140 5680
rect 5260 5600 5340 5680
rect 5460 5600 5540 5680
rect 5660 5600 5740 5680
rect 5860 5600 5940 5680
rect 6060 5600 6140 5680
rect 6260 5600 6340 5680
rect 6460 5600 6540 5680
rect -140 5415 -60 5495
rect 60 5415 140 5495
rect 260 5415 340 5495
rect 460 5415 540 5495
rect 660 5415 740 5495
rect 860 5415 940 5495
rect 1060 5415 1140 5495
rect 1260 5415 1340 5495
rect 1460 5415 1540 5495
rect 1660 5415 1740 5495
rect 1860 5415 1940 5495
rect 2060 5415 2140 5495
rect 2260 5415 2340 5495
rect 2460 5415 2540 5495
rect 2660 5415 2740 5495
rect 2860 5415 2940 5495
rect 3060 5415 3140 5495
rect 3260 5415 3340 5495
rect 3460 5415 3540 5495
rect 3660 5415 3740 5495
rect 3860 5415 3940 5495
rect 4060 5415 4140 5495
rect 4260 5415 4340 5495
rect 4460 5415 4540 5495
rect 4660 5415 4740 5495
rect 4860 5415 4940 5495
rect 5060 5415 5140 5495
rect 5260 5415 5340 5495
rect 5460 5415 5540 5495
rect 5660 5415 5740 5495
rect 5860 5415 5940 5495
rect 6060 5415 6140 5495
rect 6260 5415 6340 5495
rect 6460 5415 6540 5495
rect -140 5230 -60 5310
rect 60 5230 140 5310
rect 260 5230 340 5310
rect 460 5230 540 5310
rect 660 5230 740 5310
rect 860 5230 940 5310
rect 1060 5230 1140 5310
rect 1260 5230 1340 5310
rect 1460 5230 1540 5310
rect 1660 5230 1740 5310
rect 1860 5230 1940 5310
rect 2060 5230 2140 5310
rect 2260 5230 2340 5310
rect 2460 5230 2540 5310
rect 2660 5230 2740 5310
rect 2860 5230 2940 5310
rect 3060 5230 3140 5310
rect 3260 5230 3340 5310
rect 3460 5230 3540 5310
rect 3660 5230 3740 5310
rect 3860 5230 3940 5310
rect 4060 5230 4140 5310
rect 4260 5230 4340 5310
rect 4460 5230 4540 5310
rect 4660 5230 4740 5310
rect 4860 5230 4940 5310
rect 5060 5230 5140 5310
rect 5260 5230 5340 5310
rect 5460 5230 5540 5310
rect 5660 5230 5740 5310
rect 5860 5230 5940 5310
rect 6060 5230 6140 5310
rect 6260 5230 6340 5310
rect 6460 5230 6540 5310
rect -140 5045 -60 5125
rect 60 5045 140 5125
rect 260 5045 340 5125
rect 460 5045 540 5125
rect 660 5045 740 5125
rect 860 5045 940 5125
rect 1060 5045 1140 5125
rect 1260 5045 1340 5125
rect 1460 5045 1540 5125
rect 1660 5045 1740 5125
rect 1860 5045 1940 5125
rect 2060 5045 2140 5125
rect 2260 5045 2340 5125
rect 2460 5045 2540 5125
rect 2660 5045 2740 5125
rect 2860 5045 2940 5125
rect 3060 5045 3140 5125
rect 3260 5045 3340 5125
rect 3460 5045 3540 5125
rect 3660 5045 3740 5125
rect 3860 5045 3940 5125
rect 4060 5045 4140 5125
rect 4260 5045 4340 5125
rect 4460 5045 4540 5125
rect 4660 5045 4740 5125
rect 4860 5045 4940 5125
rect 5060 5045 5140 5125
rect 5260 5045 5340 5125
rect 5460 5045 5540 5125
rect 5660 5045 5740 5125
rect 5860 5045 5940 5125
rect 6060 5045 6140 5125
rect 6260 5045 6340 5125
rect 6460 5045 6540 5125
rect -140 4860 -60 4940
rect 60 4860 140 4940
rect 260 4860 340 4940
rect 460 4860 540 4940
rect 660 4860 740 4940
rect 860 4860 940 4940
rect 1060 4860 1140 4940
rect 1260 4860 1340 4940
rect 1460 4860 1540 4940
rect 1660 4860 1740 4940
rect 1860 4860 1940 4940
rect 2060 4860 2140 4940
rect 2260 4860 2340 4940
rect 2460 4860 2540 4940
rect 2660 4860 2740 4940
rect 2860 4860 2940 4940
rect 3060 4860 3140 4940
rect 3260 4860 3340 4940
rect 3460 4860 3540 4940
rect 3660 4860 3740 4940
rect 3860 4860 3940 4940
rect 4060 4860 4140 4940
rect 4260 4860 4340 4940
rect 4460 4860 4540 4940
rect 4660 4860 4740 4940
rect 4860 4860 4940 4940
rect 5060 4860 5140 4940
rect 5260 4860 5340 4940
rect 5460 4860 5540 4940
rect 5660 4860 5740 4940
rect 5860 4860 5940 4940
rect 6060 4860 6140 4940
rect 6260 4860 6340 4940
rect 6460 4860 6540 4940
rect -140 4675 -60 4755
rect 60 4675 140 4755
rect 260 4675 340 4755
rect 460 4675 540 4755
rect 660 4675 740 4755
rect 860 4675 940 4755
rect 1060 4675 1140 4755
rect 1260 4675 1340 4755
rect 1460 4675 1540 4755
rect 1660 4675 1740 4755
rect 1860 4675 1940 4755
rect 2060 4675 2140 4755
rect 2260 4675 2340 4755
rect 2460 4675 2540 4755
rect 2660 4675 2740 4755
rect 2860 4675 2940 4755
rect 3060 4675 3140 4755
rect 3260 4675 3340 4755
rect 3460 4675 3540 4755
rect 3660 4675 3740 4755
rect 3860 4675 3940 4755
rect 4060 4675 4140 4755
rect 4260 4675 4340 4755
rect 4460 4675 4540 4755
rect 4660 4675 4740 4755
rect 4860 4675 4940 4755
rect 5060 4675 5140 4755
rect 5260 4675 5340 4755
rect 5460 4675 5540 4755
rect 5660 4675 5740 4755
rect 5860 4675 5940 4755
rect 6060 4675 6140 4755
rect 6260 4675 6340 4755
rect 6460 4675 6540 4755
rect -140 4490 -60 4570
rect 60 4490 140 4570
rect 260 4490 340 4570
rect 460 4490 540 4570
rect 660 4490 740 4570
rect 860 4490 940 4570
rect 1060 4490 1140 4570
rect 1260 4490 1340 4570
rect 1460 4490 1540 4570
rect 1660 4490 1740 4570
rect 1860 4490 1940 4570
rect 2060 4490 2140 4570
rect 2260 4490 2340 4570
rect 2460 4490 2540 4570
rect 2660 4490 2740 4570
rect 2860 4490 2940 4570
rect 3060 4490 3140 4570
rect 3260 4490 3340 4570
rect 3460 4490 3540 4570
rect 3660 4490 3740 4570
rect 3860 4490 3940 4570
rect 4060 4490 4140 4570
rect 4260 4490 4340 4570
rect 4460 4490 4540 4570
rect 4660 4490 4740 4570
rect 4860 4490 4940 4570
rect 5060 4490 5140 4570
rect 5260 4490 5340 4570
rect 5460 4490 5540 4570
rect 5660 4490 5740 4570
rect 5860 4490 5940 4570
rect 6060 4490 6140 4570
rect 6260 4490 6340 4570
rect 6460 4490 6540 4570
rect -140 4305 -60 4385
rect 60 4305 140 4385
rect 260 4305 340 4385
rect 460 4305 540 4385
rect 660 4305 740 4385
rect 860 4305 940 4385
rect 1060 4305 1140 4385
rect 1260 4305 1340 4385
rect 1460 4305 1540 4385
rect 1660 4305 1740 4385
rect 1860 4305 1940 4385
rect 2060 4305 2140 4385
rect 2260 4305 2340 4385
rect 2460 4305 2540 4385
rect 2660 4305 2740 4385
rect 2860 4305 2940 4385
rect 3060 4305 3140 4385
rect 3260 4305 3340 4385
rect 3460 4305 3540 4385
rect 3660 4305 3740 4385
rect 3860 4305 3940 4385
rect 4060 4305 4140 4385
rect 4260 4305 4340 4385
rect 4460 4305 4540 4385
rect 4660 4305 4740 4385
rect 4860 4305 4940 4385
rect 5060 4305 5140 4385
rect 5260 4305 5340 4385
rect 5460 4305 5540 4385
rect 5660 4305 5740 4385
rect 5860 4305 5940 4385
rect 6060 4305 6140 4385
rect 6260 4305 6340 4385
rect 6460 4305 6540 4385
rect -140 4120 -60 4200
rect 60 4120 140 4200
rect 260 4120 340 4200
rect 460 4120 540 4200
rect 660 4120 740 4200
rect 860 4120 940 4200
rect 1060 4120 1140 4200
rect 1260 4120 1340 4200
rect 1460 4120 1540 4200
rect 1660 4120 1740 4200
rect 1860 4120 1940 4200
rect 2060 4120 2140 4200
rect 2260 4120 2340 4200
rect 2460 4120 2540 4200
rect 2660 4120 2740 4200
rect 2860 4120 2940 4200
rect 3060 4120 3140 4200
rect 3260 4120 3340 4200
rect 3460 4120 3540 4200
rect 3660 4120 3740 4200
rect 3860 4120 3940 4200
rect 4060 4120 4140 4200
rect 4260 4120 4340 4200
rect 4460 4120 4540 4200
rect 4660 4120 4740 4200
rect 4860 4120 4940 4200
rect 5060 4120 5140 4200
rect 5260 4120 5340 4200
rect 5460 4120 5540 4200
rect 5660 4120 5740 4200
rect 5860 4120 5940 4200
rect 6060 4120 6140 4200
rect 6260 4120 6340 4200
rect 6460 4120 6540 4200
rect -140 3935 -60 4015
rect 60 3935 140 4015
rect 260 3935 340 4015
rect 460 3935 540 4015
rect 660 3935 740 4015
rect 860 3935 940 4015
rect 1060 3935 1140 4015
rect 1260 3935 1340 4015
rect 1460 3935 1540 4015
rect 1660 3935 1740 4015
rect 1860 3935 1940 4015
rect 2060 3935 2140 4015
rect 2260 3935 2340 4015
rect 2460 3935 2540 4015
rect 2660 3935 2740 4015
rect 2860 3935 2940 4015
rect 3060 3935 3140 4015
rect 3260 3935 3340 4015
rect 3460 3935 3540 4015
rect 3660 3935 3740 4015
rect 3860 3935 3940 4015
rect 4060 3935 4140 4015
rect 4260 3935 4340 4015
rect 4460 3935 4540 4015
rect 4660 3935 4740 4015
rect 4860 3935 4940 4015
rect 5060 3935 5140 4015
rect 5260 3935 5340 4015
rect 5460 3935 5540 4015
rect 5660 3935 5740 4015
rect 5860 3935 5940 4015
rect 6060 3935 6140 4015
rect 6260 3935 6340 4015
rect 6460 3935 6540 4015
rect -140 3750 -60 3830
rect 60 3750 140 3830
rect 260 3750 340 3830
rect 460 3750 540 3830
rect 660 3750 740 3830
rect 860 3750 940 3830
rect 1060 3750 1140 3830
rect 1260 3750 1340 3830
rect 1460 3750 1540 3830
rect 1660 3750 1740 3830
rect 1860 3750 1940 3830
rect 2060 3750 2140 3830
rect 2260 3750 2340 3830
rect 2460 3750 2540 3830
rect 2660 3750 2740 3830
rect 2860 3750 2940 3830
rect 3060 3750 3140 3830
rect 3260 3750 3340 3830
rect 3460 3750 3540 3830
rect 3660 3750 3740 3830
rect 3860 3750 3940 3830
rect 4060 3750 4140 3830
rect 4260 3750 4340 3830
rect 4460 3750 4540 3830
rect 4660 3750 4740 3830
rect 4860 3750 4940 3830
rect 5060 3750 5140 3830
rect 5260 3750 5340 3830
rect 5460 3750 5540 3830
rect 5660 3750 5740 3830
rect 5860 3750 5940 3830
rect 6060 3750 6140 3830
rect 6260 3750 6340 3830
rect 6460 3750 6540 3830
rect -140 3565 -60 3645
rect 60 3565 140 3645
rect 260 3565 340 3645
rect 460 3565 540 3645
rect 660 3565 740 3645
rect 860 3565 940 3645
rect 1060 3565 1140 3645
rect 1260 3565 1340 3645
rect 1460 3565 1540 3645
rect 1660 3565 1740 3645
rect 1860 3565 1940 3645
rect 2060 3565 2140 3645
rect 2260 3565 2340 3645
rect 2460 3565 2540 3645
rect 2660 3565 2740 3645
rect 2860 3565 2940 3645
rect 3060 3565 3140 3645
rect 3260 3565 3340 3645
rect 3460 3565 3540 3645
rect 3660 3565 3740 3645
rect 3860 3565 3940 3645
rect 4060 3565 4140 3645
rect 4260 3565 4340 3645
rect 4460 3565 4540 3645
rect 4660 3565 4740 3645
rect 4860 3565 4940 3645
rect 5060 3565 5140 3645
rect 5260 3565 5340 3645
rect 5460 3565 5540 3645
rect 5660 3565 5740 3645
rect 5860 3565 5940 3645
rect 6060 3565 6140 3645
rect 6260 3565 6340 3645
rect 6460 3565 6540 3645
rect -140 3380 -60 3460
rect 60 3380 140 3460
rect 260 3380 340 3460
rect 460 3380 540 3460
rect 660 3380 740 3460
rect 860 3380 940 3460
rect 1060 3380 1140 3460
rect 1260 3380 1340 3460
rect 1460 3380 1540 3460
rect 1660 3380 1740 3460
rect 1860 3380 1940 3460
rect 2060 3380 2140 3460
rect 2260 3380 2340 3460
rect 2460 3380 2540 3460
rect 2660 3380 2740 3460
rect 2860 3380 2940 3460
rect 3060 3380 3140 3460
rect 3260 3380 3340 3460
rect 3460 3380 3540 3460
rect 3660 3380 3740 3460
rect 3860 3380 3940 3460
rect 4060 3380 4140 3460
rect 4260 3380 4340 3460
rect 4460 3380 4540 3460
rect 4660 3380 4740 3460
rect 4860 3380 4940 3460
rect 5060 3380 5140 3460
rect 5260 3380 5340 3460
rect 5460 3380 5540 3460
rect 5660 3380 5740 3460
rect 5860 3380 5940 3460
rect 6060 3380 6140 3460
rect 6260 3380 6340 3460
rect 6460 3380 6540 3460
rect -140 3195 -60 3275
rect 60 3195 140 3275
rect 260 3195 340 3275
rect 460 3195 540 3275
rect 660 3195 740 3275
rect 860 3195 940 3275
rect 1060 3195 1140 3275
rect 1260 3195 1340 3275
rect 1460 3195 1540 3275
rect 1660 3195 1740 3275
rect 1860 3195 1940 3275
rect 2060 3195 2140 3275
rect 2260 3195 2340 3275
rect 2460 3195 2540 3275
rect 2660 3195 2740 3275
rect 2860 3195 2940 3275
rect 3060 3195 3140 3275
rect 3260 3195 3340 3275
rect 3460 3195 3540 3275
rect 3660 3195 3740 3275
rect 3860 3195 3940 3275
rect 4060 3195 4140 3275
rect 4260 3195 4340 3275
rect 4460 3195 4540 3275
rect 4660 3195 4740 3275
rect 4860 3195 4940 3275
rect 5060 3195 5140 3275
rect 5260 3195 5340 3275
rect 5460 3195 5540 3275
rect 5660 3195 5740 3275
rect 5860 3195 5940 3275
rect 6060 3195 6140 3275
rect 6260 3195 6340 3275
rect 6460 3195 6540 3275
rect -140 3010 -60 3090
rect 60 3010 140 3090
rect 260 3010 340 3090
rect 460 3010 540 3090
rect 660 3010 740 3090
rect 860 3010 940 3090
rect 1060 3010 1140 3090
rect 1260 3010 1340 3090
rect 1460 3010 1540 3090
rect 1660 3010 1740 3090
rect 1860 3010 1940 3090
rect 2060 3010 2140 3090
rect 2260 3010 2340 3090
rect 2460 3010 2540 3090
rect 2660 3010 2740 3090
rect 2860 3010 2940 3090
rect 3060 3010 3140 3090
rect 3260 3010 3340 3090
rect 3460 3010 3540 3090
rect 3660 3010 3740 3090
rect 3860 3010 3940 3090
rect 4060 3010 4140 3090
rect 4260 3010 4340 3090
rect 4460 3010 4540 3090
rect 4660 3010 4740 3090
rect 4860 3010 4940 3090
rect 5060 3010 5140 3090
rect 5260 3010 5340 3090
rect 5460 3010 5540 3090
rect 5660 3010 5740 3090
rect 5860 3010 5940 3090
rect 6060 3010 6140 3090
rect 6260 3010 6340 3090
rect 6460 3010 6540 3090
rect -140 2825 -60 2905
rect 60 2825 140 2905
rect 260 2825 340 2905
rect 460 2825 540 2905
rect 660 2825 740 2905
rect 860 2825 940 2905
rect 1060 2825 1140 2905
rect 1260 2825 1340 2905
rect 1460 2825 1540 2905
rect 1660 2825 1740 2905
rect 1860 2825 1940 2905
rect 2060 2825 2140 2905
rect 2260 2825 2340 2905
rect 2460 2825 2540 2905
rect 2660 2825 2740 2905
rect 2860 2825 2940 2905
rect 3060 2825 3140 2905
rect 3260 2825 3340 2905
rect 3460 2825 3540 2905
rect 3660 2825 3740 2905
rect 3860 2825 3940 2905
rect 4060 2825 4140 2905
rect 4260 2825 4340 2905
rect 4460 2825 4540 2905
rect 4660 2825 4740 2905
rect 4860 2825 4940 2905
rect 5060 2825 5140 2905
rect 5260 2825 5340 2905
rect 5460 2825 5540 2905
rect 5660 2825 5740 2905
rect 5860 2825 5940 2905
rect 6060 2825 6140 2905
rect 6260 2825 6340 2905
rect 6460 2825 6540 2905
rect -140 2640 -60 2720
rect 60 2640 140 2720
rect 260 2640 340 2720
rect 460 2640 540 2720
rect 660 2640 740 2720
rect 860 2640 940 2720
rect 1060 2640 1140 2720
rect 1260 2640 1340 2720
rect 1460 2640 1540 2720
rect 1660 2640 1740 2720
rect 1860 2640 1940 2720
rect 2060 2640 2140 2720
rect 2260 2640 2340 2720
rect 2460 2640 2540 2720
rect 2660 2640 2740 2720
rect 2860 2640 2940 2720
rect 3060 2640 3140 2720
rect 3260 2640 3340 2720
rect 3460 2640 3540 2720
rect 3660 2640 3740 2720
rect 3860 2640 3940 2720
rect 4060 2640 4140 2720
rect 4260 2640 4340 2720
rect 4460 2640 4540 2720
rect 4660 2640 4740 2720
rect 4860 2640 4940 2720
rect 5060 2640 5140 2720
rect 5260 2640 5340 2720
rect 5460 2640 5540 2720
rect 5660 2640 5740 2720
rect 5860 2640 5940 2720
rect 6060 2640 6140 2720
rect 6260 2640 6340 2720
rect 6460 2640 6540 2720
rect -140 2455 -60 2535
rect 60 2455 140 2535
rect 260 2455 340 2535
rect 460 2455 540 2535
rect 660 2455 740 2535
rect 860 2455 940 2535
rect 1060 2455 1140 2535
rect 1260 2455 1340 2535
rect 1460 2455 1540 2535
rect 1660 2455 1740 2535
rect 1860 2455 1940 2535
rect 2060 2455 2140 2535
rect 2260 2455 2340 2535
rect 2460 2455 2540 2535
rect 2660 2455 2740 2535
rect 2860 2455 2940 2535
rect 3060 2455 3140 2535
rect 3260 2455 3340 2535
rect 3460 2455 3540 2535
rect 3660 2455 3740 2535
rect 3860 2455 3940 2535
rect 4060 2455 4140 2535
rect 4260 2455 4340 2535
rect 4460 2455 4540 2535
rect 4660 2455 4740 2535
rect 4860 2455 4940 2535
rect 5060 2455 5140 2535
rect 5260 2455 5340 2535
rect 5460 2455 5540 2535
rect 5660 2455 5740 2535
rect 5860 2455 5940 2535
rect 6060 2455 6140 2535
rect 6260 2455 6340 2535
rect 6460 2455 6540 2535
rect -140 2270 -60 2350
rect 60 2270 140 2350
rect 260 2270 340 2350
rect 460 2270 540 2350
rect 660 2270 740 2350
rect 860 2270 940 2350
rect 1060 2270 1140 2350
rect 1260 2270 1340 2350
rect 1460 2270 1540 2350
rect 1660 2270 1740 2350
rect 1860 2270 1940 2350
rect 2060 2270 2140 2350
rect 2260 2270 2340 2350
rect 2460 2270 2540 2350
rect 2660 2270 2740 2350
rect 2860 2270 2940 2350
rect 3060 2270 3140 2350
rect 3260 2270 3340 2350
rect 3460 2270 3540 2350
rect 3660 2270 3740 2350
rect 3860 2270 3940 2350
rect 4060 2270 4140 2350
rect 4260 2270 4340 2350
rect 4460 2270 4540 2350
rect 4660 2270 4740 2350
rect 4860 2270 4940 2350
rect 5060 2270 5140 2350
rect 5260 2270 5340 2350
rect 5460 2270 5540 2350
rect 5660 2270 5740 2350
rect 5860 2270 5940 2350
rect 6060 2270 6140 2350
rect 6260 2270 6340 2350
rect 6460 2270 6540 2350
rect -140 2085 -60 2165
rect 60 2085 140 2165
rect 260 2085 340 2165
rect 460 2085 540 2165
rect 660 2085 740 2165
rect 860 2085 940 2165
rect 1060 2085 1140 2165
rect 1260 2085 1340 2165
rect 1460 2085 1540 2165
rect 1660 2085 1740 2165
rect 1860 2085 1940 2165
rect 2060 2085 2140 2165
rect 2260 2085 2340 2165
rect 2460 2085 2540 2165
rect 2660 2085 2740 2165
rect 2860 2085 2940 2165
rect 3060 2085 3140 2165
rect 3260 2085 3340 2165
rect 3460 2085 3540 2165
rect 3660 2085 3740 2165
rect 3860 2085 3940 2165
rect 4060 2085 4140 2165
rect 4260 2085 4340 2165
rect 4460 2085 4540 2165
rect 4660 2085 4740 2165
rect 4860 2085 4940 2165
rect 5060 2085 5140 2165
rect 5260 2085 5340 2165
rect 5460 2085 5540 2165
rect 5660 2085 5740 2165
rect 5860 2085 5940 2165
rect 6060 2085 6140 2165
rect 6260 2085 6340 2165
rect 6460 2085 6540 2165
rect -140 1900 -60 1980
rect 60 1900 140 1980
rect 260 1900 340 1980
rect 460 1900 540 1980
rect 660 1900 740 1980
rect 860 1900 940 1980
rect 1060 1900 1140 1980
rect 1260 1900 1340 1980
rect 1460 1900 1540 1980
rect 1660 1900 1740 1980
rect 1860 1900 1940 1980
rect 2060 1900 2140 1980
rect 2260 1900 2340 1980
rect 2460 1900 2540 1980
rect 2660 1900 2740 1980
rect 2860 1900 2940 1980
rect 3060 1900 3140 1980
rect 3260 1900 3340 1980
rect 3460 1900 3540 1980
rect 3660 1900 3740 1980
rect 3860 1900 3940 1980
rect 4060 1900 4140 1980
rect 4260 1900 4340 1980
rect 4460 1900 4540 1980
rect 4660 1900 4740 1980
rect 4860 1900 4940 1980
rect 5060 1900 5140 1980
rect 5260 1900 5340 1980
rect 5460 1900 5540 1980
rect 5660 1900 5740 1980
rect 5860 1900 5940 1980
rect 6060 1900 6140 1980
rect 6260 1900 6340 1980
rect 6460 1900 6540 1980
rect -140 1715 -60 1795
rect 60 1715 140 1795
rect 260 1715 340 1795
rect 460 1715 540 1795
rect 660 1715 740 1795
rect 860 1715 940 1795
rect 1060 1715 1140 1795
rect 1260 1715 1340 1795
rect 1460 1715 1540 1795
rect 1660 1715 1740 1795
rect 1860 1715 1940 1795
rect 2060 1715 2140 1795
rect 2260 1715 2340 1795
rect 2460 1715 2540 1795
rect 2660 1715 2740 1795
rect 2860 1715 2940 1795
rect 3060 1715 3140 1795
rect 3260 1715 3340 1795
rect 3460 1715 3540 1795
rect 3660 1715 3740 1795
rect 3860 1715 3940 1795
rect 4060 1715 4140 1795
rect 4260 1715 4340 1795
rect 4460 1715 4540 1795
rect 4660 1715 4740 1795
rect 4860 1715 4940 1795
rect 5060 1715 5140 1795
rect 5260 1715 5340 1795
rect 5460 1715 5540 1795
rect 5660 1715 5740 1795
rect 5860 1715 5940 1795
rect 6060 1715 6140 1795
rect 6260 1715 6340 1795
rect 6460 1715 6540 1795
rect -140 1530 -60 1610
rect 60 1530 140 1610
rect 260 1530 340 1610
rect 460 1530 540 1610
rect 660 1530 740 1610
rect 860 1530 940 1610
rect 1060 1530 1140 1610
rect 1260 1530 1340 1610
rect 1460 1530 1540 1610
rect 1660 1530 1740 1610
rect 1860 1530 1940 1610
rect 2060 1530 2140 1610
rect 2260 1530 2340 1610
rect 2460 1530 2540 1610
rect 2660 1530 2740 1610
rect 2860 1530 2940 1610
rect 3060 1530 3140 1610
rect 3260 1530 3340 1610
rect 3460 1530 3540 1610
rect 3660 1530 3740 1610
rect 3860 1530 3940 1610
rect 4060 1530 4140 1610
rect 4260 1530 4340 1610
rect 4460 1530 4540 1610
rect 4660 1530 4740 1610
rect 4860 1530 4940 1610
rect 5060 1530 5140 1610
rect 5260 1530 5340 1610
rect 5460 1530 5540 1610
rect 5660 1530 5740 1610
rect 5860 1530 5940 1610
rect 6060 1530 6140 1610
rect 6260 1530 6340 1610
rect 6460 1530 6540 1610
rect -140 1345 -60 1425
rect 60 1345 140 1425
rect 260 1345 340 1425
rect 460 1345 540 1425
rect 660 1345 740 1425
rect 860 1345 940 1425
rect 1060 1345 1140 1425
rect 1260 1345 1340 1425
rect 1460 1345 1540 1425
rect 1660 1345 1740 1425
rect 1860 1345 1940 1425
rect 2060 1345 2140 1425
rect 2260 1345 2340 1425
rect 2460 1345 2540 1425
rect 2660 1345 2740 1425
rect 2860 1345 2940 1425
rect 3060 1345 3140 1425
rect 3260 1345 3340 1425
rect 3460 1345 3540 1425
rect 3660 1345 3740 1425
rect 3860 1345 3940 1425
rect 4060 1345 4140 1425
rect 4260 1345 4340 1425
rect 4460 1345 4540 1425
rect 4660 1345 4740 1425
rect 4860 1345 4940 1425
rect 5060 1345 5140 1425
rect 5260 1345 5340 1425
rect 5460 1345 5540 1425
rect 5660 1345 5740 1425
rect 5860 1345 5940 1425
rect 6060 1345 6140 1425
rect 6260 1345 6340 1425
rect 6460 1345 6540 1425
rect -140 1160 -60 1240
rect 60 1160 140 1240
rect 260 1160 340 1240
rect 460 1160 540 1240
rect 660 1160 740 1240
rect 860 1160 940 1240
rect 1060 1160 1140 1240
rect 1260 1160 1340 1240
rect 1460 1160 1540 1240
rect 1660 1160 1740 1240
rect 1860 1160 1940 1240
rect 2060 1160 2140 1240
rect 2260 1160 2340 1240
rect 2460 1160 2540 1240
rect 2660 1160 2740 1240
rect 2860 1160 2940 1240
rect 3060 1160 3140 1240
rect 3260 1160 3340 1240
rect 3460 1160 3540 1240
rect 3660 1160 3740 1240
rect 3860 1160 3940 1240
rect 4060 1160 4140 1240
rect 4260 1160 4340 1240
rect 4460 1160 4540 1240
rect 4660 1160 4740 1240
rect 4860 1160 4940 1240
rect 5060 1160 5140 1240
rect 5260 1160 5340 1240
rect 5460 1160 5540 1240
rect 5660 1160 5740 1240
rect 5860 1160 5940 1240
rect 6060 1160 6140 1240
rect 6260 1160 6340 1240
rect 6460 1160 6540 1240
rect -140 975 -60 1055
rect 60 975 140 1055
rect 260 975 340 1055
rect 460 975 540 1055
rect 660 975 740 1055
rect 860 975 940 1055
rect 1060 975 1140 1055
rect 1260 975 1340 1055
rect 1460 975 1540 1055
rect 1660 975 1740 1055
rect 1860 975 1940 1055
rect 2060 975 2140 1055
rect 2260 975 2340 1055
rect 2460 975 2540 1055
rect 2660 975 2740 1055
rect 2860 975 2940 1055
rect 3060 975 3140 1055
rect 3260 975 3340 1055
rect 3460 975 3540 1055
rect 3660 975 3740 1055
rect 3860 975 3940 1055
rect 4060 975 4140 1055
rect 4260 975 4340 1055
rect 4460 975 4540 1055
rect 4660 975 4740 1055
rect 4860 975 4940 1055
rect 5060 975 5140 1055
rect 5260 975 5340 1055
rect 5460 975 5540 1055
rect 5660 975 5740 1055
rect 5860 975 5940 1055
rect 6060 975 6140 1055
rect 6260 975 6340 1055
rect 6460 975 6540 1055
rect -140 790 -60 870
rect 60 790 140 870
rect 260 790 340 870
rect 460 790 540 870
rect 660 790 740 870
rect 860 790 940 870
rect 1060 790 1140 870
rect 1260 790 1340 870
rect 1460 790 1540 870
rect 1660 790 1740 870
rect 1860 790 1940 870
rect 2060 790 2140 870
rect 2260 790 2340 870
rect 2460 790 2540 870
rect 2660 790 2740 870
rect 2860 790 2940 870
rect 3060 790 3140 870
rect 3260 790 3340 870
rect 3460 790 3540 870
rect 3660 790 3740 870
rect 3860 790 3940 870
rect 4060 790 4140 870
rect 4260 790 4340 870
rect 4460 790 4540 870
rect 4660 790 4740 870
rect 4860 790 4940 870
rect 5060 790 5140 870
rect 5260 790 5340 870
rect 5460 790 5540 870
rect 5660 790 5740 870
rect 5860 790 5940 870
rect 6060 790 6140 870
rect 6260 790 6340 870
rect 6460 790 6540 870
rect -140 605 -60 685
rect 60 605 140 685
rect 260 605 340 685
rect 460 605 540 685
rect 660 605 740 685
rect 860 605 940 685
rect 1060 605 1140 685
rect 1260 605 1340 685
rect 1460 605 1540 685
rect 1660 605 1740 685
rect 1860 605 1940 685
rect 2060 605 2140 685
rect 2260 605 2340 685
rect 2460 605 2540 685
rect 2660 605 2740 685
rect 2860 605 2940 685
rect 3060 605 3140 685
rect 3260 605 3340 685
rect 3460 605 3540 685
rect 3660 605 3740 685
rect 3860 605 3940 685
rect 4060 605 4140 685
rect 4260 605 4340 685
rect 4460 605 4540 685
rect 4660 605 4740 685
rect 4860 605 4940 685
rect 5060 605 5140 685
rect 5260 605 5340 685
rect 5460 605 5540 685
rect 5660 605 5740 685
rect 5860 605 5940 685
rect 6060 605 6140 685
rect 6260 605 6340 685
rect 6460 605 6540 685
rect -140 420 -60 500
rect 60 420 140 500
rect 260 420 340 500
rect 460 420 540 500
rect 660 420 740 500
rect 860 420 940 500
rect 1060 420 1140 500
rect 1260 420 1340 500
rect 1460 420 1540 500
rect 1660 420 1740 500
rect 1860 420 1940 500
rect 2060 420 2140 500
rect 2260 420 2340 500
rect 2460 420 2540 500
rect 2660 420 2740 500
rect 2860 420 2940 500
rect 3060 420 3140 500
rect 3260 420 3340 500
rect 3460 420 3540 500
rect 3660 420 3740 500
rect 3860 420 3940 500
rect 4060 420 4140 500
rect 4260 420 4340 500
rect 4460 420 4540 500
rect 4660 420 4740 500
rect 4860 420 4940 500
rect 5060 420 5140 500
rect 5260 420 5340 500
rect 5460 420 5540 500
rect 5660 420 5740 500
rect 5860 420 5940 500
rect 6060 420 6140 500
rect 6260 420 6340 500
rect 6460 420 6540 500
rect -140 235 -60 315
rect 60 235 140 315
rect 260 235 340 315
rect 460 235 540 315
rect 660 235 740 315
rect 860 235 940 315
rect 1060 235 1140 315
rect 1260 235 1340 315
rect 1460 235 1540 315
rect 1660 235 1740 315
rect 1860 235 1940 315
rect 2060 235 2140 315
rect 2260 235 2340 315
rect 2460 235 2540 315
rect 2660 235 2740 315
rect 2860 235 2940 315
rect 3060 235 3140 315
rect 3260 235 3340 315
rect 3460 235 3540 315
rect 3660 235 3740 315
rect 3860 235 3940 315
rect 4060 235 4140 315
rect 4260 235 4340 315
rect 4460 235 4540 315
rect 4660 235 4740 315
rect 4860 235 4940 315
rect 5060 235 5140 315
rect 5260 235 5340 315
rect 5460 235 5540 315
rect 5660 235 5740 315
rect 5860 235 5940 315
rect 6060 235 6140 315
rect 6260 235 6340 315
rect 6460 235 6540 315
rect -140 50 -60 130
rect 60 50 140 130
rect 260 50 340 130
rect 460 50 540 130
rect 660 50 740 130
rect 860 50 940 130
rect 1060 50 1140 130
rect 1260 50 1340 130
rect 1460 50 1540 130
rect 1660 50 1740 130
rect 1860 50 1940 130
rect 2060 50 2140 130
rect 2260 50 2340 130
rect 2460 50 2540 130
rect 2660 50 2740 130
rect 2860 50 2940 130
rect 3060 50 3140 130
rect 3260 50 3340 130
rect 3460 50 3540 130
rect 3660 50 3740 130
rect 3860 50 3940 130
rect 4060 50 4140 130
rect 4260 50 4340 130
rect 4460 50 4540 130
rect 4660 50 4740 130
rect 4860 50 4940 130
rect 5060 50 5140 130
rect 5260 50 5340 130
rect 5460 50 5540 130
rect 5660 50 5740 130
rect 5860 50 5940 130
rect 6060 50 6140 130
rect 6260 50 6340 130
rect 6460 50 6540 130
rect -140 -135 -60 -55
rect 60 -135 140 -55
rect 260 -135 340 -55
rect 460 -135 540 -55
rect 660 -135 740 -55
rect 860 -135 940 -55
rect 1060 -135 1140 -55
rect 1260 -135 1340 -55
rect 1460 -135 1540 -55
rect 1660 -135 1740 -55
rect 1860 -135 1940 -55
rect 2060 -135 2140 -55
rect 2260 -135 2340 -55
rect 2460 -135 2540 -55
rect 2660 -135 2740 -55
rect 2860 -135 2940 -55
rect 3060 -135 3140 -55
rect 3260 -135 3340 -55
rect 3460 -135 3540 -55
rect 3660 -135 3740 -55
rect 3860 -135 3940 -55
rect 4060 -135 4140 -55
rect 4260 -135 4340 -55
rect 4460 -135 4540 -55
rect 4660 -135 4740 -55
rect 4860 -135 4940 -55
rect 5060 -135 5140 -55
rect 5260 -135 5340 -55
rect 5460 -135 5540 -55
rect 5660 -135 5740 -55
rect 5860 -135 5940 -55
rect 6060 -135 6140 -55
rect 6260 -135 6340 -55
rect 6460 -135 6540 -55
<< metal4 >>
rect -150 12095 -50 12100
rect -150 12055 -145 12095
rect -105 12055 -95 12095
rect -55 12055 -50 12095
rect -150 12050 -50 12055
rect -115 11980 -85 12050
rect 85 11980 115 12025
rect 285 11980 315 12025
rect 485 11980 515 12025
rect 685 11980 715 12025
rect 885 11980 915 12025
rect 1085 11980 1115 12025
rect 1285 11980 1315 12025
rect 1485 11980 1515 12025
rect 1685 11980 1715 12025
rect 1885 11980 1915 12025
rect 2085 11980 2115 12025
rect 2285 11980 2315 12025
rect 2485 11980 2515 12025
rect 2685 11980 2715 12025
rect 2885 11980 2915 12025
rect 3085 11980 3115 12025
rect 3285 11980 3315 12025
rect 3485 11980 3515 12025
rect 3685 11980 3715 12025
rect 3885 11980 3915 12025
rect 4085 11980 4115 12025
rect 4285 11980 4315 12025
rect 4485 11980 4515 12025
rect 4685 11980 4715 12025
rect 4885 11980 4915 12025
rect 5085 11980 5115 12025
rect 5285 11980 5315 12025
rect 5485 11980 5515 12025
rect 5685 11980 5715 12025
rect 5885 11980 5915 12025
rect 6085 11980 6115 12025
rect 6285 11980 6315 12075
rect 6450 12070 6550 12075
rect 6450 12030 6455 12070
rect 6495 12030 6505 12070
rect 6545 12030 6550 12070
rect 6450 12025 6550 12030
rect 6485 11980 6515 12025
rect -150 11970 -50 11980
rect -150 11890 -140 11970
rect -60 11890 -50 11970
rect -150 11880 -50 11890
rect 50 11970 150 11980
rect 50 11890 60 11970
rect 140 11945 150 11970
rect 250 11970 350 11980
rect 250 11945 260 11970
rect 140 11915 260 11945
rect 140 11890 150 11915
rect 50 11880 150 11890
rect 250 11890 260 11915
rect 340 11945 350 11970
rect 450 11970 550 11980
rect 450 11945 460 11970
rect 340 11915 460 11945
rect 340 11890 350 11915
rect 250 11880 350 11890
rect 450 11890 460 11915
rect 540 11945 550 11970
rect 650 11970 750 11980
rect 650 11945 660 11970
rect 540 11915 660 11945
rect 540 11890 550 11915
rect 450 11880 550 11890
rect 650 11890 660 11915
rect 740 11945 750 11970
rect 850 11970 950 11980
rect 850 11945 860 11970
rect 740 11915 860 11945
rect 740 11890 750 11915
rect 650 11880 750 11890
rect 850 11890 860 11915
rect 940 11945 950 11970
rect 1050 11970 1150 11980
rect 1050 11945 1060 11970
rect 940 11915 1060 11945
rect 940 11890 950 11915
rect 850 11880 950 11890
rect 1050 11890 1060 11915
rect 1140 11945 1150 11970
rect 1250 11970 1350 11980
rect 1250 11945 1260 11970
rect 1140 11915 1260 11945
rect 1140 11890 1150 11915
rect 1050 11880 1150 11890
rect 1250 11890 1260 11915
rect 1340 11945 1350 11970
rect 1450 11970 1550 11980
rect 1450 11945 1460 11970
rect 1340 11915 1460 11945
rect 1340 11890 1350 11915
rect 1250 11880 1350 11890
rect 1450 11890 1460 11915
rect 1540 11945 1550 11970
rect 1650 11970 1750 11980
rect 1650 11945 1660 11970
rect 1540 11915 1660 11945
rect 1540 11890 1550 11915
rect 1450 11880 1550 11890
rect 1650 11890 1660 11915
rect 1740 11945 1750 11970
rect 1850 11970 1950 11980
rect 1850 11945 1860 11970
rect 1740 11915 1860 11945
rect 1740 11890 1750 11915
rect 1650 11880 1750 11890
rect 1850 11890 1860 11915
rect 1940 11945 1950 11970
rect 2050 11970 2150 11980
rect 2050 11945 2060 11970
rect 1940 11915 2060 11945
rect 1940 11890 1950 11915
rect 1850 11880 1950 11890
rect 2050 11890 2060 11915
rect 2140 11945 2150 11970
rect 2250 11970 2350 11980
rect 2250 11945 2260 11970
rect 2140 11915 2260 11945
rect 2140 11890 2150 11915
rect 2050 11880 2150 11890
rect 2250 11890 2260 11915
rect 2340 11945 2350 11970
rect 2450 11970 2550 11980
rect 2450 11945 2460 11970
rect 2340 11915 2460 11945
rect 2340 11890 2350 11915
rect 2250 11880 2350 11890
rect 2450 11890 2460 11915
rect 2540 11945 2550 11970
rect 2650 11970 2750 11980
rect 2650 11945 2660 11970
rect 2540 11915 2660 11945
rect 2540 11890 2550 11915
rect 2450 11880 2550 11890
rect 2650 11890 2660 11915
rect 2740 11945 2750 11970
rect 2850 11970 2950 11980
rect 2850 11945 2860 11970
rect 2740 11915 2860 11945
rect 2740 11890 2750 11915
rect 2650 11880 2750 11890
rect 2850 11890 2860 11915
rect 2940 11945 2950 11970
rect 3050 11970 3150 11980
rect 3050 11945 3060 11970
rect 2940 11915 3060 11945
rect 2940 11890 2950 11915
rect 2850 11880 2950 11890
rect 3050 11890 3060 11915
rect 3140 11945 3150 11970
rect 3250 11970 3350 11980
rect 3250 11945 3260 11970
rect 3140 11915 3260 11945
rect 3140 11890 3150 11915
rect 3050 11880 3150 11890
rect 3250 11890 3260 11915
rect 3340 11945 3350 11970
rect 3450 11970 3550 11980
rect 3450 11945 3460 11970
rect 3340 11915 3460 11945
rect 3340 11890 3350 11915
rect 3250 11880 3350 11890
rect 3450 11890 3460 11915
rect 3540 11945 3550 11970
rect 3650 11970 3750 11980
rect 3650 11945 3660 11970
rect 3540 11915 3660 11945
rect 3540 11890 3550 11915
rect 3450 11880 3550 11890
rect 3650 11890 3660 11915
rect 3740 11945 3750 11970
rect 3850 11970 3950 11980
rect 3850 11945 3860 11970
rect 3740 11915 3860 11945
rect 3740 11890 3750 11915
rect 3650 11880 3750 11890
rect 3850 11890 3860 11915
rect 3940 11945 3950 11970
rect 4050 11970 4150 11980
rect 4050 11945 4060 11970
rect 3940 11915 4060 11945
rect 3940 11890 3950 11915
rect 3850 11880 3950 11890
rect 4050 11890 4060 11915
rect 4140 11945 4150 11970
rect 4250 11970 4350 11980
rect 4250 11945 4260 11970
rect 4140 11915 4260 11945
rect 4140 11890 4150 11915
rect 4050 11880 4150 11890
rect 4250 11890 4260 11915
rect 4340 11945 4350 11970
rect 4450 11970 4550 11980
rect 4450 11945 4460 11970
rect 4340 11915 4460 11945
rect 4340 11890 4350 11915
rect 4250 11880 4350 11890
rect 4450 11890 4460 11915
rect 4540 11945 4550 11970
rect 4650 11970 4750 11980
rect 4650 11945 4660 11970
rect 4540 11915 4660 11945
rect 4540 11890 4550 11915
rect 4450 11880 4550 11890
rect 4650 11890 4660 11915
rect 4740 11945 4750 11970
rect 4850 11970 4950 11980
rect 4850 11945 4860 11970
rect 4740 11915 4860 11945
rect 4740 11890 4750 11915
rect 4650 11880 4750 11890
rect 4850 11890 4860 11915
rect 4940 11945 4950 11970
rect 5050 11970 5150 11980
rect 5050 11945 5060 11970
rect 4940 11915 5060 11945
rect 4940 11890 4950 11915
rect 4850 11880 4950 11890
rect 5050 11890 5060 11915
rect 5140 11945 5150 11970
rect 5250 11970 5350 11980
rect 5250 11945 5260 11970
rect 5140 11915 5260 11945
rect 5140 11890 5150 11915
rect 5050 11880 5150 11890
rect 5250 11890 5260 11915
rect 5340 11945 5350 11970
rect 5450 11970 5550 11980
rect 5450 11945 5460 11970
rect 5340 11915 5460 11945
rect 5340 11890 5350 11915
rect 5250 11880 5350 11890
rect 5450 11890 5460 11915
rect 5540 11945 5550 11970
rect 5650 11970 5750 11980
rect 5650 11945 5660 11970
rect 5540 11915 5660 11945
rect 5540 11890 5550 11915
rect 5450 11880 5550 11890
rect 5650 11890 5660 11915
rect 5740 11945 5750 11970
rect 5850 11970 5950 11980
rect 5850 11945 5860 11970
rect 5740 11915 5860 11945
rect 5740 11890 5750 11915
rect 5650 11880 5750 11890
rect 5850 11890 5860 11915
rect 5940 11945 5950 11970
rect 6050 11970 6150 11980
rect 6050 11945 6060 11970
rect 5940 11915 6060 11945
rect 5940 11890 5950 11915
rect 5850 11880 5950 11890
rect 6050 11890 6060 11915
rect 6140 11945 6150 11970
rect 6250 11970 6350 11980
rect 6250 11945 6260 11970
rect 6140 11915 6260 11945
rect 6140 11890 6150 11915
rect 6050 11880 6150 11890
rect 6250 11890 6260 11915
rect 6340 11890 6350 11970
rect 6250 11880 6350 11890
rect 6450 11970 6550 11980
rect 6450 11890 6460 11970
rect 6540 11890 6550 11970
rect 6450 11880 6550 11890
rect -115 11795 -85 11880
rect 85 11795 115 11880
rect 285 11795 315 11880
rect 485 11795 515 11880
rect 685 11795 715 11880
rect 885 11795 915 11880
rect 1085 11795 1115 11880
rect 1285 11795 1315 11880
rect 1485 11795 1515 11880
rect 1685 11795 1715 11880
rect 1885 11795 1915 11880
rect 2085 11795 2115 11880
rect 2285 11795 2315 11880
rect 2485 11795 2515 11880
rect 2685 11795 2715 11880
rect 2885 11795 2915 11880
rect 3085 11795 3115 11880
rect 3285 11795 3315 11880
rect 3485 11795 3515 11880
rect 3685 11795 3715 11880
rect 3885 11795 3915 11880
rect 4085 11795 4115 11880
rect 4285 11795 4315 11880
rect 4485 11795 4515 11880
rect 4685 11795 4715 11880
rect 4885 11795 4915 11880
rect 5085 11795 5115 11880
rect 5285 11795 5315 11880
rect 5485 11795 5515 11880
rect 5685 11795 5715 11880
rect 5885 11795 5915 11880
rect 6085 11795 6115 11880
rect 6285 11795 6315 11880
rect 6485 11795 6515 11880
rect -150 11785 -50 11795
rect -150 11705 -140 11785
rect -60 11705 -50 11785
rect -150 11695 -50 11705
rect 50 11785 150 11795
rect 50 11705 60 11785
rect 140 11705 150 11785
rect 50 11695 150 11705
rect 250 11785 350 11795
rect 250 11705 260 11785
rect 340 11705 350 11785
rect 250 11695 350 11705
rect 450 11785 550 11795
rect 450 11705 460 11785
rect 540 11705 550 11785
rect 450 11695 550 11705
rect 650 11785 750 11795
rect 650 11705 660 11785
rect 740 11705 750 11785
rect 650 11695 750 11705
rect 850 11785 950 11795
rect 850 11705 860 11785
rect 940 11705 950 11785
rect 850 11695 950 11705
rect 1050 11785 1150 11795
rect 1050 11705 1060 11785
rect 1140 11705 1150 11785
rect 1050 11695 1150 11705
rect 1250 11785 1350 11795
rect 1250 11705 1260 11785
rect 1340 11705 1350 11785
rect 1250 11695 1350 11705
rect 1450 11785 1550 11795
rect 1450 11705 1460 11785
rect 1540 11705 1550 11785
rect 1450 11695 1550 11705
rect 1650 11785 1750 11795
rect 1650 11705 1660 11785
rect 1740 11705 1750 11785
rect 1650 11695 1750 11705
rect 1850 11785 1950 11795
rect 1850 11705 1860 11785
rect 1940 11705 1950 11785
rect 1850 11695 1950 11705
rect 2050 11785 2150 11795
rect 2050 11705 2060 11785
rect 2140 11705 2150 11785
rect 2050 11695 2150 11705
rect 2250 11785 2350 11795
rect 2250 11705 2260 11785
rect 2340 11705 2350 11785
rect 2250 11695 2350 11705
rect 2450 11785 2550 11795
rect 2450 11705 2460 11785
rect 2540 11705 2550 11785
rect 2450 11695 2550 11705
rect 2650 11785 2750 11795
rect 2650 11705 2660 11785
rect 2740 11705 2750 11785
rect 2650 11695 2750 11705
rect 2850 11785 2950 11795
rect 2850 11705 2860 11785
rect 2940 11705 2950 11785
rect 2850 11695 2950 11705
rect 3050 11785 3150 11795
rect 3050 11705 3060 11785
rect 3140 11705 3150 11785
rect 3050 11695 3150 11705
rect 3250 11785 3350 11795
rect 3250 11705 3260 11785
rect 3340 11705 3350 11785
rect 3250 11695 3350 11705
rect 3450 11785 3550 11795
rect 3450 11705 3460 11785
rect 3540 11705 3550 11785
rect 3450 11695 3550 11705
rect 3650 11785 3750 11795
rect 3650 11705 3660 11785
rect 3740 11705 3750 11785
rect 3650 11695 3750 11705
rect 3850 11785 3950 11795
rect 3850 11705 3860 11785
rect 3940 11705 3950 11785
rect 3850 11695 3950 11705
rect 4050 11785 4150 11795
rect 4050 11705 4060 11785
rect 4140 11705 4150 11785
rect 4050 11695 4150 11705
rect 4250 11785 4350 11795
rect 4250 11705 4260 11785
rect 4340 11705 4350 11785
rect 4250 11695 4350 11705
rect 4450 11785 4550 11795
rect 4450 11705 4460 11785
rect 4540 11705 4550 11785
rect 4450 11695 4550 11705
rect 4650 11785 4750 11795
rect 4650 11705 4660 11785
rect 4740 11705 4750 11785
rect 4650 11695 4750 11705
rect 4850 11785 4950 11795
rect 4850 11705 4860 11785
rect 4940 11705 4950 11785
rect 4850 11695 4950 11705
rect 5050 11785 5150 11795
rect 5050 11705 5060 11785
rect 5140 11705 5150 11785
rect 5050 11695 5150 11705
rect 5250 11785 5350 11795
rect 5250 11705 5260 11785
rect 5340 11705 5350 11785
rect 5250 11695 5350 11705
rect 5450 11785 5550 11795
rect 5450 11705 5460 11785
rect 5540 11705 5550 11785
rect 5450 11695 5550 11705
rect 5650 11785 5750 11795
rect 5650 11705 5660 11785
rect 5740 11705 5750 11785
rect 5650 11695 5750 11705
rect 5850 11785 5950 11795
rect 5850 11705 5860 11785
rect 5940 11705 5950 11785
rect 5850 11695 5950 11705
rect 6050 11785 6150 11795
rect 6050 11705 6060 11785
rect 6140 11705 6150 11785
rect 6050 11695 6150 11705
rect 6250 11785 6350 11795
rect 6250 11705 6260 11785
rect 6340 11705 6350 11785
rect 6250 11695 6350 11705
rect 6450 11785 6550 11795
rect 6450 11705 6460 11785
rect 6540 11705 6550 11785
rect 6450 11695 6550 11705
rect -115 11610 -85 11695
rect 85 11610 115 11695
rect 285 11610 315 11695
rect 485 11610 515 11695
rect 685 11610 715 11695
rect 885 11610 915 11695
rect 1085 11610 1115 11695
rect 1285 11610 1315 11695
rect 1485 11610 1515 11695
rect 1685 11610 1715 11695
rect 1885 11610 1915 11695
rect 2085 11610 2115 11695
rect 2285 11610 2315 11695
rect 2485 11610 2515 11695
rect 2685 11610 2715 11695
rect 2885 11610 2915 11695
rect 3085 11610 3115 11695
rect 3285 11610 3315 11695
rect 3485 11610 3515 11695
rect 3685 11610 3715 11695
rect 3885 11610 3915 11695
rect 4085 11610 4115 11695
rect 4285 11610 4315 11695
rect 4485 11610 4515 11695
rect 4685 11610 4715 11695
rect 4885 11610 4915 11695
rect 5085 11610 5115 11695
rect 5285 11610 5315 11695
rect 5485 11610 5515 11695
rect 5685 11610 5715 11695
rect 5885 11610 5915 11695
rect 6085 11610 6115 11695
rect 6285 11610 6315 11695
rect 6485 11610 6515 11695
rect -150 11600 -50 11610
rect -150 11520 -140 11600
rect -60 11520 -50 11600
rect -150 11510 -50 11520
rect 50 11600 150 11610
rect 50 11520 60 11600
rect 140 11520 150 11600
rect 50 11510 150 11520
rect 250 11600 350 11610
rect 250 11520 260 11600
rect 340 11520 350 11600
rect 250 11510 350 11520
rect 450 11600 550 11610
rect 450 11520 460 11600
rect 540 11520 550 11600
rect 450 11510 550 11520
rect 650 11600 750 11610
rect 650 11520 660 11600
rect 740 11520 750 11600
rect 650 11510 750 11520
rect 850 11600 950 11610
rect 850 11520 860 11600
rect 940 11520 950 11600
rect 850 11510 950 11520
rect 1050 11600 1150 11610
rect 1050 11520 1060 11600
rect 1140 11520 1150 11600
rect 1050 11510 1150 11520
rect 1250 11600 1350 11610
rect 1250 11520 1260 11600
rect 1340 11520 1350 11600
rect 1250 11510 1350 11520
rect 1450 11600 1550 11610
rect 1450 11520 1460 11600
rect 1540 11520 1550 11600
rect 1450 11510 1550 11520
rect 1650 11600 1750 11610
rect 1650 11520 1660 11600
rect 1740 11520 1750 11600
rect 1650 11510 1750 11520
rect 1850 11600 1950 11610
rect 1850 11520 1860 11600
rect 1940 11520 1950 11600
rect 1850 11510 1950 11520
rect 2050 11600 2150 11610
rect 2050 11520 2060 11600
rect 2140 11520 2150 11600
rect 2050 11510 2150 11520
rect 2250 11600 2350 11610
rect 2250 11520 2260 11600
rect 2340 11520 2350 11600
rect 2250 11510 2350 11520
rect 2450 11600 2550 11610
rect 2450 11520 2460 11600
rect 2540 11520 2550 11600
rect 2450 11510 2550 11520
rect 2650 11600 2750 11610
rect 2650 11520 2660 11600
rect 2740 11520 2750 11600
rect 2650 11510 2750 11520
rect 2850 11600 2950 11610
rect 2850 11520 2860 11600
rect 2940 11520 2950 11600
rect 2850 11510 2950 11520
rect 3050 11600 3150 11610
rect 3050 11520 3060 11600
rect 3140 11520 3150 11600
rect 3050 11510 3150 11520
rect 3250 11600 3350 11610
rect 3250 11520 3260 11600
rect 3340 11520 3350 11600
rect 3250 11510 3350 11520
rect 3450 11600 3550 11610
rect 3450 11520 3460 11600
rect 3540 11520 3550 11600
rect 3450 11510 3550 11520
rect 3650 11600 3750 11610
rect 3650 11520 3660 11600
rect 3740 11520 3750 11600
rect 3650 11510 3750 11520
rect 3850 11600 3950 11610
rect 3850 11520 3860 11600
rect 3940 11520 3950 11600
rect 3850 11510 3950 11520
rect 4050 11600 4150 11610
rect 4050 11520 4060 11600
rect 4140 11520 4150 11600
rect 4050 11510 4150 11520
rect 4250 11600 4350 11610
rect 4250 11520 4260 11600
rect 4340 11520 4350 11600
rect 4250 11510 4350 11520
rect 4450 11600 4550 11610
rect 4450 11520 4460 11600
rect 4540 11520 4550 11600
rect 4450 11510 4550 11520
rect 4650 11600 4750 11610
rect 4650 11520 4660 11600
rect 4740 11520 4750 11600
rect 4650 11510 4750 11520
rect 4850 11600 4950 11610
rect 4850 11520 4860 11600
rect 4940 11520 4950 11600
rect 4850 11510 4950 11520
rect 5050 11600 5150 11610
rect 5050 11520 5060 11600
rect 5140 11520 5150 11600
rect 5050 11510 5150 11520
rect 5250 11600 5350 11610
rect 5250 11520 5260 11600
rect 5340 11520 5350 11600
rect 5250 11510 5350 11520
rect 5450 11600 5550 11610
rect 5450 11520 5460 11600
rect 5540 11520 5550 11600
rect 5450 11510 5550 11520
rect 5650 11600 5750 11610
rect 5650 11520 5660 11600
rect 5740 11520 5750 11600
rect 5650 11510 5750 11520
rect 5850 11600 5950 11610
rect 5850 11520 5860 11600
rect 5940 11520 5950 11600
rect 5850 11510 5950 11520
rect 6050 11600 6150 11610
rect 6050 11520 6060 11600
rect 6140 11520 6150 11600
rect 6050 11510 6150 11520
rect 6250 11600 6350 11610
rect 6250 11520 6260 11600
rect 6340 11520 6350 11600
rect 6250 11510 6350 11520
rect 6450 11600 6550 11610
rect 6450 11520 6460 11600
rect 6540 11520 6550 11600
rect 6450 11510 6550 11520
rect -115 11425 -85 11510
rect 85 11425 115 11510
rect 285 11425 315 11510
rect 485 11425 515 11510
rect 685 11425 715 11510
rect 885 11425 915 11510
rect 1085 11425 1115 11510
rect 1285 11425 1315 11510
rect 1485 11425 1515 11510
rect 1685 11425 1715 11510
rect 1885 11425 1915 11510
rect 2085 11425 2115 11510
rect 2285 11425 2315 11510
rect 2485 11425 2515 11510
rect 2685 11425 2715 11510
rect 2885 11425 2915 11510
rect 3085 11425 3115 11510
rect 3285 11425 3315 11510
rect 3485 11425 3515 11510
rect 3685 11425 3715 11510
rect 3885 11425 3915 11510
rect 4085 11425 4115 11510
rect 4285 11425 4315 11510
rect 4485 11425 4515 11510
rect 4685 11425 4715 11510
rect 4885 11425 4915 11510
rect 5085 11425 5115 11510
rect 5285 11425 5315 11510
rect 5485 11425 5515 11510
rect 5685 11425 5715 11510
rect 5885 11425 5915 11510
rect 6085 11425 6115 11510
rect 6285 11425 6315 11510
rect 6485 11425 6515 11510
rect -150 11415 -50 11425
rect -150 11335 -140 11415
rect -60 11335 -50 11415
rect -150 11325 -50 11335
rect 50 11415 150 11425
rect 50 11335 60 11415
rect 140 11335 150 11415
rect 50 11325 150 11335
rect 250 11415 350 11425
rect 250 11335 260 11415
rect 340 11335 350 11415
rect 250 11325 350 11335
rect 450 11415 550 11425
rect 450 11335 460 11415
rect 540 11335 550 11415
rect 450 11325 550 11335
rect 650 11415 750 11425
rect 650 11335 660 11415
rect 740 11335 750 11415
rect 650 11325 750 11335
rect 850 11415 950 11425
rect 850 11335 860 11415
rect 940 11335 950 11415
rect 850 11325 950 11335
rect 1050 11415 1150 11425
rect 1050 11335 1060 11415
rect 1140 11335 1150 11415
rect 1050 11325 1150 11335
rect 1250 11415 1350 11425
rect 1250 11335 1260 11415
rect 1340 11335 1350 11415
rect 1250 11325 1350 11335
rect 1450 11415 1550 11425
rect 1450 11335 1460 11415
rect 1540 11335 1550 11415
rect 1450 11325 1550 11335
rect 1650 11415 1750 11425
rect 1650 11335 1660 11415
rect 1740 11335 1750 11415
rect 1650 11325 1750 11335
rect 1850 11415 1950 11425
rect 1850 11335 1860 11415
rect 1940 11335 1950 11415
rect 1850 11325 1950 11335
rect 2050 11415 2150 11425
rect 2050 11335 2060 11415
rect 2140 11335 2150 11415
rect 2050 11325 2150 11335
rect 2250 11415 2350 11425
rect 2250 11335 2260 11415
rect 2340 11335 2350 11415
rect 2250 11325 2350 11335
rect 2450 11415 2550 11425
rect 2450 11335 2460 11415
rect 2540 11335 2550 11415
rect 2450 11325 2550 11335
rect 2650 11415 2750 11425
rect 2650 11335 2660 11415
rect 2740 11335 2750 11415
rect 2650 11325 2750 11335
rect 2850 11415 2950 11425
rect 2850 11335 2860 11415
rect 2940 11335 2950 11415
rect 2850 11325 2950 11335
rect 3050 11415 3150 11425
rect 3050 11335 3060 11415
rect 3140 11335 3150 11415
rect 3050 11325 3150 11335
rect 3250 11415 3350 11425
rect 3250 11335 3260 11415
rect 3340 11335 3350 11415
rect 3250 11325 3350 11335
rect 3450 11415 3550 11425
rect 3450 11335 3460 11415
rect 3540 11335 3550 11415
rect 3450 11325 3550 11335
rect 3650 11415 3750 11425
rect 3650 11335 3660 11415
rect 3740 11335 3750 11415
rect 3650 11325 3750 11335
rect 3850 11415 3950 11425
rect 3850 11335 3860 11415
rect 3940 11335 3950 11415
rect 3850 11325 3950 11335
rect 4050 11415 4150 11425
rect 4050 11335 4060 11415
rect 4140 11335 4150 11415
rect 4050 11325 4150 11335
rect 4250 11415 4350 11425
rect 4250 11335 4260 11415
rect 4340 11335 4350 11415
rect 4250 11325 4350 11335
rect 4450 11415 4550 11425
rect 4450 11335 4460 11415
rect 4540 11335 4550 11415
rect 4450 11325 4550 11335
rect 4650 11415 4750 11425
rect 4650 11335 4660 11415
rect 4740 11335 4750 11415
rect 4650 11325 4750 11335
rect 4850 11415 4950 11425
rect 4850 11335 4860 11415
rect 4940 11335 4950 11415
rect 4850 11325 4950 11335
rect 5050 11415 5150 11425
rect 5050 11335 5060 11415
rect 5140 11335 5150 11415
rect 5050 11325 5150 11335
rect 5250 11415 5350 11425
rect 5250 11335 5260 11415
rect 5340 11335 5350 11415
rect 5250 11325 5350 11335
rect 5450 11415 5550 11425
rect 5450 11335 5460 11415
rect 5540 11335 5550 11415
rect 5450 11325 5550 11335
rect 5650 11415 5750 11425
rect 5650 11335 5660 11415
rect 5740 11335 5750 11415
rect 5650 11325 5750 11335
rect 5850 11415 5950 11425
rect 5850 11335 5860 11415
rect 5940 11335 5950 11415
rect 5850 11325 5950 11335
rect 6050 11415 6150 11425
rect 6050 11335 6060 11415
rect 6140 11335 6150 11415
rect 6050 11325 6150 11335
rect 6250 11415 6350 11425
rect 6250 11335 6260 11415
rect 6340 11335 6350 11415
rect 6250 11325 6350 11335
rect 6450 11415 6550 11425
rect 6450 11335 6460 11415
rect 6540 11335 6550 11415
rect 6450 11325 6550 11335
rect -115 11240 -85 11325
rect 85 11240 115 11325
rect 285 11240 315 11325
rect 485 11240 515 11325
rect 685 11240 715 11325
rect 885 11240 915 11325
rect 1085 11240 1115 11325
rect 1285 11240 1315 11325
rect 1485 11240 1515 11325
rect 1685 11240 1715 11325
rect 1885 11240 1915 11325
rect 2085 11240 2115 11325
rect 2285 11240 2315 11325
rect 2485 11240 2515 11325
rect 2685 11240 2715 11325
rect 2885 11240 2915 11325
rect 3085 11240 3115 11325
rect 3285 11240 3315 11325
rect 3485 11240 3515 11325
rect 3685 11240 3715 11325
rect 3885 11240 3915 11325
rect 4085 11240 4115 11325
rect 4285 11240 4315 11325
rect 4485 11240 4515 11325
rect 4685 11240 4715 11325
rect 4885 11240 4915 11325
rect 5085 11240 5115 11325
rect 5285 11240 5315 11325
rect 5485 11240 5515 11325
rect 5685 11240 5715 11325
rect 5885 11240 5915 11325
rect 6085 11240 6115 11325
rect 6285 11240 6315 11325
rect 6485 11240 6515 11325
rect -150 11230 -50 11240
rect -150 11150 -140 11230
rect -60 11150 -50 11230
rect -150 11140 -50 11150
rect 50 11230 150 11240
rect 50 11150 60 11230
rect 140 11150 150 11230
rect 50 11140 150 11150
rect 250 11230 350 11240
rect 250 11150 260 11230
rect 340 11150 350 11230
rect 250 11140 350 11150
rect 450 11230 550 11240
rect 450 11150 460 11230
rect 540 11150 550 11230
rect 450 11140 550 11150
rect 650 11230 750 11240
rect 650 11150 660 11230
rect 740 11150 750 11230
rect 650 11140 750 11150
rect 850 11230 950 11240
rect 850 11150 860 11230
rect 940 11150 950 11230
rect 850 11140 950 11150
rect 1050 11230 1150 11240
rect 1050 11150 1060 11230
rect 1140 11150 1150 11230
rect 1050 11140 1150 11150
rect 1250 11230 1350 11240
rect 1250 11150 1260 11230
rect 1340 11150 1350 11230
rect 1250 11140 1350 11150
rect 1450 11230 1550 11240
rect 1450 11150 1460 11230
rect 1540 11150 1550 11230
rect 1450 11140 1550 11150
rect 1650 11230 1750 11240
rect 1650 11150 1660 11230
rect 1740 11150 1750 11230
rect 1650 11140 1750 11150
rect 1850 11230 1950 11240
rect 1850 11150 1860 11230
rect 1940 11150 1950 11230
rect 1850 11140 1950 11150
rect 2050 11230 2150 11240
rect 2050 11150 2060 11230
rect 2140 11150 2150 11230
rect 2050 11140 2150 11150
rect 2250 11230 2350 11240
rect 2250 11150 2260 11230
rect 2340 11150 2350 11230
rect 2250 11140 2350 11150
rect 2450 11230 2550 11240
rect 2450 11150 2460 11230
rect 2540 11150 2550 11230
rect 2450 11140 2550 11150
rect 2650 11230 2750 11240
rect 2650 11150 2660 11230
rect 2740 11150 2750 11230
rect 2650 11140 2750 11150
rect 2850 11230 2950 11240
rect 2850 11150 2860 11230
rect 2940 11150 2950 11230
rect 2850 11140 2950 11150
rect 3050 11230 3150 11240
rect 3050 11150 3060 11230
rect 3140 11150 3150 11230
rect 3050 11140 3150 11150
rect 3250 11230 3350 11240
rect 3250 11150 3260 11230
rect 3340 11150 3350 11230
rect 3250 11140 3350 11150
rect 3450 11230 3550 11240
rect 3450 11150 3460 11230
rect 3540 11150 3550 11230
rect 3450 11140 3550 11150
rect 3650 11230 3750 11240
rect 3650 11150 3660 11230
rect 3740 11150 3750 11230
rect 3650 11140 3750 11150
rect 3850 11230 3950 11240
rect 3850 11150 3860 11230
rect 3940 11150 3950 11230
rect 3850 11140 3950 11150
rect 4050 11230 4150 11240
rect 4050 11150 4060 11230
rect 4140 11150 4150 11230
rect 4050 11140 4150 11150
rect 4250 11230 4350 11240
rect 4250 11150 4260 11230
rect 4340 11150 4350 11230
rect 4250 11140 4350 11150
rect 4450 11230 4550 11240
rect 4450 11150 4460 11230
rect 4540 11150 4550 11230
rect 4450 11140 4550 11150
rect 4650 11230 4750 11240
rect 4650 11150 4660 11230
rect 4740 11150 4750 11230
rect 4650 11140 4750 11150
rect 4850 11230 4950 11240
rect 4850 11150 4860 11230
rect 4940 11150 4950 11230
rect 4850 11140 4950 11150
rect 5050 11230 5150 11240
rect 5050 11150 5060 11230
rect 5140 11150 5150 11230
rect 5050 11140 5150 11150
rect 5250 11230 5350 11240
rect 5250 11150 5260 11230
rect 5340 11150 5350 11230
rect 5250 11140 5350 11150
rect 5450 11230 5550 11240
rect 5450 11150 5460 11230
rect 5540 11150 5550 11230
rect 5450 11140 5550 11150
rect 5650 11230 5750 11240
rect 5650 11150 5660 11230
rect 5740 11150 5750 11230
rect 5650 11140 5750 11150
rect 5850 11230 5950 11240
rect 5850 11150 5860 11230
rect 5940 11150 5950 11230
rect 5850 11140 5950 11150
rect 6050 11230 6150 11240
rect 6050 11150 6060 11230
rect 6140 11150 6150 11230
rect 6050 11140 6150 11150
rect 6250 11230 6350 11240
rect 6250 11150 6260 11230
rect 6340 11150 6350 11230
rect 6250 11140 6350 11150
rect 6450 11230 6550 11240
rect 6450 11150 6460 11230
rect 6540 11150 6550 11230
rect 6450 11140 6550 11150
rect -115 11055 -85 11140
rect 85 11055 115 11140
rect 285 11055 315 11140
rect 485 11055 515 11140
rect 685 11055 715 11140
rect 885 11055 915 11140
rect 1085 11055 1115 11140
rect 1285 11055 1315 11140
rect 1485 11055 1515 11140
rect 1685 11055 1715 11140
rect 1885 11055 1915 11140
rect 2085 11055 2115 11140
rect 2285 11055 2315 11140
rect 2485 11055 2515 11140
rect 2685 11055 2715 11140
rect 2885 11055 2915 11140
rect 3085 11055 3115 11140
rect 3285 11055 3315 11140
rect 3485 11055 3515 11140
rect 3685 11055 3715 11140
rect 3885 11055 3915 11140
rect 4085 11055 4115 11140
rect 4285 11055 4315 11140
rect 4485 11055 4515 11140
rect 4685 11055 4715 11140
rect 4885 11055 4915 11140
rect 5085 11055 5115 11140
rect 5285 11055 5315 11140
rect 5485 11055 5515 11140
rect 5685 11055 5715 11140
rect 5885 11055 5915 11140
rect 6085 11055 6115 11140
rect 6285 11055 6315 11140
rect 6485 11055 6515 11140
rect -150 11045 -50 11055
rect -150 10965 -140 11045
rect -60 10965 -50 11045
rect -150 10955 -50 10965
rect 50 11045 150 11055
rect 50 10965 60 11045
rect 140 10965 150 11045
rect 50 10955 150 10965
rect 250 11045 350 11055
rect 250 10965 260 11045
rect 340 10965 350 11045
rect 250 10955 350 10965
rect 450 11045 550 11055
rect 450 10965 460 11045
rect 540 10965 550 11045
rect 450 10955 550 10965
rect 650 11045 750 11055
rect 650 10965 660 11045
rect 740 10965 750 11045
rect 650 10955 750 10965
rect 850 11045 950 11055
rect 850 10965 860 11045
rect 940 10965 950 11045
rect 850 10955 950 10965
rect 1050 11045 1150 11055
rect 1050 10965 1060 11045
rect 1140 10965 1150 11045
rect 1050 10955 1150 10965
rect 1250 11045 1350 11055
rect 1250 10965 1260 11045
rect 1340 10965 1350 11045
rect 1250 10955 1350 10965
rect 1450 11045 1550 11055
rect 1450 10965 1460 11045
rect 1540 10965 1550 11045
rect 1450 10955 1550 10965
rect 1650 11045 1750 11055
rect 1650 10965 1660 11045
rect 1740 10965 1750 11045
rect 1650 10955 1750 10965
rect 1850 11045 1950 11055
rect 1850 10965 1860 11045
rect 1940 10965 1950 11045
rect 1850 10955 1950 10965
rect 2050 11045 2150 11055
rect 2050 10965 2060 11045
rect 2140 10965 2150 11045
rect 2050 10955 2150 10965
rect 2250 11045 2350 11055
rect 2250 10965 2260 11045
rect 2340 10965 2350 11045
rect 2250 10955 2350 10965
rect 2450 11045 2550 11055
rect 2450 10965 2460 11045
rect 2540 10965 2550 11045
rect 2450 10955 2550 10965
rect 2650 11045 2750 11055
rect 2650 10965 2660 11045
rect 2740 10965 2750 11045
rect 2650 10955 2750 10965
rect 2850 11045 2950 11055
rect 2850 10965 2860 11045
rect 2940 10965 2950 11045
rect 2850 10955 2950 10965
rect 3050 11045 3150 11055
rect 3050 10965 3060 11045
rect 3140 10965 3150 11045
rect 3050 10955 3150 10965
rect 3250 11045 3350 11055
rect 3250 10965 3260 11045
rect 3340 10965 3350 11045
rect 3250 10955 3350 10965
rect 3450 11045 3550 11055
rect 3450 10965 3460 11045
rect 3540 10965 3550 11045
rect 3450 10955 3550 10965
rect 3650 11045 3750 11055
rect 3650 10965 3660 11045
rect 3740 10965 3750 11045
rect 3650 10955 3750 10965
rect 3850 11045 3950 11055
rect 3850 10965 3860 11045
rect 3940 10965 3950 11045
rect 3850 10955 3950 10965
rect 4050 11045 4150 11055
rect 4050 10965 4060 11045
rect 4140 10965 4150 11045
rect 4050 10955 4150 10965
rect 4250 11045 4350 11055
rect 4250 10965 4260 11045
rect 4340 10965 4350 11045
rect 4250 10955 4350 10965
rect 4450 11045 4550 11055
rect 4450 10965 4460 11045
rect 4540 10965 4550 11045
rect 4450 10955 4550 10965
rect 4650 11045 4750 11055
rect 4650 10965 4660 11045
rect 4740 10965 4750 11045
rect 4650 10955 4750 10965
rect 4850 11045 4950 11055
rect 4850 10965 4860 11045
rect 4940 10965 4950 11045
rect 4850 10955 4950 10965
rect 5050 11045 5150 11055
rect 5050 10965 5060 11045
rect 5140 10965 5150 11045
rect 5050 10955 5150 10965
rect 5250 11045 5350 11055
rect 5250 10965 5260 11045
rect 5340 10965 5350 11045
rect 5250 10955 5350 10965
rect 5450 11045 5550 11055
rect 5450 10965 5460 11045
rect 5540 10965 5550 11045
rect 5450 10955 5550 10965
rect 5650 11045 5750 11055
rect 5650 10965 5660 11045
rect 5740 10965 5750 11045
rect 5650 10955 5750 10965
rect 5850 11045 5950 11055
rect 5850 10965 5860 11045
rect 5940 10965 5950 11045
rect 5850 10955 5950 10965
rect 6050 11045 6150 11055
rect 6050 10965 6060 11045
rect 6140 10965 6150 11045
rect 6050 10955 6150 10965
rect 6250 11045 6350 11055
rect 6250 10965 6260 11045
rect 6340 10965 6350 11045
rect 6250 10955 6350 10965
rect 6450 11045 6550 11055
rect 6450 10965 6460 11045
rect 6540 10965 6550 11045
rect 6450 10955 6550 10965
rect -115 10870 -85 10955
rect 85 10870 115 10955
rect 285 10870 315 10955
rect 485 10870 515 10955
rect 685 10870 715 10955
rect 885 10870 915 10955
rect 1085 10870 1115 10955
rect 1285 10870 1315 10955
rect 1485 10870 1515 10955
rect 1685 10870 1715 10955
rect 1885 10870 1915 10955
rect 2085 10870 2115 10955
rect 2285 10870 2315 10955
rect 2485 10870 2515 10955
rect 2685 10870 2715 10955
rect 2885 10870 2915 10955
rect 3085 10870 3115 10955
rect 3285 10870 3315 10955
rect 3485 10870 3515 10955
rect 3685 10870 3715 10955
rect 3885 10870 3915 10955
rect 4085 10870 4115 10955
rect 4285 10870 4315 10955
rect 4485 10870 4515 10955
rect 4685 10870 4715 10955
rect 4885 10870 4915 10955
rect 5085 10870 5115 10955
rect 5285 10870 5315 10955
rect 5485 10870 5515 10955
rect 5685 10870 5715 10955
rect 5885 10870 5915 10955
rect 6085 10870 6115 10955
rect 6285 10870 6315 10955
rect 6485 10870 6515 10955
rect -150 10860 -50 10870
rect -150 10780 -140 10860
rect -60 10780 -50 10860
rect -150 10770 -50 10780
rect 50 10860 150 10870
rect 50 10780 60 10860
rect 140 10780 150 10860
rect 50 10770 150 10780
rect 250 10860 350 10870
rect 250 10780 260 10860
rect 340 10780 350 10860
rect 250 10770 350 10780
rect 450 10860 550 10870
rect 450 10780 460 10860
rect 540 10780 550 10860
rect 450 10770 550 10780
rect 650 10860 750 10870
rect 650 10780 660 10860
rect 740 10780 750 10860
rect 650 10770 750 10780
rect 850 10860 950 10870
rect 850 10780 860 10860
rect 940 10780 950 10860
rect 850 10770 950 10780
rect 1050 10860 1150 10870
rect 1050 10780 1060 10860
rect 1140 10780 1150 10860
rect 1050 10770 1150 10780
rect 1250 10860 1350 10870
rect 1250 10780 1260 10860
rect 1340 10780 1350 10860
rect 1250 10770 1350 10780
rect 1450 10860 1550 10870
rect 1450 10780 1460 10860
rect 1540 10780 1550 10860
rect 1450 10770 1550 10780
rect 1650 10860 1750 10870
rect 1650 10780 1660 10860
rect 1740 10780 1750 10860
rect 1650 10770 1750 10780
rect 1850 10860 1950 10870
rect 1850 10780 1860 10860
rect 1940 10780 1950 10860
rect 1850 10770 1950 10780
rect 2050 10860 2150 10870
rect 2050 10780 2060 10860
rect 2140 10780 2150 10860
rect 2050 10770 2150 10780
rect 2250 10860 2350 10870
rect 2250 10780 2260 10860
rect 2340 10780 2350 10860
rect 2250 10770 2350 10780
rect 2450 10860 2550 10870
rect 2450 10780 2460 10860
rect 2540 10780 2550 10860
rect 2450 10770 2550 10780
rect 2650 10860 2750 10870
rect 2650 10780 2660 10860
rect 2740 10780 2750 10860
rect 2650 10770 2750 10780
rect 2850 10860 2950 10870
rect 2850 10780 2860 10860
rect 2940 10780 2950 10860
rect 2850 10770 2950 10780
rect 3050 10860 3150 10870
rect 3050 10780 3060 10860
rect 3140 10780 3150 10860
rect 3050 10770 3150 10780
rect 3250 10860 3350 10870
rect 3250 10780 3260 10860
rect 3340 10780 3350 10860
rect 3250 10770 3350 10780
rect 3450 10860 3550 10870
rect 3450 10780 3460 10860
rect 3540 10780 3550 10860
rect 3450 10770 3550 10780
rect 3650 10860 3750 10870
rect 3650 10780 3660 10860
rect 3740 10780 3750 10860
rect 3650 10770 3750 10780
rect 3850 10860 3950 10870
rect 3850 10780 3860 10860
rect 3940 10780 3950 10860
rect 3850 10770 3950 10780
rect 4050 10860 4150 10870
rect 4050 10780 4060 10860
rect 4140 10780 4150 10860
rect 4050 10770 4150 10780
rect 4250 10860 4350 10870
rect 4250 10780 4260 10860
rect 4340 10780 4350 10860
rect 4250 10770 4350 10780
rect 4450 10860 4550 10870
rect 4450 10780 4460 10860
rect 4540 10780 4550 10860
rect 4450 10770 4550 10780
rect 4650 10860 4750 10870
rect 4650 10780 4660 10860
rect 4740 10780 4750 10860
rect 4650 10770 4750 10780
rect 4850 10860 4950 10870
rect 4850 10780 4860 10860
rect 4940 10780 4950 10860
rect 4850 10770 4950 10780
rect 5050 10860 5150 10870
rect 5050 10780 5060 10860
rect 5140 10780 5150 10860
rect 5050 10770 5150 10780
rect 5250 10860 5350 10870
rect 5250 10780 5260 10860
rect 5340 10780 5350 10860
rect 5250 10770 5350 10780
rect 5450 10860 5550 10870
rect 5450 10780 5460 10860
rect 5540 10780 5550 10860
rect 5450 10770 5550 10780
rect 5650 10860 5750 10870
rect 5650 10780 5660 10860
rect 5740 10780 5750 10860
rect 5650 10770 5750 10780
rect 5850 10860 5950 10870
rect 5850 10780 5860 10860
rect 5940 10780 5950 10860
rect 5850 10770 5950 10780
rect 6050 10860 6150 10870
rect 6050 10780 6060 10860
rect 6140 10780 6150 10860
rect 6050 10770 6150 10780
rect 6250 10860 6350 10870
rect 6250 10780 6260 10860
rect 6340 10780 6350 10860
rect 6250 10770 6350 10780
rect 6450 10860 6550 10870
rect 6450 10780 6460 10860
rect 6540 10780 6550 10860
rect 6450 10770 6550 10780
rect -115 10685 -85 10770
rect 85 10685 115 10770
rect 285 10685 315 10770
rect 485 10685 515 10770
rect 685 10685 715 10770
rect 885 10685 915 10770
rect 1085 10685 1115 10770
rect 1285 10685 1315 10770
rect 1485 10685 1515 10770
rect 1685 10685 1715 10770
rect 1885 10685 1915 10770
rect 2085 10685 2115 10770
rect 2285 10685 2315 10770
rect 2485 10685 2515 10770
rect 2685 10685 2715 10770
rect 2885 10685 2915 10770
rect 3085 10685 3115 10770
rect 3285 10685 3315 10770
rect 3485 10685 3515 10770
rect 3685 10685 3715 10770
rect 3885 10685 3915 10770
rect 4085 10685 4115 10770
rect 4285 10685 4315 10770
rect 4485 10685 4515 10770
rect 4685 10685 4715 10770
rect 4885 10685 4915 10770
rect 5085 10685 5115 10770
rect 5285 10685 5315 10770
rect 5485 10685 5515 10770
rect 5685 10685 5715 10770
rect 5885 10685 5915 10770
rect 6085 10685 6115 10770
rect 6285 10685 6315 10770
rect 6485 10685 6515 10770
rect -150 10675 -50 10685
rect -150 10595 -140 10675
rect -60 10595 -50 10675
rect -150 10585 -50 10595
rect 50 10675 150 10685
rect 50 10595 60 10675
rect 140 10595 150 10675
rect 50 10585 150 10595
rect 250 10675 350 10685
rect 250 10595 260 10675
rect 340 10595 350 10675
rect 250 10585 350 10595
rect 450 10675 550 10685
rect 450 10595 460 10675
rect 540 10595 550 10675
rect 450 10585 550 10595
rect 650 10675 750 10685
rect 650 10595 660 10675
rect 740 10595 750 10675
rect 650 10585 750 10595
rect 850 10675 950 10685
rect 850 10595 860 10675
rect 940 10595 950 10675
rect 850 10585 950 10595
rect 1050 10675 1150 10685
rect 1050 10595 1060 10675
rect 1140 10595 1150 10675
rect 1050 10585 1150 10595
rect 1250 10675 1350 10685
rect 1250 10595 1260 10675
rect 1340 10595 1350 10675
rect 1250 10585 1350 10595
rect 1450 10675 1550 10685
rect 1450 10595 1460 10675
rect 1540 10595 1550 10675
rect 1450 10585 1550 10595
rect 1650 10675 1750 10685
rect 1650 10595 1660 10675
rect 1740 10595 1750 10675
rect 1650 10585 1750 10595
rect 1850 10675 1950 10685
rect 1850 10595 1860 10675
rect 1940 10595 1950 10675
rect 1850 10585 1950 10595
rect 2050 10675 2150 10685
rect 2050 10595 2060 10675
rect 2140 10595 2150 10675
rect 2050 10585 2150 10595
rect 2250 10675 2350 10685
rect 2250 10595 2260 10675
rect 2340 10595 2350 10675
rect 2250 10585 2350 10595
rect 2450 10675 2550 10685
rect 2450 10595 2460 10675
rect 2540 10595 2550 10675
rect 2450 10585 2550 10595
rect 2650 10675 2750 10685
rect 2650 10595 2660 10675
rect 2740 10595 2750 10675
rect 2650 10585 2750 10595
rect 2850 10675 2950 10685
rect 2850 10595 2860 10675
rect 2940 10595 2950 10675
rect 2850 10585 2950 10595
rect 3050 10675 3150 10685
rect 3050 10595 3060 10675
rect 3140 10595 3150 10675
rect 3050 10585 3150 10595
rect 3250 10675 3350 10685
rect 3250 10595 3260 10675
rect 3340 10595 3350 10675
rect 3250 10585 3350 10595
rect 3450 10675 3550 10685
rect 3450 10595 3460 10675
rect 3540 10595 3550 10675
rect 3450 10585 3550 10595
rect 3650 10675 3750 10685
rect 3650 10595 3660 10675
rect 3740 10595 3750 10675
rect 3650 10585 3750 10595
rect 3850 10675 3950 10685
rect 3850 10595 3860 10675
rect 3940 10595 3950 10675
rect 3850 10585 3950 10595
rect 4050 10675 4150 10685
rect 4050 10595 4060 10675
rect 4140 10595 4150 10675
rect 4050 10585 4150 10595
rect 4250 10675 4350 10685
rect 4250 10595 4260 10675
rect 4340 10595 4350 10675
rect 4250 10585 4350 10595
rect 4450 10675 4550 10685
rect 4450 10595 4460 10675
rect 4540 10595 4550 10675
rect 4450 10585 4550 10595
rect 4650 10675 4750 10685
rect 4650 10595 4660 10675
rect 4740 10595 4750 10675
rect 4650 10585 4750 10595
rect 4850 10675 4950 10685
rect 4850 10595 4860 10675
rect 4940 10595 4950 10675
rect 4850 10585 4950 10595
rect 5050 10675 5150 10685
rect 5050 10595 5060 10675
rect 5140 10595 5150 10675
rect 5050 10585 5150 10595
rect 5250 10675 5350 10685
rect 5250 10595 5260 10675
rect 5340 10595 5350 10675
rect 5250 10585 5350 10595
rect 5450 10675 5550 10685
rect 5450 10595 5460 10675
rect 5540 10595 5550 10675
rect 5450 10585 5550 10595
rect 5650 10675 5750 10685
rect 5650 10595 5660 10675
rect 5740 10595 5750 10675
rect 5650 10585 5750 10595
rect 5850 10675 5950 10685
rect 5850 10595 5860 10675
rect 5940 10595 5950 10675
rect 5850 10585 5950 10595
rect 6050 10675 6150 10685
rect 6050 10595 6060 10675
rect 6140 10595 6150 10675
rect 6050 10585 6150 10595
rect 6250 10675 6350 10685
rect 6250 10595 6260 10675
rect 6340 10595 6350 10675
rect 6250 10585 6350 10595
rect 6450 10675 6550 10685
rect 6450 10595 6460 10675
rect 6540 10595 6550 10675
rect 6450 10585 6550 10595
rect -115 10500 -85 10585
rect 85 10500 115 10585
rect 285 10500 315 10585
rect 485 10500 515 10585
rect 685 10500 715 10585
rect 885 10500 915 10585
rect 1085 10500 1115 10585
rect 1285 10500 1315 10585
rect 1485 10500 1515 10585
rect 1685 10500 1715 10585
rect 1885 10500 1915 10585
rect 2085 10500 2115 10585
rect 2285 10500 2315 10585
rect 2485 10500 2515 10585
rect 2685 10500 2715 10585
rect 2885 10500 2915 10585
rect 3085 10500 3115 10585
rect 3285 10500 3315 10585
rect 3485 10500 3515 10585
rect 3685 10500 3715 10585
rect 3885 10500 3915 10585
rect 4085 10500 4115 10585
rect 4285 10500 4315 10585
rect 4485 10500 4515 10585
rect 4685 10500 4715 10585
rect 4885 10500 4915 10585
rect 5085 10500 5115 10585
rect 5285 10500 5315 10585
rect 5485 10500 5515 10585
rect 5685 10500 5715 10585
rect 5885 10500 5915 10585
rect 6085 10500 6115 10585
rect 6285 10500 6315 10585
rect 6485 10500 6515 10585
rect -150 10490 -50 10500
rect -150 10410 -140 10490
rect -60 10410 -50 10490
rect -150 10400 -50 10410
rect 50 10490 150 10500
rect 50 10410 60 10490
rect 140 10410 150 10490
rect 50 10400 150 10410
rect 250 10490 350 10500
rect 250 10410 260 10490
rect 340 10410 350 10490
rect 250 10400 350 10410
rect 450 10490 550 10500
rect 450 10410 460 10490
rect 540 10410 550 10490
rect 450 10400 550 10410
rect 650 10490 750 10500
rect 650 10410 660 10490
rect 740 10410 750 10490
rect 650 10400 750 10410
rect 850 10490 950 10500
rect 850 10410 860 10490
rect 940 10410 950 10490
rect 850 10400 950 10410
rect 1050 10490 1150 10500
rect 1050 10410 1060 10490
rect 1140 10410 1150 10490
rect 1050 10400 1150 10410
rect 1250 10490 1350 10500
rect 1250 10410 1260 10490
rect 1340 10410 1350 10490
rect 1250 10400 1350 10410
rect 1450 10490 1550 10500
rect 1450 10410 1460 10490
rect 1540 10410 1550 10490
rect 1450 10400 1550 10410
rect 1650 10490 1750 10500
rect 1650 10410 1660 10490
rect 1740 10410 1750 10490
rect 1650 10400 1750 10410
rect 1850 10490 1950 10500
rect 1850 10410 1860 10490
rect 1940 10410 1950 10490
rect 1850 10400 1950 10410
rect 2050 10490 2150 10500
rect 2050 10410 2060 10490
rect 2140 10410 2150 10490
rect 2050 10400 2150 10410
rect 2250 10490 2350 10500
rect 2250 10410 2260 10490
rect 2340 10410 2350 10490
rect 2250 10400 2350 10410
rect 2450 10490 2550 10500
rect 2450 10410 2460 10490
rect 2540 10410 2550 10490
rect 2450 10400 2550 10410
rect 2650 10490 2750 10500
rect 2650 10410 2660 10490
rect 2740 10410 2750 10490
rect 2650 10400 2750 10410
rect 2850 10490 2950 10500
rect 2850 10410 2860 10490
rect 2940 10410 2950 10490
rect 2850 10400 2950 10410
rect 3050 10490 3150 10500
rect 3050 10410 3060 10490
rect 3140 10410 3150 10490
rect 3050 10400 3150 10410
rect 3250 10490 3350 10500
rect 3250 10410 3260 10490
rect 3340 10410 3350 10490
rect 3250 10400 3350 10410
rect 3450 10490 3550 10500
rect 3450 10410 3460 10490
rect 3540 10410 3550 10490
rect 3450 10400 3550 10410
rect 3650 10490 3750 10500
rect 3650 10410 3660 10490
rect 3740 10410 3750 10490
rect 3650 10400 3750 10410
rect 3850 10490 3950 10500
rect 3850 10410 3860 10490
rect 3940 10410 3950 10490
rect 3850 10400 3950 10410
rect 4050 10490 4150 10500
rect 4050 10410 4060 10490
rect 4140 10410 4150 10490
rect 4050 10400 4150 10410
rect 4250 10490 4350 10500
rect 4250 10410 4260 10490
rect 4340 10410 4350 10490
rect 4250 10400 4350 10410
rect 4450 10490 4550 10500
rect 4450 10410 4460 10490
rect 4540 10410 4550 10490
rect 4450 10400 4550 10410
rect 4650 10490 4750 10500
rect 4650 10410 4660 10490
rect 4740 10410 4750 10490
rect 4650 10400 4750 10410
rect 4850 10490 4950 10500
rect 4850 10410 4860 10490
rect 4940 10410 4950 10490
rect 4850 10400 4950 10410
rect 5050 10490 5150 10500
rect 5050 10410 5060 10490
rect 5140 10410 5150 10490
rect 5050 10400 5150 10410
rect 5250 10490 5350 10500
rect 5250 10410 5260 10490
rect 5340 10410 5350 10490
rect 5250 10400 5350 10410
rect 5450 10490 5550 10500
rect 5450 10410 5460 10490
rect 5540 10410 5550 10490
rect 5450 10400 5550 10410
rect 5650 10490 5750 10500
rect 5650 10410 5660 10490
rect 5740 10410 5750 10490
rect 5650 10400 5750 10410
rect 5850 10490 5950 10500
rect 5850 10410 5860 10490
rect 5940 10410 5950 10490
rect 5850 10400 5950 10410
rect 6050 10490 6150 10500
rect 6050 10410 6060 10490
rect 6140 10410 6150 10490
rect 6050 10400 6150 10410
rect 6250 10490 6350 10500
rect 6250 10410 6260 10490
rect 6340 10410 6350 10490
rect 6250 10400 6350 10410
rect 6450 10490 6550 10500
rect 6450 10410 6460 10490
rect 6540 10410 6550 10490
rect 6450 10400 6550 10410
rect -115 10315 -85 10400
rect 85 10315 115 10400
rect 285 10315 315 10400
rect 485 10315 515 10400
rect 685 10315 715 10400
rect 885 10315 915 10400
rect 1085 10315 1115 10400
rect 1285 10315 1315 10400
rect 1485 10315 1515 10400
rect 1685 10315 1715 10400
rect 1885 10315 1915 10400
rect 2085 10315 2115 10400
rect 2285 10315 2315 10400
rect 2485 10315 2515 10400
rect 2685 10315 2715 10400
rect 2885 10315 2915 10400
rect 3085 10315 3115 10400
rect 3285 10315 3315 10400
rect 3485 10315 3515 10400
rect 3685 10315 3715 10400
rect 3885 10315 3915 10400
rect 4085 10315 4115 10400
rect 4285 10315 4315 10400
rect 4485 10315 4515 10400
rect 4685 10315 4715 10400
rect 4885 10315 4915 10400
rect 5085 10315 5115 10400
rect 5285 10315 5315 10400
rect 5485 10315 5515 10400
rect 5685 10315 5715 10400
rect 5885 10315 5915 10400
rect 6085 10315 6115 10400
rect 6285 10315 6315 10400
rect 6485 10315 6515 10400
rect -150 10305 -50 10315
rect -150 10225 -140 10305
rect -60 10225 -50 10305
rect -150 10215 -50 10225
rect 50 10305 150 10315
rect 50 10225 60 10305
rect 140 10225 150 10305
rect 50 10215 150 10225
rect 250 10305 350 10315
rect 250 10225 260 10305
rect 340 10225 350 10305
rect 250 10215 350 10225
rect 450 10305 550 10315
rect 450 10225 460 10305
rect 540 10225 550 10305
rect 450 10215 550 10225
rect 650 10305 750 10315
rect 650 10225 660 10305
rect 740 10225 750 10305
rect 650 10215 750 10225
rect 850 10305 950 10315
rect 850 10225 860 10305
rect 940 10225 950 10305
rect 850 10215 950 10225
rect 1050 10305 1150 10315
rect 1050 10225 1060 10305
rect 1140 10225 1150 10305
rect 1050 10215 1150 10225
rect 1250 10305 1350 10315
rect 1250 10225 1260 10305
rect 1340 10225 1350 10305
rect 1250 10215 1350 10225
rect 1450 10305 1550 10315
rect 1450 10225 1460 10305
rect 1540 10225 1550 10305
rect 1450 10215 1550 10225
rect 1650 10305 1750 10315
rect 1650 10225 1660 10305
rect 1740 10225 1750 10305
rect 1650 10215 1750 10225
rect 1850 10305 1950 10315
rect 1850 10225 1860 10305
rect 1940 10225 1950 10305
rect 1850 10215 1950 10225
rect 2050 10305 2150 10315
rect 2050 10225 2060 10305
rect 2140 10225 2150 10305
rect 2050 10215 2150 10225
rect 2250 10305 2350 10315
rect 2250 10225 2260 10305
rect 2340 10225 2350 10305
rect 2250 10215 2350 10225
rect 2450 10305 2550 10315
rect 2450 10225 2460 10305
rect 2540 10225 2550 10305
rect 2450 10215 2550 10225
rect 2650 10305 2750 10315
rect 2650 10225 2660 10305
rect 2740 10225 2750 10305
rect 2650 10215 2750 10225
rect 2850 10305 2950 10315
rect 2850 10225 2860 10305
rect 2940 10225 2950 10305
rect 2850 10215 2950 10225
rect 3050 10305 3150 10315
rect 3050 10225 3060 10305
rect 3140 10225 3150 10305
rect 3050 10215 3150 10225
rect 3250 10305 3350 10315
rect 3250 10225 3260 10305
rect 3340 10225 3350 10305
rect 3250 10215 3350 10225
rect 3450 10305 3550 10315
rect 3450 10225 3460 10305
rect 3540 10225 3550 10305
rect 3450 10215 3550 10225
rect 3650 10305 3750 10315
rect 3650 10225 3660 10305
rect 3740 10225 3750 10305
rect 3650 10215 3750 10225
rect 3850 10305 3950 10315
rect 3850 10225 3860 10305
rect 3940 10225 3950 10305
rect 3850 10215 3950 10225
rect 4050 10305 4150 10315
rect 4050 10225 4060 10305
rect 4140 10225 4150 10305
rect 4050 10215 4150 10225
rect 4250 10305 4350 10315
rect 4250 10225 4260 10305
rect 4340 10225 4350 10305
rect 4250 10215 4350 10225
rect 4450 10305 4550 10315
rect 4450 10225 4460 10305
rect 4540 10225 4550 10305
rect 4450 10215 4550 10225
rect 4650 10305 4750 10315
rect 4650 10225 4660 10305
rect 4740 10225 4750 10305
rect 4650 10215 4750 10225
rect 4850 10305 4950 10315
rect 4850 10225 4860 10305
rect 4940 10225 4950 10305
rect 4850 10215 4950 10225
rect 5050 10305 5150 10315
rect 5050 10225 5060 10305
rect 5140 10225 5150 10305
rect 5050 10215 5150 10225
rect 5250 10305 5350 10315
rect 5250 10225 5260 10305
rect 5340 10225 5350 10305
rect 5250 10215 5350 10225
rect 5450 10305 5550 10315
rect 5450 10225 5460 10305
rect 5540 10225 5550 10305
rect 5450 10215 5550 10225
rect 5650 10305 5750 10315
rect 5650 10225 5660 10305
rect 5740 10225 5750 10305
rect 5650 10215 5750 10225
rect 5850 10305 5950 10315
rect 5850 10225 5860 10305
rect 5940 10225 5950 10305
rect 5850 10215 5950 10225
rect 6050 10305 6150 10315
rect 6050 10225 6060 10305
rect 6140 10225 6150 10305
rect 6050 10215 6150 10225
rect 6250 10305 6350 10315
rect 6250 10225 6260 10305
rect 6340 10225 6350 10305
rect 6250 10215 6350 10225
rect 6450 10305 6550 10315
rect 6450 10225 6460 10305
rect 6540 10225 6550 10305
rect 6450 10215 6550 10225
rect -115 10130 -85 10215
rect 85 10130 115 10215
rect 285 10130 315 10215
rect 485 10130 515 10215
rect 685 10130 715 10215
rect 885 10130 915 10215
rect 1085 10130 1115 10215
rect 1285 10130 1315 10215
rect 1485 10130 1515 10215
rect 1685 10130 1715 10215
rect 1885 10130 1915 10215
rect 2085 10130 2115 10215
rect 2285 10130 2315 10215
rect 2485 10130 2515 10215
rect 2685 10130 2715 10215
rect 2885 10130 2915 10215
rect 3085 10130 3115 10215
rect 3285 10130 3315 10215
rect 3485 10130 3515 10215
rect 3685 10130 3715 10215
rect 3885 10130 3915 10215
rect 4085 10130 4115 10215
rect 4285 10130 4315 10215
rect 4485 10130 4515 10215
rect 4685 10130 4715 10215
rect 4885 10130 4915 10215
rect 5085 10130 5115 10215
rect 5285 10130 5315 10215
rect 5485 10130 5515 10215
rect 5685 10130 5715 10215
rect 5885 10130 5915 10215
rect 6085 10130 6115 10215
rect 6285 10130 6315 10215
rect 6485 10130 6515 10215
rect -150 10120 -50 10130
rect -150 10040 -140 10120
rect -60 10040 -50 10120
rect -150 10030 -50 10040
rect 50 10120 150 10130
rect 50 10040 60 10120
rect 140 10040 150 10120
rect 50 10030 150 10040
rect 250 10120 350 10130
rect 250 10040 260 10120
rect 340 10040 350 10120
rect 250 10030 350 10040
rect 450 10120 550 10130
rect 450 10040 460 10120
rect 540 10040 550 10120
rect 450 10030 550 10040
rect 650 10120 750 10130
rect 650 10040 660 10120
rect 740 10040 750 10120
rect 650 10030 750 10040
rect 850 10120 950 10130
rect 850 10040 860 10120
rect 940 10040 950 10120
rect 850 10030 950 10040
rect 1050 10120 1150 10130
rect 1050 10040 1060 10120
rect 1140 10040 1150 10120
rect 1050 10030 1150 10040
rect 1250 10120 1350 10130
rect 1250 10040 1260 10120
rect 1340 10040 1350 10120
rect 1250 10030 1350 10040
rect 1450 10120 1550 10130
rect 1450 10040 1460 10120
rect 1540 10040 1550 10120
rect 1450 10030 1550 10040
rect 1650 10120 1750 10130
rect 1650 10040 1660 10120
rect 1740 10040 1750 10120
rect 1650 10030 1750 10040
rect 1850 10120 1950 10130
rect 1850 10040 1860 10120
rect 1940 10040 1950 10120
rect 1850 10030 1950 10040
rect 2050 10120 2150 10130
rect 2050 10040 2060 10120
rect 2140 10040 2150 10120
rect 2050 10030 2150 10040
rect 2250 10120 2350 10130
rect 2250 10040 2260 10120
rect 2340 10040 2350 10120
rect 2250 10030 2350 10040
rect 2450 10120 2550 10130
rect 2450 10040 2460 10120
rect 2540 10040 2550 10120
rect 2450 10030 2550 10040
rect 2650 10120 2750 10130
rect 2650 10040 2660 10120
rect 2740 10040 2750 10120
rect 2650 10030 2750 10040
rect 2850 10120 2950 10130
rect 2850 10040 2860 10120
rect 2940 10040 2950 10120
rect 2850 10030 2950 10040
rect 3050 10120 3150 10130
rect 3050 10040 3060 10120
rect 3140 10040 3150 10120
rect 3050 10030 3150 10040
rect 3250 10120 3350 10130
rect 3250 10040 3260 10120
rect 3340 10040 3350 10120
rect 3250 10030 3350 10040
rect 3450 10120 3550 10130
rect 3450 10040 3460 10120
rect 3540 10040 3550 10120
rect 3450 10030 3550 10040
rect 3650 10120 3750 10130
rect 3650 10040 3660 10120
rect 3740 10040 3750 10120
rect 3650 10030 3750 10040
rect 3850 10120 3950 10130
rect 3850 10040 3860 10120
rect 3940 10040 3950 10120
rect 3850 10030 3950 10040
rect 4050 10120 4150 10130
rect 4050 10040 4060 10120
rect 4140 10040 4150 10120
rect 4050 10030 4150 10040
rect 4250 10120 4350 10130
rect 4250 10040 4260 10120
rect 4340 10040 4350 10120
rect 4250 10030 4350 10040
rect 4450 10120 4550 10130
rect 4450 10040 4460 10120
rect 4540 10040 4550 10120
rect 4450 10030 4550 10040
rect 4650 10120 4750 10130
rect 4650 10040 4660 10120
rect 4740 10040 4750 10120
rect 4650 10030 4750 10040
rect 4850 10120 4950 10130
rect 4850 10040 4860 10120
rect 4940 10040 4950 10120
rect 4850 10030 4950 10040
rect 5050 10120 5150 10130
rect 5050 10040 5060 10120
rect 5140 10040 5150 10120
rect 5050 10030 5150 10040
rect 5250 10120 5350 10130
rect 5250 10040 5260 10120
rect 5340 10040 5350 10120
rect 5250 10030 5350 10040
rect 5450 10120 5550 10130
rect 5450 10040 5460 10120
rect 5540 10040 5550 10120
rect 5450 10030 5550 10040
rect 5650 10120 5750 10130
rect 5650 10040 5660 10120
rect 5740 10040 5750 10120
rect 5650 10030 5750 10040
rect 5850 10120 5950 10130
rect 5850 10040 5860 10120
rect 5940 10040 5950 10120
rect 5850 10030 5950 10040
rect 6050 10120 6150 10130
rect 6050 10040 6060 10120
rect 6140 10040 6150 10120
rect 6050 10030 6150 10040
rect 6250 10120 6350 10130
rect 6250 10040 6260 10120
rect 6340 10040 6350 10120
rect 6250 10030 6350 10040
rect 6450 10120 6550 10130
rect 6450 10040 6460 10120
rect 6540 10040 6550 10120
rect 6450 10030 6550 10040
rect -115 9945 -85 10030
rect 85 9945 115 10030
rect 285 9945 315 10030
rect 485 9945 515 10030
rect 685 9945 715 10030
rect 885 9945 915 10030
rect 1085 9945 1115 10030
rect 1285 9945 1315 10030
rect 1485 9945 1515 10030
rect 1685 9945 1715 10030
rect 1885 9945 1915 10030
rect 2085 9945 2115 10030
rect 2285 9945 2315 10030
rect 2485 9945 2515 10030
rect 2685 9945 2715 10030
rect 2885 9945 2915 10030
rect 3085 9945 3115 10030
rect 3285 9945 3315 10030
rect 3485 9945 3515 10030
rect 3685 9945 3715 10030
rect 3885 9945 3915 10030
rect 4085 9945 4115 10030
rect 4285 9945 4315 10030
rect 4485 9945 4515 10030
rect 4685 9945 4715 10030
rect 4885 9945 4915 10030
rect 5085 9945 5115 10030
rect 5285 9945 5315 10030
rect 5485 9945 5515 10030
rect 5685 9945 5715 10030
rect 5885 9945 5915 10030
rect 6085 9945 6115 10030
rect 6285 9945 6315 10030
rect 6485 9945 6515 10030
rect -150 9935 -50 9945
rect -150 9855 -140 9935
rect -60 9855 -50 9935
rect -150 9845 -50 9855
rect 50 9935 150 9945
rect 50 9855 60 9935
rect 140 9855 150 9935
rect 50 9845 150 9855
rect 250 9935 350 9945
rect 250 9855 260 9935
rect 340 9855 350 9935
rect 250 9845 350 9855
rect 450 9935 550 9945
rect 450 9855 460 9935
rect 540 9855 550 9935
rect 450 9845 550 9855
rect 650 9935 750 9945
rect 650 9855 660 9935
rect 740 9855 750 9935
rect 650 9845 750 9855
rect 850 9935 950 9945
rect 850 9855 860 9935
rect 940 9855 950 9935
rect 850 9845 950 9855
rect 1050 9935 1150 9945
rect 1050 9855 1060 9935
rect 1140 9855 1150 9935
rect 1050 9845 1150 9855
rect 1250 9935 1350 9945
rect 1250 9855 1260 9935
rect 1340 9855 1350 9935
rect 1250 9845 1350 9855
rect 1450 9935 1550 9945
rect 1450 9855 1460 9935
rect 1540 9855 1550 9935
rect 1450 9845 1550 9855
rect 1650 9935 1750 9945
rect 1650 9855 1660 9935
rect 1740 9855 1750 9935
rect 1650 9845 1750 9855
rect 1850 9935 1950 9945
rect 1850 9855 1860 9935
rect 1940 9855 1950 9935
rect 1850 9845 1950 9855
rect 2050 9935 2150 9945
rect 2050 9855 2060 9935
rect 2140 9855 2150 9935
rect 2050 9845 2150 9855
rect 2250 9935 2350 9945
rect 2250 9855 2260 9935
rect 2340 9855 2350 9935
rect 2250 9845 2350 9855
rect 2450 9935 2550 9945
rect 2450 9855 2460 9935
rect 2540 9855 2550 9935
rect 2450 9845 2550 9855
rect 2650 9935 2750 9945
rect 2650 9855 2660 9935
rect 2740 9855 2750 9935
rect 2650 9845 2750 9855
rect 2850 9935 2950 9945
rect 2850 9855 2860 9935
rect 2940 9855 2950 9935
rect 2850 9845 2950 9855
rect 3050 9935 3150 9945
rect 3050 9855 3060 9935
rect 3140 9855 3150 9935
rect 3050 9845 3150 9855
rect 3250 9935 3350 9945
rect 3250 9855 3260 9935
rect 3340 9855 3350 9935
rect 3250 9845 3350 9855
rect 3450 9935 3550 9945
rect 3450 9855 3460 9935
rect 3540 9855 3550 9935
rect 3450 9845 3550 9855
rect 3650 9935 3750 9945
rect 3650 9855 3660 9935
rect 3740 9855 3750 9935
rect 3650 9845 3750 9855
rect 3850 9935 3950 9945
rect 3850 9855 3860 9935
rect 3940 9855 3950 9935
rect 3850 9845 3950 9855
rect 4050 9935 4150 9945
rect 4050 9855 4060 9935
rect 4140 9855 4150 9935
rect 4050 9845 4150 9855
rect 4250 9935 4350 9945
rect 4250 9855 4260 9935
rect 4340 9855 4350 9935
rect 4250 9845 4350 9855
rect 4450 9935 4550 9945
rect 4450 9855 4460 9935
rect 4540 9855 4550 9935
rect 4450 9845 4550 9855
rect 4650 9935 4750 9945
rect 4650 9855 4660 9935
rect 4740 9855 4750 9935
rect 4650 9845 4750 9855
rect 4850 9935 4950 9945
rect 4850 9855 4860 9935
rect 4940 9855 4950 9935
rect 4850 9845 4950 9855
rect 5050 9935 5150 9945
rect 5050 9855 5060 9935
rect 5140 9855 5150 9935
rect 5050 9845 5150 9855
rect 5250 9935 5350 9945
rect 5250 9855 5260 9935
rect 5340 9855 5350 9935
rect 5250 9845 5350 9855
rect 5450 9935 5550 9945
rect 5450 9855 5460 9935
rect 5540 9855 5550 9935
rect 5450 9845 5550 9855
rect 5650 9935 5750 9945
rect 5650 9855 5660 9935
rect 5740 9855 5750 9935
rect 5650 9845 5750 9855
rect 5850 9935 5950 9945
rect 5850 9855 5860 9935
rect 5940 9855 5950 9935
rect 5850 9845 5950 9855
rect 6050 9935 6150 9945
rect 6050 9855 6060 9935
rect 6140 9855 6150 9935
rect 6050 9845 6150 9855
rect 6250 9935 6350 9945
rect 6250 9855 6260 9935
rect 6340 9855 6350 9935
rect 6250 9845 6350 9855
rect 6450 9935 6550 9945
rect 6450 9855 6460 9935
rect 6540 9855 6550 9935
rect 6450 9845 6550 9855
rect -115 9760 -85 9845
rect 85 9760 115 9845
rect 285 9760 315 9845
rect 485 9760 515 9845
rect 685 9760 715 9845
rect 885 9760 915 9845
rect 1085 9760 1115 9845
rect 1285 9760 1315 9845
rect 1485 9760 1515 9845
rect 1685 9760 1715 9845
rect 1885 9760 1915 9845
rect 2085 9760 2115 9845
rect 2285 9760 2315 9845
rect 2485 9760 2515 9845
rect 2685 9760 2715 9845
rect 2885 9760 2915 9845
rect 3085 9760 3115 9845
rect 3285 9760 3315 9845
rect 3485 9760 3515 9845
rect 3685 9760 3715 9845
rect 3885 9760 3915 9845
rect 4085 9760 4115 9845
rect 4285 9760 4315 9845
rect 4485 9760 4515 9845
rect 4685 9760 4715 9845
rect 4885 9760 4915 9845
rect 5085 9760 5115 9845
rect 5285 9760 5315 9845
rect 5485 9760 5515 9845
rect 5685 9760 5715 9845
rect 5885 9760 5915 9845
rect 6085 9760 6115 9845
rect 6285 9760 6315 9845
rect 6485 9760 6515 9845
rect -150 9750 -50 9760
rect -150 9670 -140 9750
rect -60 9670 -50 9750
rect -150 9660 -50 9670
rect 50 9750 150 9760
rect 50 9670 60 9750
rect 140 9670 150 9750
rect 50 9660 150 9670
rect 250 9750 350 9760
rect 250 9670 260 9750
rect 340 9670 350 9750
rect 250 9660 350 9670
rect 450 9750 550 9760
rect 450 9670 460 9750
rect 540 9670 550 9750
rect 450 9660 550 9670
rect 650 9750 750 9760
rect 650 9670 660 9750
rect 740 9670 750 9750
rect 650 9660 750 9670
rect 850 9750 950 9760
rect 850 9670 860 9750
rect 940 9670 950 9750
rect 850 9660 950 9670
rect 1050 9750 1150 9760
rect 1050 9670 1060 9750
rect 1140 9670 1150 9750
rect 1050 9660 1150 9670
rect 1250 9750 1350 9760
rect 1250 9670 1260 9750
rect 1340 9670 1350 9750
rect 1250 9660 1350 9670
rect 1450 9750 1550 9760
rect 1450 9670 1460 9750
rect 1540 9670 1550 9750
rect 1450 9660 1550 9670
rect 1650 9750 1750 9760
rect 1650 9670 1660 9750
rect 1740 9670 1750 9750
rect 1650 9660 1750 9670
rect 1850 9750 1950 9760
rect 1850 9670 1860 9750
rect 1940 9670 1950 9750
rect 1850 9660 1950 9670
rect 2050 9750 2150 9760
rect 2050 9670 2060 9750
rect 2140 9670 2150 9750
rect 2050 9660 2150 9670
rect 2250 9750 2350 9760
rect 2250 9670 2260 9750
rect 2340 9670 2350 9750
rect 2250 9660 2350 9670
rect 2450 9750 2550 9760
rect 2450 9670 2460 9750
rect 2540 9670 2550 9750
rect 2450 9660 2550 9670
rect 2650 9750 2750 9760
rect 2650 9670 2660 9750
rect 2740 9670 2750 9750
rect 2650 9660 2750 9670
rect 2850 9750 2950 9760
rect 2850 9670 2860 9750
rect 2940 9670 2950 9750
rect 2850 9660 2950 9670
rect 3050 9750 3150 9760
rect 3050 9670 3060 9750
rect 3140 9670 3150 9750
rect 3050 9660 3150 9670
rect 3250 9750 3350 9760
rect 3250 9670 3260 9750
rect 3340 9670 3350 9750
rect 3250 9660 3350 9670
rect 3450 9750 3550 9760
rect 3450 9670 3460 9750
rect 3540 9670 3550 9750
rect 3450 9660 3550 9670
rect 3650 9750 3750 9760
rect 3650 9670 3660 9750
rect 3740 9670 3750 9750
rect 3650 9660 3750 9670
rect 3850 9750 3950 9760
rect 3850 9670 3860 9750
rect 3940 9670 3950 9750
rect 3850 9660 3950 9670
rect 4050 9750 4150 9760
rect 4050 9670 4060 9750
rect 4140 9670 4150 9750
rect 4050 9660 4150 9670
rect 4250 9750 4350 9760
rect 4250 9670 4260 9750
rect 4340 9670 4350 9750
rect 4250 9660 4350 9670
rect 4450 9750 4550 9760
rect 4450 9670 4460 9750
rect 4540 9670 4550 9750
rect 4450 9660 4550 9670
rect 4650 9750 4750 9760
rect 4650 9670 4660 9750
rect 4740 9670 4750 9750
rect 4650 9660 4750 9670
rect 4850 9750 4950 9760
rect 4850 9670 4860 9750
rect 4940 9670 4950 9750
rect 4850 9660 4950 9670
rect 5050 9750 5150 9760
rect 5050 9670 5060 9750
rect 5140 9670 5150 9750
rect 5050 9660 5150 9670
rect 5250 9750 5350 9760
rect 5250 9670 5260 9750
rect 5340 9670 5350 9750
rect 5250 9660 5350 9670
rect 5450 9750 5550 9760
rect 5450 9670 5460 9750
rect 5540 9670 5550 9750
rect 5450 9660 5550 9670
rect 5650 9750 5750 9760
rect 5650 9670 5660 9750
rect 5740 9670 5750 9750
rect 5650 9660 5750 9670
rect 5850 9750 5950 9760
rect 5850 9670 5860 9750
rect 5940 9670 5950 9750
rect 5850 9660 5950 9670
rect 6050 9750 6150 9760
rect 6050 9670 6060 9750
rect 6140 9670 6150 9750
rect 6050 9660 6150 9670
rect 6250 9750 6350 9760
rect 6250 9670 6260 9750
rect 6340 9670 6350 9750
rect 6250 9660 6350 9670
rect 6450 9750 6550 9760
rect 6450 9670 6460 9750
rect 6540 9670 6550 9750
rect 6450 9660 6550 9670
rect -115 9575 -85 9660
rect 85 9575 115 9660
rect 285 9575 315 9660
rect 485 9575 515 9660
rect 685 9575 715 9660
rect 885 9575 915 9660
rect 1085 9575 1115 9660
rect 1285 9575 1315 9660
rect 1485 9575 1515 9660
rect 1685 9575 1715 9660
rect 1885 9575 1915 9660
rect 2085 9575 2115 9660
rect 2285 9575 2315 9660
rect 2485 9575 2515 9660
rect 2685 9575 2715 9660
rect 2885 9575 2915 9660
rect 3085 9575 3115 9660
rect 3285 9575 3315 9660
rect 3485 9575 3515 9660
rect 3685 9575 3715 9660
rect 3885 9575 3915 9660
rect 4085 9575 4115 9660
rect 4285 9575 4315 9660
rect 4485 9575 4515 9660
rect 4685 9575 4715 9660
rect 4885 9575 4915 9660
rect 5085 9575 5115 9660
rect 5285 9575 5315 9660
rect 5485 9575 5515 9660
rect 5685 9575 5715 9660
rect 5885 9575 5915 9660
rect 6085 9575 6115 9660
rect 6285 9575 6315 9660
rect 6485 9575 6515 9660
rect -150 9565 -50 9575
rect -150 9485 -140 9565
rect -60 9485 -50 9565
rect -150 9475 -50 9485
rect 50 9565 150 9575
rect 50 9485 60 9565
rect 140 9485 150 9565
rect 50 9475 150 9485
rect 250 9565 350 9575
rect 250 9485 260 9565
rect 340 9485 350 9565
rect 250 9475 350 9485
rect 450 9565 550 9575
rect 450 9485 460 9565
rect 540 9485 550 9565
rect 450 9475 550 9485
rect 650 9565 750 9575
rect 650 9485 660 9565
rect 740 9485 750 9565
rect 650 9475 750 9485
rect 850 9565 950 9575
rect 850 9485 860 9565
rect 940 9485 950 9565
rect 850 9475 950 9485
rect 1050 9565 1150 9575
rect 1050 9485 1060 9565
rect 1140 9485 1150 9565
rect 1050 9475 1150 9485
rect 1250 9565 1350 9575
rect 1250 9485 1260 9565
rect 1340 9485 1350 9565
rect 1250 9475 1350 9485
rect 1450 9565 1550 9575
rect 1450 9485 1460 9565
rect 1540 9485 1550 9565
rect 1450 9475 1550 9485
rect 1650 9565 1750 9575
rect 1650 9485 1660 9565
rect 1740 9485 1750 9565
rect 1650 9475 1750 9485
rect 1850 9565 1950 9575
rect 1850 9485 1860 9565
rect 1940 9485 1950 9565
rect 1850 9475 1950 9485
rect 2050 9565 2150 9575
rect 2050 9485 2060 9565
rect 2140 9485 2150 9565
rect 2050 9475 2150 9485
rect 2250 9565 2350 9575
rect 2250 9485 2260 9565
rect 2340 9485 2350 9565
rect 2250 9475 2350 9485
rect 2450 9565 2550 9575
rect 2450 9485 2460 9565
rect 2540 9485 2550 9565
rect 2450 9475 2550 9485
rect 2650 9565 2750 9575
rect 2650 9485 2660 9565
rect 2740 9485 2750 9565
rect 2650 9475 2750 9485
rect 2850 9565 2950 9575
rect 2850 9485 2860 9565
rect 2940 9485 2950 9565
rect 2850 9475 2950 9485
rect 3050 9565 3150 9575
rect 3050 9485 3060 9565
rect 3140 9485 3150 9565
rect 3050 9475 3150 9485
rect 3250 9565 3350 9575
rect 3250 9485 3260 9565
rect 3340 9485 3350 9565
rect 3250 9475 3350 9485
rect 3450 9565 3550 9575
rect 3450 9485 3460 9565
rect 3540 9485 3550 9565
rect 3450 9475 3550 9485
rect 3650 9565 3750 9575
rect 3650 9485 3660 9565
rect 3740 9485 3750 9565
rect 3650 9475 3750 9485
rect 3850 9565 3950 9575
rect 3850 9485 3860 9565
rect 3940 9485 3950 9565
rect 3850 9475 3950 9485
rect 4050 9565 4150 9575
rect 4050 9485 4060 9565
rect 4140 9485 4150 9565
rect 4050 9475 4150 9485
rect 4250 9565 4350 9575
rect 4250 9485 4260 9565
rect 4340 9485 4350 9565
rect 4250 9475 4350 9485
rect 4450 9565 4550 9575
rect 4450 9485 4460 9565
rect 4540 9485 4550 9565
rect 4450 9475 4550 9485
rect 4650 9565 4750 9575
rect 4650 9485 4660 9565
rect 4740 9485 4750 9565
rect 4650 9475 4750 9485
rect 4850 9565 4950 9575
rect 4850 9485 4860 9565
rect 4940 9485 4950 9565
rect 4850 9475 4950 9485
rect 5050 9565 5150 9575
rect 5050 9485 5060 9565
rect 5140 9485 5150 9565
rect 5050 9475 5150 9485
rect 5250 9565 5350 9575
rect 5250 9485 5260 9565
rect 5340 9485 5350 9565
rect 5250 9475 5350 9485
rect 5450 9565 5550 9575
rect 5450 9485 5460 9565
rect 5540 9485 5550 9565
rect 5450 9475 5550 9485
rect 5650 9565 5750 9575
rect 5650 9485 5660 9565
rect 5740 9485 5750 9565
rect 5650 9475 5750 9485
rect 5850 9565 5950 9575
rect 5850 9485 5860 9565
rect 5940 9485 5950 9565
rect 5850 9475 5950 9485
rect 6050 9565 6150 9575
rect 6050 9485 6060 9565
rect 6140 9485 6150 9565
rect 6050 9475 6150 9485
rect 6250 9565 6350 9575
rect 6250 9485 6260 9565
rect 6340 9485 6350 9565
rect 6250 9475 6350 9485
rect 6450 9565 6550 9575
rect 6450 9485 6460 9565
rect 6540 9485 6550 9565
rect 6450 9475 6550 9485
rect -115 9390 -85 9475
rect 85 9390 115 9475
rect 285 9390 315 9475
rect 485 9390 515 9475
rect 685 9390 715 9475
rect 885 9390 915 9475
rect 1085 9390 1115 9475
rect 1285 9390 1315 9475
rect 1485 9390 1515 9475
rect 1685 9390 1715 9475
rect 1885 9390 1915 9475
rect 2085 9390 2115 9475
rect 2285 9390 2315 9475
rect 2485 9390 2515 9475
rect 2685 9390 2715 9475
rect 2885 9390 2915 9475
rect 3085 9390 3115 9475
rect 3285 9390 3315 9475
rect 3485 9390 3515 9475
rect 3685 9390 3715 9475
rect 3885 9390 3915 9475
rect 4085 9390 4115 9475
rect 4285 9390 4315 9475
rect 4485 9390 4515 9475
rect 4685 9390 4715 9475
rect 4885 9390 4915 9475
rect 5085 9390 5115 9475
rect 5285 9390 5315 9475
rect 5485 9390 5515 9475
rect 5685 9390 5715 9475
rect 5885 9390 5915 9475
rect 6085 9390 6115 9475
rect 6285 9390 6315 9475
rect 6485 9390 6515 9475
rect -150 9380 -50 9390
rect -150 9300 -140 9380
rect -60 9300 -50 9380
rect -150 9290 -50 9300
rect 50 9380 150 9390
rect 50 9300 60 9380
rect 140 9300 150 9380
rect 50 9290 150 9300
rect 250 9380 350 9390
rect 250 9300 260 9380
rect 340 9300 350 9380
rect 250 9290 350 9300
rect 450 9380 550 9390
rect 450 9300 460 9380
rect 540 9300 550 9380
rect 450 9290 550 9300
rect 650 9380 750 9390
rect 650 9300 660 9380
rect 740 9300 750 9380
rect 650 9290 750 9300
rect 850 9380 950 9390
rect 850 9300 860 9380
rect 940 9300 950 9380
rect 850 9290 950 9300
rect 1050 9380 1150 9390
rect 1050 9300 1060 9380
rect 1140 9300 1150 9380
rect 1050 9290 1150 9300
rect 1250 9380 1350 9390
rect 1250 9300 1260 9380
rect 1340 9300 1350 9380
rect 1250 9290 1350 9300
rect 1450 9380 1550 9390
rect 1450 9300 1460 9380
rect 1540 9300 1550 9380
rect 1450 9290 1550 9300
rect 1650 9380 1750 9390
rect 1650 9300 1660 9380
rect 1740 9300 1750 9380
rect 1650 9290 1750 9300
rect 1850 9380 1950 9390
rect 1850 9300 1860 9380
rect 1940 9300 1950 9380
rect 1850 9290 1950 9300
rect 2050 9380 2150 9390
rect 2050 9300 2060 9380
rect 2140 9300 2150 9380
rect 2050 9290 2150 9300
rect 2250 9380 2350 9390
rect 2250 9300 2260 9380
rect 2340 9300 2350 9380
rect 2250 9290 2350 9300
rect 2450 9380 2550 9390
rect 2450 9300 2460 9380
rect 2540 9300 2550 9380
rect 2450 9290 2550 9300
rect 2650 9380 2750 9390
rect 2650 9300 2660 9380
rect 2740 9300 2750 9380
rect 2650 9290 2750 9300
rect 2850 9380 2950 9390
rect 2850 9300 2860 9380
rect 2940 9300 2950 9380
rect 2850 9290 2950 9300
rect 3050 9380 3150 9390
rect 3050 9300 3060 9380
rect 3140 9300 3150 9380
rect 3050 9290 3150 9300
rect 3250 9380 3350 9390
rect 3250 9300 3260 9380
rect 3340 9300 3350 9380
rect 3250 9290 3350 9300
rect 3450 9380 3550 9390
rect 3450 9300 3460 9380
rect 3540 9300 3550 9380
rect 3450 9290 3550 9300
rect 3650 9380 3750 9390
rect 3650 9300 3660 9380
rect 3740 9300 3750 9380
rect 3650 9290 3750 9300
rect 3850 9380 3950 9390
rect 3850 9300 3860 9380
rect 3940 9300 3950 9380
rect 3850 9290 3950 9300
rect 4050 9380 4150 9390
rect 4050 9300 4060 9380
rect 4140 9300 4150 9380
rect 4050 9290 4150 9300
rect 4250 9380 4350 9390
rect 4250 9300 4260 9380
rect 4340 9300 4350 9380
rect 4250 9290 4350 9300
rect 4450 9380 4550 9390
rect 4450 9300 4460 9380
rect 4540 9300 4550 9380
rect 4450 9290 4550 9300
rect 4650 9380 4750 9390
rect 4650 9300 4660 9380
rect 4740 9300 4750 9380
rect 4650 9290 4750 9300
rect 4850 9380 4950 9390
rect 4850 9300 4860 9380
rect 4940 9300 4950 9380
rect 4850 9290 4950 9300
rect 5050 9380 5150 9390
rect 5050 9300 5060 9380
rect 5140 9300 5150 9380
rect 5050 9290 5150 9300
rect 5250 9380 5350 9390
rect 5250 9300 5260 9380
rect 5340 9300 5350 9380
rect 5250 9290 5350 9300
rect 5450 9380 5550 9390
rect 5450 9300 5460 9380
rect 5540 9300 5550 9380
rect 5450 9290 5550 9300
rect 5650 9380 5750 9390
rect 5650 9300 5660 9380
rect 5740 9300 5750 9380
rect 5650 9290 5750 9300
rect 5850 9380 5950 9390
rect 5850 9300 5860 9380
rect 5940 9300 5950 9380
rect 5850 9290 5950 9300
rect 6050 9380 6150 9390
rect 6050 9300 6060 9380
rect 6140 9300 6150 9380
rect 6050 9290 6150 9300
rect 6250 9380 6350 9390
rect 6250 9300 6260 9380
rect 6340 9300 6350 9380
rect 6250 9290 6350 9300
rect 6450 9380 6550 9390
rect 6450 9300 6460 9380
rect 6540 9300 6550 9380
rect 6450 9290 6550 9300
rect -115 9205 -85 9290
rect 85 9205 115 9290
rect 285 9205 315 9290
rect 485 9205 515 9290
rect 685 9205 715 9290
rect 885 9205 915 9290
rect 1085 9205 1115 9290
rect 1285 9205 1315 9290
rect 1485 9205 1515 9290
rect 1685 9205 1715 9290
rect 1885 9205 1915 9290
rect 2085 9205 2115 9290
rect 2285 9205 2315 9290
rect 2485 9205 2515 9290
rect 2685 9205 2715 9290
rect 2885 9205 2915 9290
rect 3085 9205 3115 9290
rect 3285 9205 3315 9290
rect 3485 9205 3515 9290
rect 3685 9205 3715 9290
rect 3885 9205 3915 9290
rect 4085 9205 4115 9290
rect 4285 9205 4315 9290
rect 4485 9205 4515 9290
rect 4685 9205 4715 9290
rect 4885 9205 4915 9290
rect 5085 9205 5115 9290
rect 5285 9205 5315 9290
rect 5485 9205 5515 9290
rect 5685 9205 5715 9290
rect 5885 9205 5915 9290
rect 6085 9205 6115 9290
rect 6285 9205 6315 9290
rect 6485 9205 6515 9290
rect -150 9195 -50 9205
rect -150 9115 -140 9195
rect -60 9115 -50 9195
rect -150 9105 -50 9115
rect 50 9195 150 9205
rect 50 9115 60 9195
rect 140 9115 150 9195
rect 50 9105 150 9115
rect 250 9195 350 9205
rect 250 9115 260 9195
rect 340 9115 350 9195
rect 250 9105 350 9115
rect 450 9195 550 9205
rect 450 9115 460 9195
rect 540 9115 550 9195
rect 450 9105 550 9115
rect 650 9195 750 9205
rect 650 9115 660 9195
rect 740 9115 750 9195
rect 650 9105 750 9115
rect 850 9195 950 9205
rect 850 9115 860 9195
rect 940 9115 950 9195
rect 850 9105 950 9115
rect 1050 9195 1150 9205
rect 1050 9115 1060 9195
rect 1140 9115 1150 9195
rect 1050 9105 1150 9115
rect 1250 9195 1350 9205
rect 1250 9115 1260 9195
rect 1340 9115 1350 9195
rect 1250 9105 1350 9115
rect 1450 9195 1550 9205
rect 1450 9115 1460 9195
rect 1540 9115 1550 9195
rect 1450 9105 1550 9115
rect 1650 9195 1750 9205
rect 1650 9115 1660 9195
rect 1740 9115 1750 9195
rect 1650 9105 1750 9115
rect 1850 9195 1950 9205
rect 1850 9115 1860 9195
rect 1940 9115 1950 9195
rect 1850 9105 1950 9115
rect 2050 9195 2150 9205
rect 2050 9115 2060 9195
rect 2140 9115 2150 9195
rect 2050 9105 2150 9115
rect 2250 9195 2350 9205
rect 2250 9115 2260 9195
rect 2340 9115 2350 9195
rect 2250 9105 2350 9115
rect 2450 9195 2550 9205
rect 2450 9115 2460 9195
rect 2540 9115 2550 9195
rect 2450 9105 2550 9115
rect 2650 9195 2750 9205
rect 2650 9115 2660 9195
rect 2740 9115 2750 9195
rect 2650 9105 2750 9115
rect 2850 9195 2950 9205
rect 2850 9115 2860 9195
rect 2940 9115 2950 9195
rect 2850 9105 2950 9115
rect 3050 9195 3150 9205
rect 3050 9115 3060 9195
rect 3140 9115 3150 9195
rect 3050 9105 3150 9115
rect 3250 9195 3350 9205
rect 3250 9115 3260 9195
rect 3340 9115 3350 9195
rect 3250 9105 3350 9115
rect 3450 9195 3550 9205
rect 3450 9115 3460 9195
rect 3540 9115 3550 9195
rect 3450 9105 3550 9115
rect 3650 9195 3750 9205
rect 3650 9115 3660 9195
rect 3740 9115 3750 9195
rect 3650 9105 3750 9115
rect 3850 9195 3950 9205
rect 3850 9115 3860 9195
rect 3940 9115 3950 9195
rect 3850 9105 3950 9115
rect 4050 9195 4150 9205
rect 4050 9115 4060 9195
rect 4140 9115 4150 9195
rect 4050 9105 4150 9115
rect 4250 9195 4350 9205
rect 4250 9115 4260 9195
rect 4340 9115 4350 9195
rect 4250 9105 4350 9115
rect 4450 9195 4550 9205
rect 4450 9115 4460 9195
rect 4540 9115 4550 9195
rect 4450 9105 4550 9115
rect 4650 9195 4750 9205
rect 4650 9115 4660 9195
rect 4740 9115 4750 9195
rect 4650 9105 4750 9115
rect 4850 9195 4950 9205
rect 4850 9115 4860 9195
rect 4940 9115 4950 9195
rect 4850 9105 4950 9115
rect 5050 9195 5150 9205
rect 5050 9115 5060 9195
rect 5140 9115 5150 9195
rect 5050 9105 5150 9115
rect 5250 9195 5350 9205
rect 5250 9115 5260 9195
rect 5340 9115 5350 9195
rect 5250 9105 5350 9115
rect 5450 9195 5550 9205
rect 5450 9115 5460 9195
rect 5540 9115 5550 9195
rect 5450 9105 5550 9115
rect 5650 9195 5750 9205
rect 5650 9115 5660 9195
rect 5740 9115 5750 9195
rect 5650 9105 5750 9115
rect 5850 9195 5950 9205
rect 5850 9115 5860 9195
rect 5940 9115 5950 9195
rect 5850 9105 5950 9115
rect 6050 9195 6150 9205
rect 6050 9115 6060 9195
rect 6140 9115 6150 9195
rect 6050 9105 6150 9115
rect 6250 9195 6350 9205
rect 6250 9115 6260 9195
rect 6340 9115 6350 9195
rect 6250 9105 6350 9115
rect 6450 9195 6550 9205
rect 6450 9115 6460 9195
rect 6540 9115 6550 9195
rect 6450 9105 6550 9115
rect -115 9020 -85 9105
rect 85 9020 115 9105
rect 285 9020 315 9105
rect 485 9020 515 9105
rect 685 9020 715 9105
rect 885 9020 915 9105
rect 1085 9020 1115 9105
rect 1285 9020 1315 9105
rect 1485 9020 1515 9105
rect 1685 9020 1715 9105
rect 1885 9020 1915 9105
rect 2085 9020 2115 9105
rect 2285 9020 2315 9105
rect 2485 9020 2515 9105
rect 2685 9020 2715 9105
rect 2885 9020 2915 9105
rect 3085 9020 3115 9105
rect 3285 9020 3315 9105
rect 3485 9020 3515 9105
rect 3685 9020 3715 9105
rect 3885 9020 3915 9105
rect 4085 9020 4115 9105
rect 4285 9020 4315 9105
rect 4485 9020 4515 9105
rect 4685 9020 4715 9105
rect 4885 9020 4915 9105
rect 5085 9020 5115 9105
rect 5285 9020 5315 9105
rect 5485 9020 5515 9105
rect 5685 9020 5715 9105
rect 5885 9020 5915 9105
rect 6085 9020 6115 9105
rect 6285 9020 6315 9105
rect 6485 9020 6515 9105
rect -150 9010 -50 9020
rect -150 8930 -140 9010
rect -60 8930 -50 9010
rect -150 8920 -50 8930
rect 50 9010 150 9020
rect 50 8930 60 9010
rect 140 8930 150 9010
rect 50 8920 150 8930
rect 250 9010 350 9020
rect 250 8930 260 9010
rect 340 8930 350 9010
rect 250 8920 350 8930
rect 450 9010 550 9020
rect 450 8930 460 9010
rect 540 8930 550 9010
rect 450 8920 550 8930
rect 650 9010 750 9020
rect 650 8930 660 9010
rect 740 8930 750 9010
rect 650 8920 750 8930
rect 850 9010 950 9020
rect 850 8930 860 9010
rect 940 8930 950 9010
rect 850 8920 950 8930
rect 1050 9010 1150 9020
rect 1050 8930 1060 9010
rect 1140 8930 1150 9010
rect 1050 8920 1150 8930
rect 1250 9010 1350 9020
rect 1250 8930 1260 9010
rect 1340 8930 1350 9010
rect 1250 8920 1350 8930
rect 1450 9010 1550 9020
rect 1450 8930 1460 9010
rect 1540 8930 1550 9010
rect 1450 8920 1550 8930
rect 1650 9010 1750 9020
rect 1650 8930 1660 9010
rect 1740 8930 1750 9010
rect 1650 8920 1750 8930
rect 1850 9010 1950 9020
rect 1850 8930 1860 9010
rect 1940 8930 1950 9010
rect 1850 8920 1950 8930
rect 2050 9010 2150 9020
rect 2050 8930 2060 9010
rect 2140 8930 2150 9010
rect 2050 8920 2150 8930
rect 2250 9010 2350 9020
rect 2250 8930 2260 9010
rect 2340 8930 2350 9010
rect 2250 8920 2350 8930
rect 2450 9010 2550 9020
rect 2450 8930 2460 9010
rect 2540 8930 2550 9010
rect 2450 8920 2550 8930
rect 2650 9010 2750 9020
rect 2650 8930 2660 9010
rect 2740 8930 2750 9010
rect 2650 8920 2750 8930
rect 2850 9010 2950 9020
rect 2850 8930 2860 9010
rect 2940 8930 2950 9010
rect 2850 8920 2950 8930
rect 3050 9010 3150 9020
rect 3050 8930 3060 9010
rect 3140 8930 3150 9010
rect 3050 8920 3150 8930
rect 3250 9010 3350 9020
rect 3250 8930 3260 9010
rect 3340 8930 3350 9010
rect 3250 8920 3350 8930
rect 3450 9010 3550 9020
rect 3450 8930 3460 9010
rect 3540 8930 3550 9010
rect 3450 8920 3550 8930
rect 3650 9010 3750 9020
rect 3650 8930 3660 9010
rect 3740 8930 3750 9010
rect 3650 8920 3750 8930
rect 3850 9010 3950 9020
rect 3850 8930 3860 9010
rect 3940 8930 3950 9010
rect 3850 8920 3950 8930
rect 4050 9010 4150 9020
rect 4050 8930 4060 9010
rect 4140 8930 4150 9010
rect 4050 8920 4150 8930
rect 4250 9010 4350 9020
rect 4250 8930 4260 9010
rect 4340 8930 4350 9010
rect 4250 8920 4350 8930
rect 4450 9010 4550 9020
rect 4450 8930 4460 9010
rect 4540 8930 4550 9010
rect 4450 8920 4550 8930
rect 4650 9010 4750 9020
rect 4650 8930 4660 9010
rect 4740 8930 4750 9010
rect 4650 8920 4750 8930
rect 4850 9010 4950 9020
rect 4850 8930 4860 9010
rect 4940 8930 4950 9010
rect 4850 8920 4950 8930
rect 5050 9010 5150 9020
rect 5050 8930 5060 9010
rect 5140 8930 5150 9010
rect 5050 8920 5150 8930
rect 5250 9010 5350 9020
rect 5250 8930 5260 9010
rect 5340 8930 5350 9010
rect 5250 8920 5350 8930
rect 5450 9010 5550 9020
rect 5450 8930 5460 9010
rect 5540 8930 5550 9010
rect 5450 8920 5550 8930
rect 5650 9010 5750 9020
rect 5650 8930 5660 9010
rect 5740 8930 5750 9010
rect 5650 8920 5750 8930
rect 5850 9010 5950 9020
rect 5850 8930 5860 9010
rect 5940 8930 5950 9010
rect 5850 8920 5950 8930
rect 6050 9010 6150 9020
rect 6050 8930 6060 9010
rect 6140 8930 6150 9010
rect 6050 8920 6150 8930
rect 6250 9010 6350 9020
rect 6250 8930 6260 9010
rect 6340 8930 6350 9010
rect 6250 8920 6350 8930
rect 6450 9010 6550 9020
rect 6450 8930 6460 9010
rect 6540 8930 6550 9010
rect 6450 8920 6550 8930
rect -115 8835 -85 8920
rect 85 8835 115 8920
rect 285 8835 315 8920
rect 485 8835 515 8920
rect 685 8835 715 8920
rect 885 8835 915 8920
rect 1085 8835 1115 8920
rect 1285 8835 1315 8920
rect 1485 8835 1515 8920
rect 1685 8835 1715 8920
rect 1885 8835 1915 8920
rect 2085 8835 2115 8920
rect 2285 8835 2315 8920
rect 2485 8835 2515 8920
rect 2685 8835 2715 8920
rect 2885 8835 2915 8920
rect 3085 8835 3115 8920
rect 3285 8835 3315 8920
rect 3485 8835 3515 8920
rect 3685 8835 3715 8920
rect 3885 8835 3915 8920
rect 4085 8835 4115 8920
rect 4285 8835 4315 8920
rect 4485 8835 4515 8920
rect 4685 8835 4715 8920
rect 4885 8835 4915 8920
rect 5085 8835 5115 8920
rect 5285 8835 5315 8920
rect 5485 8835 5515 8920
rect 5685 8835 5715 8920
rect 5885 8835 5915 8920
rect 6085 8835 6115 8920
rect 6285 8835 6315 8920
rect 6485 8835 6515 8920
rect -150 8825 -50 8835
rect -150 8745 -140 8825
rect -60 8745 -50 8825
rect -150 8735 -50 8745
rect 50 8825 150 8835
rect 50 8745 60 8825
rect 140 8745 150 8825
rect 50 8735 150 8745
rect 250 8825 350 8835
rect 250 8745 260 8825
rect 340 8745 350 8825
rect 250 8735 350 8745
rect 450 8825 550 8835
rect 450 8745 460 8825
rect 540 8745 550 8825
rect 450 8735 550 8745
rect 650 8825 750 8835
rect 650 8745 660 8825
rect 740 8745 750 8825
rect 650 8735 750 8745
rect 850 8825 950 8835
rect 850 8745 860 8825
rect 940 8745 950 8825
rect 850 8735 950 8745
rect 1050 8825 1150 8835
rect 1050 8745 1060 8825
rect 1140 8745 1150 8825
rect 1050 8735 1150 8745
rect 1250 8825 1350 8835
rect 1250 8745 1260 8825
rect 1340 8745 1350 8825
rect 1250 8735 1350 8745
rect 1450 8825 1550 8835
rect 1450 8745 1460 8825
rect 1540 8745 1550 8825
rect 1450 8735 1550 8745
rect 1650 8825 1750 8835
rect 1650 8745 1660 8825
rect 1740 8745 1750 8825
rect 1650 8735 1750 8745
rect 1850 8825 1950 8835
rect 1850 8745 1860 8825
rect 1940 8745 1950 8825
rect 1850 8735 1950 8745
rect 2050 8825 2150 8835
rect 2050 8745 2060 8825
rect 2140 8745 2150 8825
rect 2050 8735 2150 8745
rect 2250 8825 2350 8835
rect 2250 8745 2260 8825
rect 2340 8745 2350 8825
rect 2250 8735 2350 8745
rect 2450 8825 2550 8835
rect 2450 8745 2460 8825
rect 2540 8745 2550 8825
rect 2450 8735 2550 8745
rect 2650 8825 2750 8835
rect 2650 8745 2660 8825
rect 2740 8745 2750 8825
rect 2650 8735 2750 8745
rect 2850 8825 2950 8835
rect 2850 8745 2860 8825
rect 2940 8745 2950 8825
rect 2850 8735 2950 8745
rect 3050 8825 3150 8835
rect 3050 8745 3060 8825
rect 3140 8745 3150 8825
rect 3050 8735 3150 8745
rect 3250 8825 3350 8835
rect 3250 8745 3260 8825
rect 3340 8745 3350 8825
rect 3250 8735 3350 8745
rect 3450 8825 3550 8835
rect 3450 8745 3460 8825
rect 3540 8745 3550 8825
rect 3450 8735 3550 8745
rect 3650 8825 3750 8835
rect 3650 8745 3660 8825
rect 3740 8745 3750 8825
rect 3650 8735 3750 8745
rect 3850 8825 3950 8835
rect 3850 8745 3860 8825
rect 3940 8745 3950 8825
rect 3850 8735 3950 8745
rect 4050 8825 4150 8835
rect 4050 8745 4060 8825
rect 4140 8745 4150 8825
rect 4050 8735 4150 8745
rect 4250 8825 4350 8835
rect 4250 8745 4260 8825
rect 4340 8745 4350 8825
rect 4250 8735 4350 8745
rect 4450 8825 4550 8835
rect 4450 8745 4460 8825
rect 4540 8745 4550 8825
rect 4450 8735 4550 8745
rect 4650 8825 4750 8835
rect 4650 8745 4660 8825
rect 4740 8745 4750 8825
rect 4650 8735 4750 8745
rect 4850 8825 4950 8835
rect 4850 8745 4860 8825
rect 4940 8745 4950 8825
rect 4850 8735 4950 8745
rect 5050 8825 5150 8835
rect 5050 8745 5060 8825
rect 5140 8745 5150 8825
rect 5050 8735 5150 8745
rect 5250 8825 5350 8835
rect 5250 8745 5260 8825
rect 5340 8745 5350 8825
rect 5250 8735 5350 8745
rect 5450 8825 5550 8835
rect 5450 8745 5460 8825
rect 5540 8745 5550 8825
rect 5450 8735 5550 8745
rect 5650 8825 5750 8835
rect 5650 8745 5660 8825
rect 5740 8745 5750 8825
rect 5650 8735 5750 8745
rect 5850 8825 5950 8835
rect 5850 8745 5860 8825
rect 5940 8745 5950 8825
rect 5850 8735 5950 8745
rect 6050 8825 6150 8835
rect 6050 8745 6060 8825
rect 6140 8745 6150 8825
rect 6050 8735 6150 8745
rect 6250 8825 6350 8835
rect 6250 8745 6260 8825
rect 6340 8745 6350 8825
rect 6250 8735 6350 8745
rect 6450 8825 6550 8835
rect 6450 8745 6460 8825
rect 6540 8745 6550 8825
rect 6450 8735 6550 8745
rect -115 8650 -85 8735
rect 85 8650 115 8735
rect 285 8650 315 8735
rect 485 8650 515 8735
rect 685 8650 715 8735
rect 885 8650 915 8735
rect 1085 8650 1115 8735
rect 1285 8650 1315 8735
rect 1485 8650 1515 8735
rect 1685 8650 1715 8735
rect 1885 8650 1915 8735
rect 2085 8650 2115 8735
rect 2285 8650 2315 8735
rect 2485 8650 2515 8735
rect 2685 8650 2715 8735
rect 2885 8650 2915 8735
rect 3085 8650 3115 8735
rect 3285 8650 3315 8735
rect 3485 8650 3515 8735
rect 3685 8650 3715 8735
rect 3885 8650 3915 8735
rect 4085 8650 4115 8735
rect 4285 8650 4315 8735
rect 4485 8650 4515 8735
rect 4685 8650 4715 8735
rect 4885 8650 4915 8735
rect 5085 8650 5115 8735
rect 5285 8650 5315 8735
rect 5485 8650 5515 8735
rect 5685 8650 5715 8735
rect 5885 8650 5915 8735
rect 6085 8650 6115 8735
rect 6285 8650 6315 8735
rect 6485 8650 6515 8735
rect -150 8640 -50 8650
rect -150 8560 -140 8640
rect -60 8560 -50 8640
rect -150 8550 -50 8560
rect 50 8640 150 8650
rect 50 8560 60 8640
rect 140 8560 150 8640
rect 50 8550 150 8560
rect 250 8640 350 8650
rect 250 8560 260 8640
rect 340 8560 350 8640
rect 250 8550 350 8560
rect 450 8640 550 8650
rect 450 8560 460 8640
rect 540 8560 550 8640
rect 450 8550 550 8560
rect 650 8640 750 8650
rect 650 8560 660 8640
rect 740 8560 750 8640
rect 650 8550 750 8560
rect 850 8640 950 8650
rect 850 8560 860 8640
rect 940 8560 950 8640
rect 850 8550 950 8560
rect 1050 8640 1150 8650
rect 1050 8560 1060 8640
rect 1140 8560 1150 8640
rect 1050 8550 1150 8560
rect 1250 8640 1350 8650
rect 1250 8560 1260 8640
rect 1340 8560 1350 8640
rect 1250 8550 1350 8560
rect 1450 8640 1550 8650
rect 1450 8560 1460 8640
rect 1540 8560 1550 8640
rect 1450 8550 1550 8560
rect 1650 8640 1750 8650
rect 1650 8560 1660 8640
rect 1740 8560 1750 8640
rect 1650 8550 1750 8560
rect 1850 8640 1950 8650
rect 1850 8560 1860 8640
rect 1940 8560 1950 8640
rect 1850 8550 1950 8560
rect 2050 8640 2150 8650
rect 2050 8560 2060 8640
rect 2140 8560 2150 8640
rect 2050 8550 2150 8560
rect 2250 8640 2350 8650
rect 2250 8560 2260 8640
rect 2340 8560 2350 8640
rect 2250 8550 2350 8560
rect 2450 8640 2550 8650
rect 2450 8560 2460 8640
rect 2540 8560 2550 8640
rect 2450 8550 2550 8560
rect 2650 8640 2750 8650
rect 2650 8560 2660 8640
rect 2740 8560 2750 8640
rect 2650 8550 2750 8560
rect 2850 8640 2950 8650
rect 2850 8560 2860 8640
rect 2940 8560 2950 8640
rect 2850 8550 2950 8560
rect 3050 8640 3150 8650
rect 3050 8560 3060 8640
rect 3140 8560 3150 8640
rect 3050 8550 3150 8560
rect 3250 8640 3350 8650
rect 3250 8560 3260 8640
rect 3340 8560 3350 8640
rect 3250 8550 3350 8560
rect 3450 8640 3550 8650
rect 3450 8560 3460 8640
rect 3540 8560 3550 8640
rect 3450 8550 3550 8560
rect 3650 8640 3750 8650
rect 3650 8560 3660 8640
rect 3740 8560 3750 8640
rect 3650 8550 3750 8560
rect 3850 8640 3950 8650
rect 3850 8560 3860 8640
rect 3940 8560 3950 8640
rect 3850 8550 3950 8560
rect 4050 8640 4150 8650
rect 4050 8560 4060 8640
rect 4140 8560 4150 8640
rect 4050 8550 4150 8560
rect 4250 8640 4350 8650
rect 4250 8560 4260 8640
rect 4340 8560 4350 8640
rect 4250 8550 4350 8560
rect 4450 8640 4550 8650
rect 4450 8560 4460 8640
rect 4540 8560 4550 8640
rect 4450 8550 4550 8560
rect 4650 8640 4750 8650
rect 4650 8560 4660 8640
rect 4740 8560 4750 8640
rect 4650 8550 4750 8560
rect 4850 8640 4950 8650
rect 4850 8560 4860 8640
rect 4940 8560 4950 8640
rect 4850 8550 4950 8560
rect 5050 8640 5150 8650
rect 5050 8560 5060 8640
rect 5140 8560 5150 8640
rect 5050 8550 5150 8560
rect 5250 8640 5350 8650
rect 5250 8560 5260 8640
rect 5340 8560 5350 8640
rect 5250 8550 5350 8560
rect 5450 8640 5550 8650
rect 5450 8560 5460 8640
rect 5540 8560 5550 8640
rect 5450 8550 5550 8560
rect 5650 8640 5750 8650
rect 5650 8560 5660 8640
rect 5740 8560 5750 8640
rect 5650 8550 5750 8560
rect 5850 8640 5950 8650
rect 5850 8560 5860 8640
rect 5940 8560 5950 8640
rect 5850 8550 5950 8560
rect 6050 8640 6150 8650
rect 6050 8560 6060 8640
rect 6140 8560 6150 8640
rect 6050 8550 6150 8560
rect 6250 8640 6350 8650
rect 6250 8560 6260 8640
rect 6340 8560 6350 8640
rect 6250 8550 6350 8560
rect 6450 8640 6550 8650
rect 6450 8560 6460 8640
rect 6540 8560 6550 8640
rect 6450 8550 6550 8560
rect -115 8465 -85 8550
rect 85 8465 115 8550
rect 285 8465 315 8550
rect 485 8465 515 8550
rect 685 8465 715 8550
rect 885 8465 915 8550
rect 1085 8465 1115 8550
rect 1285 8465 1315 8550
rect 1485 8465 1515 8550
rect 1685 8465 1715 8550
rect 1885 8465 1915 8550
rect 2085 8465 2115 8550
rect 2285 8465 2315 8550
rect 2485 8465 2515 8550
rect 2685 8465 2715 8550
rect 2885 8465 2915 8550
rect 3085 8465 3115 8550
rect 3285 8465 3315 8550
rect 3485 8465 3515 8550
rect 3685 8465 3715 8550
rect 3885 8465 3915 8550
rect 4085 8465 4115 8550
rect 4285 8465 4315 8550
rect 4485 8465 4515 8550
rect 4685 8465 4715 8550
rect 4885 8465 4915 8550
rect 5085 8465 5115 8550
rect 5285 8465 5315 8550
rect 5485 8465 5515 8550
rect 5685 8465 5715 8550
rect 5885 8465 5915 8550
rect 6085 8465 6115 8550
rect 6285 8465 6315 8550
rect 6485 8465 6515 8550
rect -150 8455 -50 8465
rect -150 8375 -140 8455
rect -60 8375 -50 8455
rect -150 8365 -50 8375
rect 50 8455 150 8465
rect 50 8375 60 8455
rect 140 8375 150 8455
rect 50 8365 150 8375
rect 250 8455 350 8465
rect 250 8375 260 8455
rect 340 8375 350 8455
rect 250 8365 350 8375
rect 450 8455 550 8465
rect 450 8375 460 8455
rect 540 8375 550 8455
rect 450 8365 550 8375
rect 650 8455 750 8465
rect 650 8375 660 8455
rect 740 8375 750 8455
rect 650 8365 750 8375
rect 850 8455 950 8465
rect 850 8375 860 8455
rect 940 8375 950 8455
rect 850 8365 950 8375
rect 1050 8455 1150 8465
rect 1050 8375 1060 8455
rect 1140 8375 1150 8455
rect 1050 8365 1150 8375
rect 1250 8455 1350 8465
rect 1250 8375 1260 8455
rect 1340 8375 1350 8455
rect 1250 8365 1350 8375
rect 1450 8455 1550 8465
rect 1450 8375 1460 8455
rect 1540 8375 1550 8455
rect 1450 8365 1550 8375
rect 1650 8455 1750 8465
rect 1650 8375 1660 8455
rect 1740 8375 1750 8455
rect 1650 8365 1750 8375
rect 1850 8455 1950 8465
rect 1850 8375 1860 8455
rect 1940 8375 1950 8455
rect 1850 8365 1950 8375
rect 2050 8455 2150 8465
rect 2050 8375 2060 8455
rect 2140 8375 2150 8455
rect 2050 8365 2150 8375
rect 2250 8455 2350 8465
rect 2250 8375 2260 8455
rect 2340 8375 2350 8455
rect 2250 8365 2350 8375
rect 2450 8455 2550 8465
rect 2450 8375 2460 8455
rect 2540 8375 2550 8455
rect 2450 8365 2550 8375
rect 2650 8455 2750 8465
rect 2650 8375 2660 8455
rect 2740 8375 2750 8455
rect 2650 8365 2750 8375
rect 2850 8455 2950 8465
rect 2850 8375 2860 8455
rect 2940 8375 2950 8455
rect 2850 8365 2950 8375
rect 3050 8455 3150 8465
rect 3050 8375 3060 8455
rect 3140 8375 3150 8455
rect 3050 8365 3150 8375
rect 3250 8455 3350 8465
rect 3250 8375 3260 8455
rect 3340 8375 3350 8455
rect 3250 8365 3350 8375
rect 3450 8455 3550 8465
rect 3450 8375 3460 8455
rect 3540 8375 3550 8455
rect 3450 8365 3550 8375
rect 3650 8455 3750 8465
rect 3650 8375 3660 8455
rect 3740 8375 3750 8455
rect 3650 8365 3750 8375
rect 3850 8455 3950 8465
rect 3850 8375 3860 8455
rect 3940 8375 3950 8455
rect 3850 8365 3950 8375
rect 4050 8455 4150 8465
rect 4050 8375 4060 8455
rect 4140 8375 4150 8455
rect 4050 8365 4150 8375
rect 4250 8455 4350 8465
rect 4250 8375 4260 8455
rect 4340 8375 4350 8455
rect 4250 8365 4350 8375
rect 4450 8455 4550 8465
rect 4450 8375 4460 8455
rect 4540 8375 4550 8455
rect 4450 8365 4550 8375
rect 4650 8455 4750 8465
rect 4650 8375 4660 8455
rect 4740 8375 4750 8455
rect 4650 8365 4750 8375
rect 4850 8455 4950 8465
rect 4850 8375 4860 8455
rect 4940 8375 4950 8455
rect 4850 8365 4950 8375
rect 5050 8455 5150 8465
rect 5050 8375 5060 8455
rect 5140 8375 5150 8455
rect 5050 8365 5150 8375
rect 5250 8455 5350 8465
rect 5250 8375 5260 8455
rect 5340 8375 5350 8455
rect 5250 8365 5350 8375
rect 5450 8455 5550 8465
rect 5450 8375 5460 8455
rect 5540 8375 5550 8455
rect 5450 8365 5550 8375
rect 5650 8455 5750 8465
rect 5650 8375 5660 8455
rect 5740 8375 5750 8455
rect 5650 8365 5750 8375
rect 5850 8455 5950 8465
rect 5850 8375 5860 8455
rect 5940 8375 5950 8455
rect 5850 8365 5950 8375
rect 6050 8455 6150 8465
rect 6050 8375 6060 8455
rect 6140 8375 6150 8455
rect 6050 8365 6150 8375
rect 6250 8455 6350 8465
rect 6250 8375 6260 8455
rect 6340 8375 6350 8455
rect 6250 8365 6350 8375
rect 6450 8455 6550 8465
rect 6450 8375 6460 8455
rect 6540 8375 6550 8455
rect 6450 8365 6550 8375
rect -115 8280 -85 8365
rect 85 8280 115 8365
rect 285 8280 315 8365
rect 485 8280 515 8365
rect 685 8280 715 8365
rect 885 8280 915 8365
rect 1085 8280 1115 8365
rect 1285 8280 1315 8365
rect 1485 8280 1515 8365
rect 1685 8280 1715 8365
rect 1885 8280 1915 8365
rect 2085 8280 2115 8365
rect 2285 8280 2315 8365
rect 2485 8280 2515 8365
rect 2685 8280 2715 8365
rect 2885 8280 2915 8365
rect 3085 8280 3115 8365
rect 3285 8280 3315 8365
rect 3485 8280 3515 8365
rect 3685 8280 3715 8365
rect 3885 8280 3915 8365
rect 4085 8280 4115 8365
rect 4285 8280 4315 8365
rect 4485 8280 4515 8365
rect 4685 8280 4715 8365
rect 4885 8280 4915 8365
rect 5085 8280 5115 8365
rect 5285 8280 5315 8365
rect 5485 8280 5515 8365
rect 5685 8280 5715 8365
rect 5885 8280 5915 8365
rect 6085 8280 6115 8365
rect 6285 8280 6315 8365
rect 6485 8280 6515 8365
rect -150 8270 -50 8280
rect -150 8190 -140 8270
rect -60 8190 -50 8270
rect -150 8180 -50 8190
rect 50 8270 150 8280
rect 50 8190 60 8270
rect 140 8190 150 8270
rect 50 8180 150 8190
rect 250 8270 350 8280
rect 250 8190 260 8270
rect 340 8190 350 8270
rect 250 8180 350 8190
rect 450 8270 550 8280
rect 450 8190 460 8270
rect 540 8190 550 8270
rect 450 8180 550 8190
rect 650 8270 750 8280
rect 650 8190 660 8270
rect 740 8190 750 8270
rect 650 8180 750 8190
rect 850 8270 950 8280
rect 850 8190 860 8270
rect 940 8190 950 8270
rect 850 8180 950 8190
rect 1050 8270 1150 8280
rect 1050 8190 1060 8270
rect 1140 8190 1150 8270
rect 1050 8180 1150 8190
rect 1250 8270 1350 8280
rect 1250 8190 1260 8270
rect 1340 8190 1350 8270
rect 1250 8180 1350 8190
rect 1450 8270 1550 8280
rect 1450 8190 1460 8270
rect 1540 8190 1550 8270
rect 1450 8180 1550 8190
rect 1650 8270 1750 8280
rect 1650 8190 1660 8270
rect 1740 8190 1750 8270
rect 1650 8180 1750 8190
rect 1850 8270 1950 8280
rect 1850 8190 1860 8270
rect 1940 8190 1950 8270
rect 1850 8180 1950 8190
rect 2050 8270 2150 8280
rect 2050 8190 2060 8270
rect 2140 8190 2150 8270
rect 2050 8180 2150 8190
rect 2250 8270 2350 8280
rect 2250 8190 2260 8270
rect 2340 8190 2350 8270
rect 2250 8180 2350 8190
rect 2450 8270 2550 8280
rect 2450 8190 2460 8270
rect 2540 8190 2550 8270
rect 2450 8180 2550 8190
rect 2650 8270 2750 8280
rect 2650 8190 2660 8270
rect 2740 8190 2750 8270
rect 2650 8180 2750 8190
rect 2850 8270 2950 8280
rect 2850 8190 2860 8270
rect 2940 8190 2950 8270
rect 2850 8180 2950 8190
rect 3050 8270 3150 8280
rect 3050 8190 3060 8270
rect 3140 8190 3150 8270
rect 3050 8180 3150 8190
rect 3250 8270 3350 8280
rect 3250 8190 3260 8270
rect 3340 8190 3350 8270
rect 3250 8180 3350 8190
rect 3450 8270 3550 8280
rect 3450 8190 3460 8270
rect 3540 8190 3550 8270
rect 3450 8180 3550 8190
rect 3650 8270 3750 8280
rect 3650 8190 3660 8270
rect 3740 8190 3750 8270
rect 3650 8180 3750 8190
rect 3850 8270 3950 8280
rect 3850 8190 3860 8270
rect 3940 8190 3950 8270
rect 3850 8180 3950 8190
rect 4050 8270 4150 8280
rect 4050 8190 4060 8270
rect 4140 8190 4150 8270
rect 4050 8180 4150 8190
rect 4250 8270 4350 8280
rect 4250 8190 4260 8270
rect 4340 8190 4350 8270
rect 4250 8180 4350 8190
rect 4450 8270 4550 8280
rect 4450 8190 4460 8270
rect 4540 8190 4550 8270
rect 4450 8180 4550 8190
rect 4650 8270 4750 8280
rect 4650 8190 4660 8270
rect 4740 8190 4750 8270
rect 4650 8180 4750 8190
rect 4850 8270 4950 8280
rect 4850 8190 4860 8270
rect 4940 8190 4950 8270
rect 4850 8180 4950 8190
rect 5050 8270 5150 8280
rect 5050 8190 5060 8270
rect 5140 8190 5150 8270
rect 5050 8180 5150 8190
rect 5250 8270 5350 8280
rect 5250 8190 5260 8270
rect 5340 8190 5350 8270
rect 5250 8180 5350 8190
rect 5450 8270 5550 8280
rect 5450 8190 5460 8270
rect 5540 8190 5550 8270
rect 5450 8180 5550 8190
rect 5650 8270 5750 8280
rect 5650 8190 5660 8270
rect 5740 8190 5750 8270
rect 5650 8180 5750 8190
rect 5850 8270 5950 8280
rect 5850 8190 5860 8270
rect 5940 8190 5950 8270
rect 5850 8180 5950 8190
rect 6050 8270 6150 8280
rect 6050 8190 6060 8270
rect 6140 8190 6150 8270
rect 6050 8180 6150 8190
rect 6250 8270 6350 8280
rect 6250 8190 6260 8270
rect 6340 8190 6350 8270
rect 6250 8180 6350 8190
rect 6450 8270 6550 8280
rect 6450 8190 6460 8270
rect 6540 8190 6550 8270
rect 6450 8180 6550 8190
rect -115 8095 -85 8180
rect 85 8095 115 8180
rect 285 8095 315 8180
rect 485 8095 515 8180
rect 685 8095 715 8180
rect 885 8095 915 8180
rect 1085 8095 1115 8180
rect 1285 8095 1315 8180
rect 1485 8095 1515 8180
rect 1685 8095 1715 8180
rect 1885 8095 1915 8180
rect 2085 8095 2115 8180
rect 2285 8095 2315 8180
rect 2485 8095 2515 8180
rect 2685 8095 2715 8180
rect 2885 8095 2915 8180
rect 3085 8095 3115 8180
rect 3285 8095 3315 8180
rect 3485 8095 3515 8180
rect 3685 8095 3715 8180
rect 3885 8095 3915 8180
rect 4085 8095 4115 8180
rect 4285 8095 4315 8180
rect 4485 8095 4515 8180
rect 4685 8095 4715 8180
rect 4885 8095 4915 8180
rect 5085 8095 5115 8180
rect 5285 8095 5315 8180
rect 5485 8095 5515 8180
rect 5685 8095 5715 8180
rect 5885 8095 5915 8180
rect 6085 8095 6115 8180
rect 6285 8095 6315 8180
rect 6485 8095 6515 8180
rect -150 8085 -50 8095
rect -150 8005 -140 8085
rect -60 8005 -50 8085
rect -150 7995 -50 8005
rect 50 8085 150 8095
rect 50 8005 60 8085
rect 140 8005 150 8085
rect 50 7995 150 8005
rect 250 8085 350 8095
rect 250 8005 260 8085
rect 340 8005 350 8085
rect 250 7995 350 8005
rect 450 8085 550 8095
rect 450 8005 460 8085
rect 540 8005 550 8085
rect 450 7995 550 8005
rect 650 8085 750 8095
rect 650 8005 660 8085
rect 740 8005 750 8085
rect 650 7995 750 8005
rect 850 8085 950 8095
rect 850 8005 860 8085
rect 940 8005 950 8085
rect 850 7995 950 8005
rect 1050 8085 1150 8095
rect 1050 8005 1060 8085
rect 1140 8005 1150 8085
rect 1050 7995 1150 8005
rect 1250 8085 1350 8095
rect 1250 8005 1260 8085
rect 1340 8005 1350 8085
rect 1250 7995 1350 8005
rect 1450 8085 1550 8095
rect 1450 8005 1460 8085
rect 1540 8005 1550 8085
rect 1450 7995 1550 8005
rect 1650 8085 1750 8095
rect 1650 8005 1660 8085
rect 1740 8005 1750 8085
rect 1650 7995 1750 8005
rect 1850 8085 1950 8095
rect 1850 8005 1860 8085
rect 1940 8005 1950 8085
rect 1850 7995 1950 8005
rect 2050 8085 2150 8095
rect 2050 8005 2060 8085
rect 2140 8005 2150 8085
rect 2050 7995 2150 8005
rect 2250 8085 2350 8095
rect 2250 8005 2260 8085
rect 2340 8005 2350 8085
rect 2250 7995 2350 8005
rect 2450 8085 2550 8095
rect 2450 8005 2460 8085
rect 2540 8005 2550 8085
rect 2450 7995 2550 8005
rect 2650 8085 2750 8095
rect 2650 8005 2660 8085
rect 2740 8005 2750 8085
rect 2650 7995 2750 8005
rect 2850 8085 2950 8095
rect 2850 8005 2860 8085
rect 2940 8005 2950 8085
rect 2850 7995 2950 8005
rect 3050 8085 3150 8095
rect 3050 8005 3060 8085
rect 3140 8005 3150 8085
rect 3050 7995 3150 8005
rect 3250 8085 3350 8095
rect 3250 8005 3260 8085
rect 3340 8005 3350 8085
rect 3250 7995 3350 8005
rect 3450 8085 3550 8095
rect 3450 8005 3460 8085
rect 3540 8005 3550 8085
rect 3450 7995 3550 8005
rect 3650 8085 3750 8095
rect 3650 8005 3660 8085
rect 3740 8005 3750 8085
rect 3650 7995 3750 8005
rect 3850 8085 3950 8095
rect 3850 8005 3860 8085
rect 3940 8005 3950 8085
rect 3850 7995 3950 8005
rect 4050 8085 4150 8095
rect 4050 8005 4060 8085
rect 4140 8005 4150 8085
rect 4050 7995 4150 8005
rect 4250 8085 4350 8095
rect 4250 8005 4260 8085
rect 4340 8005 4350 8085
rect 4250 7995 4350 8005
rect 4450 8085 4550 8095
rect 4450 8005 4460 8085
rect 4540 8005 4550 8085
rect 4450 7995 4550 8005
rect 4650 8085 4750 8095
rect 4650 8005 4660 8085
rect 4740 8005 4750 8085
rect 4650 7995 4750 8005
rect 4850 8085 4950 8095
rect 4850 8005 4860 8085
rect 4940 8005 4950 8085
rect 4850 7995 4950 8005
rect 5050 8085 5150 8095
rect 5050 8005 5060 8085
rect 5140 8005 5150 8085
rect 5050 7995 5150 8005
rect 5250 8085 5350 8095
rect 5250 8005 5260 8085
rect 5340 8005 5350 8085
rect 5250 7995 5350 8005
rect 5450 8085 5550 8095
rect 5450 8005 5460 8085
rect 5540 8005 5550 8085
rect 5450 7995 5550 8005
rect 5650 8085 5750 8095
rect 5650 8005 5660 8085
rect 5740 8005 5750 8085
rect 5650 7995 5750 8005
rect 5850 8085 5950 8095
rect 5850 8005 5860 8085
rect 5940 8005 5950 8085
rect 5850 7995 5950 8005
rect 6050 8085 6150 8095
rect 6050 8005 6060 8085
rect 6140 8005 6150 8085
rect 6050 7995 6150 8005
rect 6250 8085 6350 8095
rect 6250 8005 6260 8085
rect 6340 8005 6350 8085
rect 6250 7995 6350 8005
rect 6450 8085 6550 8095
rect 6450 8005 6460 8085
rect 6540 8005 6550 8085
rect 6450 7995 6550 8005
rect -115 7910 -85 7995
rect 85 7910 115 7995
rect 285 7910 315 7995
rect 485 7910 515 7995
rect 685 7910 715 7995
rect 885 7910 915 7995
rect 1085 7910 1115 7995
rect 1285 7910 1315 7995
rect 1485 7910 1515 7995
rect 1685 7910 1715 7995
rect 1885 7910 1915 7995
rect 2085 7910 2115 7995
rect 2285 7910 2315 7995
rect 2485 7910 2515 7995
rect 2685 7910 2715 7995
rect 2885 7910 2915 7995
rect 3085 7910 3115 7995
rect 3285 7910 3315 7995
rect 3485 7910 3515 7995
rect 3685 7910 3715 7995
rect 3885 7910 3915 7995
rect 4085 7910 4115 7995
rect 4285 7910 4315 7995
rect 4485 7910 4515 7995
rect 4685 7910 4715 7995
rect 4885 7910 4915 7995
rect 5085 7910 5115 7995
rect 5285 7910 5315 7995
rect 5485 7910 5515 7995
rect 5685 7910 5715 7995
rect 5885 7910 5915 7995
rect 6085 7910 6115 7995
rect 6285 7910 6315 7995
rect 6485 7910 6515 7995
rect -150 7900 -50 7910
rect -150 7820 -140 7900
rect -60 7820 -50 7900
rect -150 7810 -50 7820
rect 50 7900 150 7910
rect 50 7820 60 7900
rect 140 7820 150 7900
rect 50 7810 150 7820
rect 250 7900 350 7910
rect 250 7820 260 7900
rect 340 7820 350 7900
rect 250 7810 350 7820
rect 450 7900 550 7910
rect 450 7820 460 7900
rect 540 7820 550 7900
rect 450 7810 550 7820
rect 650 7900 750 7910
rect 650 7820 660 7900
rect 740 7820 750 7900
rect 650 7810 750 7820
rect 850 7900 950 7910
rect 850 7820 860 7900
rect 940 7820 950 7900
rect 850 7810 950 7820
rect 1050 7900 1150 7910
rect 1050 7820 1060 7900
rect 1140 7820 1150 7900
rect 1050 7810 1150 7820
rect 1250 7900 1350 7910
rect 1250 7820 1260 7900
rect 1340 7820 1350 7900
rect 1250 7810 1350 7820
rect 1450 7900 1550 7910
rect 1450 7820 1460 7900
rect 1540 7820 1550 7900
rect 1450 7810 1550 7820
rect 1650 7900 1750 7910
rect 1650 7820 1660 7900
rect 1740 7820 1750 7900
rect 1650 7810 1750 7820
rect 1850 7900 1950 7910
rect 1850 7820 1860 7900
rect 1940 7820 1950 7900
rect 1850 7810 1950 7820
rect 2050 7900 2150 7910
rect 2050 7820 2060 7900
rect 2140 7820 2150 7900
rect 2050 7810 2150 7820
rect 2250 7900 2350 7910
rect 2250 7820 2260 7900
rect 2340 7820 2350 7900
rect 2250 7810 2350 7820
rect 2450 7900 2550 7910
rect 2450 7820 2460 7900
rect 2540 7820 2550 7900
rect 2450 7810 2550 7820
rect 2650 7900 2750 7910
rect 2650 7820 2660 7900
rect 2740 7820 2750 7900
rect 2650 7810 2750 7820
rect 2850 7900 2950 7910
rect 2850 7820 2860 7900
rect 2940 7820 2950 7900
rect 2850 7810 2950 7820
rect 3050 7900 3150 7910
rect 3050 7820 3060 7900
rect 3140 7820 3150 7900
rect 3050 7810 3150 7820
rect 3250 7900 3350 7910
rect 3250 7820 3260 7900
rect 3340 7820 3350 7900
rect 3250 7810 3350 7820
rect 3450 7900 3550 7910
rect 3450 7820 3460 7900
rect 3540 7820 3550 7900
rect 3450 7810 3550 7820
rect 3650 7900 3750 7910
rect 3650 7820 3660 7900
rect 3740 7820 3750 7900
rect 3650 7810 3750 7820
rect 3850 7900 3950 7910
rect 3850 7820 3860 7900
rect 3940 7820 3950 7900
rect 3850 7810 3950 7820
rect 4050 7900 4150 7910
rect 4050 7820 4060 7900
rect 4140 7820 4150 7900
rect 4050 7810 4150 7820
rect 4250 7900 4350 7910
rect 4250 7820 4260 7900
rect 4340 7820 4350 7900
rect 4250 7810 4350 7820
rect 4450 7900 4550 7910
rect 4450 7820 4460 7900
rect 4540 7820 4550 7900
rect 4450 7810 4550 7820
rect 4650 7900 4750 7910
rect 4650 7820 4660 7900
rect 4740 7820 4750 7900
rect 4650 7810 4750 7820
rect 4850 7900 4950 7910
rect 4850 7820 4860 7900
rect 4940 7820 4950 7900
rect 4850 7810 4950 7820
rect 5050 7900 5150 7910
rect 5050 7820 5060 7900
rect 5140 7820 5150 7900
rect 5050 7810 5150 7820
rect 5250 7900 5350 7910
rect 5250 7820 5260 7900
rect 5340 7820 5350 7900
rect 5250 7810 5350 7820
rect 5450 7900 5550 7910
rect 5450 7820 5460 7900
rect 5540 7820 5550 7900
rect 5450 7810 5550 7820
rect 5650 7900 5750 7910
rect 5650 7820 5660 7900
rect 5740 7820 5750 7900
rect 5650 7810 5750 7820
rect 5850 7900 5950 7910
rect 5850 7820 5860 7900
rect 5940 7820 5950 7900
rect 5850 7810 5950 7820
rect 6050 7900 6150 7910
rect 6050 7820 6060 7900
rect 6140 7820 6150 7900
rect 6050 7810 6150 7820
rect 6250 7900 6350 7910
rect 6250 7820 6260 7900
rect 6340 7820 6350 7900
rect 6250 7810 6350 7820
rect 6450 7900 6550 7910
rect 6450 7820 6460 7900
rect 6540 7820 6550 7900
rect 6450 7810 6550 7820
rect -115 7725 -85 7810
rect 85 7725 115 7810
rect 285 7725 315 7810
rect 485 7725 515 7810
rect 685 7725 715 7810
rect 885 7725 915 7810
rect 1085 7725 1115 7810
rect 1285 7725 1315 7810
rect 1485 7725 1515 7810
rect 1685 7725 1715 7810
rect 1885 7725 1915 7810
rect 2085 7725 2115 7810
rect 2285 7725 2315 7810
rect 2485 7725 2515 7810
rect 2685 7725 2715 7810
rect 2885 7725 2915 7810
rect 3085 7725 3115 7810
rect 3285 7725 3315 7810
rect 3485 7725 3515 7810
rect 3685 7725 3715 7810
rect 3885 7725 3915 7810
rect 4085 7725 4115 7810
rect 4285 7725 4315 7810
rect 4485 7725 4515 7810
rect 4685 7725 4715 7810
rect 4885 7725 4915 7810
rect 5085 7725 5115 7810
rect 5285 7725 5315 7810
rect 5485 7725 5515 7810
rect 5685 7725 5715 7810
rect 5885 7725 5915 7810
rect 6085 7725 6115 7810
rect 6285 7725 6315 7810
rect 6485 7725 6515 7810
rect -150 7715 -50 7725
rect -150 7635 -140 7715
rect -60 7635 -50 7715
rect -150 7625 -50 7635
rect 50 7715 150 7725
rect 50 7635 60 7715
rect 140 7635 150 7715
rect 50 7625 150 7635
rect 250 7715 350 7725
rect 250 7635 260 7715
rect 340 7635 350 7715
rect 250 7625 350 7635
rect 450 7715 550 7725
rect 450 7635 460 7715
rect 540 7635 550 7715
rect 450 7625 550 7635
rect 650 7715 750 7725
rect 650 7635 660 7715
rect 740 7635 750 7715
rect 650 7625 750 7635
rect 850 7715 950 7725
rect 850 7635 860 7715
rect 940 7635 950 7715
rect 850 7625 950 7635
rect 1050 7715 1150 7725
rect 1050 7635 1060 7715
rect 1140 7635 1150 7715
rect 1050 7625 1150 7635
rect 1250 7715 1350 7725
rect 1250 7635 1260 7715
rect 1340 7635 1350 7715
rect 1250 7625 1350 7635
rect 1450 7715 1550 7725
rect 1450 7635 1460 7715
rect 1540 7635 1550 7715
rect 1450 7625 1550 7635
rect 1650 7715 1750 7725
rect 1650 7635 1660 7715
rect 1740 7635 1750 7715
rect 1650 7625 1750 7635
rect 1850 7715 1950 7725
rect 1850 7635 1860 7715
rect 1940 7635 1950 7715
rect 1850 7625 1950 7635
rect 2050 7715 2150 7725
rect 2050 7635 2060 7715
rect 2140 7635 2150 7715
rect 2050 7625 2150 7635
rect 2250 7715 2350 7725
rect 2250 7635 2260 7715
rect 2340 7635 2350 7715
rect 2250 7625 2350 7635
rect 2450 7715 2550 7725
rect 2450 7635 2460 7715
rect 2540 7635 2550 7715
rect 2450 7625 2550 7635
rect 2650 7715 2750 7725
rect 2650 7635 2660 7715
rect 2740 7635 2750 7715
rect 2650 7625 2750 7635
rect 2850 7715 2950 7725
rect 2850 7635 2860 7715
rect 2940 7635 2950 7715
rect 2850 7625 2950 7635
rect 3050 7715 3150 7725
rect 3050 7635 3060 7715
rect 3140 7635 3150 7715
rect 3050 7625 3150 7635
rect 3250 7715 3350 7725
rect 3250 7635 3260 7715
rect 3340 7635 3350 7715
rect 3250 7625 3350 7635
rect 3450 7715 3550 7725
rect 3450 7635 3460 7715
rect 3540 7635 3550 7715
rect 3450 7625 3550 7635
rect 3650 7715 3750 7725
rect 3650 7635 3660 7715
rect 3740 7635 3750 7715
rect 3650 7625 3750 7635
rect 3850 7715 3950 7725
rect 3850 7635 3860 7715
rect 3940 7635 3950 7715
rect 3850 7625 3950 7635
rect 4050 7715 4150 7725
rect 4050 7635 4060 7715
rect 4140 7635 4150 7715
rect 4050 7625 4150 7635
rect 4250 7715 4350 7725
rect 4250 7635 4260 7715
rect 4340 7635 4350 7715
rect 4250 7625 4350 7635
rect 4450 7715 4550 7725
rect 4450 7635 4460 7715
rect 4540 7635 4550 7715
rect 4450 7625 4550 7635
rect 4650 7715 4750 7725
rect 4650 7635 4660 7715
rect 4740 7635 4750 7715
rect 4650 7625 4750 7635
rect 4850 7715 4950 7725
rect 4850 7635 4860 7715
rect 4940 7635 4950 7715
rect 4850 7625 4950 7635
rect 5050 7715 5150 7725
rect 5050 7635 5060 7715
rect 5140 7635 5150 7715
rect 5050 7625 5150 7635
rect 5250 7715 5350 7725
rect 5250 7635 5260 7715
rect 5340 7635 5350 7715
rect 5250 7625 5350 7635
rect 5450 7715 5550 7725
rect 5450 7635 5460 7715
rect 5540 7635 5550 7715
rect 5450 7625 5550 7635
rect 5650 7715 5750 7725
rect 5650 7635 5660 7715
rect 5740 7635 5750 7715
rect 5650 7625 5750 7635
rect 5850 7715 5950 7725
rect 5850 7635 5860 7715
rect 5940 7635 5950 7715
rect 5850 7625 5950 7635
rect 6050 7715 6150 7725
rect 6050 7635 6060 7715
rect 6140 7635 6150 7715
rect 6050 7625 6150 7635
rect 6250 7715 6350 7725
rect 6250 7635 6260 7715
rect 6340 7635 6350 7715
rect 6250 7625 6350 7635
rect 6450 7715 6550 7725
rect 6450 7635 6460 7715
rect 6540 7635 6550 7715
rect 6450 7625 6550 7635
rect -115 7540 -85 7625
rect 85 7540 115 7625
rect 285 7540 315 7625
rect 485 7540 515 7625
rect 685 7540 715 7625
rect 885 7540 915 7625
rect 1085 7540 1115 7625
rect 1285 7540 1315 7625
rect 1485 7540 1515 7625
rect 1685 7540 1715 7625
rect 1885 7540 1915 7625
rect 2085 7540 2115 7625
rect 2285 7540 2315 7625
rect 2485 7540 2515 7625
rect 2685 7540 2715 7625
rect 2885 7540 2915 7625
rect 3085 7540 3115 7625
rect 3285 7540 3315 7625
rect 3485 7540 3515 7625
rect 3685 7540 3715 7625
rect 3885 7540 3915 7625
rect 4085 7540 4115 7625
rect 4285 7540 4315 7625
rect 4485 7540 4515 7625
rect 4685 7540 4715 7625
rect 4885 7540 4915 7625
rect 5085 7540 5115 7625
rect 5285 7540 5315 7625
rect 5485 7540 5515 7625
rect 5685 7540 5715 7625
rect 5885 7540 5915 7625
rect 6085 7540 6115 7625
rect 6285 7540 6315 7625
rect 6485 7540 6515 7625
rect -150 7530 -50 7540
rect -150 7450 -140 7530
rect -60 7450 -50 7530
rect -150 7440 -50 7450
rect 50 7530 150 7540
rect 50 7450 60 7530
rect 140 7450 150 7530
rect 50 7440 150 7450
rect 250 7530 350 7540
rect 250 7450 260 7530
rect 340 7450 350 7530
rect 250 7440 350 7450
rect 450 7530 550 7540
rect 450 7450 460 7530
rect 540 7450 550 7530
rect 450 7440 550 7450
rect 650 7530 750 7540
rect 650 7450 660 7530
rect 740 7450 750 7530
rect 650 7440 750 7450
rect 850 7530 950 7540
rect 850 7450 860 7530
rect 940 7450 950 7530
rect 850 7440 950 7450
rect 1050 7530 1150 7540
rect 1050 7450 1060 7530
rect 1140 7450 1150 7530
rect 1050 7440 1150 7450
rect 1250 7530 1350 7540
rect 1250 7450 1260 7530
rect 1340 7450 1350 7530
rect 1250 7440 1350 7450
rect 1450 7530 1550 7540
rect 1450 7450 1460 7530
rect 1540 7450 1550 7530
rect 1450 7440 1550 7450
rect 1650 7530 1750 7540
rect 1650 7450 1660 7530
rect 1740 7450 1750 7530
rect 1650 7440 1750 7450
rect 1850 7530 1950 7540
rect 1850 7450 1860 7530
rect 1940 7450 1950 7530
rect 1850 7440 1950 7450
rect 2050 7530 2150 7540
rect 2050 7450 2060 7530
rect 2140 7450 2150 7530
rect 2050 7440 2150 7450
rect 2250 7530 2350 7540
rect 2250 7450 2260 7530
rect 2340 7450 2350 7530
rect 2250 7440 2350 7450
rect 2450 7530 2550 7540
rect 2450 7450 2460 7530
rect 2540 7450 2550 7530
rect 2450 7440 2550 7450
rect 2650 7530 2750 7540
rect 2650 7450 2660 7530
rect 2740 7450 2750 7530
rect 2650 7440 2750 7450
rect 2850 7530 2950 7540
rect 2850 7450 2860 7530
rect 2940 7450 2950 7530
rect 2850 7440 2950 7450
rect 3050 7530 3150 7540
rect 3050 7450 3060 7530
rect 3140 7450 3150 7530
rect 3050 7440 3150 7450
rect 3250 7530 3350 7540
rect 3250 7450 3260 7530
rect 3340 7450 3350 7530
rect 3250 7440 3350 7450
rect 3450 7530 3550 7540
rect 3450 7450 3460 7530
rect 3540 7450 3550 7530
rect 3450 7440 3550 7450
rect 3650 7530 3750 7540
rect 3650 7450 3660 7530
rect 3740 7450 3750 7530
rect 3650 7440 3750 7450
rect 3850 7530 3950 7540
rect 3850 7450 3860 7530
rect 3940 7450 3950 7530
rect 3850 7440 3950 7450
rect 4050 7530 4150 7540
rect 4050 7450 4060 7530
rect 4140 7450 4150 7530
rect 4050 7440 4150 7450
rect 4250 7530 4350 7540
rect 4250 7450 4260 7530
rect 4340 7450 4350 7530
rect 4250 7440 4350 7450
rect 4450 7530 4550 7540
rect 4450 7450 4460 7530
rect 4540 7450 4550 7530
rect 4450 7440 4550 7450
rect 4650 7530 4750 7540
rect 4650 7450 4660 7530
rect 4740 7450 4750 7530
rect 4650 7440 4750 7450
rect 4850 7530 4950 7540
rect 4850 7450 4860 7530
rect 4940 7450 4950 7530
rect 4850 7440 4950 7450
rect 5050 7530 5150 7540
rect 5050 7450 5060 7530
rect 5140 7450 5150 7530
rect 5050 7440 5150 7450
rect 5250 7530 5350 7540
rect 5250 7450 5260 7530
rect 5340 7450 5350 7530
rect 5250 7440 5350 7450
rect 5450 7530 5550 7540
rect 5450 7450 5460 7530
rect 5540 7450 5550 7530
rect 5450 7440 5550 7450
rect 5650 7530 5750 7540
rect 5650 7450 5660 7530
rect 5740 7450 5750 7530
rect 5650 7440 5750 7450
rect 5850 7530 5950 7540
rect 5850 7450 5860 7530
rect 5940 7450 5950 7530
rect 5850 7440 5950 7450
rect 6050 7530 6150 7540
rect 6050 7450 6060 7530
rect 6140 7450 6150 7530
rect 6050 7440 6150 7450
rect 6250 7530 6350 7540
rect 6250 7450 6260 7530
rect 6340 7450 6350 7530
rect 6250 7440 6350 7450
rect 6450 7530 6550 7540
rect 6450 7450 6460 7530
rect 6540 7450 6550 7530
rect 6450 7440 6550 7450
rect -115 7355 -85 7440
rect 85 7355 115 7440
rect 285 7355 315 7440
rect 485 7355 515 7440
rect 685 7355 715 7440
rect 885 7355 915 7440
rect 1085 7355 1115 7440
rect 1285 7355 1315 7440
rect 1485 7355 1515 7440
rect 1685 7355 1715 7440
rect 1885 7355 1915 7440
rect 2085 7355 2115 7440
rect 2285 7355 2315 7440
rect 2485 7355 2515 7440
rect 2685 7355 2715 7440
rect 2885 7355 2915 7440
rect 3085 7355 3115 7440
rect 3285 7355 3315 7440
rect 3485 7355 3515 7440
rect 3685 7355 3715 7440
rect 3885 7355 3915 7440
rect 4085 7355 4115 7440
rect 4285 7355 4315 7440
rect 4485 7355 4515 7440
rect 4685 7355 4715 7440
rect 4885 7355 4915 7440
rect 5085 7355 5115 7440
rect 5285 7355 5315 7440
rect 5485 7355 5515 7440
rect 5685 7355 5715 7440
rect 5885 7355 5915 7440
rect 6085 7355 6115 7440
rect 6285 7355 6315 7440
rect 6485 7355 6515 7440
rect -150 7345 -50 7355
rect -150 7265 -140 7345
rect -60 7265 -50 7345
rect -150 7255 -50 7265
rect 50 7345 150 7355
rect 50 7265 60 7345
rect 140 7265 150 7345
rect 50 7255 150 7265
rect 250 7345 350 7355
rect 250 7265 260 7345
rect 340 7265 350 7345
rect 250 7255 350 7265
rect 450 7345 550 7355
rect 450 7265 460 7345
rect 540 7265 550 7345
rect 450 7255 550 7265
rect 650 7345 750 7355
rect 650 7265 660 7345
rect 740 7265 750 7345
rect 650 7255 750 7265
rect 850 7345 950 7355
rect 850 7265 860 7345
rect 940 7265 950 7345
rect 850 7255 950 7265
rect 1050 7345 1150 7355
rect 1050 7265 1060 7345
rect 1140 7265 1150 7345
rect 1050 7255 1150 7265
rect 1250 7345 1350 7355
rect 1250 7265 1260 7345
rect 1340 7265 1350 7345
rect 1250 7255 1350 7265
rect 1450 7345 1550 7355
rect 1450 7265 1460 7345
rect 1540 7265 1550 7345
rect 1450 7255 1550 7265
rect 1650 7345 1750 7355
rect 1650 7265 1660 7345
rect 1740 7265 1750 7345
rect 1650 7255 1750 7265
rect 1850 7345 1950 7355
rect 1850 7265 1860 7345
rect 1940 7265 1950 7345
rect 1850 7255 1950 7265
rect 2050 7345 2150 7355
rect 2050 7265 2060 7345
rect 2140 7265 2150 7345
rect 2050 7255 2150 7265
rect 2250 7345 2350 7355
rect 2250 7265 2260 7345
rect 2340 7265 2350 7345
rect 2250 7255 2350 7265
rect 2450 7345 2550 7355
rect 2450 7265 2460 7345
rect 2540 7265 2550 7345
rect 2450 7255 2550 7265
rect 2650 7345 2750 7355
rect 2650 7265 2660 7345
rect 2740 7265 2750 7345
rect 2650 7255 2750 7265
rect 2850 7345 2950 7355
rect 2850 7265 2860 7345
rect 2940 7265 2950 7345
rect 2850 7255 2950 7265
rect 3050 7345 3150 7355
rect 3050 7265 3060 7345
rect 3140 7265 3150 7345
rect 3050 7255 3150 7265
rect 3250 7345 3350 7355
rect 3250 7265 3260 7345
rect 3340 7265 3350 7345
rect 3250 7255 3350 7265
rect 3450 7345 3550 7355
rect 3450 7265 3460 7345
rect 3540 7265 3550 7345
rect 3450 7255 3550 7265
rect 3650 7345 3750 7355
rect 3650 7265 3660 7345
rect 3740 7265 3750 7345
rect 3650 7255 3750 7265
rect 3850 7345 3950 7355
rect 3850 7265 3860 7345
rect 3940 7265 3950 7345
rect 3850 7255 3950 7265
rect 4050 7345 4150 7355
rect 4050 7265 4060 7345
rect 4140 7265 4150 7345
rect 4050 7255 4150 7265
rect 4250 7345 4350 7355
rect 4250 7265 4260 7345
rect 4340 7265 4350 7345
rect 4250 7255 4350 7265
rect 4450 7345 4550 7355
rect 4450 7265 4460 7345
rect 4540 7265 4550 7345
rect 4450 7255 4550 7265
rect 4650 7345 4750 7355
rect 4650 7265 4660 7345
rect 4740 7265 4750 7345
rect 4650 7255 4750 7265
rect 4850 7345 4950 7355
rect 4850 7265 4860 7345
rect 4940 7265 4950 7345
rect 4850 7255 4950 7265
rect 5050 7345 5150 7355
rect 5050 7265 5060 7345
rect 5140 7265 5150 7345
rect 5050 7255 5150 7265
rect 5250 7345 5350 7355
rect 5250 7265 5260 7345
rect 5340 7265 5350 7345
rect 5250 7255 5350 7265
rect 5450 7345 5550 7355
rect 5450 7265 5460 7345
rect 5540 7265 5550 7345
rect 5450 7255 5550 7265
rect 5650 7345 5750 7355
rect 5650 7265 5660 7345
rect 5740 7265 5750 7345
rect 5650 7255 5750 7265
rect 5850 7345 5950 7355
rect 5850 7265 5860 7345
rect 5940 7265 5950 7345
rect 5850 7255 5950 7265
rect 6050 7345 6150 7355
rect 6050 7265 6060 7345
rect 6140 7265 6150 7345
rect 6050 7255 6150 7265
rect 6250 7345 6350 7355
rect 6250 7265 6260 7345
rect 6340 7265 6350 7345
rect 6250 7255 6350 7265
rect 6450 7345 6550 7355
rect 6450 7265 6460 7345
rect 6540 7265 6550 7345
rect 6450 7255 6550 7265
rect -115 7170 -85 7255
rect 85 7170 115 7255
rect 285 7170 315 7255
rect 485 7170 515 7255
rect 685 7170 715 7255
rect 885 7170 915 7255
rect 1085 7170 1115 7255
rect 1285 7170 1315 7255
rect 1485 7170 1515 7255
rect 1685 7170 1715 7255
rect 1885 7170 1915 7255
rect 2085 7170 2115 7255
rect 2285 7170 2315 7255
rect 2485 7170 2515 7255
rect 2685 7170 2715 7255
rect 2885 7170 2915 7255
rect 3085 7170 3115 7255
rect 3285 7170 3315 7255
rect 3485 7170 3515 7255
rect 3685 7170 3715 7255
rect 3885 7170 3915 7255
rect 4085 7170 4115 7255
rect 4285 7170 4315 7255
rect 4485 7170 4515 7255
rect 4685 7170 4715 7255
rect 4885 7170 4915 7255
rect 5085 7170 5115 7255
rect 5285 7170 5315 7255
rect 5485 7170 5515 7255
rect 5685 7170 5715 7255
rect 5885 7170 5915 7255
rect 6085 7170 6115 7255
rect 6285 7170 6315 7255
rect 6485 7170 6515 7255
rect -150 7160 -50 7170
rect -150 7080 -140 7160
rect -60 7080 -50 7160
rect -150 7070 -50 7080
rect 50 7160 150 7170
rect 50 7080 60 7160
rect 140 7080 150 7160
rect 50 7070 150 7080
rect 250 7160 350 7170
rect 250 7080 260 7160
rect 340 7080 350 7160
rect 250 7070 350 7080
rect 450 7160 550 7170
rect 450 7080 460 7160
rect 540 7080 550 7160
rect 450 7070 550 7080
rect 650 7160 750 7170
rect 650 7080 660 7160
rect 740 7080 750 7160
rect 650 7070 750 7080
rect 850 7160 950 7170
rect 850 7080 860 7160
rect 940 7080 950 7160
rect 850 7070 950 7080
rect 1050 7160 1150 7170
rect 1050 7080 1060 7160
rect 1140 7080 1150 7160
rect 1050 7070 1150 7080
rect 1250 7160 1350 7170
rect 1250 7080 1260 7160
rect 1340 7080 1350 7160
rect 1250 7070 1350 7080
rect 1450 7160 1550 7170
rect 1450 7080 1460 7160
rect 1540 7080 1550 7160
rect 1450 7070 1550 7080
rect 1650 7160 1750 7170
rect 1650 7080 1660 7160
rect 1740 7080 1750 7160
rect 1650 7070 1750 7080
rect 1850 7160 1950 7170
rect 1850 7080 1860 7160
rect 1940 7080 1950 7160
rect 1850 7070 1950 7080
rect 2050 7160 2150 7170
rect 2050 7080 2060 7160
rect 2140 7080 2150 7160
rect 2050 7070 2150 7080
rect 2250 7160 2350 7170
rect 2250 7080 2260 7160
rect 2340 7080 2350 7160
rect 2250 7070 2350 7080
rect 2450 7160 2550 7170
rect 2450 7080 2460 7160
rect 2540 7080 2550 7160
rect 2450 7070 2550 7080
rect 2650 7160 2750 7170
rect 2650 7080 2660 7160
rect 2740 7080 2750 7160
rect 2650 7070 2750 7080
rect 2850 7160 2950 7170
rect 2850 7080 2860 7160
rect 2940 7080 2950 7160
rect 2850 7070 2950 7080
rect 3050 7160 3150 7170
rect 3050 7080 3060 7160
rect 3140 7080 3150 7160
rect 3050 7070 3150 7080
rect 3250 7160 3350 7170
rect 3250 7080 3260 7160
rect 3340 7080 3350 7160
rect 3250 7070 3350 7080
rect 3450 7160 3550 7170
rect 3450 7080 3460 7160
rect 3540 7080 3550 7160
rect 3450 7070 3550 7080
rect 3650 7160 3750 7170
rect 3650 7080 3660 7160
rect 3740 7080 3750 7160
rect 3650 7070 3750 7080
rect 3850 7160 3950 7170
rect 3850 7080 3860 7160
rect 3940 7080 3950 7160
rect 3850 7070 3950 7080
rect 4050 7160 4150 7170
rect 4050 7080 4060 7160
rect 4140 7080 4150 7160
rect 4050 7070 4150 7080
rect 4250 7160 4350 7170
rect 4250 7080 4260 7160
rect 4340 7080 4350 7160
rect 4250 7070 4350 7080
rect 4450 7160 4550 7170
rect 4450 7080 4460 7160
rect 4540 7080 4550 7160
rect 4450 7070 4550 7080
rect 4650 7160 4750 7170
rect 4650 7080 4660 7160
rect 4740 7080 4750 7160
rect 4650 7070 4750 7080
rect 4850 7160 4950 7170
rect 4850 7080 4860 7160
rect 4940 7080 4950 7160
rect 4850 7070 4950 7080
rect 5050 7160 5150 7170
rect 5050 7080 5060 7160
rect 5140 7080 5150 7160
rect 5050 7070 5150 7080
rect 5250 7160 5350 7170
rect 5250 7080 5260 7160
rect 5340 7080 5350 7160
rect 5250 7070 5350 7080
rect 5450 7160 5550 7170
rect 5450 7080 5460 7160
rect 5540 7080 5550 7160
rect 5450 7070 5550 7080
rect 5650 7160 5750 7170
rect 5650 7080 5660 7160
rect 5740 7080 5750 7160
rect 5650 7070 5750 7080
rect 5850 7160 5950 7170
rect 5850 7080 5860 7160
rect 5940 7080 5950 7160
rect 5850 7070 5950 7080
rect 6050 7160 6150 7170
rect 6050 7080 6060 7160
rect 6140 7080 6150 7160
rect 6050 7070 6150 7080
rect 6250 7160 6350 7170
rect 6250 7080 6260 7160
rect 6340 7080 6350 7160
rect 6250 7070 6350 7080
rect 6450 7160 6550 7170
rect 6450 7080 6460 7160
rect 6540 7080 6550 7160
rect 6450 7070 6550 7080
rect -115 6985 -85 7070
rect 85 6985 115 7070
rect 285 6985 315 7070
rect 485 6985 515 7070
rect 685 6985 715 7070
rect 885 6985 915 7070
rect 1085 6985 1115 7070
rect 1285 6985 1315 7070
rect 1485 6985 1515 7070
rect 1685 6985 1715 7070
rect 1885 6985 1915 7070
rect 2085 6985 2115 7070
rect 2285 6985 2315 7070
rect 2485 6985 2515 7070
rect 2685 6985 2715 7070
rect 2885 6985 2915 7070
rect 3085 6985 3115 7070
rect 3285 6985 3315 7070
rect 3485 6985 3515 7070
rect 3685 6985 3715 7070
rect 3885 6985 3915 7070
rect 4085 6985 4115 7070
rect 4285 6985 4315 7070
rect 4485 6985 4515 7070
rect 4685 6985 4715 7070
rect 4885 6985 4915 7070
rect 5085 6985 5115 7070
rect 5285 6985 5315 7070
rect 5485 6985 5515 7070
rect 5685 6985 5715 7070
rect 5885 6985 5915 7070
rect 6085 6985 6115 7070
rect 6285 6985 6315 7070
rect 6485 6985 6515 7070
rect -150 6975 -50 6985
rect -150 6895 -140 6975
rect -60 6895 -50 6975
rect -150 6885 -50 6895
rect 50 6975 150 6985
rect 50 6895 60 6975
rect 140 6895 150 6975
rect 50 6885 150 6895
rect 250 6975 350 6985
rect 250 6895 260 6975
rect 340 6895 350 6975
rect 250 6885 350 6895
rect 450 6975 550 6985
rect 450 6895 460 6975
rect 540 6895 550 6975
rect 450 6885 550 6895
rect 650 6975 750 6985
rect 650 6895 660 6975
rect 740 6895 750 6975
rect 650 6885 750 6895
rect 850 6975 950 6985
rect 850 6895 860 6975
rect 940 6895 950 6975
rect 850 6885 950 6895
rect 1050 6975 1150 6985
rect 1050 6895 1060 6975
rect 1140 6895 1150 6975
rect 1050 6885 1150 6895
rect 1250 6975 1350 6985
rect 1250 6895 1260 6975
rect 1340 6895 1350 6975
rect 1250 6885 1350 6895
rect 1450 6975 1550 6985
rect 1450 6895 1460 6975
rect 1540 6895 1550 6975
rect 1450 6885 1550 6895
rect 1650 6975 1750 6985
rect 1650 6895 1660 6975
rect 1740 6895 1750 6975
rect 1650 6885 1750 6895
rect 1850 6975 1950 6985
rect 1850 6895 1860 6975
rect 1940 6895 1950 6975
rect 1850 6885 1950 6895
rect 2050 6975 2150 6985
rect 2050 6895 2060 6975
rect 2140 6895 2150 6975
rect 2050 6885 2150 6895
rect 2250 6975 2350 6985
rect 2250 6895 2260 6975
rect 2340 6895 2350 6975
rect 2250 6885 2350 6895
rect 2450 6975 2550 6985
rect 2450 6895 2460 6975
rect 2540 6895 2550 6975
rect 2450 6885 2550 6895
rect 2650 6975 2750 6985
rect 2650 6895 2660 6975
rect 2740 6895 2750 6975
rect 2650 6885 2750 6895
rect 2850 6975 2950 6985
rect 2850 6895 2860 6975
rect 2940 6895 2950 6975
rect 2850 6885 2950 6895
rect 3050 6975 3150 6985
rect 3050 6895 3060 6975
rect 3140 6895 3150 6975
rect 3050 6885 3150 6895
rect 3250 6975 3350 6985
rect 3250 6895 3260 6975
rect 3340 6895 3350 6975
rect 3250 6885 3350 6895
rect 3450 6975 3550 6985
rect 3450 6895 3460 6975
rect 3540 6895 3550 6975
rect 3450 6885 3550 6895
rect 3650 6975 3750 6985
rect 3650 6895 3660 6975
rect 3740 6895 3750 6975
rect 3650 6885 3750 6895
rect 3850 6975 3950 6985
rect 3850 6895 3860 6975
rect 3940 6895 3950 6975
rect 3850 6885 3950 6895
rect 4050 6975 4150 6985
rect 4050 6895 4060 6975
rect 4140 6895 4150 6975
rect 4050 6885 4150 6895
rect 4250 6975 4350 6985
rect 4250 6895 4260 6975
rect 4340 6895 4350 6975
rect 4250 6885 4350 6895
rect 4450 6975 4550 6985
rect 4450 6895 4460 6975
rect 4540 6895 4550 6975
rect 4450 6885 4550 6895
rect 4650 6975 4750 6985
rect 4650 6895 4660 6975
rect 4740 6895 4750 6975
rect 4650 6885 4750 6895
rect 4850 6975 4950 6985
rect 4850 6895 4860 6975
rect 4940 6895 4950 6975
rect 4850 6885 4950 6895
rect 5050 6975 5150 6985
rect 5050 6895 5060 6975
rect 5140 6895 5150 6975
rect 5050 6885 5150 6895
rect 5250 6975 5350 6985
rect 5250 6895 5260 6975
rect 5340 6895 5350 6975
rect 5250 6885 5350 6895
rect 5450 6975 5550 6985
rect 5450 6895 5460 6975
rect 5540 6895 5550 6975
rect 5450 6885 5550 6895
rect 5650 6975 5750 6985
rect 5650 6895 5660 6975
rect 5740 6895 5750 6975
rect 5650 6885 5750 6895
rect 5850 6975 5950 6985
rect 5850 6895 5860 6975
rect 5940 6895 5950 6975
rect 5850 6885 5950 6895
rect 6050 6975 6150 6985
rect 6050 6895 6060 6975
rect 6140 6895 6150 6975
rect 6050 6885 6150 6895
rect 6250 6975 6350 6985
rect 6250 6895 6260 6975
rect 6340 6895 6350 6975
rect 6250 6885 6350 6895
rect 6450 6975 6550 6985
rect 6450 6895 6460 6975
rect 6540 6895 6550 6975
rect 6450 6885 6550 6895
rect -115 6800 -85 6885
rect 85 6800 115 6885
rect 285 6800 315 6885
rect 485 6800 515 6885
rect 685 6800 715 6885
rect 885 6800 915 6885
rect 1085 6800 1115 6885
rect 1285 6800 1315 6885
rect 1485 6800 1515 6885
rect 1685 6800 1715 6885
rect 1885 6800 1915 6885
rect 2085 6800 2115 6885
rect 2285 6800 2315 6885
rect 2485 6800 2515 6885
rect 2685 6800 2715 6885
rect 2885 6800 2915 6885
rect 3085 6800 3115 6885
rect 3285 6800 3315 6885
rect 3485 6800 3515 6885
rect 3685 6800 3715 6885
rect 3885 6800 3915 6885
rect 4085 6800 4115 6885
rect 4285 6800 4315 6885
rect 4485 6800 4515 6885
rect 4685 6800 4715 6885
rect 4885 6800 4915 6885
rect 5085 6800 5115 6885
rect 5285 6800 5315 6885
rect 5485 6800 5515 6885
rect 5685 6800 5715 6885
rect 5885 6800 5915 6885
rect 6085 6800 6115 6885
rect 6285 6800 6315 6885
rect 6485 6800 6515 6885
rect -150 6790 -50 6800
rect -150 6710 -140 6790
rect -60 6710 -50 6790
rect -150 6700 -50 6710
rect 50 6790 150 6800
rect 50 6710 60 6790
rect 140 6710 150 6790
rect 50 6700 150 6710
rect 250 6790 350 6800
rect 250 6710 260 6790
rect 340 6710 350 6790
rect 250 6700 350 6710
rect 450 6790 550 6800
rect 450 6710 460 6790
rect 540 6710 550 6790
rect 450 6700 550 6710
rect 650 6790 750 6800
rect 650 6710 660 6790
rect 740 6710 750 6790
rect 650 6700 750 6710
rect 850 6790 950 6800
rect 850 6710 860 6790
rect 940 6710 950 6790
rect 850 6700 950 6710
rect 1050 6790 1150 6800
rect 1050 6710 1060 6790
rect 1140 6710 1150 6790
rect 1050 6700 1150 6710
rect 1250 6790 1350 6800
rect 1250 6710 1260 6790
rect 1340 6710 1350 6790
rect 1250 6700 1350 6710
rect 1450 6790 1550 6800
rect 1450 6710 1460 6790
rect 1540 6710 1550 6790
rect 1450 6700 1550 6710
rect 1650 6790 1750 6800
rect 1650 6710 1660 6790
rect 1740 6710 1750 6790
rect 1650 6700 1750 6710
rect 1850 6790 1950 6800
rect 1850 6710 1860 6790
rect 1940 6710 1950 6790
rect 1850 6700 1950 6710
rect 2050 6790 2150 6800
rect 2050 6710 2060 6790
rect 2140 6710 2150 6790
rect 2050 6700 2150 6710
rect 2250 6790 2350 6800
rect 2250 6710 2260 6790
rect 2340 6710 2350 6790
rect 2250 6700 2350 6710
rect 2450 6790 2550 6800
rect 2450 6710 2460 6790
rect 2540 6710 2550 6790
rect 2450 6700 2550 6710
rect 2650 6790 2750 6800
rect 2650 6710 2660 6790
rect 2740 6710 2750 6790
rect 2650 6700 2750 6710
rect 2850 6790 2950 6800
rect 2850 6710 2860 6790
rect 2940 6710 2950 6790
rect 2850 6700 2950 6710
rect 3050 6790 3150 6800
rect 3050 6710 3060 6790
rect 3140 6710 3150 6790
rect 3050 6700 3150 6710
rect 3250 6790 3350 6800
rect 3250 6710 3260 6790
rect 3340 6710 3350 6790
rect 3250 6700 3350 6710
rect 3450 6790 3550 6800
rect 3450 6710 3460 6790
rect 3540 6710 3550 6790
rect 3450 6700 3550 6710
rect 3650 6790 3750 6800
rect 3650 6710 3660 6790
rect 3740 6710 3750 6790
rect 3650 6700 3750 6710
rect 3850 6790 3950 6800
rect 3850 6710 3860 6790
rect 3940 6710 3950 6790
rect 3850 6700 3950 6710
rect 4050 6790 4150 6800
rect 4050 6710 4060 6790
rect 4140 6710 4150 6790
rect 4050 6700 4150 6710
rect 4250 6790 4350 6800
rect 4250 6710 4260 6790
rect 4340 6710 4350 6790
rect 4250 6700 4350 6710
rect 4450 6790 4550 6800
rect 4450 6710 4460 6790
rect 4540 6710 4550 6790
rect 4450 6700 4550 6710
rect 4650 6790 4750 6800
rect 4650 6710 4660 6790
rect 4740 6710 4750 6790
rect 4650 6700 4750 6710
rect 4850 6790 4950 6800
rect 4850 6710 4860 6790
rect 4940 6710 4950 6790
rect 4850 6700 4950 6710
rect 5050 6790 5150 6800
rect 5050 6710 5060 6790
rect 5140 6710 5150 6790
rect 5050 6700 5150 6710
rect 5250 6790 5350 6800
rect 5250 6710 5260 6790
rect 5340 6710 5350 6790
rect 5250 6700 5350 6710
rect 5450 6790 5550 6800
rect 5450 6710 5460 6790
rect 5540 6710 5550 6790
rect 5450 6700 5550 6710
rect 5650 6790 5750 6800
rect 5650 6710 5660 6790
rect 5740 6710 5750 6790
rect 5650 6700 5750 6710
rect 5850 6790 5950 6800
rect 5850 6710 5860 6790
rect 5940 6710 5950 6790
rect 5850 6700 5950 6710
rect 6050 6790 6150 6800
rect 6050 6710 6060 6790
rect 6140 6710 6150 6790
rect 6050 6700 6150 6710
rect 6250 6790 6350 6800
rect 6250 6710 6260 6790
rect 6340 6710 6350 6790
rect 6250 6700 6350 6710
rect 6450 6790 6550 6800
rect 6450 6710 6460 6790
rect 6540 6710 6550 6790
rect 6450 6700 6550 6710
rect -115 6615 -85 6700
rect 85 6615 115 6700
rect 285 6615 315 6700
rect 485 6615 515 6700
rect 685 6615 715 6700
rect 885 6615 915 6700
rect 1085 6615 1115 6700
rect 1285 6615 1315 6700
rect 1485 6615 1515 6700
rect 1685 6615 1715 6700
rect 1885 6615 1915 6700
rect 2085 6615 2115 6700
rect 2285 6615 2315 6700
rect 2485 6615 2515 6700
rect 2685 6615 2715 6700
rect 2885 6615 2915 6700
rect 3085 6615 3115 6700
rect 3285 6615 3315 6700
rect 3485 6615 3515 6700
rect 3685 6615 3715 6700
rect 3885 6615 3915 6700
rect 4085 6615 4115 6700
rect 4285 6615 4315 6700
rect 4485 6615 4515 6700
rect 4685 6615 4715 6700
rect 4885 6615 4915 6700
rect 5085 6615 5115 6700
rect 5285 6615 5315 6700
rect 5485 6615 5515 6700
rect 5685 6615 5715 6700
rect 5885 6615 5915 6700
rect 6085 6615 6115 6700
rect 6285 6615 6315 6700
rect 6485 6615 6515 6700
rect -150 6605 -50 6615
rect -150 6525 -140 6605
rect -60 6525 -50 6605
rect -150 6515 -50 6525
rect 50 6605 150 6615
rect 50 6525 60 6605
rect 140 6525 150 6605
rect 50 6515 150 6525
rect 250 6605 350 6615
rect 250 6525 260 6605
rect 340 6525 350 6605
rect 250 6515 350 6525
rect 450 6605 550 6615
rect 450 6525 460 6605
rect 540 6525 550 6605
rect 450 6515 550 6525
rect 650 6605 750 6615
rect 650 6525 660 6605
rect 740 6525 750 6605
rect 650 6515 750 6525
rect 850 6605 950 6615
rect 850 6525 860 6605
rect 940 6525 950 6605
rect 850 6515 950 6525
rect 1050 6605 1150 6615
rect 1050 6525 1060 6605
rect 1140 6525 1150 6605
rect 1050 6515 1150 6525
rect 1250 6605 1350 6615
rect 1250 6525 1260 6605
rect 1340 6525 1350 6605
rect 1250 6515 1350 6525
rect 1450 6605 1550 6615
rect 1450 6525 1460 6605
rect 1540 6525 1550 6605
rect 1450 6515 1550 6525
rect 1650 6605 1750 6615
rect 1650 6525 1660 6605
rect 1740 6525 1750 6605
rect 1650 6515 1750 6525
rect 1850 6605 1950 6615
rect 1850 6525 1860 6605
rect 1940 6525 1950 6605
rect 1850 6515 1950 6525
rect 2050 6605 2150 6615
rect 2050 6525 2060 6605
rect 2140 6525 2150 6605
rect 2050 6515 2150 6525
rect 2250 6605 2350 6615
rect 2250 6525 2260 6605
rect 2340 6525 2350 6605
rect 2250 6515 2350 6525
rect 2450 6605 2550 6615
rect 2450 6525 2460 6605
rect 2540 6525 2550 6605
rect 2450 6515 2550 6525
rect 2650 6605 2750 6615
rect 2650 6525 2660 6605
rect 2740 6525 2750 6605
rect 2650 6515 2750 6525
rect 2850 6605 2950 6615
rect 2850 6525 2860 6605
rect 2940 6525 2950 6605
rect 2850 6515 2950 6525
rect 3050 6605 3150 6615
rect 3050 6525 3060 6605
rect 3140 6525 3150 6605
rect 3050 6515 3150 6525
rect 3250 6605 3350 6615
rect 3250 6525 3260 6605
rect 3340 6525 3350 6605
rect 3250 6515 3350 6525
rect 3450 6605 3550 6615
rect 3450 6525 3460 6605
rect 3540 6525 3550 6605
rect 3450 6515 3550 6525
rect 3650 6605 3750 6615
rect 3650 6525 3660 6605
rect 3740 6525 3750 6605
rect 3650 6515 3750 6525
rect 3850 6605 3950 6615
rect 3850 6525 3860 6605
rect 3940 6525 3950 6605
rect 3850 6515 3950 6525
rect 4050 6605 4150 6615
rect 4050 6525 4060 6605
rect 4140 6525 4150 6605
rect 4050 6515 4150 6525
rect 4250 6605 4350 6615
rect 4250 6525 4260 6605
rect 4340 6525 4350 6605
rect 4250 6515 4350 6525
rect 4450 6605 4550 6615
rect 4450 6525 4460 6605
rect 4540 6525 4550 6605
rect 4450 6515 4550 6525
rect 4650 6605 4750 6615
rect 4650 6525 4660 6605
rect 4740 6525 4750 6605
rect 4650 6515 4750 6525
rect 4850 6605 4950 6615
rect 4850 6525 4860 6605
rect 4940 6525 4950 6605
rect 4850 6515 4950 6525
rect 5050 6605 5150 6615
rect 5050 6525 5060 6605
rect 5140 6525 5150 6605
rect 5050 6515 5150 6525
rect 5250 6605 5350 6615
rect 5250 6525 5260 6605
rect 5340 6525 5350 6605
rect 5250 6515 5350 6525
rect 5450 6605 5550 6615
rect 5450 6525 5460 6605
rect 5540 6525 5550 6605
rect 5450 6515 5550 6525
rect 5650 6605 5750 6615
rect 5650 6525 5660 6605
rect 5740 6525 5750 6605
rect 5650 6515 5750 6525
rect 5850 6605 5950 6615
rect 5850 6525 5860 6605
rect 5940 6525 5950 6605
rect 5850 6515 5950 6525
rect 6050 6605 6150 6615
rect 6050 6525 6060 6605
rect 6140 6525 6150 6605
rect 6050 6515 6150 6525
rect 6250 6605 6350 6615
rect 6250 6525 6260 6605
rect 6340 6525 6350 6605
rect 6250 6515 6350 6525
rect 6450 6605 6550 6615
rect 6450 6525 6460 6605
rect 6540 6525 6550 6605
rect 6450 6515 6550 6525
rect -115 6430 -85 6515
rect 85 6430 115 6515
rect 285 6430 315 6515
rect 485 6430 515 6515
rect 685 6430 715 6515
rect 885 6430 915 6515
rect 1085 6430 1115 6515
rect 1285 6430 1315 6515
rect 1485 6430 1515 6515
rect 1685 6430 1715 6515
rect 1885 6430 1915 6515
rect 2085 6430 2115 6515
rect 2285 6430 2315 6515
rect 2485 6430 2515 6515
rect 2685 6430 2715 6515
rect 2885 6430 2915 6515
rect 3085 6430 3115 6515
rect 3285 6430 3315 6515
rect 3485 6430 3515 6515
rect 3685 6430 3715 6515
rect 3885 6430 3915 6515
rect 4085 6430 4115 6515
rect 4285 6430 4315 6515
rect 4485 6430 4515 6515
rect 4685 6430 4715 6515
rect 4885 6430 4915 6515
rect 5085 6430 5115 6515
rect 5285 6430 5315 6515
rect 5485 6430 5515 6515
rect 5685 6430 5715 6515
rect 5885 6430 5915 6515
rect 6085 6430 6115 6515
rect 6285 6430 6315 6515
rect 6485 6430 6515 6515
rect -150 6420 -50 6430
rect -150 6340 -140 6420
rect -60 6340 -50 6420
rect -150 6330 -50 6340
rect 50 6420 150 6430
rect 50 6340 60 6420
rect 140 6340 150 6420
rect 50 6330 150 6340
rect 250 6420 350 6430
rect 250 6340 260 6420
rect 340 6340 350 6420
rect 250 6330 350 6340
rect 450 6420 550 6430
rect 450 6340 460 6420
rect 540 6340 550 6420
rect 450 6330 550 6340
rect 650 6420 750 6430
rect 650 6340 660 6420
rect 740 6340 750 6420
rect 650 6330 750 6340
rect 850 6420 950 6430
rect 850 6340 860 6420
rect 940 6340 950 6420
rect 850 6330 950 6340
rect 1050 6420 1150 6430
rect 1050 6340 1060 6420
rect 1140 6340 1150 6420
rect 1050 6330 1150 6340
rect 1250 6420 1350 6430
rect 1250 6340 1260 6420
rect 1340 6340 1350 6420
rect 1250 6330 1350 6340
rect 1450 6420 1550 6430
rect 1450 6340 1460 6420
rect 1540 6340 1550 6420
rect 1450 6330 1550 6340
rect 1650 6420 1750 6430
rect 1650 6340 1660 6420
rect 1740 6340 1750 6420
rect 1650 6330 1750 6340
rect 1850 6420 1950 6430
rect 1850 6340 1860 6420
rect 1940 6340 1950 6420
rect 1850 6330 1950 6340
rect 2050 6420 2150 6430
rect 2050 6340 2060 6420
rect 2140 6340 2150 6420
rect 2050 6330 2150 6340
rect 2250 6420 2350 6430
rect 2250 6340 2260 6420
rect 2340 6340 2350 6420
rect 2250 6330 2350 6340
rect 2450 6420 2550 6430
rect 2450 6340 2460 6420
rect 2540 6340 2550 6420
rect 2450 6330 2550 6340
rect 2650 6420 2750 6430
rect 2650 6340 2660 6420
rect 2740 6340 2750 6420
rect 2650 6330 2750 6340
rect 2850 6420 2950 6430
rect 2850 6340 2860 6420
rect 2940 6340 2950 6420
rect 2850 6330 2950 6340
rect 3050 6420 3150 6430
rect 3050 6340 3060 6420
rect 3140 6340 3150 6420
rect 3050 6330 3150 6340
rect 3250 6420 3350 6430
rect 3250 6340 3260 6420
rect 3340 6340 3350 6420
rect 3250 6330 3350 6340
rect 3450 6420 3550 6430
rect 3450 6340 3460 6420
rect 3540 6340 3550 6420
rect 3450 6330 3550 6340
rect 3650 6420 3750 6430
rect 3650 6340 3660 6420
rect 3740 6340 3750 6420
rect 3650 6330 3750 6340
rect 3850 6420 3950 6430
rect 3850 6340 3860 6420
rect 3940 6340 3950 6420
rect 3850 6330 3950 6340
rect 4050 6420 4150 6430
rect 4050 6340 4060 6420
rect 4140 6340 4150 6420
rect 4050 6330 4150 6340
rect 4250 6420 4350 6430
rect 4250 6340 4260 6420
rect 4340 6340 4350 6420
rect 4250 6330 4350 6340
rect 4450 6420 4550 6430
rect 4450 6340 4460 6420
rect 4540 6340 4550 6420
rect 4450 6330 4550 6340
rect 4650 6420 4750 6430
rect 4650 6340 4660 6420
rect 4740 6340 4750 6420
rect 4650 6330 4750 6340
rect 4850 6420 4950 6430
rect 4850 6340 4860 6420
rect 4940 6340 4950 6420
rect 4850 6330 4950 6340
rect 5050 6420 5150 6430
rect 5050 6340 5060 6420
rect 5140 6340 5150 6420
rect 5050 6330 5150 6340
rect 5250 6420 5350 6430
rect 5250 6340 5260 6420
rect 5340 6340 5350 6420
rect 5250 6330 5350 6340
rect 5450 6420 5550 6430
rect 5450 6340 5460 6420
rect 5540 6340 5550 6420
rect 5450 6330 5550 6340
rect 5650 6420 5750 6430
rect 5650 6340 5660 6420
rect 5740 6340 5750 6420
rect 5650 6330 5750 6340
rect 5850 6420 5950 6430
rect 5850 6340 5860 6420
rect 5940 6340 5950 6420
rect 5850 6330 5950 6340
rect 6050 6420 6150 6430
rect 6050 6340 6060 6420
rect 6140 6340 6150 6420
rect 6050 6330 6150 6340
rect 6250 6420 6350 6430
rect 6250 6340 6260 6420
rect 6340 6340 6350 6420
rect 6250 6330 6350 6340
rect 6450 6420 6550 6430
rect 6450 6340 6460 6420
rect 6540 6340 6550 6420
rect 6450 6330 6550 6340
rect -115 6245 -85 6330
rect 85 6245 115 6330
rect 285 6245 315 6330
rect 485 6245 515 6330
rect 685 6245 715 6330
rect 885 6245 915 6330
rect 1085 6245 1115 6330
rect 1285 6245 1315 6330
rect 1485 6245 1515 6330
rect 1685 6245 1715 6330
rect 1885 6245 1915 6330
rect 2085 6245 2115 6330
rect 2285 6245 2315 6330
rect 2485 6245 2515 6330
rect 2685 6245 2715 6330
rect 2885 6245 2915 6330
rect 3085 6245 3115 6330
rect 3285 6245 3315 6330
rect 3485 6245 3515 6330
rect 3685 6245 3715 6330
rect 3885 6245 3915 6330
rect 4085 6245 4115 6330
rect 4285 6245 4315 6330
rect 4485 6245 4515 6330
rect 4685 6245 4715 6330
rect 4885 6245 4915 6330
rect 5085 6245 5115 6330
rect 5285 6245 5315 6330
rect 5485 6245 5515 6330
rect 5685 6245 5715 6330
rect 5885 6245 5915 6330
rect 6085 6245 6115 6330
rect 6285 6245 6315 6330
rect 6485 6245 6515 6330
rect -150 6235 -50 6245
rect -150 6155 -140 6235
rect -60 6155 -50 6235
rect -150 6145 -50 6155
rect 50 6235 150 6245
rect 50 6155 60 6235
rect 140 6155 150 6235
rect 50 6145 150 6155
rect 250 6235 350 6245
rect 250 6155 260 6235
rect 340 6155 350 6235
rect 250 6145 350 6155
rect 450 6235 550 6245
rect 450 6155 460 6235
rect 540 6155 550 6235
rect 450 6145 550 6155
rect 650 6235 750 6245
rect 650 6155 660 6235
rect 740 6155 750 6235
rect 650 6145 750 6155
rect 850 6235 950 6245
rect 850 6155 860 6235
rect 940 6155 950 6235
rect 850 6145 950 6155
rect 1050 6235 1150 6245
rect 1050 6155 1060 6235
rect 1140 6155 1150 6235
rect 1050 6145 1150 6155
rect 1250 6235 1350 6245
rect 1250 6155 1260 6235
rect 1340 6155 1350 6235
rect 1250 6145 1350 6155
rect 1450 6235 1550 6245
rect 1450 6155 1460 6235
rect 1540 6155 1550 6235
rect 1450 6145 1550 6155
rect 1650 6235 1750 6245
rect 1650 6155 1660 6235
rect 1740 6155 1750 6235
rect 1650 6145 1750 6155
rect 1850 6235 1950 6245
rect 1850 6155 1860 6235
rect 1940 6155 1950 6235
rect 1850 6145 1950 6155
rect 2050 6235 2150 6245
rect 2050 6155 2060 6235
rect 2140 6155 2150 6235
rect 2050 6145 2150 6155
rect 2250 6235 2350 6245
rect 2250 6155 2260 6235
rect 2340 6155 2350 6235
rect 2250 6145 2350 6155
rect 2450 6235 2550 6245
rect 2450 6155 2460 6235
rect 2540 6155 2550 6235
rect 2450 6145 2550 6155
rect 2650 6235 2750 6245
rect 2650 6155 2660 6235
rect 2740 6155 2750 6235
rect 2650 6145 2750 6155
rect 2850 6235 2950 6245
rect 2850 6155 2860 6235
rect 2940 6155 2950 6235
rect 2850 6145 2950 6155
rect 3050 6235 3150 6245
rect 3050 6155 3060 6235
rect 3140 6155 3150 6235
rect 3050 6145 3150 6155
rect 3250 6235 3350 6245
rect 3250 6155 3260 6235
rect 3340 6155 3350 6235
rect 3250 6145 3350 6155
rect 3450 6235 3550 6245
rect 3450 6155 3460 6235
rect 3540 6155 3550 6235
rect 3450 6145 3550 6155
rect 3650 6235 3750 6245
rect 3650 6155 3660 6235
rect 3740 6155 3750 6235
rect 3650 6145 3750 6155
rect 3850 6235 3950 6245
rect 3850 6155 3860 6235
rect 3940 6155 3950 6235
rect 3850 6145 3950 6155
rect 4050 6235 4150 6245
rect 4050 6155 4060 6235
rect 4140 6155 4150 6235
rect 4050 6145 4150 6155
rect 4250 6235 4350 6245
rect 4250 6155 4260 6235
rect 4340 6155 4350 6235
rect 4250 6145 4350 6155
rect 4450 6235 4550 6245
rect 4450 6155 4460 6235
rect 4540 6155 4550 6235
rect 4450 6145 4550 6155
rect 4650 6235 4750 6245
rect 4650 6155 4660 6235
rect 4740 6155 4750 6235
rect 4650 6145 4750 6155
rect 4850 6235 4950 6245
rect 4850 6155 4860 6235
rect 4940 6155 4950 6235
rect 4850 6145 4950 6155
rect 5050 6235 5150 6245
rect 5050 6155 5060 6235
rect 5140 6155 5150 6235
rect 5050 6145 5150 6155
rect 5250 6235 5350 6245
rect 5250 6155 5260 6235
rect 5340 6155 5350 6235
rect 5250 6145 5350 6155
rect 5450 6235 5550 6245
rect 5450 6155 5460 6235
rect 5540 6155 5550 6235
rect 5450 6145 5550 6155
rect 5650 6235 5750 6245
rect 5650 6155 5660 6235
rect 5740 6155 5750 6235
rect 5650 6145 5750 6155
rect 5850 6235 5950 6245
rect 5850 6155 5860 6235
rect 5940 6155 5950 6235
rect 5850 6145 5950 6155
rect 6050 6235 6150 6245
rect 6050 6155 6060 6235
rect 6140 6155 6150 6235
rect 6050 6145 6150 6155
rect 6250 6235 6350 6245
rect 6250 6155 6260 6235
rect 6340 6155 6350 6235
rect 6250 6145 6350 6155
rect 6450 6235 6550 6245
rect 6450 6155 6460 6235
rect 6540 6155 6550 6235
rect 6450 6145 6550 6155
rect -115 6060 -85 6145
rect 85 6060 115 6145
rect 285 6060 315 6145
rect 485 6060 515 6145
rect 685 6060 715 6145
rect 885 6060 915 6145
rect 1085 6060 1115 6145
rect 1285 6060 1315 6145
rect 1485 6060 1515 6145
rect 1685 6060 1715 6145
rect 1885 6060 1915 6145
rect 2085 6060 2115 6145
rect 2285 6060 2315 6145
rect 2485 6060 2515 6145
rect 2685 6060 2715 6145
rect 2885 6060 2915 6145
rect 3085 6060 3115 6145
rect 3285 6060 3315 6145
rect 3485 6060 3515 6145
rect 3685 6060 3715 6145
rect 3885 6060 3915 6145
rect 4085 6060 4115 6145
rect 4285 6060 4315 6145
rect 4485 6060 4515 6145
rect 4685 6060 4715 6145
rect 4885 6060 4915 6145
rect 5085 6060 5115 6145
rect 5285 6060 5315 6145
rect 5485 6060 5515 6145
rect 5685 6060 5715 6145
rect 5885 6060 5915 6145
rect 6085 6060 6115 6145
rect 6285 6060 6315 6145
rect 6485 6060 6515 6145
rect -150 6050 -50 6060
rect -150 5970 -140 6050
rect -60 5970 -50 6050
rect -150 5960 -50 5970
rect 50 6050 150 6060
rect 50 5970 60 6050
rect 140 5970 150 6050
rect 50 5960 150 5970
rect 250 6050 350 6060
rect 250 5970 260 6050
rect 340 5970 350 6050
rect 250 5960 350 5970
rect 450 6050 550 6060
rect 450 5970 460 6050
rect 540 5970 550 6050
rect 450 5960 550 5970
rect 650 6050 750 6060
rect 650 5970 660 6050
rect 740 5970 750 6050
rect 650 5960 750 5970
rect 850 6050 950 6060
rect 850 5970 860 6050
rect 940 5970 950 6050
rect 850 5960 950 5970
rect 1050 6050 1150 6060
rect 1050 5970 1060 6050
rect 1140 5970 1150 6050
rect 1050 5960 1150 5970
rect 1250 6050 1350 6060
rect 1250 5970 1260 6050
rect 1340 5970 1350 6050
rect 1250 5960 1350 5970
rect 1450 6050 1550 6060
rect 1450 5970 1460 6050
rect 1540 5970 1550 6050
rect 1450 5960 1550 5970
rect 1650 6050 1750 6060
rect 1650 5970 1660 6050
rect 1740 5970 1750 6050
rect 1650 5960 1750 5970
rect 1850 6050 1950 6060
rect 1850 5970 1860 6050
rect 1940 5970 1950 6050
rect 1850 5960 1950 5970
rect 2050 6050 2150 6060
rect 2050 5970 2060 6050
rect 2140 5970 2150 6050
rect 2050 5960 2150 5970
rect 2250 6050 2350 6060
rect 2250 5970 2260 6050
rect 2340 5970 2350 6050
rect 2250 5960 2350 5970
rect 2450 6050 2550 6060
rect 2450 5970 2460 6050
rect 2540 5970 2550 6050
rect 2450 5960 2550 5970
rect 2650 6050 2750 6060
rect 2650 5970 2660 6050
rect 2740 5970 2750 6050
rect 2650 5960 2750 5970
rect 2850 6050 2950 6060
rect 2850 5970 2860 6050
rect 2940 5970 2950 6050
rect 2850 5960 2950 5970
rect 3050 6050 3150 6060
rect 3050 5970 3060 6050
rect 3140 5970 3150 6050
rect 3050 5960 3150 5970
rect 3250 6050 3350 6060
rect 3250 5970 3260 6050
rect 3340 5970 3350 6050
rect 3250 5960 3350 5970
rect 3450 6050 3550 6060
rect 3450 5970 3460 6050
rect 3540 5970 3550 6050
rect 3450 5960 3550 5970
rect 3650 6050 3750 6060
rect 3650 5970 3660 6050
rect 3740 5970 3750 6050
rect 3650 5960 3750 5970
rect 3850 6050 3950 6060
rect 3850 5970 3860 6050
rect 3940 5970 3950 6050
rect 3850 5960 3950 5970
rect 4050 6050 4150 6060
rect 4050 5970 4060 6050
rect 4140 5970 4150 6050
rect 4050 5960 4150 5970
rect 4250 6050 4350 6060
rect 4250 5970 4260 6050
rect 4340 5970 4350 6050
rect 4250 5960 4350 5970
rect 4450 6050 4550 6060
rect 4450 5970 4460 6050
rect 4540 5970 4550 6050
rect 4450 5960 4550 5970
rect 4650 6050 4750 6060
rect 4650 5970 4660 6050
rect 4740 5970 4750 6050
rect 4650 5960 4750 5970
rect 4850 6050 4950 6060
rect 4850 5970 4860 6050
rect 4940 5970 4950 6050
rect 4850 5960 4950 5970
rect 5050 6050 5150 6060
rect 5050 5970 5060 6050
rect 5140 5970 5150 6050
rect 5050 5960 5150 5970
rect 5250 6050 5350 6060
rect 5250 5970 5260 6050
rect 5340 5970 5350 6050
rect 5250 5960 5350 5970
rect 5450 6050 5550 6060
rect 5450 5970 5460 6050
rect 5540 5970 5550 6050
rect 5450 5960 5550 5970
rect 5650 6050 5750 6060
rect 5650 5970 5660 6050
rect 5740 5970 5750 6050
rect 5650 5960 5750 5970
rect 5850 6050 5950 6060
rect 5850 5970 5860 6050
rect 5940 5970 5950 6050
rect 5850 5960 5950 5970
rect 6050 6050 6150 6060
rect 6050 5970 6060 6050
rect 6140 5970 6150 6050
rect 6050 5960 6150 5970
rect 6250 6050 6350 6060
rect 6250 5970 6260 6050
rect 6340 5970 6350 6050
rect 6250 5960 6350 5970
rect 6450 6050 6550 6060
rect 6450 5970 6460 6050
rect 6540 5970 6550 6050
rect 6450 5960 6550 5970
rect -115 5875 -85 5960
rect 85 5875 115 5960
rect 285 5875 315 5960
rect 485 5875 515 5960
rect 685 5875 715 5960
rect 885 5875 915 5960
rect 1085 5875 1115 5960
rect 1285 5875 1315 5960
rect 1485 5875 1515 5960
rect 1685 5875 1715 5960
rect 1885 5875 1915 5960
rect 2085 5875 2115 5960
rect 2285 5875 2315 5960
rect 2485 5875 2515 5960
rect 2685 5875 2715 5960
rect 2885 5875 2915 5960
rect 3085 5875 3115 5960
rect 3285 5875 3315 5960
rect 3485 5875 3515 5960
rect 3685 5875 3715 5960
rect 3885 5875 3915 5960
rect 4085 5875 4115 5960
rect 4285 5875 4315 5960
rect 4485 5875 4515 5960
rect 4685 5875 4715 5960
rect 4885 5875 4915 5960
rect 5085 5875 5115 5960
rect 5285 5875 5315 5960
rect 5485 5875 5515 5960
rect 5685 5875 5715 5960
rect 5885 5875 5915 5960
rect 6085 5875 6115 5960
rect 6285 5875 6315 5960
rect 6485 5875 6515 5960
rect -150 5865 -50 5875
rect -150 5785 -140 5865
rect -60 5785 -50 5865
rect -150 5775 -50 5785
rect 50 5865 150 5875
rect 50 5785 60 5865
rect 140 5785 150 5865
rect 50 5775 150 5785
rect 250 5865 350 5875
rect 250 5785 260 5865
rect 340 5785 350 5865
rect 250 5775 350 5785
rect 450 5865 550 5875
rect 450 5785 460 5865
rect 540 5785 550 5865
rect 450 5775 550 5785
rect 650 5865 750 5875
rect 650 5785 660 5865
rect 740 5785 750 5865
rect 650 5775 750 5785
rect 850 5865 950 5875
rect 850 5785 860 5865
rect 940 5785 950 5865
rect 850 5775 950 5785
rect 1050 5865 1150 5875
rect 1050 5785 1060 5865
rect 1140 5785 1150 5865
rect 1050 5775 1150 5785
rect 1250 5865 1350 5875
rect 1250 5785 1260 5865
rect 1340 5785 1350 5865
rect 1250 5775 1350 5785
rect 1450 5865 1550 5875
rect 1450 5785 1460 5865
rect 1540 5785 1550 5865
rect 1450 5775 1550 5785
rect 1650 5865 1750 5875
rect 1650 5785 1660 5865
rect 1740 5785 1750 5865
rect 1650 5775 1750 5785
rect 1850 5865 1950 5875
rect 1850 5785 1860 5865
rect 1940 5785 1950 5865
rect 1850 5775 1950 5785
rect 2050 5865 2150 5875
rect 2050 5785 2060 5865
rect 2140 5785 2150 5865
rect 2050 5775 2150 5785
rect 2250 5865 2350 5875
rect 2250 5785 2260 5865
rect 2340 5785 2350 5865
rect 2250 5775 2350 5785
rect 2450 5865 2550 5875
rect 2450 5785 2460 5865
rect 2540 5785 2550 5865
rect 2450 5775 2550 5785
rect 2650 5865 2750 5875
rect 2650 5785 2660 5865
rect 2740 5785 2750 5865
rect 2650 5775 2750 5785
rect 2850 5865 2950 5875
rect 2850 5785 2860 5865
rect 2940 5785 2950 5865
rect 2850 5775 2950 5785
rect 3050 5865 3150 5875
rect 3050 5785 3060 5865
rect 3140 5785 3150 5865
rect 3050 5775 3150 5785
rect 3250 5865 3350 5875
rect 3250 5785 3260 5865
rect 3340 5785 3350 5865
rect 3250 5775 3350 5785
rect 3450 5865 3550 5875
rect 3450 5785 3460 5865
rect 3540 5785 3550 5865
rect 3450 5775 3550 5785
rect 3650 5865 3750 5875
rect 3650 5785 3660 5865
rect 3740 5785 3750 5865
rect 3650 5775 3750 5785
rect 3850 5865 3950 5875
rect 3850 5785 3860 5865
rect 3940 5785 3950 5865
rect 3850 5775 3950 5785
rect 4050 5865 4150 5875
rect 4050 5785 4060 5865
rect 4140 5785 4150 5865
rect 4050 5775 4150 5785
rect 4250 5865 4350 5875
rect 4250 5785 4260 5865
rect 4340 5785 4350 5865
rect 4250 5775 4350 5785
rect 4450 5865 4550 5875
rect 4450 5785 4460 5865
rect 4540 5785 4550 5865
rect 4450 5775 4550 5785
rect 4650 5865 4750 5875
rect 4650 5785 4660 5865
rect 4740 5785 4750 5865
rect 4650 5775 4750 5785
rect 4850 5865 4950 5875
rect 4850 5785 4860 5865
rect 4940 5785 4950 5865
rect 4850 5775 4950 5785
rect 5050 5865 5150 5875
rect 5050 5785 5060 5865
rect 5140 5785 5150 5865
rect 5050 5775 5150 5785
rect 5250 5865 5350 5875
rect 5250 5785 5260 5865
rect 5340 5785 5350 5865
rect 5250 5775 5350 5785
rect 5450 5865 5550 5875
rect 5450 5785 5460 5865
rect 5540 5785 5550 5865
rect 5450 5775 5550 5785
rect 5650 5865 5750 5875
rect 5650 5785 5660 5865
rect 5740 5785 5750 5865
rect 5650 5775 5750 5785
rect 5850 5865 5950 5875
rect 5850 5785 5860 5865
rect 5940 5785 5950 5865
rect 5850 5775 5950 5785
rect 6050 5865 6150 5875
rect 6050 5785 6060 5865
rect 6140 5785 6150 5865
rect 6050 5775 6150 5785
rect 6250 5865 6350 5875
rect 6250 5785 6260 5865
rect 6340 5785 6350 5865
rect 6250 5775 6350 5785
rect 6450 5865 6550 5875
rect 6450 5785 6460 5865
rect 6540 5785 6550 5865
rect 6450 5775 6550 5785
rect -115 5690 -85 5775
rect 85 5690 115 5775
rect 285 5690 315 5775
rect 485 5690 515 5775
rect 685 5690 715 5775
rect 885 5690 915 5775
rect 1085 5690 1115 5775
rect 1285 5690 1315 5775
rect 1485 5690 1515 5775
rect 1685 5690 1715 5775
rect 1885 5690 1915 5775
rect 2085 5690 2115 5775
rect 2285 5690 2315 5775
rect 2485 5690 2515 5775
rect 2685 5690 2715 5775
rect 2885 5690 2915 5775
rect 3085 5690 3115 5775
rect 3285 5690 3315 5775
rect 3485 5690 3515 5775
rect 3685 5690 3715 5775
rect 3885 5690 3915 5775
rect 4085 5690 4115 5775
rect 4285 5690 4315 5775
rect 4485 5690 4515 5775
rect 4685 5690 4715 5775
rect 4885 5690 4915 5775
rect 5085 5690 5115 5775
rect 5285 5690 5315 5775
rect 5485 5690 5515 5775
rect 5685 5690 5715 5775
rect 5885 5690 5915 5775
rect 6085 5690 6115 5775
rect 6285 5690 6315 5775
rect 6485 5690 6515 5775
rect -150 5680 -50 5690
rect -150 5600 -140 5680
rect -60 5600 -50 5680
rect -150 5590 -50 5600
rect 50 5680 150 5690
rect 50 5600 60 5680
rect 140 5600 150 5680
rect 50 5590 150 5600
rect 250 5680 350 5690
rect 250 5600 260 5680
rect 340 5600 350 5680
rect 250 5590 350 5600
rect 450 5680 550 5690
rect 450 5600 460 5680
rect 540 5600 550 5680
rect 450 5590 550 5600
rect 650 5680 750 5690
rect 650 5600 660 5680
rect 740 5600 750 5680
rect 650 5590 750 5600
rect 850 5680 950 5690
rect 850 5600 860 5680
rect 940 5600 950 5680
rect 850 5590 950 5600
rect 1050 5680 1150 5690
rect 1050 5600 1060 5680
rect 1140 5600 1150 5680
rect 1050 5590 1150 5600
rect 1250 5680 1350 5690
rect 1250 5600 1260 5680
rect 1340 5600 1350 5680
rect 1250 5590 1350 5600
rect 1450 5680 1550 5690
rect 1450 5600 1460 5680
rect 1540 5600 1550 5680
rect 1450 5590 1550 5600
rect 1650 5680 1750 5690
rect 1650 5600 1660 5680
rect 1740 5600 1750 5680
rect 1650 5590 1750 5600
rect 1850 5680 1950 5690
rect 1850 5600 1860 5680
rect 1940 5600 1950 5680
rect 1850 5590 1950 5600
rect 2050 5680 2150 5690
rect 2050 5600 2060 5680
rect 2140 5600 2150 5680
rect 2050 5590 2150 5600
rect 2250 5680 2350 5690
rect 2250 5600 2260 5680
rect 2340 5600 2350 5680
rect 2250 5590 2350 5600
rect 2450 5680 2550 5690
rect 2450 5600 2460 5680
rect 2540 5600 2550 5680
rect 2450 5590 2550 5600
rect 2650 5680 2750 5690
rect 2650 5600 2660 5680
rect 2740 5600 2750 5680
rect 2650 5590 2750 5600
rect 2850 5680 2950 5690
rect 2850 5600 2860 5680
rect 2940 5600 2950 5680
rect 2850 5590 2950 5600
rect 3050 5680 3150 5690
rect 3050 5600 3060 5680
rect 3140 5600 3150 5680
rect 3050 5590 3150 5600
rect 3250 5680 3350 5690
rect 3250 5600 3260 5680
rect 3340 5600 3350 5680
rect 3250 5590 3350 5600
rect 3450 5680 3550 5690
rect 3450 5600 3460 5680
rect 3540 5600 3550 5680
rect 3450 5590 3550 5600
rect 3650 5680 3750 5690
rect 3650 5600 3660 5680
rect 3740 5600 3750 5680
rect 3650 5590 3750 5600
rect 3850 5680 3950 5690
rect 3850 5600 3860 5680
rect 3940 5600 3950 5680
rect 3850 5590 3950 5600
rect 4050 5680 4150 5690
rect 4050 5600 4060 5680
rect 4140 5600 4150 5680
rect 4050 5590 4150 5600
rect 4250 5680 4350 5690
rect 4250 5600 4260 5680
rect 4340 5600 4350 5680
rect 4250 5590 4350 5600
rect 4450 5680 4550 5690
rect 4450 5600 4460 5680
rect 4540 5600 4550 5680
rect 4450 5590 4550 5600
rect 4650 5680 4750 5690
rect 4650 5600 4660 5680
rect 4740 5600 4750 5680
rect 4650 5590 4750 5600
rect 4850 5680 4950 5690
rect 4850 5600 4860 5680
rect 4940 5600 4950 5680
rect 4850 5590 4950 5600
rect 5050 5680 5150 5690
rect 5050 5600 5060 5680
rect 5140 5600 5150 5680
rect 5050 5590 5150 5600
rect 5250 5680 5350 5690
rect 5250 5600 5260 5680
rect 5340 5600 5350 5680
rect 5250 5590 5350 5600
rect 5450 5680 5550 5690
rect 5450 5600 5460 5680
rect 5540 5600 5550 5680
rect 5450 5590 5550 5600
rect 5650 5680 5750 5690
rect 5650 5600 5660 5680
rect 5740 5600 5750 5680
rect 5650 5590 5750 5600
rect 5850 5680 5950 5690
rect 5850 5600 5860 5680
rect 5940 5600 5950 5680
rect 5850 5590 5950 5600
rect 6050 5680 6150 5690
rect 6050 5600 6060 5680
rect 6140 5600 6150 5680
rect 6050 5590 6150 5600
rect 6250 5680 6350 5690
rect 6250 5600 6260 5680
rect 6340 5600 6350 5680
rect 6250 5590 6350 5600
rect 6450 5680 6550 5690
rect 6450 5600 6460 5680
rect 6540 5600 6550 5680
rect 6450 5590 6550 5600
rect -115 5505 -85 5590
rect 85 5505 115 5590
rect 285 5505 315 5590
rect 485 5505 515 5590
rect 685 5505 715 5590
rect 885 5505 915 5590
rect 1085 5505 1115 5590
rect 1285 5505 1315 5590
rect 1485 5505 1515 5590
rect 1685 5505 1715 5590
rect 1885 5505 1915 5590
rect 2085 5505 2115 5590
rect 2285 5505 2315 5590
rect 2485 5505 2515 5590
rect 2685 5505 2715 5590
rect 2885 5505 2915 5590
rect 3085 5505 3115 5590
rect 3285 5505 3315 5590
rect 3485 5505 3515 5590
rect 3685 5505 3715 5590
rect 3885 5505 3915 5590
rect 4085 5505 4115 5590
rect 4285 5505 4315 5590
rect 4485 5505 4515 5590
rect 4685 5505 4715 5590
rect 4885 5505 4915 5590
rect 5085 5505 5115 5590
rect 5285 5505 5315 5590
rect 5485 5505 5515 5590
rect 5685 5505 5715 5590
rect 5885 5505 5915 5590
rect 6085 5505 6115 5590
rect 6285 5505 6315 5590
rect 6485 5505 6515 5590
rect -150 5495 -50 5505
rect -150 5415 -140 5495
rect -60 5415 -50 5495
rect -150 5405 -50 5415
rect 50 5495 150 5505
rect 50 5415 60 5495
rect 140 5415 150 5495
rect 50 5405 150 5415
rect 250 5495 350 5505
rect 250 5415 260 5495
rect 340 5415 350 5495
rect 250 5405 350 5415
rect 450 5495 550 5505
rect 450 5415 460 5495
rect 540 5415 550 5495
rect 450 5405 550 5415
rect 650 5495 750 5505
rect 650 5415 660 5495
rect 740 5415 750 5495
rect 650 5405 750 5415
rect 850 5495 950 5505
rect 850 5415 860 5495
rect 940 5415 950 5495
rect 850 5405 950 5415
rect 1050 5495 1150 5505
rect 1050 5415 1060 5495
rect 1140 5415 1150 5495
rect 1050 5405 1150 5415
rect 1250 5495 1350 5505
rect 1250 5415 1260 5495
rect 1340 5415 1350 5495
rect 1250 5405 1350 5415
rect 1450 5495 1550 5505
rect 1450 5415 1460 5495
rect 1540 5415 1550 5495
rect 1450 5405 1550 5415
rect 1650 5495 1750 5505
rect 1650 5415 1660 5495
rect 1740 5415 1750 5495
rect 1650 5405 1750 5415
rect 1850 5495 1950 5505
rect 1850 5415 1860 5495
rect 1940 5415 1950 5495
rect 1850 5405 1950 5415
rect 2050 5495 2150 5505
rect 2050 5415 2060 5495
rect 2140 5415 2150 5495
rect 2050 5405 2150 5415
rect 2250 5495 2350 5505
rect 2250 5415 2260 5495
rect 2340 5415 2350 5495
rect 2250 5405 2350 5415
rect 2450 5495 2550 5505
rect 2450 5415 2460 5495
rect 2540 5415 2550 5495
rect 2450 5405 2550 5415
rect 2650 5495 2750 5505
rect 2650 5415 2660 5495
rect 2740 5415 2750 5495
rect 2650 5405 2750 5415
rect 2850 5495 2950 5505
rect 2850 5415 2860 5495
rect 2940 5415 2950 5495
rect 2850 5405 2950 5415
rect 3050 5495 3150 5505
rect 3050 5415 3060 5495
rect 3140 5415 3150 5495
rect 3050 5405 3150 5415
rect 3250 5495 3350 5505
rect 3250 5415 3260 5495
rect 3340 5415 3350 5495
rect 3250 5405 3350 5415
rect 3450 5495 3550 5505
rect 3450 5415 3460 5495
rect 3540 5415 3550 5495
rect 3450 5405 3550 5415
rect 3650 5495 3750 5505
rect 3650 5415 3660 5495
rect 3740 5415 3750 5495
rect 3650 5405 3750 5415
rect 3850 5495 3950 5505
rect 3850 5415 3860 5495
rect 3940 5415 3950 5495
rect 3850 5405 3950 5415
rect 4050 5495 4150 5505
rect 4050 5415 4060 5495
rect 4140 5415 4150 5495
rect 4050 5405 4150 5415
rect 4250 5495 4350 5505
rect 4250 5415 4260 5495
rect 4340 5415 4350 5495
rect 4250 5405 4350 5415
rect 4450 5495 4550 5505
rect 4450 5415 4460 5495
rect 4540 5415 4550 5495
rect 4450 5405 4550 5415
rect 4650 5495 4750 5505
rect 4650 5415 4660 5495
rect 4740 5415 4750 5495
rect 4650 5405 4750 5415
rect 4850 5495 4950 5505
rect 4850 5415 4860 5495
rect 4940 5415 4950 5495
rect 4850 5405 4950 5415
rect 5050 5495 5150 5505
rect 5050 5415 5060 5495
rect 5140 5415 5150 5495
rect 5050 5405 5150 5415
rect 5250 5495 5350 5505
rect 5250 5415 5260 5495
rect 5340 5415 5350 5495
rect 5250 5405 5350 5415
rect 5450 5495 5550 5505
rect 5450 5415 5460 5495
rect 5540 5415 5550 5495
rect 5450 5405 5550 5415
rect 5650 5495 5750 5505
rect 5650 5415 5660 5495
rect 5740 5415 5750 5495
rect 5650 5405 5750 5415
rect 5850 5495 5950 5505
rect 5850 5415 5860 5495
rect 5940 5415 5950 5495
rect 5850 5405 5950 5415
rect 6050 5495 6150 5505
rect 6050 5415 6060 5495
rect 6140 5415 6150 5495
rect 6050 5405 6150 5415
rect 6250 5495 6350 5505
rect 6250 5415 6260 5495
rect 6340 5415 6350 5495
rect 6250 5405 6350 5415
rect 6450 5495 6550 5505
rect 6450 5415 6460 5495
rect 6540 5415 6550 5495
rect 6450 5405 6550 5415
rect -115 5320 -85 5405
rect 85 5320 115 5405
rect 285 5320 315 5405
rect 485 5320 515 5405
rect 685 5320 715 5405
rect 885 5320 915 5405
rect 1085 5320 1115 5405
rect 1285 5320 1315 5405
rect 1485 5320 1515 5405
rect 1685 5320 1715 5405
rect 1885 5320 1915 5405
rect 2085 5320 2115 5405
rect 2285 5320 2315 5405
rect 2485 5320 2515 5405
rect 2685 5320 2715 5405
rect 2885 5320 2915 5405
rect 3085 5320 3115 5405
rect 3285 5320 3315 5405
rect 3485 5320 3515 5405
rect 3685 5320 3715 5405
rect 3885 5320 3915 5405
rect 4085 5320 4115 5405
rect 4285 5320 4315 5405
rect 4485 5320 4515 5405
rect 4685 5320 4715 5405
rect 4885 5320 4915 5405
rect 5085 5320 5115 5405
rect 5285 5320 5315 5405
rect 5485 5320 5515 5405
rect 5685 5320 5715 5405
rect 5885 5320 5915 5405
rect 6085 5320 6115 5405
rect 6285 5320 6315 5405
rect 6485 5320 6515 5405
rect -150 5310 -50 5320
rect -150 5230 -140 5310
rect -60 5230 -50 5310
rect -150 5220 -50 5230
rect 50 5310 150 5320
rect 50 5230 60 5310
rect 140 5230 150 5310
rect 50 5220 150 5230
rect 250 5310 350 5320
rect 250 5230 260 5310
rect 340 5230 350 5310
rect 250 5220 350 5230
rect 450 5310 550 5320
rect 450 5230 460 5310
rect 540 5230 550 5310
rect 450 5220 550 5230
rect 650 5310 750 5320
rect 650 5230 660 5310
rect 740 5230 750 5310
rect 650 5220 750 5230
rect 850 5310 950 5320
rect 850 5230 860 5310
rect 940 5230 950 5310
rect 850 5220 950 5230
rect 1050 5310 1150 5320
rect 1050 5230 1060 5310
rect 1140 5230 1150 5310
rect 1050 5220 1150 5230
rect 1250 5310 1350 5320
rect 1250 5230 1260 5310
rect 1340 5230 1350 5310
rect 1250 5220 1350 5230
rect 1450 5310 1550 5320
rect 1450 5230 1460 5310
rect 1540 5230 1550 5310
rect 1450 5220 1550 5230
rect 1650 5310 1750 5320
rect 1650 5230 1660 5310
rect 1740 5230 1750 5310
rect 1650 5220 1750 5230
rect 1850 5310 1950 5320
rect 1850 5230 1860 5310
rect 1940 5230 1950 5310
rect 1850 5220 1950 5230
rect 2050 5310 2150 5320
rect 2050 5230 2060 5310
rect 2140 5230 2150 5310
rect 2050 5220 2150 5230
rect 2250 5310 2350 5320
rect 2250 5230 2260 5310
rect 2340 5230 2350 5310
rect 2250 5220 2350 5230
rect 2450 5310 2550 5320
rect 2450 5230 2460 5310
rect 2540 5230 2550 5310
rect 2450 5220 2550 5230
rect 2650 5310 2750 5320
rect 2650 5230 2660 5310
rect 2740 5230 2750 5310
rect 2650 5220 2750 5230
rect 2850 5310 2950 5320
rect 2850 5230 2860 5310
rect 2940 5230 2950 5310
rect 2850 5220 2950 5230
rect 3050 5310 3150 5320
rect 3050 5230 3060 5310
rect 3140 5230 3150 5310
rect 3050 5220 3150 5230
rect 3250 5310 3350 5320
rect 3250 5230 3260 5310
rect 3340 5230 3350 5310
rect 3250 5220 3350 5230
rect 3450 5310 3550 5320
rect 3450 5230 3460 5310
rect 3540 5230 3550 5310
rect 3450 5220 3550 5230
rect 3650 5310 3750 5320
rect 3650 5230 3660 5310
rect 3740 5230 3750 5310
rect 3650 5220 3750 5230
rect 3850 5310 3950 5320
rect 3850 5230 3860 5310
rect 3940 5230 3950 5310
rect 3850 5220 3950 5230
rect 4050 5310 4150 5320
rect 4050 5230 4060 5310
rect 4140 5230 4150 5310
rect 4050 5220 4150 5230
rect 4250 5310 4350 5320
rect 4250 5230 4260 5310
rect 4340 5230 4350 5310
rect 4250 5220 4350 5230
rect 4450 5310 4550 5320
rect 4450 5230 4460 5310
rect 4540 5230 4550 5310
rect 4450 5220 4550 5230
rect 4650 5310 4750 5320
rect 4650 5230 4660 5310
rect 4740 5230 4750 5310
rect 4650 5220 4750 5230
rect 4850 5310 4950 5320
rect 4850 5230 4860 5310
rect 4940 5230 4950 5310
rect 4850 5220 4950 5230
rect 5050 5310 5150 5320
rect 5050 5230 5060 5310
rect 5140 5230 5150 5310
rect 5050 5220 5150 5230
rect 5250 5310 5350 5320
rect 5250 5230 5260 5310
rect 5340 5230 5350 5310
rect 5250 5220 5350 5230
rect 5450 5310 5550 5320
rect 5450 5230 5460 5310
rect 5540 5230 5550 5310
rect 5450 5220 5550 5230
rect 5650 5310 5750 5320
rect 5650 5230 5660 5310
rect 5740 5230 5750 5310
rect 5650 5220 5750 5230
rect 5850 5310 5950 5320
rect 5850 5230 5860 5310
rect 5940 5230 5950 5310
rect 5850 5220 5950 5230
rect 6050 5310 6150 5320
rect 6050 5230 6060 5310
rect 6140 5230 6150 5310
rect 6050 5220 6150 5230
rect 6250 5310 6350 5320
rect 6250 5230 6260 5310
rect 6340 5230 6350 5310
rect 6250 5220 6350 5230
rect 6450 5310 6550 5320
rect 6450 5230 6460 5310
rect 6540 5230 6550 5310
rect 6450 5220 6550 5230
rect -115 5135 -85 5220
rect 85 5135 115 5220
rect 285 5135 315 5220
rect 485 5135 515 5220
rect 685 5135 715 5220
rect 885 5135 915 5220
rect 1085 5135 1115 5220
rect 1285 5135 1315 5220
rect 1485 5135 1515 5220
rect 1685 5135 1715 5220
rect 1885 5135 1915 5220
rect 2085 5135 2115 5220
rect 2285 5135 2315 5220
rect 2485 5135 2515 5220
rect 2685 5135 2715 5220
rect 2885 5135 2915 5220
rect 3085 5135 3115 5220
rect 3285 5135 3315 5220
rect 3485 5135 3515 5220
rect 3685 5135 3715 5220
rect 3885 5135 3915 5220
rect 4085 5135 4115 5220
rect 4285 5135 4315 5220
rect 4485 5135 4515 5220
rect 4685 5135 4715 5220
rect 4885 5135 4915 5220
rect 5085 5135 5115 5220
rect 5285 5135 5315 5220
rect 5485 5135 5515 5220
rect 5685 5135 5715 5220
rect 5885 5135 5915 5220
rect 6085 5135 6115 5220
rect 6285 5135 6315 5220
rect 6485 5135 6515 5220
rect -150 5125 -50 5135
rect -150 5045 -140 5125
rect -60 5045 -50 5125
rect -150 5035 -50 5045
rect 50 5125 150 5135
rect 50 5045 60 5125
rect 140 5045 150 5125
rect 50 5035 150 5045
rect 250 5125 350 5135
rect 250 5045 260 5125
rect 340 5045 350 5125
rect 250 5035 350 5045
rect 450 5125 550 5135
rect 450 5045 460 5125
rect 540 5045 550 5125
rect 450 5035 550 5045
rect 650 5125 750 5135
rect 650 5045 660 5125
rect 740 5045 750 5125
rect 650 5035 750 5045
rect 850 5125 950 5135
rect 850 5045 860 5125
rect 940 5045 950 5125
rect 850 5035 950 5045
rect 1050 5125 1150 5135
rect 1050 5045 1060 5125
rect 1140 5045 1150 5125
rect 1050 5035 1150 5045
rect 1250 5125 1350 5135
rect 1250 5045 1260 5125
rect 1340 5045 1350 5125
rect 1250 5035 1350 5045
rect 1450 5125 1550 5135
rect 1450 5045 1460 5125
rect 1540 5045 1550 5125
rect 1450 5035 1550 5045
rect 1650 5125 1750 5135
rect 1650 5045 1660 5125
rect 1740 5045 1750 5125
rect 1650 5035 1750 5045
rect 1850 5125 1950 5135
rect 1850 5045 1860 5125
rect 1940 5045 1950 5125
rect 1850 5035 1950 5045
rect 2050 5125 2150 5135
rect 2050 5045 2060 5125
rect 2140 5045 2150 5125
rect 2050 5035 2150 5045
rect 2250 5125 2350 5135
rect 2250 5045 2260 5125
rect 2340 5045 2350 5125
rect 2250 5035 2350 5045
rect 2450 5125 2550 5135
rect 2450 5045 2460 5125
rect 2540 5045 2550 5125
rect 2450 5035 2550 5045
rect 2650 5125 2750 5135
rect 2650 5045 2660 5125
rect 2740 5045 2750 5125
rect 2650 5035 2750 5045
rect 2850 5125 2950 5135
rect 2850 5045 2860 5125
rect 2940 5045 2950 5125
rect 2850 5035 2950 5045
rect 3050 5125 3150 5135
rect 3050 5045 3060 5125
rect 3140 5045 3150 5125
rect 3050 5035 3150 5045
rect 3250 5125 3350 5135
rect 3250 5045 3260 5125
rect 3340 5045 3350 5125
rect 3250 5035 3350 5045
rect 3450 5125 3550 5135
rect 3450 5045 3460 5125
rect 3540 5045 3550 5125
rect 3450 5035 3550 5045
rect 3650 5125 3750 5135
rect 3650 5045 3660 5125
rect 3740 5045 3750 5125
rect 3650 5035 3750 5045
rect 3850 5125 3950 5135
rect 3850 5045 3860 5125
rect 3940 5045 3950 5125
rect 3850 5035 3950 5045
rect 4050 5125 4150 5135
rect 4050 5045 4060 5125
rect 4140 5045 4150 5125
rect 4050 5035 4150 5045
rect 4250 5125 4350 5135
rect 4250 5045 4260 5125
rect 4340 5045 4350 5125
rect 4250 5035 4350 5045
rect 4450 5125 4550 5135
rect 4450 5045 4460 5125
rect 4540 5045 4550 5125
rect 4450 5035 4550 5045
rect 4650 5125 4750 5135
rect 4650 5045 4660 5125
rect 4740 5045 4750 5125
rect 4650 5035 4750 5045
rect 4850 5125 4950 5135
rect 4850 5045 4860 5125
rect 4940 5045 4950 5125
rect 4850 5035 4950 5045
rect 5050 5125 5150 5135
rect 5050 5045 5060 5125
rect 5140 5045 5150 5125
rect 5050 5035 5150 5045
rect 5250 5125 5350 5135
rect 5250 5045 5260 5125
rect 5340 5045 5350 5125
rect 5250 5035 5350 5045
rect 5450 5125 5550 5135
rect 5450 5045 5460 5125
rect 5540 5045 5550 5125
rect 5450 5035 5550 5045
rect 5650 5125 5750 5135
rect 5650 5045 5660 5125
rect 5740 5045 5750 5125
rect 5650 5035 5750 5045
rect 5850 5125 5950 5135
rect 5850 5045 5860 5125
rect 5940 5045 5950 5125
rect 5850 5035 5950 5045
rect 6050 5125 6150 5135
rect 6050 5045 6060 5125
rect 6140 5045 6150 5125
rect 6050 5035 6150 5045
rect 6250 5125 6350 5135
rect 6250 5045 6260 5125
rect 6340 5045 6350 5125
rect 6250 5035 6350 5045
rect 6450 5125 6550 5135
rect 6450 5045 6460 5125
rect 6540 5045 6550 5125
rect 6450 5035 6550 5045
rect -115 4950 -85 5035
rect 85 4950 115 5035
rect 285 4950 315 5035
rect 485 4950 515 5035
rect 685 4950 715 5035
rect 885 4950 915 5035
rect 1085 4950 1115 5035
rect 1285 4950 1315 5035
rect 1485 4950 1515 5035
rect 1685 4950 1715 5035
rect 1885 4950 1915 5035
rect 2085 4950 2115 5035
rect 2285 4950 2315 5035
rect 2485 4950 2515 5035
rect 2685 4950 2715 5035
rect 2885 4950 2915 5035
rect 3085 4950 3115 5035
rect 3285 4950 3315 5035
rect 3485 4950 3515 5035
rect 3685 4950 3715 5035
rect 3885 4950 3915 5035
rect 4085 4950 4115 5035
rect 4285 4950 4315 5035
rect 4485 4950 4515 5035
rect 4685 4950 4715 5035
rect 4885 4950 4915 5035
rect 5085 4950 5115 5035
rect 5285 4950 5315 5035
rect 5485 4950 5515 5035
rect 5685 4950 5715 5035
rect 5885 4950 5915 5035
rect 6085 4950 6115 5035
rect 6285 4950 6315 5035
rect 6485 4950 6515 5035
rect -150 4940 -50 4950
rect -150 4860 -140 4940
rect -60 4860 -50 4940
rect -150 4850 -50 4860
rect 50 4940 150 4950
rect 50 4860 60 4940
rect 140 4860 150 4940
rect 50 4850 150 4860
rect 250 4940 350 4950
rect 250 4860 260 4940
rect 340 4860 350 4940
rect 250 4850 350 4860
rect 450 4940 550 4950
rect 450 4860 460 4940
rect 540 4860 550 4940
rect 450 4850 550 4860
rect 650 4940 750 4950
rect 650 4860 660 4940
rect 740 4860 750 4940
rect 650 4850 750 4860
rect 850 4940 950 4950
rect 850 4860 860 4940
rect 940 4860 950 4940
rect 850 4850 950 4860
rect 1050 4940 1150 4950
rect 1050 4860 1060 4940
rect 1140 4860 1150 4940
rect 1050 4850 1150 4860
rect 1250 4940 1350 4950
rect 1250 4860 1260 4940
rect 1340 4860 1350 4940
rect 1250 4850 1350 4860
rect 1450 4940 1550 4950
rect 1450 4860 1460 4940
rect 1540 4860 1550 4940
rect 1450 4850 1550 4860
rect 1650 4940 1750 4950
rect 1650 4860 1660 4940
rect 1740 4860 1750 4940
rect 1650 4850 1750 4860
rect 1850 4940 1950 4950
rect 1850 4860 1860 4940
rect 1940 4860 1950 4940
rect 1850 4850 1950 4860
rect 2050 4940 2150 4950
rect 2050 4860 2060 4940
rect 2140 4860 2150 4940
rect 2050 4850 2150 4860
rect 2250 4940 2350 4950
rect 2250 4860 2260 4940
rect 2340 4860 2350 4940
rect 2250 4850 2350 4860
rect 2450 4940 2550 4950
rect 2450 4860 2460 4940
rect 2540 4860 2550 4940
rect 2450 4850 2550 4860
rect 2650 4940 2750 4950
rect 2650 4860 2660 4940
rect 2740 4860 2750 4940
rect 2650 4850 2750 4860
rect 2850 4940 2950 4950
rect 2850 4860 2860 4940
rect 2940 4860 2950 4940
rect 2850 4850 2950 4860
rect 3050 4940 3150 4950
rect 3050 4860 3060 4940
rect 3140 4860 3150 4940
rect 3050 4850 3150 4860
rect 3250 4940 3350 4950
rect 3250 4860 3260 4940
rect 3340 4860 3350 4940
rect 3250 4850 3350 4860
rect 3450 4940 3550 4950
rect 3450 4860 3460 4940
rect 3540 4860 3550 4940
rect 3450 4850 3550 4860
rect 3650 4940 3750 4950
rect 3650 4860 3660 4940
rect 3740 4860 3750 4940
rect 3650 4850 3750 4860
rect 3850 4940 3950 4950
rect 3850 4860 3860 4940
rect 3940 4860 3950 4940
rect 3850 4850 3950 4860
rect 4050 4940 4150 4950
rect 4050 4860 4060 4940
rect 4140 4860 4150 4940
rect 4050 4850 4150 4860
rect 4250 4940 4350 4950
rect 4250 4860 4260 4940
rect 4340 4860 4350 4940
rect 4250 4850 4350 4860
rect 4450 4940 4550 4950
rect 4450 4860 4460 4940
rect 4540 4860 4550 4940
rect 4450 4850 4550 4860
rect 4650 4940 4750 4950
rect 4650 4860 4660 4940
rect 4740 4860 4750 4940
rect 4650 4850 4750 4860
rect 4850 4940 4950 4950
rect 4850 4860 4860 4940
rect 4940 4860 4950 4940
rect 4850 4850 4950 4860
rect 5050 4940 5150 4950
rect 5050 4860 5060 4940
rect 5140 4860 5150 4940
rect 5050 4850 5150 4860
rect 5250 4940 5350 4950
rect 5250 4860 5260 4940
rect 5340 4860 5350 4940
rect 5250 4850 5350 4860
rect 5450 4940 5550 4950
rect 5450 4860 5460 4940
rect 5540 4860 5550 4940
rect 5450 4850 5550 4860
rect 5650 4940 5750 4950
rect 5650 4860 5660 4940
rect 5740 4860 5750 4940
rect 5650 4850 5750 4860
rect 5850 4940 5950 4950
rect 5850 4860 5860 4940
rect 5940 4860 5950 4940
rect 5850 4850 5950 4860
rect 6050 4940 6150 4950
rect 6050 4860 6060 4940
rect 6140 4860 6150 4940
rect 6050 4850 6150 4860
rect 6250 4940 6350 4950
rect 6250 4860 6260 4940
rect 6340 4860 6350 4940
rect 6250 4850 6350 4860
rect 6450 4940 6550 4950
rect 6450 4860 6460 4940
rect 6540 4860 6550 4940
rect 6450 4850 6550 4860
rect -115 4765 -85 4850
rect 85 4765 115 4850
rect 285 4765 315 4850
rect 485 4765 515 4850
rect 685 4765 715 4850
rect 885 4765 915 4850
rect 1085 4765 1115 4850
rect 1285 4765 1315 4850
rect 1485 4765 1515 4850
rect 1685 4765 1715 4850
rect 1885 4765 1915 4850
rect 2085 4765 2115 4850
rect 2285 4765 2315 4850
rect 2485 4765 2515 4850
rect 2685 4765 2715 4850
rect 2885 4765 2915 4850
rect 3085 4765 3115 4850
rect 3285 4765 3315 4850
rect 3485 4765 3515 4850
rect 3685 4765 3715 4850
rect 3885 4765 3915 4850
rect 4085 4765 4115 4850
rect 4285 4765 4315 4850
rect 4485 4765 4515 4850
rect 4685 4765 4715 4850
rect 4885 4765 4915 4850
rect 5085 4765 5115 4850
rect 5285 4765 5315 4850
rect 5485 4765 5515 4850
rect 5685 4765 5715 4850
rect 5885 4765 5915 4850
rect 6085 4765 6115 4850
rect 6285 4765 6315 4850
rect 6485 4765 6515 4850
rect -150 4755 -50 4765
rect -150 4675 -140 4755
rect -60 4675 -50 4755
rect -150 4665 -50 4675
rect 50 4755 150 4765
rect 50 4675 60 4755
rect 140 4675 150 4755
rect 50 4665 150 4675
rect 250 4755 350 4765
rect 250 4675 260 4755
rect 340 4675 350 4755
rect 250 4665 350 4675
rect 450 4755 550 4765
rect 450 4675 460 4755
rect 540 4675 550 4755
rect 450 4665 550 4675
rect 650 4755 750 4765
rect 650 4675 660 4755
rect 740 4675 750 4755
rect 650 4665 750 4675
rect 850 4755 950 4765
rect 850 4675 860 4755
rect 940 4675 950 4755
rect 850 4665 950 4675
rect 1050 4755 1150 4765
rect 1050 4675 1060 4755
rect 1140 4675 1150 4755
rect 1050 4665 1150 4675
rect 1250 4755 1350 4765
rect 1250 4675 1260 4755
rect 1340 4675 1350 4755
rect 1250 4665 1350 4675
rect 1450 4755 1550 4765
rect 1450 4675 1460 4755
rect 1540 4675 1550 4755
rect 1450 4665 1550 4675
rect 1650 4755 1750 4765
rect 1650 4675 1660 4755
rect 1740 4675 1750 4755
rect 1650 4665 1750 4675
rect 1850 4755 1950 4765
rect 1850 4675 1860 4755
rect 1940 4675 1950 4755
rect 1850 4665 1950 4675
rect 2050 4755 2150 4765
rect 2050 4675 2060 4755
rect 2140 4675 2150 4755
rect 2050 4665 2150 4675
rect 2250 4755 2350 4765
rect 2250 4675 2260 4755
rect 2340 4675 2350 4755
rect 2250 4665 2350 4675
rect 2450 4755 2550 4765
rect 2450 4675 2460 4755
rect 2540 4675 2550 4755
rect 2450 4665 2550 4675
rect 2650 4755 2750 4765
rect 2650 4675 2660 4755
rect 2740 4675 2750 4755
rect 2650 4665 2750 4675
rect 2850 4755 2950 4765
rect 2850 4675 2860 4755
rect 2940 4675 2950 4755
rect 2850 4665 2950 4675
rect 3050 4755 3150 4765
rect 3050 4675 3060 4755
rect 3140 4675 3150 4755
rect 3050 4665 3150 4675
rect 3250 4755 3350 4765
rect 3250 4675 3260 4755
rect 3340 4675 3350 4755
rect 3250 4665 3350 4675
rect 3450 4755 3550 4765
rect 3450 4675 3460 4755
rect 3540 4675 3550 4755
rect 3450 4665 3550 4675
rect 3650 4755 3750 4765
rect 3650 4675 3660 4755
rect 3740 4675 3750 4755
rect 3650 4665 3750 4675
rect 3850 4755 3950 4765
rect 3850 4675 3860 4755
rect 3940 4675 3950 4755
rect 3850 4665 3950 4675
rect 4050 4755 4150 4765
rect 4050 4675 4060 4755
rect 4140 4675 4150 4755
rect 4050 4665 4150 4675
rect 4250 4755 4350 4765
rect 4250 4675 4260 4755
rect 4340 4675 4350 4755
rect 4250 4665 4350 4675
rect 4450 4755 4550 4765
rect 4450 4675 4460 4755
rect 4540 4675 4550 4755
rect 4450 4665 4550 4675
rect 4650 4755 4750 4765
rect 4650 4675 4660 4755
rect 4740 4675 4750 4755
rect 4650 4665 4750 4675
rect 4850 4755 4950 4765
rect 4850 4675 4860 4755
rect 4940 4675 4950 4755
rect 4850 4665 4950 4675
rect 5050 4755 5150 4765
rect 5050 4675 5060 4755
rect 5140 4675 5150 4755
rect 5050 4665 5150 4675
rect 5250 4755 5350 4765
rect 5250 4675 5260 4755
rect 5340 4675 5350 4755
rect 5250 4665 5350 4675
rect 5450 4755 5550 4765
rect 5450 4675 5460 4755
rect 5540 4675 5550 4755
rect 5450 4665 5550 4675
rect 5650 4755 5750 4765
rect 5650 4675 5660 4755
rect 5740 4675 5750 4755
rect 5650 4665 5750 4675
rect 5850 4755 5950 4765
rect 5850 4675 5860 4755
rect 5940 4675 5950 4755
rect 5850 4665 5950 4675
rect 6050 4755 6150 4765
rect 6050 4675 6060 4755
rect 6140 4675 6150 4755
rect 6050 4665 6150 4675
rect 6250 4755 6350 4765
rect 6250 4675 6260 4755
rect 6340 4675 6350 4755
rect 6250 4665 6350 4675
rect 6450 4755 6550 4765
rect 6450 4675 6460 4755
rect 6540 4675 6550 4755
rect 6450 4665 6550 4675
rect -115 4580 -85 4665
rect 85 4580 115 4665
rect 285 4580 315 4665
rect 485 4580 515 4665
rect 685 4580 715 4665
rect 885 4580 915 4665
rect 1085 4580 1115 4665
rect 1285 4580 1315 4665
rect 1485 4580 1515 4665
rect 1685 4580 1715 4665
rect 1885 4580 1915 4665
rect 2085 4580 2115 4665
rect 2285 4580 2315 4665
rect 2485 4580 2515 4665
rect 2685 4580 2715 4665
rect 2885 4580 2915 4665
rect 3085 4580 3115 4665
rect 3285 4580 3315 4665
rect 3485 4580 3515 4665
rect 3685 4580 3715 4665
rect 3885 4580 3915 4665
rect 4085 4580 4115 4665
rect 4285 4580 4315 4665
rect 4485 4580 4515 4665
rect 4685 4580 4715 4665
rect 4885 4580 4915 4665
rect 5085 4580 5115 4665
rect 5285 4580 5315 4665
rect 5485 4580 5515 4665
rect 5685 4580 5715 4665
rect 5885 4580 5915 4665
rect 6085 4580 6115 4665
rect 6285 4580 6315 4665
rect 6485 4580 6515 4665
rect -150 4570 -50 4580
rect -150 4490 -140 4570
rect -60 4490 -50 4570
rect -150 4480 -50 4490
rect 50 4570 150 4580
rect 50 4490 60 4570
rect 140 4490 150 4570
rect 50 4480 150 4490
rect 250 4570 350 4580
rect 250 4490 260 4570
rect 340 4490 350 4570
rect 250 4480 350 4490
rect 450 4570 550 4580
rect 450 4490 460 4570
rect 540 4490 550 4570
rect 450 4480 550 4490
rect 650 4570 750 4580
rect 650 4490 660 4570
rect 740 4490 750 4570
rect 650 4480 750 4490
rect 850 4570 950 4580
rect 850 4490 860 4570
rect 940 4490 950 4570
rect 850 4480 950 4490
rect 1050 4570 1150 4580
rect 1050 4490 1060 4570
rect 1140 4490 1150 4570
rect 1050 4480 1150 4490
rect 1250 4570 1350 4580
rect 1250 4490 1260 4570
rect 1340 4490 1350 4570
rect 1250 4480 1350 4490
rect 1450 4570 1550 4580
rect 1450 4490 1460 4570
rect 1540 4490 1550 4570
rect 1450 4480 1550 4490
rect 1650 4570 1750 4580
rect 1650 4490 1660 4570
rect 1740 4490 1750 4570
rect 1650 4480 1750 4490
rect 1850 4570 1950 4580
rect 1850 4490 1860 4570
rect 1940 4490 1950 4570
rect 1850 4480 1950 4490
rect 2050 4570 2150 4580
rect 2050 4490 2060 4570
rect 2140 4490 2150 4570
rect 2050 4480 2150 4490
rect 2250 4570 2350 4580
rect 2250 4490 2260 4570
rect 2340 4490 2350 4570
rect 2250 4480 2350 4490
rect 2450 4570 2550 4580
rect 2450 4490 2460 4570
rect 2540 4490 2550 4570
rect 2450 4480 2550 4490
rect 2650 4570 2750 4580
rect 2650 4490 2660 4570
rect 2740 4490 2750 4570
rect 2650 4480 2750 4490
rect 2850 4570 2950 4580
rect 2850 4490 2860 4570
rect 2940 4490 2950 4570
rect 2850 4480 2950 4490
rect 3050 4570 3150 4580
rect 3050 4490 3060 4570
rect 3140 4490 3150 4570
rect 3050 4480 3150 4490
rect 3250 4570 3350 4580
rect 3250 4490 3260 4570
rect 3340 4490 3350 4570
rect 3250 4480 3350 4490
rect 3450 4570 3550 4580
rect 3450 4490 3460 4570
rect 3540 4490 3550 4570
rect 3450 4480 3550 4490
rect 3650 4570 3750 4580
rect 3650 4490 3660 4570
rect 3740 4490 3750 4570
rect 3650 4480 3750 4490
rect 3850 4570 3950 4580
rect 3850 4490 3860 4570
rect 3940 4490 3950 4570
rect 3850 4480 3950 4490
rect 4050 4570 4150 4580
rect 4050 4490 4060 4570
rect 4140 4490 4150 4570
rect 4050 4480 4150 4490
rect 4250 4570 4350 4580
rect 4250 4490 4260 4570
rect 4340 4490 4350 4570
rect 4250 4480 4350 4490
rect 4450 4570 4550 4580
rect 4450 4490 4460 4570
rect 4540 4490 4550 4570
rect 4450 4480 4550 4490
rect 4650 4570 4750 4580
rect 4650 4490 4660 4570
rect 4740 4490 4750 4570
rect 4650 4480 4750 4490
rect 4850 4570 4950 4580
rect 4850 4490 4860 4570
rect 4940 4490 4950 4570
rect 4850 4480 4950 4490
rect 5050 4570 5150 4580
rect 5050 4490 5060 4570
rect 5140 4490 5150 4570
rect 5050 4480 5150 4490
rect 5250 4570 5350 4580
rect 5250 4490 5260 4570
rect 5340 4490 5350 4570
rect 5250 4480 5350 4490
rect 5450 4570 5550 4580
rect 5450 4490 5460 4570
rect 5540 4490 5550 4570
rect 5450 4480 5550 4490
rect 5650 4570 5750 4580
rect 5650 4490 5660 4570
rect 5740 4490 5750 4570
rect 5650 4480 5750 4490
rect 5850 4570 5950 4580
rect 5850 4490 5860 4570
rect 5940 4490 5950 4570
rect 5850 4480 5950 4490
rect 6050 4570 6150 4580
rect 6050 4490 6060 4570
rect 6140 4490 6150 4570
rect 6050 4480 6150 4490
rect 6250 4570 6350 4580
rect 6250 4490 6260 4570
rect 6340 4490 6350 4570
rect 6250 4480 6350 4490
rect 6450 4570 6550 4580
rect 6450 4490 6460 4570
rect 6540 4490 6550 4570
rect 6450 4480 6550 4490
rect -115 4395 -85 4480
rect 85 4395 115 4480
rect 285 4395 315 4480
rect 485 4395 515 4480
rect 685 4395 715 4480
rect 885 4395 915 4480
rect 1085 4395 1115 4480
rect 1285 4395 1315 4480
rect 1485 4395 1515 4480
rect 1685 4395 1715 4480
rect 1885 4395 1915 4480
rect 2085 4395 2115 4480
rect 2285 4395 2315 4480
rect 2485 4395 2515 4480
rect 2685 4395 2715 4480
rect 2885 4395 2915 4480
rect 3085 4395 3115 4480
rect 3285 4395 3315 4480
rect 3485 4395 3515 4480
rect 3685 4395 3715 4480
rect 3885 4395 3915 4480
rect 4085 4395 4115 4480
rect 4285 4395 4315 4480
rect 4485 4395 4515 4480
rect 4685 4395 4715 4480
rect 4885 4395 4915 4480
rect 5085 4395 5115 4480
rect 5285 4395 5315 4480
rect 5485 4395 5515 4480
rect 5685 4395 5715 4480
rect 5885 4395 5915 4480
rect 6085 4395 6115 4480
rect 6285 4395 6315 4480
rect 6485 4395 6515 4480
rect -150 4385 -50 4395
rect -150 4305 -140 4385
rect -60 4305 -50 4385
rect -150 4295 -50 4305
rect 50 4385 150 4395
rect 50 4305 60 4385
rect 140 4305 150 4385
rect 50 4295 150 4305
rect 250 4385 350 4395
rect 250 4305 260 4385
rect 340 4305 350 4385
rect 250 4295 350 4305
rect 450 4385 550 4395
rect 450 4305 460 4385
rect 540 4305 550 4385
rect 450 4295 550 4305
rect 650 4385 750 4395
rect 650 4305 660 4385
rect 740 4305 750 4385
rect 650 4295 750 4305
rect 850 4385 950 4395
rect 850 4305 860 4385
rect 940 4305 950 4385
rect 850 4295 950 4305
rect 1050 4385 1150 4395
rect 1050 4305 1060 4385
rect 1140 4305 1150 4385
rect 1050 4295 1150 4305
rect 1250 4385 1350 4395
rect 1250 4305 1260 4385
rect 1340 4305 1350 4385
rect 1250 4295 1350 4305
rect 1450 4385 1550 4395
rect 1450 4305 1460 4385
rect 1540 4305 1550 4385
rect 1450 4295 1550 4305
rect 1650 4385 1750 4395
rect 1650 4305 1660 4385
rect 1740 4305 1750 4385
rect 1650 4295 1750 4305
rect 1850 4385 1950 4395
rect 1850 4305 1860 4385
rect 1940 4305 1950 4385
rect 1850 4295 1950 4305
rect 2050 4385 2150 4395
rect 2050 4305 2060 4385
rect 2140 4305 2150 4385
rect 2050 4295 2150 4305
rect 2250 4385 2350 4395
rect 2250 4305 2260 4385
rect 2340 4305 2350 4385
rect 2250 4295 2350 4305
rect 2450 4385 2550 4395
rect 2450 4305 2460 4385
rect 2540 4305 2550 4385
rect 2450 4295 2550 4305
rect 2650 4385 2750 4395
rect 2650 4305 2660 4385
rect 2740 4305 2750 4385
rect 2650 4295 2750 4305
rect 2850 4385 2950 4395
rect 2850 4305 2860 4385
rect 2940 4305 2950 4385
rect 2850 4295 2950 4305
rect 3050 4385 3150 4395
rect 3050 4305 3060 4385
rect 3140 4305 3150 4385
rect 3050 4295 3150 4305
rect 3250 4385 3350 4395
rect 3250 4305 3260 4385
rect 3340 4305 3350 4385
rect 3250 4295 3350 4305
rect 3450 4385 3550 4395
rect 3450 4305 3460 4385
rect 3540 4305 3550 4385
rect 3450 4295 3550 4305
rect 3650 4385 3750 4395
rect 3650 4305 3660 4385
rect 3740 4305 3750 4385
rect 3650 4295 3750 4305
rect 3850 4385 3950 4395
rect 3850 4305 3860 4385
rect 3940 4305 3950 4385
rect 3850 4295 3950 4305
rect 4050 4385 4150 4395
rect 4050 4305 4060 4385
rect 4140 4305 4150 4385
rect 4050 4295 4150 4305
rect 4250 4385 4350 4395
rect 4250 4305 4260 4385
rect 4340 4305 4350 4385
rect 4250 4295 4350 4305
rect 4450 4385 4550 4395
rect 4450 4305 4460 4385
rect 4540 4305 4550 4385
rect 4450 4295 4550 4305
rect 4650 4385 4750 4395
rect 4650 4305 4660 4385
rect 4740 4305 4750 4385
rect 4650 4295 4750 4305
rect 4850 4385 4950 4395
rect 4850 4305 4860 4385
rect 4940 4305 4950 4385
rect 4850 4295 4950 4305
rect 5050 4385 5150 4395
rect 5050 4305 5060 4385
rect 5140 4305 5150 4385
rect 5050 4295 5150 4305
rect 5250 4385 5350 4395
rect 5250 4305 5260 4385
rect 5340 4305 5350 4385
rect 5250 4295 5350 4305
rect 5450 4385 5550 4395
rect 5450 4305 5460 4385
rect 5540 4305 5550 4385
rect 5450 4295 5550 4305
rect 5650 4385 5750 4395
rect 5650 4305 5660 4385
rect 5740 4305 5750 4385
rect 5650 4295 5750 4305
rect 5850 4385 5950 4395
rect 5850 4305 5860 4385
rect 5940 4305 5950 4385
rect 5850 4295 5950 4305
rect 6050 4385 6150 4395
rect 6050 4305 6060 4385
rect 6140 4305 6150 4385
rect 6050 4295 6150 4305
rect 6250 4385 6350 4395
rect 6250 4305 6260 4385
rect 6340 4305 6350 4385
rect 6250 4295 6350 4305
rect 6450 4385 6550 4395
rect 6450 4305 6460 4385
rect 6540 4305 6550 4385
rect 6450 4295 6550 4305
rect -115 4210 -85 4295
rect 85 4210 115 4295
rect 285 4210 315 4295
rect 485 4210 515 4295
rect 685 4210 715 4295
rect 885 4210 915 4295
rect 1085 4210 1115 4295
rect 1285 4210 1315 4295
rect 1485 4210 1515 4295
rect 1685 4210 1715 4295
rect 1885 4210 1915 4295
rect 2085 4210 2115 4295
rect 2285 4210 2315 4295
rect 2485 4210 2515 4295
rect 2685 4210 2715 4295
rect 2885 4210 2915 4295
rect 3085 4210 3115 4295
rect 3285 4210 3315 4295
rect 3485 4210 3515 4295
rect 3685 4210 3715 4295
rect 3885 4210 3915 4295
rect 4085 4210 4115 4295
rect 4285 4210 4315 4295
rect 4485 4210 4515 4295
rect 4685 4210 4715 4295
rect 4885 4210 4915 4295
rect 5085 4210 5115 4295
rect 5285 4210 5315 4295
rect 5485 4210 5515 4295
rect 5685 4210 5715 4295
rect 5885 4210 5915 4295
rect 6085 4210 6115 4295
rect 6285 4210 6315 4295
rect 6485 4210 6515 4295
rect -150 4200 -50 4210
rect -150 4120 -140 4200
rect -60 4120 -50 4200
rect -150 4110 -50 4120
rect 50 4200 150 4210
rect 50 4120 60 4200
rect 140 4120 150 4200
rect 50 4110 150 4120
rect 250 4200 350 4210
rect 250 4120 260 4200
rect 340 4120 350 4200
rect 250 4110 350 4120
rect 450 4200 550 4210
rect 450 4120 460 4200
rect 540 4120 550 4200
rect 450 4110 550 4120
rect 650 4200 750 4210
rect 650 4120 660 4200
rect 740 4120 750 4200
rect 650 4110 750 4120
rect 850 4200 950 4210
rect 850 4120 860 4200
rect 940 4120 950 4200
rect 850 4110 950 4120
rect 1050 4200 1150 4210
rect 1050 4120 1060 4200
rect 1140 4120 1150 4200
rect 1050 4110 1150 4120
rect 1250 4200 1350 4210
rect 1250 4120 1260 4200
rect 1340 4120 1350 4200
rect 1250 4110 1350 4120
rect 1450 4200 1550 4210
rect 1450 4120 1460 4200
rect 1540 4120 1550 4200
rect 1450 4110 1550 4120
rect 1650 4200 1750 4210
rect 1650 4120 1660 4200
rect 1740 4120 1750 4200
rect 1650 4110 1750 4120
rect 1850 4200 1950 4210
rect 1850 4120 1860 4200
rect 1940 4120 1950 4200
rect 1850 4110 1950 4120
rect 2050 4200 2150 4210
rect 2050 4120 2060 4200
rect 2140 4120 2150 4200
rect 2050 4110 2150 4120
rect 2250 4200 2350 4210
rect 2250 4120 2260 4200
rect 2340 4120 2350 4200
rect 2250 4110 2350 4120
rect 2450 4200 2550 4210
rect 2450 4120 2460 4200
rect 2540 4120 2550 4200
rect 2450 4110 2550 4120
rect 2650 4200 2750 4210
rect 2650 4120 2660 4200
rect 2740 4120 2750 4200
rect 2650 4110 2750 4120
rect 2850 4200 2950 4210
rect 2850 4120 2860 4200
rect 2940 4120 2950 4200
rect 2850 4110 2950 4120
rect 3050 4200 3150 4210
rect 3050 4120 3060 4200
rect 3140 4120 3150 4200
rect 3050 4110 3150 4120
rect 3250 4200 3350 4210
rect 3250 4120 3260 4200
rect 3340 4120 3350 4200
rect 3250 4110 3350 4120
rect 3450 4200 3550 4210
rect 3450 4120 3460 4200
rect 3540 4120 3550 4200
rect 3450 4110 3550 4120
rect 3650 4200 3750 4210
rect 3650 4120 3660 4200
rect 3740 4120 3750 4200
rect 3650 4110 3750 4120
rect 3850 4200 3950 4210
rect 3850 4120 3860 4200
rect 3940 4120 3950 4200
rect 3850 4110 3950 4120
rect 4050 4200 4150 4210
rect 4050 4120 4060 4200
rect 4140 4120 4150 4200
rect 4050 4110 4150 4120
rect 4250 4200 4350 4210
rect 4250 4120 4260 4200
rect 4340 4120 4350 4200
rect 4250 4110 4350 4120
rect 4450 4200 4550 4210
rect 4450 4120 4460 4200
rect 4540 4120 4550 4200
rect 4450 4110 4550 4120
rect 4650 4200 4750 4210
rect 4650 4120 4660 4200
rect 4740 4120 4750 4200
rect 4650 4110 4750 4120
rect 4850 4200 4950 4210
rect 4850 4120 4860 4200
rect 4940 4120 4950 4200
rect 4850 4110 4950 4120
rect 5050 4200 5150 4210
rect 5050 4120 5060 4200
rect 5140 4120 5150 4200
rect 5050 4110 5150 4120
rect 5250 4200 5350 4210
rect 5250 4120 5260 4200
rect 5340 4120 5350 4200
rect 5250 4110 5350 4120
rect 5450 4200 5550 4210
rect 5450 4120 5460 4200
rect 5540 4120 5550 4200
rect 5450 4110 5550 4120
rect 5650 4200 5750 4210
rect 5650 4120 5660 4200
rect 5740 4120 5750 4200
rect 5650 4110 5750 4120
rect 5850 4200 5950 4210
rect 5850 4120 5860 4200
rect 5940 4120 5950 4200
rect 5850 4110 5950 4120
rect 6050 4200 6150 4210
rect 6050 4120 6060 4200
rect 6140 4120 6150 4200
rect 6050 4110 6150 4120
rect 6250 4200 6350 4210
rect 6250 4120 6260 4200
rect 6340 4120 6350 4200
rect 6250 4110 6350 4120
rect 6450 4200 6550 4210
rect 6450 4120 6460 4200
rect 6540 4120 6550 4200
rect 6450 4110 6550 4120
rect -115 4025 -85 4110
rect 85 4025 115 4110
rect 285 4025 315 4110
rect 485 4025 515 4110
rect 685 4025 715 4110
rect 885 4025 915 4110
rect 1085 4025 1115 4110
rect 1285 4025 1315 4110
rect 1485 4025 1515 4110
rect 1685 4025 1715 4110
rect 1885 4025 1915 4110
rect 2085 4025 2115 4110
rect 2285 4025 2315 4110
rect 2485 4025 2515 4110
rect 2685 4025 2715 4110
rect 2885 4025 2915 4110
rect 3085 4025 3115 4110
rect 3285 4025 3315 4110
rect 3485 4025 3515 4110
rect 3685 4025 3715 4110
rect 3885 4025 3915 4110
rect 4085 4025 4115 4110
rect 4285 4025 4315 4110
rect 4485 4025 4515 4110
rect 4685 4025 4715 4110
rect 4885 4025 4915 4110
rect 5085 4025 5115 4110
rect 5285 4025 5315 4110
rect 5485 4025 5515 4110
rect 5685 4025 5715 4110
rect 5885 4025 5915 4110
rect 6085 4025 6115 4110
rect 6285 4025 6315 4110
rect 6485 4025 6515 4110
rect -150 4015 -50 4025
rect -150 3935 -140 4015
rect -60 3935 -50 4015
rect -150 3925 -50 3935
rect 50 4015 150 4025
rect 50 3935 60 4015
rect 140 3935 150 4015
rect 50 3925 150 3935
rect 250 4015 350 4025
rect 250 3935 260 4015
rect 340 3935 350 4015
rect 250 3925 350 3935
rect 450 4015 550 4025
rect 450 3935 460 4015
rect 540 3935 550 4015
rect 450 3925 550 3935
rect 650 4015 750 4025
rect 650 3935 660 4015
rect 740 3935 750 4015
rect 650 3925 750 3935
rect 850 4015 950 4025
rect 850 3935 860 4015
rect 940 3935 950 4015
rect 850 3925 950 3935
rect 1050 4015 1150 4025
rect 1050 3935 1060 4015
rect 1140 3935 1150 4015
rect 1050 3925 1150 3935
rect 1250 4015 1350 4025
rect 1250 3935 1260 4015
rect 1340 3935 1350 4015
rect 1250 3925 1350 3935
rect 1450 4015 1550 4025
rect 1450 3935 1460 4015
rect 1540 3935 1550 4015
rect 1450 3925 1550 3935
rect 1650 4015 1750 4025
rect 1650 3935 1660 4015
rect 1740 3935 1750 4015
rect 1650 3925 1750 3935
rect 1850 4015 1950 4025
rect 1850 3935 1860 4015
rect 1940 3935 1950 4015
rect 1850 3925 1950 3935
rect 2050 4015 2150 4025
rect 2050 3935 2060 4015
rect 2140 3935 2150 4015
rect 2050 3925 2150 3935
rect 2250 4015 2350 4025
rect 2250 3935 2260 4015
rect 2340 3935 2350 4015
rect 2250 3925 2350 3935
rect 2450 4015 2550 4025
rect 2450 3935 2460 4015
rect 2540 3935 2550 4015
rect 2450 3925 2550 3935
rect 2650 4015 2750 4025
rect 2650 3935 2660 4015
rect 2740 3935 2750 4015
rect 2650 3925 2750 3935
rect 2850 4015 2950 4025
rect 2850 3935 2860 4015
rect 2940 3935 2950 4015
rect 2850 3925 2950 3935
rect 3050 4015 3150 4025
rect 3050 3935 3060 4015
rect 3140 3935 3150 4015
rect 3050 3925 3150 3935
rect 3250 4015 3350 4025
rect 3250 3935 3260 4015
rect 3340 3935 3350 4015
rect 3250 3925 3350 3935
rect 3450 4015 3550 4025
rect 3450 3935 3460 4015
rect 3540 3935 3550 4015
rect 3450 3925 3550 3935
rect 3650 4015 3750 4025
rect 3650 3935 3660 4015
rect 3740 3935 3750 4015
rect 3650 3925 3750 3935
rect 3850 4015 3950 4025
rect 3850 3935 3860 4015
rect 3940 3935 3950 4015
rect 3850 3925 3950 3935
rect 4050 4015 4150 4025
rect 4050 3935 4060 4015
rect 4140 3935 4150 4015
rect 4050 3925 4150 3935
rect 4250 4015 4350 4025
rect 4250 3935 4260 4015
rect 4340 3935 4350 4015
rect 4250 3925 4350 3935
rect 4450 4015 4550 4025
rect 4450 3935 4460 4015
rect 4540 3935 4550 4015
rect 4450 3925 4550 3935
rect 4650 4015 4750 4025
rect 4650 3935 4660 4015
rect 4740 3935 4750 4015
rect 4650 3925 4750 3935
rect 4850 4015 4950 4025
rect 4850 3935 4860 4015
rect 4940 3935 4950 4015
rect 4850 3925 4950 3935
rect 5050 4015 5150 4025
rect 5050 3935 5060 4015
rect 5140 3935 5150 4015
rect 5050 3925 5150 3935
rect 5250 4015 5350 4025
rect 5250 3935 5260 4015
rect 5340 3935 5350 4015
rect 5250 3925 5350 3935
rect 5450 4015 5550 4025
rect 5450 3935 5460 4015
rect 5540 3935 5550 4015
rect 5450 3925 5550 3935
rect 5650 4015 5750 4025
rect 5650 3935 5660 4015
rect 5740 3935 5750 4015
rect 5650 3925 5750 3935
rect 5850 4015 5950 4025
rect 5850 3935 5860 4015
rect 5940 3935 5950 4015
rect 5850 3925 5950 3935
rect 6050 4015 6150 4025
rect 6050 3935 6060 4015
rect 6140 3935 6150 4015
rect 6050 3925 6150 3935
rect 6250 4015 6350 4025
rect 6250 3935 6260 4015
rect 6340 3935 6350 4015
rect 6250 3925 6350 3935
rect 6450 4015 6550 4025
rect 6450 3935 6460 4015
rect 6540 3935 6550 4015
rect 6450 3925 6550 3935
rect -115 3840 -85 3925
rect 85 3840 115 3925
rect 285 3840 315 3925
rect 485 3840 515 3925
rect 685 3840 715 3925
rect 885 3840 915 3925
rect 1085 3840 1115 3925
rect 1285 3840 1315 3925
rect 1485 3840 1515 3925
rect 1685 3840 1715 3925
rect 1885 3840 1915 3925
rect 2085 3840 2115 3925
rect 2285 3840 2315 3925
rect 2485 3840 2515 3925
rect 2685 3840 2715 3925
rect 2885 3840 2915 3925
rect 3085 3840 3115 3925
rect 3285 3840 3315 3925
rect 3485 3840 3515 3925
rect 3685 3840 3715 3925
rect 3885 3840 3915 3925
rect 4085 3840 4115 3925
rect 4285 3840 4315 3925
rect 4485 3840 4515 3925
rect 4685 3840 4715 3925
rect 4885 3840 4915 3925
rect 5085 3840 5115 3925
rect 5285 3840 5315 3925
rect 5485 3840 5515 3925
rect 5685 3840 5715 3925
rect 5885 3840 5915 3925
rect 6085 3840 6115 3925
rect 6285 3840 6315 3925
rect 6485 3840 6515 3925
rect -150 3830 -50 3840
rect -150 3750 -140 3830
rect -60 3750 -50 3830
rect -150 3740 -50 3750
rect 50 3830 150 3840
rect 50 3750 60 3830
rect 140 3750 150 3830
rect 50 3740 150 3750
rect 250 3830 350 3840
rect 250 3750 260 3830
rect 340 3750 350 3830
rect 250 3740 350 3750
rect 450 3830 550 3840
rect 450 3750 460 3830
rect 540 3750 550 3830
rect 450 3740 550 3750
rect 650 3830 750 3840
rect 650 3750 660 3830
rect 740 3750 750 3830
rect 650 3740 750 3750
rect 850 3830 950 3840
rect 850 3750 860 3830
rect 940 3750 950 3830
rect 850 3740 950 3750
rect 1050 3830 1150 3840
rect 1050 3750 1060 3830
rect 1140 3750 1150 3830
rect 1050 3740 1150 3750
rect 1250 3830 1350 3840
rect 1250 3750 1260 3830
rect 1340 3750 1350 3830
rect 1250 3740 1350 3750
rect 1450 3830 1550 3840
rect 1450 3750 1460 3830
rect 1540 3750 1550 3830
rect 1450 3740 1550 3750
rect 1650 3830 1750 3840
rect 1650 3750 1660 3830
rect 1740 3750 1750 3830
rect 1650 3740 1750 3750
rect 1850 3830 1950 3840
rect 1850 3750 1860 3830
rect 1940 3750 1950 3830
rect 1850 3740 1950 3750
rect 2050 3830 2150 3840
rect 2050 3750 2060 3830
rect 2140 3750 2150 3830
rect 2050 3740 2150 3750
rect 2250 3830 2350 3840
rect 2250 3750 2260 3830
rect 2340 3750 2350 3830
rect 2250 3740 2350 3750
rect 2450 3830 2550 3840
rect 2450 3750 2460 3830
rect 2540 3750 2550 3830
rect 2450 3740 2550 3750
rect 2650 3830 2750 3840
rect 2650 3750 2660 3830
rect 2740 3750 2750 3830
rect 2650 3740 2750 3750
rect 2850 3830 2950 3840
rect 2850 3750 2860 3830
rect 2940 3750 2950 3830
rect 2850 3740 2950 3750
rect 3050 3830 3150 3840
rect 3050 3750 3060 3830
rect 3140 3750 3150 3830
rect 3050 3740 3150 3750
rect 3250 3830 3350 3840
rect 3250 3750 3260 3830
rect 3340 3750 3350 3830
rect 3250 3740 3350 3750
rect 3450 3830 3550 3840
rect 3450 3750 3460 3830
rect 3540 3750 3550 3830
rect 3450 3740 3550 3750
rect 3650 3830 3750 3840
rect 3650 3750 3660 3830
rect 3740 3750 3750 3830
rect 3650 3740 3750 3750
rect 3850 3830 3950 3840
rect 3850 3750 3860 3830
rect 3940 3750 3950 3830
rect 3850 3740 3950 3750
rect 4050 3830 4150 3840
rect 4050 3750 4060 3830
rect 4140 3750 4150 3830
rect 4050 3740 4150 3750
rect 4250 3830 4350 3840
rect 4250 3750 4260 3830
rect 4340 3750 4350 3830
rect 4250 3740 4350 3750
rect 4450 3830 4550 3840
rect 4450 3750 4460 3830
rect 4540 3750 4550 3830
rect 4450 3740 4550 3750
rect 4650 3830 4750 3840
rect 4650 3750 4660 3830
rect 4740 3750 4750 3830
rect 4650 3740 4750 3750
rect 4850 3830 4950 3840
rect 4850 3750 4860 3830
rect 4940 3750 4950 3830
rect 4850 3740 4950 3750
rect 5050 3830 5150 3840
rect 5050 3750 5060 3830
rect 5140 3750 5150 3830
rect 5050 3740 5150 3750
rect 5250 3830 5350 3840
rect 5250 3750 5260 3830
rect 5340 3750 5350 3830
rect 5250 3740 5350 3750
rect 5450 3830 5550 3840
rect 5450 3750 5460 3830
rect 5540 3750 5550 3830
rect 5450 3740 5550 3750
rect 5650 3830 5750 3840
rect 5650 3750 5660 3830
rect 5740 3750 5750 3830
rect 5650 3740 5750 3750
rect 5850 3830 5950 3840
rect 5850 3750 5860 3830
rect 5940 3750 5950 3830
rect 5850 3740 5950 3750
rect 6050 3830 6150 3840
rect 6050 3750 6060 3830
rect 6140 3750 6150 3830
rect 6050 3740 6150 3750
rect 6250 3830 6350 3840
rect 6250 3750 6260 3830
rect 6340 3750 6350 3830
rect 6250 3740 6350 3750
rect 6450 3830 6550 3840
rect 6450 3750 6460 3830
rect 6540 3750 6550 3830
rect 6450 3740 6550 3750
rect -115 3655 -85 3740
rect 85 3655 115 3740
rect 285 3655 315 3740
rect 485 3655 515 3740
rect 685 3655 715 3740
rect 885 3655 915 3740
rect 1085 3655 1115 3740
rect 1285 3655 1315 3740
rect 1485 3655 1515 3740
rect 1685 3655 1715 3740
rect 1885 3655 1915 3740
rect 2085 3655 2115 3740
rect 2285 3655 2315 3740
rect 2485 3655 2515 3740
rect 2685 3655 2715 3740
rect 2885 3655 2915 3740
rect 3085 3655 3115 3740
rect 3285 3655 3315 3740
rect 3485 3655 3515 3740
rect 3685 3655 3715 3740
rect 3885 3655 3915 3740
rect 4085 3655 4115 3740
rect 4285 3655 4315 3740
rect 4485 3655 4515 3740
rect 4685 3655 4715 3740
rect 4885 3655 4915 3740
rect 5085 3655 5115 3740
rect 5285 3655 5315 3740
rect 5485 3655 5515 3740
rect 5685 3655 5715 3740
rect 5885 3655 5915 3740
rect 6085 3655 6115 3740
rect 6285 3655 6315 3740
rect 6485 3655 6515 3740
rect -150 3645 -50 3655
rect -150 3565 -140 3645
rect -60 3565 -50 3645
rect -150 3555 -50 3565
rect 50 3645 150 3655
rect 50 3565 60 3645
rect 140 3565 150 3645
rect 50 3555 150 3565
rect 250 3645 350 3655
rect 250 3565 260 3645
rect 340 3565 350 3645
rect 250 3555 350 3565
rect 450 3645 550 3655
rect 450 3565 460 3645
rect 540 3565 550 3645
rect 450 3555 550 3565
rect 650 3645 750 3655
rect 650 3565 660 3645
rect 740 3565 750 3645
rect 650 3555 750 3565
rect 850 3645 950 3655
rect 850 3565 860 3645
rect 940 3565 950 3645
rect 850 3555 950 3565
rect 1050 3645 1150 3655
rect 1050 3565 1060 3645
rect 1140 3565 1150 3645
rect 1050 3555 1150 3565
rect 1250 3645 1350 3655
rect 1250 3565 1260 3645
rect 1340 3565 1350 3645
rect 1250 3555 1350 3565
rect 1450 3645 1550 3655
rect 1450 3565 1460 3645
rect 1540 3565 1550 3645
rect 1450 3555 1550 3565
rect 1650 3645 1750 3655
rect 1650 3565 1660 3645
rect 1740 3565 1750 3645
rect 1650 3555 1750 3565
rect 1850 3645 1950 3655
rect 1850 3565 1860 3645
rect 1940 3565 1950 3645
rect 1850 3555 1950 3565
rect 2050 3645 2150 3655
rect 2050 3565 2060 3645
rect 2140 3565 2150 3645
rect 2050 3555 2150 3565
rect 2250 3645 2350 3655
rect 2250 3565 2260 3645
rect 2340 3565 2350 3645
rect 2250 3555 2350 3565
rect 2450 3645 2550 3655
rect 2450 3565 2460 3645
rect 2540 3565 2550 3645
rect 2450 3555 2550 3565
rect 2650 3645 2750 3655
rect 2650 3565 2660 3645
rect 2740 3565 2750 3645
rect 2650 3555 2750 3565
rect 2850 3645 2950 3655
rect 2850 3565 2860 3645
rect 2940 3565 2950 3645
rect 2850 3555 2950 3565
rect 3050 3645 3150 3655
rect 3050 3565 3060 3645
rect 3140 3565 3150 3645
rect 3050 3555 3150 3565
rect 3250 3645 3350 3655
rect 3250 3565 3260 3645
rect 3340 3565 3350 3645
rect 3250 3555 3350 3565
rect 3450 3645 3550 3655
rect 3450 3565 3460 3645
rect 3540 3565 3550 3645
rect 3450 3555 3550 3565
rect 3650 3645 3750 3655
rect 3650 3565 3660 3645
rect 3740 3565 3750 3645
rect 3650 3555 3750 3565
rect 3850 3645 3950 3655
rect 3850 3565 3860 3645
rect 3940 3565 3950 3645
rect 3850 3555 3950 3565
rect 4050 3645 4150 3655
rect 4050 3565 4060 3645
rect 4140 3565 4150 3645
rect 4050 3555 4150 3565
rect 4250 3645 4350 3655
rect 4250 3565 4260 3645
rect 4340 3565 4350 3645
rect 4250 3555 4350 3565
rect 4450 3645 4550 3655
rect 4450 3565 4460 3645
rect 4540 3565 4550 3645
rect 4450 3555 4550 3565
rect 4650 3645 4750 3655
rect 4650 3565 4660 3645
rect 4740 3565 4750 3645
rect 4650 3555 4750 3565
rect 4850 3645 4950 3655
rect 4850 3565 4860 3645
rect 4940 3565 4950 3645
rect 4850 3555 4950 3565
rect 5050 3645 5150 3655
rect 5050 3565 5060 3645
rect 5140 3565 5150 3645
rect 5050 3555 5150 3565
rect 5250 3645 5350 3655
rect 5250 3565 5260 3645
rect 5340 3565 5350 3645
rect 5250 3555 5350 3565
rect 5450 3645 5550 3655
rect 5450 3565 5460 3645
rect 5540 3565 5550 3645
rect 5450 3555 5550 3565
rect 5650 3645 5750 3655
rect 5650 3565 5660 3645
rect 5740 3565 5750 3645
rect 5650 3555 5750 3565
rect 5850 3645 5950 3655
rect 5850 3565 5860 3645
rect 5940 3565 5950 3645
rect 5850 3555 5950 3565
rect 6050 3645 6150 3655
rect 6050 3565 6060 3645
rect 6140 3565 6150 3645
rect 6050 3555 6150 3565
rect 6250 3645 6350 3655
rect 6250 3565 6260 3645
rect 6340 3565 6350 3645
rect 6250 3555 6350 3565
rect 6450 3645 6550 3655
rect 6450 3565 6460 3645
rect 6540 3565 6550 3645
rect 6450 3555 6550 3565
rect -115 3470 -85 3555
rect 85 3470 115 3555
rect 285 3470 315 3555
rect 485 3470 515 3555
rect 685 3470 715 3555
rect 885 3470 915 3555
rect 1085 3470 1115 3555
rect 1285 3470 1315 3555
rect 1485 3470 1515 3555
rect 1685 3470 1715 3555
rect 1885 3470 1915 3555
rect 2085 3470 2115 3555
rect 2285 3470 2315 3555
rect 2485 3470 2515 3555
rect 2685 3470 2715 3555
rect 2885 3470 2915 3555
rect 3085 3470 3115 3555
rect 3285 3470 3315 3555
rect 3485 3470 3515 3555
rect 3685 3470 3715 3555
rect 3885 3470 3915 3555
rect 4085 3470 4115 3555
rect 4285 3470 4315 3555
rect 4485 3470 4515 3555
rect 4685 3470 4715 3555
rect 4885 3470 4915 3555
rect 5085 3470 5115 3555
rect 5285 3470 5315 3555
rect 5485 3470 5515 3555
rect 5685 3470 5715 3555
rect 5885 3470 5915 3555
rect 6085 3470 6115 3555
rect 6285 3470 6315 3555
rect 6485 3470 6515 3555
rect -150 3460 -50 3470
rect -150 3380 -140 3460
rect -60 3380 -50 3460
rect -150 3370 -50 3380
rect 50 3460 150 3470
rect 50 3380 60 3460
rect 140 3380 150 3460
rect 50 3370 150 3380
rect 250 3460 350 3470
rect 250 3380 260 3460
rect 340 3380 350 3460
rect 250 3370 350 3380
rect 450 3460 550 3470
rect 450 3380 460 3460
rect 540 3380 550 3460
rect 450 3370 550 3380
rect 650 3460 750 3470
rect 650 3380 660 3460
rect 740 3380 750 3460
rect 650 3370 750 3380
rect 850 3460 950 3470
rect 850 3380 860 3460
rect 940 3380 950 3460
rect 850 3370 950 3380
rect 1050 3460 1150 3470
rect 1050 3380 1060 3460
rect 1140 3380 1150 3460
rect 1050 3370 1150 3380
rect 1250 3460 1350 3470
rect 1250 3380 1260 3460
rect 1340 3380 1350 3460
rect 1250 3370 1350 3380
rect 1450 3460 1550 3470
rect 1450 3380 1460 3460
rect 1540 3380 1550 3460
rect 1450 3370 1550 3380
rect 1650 3460 1750 3470
rect 1650 3380 1660 3460
rect 1740 3380 1750 3460
rect 1650 3370 1750 3380
rect 1850 3460 1950 3470
rect 1850 3380 1860 3460
rect 1940 3380 1950 3460
rect 1850 3370 1950 3380
rect 2050 3460 2150 3470
rect 2050 3380 2060 3460
rect 2140 3380 2150 3460
rect 2050 3370 2150 3380
rect 2250 3460 2350 3470
rect 2250 3380 2260 3460
rect 2340 3380 2350 3460
rect 2250 3370 2350 3380
rect 2450 3460 2550 3470
rect 2450 3380 2460 3460
rect 2540 3380 2550 3460
rect 2450 3370 2550 3380
rect 2650 3460 2750 3470
rect 2650 3380 2660 3460
rect 2740 3380 2750 3460
rect 2650 3370 2750 3380
rect 2850 3460 2950 3470
rect 2850 3380 2860 3460
rect 2940 3380 2950 3460
rect 2850 3370 2950 3380
rect 3050 3460 3150 3470
rect 3050 3380 3060 3460
rect 3140 3380 3150 3460
rect 3050 3370 3150 3380
rect 3250 3460 3350 3470
rect 3250 3380 3260 3460
rect 3340 3380 3350 3460
rect 3250 3370 3350 3380
rect 3450 3460 3550 3470
rect 3450 3380 3460 3460
rect 3540 3380 3550 3460
rect 3450 3370 3550 3380
rect 3650 3460 3750 3470
rect 3650 3380 3660 3460
rect 3740 3380 3750 3460
rect 3650 3370 3750 3380
rect 3850 3460 3950 3470
rect 3850 3380 3860 3460
rect 3940 3380 3950 3460
rect 3850 3370 3950 3380
rect 4050 3460 4150 3470
rect 4050 3380 4060 3460
rect 4140 3380 4150 3460
rect 4050 3370 4150 3380
rect 4250 3460 4350 3470
rect 4250 3380 4260 3460
rect 4340 3380 4350 3460
rect 4250 3370 4350 3380
rect 4450 3460 4550 3470
rect 4450 3380 4460 3460
rect 4540 3380 4550 3460
rect 4450 3370 4550 3380
rect 4650 3460 4750 3470
rect 4650 3380 4660 3460
rect 4740 3380 4750 3460
rect 4650 3370 4750 3380
rect 4850 3460 4950 3470
rect 4850 3380 4860 3460
rect 4940 3380 4950 3460
rect 4850 3370 4950 3380
rect 5050 3460 5150 3470
rect 5050 3380 5060 3460
rect 5140 3380 5150 3460
rect 5050 3370 5150 3380
rect 5250 3460 5350 3470
rect 5250 3380 5260 3460
rect 5340 3380 5350 3460
rect 5250 3370 5350 3380
rect 5450 3460 5550 3470
rect 5450 3380 5460 3460
rect 5540 3380 5550 3460
rect 5450 3370 5550 3380
rect 5650 3460 5750 3470
rect 5650 3380 5660 3460
rect 5740 3380 5750 3460
rect 5650 3370 5750 3380
rect 5850 3460 5950 3470
rect 5850 3380 5860 3460
rect 5940 3380 5950 3460
rect 5850 3370 5950 3380
rect 6050 3460 6150 3470
rect 6050 3380 6060 3460
rect 6140 3380 6150 3460
rect 6050 3370 6150 3380
rect 6250 3460 6350 3470
rect 6250 3380 6260 3460
rect 6340 3380 6350 3460
rect 6250 3370 6350 3380
rect 6450 3460 6550 3470
rect 6450 3380 6460 3460
rect 6540 3380 6550 3460
rect 6450 3370 6550 3380
rect -115 3285 -85 3370
rect 85 3285 115 3370
rect 285 3285 315 3370
rect 485 3285 515 3370
rect 685 3285 715 3370
rect 885 3285 915 3370
rect 1085 3285 1115 3370
rect 1285 3285 1315 3370
rect 1485 3285 1515 3370
rect 1685 3285 1715 3370
rect 1885 3285 1915 3370
rect 2085 3285 2115 3370
rect 2285 3285 2315 3370
rect 2485 3285 2515 3370
rect 2685 3285 2715 3370
rect 2885 3285 2915 3370
rect 3085 3285 3115 3370
rect 3285 3285 3315 3370
rect 3485 3285 3515 3370
rect 3685 3285 3715 3370
rect 3885 3285 3915 3370
rect 4085 3285 4115 3370
rect 4285 3285 4315 3370
rect 4485 3285 4515 3370
rect 4685 3285 4715 3370
rect 4885 3285 4915 3370
rect 5085 3285 5115 3370
rect 5285 3285 5315 3370
rect 5485 3285 5515 3370
rect 5685 3285 5715 3370
rect 5885 3285 5915 3370
rect 6085 3285 6115 3370
rect 6285 3285 6315 3370
rect 6485 3285 6515 3370
rect -150 3275 -50 3285
rect -150 3195 -140 3275
rect -60 3195 -50 3275
rect -150 3185 -50 3195
rect 50 3275 150 3285
rect 50 3195 60 3275
rect 140 3195 150 3275
rect 50 3185 150 3195
rect 250 3275 350 3285
rect 250 3195 260 3275
rect 340 3195 350 3275
rect 250 3185 350 3195
rect 450 3275 550 3285
rect 450 3195 460 3275
rect 540 3195 550 3275
rect 450 3185 550 3195
rect 650 3275 750 3285
rect 650 3195 660 3275
rect 740 3195 750 3275
rect 650 3185 750 3195
rect 850 3275 950 3285
rect 850 3195 860 3275
rect 940 3195 950 3275
rect 850 3185 950 3195
rect 1050 3275 1150 3285
rect 1050 3195 1060 3275
rect 1140 3195 1150 3275
rect 1050 3185 1150 3195
rect 1250 3275 1350 3285
rect 1250 3195 1260 3275
rect 1340 3195 1350 3275
rect 1250 3185 1350 3195
rect 1450 3275 1550 3285
rect 1450 3195 1460 3275
rect 1540 3195 1550 3275
rect 1450 3185 1550 3195
rect 1650 3275 1750 3285
rect 1650 3195 1660 3275
rect 1740 3195 1750 3275
rect 1650 3185 1750 3195
rect 1850 3275 1950 3285
rect 1850 3195 1860 3275
rect 1940 3195 1950 3275
rect 1850 3185 1950 3195
rect 2050 3275 2150 3285
rect 2050 3195 2060 3275
rect 2140 3195 2150 3275
rect 2050 3185 2150 3195
rect 2250 3275 2350 3285
rect 2250 3195 2260 3275
rect 2340 3195 2350 3275
rect 2250 3185 2350 3195
rect 2450 3275 2550 3285
rect 2450 3195 2460 3275
rect 2540 3195 2550 3275
rect 2450 3185 2550 3195
rect 2650 3275 2750 3285
rect 2650 3195 2660 3275
rect 2740 3195 2750 3275
rect 2650 3185 2750 3195
rect 2850 3275 2950 3285
rect 2850 3195 2860 3275
rect 2940 3195 2950 3275
rect 2850 3185 2950 3195
rect 3050 3275 3150 3285
rect 3050 3195 3060 3275
rect 3140 3195 3150 3275
rect 3050 3185 3150 3195
rect 3250 3275 3350 3285
rect 3250 3195 3260 3275
rect 3340 3195 3350 3275
rect 3250 3185 3350 3195
rect 3450 3275 3550 3285
rect 3450 3195 3460 3275
rect 3540 3195 3550 3275
rect 3450 3185 3550 3195
rect 3650 3275 3750 3285
rect 3650 3195 3660 3275
rect 3740 3195 3750 3275
rect 3650 3185 3750 3195
rect 3850 3275 3950 3285
rect 3850 3195 3860 3275
rect 3940 3195 3950 3275
rect 3850 3185 3950 3195
rect 4050 3275 4150 3285
rect 4050 3195 4060 3275
rect 4140 3195 4150 3275
rect 4050 3185 4150 3195
rect 4250 3275 4350 3285
rect 4250 3195 4260 3275
rect 4340 3195 4350 3275
rect 4250 3185 4350 3195
rect 4450 3275 4550 3285
rect 4450 3195 4460 3275
rect 4540 3195 4550 3275
rect 4450 3185 4550 3195
rect 4650 3275 4750 3285
rect 4650 3195 4660 3275
rect 4740 3195 4750 3275
rect 4650 3185 4750 3195
rect 4850 3275 4950 3285
rect 4850 3195 4860 3275
rect 4940 3195 4950 3275
rect 4850 3185 4950 3195
rect 5050 3275 5150 3285
rect 5050 3195 5060 3275
rect 5140 3195 5150 3275
rect 5050 3185 5150 3195
rect 5250 3275 5350 3285
rect 5250 3195 5260 3275
rect 5340 3195 5350 3275
rect 5250 3185 5350 3195
rect 5450 3275 5550 3285
rect 5450 3195 5460 3275
rect 5540 3195 5550 3275
rect 5450 3185 5550 3195
rect 5650 3275 5750 3285
rect 5650 3195 5660 3275
rect 5740 3195 5750 3275
rect 5650 3185 5750 3195
rect 5850 3275 5950 3285
rect 5850 3195 5860 3275
rect 5940 3195 5950 3275
rect 5850 3185 5950 3195
rect 6050 3275 6150 3285
rect 6050 3195 6060 3275
rect 6140 3195 6150 3275
rect 6050 3185 6150 3195
rect 6250 3275 6350 3285
rect 6250 3195 6260 3275
rect 6340 3195 6350 3275
rect 6250 3185 6350 3195
rect 6450 3275 6550 3285
rect 6450 3195 6460 3275
rect 6540 3195 6550 3275
rect 6450 3185 6550 3195
rect -115 3100 -85 3185
rect 85 3100 115 3185
rect 285 3100 315 3185
rect 485 3100 515 3185
rect 685 3100 715 3185
rect 885 3100 915 3185
rect 1085 3100 1115 3185
rect 1285 3100 1315 3185
rect 1485 3100 1515 3185
rect 1685 3100 1715 3185
rect 1885 3100 1915 3185
rect 2085 3100 2115 3185
rect 2285 3100 2315 3185
rect 2485 3100 2515 3185
rect 2685 3100 2715 3185
rect 2885 3100 2915 3185
rect 3085 3100 3115 3185
rect 3285 3100 3315 3185
rect 3485 3100 3515 3185
rect 3685 3100 3715 3185
rect 3885 3100 3915 3185
rect 4085 3100 4115 3185
rect 4285 3100 4315 3185
rect 4485 3100 4515 3185
rect 4685 3100 4715 3185
rect 4885 3100 4915 3185
rect 5085 3100 5115 3185
rect 5285 3100 5315 3185
rect 5485 3100 5515 3185
rect 5685 3100 5715 3185
rect 5885 3100 5915 3185
rect 6085 3100 6115 3185
rect 6285 3100 6315 3185
rect 6485 3100 6515 3185
rect -150 3090 -50 3100
rect -150 3010 -140 3090
rect -60 3010 -50 3090
rect -150 3000 -50 3010
rect 50 3090 150 3100
rect 50 3010 60 3090
rect 140 3010 150 3090
rect 50 3000 150 3010
rect 250 3090 350 3100
rect 250 3010 260 3090
rect 340 3010 350 3090
rect 250 3000 350 3010
rect 450 3090 550 3100
rect 450 3010 460 3090
rect 540 3010 550 3090
rect 450 3000 550 3010
rect 650 3090 750 3100
rect 650 3010 660 3090
rect 740 3010 750 3090
rect 650 3000 750 3010
rect 850 3090 950 3100
rect 850 3010 860 3090
rect 940 3010 950 3090
rect 850 3000 950 3010
rect 1050 3090 1150 3100
rect 1050 3010 1060 3090
rect 1140 3010 1150 3090
rect 1050 3000 1150 3010
rect 1250 3090 1350 3100
rect 1250 3010 1260 3090
rect 1340 3010 1350 3090
rect 1250 3000 1350 3010
rect 1450 3090 1550 3100
rect 1450 3010 1460 3090
rect 1540 3010 1550 3090
rect 1450 3000 1550 3010
rect 1650 3090 1750 3100
rect 1650 3010 1660 3090
rect 1740 3010 1750 3090
rect 1650 3000 1750 3010
rect 1850 3090 1950 3100
rect 1850 3010 1860 3090
rect 1940 3010 1950 3090
rect 1850 3000 1950 3010
rect 2050 3090 2150 3100
rect 2050 3010 2060 3090
rect 2140 3010 2150 3090
rect 2050 3000 2150 3010
rect 2250 3090 2350 3100
rect 2250 3010 2260 3090
rect 2340 3010 2350 3090
rect 2250 3000 2350 3010
rect 2450 3090 2550 3100
rect 2450 3010 2460 3090
rect 2540 3010 2550 3090
rect 2450 3000 2550 3010
rect 2650 3090 2750 3100
rect 2650 3010 2660 3090
rect 2740 3010 2750 3090
rect 2650 3000 2750 3010
rect 2850 3090 2950 3100
rect 2850 3010 2860 3090
rect 2940 3010 2950 3090
rect 2850 3000 2950 3010
rect 3050 3090 3150 3100
rect 3050 3010 3060 3090
rect 3140 3010 3150 3090
rect 3050 3000 3150 3010
rect 3250 3090 3350 3100
rect 3250 3010 3260 3090
rect 3340 3010 3350 3090
rect 3250 3000 3350 3010
rect 3450 3090 3550 3100
rect 3450 3010 3460 3090
rect 3540 3010 3550 3090
rect 3450 3000 3550 3010
rect 3650 3090 3750 3100
rect 3650 3010 3660 3090
rect 3740 3010 3750 3090
rect 3650 3000 3750 3010
rect 3850 3090 3950 3100
rect 3850 3010 3860 3090
rect 3940 3010 3950 3090
rect 3850 3000 3950 3010
rect 4050 3090 4150 3100
rect 4050 3010 4060 3090
rect 4140 3010 4150 3090
rect 4050 3000 4150 3010
rect 4250 3090 4350 3100
rect 4250 3010 4260 3090
rect 4340 3010 4350 3090
rect 4250 3000 4350 3010
rect 4450 3090 4550 3100
rect 4450 3010 4460 3090
rect 4540 3010 4550 3090
rect 4450 3000 4550 3010
rect 4650 3090 4750 3100
rect 4650 3010 4660 3090
rect 4740 3010 4750 3090
rect 4650 3000 4750 3010
rect 4850 3090 4950 3100
rect 4850 3010 4860 3090
rect 4940 3010 4950 3090
rect 4850 3000 4950 3010
rect 5050 3090 5150 3100
rect 5050 3010 5060 3090
rect 5140 3010 5150 3090
rect 5050 3000 5150 3010
rect 5250 3090 5350 3100
rect 5250 3010 5260 3090
rect 5340 3010 5350 3090
rect 5250 3000 5350 3010
rect 5450 3090 5550 3100
rect 5450 3010 5460 3090
rect 5540 3010 5550 3090
rect 5450 3000 5550 3010
rect 5650 3090 5750 3100
rect 5650 3010 5660 3090
rect 5740 3010 5750 3090
rect 5650 3000 5750 3010
rect 5850 3090 5950 3100
rect 5850 3010 5860 3090
rect 5940 3010 5950 3090
rect 5850 3000 5950 3010
rect 6050 3090 6150 3100
rect 6050 3010 6060 3090
rect 6140 3010 6150 3090
rect 6050 3000 6150 3010
rect 6250 3090 6350 3100
rect 6250 3010 6260 3090
rect 6340 3010 6350 3090
rect 6250 3000 6350 3010
rect 6450 3090 6550 3100
rect 6450 3010 6460 3090
rect 6540 3010 6550 3090
rect 6450 3000 6550 3010
rect -115 2915 -85 3000
rect 85 2915 115 3000
rect 285 2915 315 3000
rect 485 2915 515 3000
rect 685 2915 715 3000
rect 885 2915 915 3000
rect 1085 2915 1115 3000
rect 1285 2915 1315 3000
rect 1485 2915 1515 3000
rect 1685 2915 1715 3000
rect 1885 2915 1915 3000
rect 2085 2915 2115 3000
rect 2285 2915 2315 3000
rect 2485 2915 2515 3000
rect 2685 2915 2715 3000
rect 2885 2915 2915 3000
rect 3085 2915 3115 3000
rect 3285 2915 3315 3000
rect 3485 2915 3515 3000
rect 3685 2915 3715 3000
rect 3885 2915 3915 3000
rect 4085 2915 4115 3000
rect 4285 2915 4315 3000
rect 4485 2915 4515 3000
rect 4685 2915 4715 3000
rect 4885 2915 4915 3000
rect 5085 2915 5115 3000
rect 5285 2915 5315 3000
rect 5485 2915 5515 3000
rect 5685 2915 5715 3000
rect 5885 2915 5915 3000
rect 6085 2915 6115 3000
rect 6285 2915 6315 3000
rect 6485 2915 6515 3000
rect -150 2905 -50 2915
rect -150 2825 -140 2905
rect -60 2825 -50 2905
rect -150 2815 -50 2825
rect 50 2905 150 2915
rect 50 2825 60 2905
rect 140 2825 150 2905
rect 50 2815 150 2825
rect 250 2905 350 2915
rect 250 2825 260 2905
rect 340 2825 350 2905
rect 250 2815 350 2825
rect 450 2905 550 2915
rect 450 2825 460 2905
rect 540 2825 550 2905
rect 450 2815 550 2825
rect 650 2905 750 2915
rect 650 2825 660 2905
rect 740 2825 750 2905
rect 650 2815 750 2825
rect 850 2905 950 2915
rect 850 2825 860 2905
rect 940 2825 950 2905
rect 850 2815 950 2825
rect 1050 2905 1150 2915
rect 1050 2825 1060 2905
rect 1140 2825 1150 2905
rect 1050 2815 1150 2825
rect 1250 2905 1350 2915
rect 1250 2825 1260 2905
rect 1340 2825 1350 2905
rect 1250 2815 1350 2825
rect 1450 2905 1550 2915
rect 1450 2825 1460 2905
rect 1540 2825 1550 2905
rect 1450 2815 1550 2825
rect 1650 2905 1750 2915
rect 1650 2825 1660 2905
rect 1740 2825 1750 2905
rect 1650 2815 1750 2825
rect 1850 2905 1950 2915
rect 1850 2825 1860 2905
rect 1940 2825 1950 2905
rect 1850 2815 1950 2825
rect 2050 2905 2150 2915
rect 2050 2825 2060 2905
rect 2140 2825 2150 2905
rect 2050 2815 2150 2825
rect 2250 2905 2350 2915
rect 2250 2825 2260 2905
rect 2340 2825 2350 2905
rect 2250 2815 2350 2825
rect 2450 2905 2550 2915
rect 2450 2825 2460 2905
rect 2540 2825 2550 2905
rect 2450 2815 2550 2825
rect 2650 2905 2750 2915
rect 2650 2825 2660 2905
rect 2740 2825 2750 2905
rect 2650 2815 2750 2825
rect 2850 2905 2950 2915
rect 2850 2825 2860 2905
rect 2940 2825 2950 2905
rect 2850 2815 2950 2825
rect 3050 2905 3150 2915
rect 3050 2825 3060 2905
rect 3140 2825 3150 2905
rect 3050 2815 3150 2825
rect 3250 2905 3350 2915
rect 3250 2825 3260 2905
rect 3340 2825 3350 2905
rect 3250 2815 3350 2825
rect 3450 2905 3550 2915
rect 3450 2825 3460 2905
rect 3540 2825 3550 2905
rect 3450 2815 3550 2825
rect 3650 2905 3750 2915
rect 3650 2825 3660 2905
rect 3740 2825 3750 2905
rect 3650 2815 3750 2825
rect 3850 2905 3950 2915
rect 3850 2825 3860 2905
rect 3940 2825 3950 2905
rect 3850 2815 3950 2825
rect 4050 2905 4150 2915
rect 4050 2825 4060 2905
rect 4140 2825 4150 2905
rect 4050 2815 4150 2825
rect 4250 2905 4350 2915
rect 4250 2825 4260 2905
rect 4340 2825 4350 2905
rect 4250 2815 4350 2825
rect 4450 2905 4550 2915
rect 4450 2825 4460 2905
rect 4540 2825 4550 2905
rect 4450 2815 4550 2825
rect 4650 2905 4750 2915
rect 4650 2825 4660 2905
rect 4740 2825 4750 2905
rect 4650 2815 4750 2825
rect 4850 2905 4950 2915
rect 4850 2825 4860 2905
rect 4940 2825 4950 2905
rect 4850 2815 4950 2825
rect 5050 2905 5150 2915
rect 5050 2825 5060 2905
rect 5140 2825 5150 2905
rect 5050 2815 5150 2825
rect 5250 2905 5350 2915
rect 5250 2825 5260 2905
rect 5340 2825 5350 2905
rect 5250 2815 5350 2825
rect 5450 2905 5550 2915
rect 5450 2825 5460 2905
rect 5540 2825 5550 2905
rect 5450 2815 5550 2825
rect 5650 2905 5750 2915
rect 5650 2825 5660 2905
rect 5740 2825 5750 2905
rect 5650 2815 5750 2825
rect 5850 2905 5950 2915
rect 5850 2825 5860 2905
rect 5940 2825 5950 2905
rect 5850 2815 5950 2825
rect 6050 2905 6150 2915
rect 6050 2825 6060 2905
rect 6140 2825 6150 2905
rect 6050 2815 6150 2825
rect 6250 2905 6350 2915
rect 6250 2825 6260 2905
rect 6340 2825 6350 2905
rect 6250 2815 6350 2825
rect 6450 2905 6550 2915
rect 6450 2825 6460 2905
rect 6540 2825 6550 2905
rect 6450 2815 6550 2825
rect -115 2730 -85 2815
rect 85 2730 115 2815
rect 285 2730 315 2815
rect 485 2730 515 2815
rect 685 2730 715 2815
rect 885 2730 915 2815
rect 1085 2730 1115 2815
rect 1285 2730 1315 2815
rect 1485 2730 1515 2815
rect 1685 2730 1715 2815
rect 1885 2730 1915 2815
rect 2085 2730 2115 2815
rect 2285 2730 2315 2815
rect 2485 2730 2515 2815
rect 2685 2730 2715 2815
rect 2885 2730 2915 2815
rect 3085 2730 3115 2815
rect 3285 2730 3315 2815
rect 3485 2730 3515 2815
rect 3685 2730 3715 2815
rect 3885 2730 3915 2815
rect 4085 2730 4115 2815
rect 4285 2730 4315 2815
rect 4485 2730 4515 2815
rect 4685 2730 4715 2815
rect 4885 2730 4915 2815
rect 5085 2730 5115 2815
rect 5285 2730 5315 2815
rect 5485 2730 5515 2815
rect 5685 2730 5715 2815
rect 5885 2730 5915 2815
rect 6085 2730 6115 2815
rect 6285 2730 6315 2815
rect 6485 2730 6515 2815
rect -150 2720 -50 2730
rect -150 2640 -140 2720
rect -60 2640 -50 2720
rect -150 2630 -50 2640
rect 50 2720 150 2730
rect 50 2640 60 2720
rect 140 2640 150 2720
rect 50 2630 150 2640
rect 250 2720 350 2730
rect 250 2640 260 2720
rect 340 2640 350 2720
rect 250 2630 350 2640
rect 450 2720 550 2730
rect 450 2640 460 2720
rect 540 2640 550 2720
rect 450 2630 550 2640
rect 650 2720 750 2730
rect 650 2640 660 2720
rect 740 2640 750 2720
rect 650 2630 750 2640
rect 850 2720 950 2730
rect 850 2640 860 2720
rect 940 2640 950 2720
rect 850 2630 950 2640
rect 1050 2720 1150 2730
rect 1050 2640 1060 2720
rect 1140 2640 1150 2720
rect 1050 2630 1150 2640
rect 1250 2720 1350 2730
rect 1250 2640 1260 2720
rect 1340 2640 1350 2720
rect 1250 2630 1350 2640
rect 1450 2720 1550 2730
rect 1450 2640 1460 2720
rect 1540 2640 1550 2720
rect 1450 2630 1550 2640
rect 1650 2720 1750 2730
rect 1650 2640 1660 2720
rect 1740 2640 1750 2720
rect 1650 2630 1750 2640
rect 1850 2720 1950 2730
rect 1850 2640 1860 2720
rect 1940 2640 1950 2720
rect 1850 2630 1950 2640
rect 2050 2720 2150 2730
rect 2050 2640 2060 2720
rect 2140 2640 2150 2720
rect 2050 2630 2150 2640
rect 2250 2720 2350 2730
rect 2250 2640 2260 2720
rect 2340 2640 2350 2720
rect 2250 2630 2350 2640
rect 2450 2720 2550 2730
rect 2450 2640 2460 2720
rect 2540 2640 2550 2720
rect 2450 2630 2550 2640
rect 2650 2720 2750 2730
rect 2650 2640 2660 2720
rect 2740 2640 2750 2720
rect 2650 2630 2750 2640
rect 2850 2720 2950 2730
rect 2850 2640 2860 2720
rect 2940 2640 2950 2720
rect 2850 2630 2950 2640
rect 3050 2720 3150 2730
rect 3050 2640 3060 2720
rect 3140 2640 3150 2720
rect 3050 2630 3150 2640
rect 3250 2720 3350 2730
rect 3250 2640 3260 2720
rect 3340 2640 3350 2720
rect 3250 2630 3350 2640
rect 3450 2720 3550 2730
rect 3450 2640 3460 2720
rect 3540 2640 3550 2720
rect 3450 2630 3550 2640
rect 3650 2720 3750 2730
rect 3650 2640 3660 2720
rect 3740 2640 3750 2720
rect 3650 2630 3750 2640
rect 3850 2720 3950 2730
rect 3850 2640 3860 2720
rect 3940 2640 3950 2720
rect 3850 2630 3950 2640
rect 4050 2720 4150 2730
rect 4050 2640 4060 2720
rect 4140 2640 4150 2720
rect 4050 2630 4150 2640
rect 4250 2720 4350 2730
rect 4250 2640 4260 2720
rect 4340 2640 4350 2720
rect 4250 2630 4350 2640
rect 4450 2720 4550 2730
rect 4450 2640 4460 2720
rect 4540 2640 4550 2720
rect 4450 2630 4550 2640
rect 4650 2720 4750 2730
rect 4650 2640 4660 2720
rect 4740 2640 4750 2720
rect 4650 2630 4750 2640
rect 4850 2720 4950 2730
rect 4850 2640 4860 2720
rect 4940 2640 4950 2720
rect 4850 2630 4950 2640
rect 5050 2720 5150 2730
rect 5050 2640 5060 2720
rect 5140 2640 5150 2720
rect 5050 2630 5150 2640
rect 5250 2720 5350 2730
rect 5250 2640 5260 2720
rect 5340 2640 5350 2720
rect 5250 2630 5350 2640
rect 5450 2720 5550 2730
rect 5450 2640 5460 2720
rect 5540 2640 5550 2720
rect 5450 2630 5550 2640
rect 5650 2720 5750 2730
rect 5650 2640 5660 2720
rect 5740 2640 5750 2720
rect 5650 2630 5750 2640
rect 5850 2720 5950 2730
rect 5850 2640 5860 2720
rect 5940 2640 5950 2720
rect 5850 2630 5950 2640
rect 6050 2720 6150 2730
rect 6050 2640 6060 2720
rect 6140 2640 6150 2720
rect 6050 2630 6150 2640
rect 6250 2720 6350 2730
rect 6250 2640 6260 2720
rect 6340 2640 6350 2720
rect 6250 2630 6350 2640
rect 6450 2720 6550 2730
rect 6450 2640 6460 2720
rect 6540 2640 6550 2720
rect 6450 2630 6550 2640
rect -115 2545 -85 2630
rect 85 2545 115 2630
rect 285 2545 315 2630
rect 485 2545 515 2630
rect 685 2545 715 2630
rect 885 2545 915 2630
rect 1085 2545 1115 2630
rect 1285 2545 1315 2630
rect 1485 2545 1515 2630
rect 1685 2545 1715 2630
rect 1885 2545 1915 2630
rect 2085 2545 2115 2630
rect 2285 2545 2315 2630
rect 2485 2545 2515 2630
rect 2685 2545 2715 2630
rect 2885 2545 2915 2630
rect 3085 2545 3115 2630
rect 3285 2545 3315 2630
rect 3485 2545 3515 2630
rect 3685 2545 3715 2630
rect 3885 2545 3915 2630
rect 4085 2545 4115 2630
rect 4285 2545 4315 2630
rect 4485 2545 4515 2630
rect 4685 2545 4715 2630
rect 4885 2545 4915 2630
rect 5085 2545 5115 2630
rect 5285 2545 5315 2630
rect 5485 2545 5515 2630
rect 5685 2545 5715 2630
rect 5885 2545 5915 2630
rect 6085 2545 6115 2630
rect 6285 2545 6315 2630
rect 6485 2545 6515 2630
rect -150 2535 -50 2545
rect -150 2455 -140 2535
rect -60 2455 -50 2535
rect -150 2445 -50 2455
rect 50 2535 150 2545
rect 50 2455 60 2535
rect 140 2455 150 2535
rect 50 2445 150 2455
rect 250 2535 350 2545
rect 250 2455 260 2535
rect 340 2455 350 2535
rect 250 2445 350 2455
rect 450 2535 550 2545
rect 450 2455 460 2535
rect 540 2455 550 2535
rect 450 2445 550 2455
rect 650 2535 750 2545
rect 650 2455 660 2535
rect 740 2455 750 2535
rect 650 2445 750 2455
rect 850 2535 950 2545
rect 850 2455 860 2535
rect 940 2455 950 2535
rect 850 2445 950 2455
rect 1050 2535 1150 2545
rect 1050 2455 1060 2535
rect 1140 2455 1150 2535
rect 1050 2445 1150 2455
rect 1250 2535 1350 2545
rect 1250 2455 1260 2535
rect 1340 2455 1350 2535
rect 1250 2445 1350 2455
rect 1450 2535 1550 2545
rect 1450 2455 1460 2535
rect 1540 2455 1550 2535
rect 1450 2445 1550 2455
rect 1650 2535 1750 2545
rect 1650 2455 1660 2535
rect 1740 2455 1750 2535
rect 1650 2445 1750 2455
rect 1850 2535 1950 2545
rect 1850 2455 1860 2535
rect 1940 2455 1950 2535
rect 1850 2445 1950 2455
rect 2050 2535 2150 2545
rect 2050 2455 2060 2535
rect 2140 2455 2150 2535
rect 2050 2445 2150 2455
rect 2250 2535 2350 2545
rect 2250 2455 2260 2535
rect 2340 2455 2350 2535
rect 2250 2445 2350 2455
rect 2450 2535 2550 2545
rect 2450 2455 2460 2535
rect 2540 2455 2550 2535
rect 2450 2445 2550 2455
rect 2650 2535 2750 2545
rect 2650 2455 2660 2535
rect 2740 2455 2750 2535
rect 2650 2445 2750 2455
rect 2850 2535 2950 2545
rect 2850 2455 2860 2535
rect 2940 2455 2950 2535
rect 2850 2445 2950 2455
rect 3050 2535 3150 2545
rect 3050 2455 3060 2535
rect 3140 2455 3150 2535
rect 3050 2445 3150 2455
rect 3250 2535 3350 2545
rect 3250 2455 3260 2535
rect 3340 2455 3350 2535
rect 3250 2445 3350 2455
rect 3450 2535 3550 2545
rect 3450 2455 3460 2535
rect 3540 2455 3550 2535
rect 3450 2445 3550 2455
rect 3650 2535 3750 2545
rect 3650 2455 3660 2535
rect 3740 2455 3750 2535
rect 3650 2445 3750 2455
rect 3850 2535 3950 2545
rect 3850 2455 3860 2535
rect 3940 2455 3950 2535
rect 3850 2445 3950 2455
rect 4050 2535 4150 2545
rect 4050 2455 4060 2535
rect 4140 2455 4150 2535
rect 4050 2445 4150 2455
rect 4250 2535 4350 2545
rect 4250 2455 4260 2535
rect 4340 2455 4350 2535
rect 4250 2445 4350 2455
rect 4450 2535 4550 2545
rect 4450 2455 4460 2535
rect 4540 2455 4550 2535
rect 4450 2445 4550 2455
rect 4650 2535 4750 2545
rect 4650 2455 4660 2535
rect 4740 2455 4750 2535
rect 4650 2445 4750 2455
rect 4850 2535 4950 2545
rect 4850 2455 4860 2535
rect 4940 2455 4950 2535
rect 4850 2445 4950 2455
rect 5050 2535 5150 2545
rect 5050 2455 5060 2535
rect 5140 2455 5150 2535
rect 5050 2445 5150 2455
rect 5250 2535 5350 2545
rect 5250 2455 5260 2535
rect 5340 2455 5350 2535
rect 5250 2445 5350 2455
rect 5450 2535 5550 2545
rect 5450 2455 5460 2535
rect 5540 2455 5550 2535
rect 5450 2445 5550 2455
rect 5650 2535 5750 2545
rect 5650 2455 5660 2535
rect 5740 2455 5750 2535
rect 5650 2445 5750 2455
rect 5850 2535 5950 2545
rect 5850 2455 5860 2535
rect 5940 2455 5950 2535
rect 5850 2445 5950 2455
rect 6050 2535 6150 2545
rect 6050 2455 6060 2535
rect 6140 2455 6150 2535
rect 6050 2445 6150 2455
rect 6250 2535 6350 2545
rect 6250 2455 6260 2535
rect 6340 2455 6350 2535
rect 6250 2445 6350 2455
rect 6450 2535 6550 2545
rect 6450 2455 6460 2535
rect 6540 2455 6550 2535
rect 6450 2445 6550 2455
rect -115 2360 -85 2445
rect 85 2360 115 2445
rect 285 2360 315 2445
rect 485 2360 515 2445
rect 685 2360 715 2445
rect 885 2360 915 2445
rect 1085 2360 1115 2445
rect 1285 2360 1315 2445
rect 1485 2360 1515 2445
rect 1685 2360 1715 2445
rect 1885 2360 1915 2445
rect 2085 2360 2115 2445
rect 2285 2360 2315 2445
rect 2485 2360 2515 2445
rect 2685 2360 2715 2445
rect 2885 2360 2915 2445
rect 3085 2360 3115 2445
rect 3285 2360 3315 2445
rect 3485 2360 3515 2445
rect 3685 2360 3715 2445
rect 3885 2360 3915 2445
rect 4085 2360 4115 2445
rect 4285 2360 4315 2445
rect 4485 2360 4515 2445
rect 4685 2360 4715 2445
rect 4885 2360 4915 2445
rect 5085 2360 5115 2445
rect 5285 2360 5315 2445
rect 5485 2360 5515 2445
rect 5685 2360 5715 2445
rect 5885 2360 5915 2445
rect 6085 2360 6115 2445
rect 6285 2360 6315 2445
rect 6485 2360 6515 2445
rect -150 2350 -50 2360
rect -150 2270 -140 2350
rect -60 2270 -50 2350
rect -150 2260 -50 2270
rect 50 2350 150 2360
rect 50 2270 60 2350
rect 140 2270 150 2350
rect 50 2260 150 2270
rect 250 2350 350 2360
rect 250 2270 260 2350
rect 340 2270 350 2350
rect 250 2260 350 2270
rect 450 2350 550 2360
rect 450 2270 460 2350
rect 540 2270 550 2350
rect 450 2260 550 2270
rect 650 2350 750 2360
rect 650 2270 660 2350
rect 740 2270 750 2350
rect 650 2260 750 2270
rect 850 2350 950 2360
rect 850 2270 860 2350
rect 940 2270 950 2350
rect 850 2260 950 2270
rect 1050 2350 1150 2360
rect 1050 2270 1060 2350
rect 1140 2270 1150 2350
rect 1050 2260 1150 2270
rect 1250 2350 1350 2360
rect 1250 2270 1260 2350
rect 1340 2270 1350 2350
rect 1250 2260 1350 2270
rect 1450 2350 1550 2360
rect 1450 2270 1460 2350
rect 1540 2270 1550 2350
rect 1450 2260 1550 2270
rect 1650 2350 1750 2360
rect 1650 2270 1660 2350
rect 1740 2270 1750 2350
rect 1650 2260 1750 2270
rect 1850 2350 1950 2360
rect 1850 2270 1860 2350
rect 1940 2270 1950 2350
rect 1850 2260 1950 2270
rect 2050 2350 2150 2360
rect 2050 2270 2060 2350
rect 2140 2270 2150 2350
rect 2050 2260 2150 2270
rect 2250 2350 2350 2360
rect 2250 2270 2260 2350
rect 2340 2270 2350 2350
rect 2250 2260 2350 2270
rect 2450 2350 2550 2360
rect 2450 2270 2460 2350
rect 2540 2270 2550 2350
rect 2450 2260 2550 2270
rect 2650 2350 2750 2360
rect 2650 2270 2660 2350
rect 2740 2270 2750 2350
rect 2650 2260 2750 2270
rect 2850 2350 2950 2360
rect 2850 2270 2860 2350
rect 2940 2270 2950 2350
rect 2850 2260 2950 2270
rect 3050 2350 3150 2360
rect 3050 2270 3060 2350
rect 3140 2270 3150 2350
rect 3050 2260 3150 2270
rect 3250 2350 3350 2360
rect 3250 2270 3260 2350
rect 3340 2270 3350 2350
rect 3250 2260 3350 2270
rect 3450 2350 3550 2360
rect 3450 2270 3460 2350
rect 3540 2270 3550 2350
rect 3450 2260 3550 2270
rect 3650 2350 3750 2360
rect 3650 2270 3660 2350
rect 3740 2270 3750 2350
rect 3650 2260 3750 2270
rect 3850 2350 3950 2360
rect 3850 2270 3860 2350
rect 3940 2270 3950 2350
rect 3850 2260 3950 2270
rect 4050 2350 4150 2360
rect 4050 2270 4060 2350
rect 4140 2270 4150 2350
rect 4050 2260 4150 2270
rect 4250 2350 4350 2360
rect 4250 2270 4260 2350
rect 4340 2270 4350 2350
rect 4250 2260 4350 2270
rect 4450 2350 4550 2360
rect 4450 2270 4460 2350
rect 4540 2270 4550 2350
rect 4450 2260 4550 2270
rect 4650 2350 4750 2360
rect 4650 2270 4660 2350
rect 4740 2270 4750 2350
rect 4650 2260 4750 2270
rect 4850 2350 4950 2360
rect 4850 2270 4860 2350
rect 4940 2270 4950 2350
rect 4850 2260 4950 2270
rect 5050 2350 5150 2360
rect 5050 2270 5060 2350
rect 5140 2270 5150 2350
rect 5050 2260 5150 2270
rect 5250 2350 5350 2360
rect 5250 2270 5260 2350
rect 5340 2270 5350 2350
rect 5250 2260 5350 2270
rect 5450 2350 5550 2360
rect 5450 2270 5460 2350
rect 5540 2270 5550 2350
rect 5450 2260 5550 2270
rect 5650 2350 5750 2360
rect 5650 2270 5660 2350
rect 5740 2270 5750 2350
rect 5650 2260 5750 2270
rect 5850 2350 5950 2360
rect 5850 2270 5860 2350
rect 5940 2270 5950 2350
rect 5850 2260 5950 2270
rect 6050 2350 6150 2360
rect 6050 2270 6060 2350
rect 6140 2270 6150 2350
rect 6050 2260 6150 2270
rect 6250 2350 6350 2360
rect 6250 2270 6260 2350
rect 6340 2270 6350 2350
rect 6250 2260 6350 2270
rect 6450 2350 6550 2360
rect 6450 2270 6460 2350
rect 6540 2270 6550 2350
rect 6450 2260 6550 2270
rect -115 2175 -85 2260
rect 85 2175 115 2260
rect 285 2175 315 2260
rect 485 2175 515 2260
rect 685 2175 715 2260
rect 885 2175 915 2260
rect 1085 2175 1115 2260
rect 1285 2175 1315 2260
rect 1485 2175 1515 2260
rect 1685 2175 1715 2260
rect 1885 2175 1915 2260
rect 2085 2175 2115 2260
rect 2285 2175 2315 2260
rect 2485 2175 2515 2260
rect 2685 2175 2715 2260
rect 2885 2175 2915 2260
rect 3085 2175 3115 2260
rect 3285 2175 3315 2260
rect 3485 2175 3515 2260
rect 3685 2175 3715 2260
rect 3885 2175 3915 2260
rect 4085 2175 4115 2260
rect 4285 2175 4315 2260
rect 4485 2175 4515 2260
rect 4685 2175 4715 2260
rect 4885 2175 4915 2260
rect 5085 2175 5115 2260
rect 5285 2175 5315 2260
rect 5485 2175 5515 2260
rect 5685 2175 5715 2260
rect 5885 2175 5915 2260
rect 6085 2175 6115 2260
rect 6285 2175 6315 2260
rect 6485 2175 6515 2260
rect -150 2165 -50 2175
rect -150 2085 -140 2165
rect -60 2085 -50 2165
rect -150 2075 -50 2085
rect 50 2165 150 2175
rect 50 2085 60 2165
rect 140 2085 150 2165
rect 50 2075 150 2085
rect 250 2165 350 2175
rect 250 2085 260 2165
rect 340 2085 350 2165
rect 250 2075 350 2085
rect 450 2165 550 2175
rect 450 2085 460 2165
rect 540 2085 550 2165
rect 450 2075 550 2085
rect 650 2165 750 2175
rect 650 2085 660 2165
rect 740 2085 750 2165
rect 650 2075 750 2085
rect 850 2165 950 2175
rect 850 2085 860 2165
rect 940 2085 950 2165
rect 850 2075 950 2085
rect 1050 2165 1150 2175
rect 1050 2085 1060 2165
rect 1140 2085 1150 2165
rect 1050 2075 1150 2085
rect 1250 2165 1350 2175
rect 1250 2085 1260 2165
rect 1340 2085 1350 2165
rect 1250 2075 1350 2085
rect 1450 2165 1550 2175
rect 1450 2085 1460 2165
rect 1540 2085 1550 2165
rect 1450 2075 1550 2085
rect 1650 2165 1750 2175
rect 1650 2085 1660 2165
rect 1740 2085 1750 2165
rect 1650 2075 1750 2085
rect 1850 2165 1950 2175
rect 1850 2085 1860 2165
rect 1940 2085 1950 2165
rect 1850 2075 1950 2085
rect 2050 2165 2150 2175
rect 2050 2085 2060 2165
rect 2140 2085 2150 2165
rect 2050 2075 2150 2085
rect 2250 2165 2350 2175
rect 2250 2085 2260 2165
rect 2340 2085 2350 2165
rect 2250 2075 2350 2085
rect 2450 2165 2550 2175
rect 2450 2085 2460 2165
rect 2540 2085 2550 2165
rect 2450 2075 2550 2085
rect 2650 2165 2750 2175
rect 2650 2085 2660 2165
rect 2740 2085 2750 2165
rect 2650 2075 2750 2085
rect 2850 2165 2950 2175
rect 2850 2085 2860 2165
rect 2940 2085 2950 2165
rect 2850 2075 2950 2085
rect 3050 2165 3150 2175
rect 3050 2085 3060 2165
rect 3140 2085 3150 2165
rect 3050 2075 3150 2085
rect 3250 2165 3350 2175
rect 3250 2085 3260 2165
rect 3340 2085 3350 2165
rect 3250 2075 3350 2085
rect 3450 2165 3550 2175
rect 3450 2085 3460 2165
rect 3540 2085 3550 2165
rect 3450 2075 3550 2085
rect 3650 2165 3750 2175
rect 3650 2085 3660 2165
rect 3740 2085 3750 2165
rect 3650 2075 3750 2085
rect 3850 2165 3950 2175
rect 3850 2085 3860 2165
rect 3940 2085 3950 2165
rect 3850 2075 3950 2085
rect 4050 2165 4150 2175
rect 4050 2085 4060 2165
rect 4140 2085 4150 2165
rect 4050 2075 4150 2085
rect 4250 2165 4350 2175
rect 4250 2085 4260 2165
rect 4340 2085 4350 2165
rect 4250 2075 4350 2085
rect 4450 2165 4550 2175
rect 4450 2085 4460 2165
rect 4540 2085 4550 2165
rect 4450 2075 4550 2085
rect 4650 2165 4750 2175
rect 4650 2085 4660 2165
rect 4740 2085 4750 2165
rect 4650 2075 4750 2085
rect 4850 2165 4950 2175
rect 4850 2085 4860 2165
rect 4940 2085 4950 2165
rect 4850 2075 4950 2085
rect 5050 2165 5150 2175
rect 5050 2085 5060 2165
rect 5140 2085 5150 2165
rect 5050 2075 5150 2085
rect 5250 2165 5350 2175
rect 5250 2085 5260 2165
rect 5340 2085 5350 2165
rect 5250 2075 5350 2085
rect 5450 2165 5550 2175
rect 5450 2085 5460 2165
rect 5540 2085 5550 2165
rect 5450 2075 5550 2085
rect 5650 2165 5750 2175
rect 5650 2085 5660 2165
rect 5740 2085 5750 2165
rect 5650 2075 5750 2085
rect 5850 2165 5950 2175
rect 5850 2085 5860 2165
rect 5940 2085 5950 2165
rect 5850 2075 5950 2085
rect 6050 2165 6150 2175
rect 6050 2085 6060 2165
rect 6140 2085 6150 2165
rect 6050 2075 6150 2085
rect 6250 2165 6350 2175
rect 6250 2085 6260 2165
rect 6340 2085 6350 2165
rect 6250 2075 6350 2085
rect 6450 2165 6550 2175
rect 6450 2085 6460 2165
rect 6540 2085 6550 2165
rect 6450 2075 6550 2085
rect -115 1990 -85 2075
rect 85 1990 115 2075
rect 285 1990 315 2075
rect 485 1990 515 2075
rect 685 1990 715 2075
rect 885 1990 915 2075
rect 1085 1990 1115 2075
rect 1285 1990 1315 2075
rect 1485 1990 1515 2075
rect 1685 1990 1715 2075
rect 1885 1990 1915 2075
rect 2085 1990 2115 2075
rect 2285 1990 2315 2075
rect 2485 1990 2515 2075
rect 2685 1990 2715 2075
rect 2885 1990 2915 2075
rect 3085 1990 3115 2075
rect 3285 1990 3315 2075
rect 3485 1990 3515 2075
rect 3685 1990 3715 2075
rect 3885 1990 3915 2075
rect 4085 1990 4115 2075
rect 4285 1990 4315 2075
rect 4485 1990 4515 2075
rect 4685 1990 4715 2075
rect 4885 1990 4915 2075
rect 5085 1990 5115 2075
rect 5285 1990 5315 2075
rect 5485 1990 5515 2075
rect 5685 1990 5715 2075
rect 5885 1990 5915 2075
rect 6085 1990 6115 2075
rect 6285 1990 6315 2075
rect 6485 1990 6515 2075
rect -150 1980 -50 1990
rect -150 1900 -140 1980
rect -60 1900 -50 1980
rect -150 1890 -50 1900
rect 50 1980 150 1990
rect 50 1900 60 1980
rect 140 1900 150 1980
rect 50 1890 150 1900
rect 250 1980 350 1990
rect 250 1900 260 1980
rect 340 1900 350 1980
rect 250 1890 350 1900
rect 450 1980 550 1990
rect 450 1900 460 1980
rect 540 1900 550 1980
rect 450 1890 550 1900
rect 650 1980 750 1990
rect 650 1900 660 1980
rect 740 1900 750 1980
rect 650 1890 750 1900
rect 850 1980 950 1990
rect 850 1900 860 1980
rect 940 1900 950 1980
rect 850 1890 950 1900
rect 1050 1980 1150 1990
rect 1050 1900 1060 1980
rect 1140 1900 1150 1980
rect 1050 1890 1150 1900
rect 1250 1980 1350 1990
rect 1250 1900 1260 1980
rect 1340 1900 1350 1980
rect 1250 1890 1350 1900
rect 1450 1980 1550 1990
rect 1450 1900 1460 1980
rect 1540 1900 1550 1980
rect 1450 1890 1550 1900
rect 1650 1980 1750 1990
rect 1650 1900 1660 1980
rect 1740 1900 1750 1980
rect 1650 1890 1750 1900
rect 1850 1980 1950 1990
rect 1850 1900 1860 1980
rect 1940 1900 1950 1980
rect 1850 1890 1950 1900
rect 2050 1980 2150 1990
rect 2050 1900 2060 1980
rect 2140 1900 2150 1980
rect 2050 1890 2150 1900
rect 2250 1980 2350 1990
rect 2250 1900 2260 1980
rect 2340 1900 2350 1980
rect 2250 1890 2350 1900
rect 2450 1980 2550 1990
rect 2450 1900 2460 1980
rect 2540 1900 2550 1980
rect 2450 1890 2550 1900
rect 2650 1980 2750 1990
rect 2650 1900 2660 1980
rect 2740 1900 2750 1980
rect 2650 1890 2750 1900
rect 2850 1980 2950 1990
rect 2850 1900 2860 1980
rect 2940 1900 2950 1980
rect 2850 1890 2950 1900
rect 3050 1980 3150 1990
rect 3050 1900 3060 1980
rect 3140 1900 3150 1980
rect 3050 1890 3150 1900
rect 3250 1980 3350 1990
rect 3250 1900 3260 1980
rect 3340 1900 3350 1980
rect 3250 1890 3350 1900
rect 3450 1980 3550 1990
rect 3450 1900 3460 1980
rect 3540 1900 3550 1980
rect 3450 1890 3550 1900
rect 3650 1980 3750 1990
rect 3650 1900 3660 1980
rect 3740 1900 3750 1980
rect 3650 1890 3750 1900
rect 3850 1980 3950 1990
rect 3850 1900 3860 1980
rect 3940 1900 3950 1980
rect 3850 1890 3950 1900
rect 4050 1980 4150 1990
rect 4050 1900 4060 1980
rect 4140 1900 4150 1980
rect 4050 1890 4150 1900
rect 4250 1980 4350 1990
rect 4250 1900 4260 1980
rect 4340 1900 4350 1980
rect 4250 1890 4350 1900
rect 4450 1980 4550 1990
rect 4450 1900 4460 1980
rect 4540 1900 4550 1980
rect 4450 1890 4550 1900
rect 4650 1980 4750 1990
rect 4650 1900 4660 1980
rect 4740 1900 4750 1980
rect 4650 1890 4750 1900
rect 4850 1980 4950 1990
rect 4850 1900 4860 1980
rect 4940 1900 4950 1980
rect 4850 1890 4950 1900
rect 5050 1980 5150 1990
rect 5050 1900 5060 1980
rect 5140 1900 5150 1980
rect 5050 1890 5150 1900
rect 5250 1980 5350 1990
rect 5250 1900 5260 1980
rect 5340 1900 5350 1980
rect 5250 1890 5350 1900
rect 5450 1980 5550 1990
rect 5450 1900 5460 1980
rect 5540 1900 5550 1980
rect 5450 1890 5550 1900
rect 5650 1980 5750 1990
rect 5650 1900 5660 1980
rect 5740 1900 5750 1980
rect 5650 1890 5750 1900
rect 5850 1980 5950 1990
rect 5850 1900 5860 1980
rect 5940 1900 5950 1980
rect 5850 1890 5950 1900
rect 6050 1980 6150 1990
rect 6050 1900 6060 1980
rect 6140 1900 6150 1980
rect 6050 1890 6150 1900
rect 6250 1980 6350 1990
rect 6250 1900 6260 1980
rect 6340 1900 6350 1980
rect 6250 1890 6350 1900
rect 6450 1980 6550 1990
rect 6450 1900 6460 1980
rect 6540 1900 6550 1980
rect 6450 1890 6550 1900
rect -115 1805 -85 1890
rect 85 1805 115 1890
rect 285 1805 315 1890
rect 485 1805 515 1890
rect 685 1805 715 1890
rect 885 1805 915 1890
rect 1085 1805 1115 1890
rect 1285 1805 1315 1890
rect 1485 1805 1515 1890
rect 1685 1805 1715 1890
rect 1885 1805 1915 1890
rect 2085 1805 2115 1890
rect 2285 1805 2315 1890
rect 2485 1805 2515 1890
rect 2685 1805 2715 1890
rect 2885 1805 2915 1890
rect 3085 1805 3115 1890
rect 3285 1805 3315 1890
rect 3485 1805 3515 1890
rect 3685 1805 3715 1890
rect 3885 1805 3915 1890
rect 4085 1805 4115 1890
rect 4285 1805 4315 1890
rect 4485 1805 4515 1890
rect 4685 1805 4715 1890
rect 4885 1805 4915 1890
rect 5085 1805 5115 1890
rect 5285 1805 5315 1890
rect 5485 1805 5515 1890
rect 5685 1805 5715 1890
rect 5885 1805 5915 1890
rect 6085 1805 6115 1890
rect 6285 1805 6315 1890
rect 6485 1805 6515 1890
rect -150 1795 -50 1805
rect -150 1715 -140 1795
rect -60 1715 -50 1795
rect -150 1705 -50 1715
rect 50 1795 150 1805
rect 50 1715 60 1795
rect 140 1715 150 1795
rect 50 1705 150 1715
rect 250 1795 350 1805
rect 250 1715 260 1795
rect 340 1715 350 1795
rect 250 1705 350 1715
rect 450 1795 550 1805
rect 450 1715 460 1795
rect 540 1715 550 1795
rect 450 1705 550 1715
rect 650 1795 750 1805
rect 650 1715 660 1795
rect 740 1715 750 1795
rect 650 1705 750 1715
rect 850 1795 950 1805
rect 850 1715 860 1795
rect 940 1715 950 1795
rect 850 1705 950 1715
rect 1050 1795 1150 1805
rect 1050 1715 1060 1795
rect 1140 1715 1150 1795
rect 1050 1705 1150 1715
rect 1250 1795 1350 1805
rect 1250 1715 1260 1795
rect 1340 1715 1350 1795
rect 1250 1705 1350 1715
rect 1450 1795 1550 1805
rect 1450 1715 1460 1795
rect 1540 1715 1550 1795
rect 1450 1705 1550 1715
rect 1650 1795 1750 1805
rect 1650 1715 1660 1795
rect 1740 1715 1750 1795
rect 1650 1705 1750 1715
rect 1850 1795 1950 1805
rect 1850 1715 1860 1795
rect 1940 1715 1950 1795
rect 1850 1705 1950 1715
rect 2050 1795 2150 1805
rect 2050 1715 2060 1795
rect 2140 1715 2150 1795
rect 2050 1705 2150 1715
rect 2250 1795 2350 1805
rect 2250 1715 2260 1795
rect 2340 1715 2350 1795
rect 2250 1705 2350 1715
rect 2450 1795 2550 1805
rect 2450 1715 2460 1795
rect 2540 1715 2550 1795
rect 2450 1705 2550 1715
rect 2650 1795 2750 1805
rect 2650 1715 2660 1795
rect 2740 1715 2750 1795
rect 2650 1705 2750 1715
rect 2850 1795 2950 1805
rect 2850 1715 2860 1795
rect 2940 1715 2950 1795
rect 2850 1705 2950 1715
rect 3050 1795 3150 1805
rect 3050 1715 3060 1795
rect 3140 1715 3150 1795
rect 3050 1705 3150 1715
rect 3250 1795 3350 1805
rect 3250 1715 3260 1795
rect 3340 1715 3350 1795
rect 3250 1705 3350 1715
rect 3450 1795 3550 1805
rect 3450 1715 3460 1795
rect 3540 1715 3550 1795
rect 3450 1705 3550 1715
rect 3650 1795 3750 1805
rect 3650 1715 3660 1795
rect 3740 1715 3750 1795
rect 3650 1705 3750 1715
rect 3850 1795 3950 1805
rect 3850 1715 3860 1795
rect 3940 1715 3950 1795
rect 3850 1705 3950 1715
rect 4050 1795 4150 1805
rect 4050 1715 4060 1795
rect 4140 1715 4150 1795
rect 4050 1705 4150 1715
rect 4250 1795 4350 1805
rect 4250 1715 4260 1795
rect 4340 1715 4350 1795
rect 4250 1705 4350 1715
rect 4450 1795 4550 1805
rect 4450 1715 4460 1795
rect 4540 1715 4550 1795
rect 4450 1705 4550 1715
rect 4650 1795 4750 1805
rect 4650 1715 4660 1795
rect 4740 1715 4750 1795
rect 4650 1705 4750 1715
rect 4850 1795 4950 1805
rect 4850 1715 4860 1795
rect 4940 1715 4950 1795
rect 4850 1705 4950 1715
rect 5050 1795 5150 1805
rect 5050 1715 5060 1795
rect 5140 1715 5150 1795
rect 5050 1705 5150 1715
rect 5250 1795 5350 1805
rect 5250 1715 5260 1795
rect 5340 1715 5350 1795
rect 5250 1705 5350 1715
rect 5450 1795 5550 1805
rect 5450 1715 5460 1795
rect 5540 1715 5550 1795
rect 5450 1705 5550 1715
rect 5650 1795 5750 1805
rect 5650 1715 5660 1795
rect 5740 1715 5750 1795
rect 5650 1705 5750 1715
rect 5850 1795 5950 1805
rect 5850 1715 5860 1795
rect 5940 1715 5950 1795
rect 5850 1705 5950 1715
rect 6050 1795 6150 1805
rect 6050 1715 6060 1795
rect 6140 1715 6150 1795
rect 6050 1705 6150 1715
rect 6250 1795 6350 1805
rect 6250 1715 6260 1795
rect 6340 1715 6350 1795
rect 6250 1705 6350 1715
rect 6450 1795 6550 1805
rect 6450 1715 6460 1795
rect 6540 1715 6550 1795
rect 6450 1705 6550 1715
rect -115 1620 -85 1705
rect 85 1620 115 1705
rect 285 1620 315 1705
rect 485 1620 515 1705
rect 685 1620 715 1705
rect 885 1620 915 1705
rect 1085 1620 1115 1705
rect 1285 1620 1315 1705
rect 1485 1620 1515 1705
rect 1685 1620 1715 1705
rect 1885 1620 1915 1705
rect 2085 1620 2115 1705
rect 2285 1620 2315 1705
rect 2485 1620 2515 1705
rect 2685 1620 2715 1705
rect 2885 1620 2915 1705
rect 3085 1620 3115 1705
rect 3285 1620 3315 1705
rect 3485 1620 3515 1705
rect 3685 1620 3715 1705
rect 3885 1620 3915 1705
rect 4085 1620 4115 1705
rect 4285 1620 4315 1705
rect 4485 1620 4515 1705
rect 4685 1620 4715 1705
rect 4885 1620 4915 1705
rect 5085 1620 5115 1705
rect 5285 1620 5315 1705
rect 5485 1620 5515 1705
rect 5685 1620 5715 1705
rect 5885 1620 5915 1705
rect 6085 1620 6115 1705
rect 6285 1620 6315 1705
rect 6485 1620 6515 1705
rect -150 1610 -50 1620
rect -150 1530 -140 1610
rect -60 1530 -50 1610
rect -150 1520 -50 1530
rect 50 1610 150 1620
rect 50 1530 60 1610
rect 140 1530 150 1610
rect 50 1520 150 1530
rect 250 1610 350 1620
rect 250 1530 260 1610
rect 340 1530 350 1610
rect 250 1520 350 1530
rect 450 1610 550 1620
rect 450 1530 460 1610
rect 540 1530 550 1610
rect 450 1520 550 1530
rect 650 1610 750 1620
rect 650 1530 660 1610
rect 740 1530 750 1610
rect 650 1520 750 1530
rect 850 1610 950 1620
rect 850 1530 860 1610
rect 940 1530 950 1610
rect 850 1520 950 1530
rect 1050 1610 1150 1620
rect 1050 1530 1060 1610
rect 1140 1530 1150 1610
rect 1050 1520 1150 1530
rect 1250 1610 1350 1620
rect 1250 1530 1260 1610
rect 1340 1530 1350 1610
rect 1250 1520 1350 1530
rect 1450 1610 1550 1620
rect 1450 1530 1460 1610
rect 1540 1530 1550 1610
rect 1450 1520 1550 1530
rect 1650 1610 1750 1620
rect 1650 1530 1660 1610
rect 1740 1530 1750 1610
rect 1650 1520 1750 1530
rect 1850 1610 1950 1620
rect 1850 1530 1860 1610
rect 1940 1530 1950 1610
rect 1850 1520 1950 1530
rect 2050 1610 2150 1620
rect 2050 1530 2060 1610
rect 2140 1530 2150 1610
rect 2050 1520 2150 1530
rect 2250 1610 2350 1620
rect 2250 1530 2260 1610
rect 2340 1530 2350 1610
rect 2250 1520 2350 1530
rect 2450 1610 2550 1620
rect 2450 1530 2460 1610
rect 2540 1530 2550 1610
rect 2450 1520 2550 1530
rect 2650 1610 2750 1620
rect 2650 1530 2660 1610
rect 2740 1530 2750 1610
rect 2650 1520 2750 1530
rect 2850 1610 2950 1620
rect 2850 1530 2860 1610
rect 2940 1530 2950 1610
rect 2850 1520 2950 1530
rect 3050 1610 3150 1620
rect 3050 1530 3060 1610
rect 3140 1530 3150 1610
rect 3050 1520 3150 1530
rect 3250 1610 3350 1620
rect 3250 1530 3260 1610
rect 3340 1530 3350 1610
rect 3250 1520 3350 1530
rect 3450 1610 3550 1620
rect 3450 1530 3460 1610
rect 3540 1530 3550 1610
rect 3450 1520 3550 1530
rect 3650 1610 3750 1620
rect 3650 1530 3660 1610
rect 3740 1530 3750 1610
rect 3650 1520 3750 1530
rect 3850 1610 3950 1620
rect 3850 1530 3860 1610
rect 3940 1530 3950 1610
rect 3850 1520 3950 1530
rect 4050 1610 4150 1620
rect 4050 1530 4060 1610
rect 4140 1530 4150 1610
rect 4050 1520 4150 1530
rect 4250 1610 4350 1620
rect 4250 1530 4260 1610
rect 4340 1530 4350 1610
rect 4250 1520 4350 1530
rect 4450 1610 4550 1620
rect 4450 1530 4460 1610
rect 4540 1530 4550 1610
rect 4450 1520 4550 1530
rect 4650 1610 4750 1620
rect 4650 1530 4660 1610
rect 4740 1530 4750 1610
rect 4650 1520 4750 1530
rect 4850 1610 4950 1620
rect 4850 1530 4860 1610
rect 4940 1530 4950 1610
rect 4850 1520 4950 1530
rect 5050 1610 5150 1620
rect 5050 1530 5060 1610
rect 5140 1530 5150 1610
rect 5050 1520 5150 1530
rect 5250 1610 5350 1620
rect 5250 1530 5260 1610
rect 5340 1530 5350 1610
rect 5250 1520 5350 1530
rect 5450 1610 5550 1620
rect 5450 1530 5460 1610
rect 5540 1530 5550 1610
rect 5450 1520 5550 1530
rect 5650 1610 5750 1620
rect 5650 1530 5660 1610
rect 5740 1530 5750 1610
rect 5650 1520 5750 1530
rect 5850 1610 5950 1620
rect 5850 1530 5860 1610
rect 5940 1530 5950 1610
rect 5850 1520 5950 1530
rect 6050 1610 6150 1620
rect 6050 1530 6060 1610
rect 6140 1530 6150 1610
rect 6050 1520 6150 1530
rect 6250 1610 6350 1620
rect 6250 1530 6260 1610
rect 6340 1530 6350 1610
rect 6250 1520 6350 1530
rect 6450 1610 6550 1620
rect 6450 1530 6460 1610
rect 6540 1530 6550 1610
rect 6450 1520 6550 1530
rect -115 1435 -85 1520
rect 85 1435 115 1520
rect 285 1435 315 1520
rect 485 1435 515 1520
rect 685 1435 715 1520
rect 885 1435 915 1520
rect 1085 1435 1115 1520
rect 1285 1435 1315 1520
rect 1485 1435 1515 1520
rect 1685 1435 1715 1520
rect 1885 1435 1915 1520
rect 2085 1435 2115 1520
rect 2285 1435 2315 1520
rect 2485 1435 2515 1520
rect 2685 1435 2715 1520
rect 2885 1435 2915 1520
rect 3085 1435 3115 1520
rect 3285 1435 3315 1520
rect 3485 1435 3515 1520
rect 3685 1435 3715 1520
rect 3885 1435 3915 1520
rect 4085 1435 4115 1520
rect 4285 1435 4315 1520
rect 4485 1435 4515 1520
rect 4685 1435 4715 1520
rect 4885 1435 4915 1520
rect 5085 1435 5115 1520
rect 5285 1435 5315 1520
rect 5485 1435 5515 1520
rect 5685 1435 5715 1520
rect 5885 1435 5915 1520
rect 6085 1435 6115 1520
rect 6285 1435 6315 1520
rect 6485 1435 6515 1520
rect -150 1425 -50 1435
rect -150 1345 -140 1425
rect -60 1345 -50 1425
rect -150 1335 -50 1345
rect 50 1425 150 1435
rect 50 1345 60 1425
rect 140 1345 150 1425
rect 50 1335 150 1345
rect 250 1425 350 1435
rect 250 1345 260 1425
rect 340 1345 350 1425
rect 250 1335 350 1345
rect 450 1425 550 1435
rect 450 1345 460 1425
rect 540 1345 550 1425
rect 450 1335 550 1345
rect 650 1425 750 1435
rect 650 1345 660 1425
rect 740 1345 750 1425
rect 650 1335 750 1345
rect 850 1425 950 1435
rect 850 1345 860 1425
rect 940 1345 950 1425
rect 850 1335 950 1345
rect 1050 1425 1150 1435
rect 1050 1345 1060 1425
rect 1140 1345 1150 1425
rect 1050 1335 1150 1345
rect 1250 1425 1350 1435
rect 1250 1345 1260 1425
rect 1340 1345 1350 1425
rect 1250 1335 1350 1345
rect 1450 1425 1550 1435
rect 1450 1345 1460 1425
rect 1540 1345 1550 1425
rect 1450 1335 1550 1345
rect 1650 1425 1750 1435
rect 1650 1345 1660 1425
rect 1740 1345 1750 1425
rect 1650 1335 1750 1345
rect 1850 1425 1950 1435
rect 1850 1345 1860 1425
rect 1940 1345 1950 1425
rect 1850 1335 1950 1345
rect 2050 1425 2150 1435
rect 2050 1345 2060 1425
rect 2140 1345 2150 1425
rect 2050 1335 2150 1345
rect 2250 1425 2350 1435
rect 2250 1345 2260 1425
rect 2340 1345 2350 1425
rect 2250 1335 2350 1345
rect 2450 1425 2550 1435
rect 2450 1345 2460 1425
rect 2540 1345 2550 1425
rect 2450 1335 2550 1345
rect 2650 1425 2750 1435
rect 2650 1345 2660 1425
rect 2740 1345 2750 1425
rect 2650 1335 2750 1345
rect 2850 1425 2950 1435
rect 2850 1345 2860 1425
rect 2940 1345 2950 1425
rect 2850 1335 2950 1345
rect 3050 1425 3150 1435
rect 3050 1345 3060 1425
rect 3140 1345 3150 1425
rect 3050 1335 3150 1345
rect 3250 1425 3350 1435
rect 3250 1345 3260 1425
rect 3340 1345 3350 1425
rect 3250 1335 3350 1345
rect 3450 1425 3550 1435
rect 3450 1345 3460 1425
rect 3540 1345 3550 1425
rect 3450 1335 3550 1345
rect 3650 1425 3750 1435
rect 3650 1345 3660 1425
rect 3740 1345 3750 1425
rect 3650 1335 3750 1345
rect 3850 1425 3950 1435
rect 3850 1345 3860 1425
rect 3940 1345 3950 1425
rect 3850 1335 3950 1345
rect 4050 1425 4150 1435
rect 4050 1345 4060 1425
rect 4140 1345 4150 1425
rect 4050 1335 4150 1345
rect 4250 1425 4350 1435
rect 4250 1345 4260 1425
rect 4340 1345 4350 1425
rect 4250 1335 4350 1345
rect 4450 1425 4550 1435
rect 4450 1345 4460 1425
rect 4540 1345 4550 1425
rect 4450 1335 4550 1345
rect 4650 1425 4750 1435
rect 4650 1345 4660 1425
rect 4740 1345 4750 1425
rect 4650 1335 4750 1345
rect 4850 1425 4950 1435
rect 4850 1345 4860 1425
rect 4940 1345 4950 1425
rect 4850 1335 4950 1345
rect 5050 1425 5150 1435
rect 5050 1345 5060 1425
rect 5140 1345 5150 1425
rect 5050 1335 5150 1345
rect 5250 1425 5350 1435
rect 5250 1345 5260 1425
rect 5340 1345 5350 1425
rect 5250 1335 5350 1345
rect 5450 1425 5550 1435
rect 5450 1345 5460 1425
rect 5540 1345 5550 1425
rect 5450 1335 5550 1345
rect 5650 1425 5750 1435
rect 5650 1345 5660 1425
rect 5740 1345 5750 1425
rect 5650 1335 5750 1345
rect 5850 1425 5950 1435
rect 5850 1345 5860 1425
rect 5940 1345 5950 1425
rect 5850 1335 5950 1345
rect 6050 1425 6150 1435
rect 6050 1345 6060 1425
rect 6140 1345 6150 1425
rect 6050 1335 6150 1345
rect 6250 1425 6350 1435
rect 6250 1345 6260 1425
rect 6340 1345 6350 1425
rect 6250 1335 6350 1345
rect 6450 1425 6550 1435
rect 6450 1345 6460 1425
rect 6540 1345 6550 1425
rect 6450 1335 6550 1345
rect -115 1250 -85 1335
rect 85 1250 115 1335
rect 285 1250 315 1335
rect 485 1250 515 1335
rect 685 1250 715 1335
rect 885 1250 915 1335
rect 1085 1250 1115 1335
rect 1285 1250 1315 1335
rect 1485 1250 1515 1335
rect 1685 1250 1715 1335
rect 1885 1250 1915 1335
rect 2085 1250 2115 1335
rect 2285 1250 2315 1335
rect 2485 1250 2515 1335
rect 2685 1250 2715 1335
rect 2885 1250 2915 1335
rect 3085 1250 3115 1335
rect 3285 1250 3315 1335
rect 3485 1250 3515 1335
rect 3685 1250 3715 1335
rect 3885 1250 3915 1335
rect 4085 1250 4115 1335
rect 4285 1250 4315 1335
rect 4485 1250 4515 1335
rect 4685 1250 4715 1335
rect 4885 1250 4915 1335
rect 5085 1250 5115 1335
rect 5285 1250 5315 1335
rect 5485 1250 5515 1335
rect 5685 1250 5715 1335
rect 5885 1250 5915 1335
rect 6085 1250 6115 1335
rect 6285 1250 6315 1335
rect 6485 1250 6515 1335
rect -150 1240 -50 1250
rect -150 1160 -140 1240
rect -60 1160 -50 1240
rect -150 1150 -50 1160
rect 50 1240 150 1250
rect 50 1160 60 1240
rect 140 1160 150 1240
rect 50 1150 150 1160
rect 250 1240 350 1250
rect 250 1160 260 1240
rect 340 1160 350 1240
rect 250 1150 350 1160
rect 450 1240 550 1250
rect 450 1160 460 1240
rect 540 1160 550 1240
rect 450 1150 550 1160
rect 650 1240 750 1250
rect 650 1160 660 1240
rect 740 1160 750 1240
rect 650 1150 750 1160
rect 850 1240 950 1250
rect 850 1160 860 1240
rect 940 1160 950 1240
rect 850 1150 950 1160
rect 1050 1240 1150 1250
rect 1050 1160 1060 1240
rect 1140 1160 1150 1240
rect 1050 1150 1150 1160
rect 1250 1240 1350 1250
rect 1250 1160 1260 1240
rect 1340 1160 1350 1240
rect 1250 1150 1350 1160
rect 1450 1240 1550 1250
rect 1450 1160 1460 1240
rect 1540 1160 1550 1240
rect 1450 1150 1550 1160
rect 1650 1240 1750 1250
rect 1650 1160 1660 1240
rect 1740 1160 1750 1240
rect 1650 1150 1750 1160
rect 1850 1240 1950 1250
rect 1850 1160 1860 1240
rect 1940 1160 1950 1240
rect 1850 1150 1950 1160
rect 2050 1240 2150 1250
rect 2050 1160 2060 1240
rect 2140 1160 2150 1240
rect 2050 1150 2150 1160
rect 2250 1240 2350 1250
rect 2250 1160 2260 1240
rect 2340 1160 2350 1240
rect 2250 1150 2350 1160
rect 2450 1240 2550 1250
rect 2450 1160 2460 1240
rect 2540 1160 2550 1240
rect 2450 1150 2550 1160
rect 2650 1240 2750 1250
rect 2650 1160 2660 1240
rect 2740 1160 2750 1240
rect 2650 1150 2750 1160
rect 2850 1240 2950 1250
rect 2850 1160 2860 1240
rect 2940 1160 2950 1240
rect 2850 1150 2950 1160
rect 3050 1240 3150 1250
rect 3050 1160 3060 1240
rect 3140 1160 3150 1240
rect 3050 1150 3150 1160
rect 3250 1240 3350 1250
rect 3250 1160 3260 1240
rect 3340 1160 3350 1240
rect 3250 1150 3350 1160
rect 3450 1240 3550 1250
rect 3450 1160 3460 1240
rect 3540 1160 3550 1240
rect 3450 1150 3550 1160
rect 3650 1240 3750 1250
rect 3650 1160 3660 1240
rect 3740 1160 3750 1240
rect 3650 1150 3750 1160
rect 3850 1240 3950 1250
rect 3850 1160 3860 1240
rect 3940 1160 3950 1240
rect 3850 1150 3950 1160
rect 4050 1240 4150 1250
rect 4050 1160 4060 1240
rect 4140 1160 4150 1240
rect 4050 1150 4150 1160
rect 4250 1240 4350 1250
rect 4250 1160 4260 1240
rect 4340 1160 4350 1240
rect 4250 1150 4350 1160
rect 4450 1240 4550 1250
rect 4450 1160 4460 1240
rect 4540 1160 4550 1240
rect 4450 1150 4550 1160
rect 4650 1240 4750 1250
rect 4650 1160 4660 1240
rect 4740 1160 4750 1240
rect 4650 1150 4750 1160
rect 4850 1240 4950 1250
rect 4850 1160 4860 1240
rect 4940 1160 4950 1240
rect 4850 1150 4950 1160
rect 5050 1240 5150 1250
rect 5050 1160 5060 1240
rect 5140 1160 5150 1240
rect 5050 1150 5150 1160
rect 5250 1240 5350 1250
rect 5250 1160 5260 1240
rect 5340 1160 5350 1240
rect 5250 1150 5350 1160
rect 5450 1240 5550 1250
rect 5450 1160 5460 1240
rect 5540 1160 5550 1240
rect 5450 1150 5550 1160
rect 5650 1240 5750 1250
rect 5650 1160 5660 1240
rect 5740 1160 5750 1240
rect 5650 1150 5750 1160
rect 5850 1240 5950 1250
rect 5850 1160 5860 1240
rect 5940 1160 5950 1240
rect 5850 1150 5950 1160
rect 6050 1240 6150 1250
rect 6050 1160 6060 1240
rect 6140 1160 6150 1240
rect 6050 1150 6150 1160
rect 6250 1240 6350 1250
rect 6250 1160 6260 1240
rect 6340 1160 6350 1240
rect 6250 1150 6350 1160
rect 6450 1240 6550 1250
rect 6450 1160 6460 1240
rect 6540 1160 6550 1240
rect 6450 1150 6550 1160
rect -115 1065 -85 1150
rect 85 1065 115 1150
rect 285 1065 315 1150
rect 485 1065 515 1150
rect 685 1065 715 1150
rect 885 1065 915 1150
rect 1085 1065 1115 1150
rect 1285 1065 1315 1150
rect 1485 1065 1515 1150
rect 1685 1065 1715 1150
rect 1885 1065 1915 1150
rect 2085 1065 2115 1150
rect 2285 1065 2315 1150
rect 2485 1065 2515 1150
rect 2685 1065 2715 1150
rect 2885 1065 2915 1150
rect 3085 1065 3115 1150
rect 3285 1065 3315 1150
rect 3485 1065 3515 1150
rect 3685 1065 3715 1150
rect 3885 1065 3915 1150
rect 4085 1065 4115 1150
rect 4285 1065 4315 1150
rect 4485 1065 4515 1150
rect 4685 1065 4715 1150
rect 4885 1065 4915 1150
rect 5085 1065 5115 1150
rect 5285 1065 5315 1150
rect 5485 1065 5515 1150
rect 5685 1065 5715 1150
rect 5885 1065 5915 1150
rect 6085 1065 6115 1150
rect 6285 1065 6315 1150
rect 6485 1065 6515 1150
rect -150 1055 -50 1065
rect -150 975 -140 1055
rect -60 975 -50 1055
rect -150 965 -50 975
rect 50 1055 150 1065
rect 50 975 60 1055
rect 140 975 150 1055
rect 50 965 150 975
rect 250 1055 350 1065
rect 250 975 260 1055
rect 340 975 350 1055
rect 250 965 350 975
rect 450 1055 550 1065
rect 450 975 460 1055
rect 540 975 550 1055
rect 450 965 550 975
rect 650 1055 750 1065
rect 650 975 660 1055
rect 740 975 750 1055
rect 650 965 750 975
rect 850 1055 950 1065
rect 850 975 860 1055
rect 940 975 950 1055
rect 850 965 950 975
rect 1050 1055 1150 1065
rect 1050 975 1060 1055
rect 1140 975 1150 1055
rect 1050 965 1150 975
rect 1250 1055 1350 1065
rect 1250 975 1260 1055
rect 1340 975 1350 1055
rect 1250 965 1350 975
rect 1450 1055 1550 1065
rect 1450 975 1460 1055
rect 1540 975 1550 1055
rect 1450 965 1550 975
rect 1650 1055 1750 1065
rect 1650 975 1660 1055
rect 1740 975 1750 1055
rect 1650 965 1750 975
rect 1850 1055 1950 1065
rect 1850 975 1860 1055
rect 1940 975 1950 1055
rect 1850 965 1950 975
rect 2050 1055 2150 1065
rect 2050 975 2060 1055
rect 2140 975 2150 1055
rect 2050 965 2150 975
rect 2250 1055 2350 1065
rect 2250 975 2260 1055
rect 2340 975 2350 1055
rect 2250 965 2350 975
rect 2450 1055 2550 1065
rect 2450 975 2460 1055
rect 2540 975 2550 1055
rect 2450 965 2550 975
rect 2650 1055 2750 1065
rect 2650 975 2660 1055
rect 2740 975 2750 1055
rect 2650 965 2750 975
rect 2850 1055 2950 1065
rect 2850 975 2860 1055
rect 2940 975 2950 1055
rect 2850 965 2950 975
rect 3050 1055 3150 1065
rect 3050 975 3060 1055
rect 3140 975 3150 1055
rect 3050 965 3150 975
rect 3250 1055 3350 1065
rect 3250 975 3260 1055
rect 3340 975 3350 1055
rect 3250 965 3350 975
rect 3450 1055 3550 1065
rect 3450 975 3460 1055
rect 3540 975 3550 1055
rect 3450 965 3550 975
rect 3650 1055 3750 1065
rect 3650 975 3660 1055
rect 3740 975 3750 1055
rect 3650 965 3750 975
rect 3850 1055 3950 1065
rect 3850 975 3860 1055
rect 3940 975 3950 1055
rect 3850 965 3950 975
rect 4050 1055 4150 1065
rect 4050 975 4060 1055
rect 4140 975 4150 1055
rect 4050 965 4150 975
rect 4250 1055 4350 1065
rect 4250 975 4260 1055
rect 4340 975 4350 1055
rect 4250 965 4350 975
rect 4450 1055 4550 1065
rect 4450 975 4460 1055
rect 4540 975 4550 1055
rect 4450 965 4550 975
rect 4650 1055 4750 1065
rect 4650 975 4660 1055
rect 4740 975 4750 1055
rect 4650 965 4750 975
rect 4850 1055 4950 1065
rect 4850 975 4860 1055
rect 4940 975 4950 1055
rect 4850 965 4950 975
rect 5050 1055 5150 1065
rect 5050 975 5060 1055
rect 5140 975 5150 1055
rect 5050 965 5150 975
rect 5250 1055 5350 1065
rect 5250 975 5260 1055
rect 5340 975 5350 1055
rect 5250 965 5350 975
rect 5450 1055 5550 1065
rect 5450 975 5460 1055
rect 5540 975 5550 1055
rect 5450 965 5550 975
rect 5650 1055 5750 1065
rect 5650 975 5660 1055
rect 5740 975 5750 1055
rect 5650 965 5750 975
rect 5850 1055 5950 1065
rect 5850 975 5860 1055
rect 5940 975 5950 1055
rect 5850 965 5950 975
rect 6050 1055 6150 1065
rect 6050 975 6060 1055
rect 6140 975 6150 1055
rect 6050 965 6150 975
rect 6250 1055 6350 1065
rect 6250 975 6260 1055
rect 6340 975 6350 1055
rect 6250 965 6350 975
rect 6450 1055 6550 1065
rect 6450 975 6460 1055
rect 6540 975 6550 1055
rect 6450 965 6550 975
rect -115 880 -85 965
rect 85 880 115 965
rect 285 880 315 965
rect 485 880 515 965
rect 685 880 715 965
rect 885 880 915 965
rect 1085 880 1115 965
rect 1285 880 1315 965
rect 1485 880 1515 965
rect 1685 880 1715 965
rect 1885 880 1915 965
rect 2085 880 2115 965
rect 2285 880 2315 965
rect 2485 880 2515 965
rect 2685 880 2715 965
rect 2885 880 2915 965
rect 3085 880 3115 965
rect 3285 880 3315 965
rect 3485 880 3515 965
rect 3685 880 3715 965
rect 3885 880 3915 965
rect 4085 880 4115 965
rect 4285 880 4315 965
rect 4485 880 4515 965
rect 4685 880 4715 965
rect 4885 880 4915 965
rect 5085 880 5115 965
rect 5285 880 5315 965
rect 5485 880 5515 965
rect 5685 880 5715 965
rect 5885 880 5915 965
rect 6085 880 6115 965
rect 6285 880 6315 965
rect 6485 880 6515 965
rect -150 870 -50 880
rect -150 790 -140 870
rect -60 790 -50 870
rect -150 780 -50 790
rect 50 870 150 880
rect 50 790 60 870
rect 140 790 150 870
rect 50 780 150 790
rect 250 870 350 880
rect 250 790 260 870
rect 340 790 350 870
rect 250 780 350 790
rect 450 870 550 880
rect 450 790 460 870
rect 540 790 550 870
rect 450 780 550 790
rect 650 870 750 880
rect 650 790 660 870
rect 740 790 750 870
rect 650 780 750 790
rect 850 870 950 880
rect 850 790 860 870
rect 940 790 950 870
rect 850 780 950 790
rect 1050 870 1150 880
rect 1050 790 1060 870
rect 1140 790 1150 870
rect 1050 780 1150 790
rect 1250 870 1350 880
rect 1250 790 1260 870
rect 1340 790 1350 870
rect 1250 780 1350 790
rect 1450 870 1550 880
rect 1450 790 1460 870
rect 1540 790 1550 870
rect 1450 780 1550 790
rect 1650 870 1750 880
rect 1650 790 1660 870
rect 1740 790 1750 870
rect 1650 780 1750 790
rect 1850 870 1950 880
rect 1850 790 1860 870
rect 1940 790 1950 870
rect 1850 780 1950 790
rect 2050 870 2150 880
rect 2050 790 2060 870
rect 2140 790 2150 870
rect 2050 780 2150 790
rect 2250 870 2350 880
rect 2250 790 2260 870
rect 2340 790 2350 870
rect 2250 780 2350 790
rect 2450 870 2550 880
rect 2450 790 2460 870
rect 2540 790 2550 870
rect 2450 780 2550 790
rect 2650 870 2750 880
rect 2650 790 2660 870
rect 2740 790 2750 870
rect 2650 780 2750 790
rect 2850 870 2950 880
rect 2850 790 2860 870
rect 2940 790 2950 870
rect 2850 780 2950 790
rect 3050 870 3150 880
rect 3050 790 3060 870
rect 3140 790 3150 870
rect 3050 780 3150 790
rect 3250 870 3350 880
rect 3250 790 3260 870
rect 3340 790 3350 870
rect 3250 780 3350 790
rect 3450 870 3550 880
rect 3450 790 3460 870
rect 3540 790 3550 870
rect 3450 780 3550 790
rect 3650 870 3750 880
rect 3650 790 3660 870
rect 3740 790 3750 870
rect 3650 780 3750 790
rect 3850 870 3950 880
rect 3850 790 3860 870
rect 3940 790 3950 870
rect 3850 780 3950 790
rect 4050 870 4150 880
rect 4050 790 4060 870
rect 4140 790 4150 870
rect 4050 780 4150 790
rect 4250 870 4350 880
rect 4250 790 4260 870
rect 4340 790 4350 870
rect 4250 780 4350 790
rect 4450 870 4550 880
rect 4450 790 4460 870
rect 4540 790 4550 870
rect 4450 780 4550 790
rect 4650 870 4750 880
rect 4650 790 4660 870
rect 4740 790 4750 870
rect 4650 780 4750 790
rect 4850 870 4950 880
rect 4850 790 4860 870
rect 4940 790 4950 870
rect 4850 780 4950 790
rect 5050 870 5150 880
rect 5050 790 5060 870
rect 5140 790 5150 870
rect 5050 780 5150 790
rect 5250 870 5350 880
rect 5250 790 5260 870
rect 5340 790 5350 870
rect 5250 780 5350 790
rect 5450 870 5550 880
rect 5450 790 5460 870
rect 5540 790 5550 870
rect 5450 780 5550 790
rect 5650 870 5750 880
rect 5650 790 5660 870
rect 5740 790 5750 870
rect 5650 780 5750 790
rect 5850 870 5950 880
rect 5850 790 5860 870
rect 5940 790 5950 870
rect 5850 780 5950 790
rect 6050 870 6150 880
rect 6050 790 6060 870
rect 6140 790 6150 870
rect 6050 780 6150 790
rect 6250 870 6350 880
rect 6250 790 6260 870
rect 6340 790 6350 870
rect 6250 780 6350 790
rect 6450 870 6550 880
rect 6450 790 6460 870
rect 6540 790 6550 870
rect 6450 780 6550 790
rect -115 695 -85 780
rect 85 695 115 780
rect 285 695 315 780
rect 485 695 515 780
rect 685 695 715 780
rect 885 695 915 780
rect 1085 695 1115 780
rect 1285 695 1315 780
rect 1485 695 1515 780
rect 1685 695 1715 780
rect 1885 695 1915 780
rect 2085 695 2115 780
rect 2285 695 2315 780
rect 2485 695 2515 780
rect 2685 695 2715 780
rect 2885 695 2915 780
rect 3085 695 3115 780
rect 3285 695 3315 780
rect 3485 695 3515 780
rect 3685 695 3715 780
rect 3885 695 3915 780
rect 4085 695 4115 780
rect 4285 695 4315 780
rect 4485 695 4515 780
rect 4685 695 4715 780
rect 4885 695 4915 780
rect 5085 695 5115 780
rect 5285 695 5315 780
rect 5485 695 5515 780
rect 5685 695 5715 780
rect 5885 695 5915 780
rect 6085 695 6115 780
rect 6285 695 6315 780
rect 6485 695 6515 780
rect -150 685 -50 695
rect -150 605 -140 685
rect -60 605 -50 685
rect -150 595 -50 605
rect 50 685 150 695
rect 50 605 60 685
rect 140 605 150 685
rect 50 595 150 605
rect 250 685 350 695
rect 250 605 260 685
rect 340 605 350 685
rect 250 595 350 605
rect 450 685 550 695
rect 450 605 460 685
rect 540 605 550 685
rect 450 595 550 605
rect 650 685 750 695
rect 650 605 660 685
rect 740 605 750 685
rect 650 595 750 605
rect 850 685 950 695
rect 850 605 860 685
rect 940 605 950 685
rect 850 595 950 605
rect 1050 685 1150 695
rect 1050 605 1060 685
rect 1140 605 1150 685
rect 1050 595 1150 605
rect 1250 685 1350 695
rect 1250 605 1260 685
rect 1340 605 1350 685
rect 1250 595 1350 605
rect 1450 685 1550 695
rect 1450 605 1460 685
rect 1540 605 1550 685
rect 1450 595 1550 605
rect 1650 685 1750 695
rect 1650 605 1660 685
rect 1740 605 1750 685
rect 1650 595 1750 605
rect 1850 685 1950 695
rect 1850 605 1860 685
rect 1940 605 1950 685
rect 1850 595 1950 605
rect 2050 685 2150 695
rect 2050 605 2060 685
rect 2140 605 2150 685
rect 2050 595 2150 605
rect 2250 685 2350 695
rect 2250 605 2260 685
rect 2340 605 2350 685
rect 2250 595 2350 605
rect 2450 685 2550 695
rect 2450 605 2460 685
rect 2540 605 2550 685
rect 2450 595 2550 605
rect 2650 685 2750 695
rect 2650 605 2660 685
rect 2740 605 2750 685
rect 2650 595 2750 605
rect 2850 685 2950 695
rect 2850 605 2860 685
rect 2940 605 2950 685
rect 2850 595 2950 605
rect 3050 685 3150 695
rect 3050 605 3060 685
rect 3140 605 3150 685
rect 3050 595 3150 605
rect 3250 685 3350 695
rect 3250 605 3260 685
rect 3340 605 3350 685
rect 3250 595 3350 605
rect 3450 685 3550 695
rect 3450 605 3460 685
rect 3540 605 3550 685
rect 3450 595 3550 605
rect 3650 685 3750 695
rect 3650 605 3660 685
rect 3740 605 3750 685
rect 3650 595 3750 605
rect 3850 685 3950 695
rect 3850 605 3860 685
rect 3940 605 3950 685
rect 3850 595 3950 605
rect 4050 685 4150 695
rect 4050 605 4060 685
rect 4140 605 4150 685
rect 4050 595 4150 605
rect 4250 685 4350 695
rect 4250 605 4260 685
rect 4340 605 4350 685
rect 4250 595 4350 605
rect 4450 685 4550 695
rect 4450 605 4460 685
rect 4540 605 4550 685
rect 4450 595 4550 605
rect 4650 685 4750 695
rect 4650 605 4660 685
rect 4740 605 4750 685
rect 4650 595 4750 605
rect 4850 685 4950 695
rect 4850 605 4860 685
rect 4940 605 4950 685
rect 4850 595 4950 605
rect 5050 685 5150 695
rect 5050 605 5060 685
rect 5140 605 5150 685
rect 5050 595 5150 605
rect 5250 685 5350 695
rect 5250 605 5260 685
rect 5340 605 5350 685
rect 5250 595 5350 605
rect 5450 685 5550 695
rect 5450 605 5460 685
rect 5540 605 5550 685
rect 5450 595 5550 605
rect 5650 685 5750 695
rect 5650 605 5660 685
rect 5740 605 5750 685
rect 5650 595 5750 605
rect 5850 685 5950 695
rect 5850 605 5860 685
rect 5940 605 5950 685
rect 5850 595 5950 605
rect 6050 685 6150 695
rect 6050 605 6060 685
rect 6140 605 6150 685
rect 6050 595 6150 605
rect 6250 685 6350 695
rect 6250 605 6260 685
rect 6340 605 6350 685
rect 6250 595 6350 605
rect 6450 685 6550 695
rect 6450 605 6460 685
rect 6540 605 6550 685
rect 6450 595 6550 605
rect -115 510 -85 595
rect 85 510 115 595
rect 285 510 315 595
rect 485 510 515 595
rect 685 510 715 595
rect 885 510 915 595
rect 1085 510 1115 595
rect 1285 510 1315 595
rect 1485 510 1515 595
rect 1685 510 1715 595
rect 1885 510 1915 595
rect 2085 510 2115 595
rect 2285 510 2315 595
rect 2485 510 2515 595
rect 2685 510 2715 595
rect 2885 510 2915 595
rect 3085 510 3115 595
rect 3285 510 3315 595
rect 3485 510 3515 595
rect 3685 510 3715 595
rect 3885 510 3915 595
rect 4085 510 4115 595
rect 4285 510 4315 595
rect 4485 510 4515 595
rect 4685 510 4715 595
rect 4885 510 4915 595
rect 5085 510 5115 595
rect 5285 510 5315 595
rect 5485 510 5515 595
rect 5685 510 5715 595
rect 5885 510 5915 595
rect 6085 510 6115 595
rect 6285 510 6315 595
rect 6485 510 6515 595
rect -150 500 -50 510
rect -150 420 -140 500
rect -60 420 -50 500
rect -150 410 -50 420
rect 50 500 150 510
rect 50 420 60 500
rect 140 420 150 500
rect 50 410 150 420
rect 250 500 350 510
rect 250 420 260 500
rect 340 420 350 500
rect 250 410 350 420
rect 450 500 550 510
rect 450 420 460 500
rect 540 420 550 500
rect 450 410 550 420
rect 650 500 750 510
rect 650 420 660 500
rect 740 420 750 500
rect 650 410 750 420
rect 850 500 950 510
rect 850 420 860 500
rect 940 420 950 500
rect 850 410 950 420
rect 1050 500 1150 510
rect 1050 420 1060 500
rect 1140 420 1150 500
rect 1050 410 1150 420
rect 1250 500 1350 510
rect 1250 420 1260 500
rect 1340 420 1350 500
rect 1250 410 1350 420
rect 1450 500 1550 510
rect 1450 420 1460 500
rect 1540 420 1550 500
rect 1450 410 1550 420
rect 1650 500 1750 510
rect 1650 420 1660 500
rect 1740 420 1750 500
rect 1650 410 1750 420
rect 1850 500 1950 510
rect 1850 420 1860 500
rect 1940 420 1950 500
rect 1850 410 1950 420
rect 2050 500 2150 510
rect 2050 420 2060 500
rect 2140 420 2150 500
rect 2050 410 2150 420
rect 2250 500 2350 510
rect 2250 420 2260 500
rect 2340 420 2350 500
rect 2250 410 2350 420
rect 2450 500 2550 510
rect 2450 420 2460 500
rect 2540 420 2550 500
rect 2450 410 2550 420
rect 2650 500 2750 510
rect 2650 420 2660 500
rect 2740 420 2750 500
rect 2650 410 2750 420
rect 2850 500 2950 510
rect 2850 420 2860 500
rect 2940 420 2950 500
rect 2850 410 2950 420
rect 3050 500 3150 510
rect 3050 420 3060 500
rect 3140 420 3150 500
rect 3050 410 3150 420
rect 3250 500 3350 510
rect 3250 420 3260 500
rect 3340 420 3350 500
rect 3250 410 3350 420
rect 3450 500 3550 510
rect 3450 420 3460 500
rect 3540 420 3550 500
rect 3450 410 3550 420
rect 3650 500 3750 510
rect 3650 420 3660 500
rect 3740 420 3750 500
rect 3650 410 3750 420
rect 3850 500 3950 510
rect 3850 420 3860 500
rect 3940 420 3950 500
rect 3850 410 3950 420
rect 4050 500 4150 510
rect 4050 420 4060 500
rect 4140 420 4150 500
rect 4050 410 4150 420
rect 4250 500 4350 510
rect 4250 420 4260 500
rect 4340 420 4350 500
rect 4250 410 4350 420
rect 4450 500 4550 510
rect 4450 420 4460 500
rect 4540 420 4550 500
rect 4450 410 4550 420
rect 4650 500 4750 510
rect 4650 420 4660 500
rect 4740 420 4750 500
rect 4650 410 4750 420
rect 4850 500 4950 510
rect 4850 420 4860 500
rect 4940 420 4950 500
rect 4850 410 4950 420
rect 5050 500 5150 510
rect 5050 420 5060 500
rect 5140 420 5150 500
rect 5050 410 5150 420
rect 5250 500 5350 510
rect 5250 420 5260 500
rect 5340 420 5350 500
rect 5250 410 5350 420
rect 5450 500 5550 510
rect 5450 420 5460 500
rect 5540 420 5550 500
rect 5450 410 5550 420
rect 5650 500 5750 510
rect 5650 420 5660 500
rect 5740 420 5750 500
rect 5650 410 5750 420
rect 5850 500 5950 510
rect 5850 420 5860 500
rect 5940 420 5950 500
rect 5850 410 5950 420
rect 6050 500 6150 510
rect 6050 420 6060 500
rect 6140 420 6150 500
rect 6050 410 6150 420
rect 6250 500 6350 510
rect 6250 420 6260 500
rect 6340 420 6350 500
rect 6250 410 6350 420
rect 6450 500 6550 510
rect 6450 420 6460 500
rect 6540 420 6550 500
rect 6450 410 6550 420
rect -115 325 -85 410
rect 85 325 115 410
rect 285 325 315 410
rect 485 325 515 410
rect 685 325 715 410
rect 885 325 915 410
rect 1085 325 1115 410
rect 1285 325 1315 410
rect 1485 325 1515 410
rect 1685 325 1715 410
rect 1885 325 1915 410
rect 2085 325 2115 410
rect 2285 325 2315 410
rect 2485 325 2515 410
rect 2685 325 2715 410
rect 2885 325 2915 410
rect 3085 325 3115 410
rect 3285 325 3315 410
rect 3485 325 3515 410
rect 3685 325 3715 410
rect 3885 325 3915 410
rect 4085 325 4115 410
rect 4285 325 4315 410
rect 4485 325 4515 410
rect 4685 325 4715 410
rect 4885 325 4915 410
rect 5085 325 5115 410
rect 5285 325 5315 410
rect 5485 325 5515 410
rect 5685 325 5715 410
rect 5885 325 5915 410
rect 6085 325 6115 410
rect 6285 325 6315 410
rect 6485 325 6515 410
rect -150 315 -50 325
rect -150 235 -140 315
rect -60 235 -50 315
rect -150 225 -50 235
rect 50 315 150 325
rect 50 235 60 315
rect 140 235 150 315
rect 50 225 150 235
rect 250 315 350 325
rect 250 235 260 315
rect 340 235 350 315
rect 250 225 350 235
rect 450 315 550 325
rect 450 235 460 315
rect 540 235 550 315
rect 450 225 550 235
rect 650 315 750 325
rect 650 235 660 315
rect 740 235 750 315
rect 650 225 750 235
rect 850 315 950 325
rect 850 235 860 315
rect 940 235 950 315
rect 850 225 950 235
rect 1050 315 1150 325
rect 1050 235 1060 315
rect 1140 235 1150 315
rect 1050 225 1150 235
rect 1250 315 1350 325
rect 1250 235 1260 315
rect 1340 235 1350 315
rect 1250 225 1350 235
rect 1450 315 1550 325
rect 1450 235 1460 315
rect 1540 235 1550 315
rect 1450 225 1550 235
rect 1650 315 1750 325
rect 1650 235 1660 315
rect 1740 235 1750 315
rect 1650 225 1750 235
rect 1850 315 1950 325
rect 1850 235 1860 315
rect 1940 235 1950 315
rect 1850 225 1950 235
rect 2050 315 2150 325
rect 2050 235 2060 315
rect 2140 235 2150 315
rect 2050 225 2150 235
rect 2250 315 2350 325
rect 2250 235 2260 315
rect 2340 235 2350 315
rect 2250 225 2350 235
rect 2450 315 2550 325
rect 2450 235 2460 315
rect 2540 235 2550 315
rect 2450 225 2550 235
rect 2650 315 2750 325
rect 2650 235 2660 315
rect 2740 235 2750 315
rect 2650 225 2750 235
rect 2850 315 2950 325
rect 2850 235 2860 315
rect 2940 235 2950 315
rect 2850 225 2950 235
rect 3050 315 3150 325
rect 3050 235 3060 315
rect 3140 235 3150 315
rect 3050 225 3150 235
rect 3250 315 3350 325
rect 3250 235 3260 315
rect 3340 235 3350 315
rect 3250 225 3350 235
rect 3450 315 3550 325
rect 3450 235 3460 315
rect 3540 235 3550 315
rect 3450 225 3550 235
rect 3650 315 3750 325
rect 3650 235 3660 315
rect 3740 235 3750 315
rect 3650 225 3750 235
rect 3850 315 3950 325
rect 3850 235 3860 315
rect 3940 235 3950 315
rect 3850 225 3950 235
rect 4050 315 4150 325
rect 4050 235 4060 315
rect 4140 235 4150 315
rect 4050 225 4150 235
rect 4250 315 4350 325
rect 4250 235 4260 315
rect 4340 235 4350 315
rect 4250 225 4350 235
rect 4450 315 4550 325
rect 4450 235 4460 315
rect 4540 235 4550 315
rect 4450 225 4550 235
rect 4650 315 4750 325
rect 4650 235 4660 315
rect 4740 235 4750 315
rect 4650 225 4750 235
rect 4850 315 4950 325
rect 4850 235 4860 315
rect 4940 235 4950 315
rect 4850 225 4950 235
rect 5050 315 5150 325
rect 5050 235 5060 315
rect 5140 235 5150 315
rect 5050 225 5150 235
rect 5250 315 5350 325
rect 5250 235 5260 315
rect 5340 235 5350 315
rect 5250 225 5350 235
rect 5450 315 5550 325
rect 5450 235 5460 315
rect 5540 235 5550 315
rect 5450 225 5550 235
rect 5650 315 5750 325
rect 5650 235 5660 315
rect 5740 235 5750 315
rect 5650 225 5750 235
rect 5850 315 5950 325
rect 5850 235 5860 315
rect 5940 235 5950 315
rect 5850 225 5950 235
rect 6050 315 6150 325
rect 6050 235 6060 315
rect 6140 235 6150 315
rect 6050 225 6150 235
rect 6250 315 6350 325
rect 6250 235 6260 315
rect 6340 235 6350 315
rect 6250 225 6350 235
rect 6450 315 6550 325
rect 6450 235 6460 315
rect 6540 235 6550 315
rect 6450 225 6550 235
rect -115 140 -85 225
rect 85 140 115 225
rect 285 140 315 225
rect 485 140 515 225
rect 685 140 715 225
rect 885 140 915 225
rect 1085 140 1115 225
rect 1285 140 1315 225
rect 1485 140 1515 225
rect 1685 140 1715 225
rect 1885 140 1915 225
rect 2085 140 2115 225
rect 2285 140 2315 225
rect 2485 140 2515 225
rect 2685 140 2715 225
rect 2885 140 2915 225
rect 3085 140 3115 225
rect 3285 140 3315 225
rect 3485 140 3515 225
rect 3685 140 3715 225
rect 3885 140 3915 225
rect 4085 140 4115 225
rect 4285 140 4315 225
rect 4485 140 4515 225
rect 4685 140 4715 225
rect 4885 140 4915 225
rect 5085 140 5115 225
rect 5285 140 5315 225
rect 5485 140 5515 225
rect 5685 140 5715 225
rect 5885 140 5915 225
rect 6085 140 6115 225
rect 6285 140 6315 225
rect 6485 140 6515 225
rect -150 130 -50 140
rect -150 50 -140 130
rect -60 50 -50 130
rect -150 40 -50 50
rect 50 130 150 140
rect 50 50 60 130
rect 140 50 150 130
rect 50 40 150 50
rect 250 130 350 140
rect 250 50 260 130
rect 340 50 350 130
rect 250 40 350 50
rect 450 130 550 140
rect 450 50 460 130
rect 540 50 550 130
rect 450 40 550 50
rect 650 130 750 140
rect 650 50 660 130
rect 740 50 750 130
rect 650 40 750 50
rect 850 130 950 140
rect 850 50 860 130
rect 940 50 950 130
rect 850 40 950 50
rect 1050 130 1150 140
rect 1050 50 1060 130
rect 1140 50 1150 130
rect 1050 40 1150 50
rect 1250 130 1350 140
rect 1250 50 1260 130
rect 1340 50 1350 130
rect 1250 40 1350 50
rect 1450 130 1550 140
rect 1450 50 1460 130
rect 1540 50 1550 130
rect 1450 40 1550 50
rect 1650 130 1750 140
rect 1650 50 1660 130
rect 1740 50 1750 130
rect 1650 40 1750 50
rect 1850 130 1950 140
rect 1850 50 1860 130
rect 1940 50 1950 130
rect 1850 40 1950 50
rect 2050 130 2150 140
rect 2050 50 2060 130
rect 2140 50 2150 130
rect 2050 40 2150 50
rect 2250 130 2350 140
rect 2250 50 2260 130
rect 2340 50 2350 130
rect 2250 40 2350 50
rect 2450 130 2550 140
rect 2450 50 2460 130
rect 2540 50 2550 130
rect 2450 40 2550 50
rect 2650 130 2750 140
rect 2650 50 2660 130
rect 2740 50 2750 130
rect 2650 40 2750 50
rect 2850 130 2950 140
rect 2850 50 2860 130
rect 2940 50 2950 130
rect 2850 40 2950 50
rect 3050 130 3150 140
rect 3050 50 3060 130
rect 3140 50 3150 130
rect 3050 40 3150 50
rect 3250 130 3350 140
rect 3250 50 3260 130
rect 3340 50 3350 130
rect 3250 40 3350 50
rect 3450 130 3550 140
rect 3450 50 3460 130
rect 3540 50 3550 130
rect 3450 40 3550 50
rect 3650 130 3750 140
rect 3650 50 3660 130
rect 3740 50 3750 130
rect 3650 40 3750 50
rect 3850 130 3950 140
rect 3850 50 3860 130
rect 3940 50 3950 130
rect 3850 40 3950 50
rect 4050 130 4150 140
rect 4050 50 4060 130
rect 4140 50 4150 130
rect 4050 40 4150 50
rect 4250 130 4350 140
rect 4250 50 4260 130
rect 4340 50 4350 130
rect 4250 40 4350 50
rect 4450 130 4550 140
rect 4450 50 4460 130
rect 4540 50 4550 130
rect 4450 40 4550 50
rect 4650 130 4750 140
rect 4650 50 4660 130
rect 4740 50 4750 130
rect 4650 40 4750 50
rect 4850 130 4950 140
rect 4850 50 4860 130
rect 4940 50 4950 130
rect 4850 40 4950 50
rect 5050 130 5150 140
rect 5050 50 5060 130
rect 5140 50 5150 130
rect 5050 40 5150 50
rect 5250 130 5350 140
rect 5250 50 5260 130
rect 5340 50 5350 130
rect 5250 40 5350 50
rect 5450 130 5550 140
rect 5450 50 5460 130
rect 5540 50 5550 130
rect 5450 40 5550 50
rect 5650 130 5750 140
rect 5650 50 5660 130
rect 5740 50 5750 130
rect 5650 40 5750 50
rect 5850 130 5950 140
rect 5850 50 5860 130
rect 5940 50 5950 130
rect 5850 40 5950 50
rect 6050 130 6150 140
rect 6050 50 6060 130
rect 6140 50 6150 130
rect 6050 40 6150 50
rect 6250 130 6350 140
rect 6250 50 6260 130
rect 6340 50 6350 130
rect 6250 40 6350 50
rect 6450 130 6550 140
rect 6450 50 6460 130
rect 6540 50 6550 130
rect 6450 40 6550 50
rect -115 -45 -85 40
rect 85 -45 115 40
rect 285 -45 315 40
rect 485 -45 515 40
rect 685 -45 715 40
rect 885 -45 915 40
rect 1085 -45 1115 40
rect 1285 -45 1315 40
rect 1485 -45 1515 40
rect 1685 -45 1715 40
rect 1885 -45 1915 40
rect 2085 -45 2115 40
rect 2285 -45 2315 40
rect 2485 -45 2515 40
rect 2685 -45 2715 40
rect 2885 -45 2915 40
rect 3085 -45 3115 40
rect 3285 -45 3315 40
rect 3485 -45 3515 40
rect 3685 -45 3715 40
rect 3885 -45 3915 40
rect 4085 -45 4115 40
rect 4285 -45 4315 40
rect 4485 -45 4515 40
rect 4685 -45 4715 40
rect 4885 -45 4915 40
rect 5085 -45 5115 40
rect 5285 -45 5315 40
rect 5485 -45 5515 40
rect 5685 -45 5715 40
rect 5885 -45 5915 40
rect 6085 -45 6115 40
rect 6285 -45 6315 40
rect 6485 -45 6515 40
rect -150 -55 -50 -45
rect -150 -135 -140 -55
rect -60 -135 -50 -55
rect -150 -145 -50 -135
rect 50 -55 150 -45
rect 50 -135 60 -55
rect 140 -80 150 -55
rect 250 -55 350 -45
rect 250 -80 260 -55
rect 140 -110 260 -80
rect 140 -135 150 -110
rect 50 -145 150 -135
rect 250 -135 260 -110
rect 340 -80 350 -55
rect 450 -55 550 -45
rect 450 -80 460 -55
rect 340 -110 460 -80
rect 340 -135 350 -110
rect 250 -145 350 -135
rect 450 -135 460 -110
rect 540 -80 550 -55
rect 650 -55 750 -45
rect 650 -80 660 -55
rect 540 -110 660 -80
rect 540 -135 550 -110
rect 450 -145 550 -135
rect 650 -135 660 -110
rect 740 -80 750 -55
rect 850 -55 950 -45
rect 850 -80 860 -55
rect 740 -110 860 -80
rect 740 -135 750 -110
rect 650 -145 750 -135
rect 850 -135 860 -110
rect 940 -80 950 -55
rect 1050 -55 1150 -45
rect 1050 -80 1060 -55
rect 940 -110 1060 -80
rect 940 -135 950 -110
rect 850 -145 950 -135
rect 1050 -135 1060 -110
rect 1140 -80 1150 -55
rect 1250 -55 1350 -45
rect 1250 -80 1260 -55
rect 1140 -110 1260 -80
rect 1140 -135 1150 -110
rect 1050 -145 1150 -135
rect 1250 -135 1260 -110
rect 1340 -80 1350 -55
rect 1450 -55 1550 -45
rect 1450 -80 1460 -55
rect 1340 -110 1460 -80
rect 1340 -135 1350 -110
rect 1250 -145 1350 -135
rect 1450 -135 1460 -110
rect 1540 -80 1550 -55
rect 1650 -55 1750 -45
rect 1650 -80 1660 -55
rect 1540 -110 1660 -80
rect 1540 -135 1550 -110
rect 1450 -145 1550 -135
rect 1650 -135 1660 -110
rect 1740 -80 1750 -55
rect 1850 -55 1950 -45
rect 1850 -80 1860 -55
rect 1740 -110 1860 -80
rect 1740 -135 1750 -110
rect 1650 -145 1750 -135
rect 1850 -135 1860 -110
rect 1940 -80 1950 -55
rect 2050 -55 2150 -45
rect 2050 -80 2060 -55
rect 1940 -110 2060 -80
rect 1940 -135 1950 -110
rect 1850 -145 1950 -135
rect 2050 -135 2060 -110
rect 2140 -80 2150 -55
rect 2250 -55 2350 -45
rect 2250 -80 2260 -55
rect 2140 -110 2260 -80
rect 2140 -135 2150 -110
rect 2050 -145 2150 -135
rect 2250 -135 2260 -110
rect 2340 -80 2350 -55
rect 2450 -55 2550 -45
rect 2450 -80 2460 -55
rect 2340 -110 2460 -80
rect 2340 -135 2350 -110
rect 2250 -145 2350 -135
rect 2450 -135 2460 -110
rect 2540 -80 2550 -55
rect 2650 -55 2750 -45
rect 2650 -80 2660 -55
rect 2540 -110 2660 -80
rect 2540 -135 2550 -110
rect 2450 -145 2550 -135
rect 2650 -135 2660 -110
rect 2740 -80 2750 -55
rect 2850 -55 2950 -45
rect 2850 -80 2860 -55
rect 2740 -110 2860 -80
rect 2740 -135 2750 -110
rect 2650 -145 2750 -135
rect 2850 -135 2860 -110
rect 2940 -80 2950 -55
rect 3050 -55 3150 -45
rect 3050 -80 3060 -55
rect 2940 -110 3060 -80
rect 2940 -135 2950 -110
rect 2850 -145 2950 -135
rect 3050 -135 3060 -110
rect 3140 -80 3150 -55
rect 3250 -55 3350 -45
rect 3250 -80 3260 -55
rect 3140 -110 3260 -80
rect 3140 -135 3150 -110
rect 3050 -145 3150 -135
rect 3250 -135 3260 -110
rect 3340 -80 3350 -55
rect 3450 -55 3550 -45
rect 3450 -80 3460 -55
rect 3340 -110 3460 -80
rect 3340 -135 3350 -110
rect 3250 -145 3350 -135
rect 3450 -135 3460 -110
rect 3540 -80 3550 -55
rect 3650 -55 3750 -45
rect 3650 -80 3660 -55
rect 3540 -110 3660 -80
rect 3540 -135 3550 -110
rect 3450 -145 3550 -135
rect 3650 -135 3660 -110
rect 3740 -80 3750 -55
rect 3850 -55 3950 -45
rect 3850 -80 3860 -55
rect 3740 -110 3860 -80
rect 3740 -135 3750 -110
rect 3650 -145 3750 -135
rect 3850 -135 3860 -110
rect 3940 -80 3950 -55
rect 4050 -55 4150 -45
rect 4050 -80 4060 -55
rect 3940 -110 4060 -80
rect 3940 -135 3950 -110
rect 3850 -145 3950 -135
rect 4050 -135 4060 -110
rect 4140 -80 4150 -55
rect 4250 -55 4350 -45
rect 4250 -80 4260 -55
rect 4140 -110 4260 -80
rect 4140 -135 4150 -110
rect 4050 -145 4150 -135
rect 4250 -135 4260 -110
rect 4340 -80 4350 -55
rect 4450 -55 4550 -45
rect 4450 -80 4460 -55
rect 4340 -110 4460 -80
rect 4340 -135 4350 -110
rect 4250 -145 4350 -135
rect 4450 -135 4460 -110
rect 4540 -80 4550 -55
rect 4650 -55 4750 -45
rect 4650 -80 4660 -55
rect 4540 -110 4660 -80
rect 4540 -135 4550 -110
rect 4450 -145 4550 -135
rect 4650 -135 4660 -110
rect 4740 -80 4750 -55
rect 4850 -55 4950 -45
rect 4850 -80 4860 -55
rect 4740 -110 4860 -80
rect 4740 -135 4750 -110
rect 4650 -145 4750 -135
rect 4850 -135 4860 -110
rect 4940 -80 4950 -55
rect 5050 -55 5150 -45
rect 5050 -80 5060 -55
rect 4940 -110 5060 -80
rect 4940 -135 4950 -110
rect 4850 -145 4950 -135
rect 5050 -135 5060 -110
rect 5140 -80 5150 -55
rect 5250 -55 5350 -45
rect 5250 -80 5260 -55
rect 5140 -110 5260 -80
rect 5140 -135 5150 -110
rect 5050 -145 5150 -135
rect 5250 -135 5260 -110
rect 5340 -80 5350 -55
rect 5450 -55 5550 -45
rect 5450 -80 5460 -55
rect 5340 -110 5460 -80
rect 5340 -135 5350 -110
rect 5250 -145 5350 -135
rect 5450 -135 5460 -110
rect 5540 -80 5550 -55
rect 5650 -55 5750 -45
rect 5650 -80 5660 -55
rect 5540 -110 5660 -80
rect 5540 -135 5550 -110
rect 5450 -145 5550 -135
rect 5650 -135 5660 -110
rect 5740 -80 5750 -55
rect 5850 -55 5950 -45
rect 5850 -80 5860 -55
rect 5740 -110 5860 -80
rect 5740 -135 5750 -110
rect 5650 -145 5750 -135
rect 5850 -135 5860 -110
rect 5940 -80 5950 -55
rect 6050 -55 6150 -45
rect 6050 -80 6060 -55
rect 5940 -110 6060 -80
rect 5940 -135 5950 -110
rect 5850 -145 5950 -135
rect 6050 -135 6060 -110
rect 6140 -80 6150 -55
rect 6250 -55 6350 -45
rect 6250 -80 6260 -55
rect 6140 -110 6260 -80
rect 6140 -135 6150 -110
rect 6050 -145 6150 -135
rect 6250 -135 6260 -110
rect 6340 -135 6350 -55
rect 6250 -145 6350 -135
rect 6450 -55 6550 -45
rect 6450 -135 6460 -55
rect 6540 -135 6550 -55
rect 6450 -145 6550 -135
rect -115 -185 -85 -145
rect 85 -185 115 -145
rect 285 -185 315 -145
rect 485 -185 515 -145
rect 685 -185 715 -145
rect 885 -185 915 -145
rect 1085 -185 1115 -145
rect 1285 -185 1315 -145
rect 1485 -185 1515 -145
rect 1685 -185 1715 -145
rect 1885 -185 1915 -145
rect 2085 -185 2115 -145
rect 2285 -185 2315 -145
rect 2485 -185 2515 -145
rect 2685 -185 2715 -145
rect 2885 -185 2915 -145
rect 3085 -185 3115 -145
rect 3285 -185 3315 -145
rect 3485 -185 3515 -145
rect 3685 -185 3715 -145
rect 3885 -185 3915 -145
rect 4085 -185 4115 -145
rect 4285 -185 4315 -145
rect 4485 -185 4515 -145
rect 4685 -185 4715 -145
rect 4885 -185 4915 -145
rect 5085 -185 5115 -145
rect 5285 -185 5315 -145
rect 5485 -185 5515 -145
rect 5685 -185 5715 -145
rect 5885 -185 5915 -145
rect 6085 -185 6115 -145
rect 6285 -185 6315 -145
rect 6485 -185 6515 -145
<< labels >>
rlabel metal1 6680 1935 6690 1945 1 C10
port 12 n
rlabel metal4 6295 12060 6305 12070 1 Ctop
port 14 n
rlabel metal4 6495 12055 6505 12065 1 VSS
port 15 n
rlabel metal1 6680 3045 6690 3055 1 C9
port 11 n
rlabel metal1 6680 3970 6690 3980 1 C8
port 10 n
rlabel metal1 6680 4525 6690 4535 1 C7
port 9 n
rlabel metal1 6680 4895 6690 4905 1 C6
port 8 n
rlabel metal1 6680 5080 6690 5090 1 C5
port 7 n
rlabel metal1 6680 5450 6690 5460 1 C4
port 6 n
rlabel metal1 6680 6375 6690 6385 1 C3
port 5 n
rlabel metal1 6680 5635 6690 5645 1 C2
port 4 n
rlabel metal1 6680 6190 6690 6200 1 C1
port 3 n
rlabel metal1 6680 6005 6690 6015 1 C0
port 2 n
rlabel metal1 6680 5820 6690 5830 1 C0_dummy
port 1 n
<< end >>
