* SPICE3 file created from preamplifier_flat.ext - technology: sky130A

.subckt preamplifier IN_N IN_P VDD EN OUT_P OUT_N VSS CAL_P CAL_N
X0 a_468_8407# IN_P a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1 a_468_8407# IN_P a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X2 a_468_6971# IN_N a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X3 a_n2304_8007# IN_P a_468_8407# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4 a_n1438_7546# a_n400_8007# OUT_P VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X5 a_2588_6962# a_6950_9426# VSS sky130_fd_pr__res_high_po_0p35 l=18
X6 a_n2304_8007# a_n3220_7910# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X7 a_n2848_8007# CAL_P a_n1954_7546# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X8 a_n624_7154# a_n882_7066# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X9 a_468_6971# IN_N a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X10 a_n2304_8007# IN_N a_468_6971# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X11 a_468_6971# IN_N a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X12 a_n2304_8007# IN_P a_468_8407# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X13 a_n1954_7546# a_n400_8007# OUT_N VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X14 VDD EN a_n3220_7910# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X15 OUT_N VSS a_468_8407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X16 a_n2848_8007# a_n3220_7910# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X17 OUT_P VSS a_468_6971# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X18 a_2588_6962# EN VSS VSS sky130_fd_pr__nfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.15
X19 a_468_8407# IN_P a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X20 a_n2304_8007# IN_N a_468_6971# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X21 a_n2304_8007# a_n3220_7910# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X22 VSS a_n882_7066# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=8.924 ps=66.62 w=2 l=0.15
X23 a_n3220_7910# a_6950_9426# VSS sky130_fd_pr__res_high_po_0p35 l=18
X24 a_2950_8762# a_6950_8928# VSS sky130_fd_pr__res_high_po_0p35 l=18
X25 OUT_P a_n400_8007# a_n1438_7546# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X26 a_n2304_8007# IN_P a_468_8407# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X27 a_n2304_8007# IN_N a_468_6971# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X28 a_468_8407# IN_P a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X29 a_n2304_8007# a_n3220_7910# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X30 VSS a_n882_7066# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X31 a_n3230_7261# EN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X32 a_468_6971# IN_N a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X33 VDD OUT_P a_n624_7154# VSS sky130_fd_pr__nfet_03v3_nvt ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X34 a_468_8407# VSS OUT_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X35 a_n1438_7546# a_n400_8007# OUT_P VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X36 a_n2304_8007# a_n3220_7910# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X37 a_n2304_8007# IN_N a_468_6971# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X38 a_n1954_7546# VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.589 ps=4.42 w=1.9 l=0.15
X39 a_2950_9094# OUT_P VSS sky130_fd_pr__res_high_po_0p35 l=18
X40 a_n1954_7546# a_n400_8007# OUT_N VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X41 a_468_8407# IN_P a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X42 VSS VSS a_n1438_7546# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.589 pd=4.42 as=0.3135 ps=2.23 w=1.9 l=0.15
X43 a_n400_8007# a_n3220_7910# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X44 a_2950_9094# a_6950_8928# VSS sky130_fd_pr__res_high_po_0p35 l=18
X45 a_n2304_8007# IN_P a_468_8407# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X46 a_468_6971# IN_N a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X47 a_n2848_8007# a_n3220_7910# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X48 a_468_6971# IN_N a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X49 a_n2304_8007# IN_P a_468_8407# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X50 a_n624_7154# OUT_N VDD VSS sky130_fd_pr__nfet_03v3_nvt ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X51 OUT_N VSS a_468_8407# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X52 a_n2304_8007# a_n3220_7910# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X53 a_2950_8762# a_6950_8596# VSS sky130_fd_pr__res_high_po_0p35 l=18
X54 OUT_N a_n400_8007# a_n1954_7546# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X55 a_n2304_8007# IN_N a_468_6971# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X56 a_n400_8007# a_n3230_7261# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X57 a_468_6971# VSS OUT_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X58 a_n3220_7910# a_n3220_7910# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X59 a_n624_7154# a_n882_7066# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X60 a_2950_8430# a_6950_8596# VSS sky130_fd_pr__res_high_po_0p35 l=18
X61 a_n1438_7546# a_n624_7154# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X62 a_468_8407# VSS OUT_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X63 a_468_8407# IN_P a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X64 a_468_6971# IN_N a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X65 a_n2304_8007# IN_N a_468_6971# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X66 a_n2304_8007# IN_P a_468_8407# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X67 a_n2304_8007# a_n3220_7910# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X68 a_468_8407# IN_P a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X69 a_n2304_8007# IN_P a_468_8407# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X70 a_n2304_8007# IN_N a_468_6971# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X71 a_2950_8430# a_6950_8264# VSS sky130_fd_pr__res_high_po_0p35 l=18
X72 VDD a_n3220_7910# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=35.35 ps=253.8 w=8 l=0.5
X73 a_n2848_8007# a_n3220_7910# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X74 a_n3230_7261# EN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X75 a_2950_8098# a_6950_8264# VSS sky130_fd_pr__res_high_po_0p35 l=18
X76 OUT_P a_n400_8007# a_n1438_7546# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X77 a_n2304_8007# IN_N a_468_6971# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X78 a_468_8407# IN_P a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X79 OUT_P VSS a_468_6971# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X80 a_n1438_7546# CAL_N a_n2848_8007# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X81 a_n882_7066# a_n882_7066# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X82 a_2950_8098# OUT_N VSS sky130_fd_pr__res_high_po_0p35 l=18
X83 VSS a_n624_7154# a_n1954_7546# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X84 OUT_N a_n400_8007# a_n1954_7546# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X85 a_n2304_8007# IN_P a_468_8407# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X86 a_468_6971# IN_N a_n2304_8007# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X87 a_n882_7066# a_n400_8007# VSS sky130_fd_pr__res_high_po_0p35 l=18
X88 a_468_6971# VSS OUT_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X89 VDD a_n3220_7910# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.5
C0 a_6950_8928# OUT_N 0.001054f
C1 a_2950_9094# a_2950_8762# 0.296258f
C2 a_6950_8928# OUT_P 0.308867f
C3 OUT_P OUT_N 3.03087f
C4 a_2588_6962# a_2950_8762# 3.86e-20
C5 a_6950_9426# OUT_N 7.07e-21
C6 a_468_6971# a_2950_8762# 2.64e-19
C7 EN OUT_N 1.24e-19
C8 a_2950_8762# VDD 0.043459f
C9 a_6950_9426# OUT_P 0.296508f
C10 EN OUT_P 0.002395f
C11 CAL_P CAL_N 0.869119f
C12 a_2950_9094# EN 0.030938f
C13 a_2588_6962# OUT_N 0.207118f
C14 IN_P OUT_N 1.02e-19
C15 EN CAL_N 0.031057f
C16 a_468_6971# OUT_N 0.079762f
C17 a_2588_6962# OUT_P 0.001576f
C18 a_2588_6962# a_2950_9094# 0.296522f
C19 EN CAL_P 0.480436f
C20 VDD OUT_N 0.288237f
C21 IN_P OUT_P 2.7e-19
C22 IN_N CAL_N 3.61e-21
C23 a_n624_7154# OUT_N 0.178275f
C24 a_468_6971# OUT_P 2.20213f
C25 IN_N CAL_P 7.22e-21
C26 VDD OUT_P 0.575696f
C27 IN_P CAL_N 3.08e-21
C28 a_2950_9094# VDD 0.196089f
C29 a_n882_7066# OUT_N 0.005657f
C30 a_n624_7154# OUT_P 0.259481f
C31 a_n3230_7261# a_2950_8762# 3.17e-19
C32 VDD CAL_N 0.33878f
C33 IN_P CAL_P 6.16e-21
C34 IN_N EN 0.149397f
C35 a_n624_7154# CAL_N 1.24e-19
C36 a_n1438_7546# OUT_N 0.640491f
C37 a_2588_6962# EN 0.843939f
C38 a_n882_7066# OUT_P 0.008396f
C39 a_468_8407# a_2950_8762# 1.3e-19
C40 IN_P EN 0.151629f
C41 VDD CAL_P 0.343729f
C42 a_n1438_7546# OUT_P 1.92365f
C43 a_n882_7066# CAL_N 3.08e-19
C44 a_n1954_7546# OUT_N 1.5258f
C45 a_n624_7154# CAL_P 0.002915f
C46 a_468_6971# EN 0.051902f
C47 a_2588_6962# IN_N 2.46e-19
C48 a_n400_8007# a_2950_8762# 0.082848f
C49 IN_P IN_N 2.70779f
C50 VDD EN 0.665966f
C51 a_n3230_7261# OUT_N 1.72e-20
C52 a_n1954_7546# OUT_P 1.17133f
C53 a_n1438_7546# CAL_N 0.052373f
C54 a_n882_7066# CAL_P 1.73e-19
C55 a_n624_7154# EN 0.031635f
C56 a_468_6971# IN_N 1.08412f
C57 a_2588_6962# IN_P 8.28e-19
C58 a_n400_8007# a_6950_8928# 7.8e-20
C59 a_468_6971# a_2588_6962# 0.095724f
C60 VDD IN_N 4.45083f
C61 a_2950_8098# OUT_N 1.97e-19
C62 a_468_8407# OUT_N 1.70462f
C63 a_n3230_7261# OUT_P 1.79e-20
C64 a_n1954_7546# CAL_N 0.036205f
C65 a_n1438_7546# CAL_P 0.00316f
C66 a_n882_7066# EN 0.034995f
C67 a_n624_7154# IN_N 0.060805f
C68 a_468_6971# IN_P 0.071587f
C69 a_2588_6962# VDD 0.8341f
C70 a_n3230_7261# a_2950_9094# 1.05e-19
C71 a_n624_7154# a_2588_6962# 0.035115f
C72 a_2950_8098# OUT_P 1.59e-19
C73 VDD IN_P 5.09118f
C74 a_6950_8264# OUT_N 0.301032f
C75 a_n400_8007# OUT_N 0.911395f
C76 a_2950_8762# a_2950_8430# 0.296258f
C77 a_468_8407# OUT_P 0.391059f
C78 a_n1954_7546# CAL_P 0.102027f
C79 a_n1438_7546# EN 0.01719f
C80 a_n882_7066# IN_N 0.100194f
C81 a_n624_7154# IN_P 0.058665f
C82 a_n3230_7261# CAL_N 0.637551f
C83 a_468_6971# VDD 1.04704f
C84 a_n882_7066# a_2588_6962# 0.241119f
C85 a_n624_7154# a_468_6971# 0.13762f
C86 a_6950_8264# OUT_P 0.00191f
C87 a_n624_7154# VDD 0.235486f
C88 a_n2304_8007# OUT_N 4.77e-20
C89 a_n3230_7261# CAL_P 0.035837f
C90 a_n400_8007# OUT_P 0.388914f
C91 a_n1954_7546# EN 1.60318f
C92 a_n1438_7546# IN_N 0.042695f
C93 a_n882_7066# IN_P 0.060633f
C94 a_n400_8007# a_2950_9094# 0.002634f
C95 a_n1438_7546# a_2588_6962# 0.021449f
C96 a_n882_7066# a_468_6971# 0.971846f
C97 a_n882_7066# VDD 0.302129f
C98 a_n3230_7261# EN 0.426226f
C99 a_6950_8928# a_6950_8596# 0.296258f
C100 a_n2304_8007# OUT_P 1.57e-19
C101 a_n1954_7546# IN_N 0.058988f
C102 a_n1438_7546# IN_P 0.034165f
C103 a_n1954_7546# a_2588_6962# 0.030605f
C104 a_n1438_7546# a_468_6971# 2.69237f
C105 a_n882_7066# a_n624_7154# 0.180842f
C106 a_2950_8430# OUT_N 1.16e-19
C107 a_n2304_8007# CAL_N 0.017398f
C108 a_n1438_7546# VDD 0.525635f
C109 a_n3230_7261# IN_N 0.061498f
C110 a_468_8407# EN 0.059771f
C111 a_n1954_7546# IN_P 0.0565f
C112 a_n1954_7546# a_468_6971# 0.574743f
C113 a_n1438_7546# a_n624_7154# 1.95816f
C114 a_n3230_7261# a_2588_6962# 9.77e-19
C115 a_6950_8596# OUT_N 0.00194f
C116 a_2950_8098# IN_N 9.38e-20
C117 a_2950_8430# OUT_P 8.23e-20
C118 a_n2848_8007# CAL_N 0.050334f
C119 a_n1954_7546# VDD 0.341303f
C120 a_n3230_7261# IN_P 0.060762f
C121 a_n2304_8007# CAL_P 0.007121f
C122 a_468_8407# IN_N 0.395477f
C123 a_n400_8007# EN 0.203816f
C124 a_2588_6962# a_2950_8098# 0.005394f
C125 a_n1954_7546# a_n624_7154# 0.702909f
C126 a_n1438_7546# a_n882_7066# 0.208284f
C127 a_n3230_7261# a_468_6971# 0.947638f
C128 a_468_8407# a_2588_6962# 0.392826f
C129 a_2950_8098# IN_P 3.34e-19
C130 a_6950_8596# OUT_P 0.012307f
C131 a_n3220_7910# CAL_N 0.050259f
C132 a_n2848_8007# CAL_P 0.23462f
C133 a_n2304_8007# EN 0.082942f
C134 a_n400_8007# IN_N 0.158832f
C135 a_468_8407# IN_P 1.12513f
C136 a_n3230_7261# VDD 0.341474f
C137 a_n1954_7546# a_n882_7066# 0.124796f
C138 a_n3230_7261# a_n624_7154# 0.616015f
C139 a_468_8407# a_468_6971# 1.48771f
C140 a_n400_8007# a_2588_6962# 0.081868f
C141 a_2950_8098# VDD 0.035277f
C142 a_n3220_7910# CAL_P 0.04831f
C143 a_n2848_8007# EN 0.268253f
C144 a_n2304_8007# IN_N 3.35861f
C145 a_n400_8007# IN_P 0.309182f
C146 a_468_8407# VDD 1.14768f
C147 a_n1954_7546# a_n1438_7546# 0.212154f
C148 a_n3230_7261# a_n882_7066# 0.143675f
C149 a_468_8407# a_n624_7154# 0.136505f
C150 a_n2304_8007# a_2588_6962# 0.003864f
C151 a_n400_8007# a_468_6971# 0.12419f
C152 a_2950_8430# EN 9.75e-19
C153 a_n2848_8007# IN_N 0.146122f
C154 a_n3220_7910# EN 0.021669f
C155 a_n2304_8007# IN_P 3.12006f
C156 a_n400_8007# VDD 2.50876f
C157 a_n882_7066# a_2950_8098# 0.296258f
C158 a_n3230_7261# a_n1438_7546# 0.093669f
C159 a_468_8407# a_n882_7066# 0.394117f
C160 a_n2304_8007# a_468_6971# 15.051701f
C161 a_n400_8007# a_n624_7154# 7.59e-20
C162 a_n3220_7910# IN_N 0.40985f
C163 a_n2848_8007# IN_P 0.101447f
C164 a_n2304_8007# VDD 18.2688f
C165 a_2588_6962# a_2950_8430# 1.48e-20
C166 a_n3230_7261# a_n1954_7546# 1.35509f
C167 a_468_8407# a_n1438_7546# 0.896828f
C168 a_n2848_8007# a_468_6971# 4.96e-20
C169 a_n2304_8007# a_n624_7154# 0.339465f
C170 a_n3220_7910# a_2588_6962# 0.301877f
C171 a_n400_8007# a_n882_7066# 3.02e-20
C172 a_n3220_7910# IN_P 0.334395f
C173 a_n2848_8007# VDD 8.74726f
C174 a_468_8407# a_n1954_7546# 0.189392f
C175 a_n400_8007# a_n1438_7546# 0.473597f
C176 a_n2304_8007# a_n882_7066# 0.575911f
C177 a_n3220_7910# a_468_6971# 0.037095f
C178 a_2950_8430# VDD 0.038604f
C179 a_n3220_7910# VDD 12.7771f
C180 a_468_8407# a_n3230_7261# 0.166912f
C181 a_n2304_8007# a_n1438_7546# 0.331796f
C182 a_n400_8007# a_n1954_7546# 0.5545f
C183 a_n2848_8007# a_n882_7066# 7.39e-19
C184 a_n3220_7910# a_n624_7154# 0.006212f
C185 a_468_8407# a_2950_8098# 0.288061f
C186 a_n2304_8007# a_n1954_7546# 0.267651f
C187 a_n2848_8007# a_n1438_7546# 0.072616f
C188 a_n3220_7910# a_n882_7066# 0.111791f
C189 a_n400_8007# a_n3230_7261# 0.059662f
C190 a_n400_8007# a_2950_8098# 0.037604f
C191 a_n2848_8007# a_n1954_7546# 0.11542f
C192 a_n3220_7910# a_n1438_7546# 0.030623f
C193 a_n2304_8007# a_n3230_7261# 0.426772f
C194 a_n400_8007# a_468_8407# 0.632585f
C195 a_n2304_8007# a_2950_8098# 5.52e-19
C196 a_n400_8007# a_6950_8264# 0.02792f
C197 a_n3220_7910# a_n1954_7546# 0.021358f
C198 a_n2848_8007# a_n3230_7261# 0.046219f
C199 a_n2304_8007# a_468_8407# 16.190699f
C200 a_n3220_7910# a_n3230_7261# 0.013981f
C201 a_n2848_8007# a_468_8407# 0.005271f
C202 a_n2304_8007# a_n400_8007# 1.88343f
C203 a_2950_8430# a_2950_8098# 0.296258f
C204 a_n3220_7910# a_468_8407# 0.036831f
C205 a_n2848_8007# a_n400_8007# 0.078412f
C206 a_n400_8007# a_2950_8430# 0.209356f
C207 a_n2848_8007# a_n2304_8007# 1.26605f
C208 a_n3220_7910# a_n400_8007# 0.191861f
C209 a_6950_8596# a_6950_8264# 0.296258f
C210 a_n2304_8007# a_2950_8430# 6.06e-19
C211 a_n400_8007# a_6950_8596# 2.48e-19
C212 a_n3220_7910# a_n2304_8007# 1.81084f
C213 a_n3220_7910# a_n2848_8007# 0.736866f
C214 OUT_N VSS 2.17977f
C215 OUT_P VSS 2.54762f
C216 CAL_N VSS 0.570553f
C217 CAL_P VSS 0.303092f
C218 EN VSS 4.22554f
C219 IN_N VSS 0.962271f
C220 IN_P VSS 0.871953f
C221 VDD VSS 61.8014f
C222 a_2950_8098# VSS 0.351821f
C223 a_6950_8264# VSS 0.389079f
C224 a_2950_8430# VSS 0.329713f
C225 a_6950_8596# VSS 0.401983f
C226 a_2950_8762# VSS 0.330267f
C227 a_6950_8928# VSS 0.401172f
C228 a_2950_9094# VSS 0.340541f
C229 a_6950_9426# VSS 0.671366f
C230 a_2588_6962# VSS 2.61317f
C231 a_468_6971# VSS 1.32264f
C232 a_n624_7154# VSS 3.39812f
C233 a_n882_7066# VSS 2.83787f
C234 a_n1438_7546# VSS 2.3787f
C235 a_n1954_7546# VSS 3.72242f
C236 a_n3230_7261# VSS 2.41539f
C237 a_468_8407# VSS 1.88486f
C238 a_n400_8007# VSS 4.47f
C239 a_n2304_8007# VSS 1.84889f
C240 a_n2848_8007# VSS 0.838443f
C241 a_n3220_7910# VSS 2.77006f
.ends
