magic
tech sky130A
magscale 1 2
timestamp 1711797897
<< error_p >>
rect -415 445 -353 451
rect -287 445 -225 451
rect -159 445 -97 451
rect -31 445 31 451
rect 97 445 159 451
rect 225 445 287 451
rect 353 445 415 451
rect -415 411 -403 445
rect -287 411 -275 445
rect -159 411 -147 445
rect -31 411 -19 445
rect 97 411 109 445
rect 225 411 237 445
rect 353 411 365 445
rect -415 405 -353 411
rect -287 405 -225 411
rect -159 405 -97 411
rect -31 405 31 411
rect 97 405 159 411
rect 225 405 287 411
rect 353 405 415 411
<< nwell >>
rect -513 -498 513 464
<< pmoslvt >>
rect -419 -436 -349 364
rect -291 -436 -221 364
rect -163 -436 -93 364
rect -35 -436 35 364
rect 93 -436 163 364
rect 221 -436 291 364
rect 349 -436 419 364
<< pdiff >>
rect -477 352 -419 364
rect -477 -424 -465 352
rect -431 -424 -419 352
rect -477 -436 -419 -424
rect -349 352 -291 364
rect -349 -424 -337 352
rect -303 -424 -291 352
rect -349 -436 -291 -424
rect -221 352 -163 364
rect -221 -424 -209 352
rect -175 -424 -163 352
rect -221 -436 -163 -424
rect -93 352 -35 364
rect -93 -424 -81 352
rect -47 -424 -35 352
rect -93 -436 -35 -424
rect 35 352 93 364
rect 35 -424 47 352
rect 81 -424 93 352
rect 35 -436 93 -424
rect 163 352 221 364
rect 163 -424 175 352
rect 209 -424 221 352
rect 163 -436 221 -424
rect 291 352 349 364
rect 291 -424 303 352
rect 337 -424 349 352
rect 291 -436 349 -424
rect 419 352 477 364
rect 419 -424 431 352
rect 465 -424 477 352
rect 419 -436 477 -424
<< pdiffc >>
rect -465 -424 -431 352
rect -337 -424 -303 352
rect -209 -424 -175 352
rect -81 -424 -47 352
rect 47 -424 81 352
rect 175 -424 209 352
rect 303 -424 337 352
rect 431 -424 465 352
<< poly >>
rect -419 445 -349 461
rect -419 411 -403 445
rect -365 411 -349 445
rect -419 364 -349 411
rect -291 445 -221 461
rect -291 411 -275 445
rect -237 411 -221 445
rect -291 364 -221 411
rect -163 445 -93 461
rect -163 411 -147 445
rect -109 411 -93 445
rect -163 364 -93 411
rect -35 445 35 461
rect -35 411 -19 445
rect 19 411 35 445
rect -35 364 35 411
rect 93 445 163 461
rect 93 411 109 445
rect 147 411 163 445
rect 93 364 163 411
rect 221 445 291 461
rect 221 411 237 445
rect 275 411 291 445
rect 221 364 291 411
rect 349 445 419 461
rect 349 411 365 445
rect 403 411 419 445
rect 349 364 419 411
rect -419 -462 -349 -436
rect -291 -462 -221 -436
rect -163 -462 -93 -436
rect -35 -462 35 -436
rect 93 -462 163 -436
rect 221 -462 291 -436
rect 349 -462 419 -436
<< polycont >>
rect -403 411 -365 445
rect -275 411 -237 445
rect -147 411 -109 445
rect -19 411 19 445
rect 109 411 147 445
rect 237 411 275 445
rect 365 411 403 445
<< locali >>
rect -419 411 -403 445
rect -365 411 -349 445
rect -291 411 -275 445
rect -237 411 -221 445
rect -163 411 -147 445
rect -109 411 -93 445
rect -35 411 -19 445
rect 19 411 35 445
rect 93 411 109 445
rect 147 411 163 445
rect 221 411 237 445
rect 275 411 291 445
rect 349 411 365 445
rect 403 411 419 445
rect -465 352 -431 368
rect -465 -440 -431 -424
rect -337 352 -303 368
rect -337 -440 -303 -424
rect -209 352 -175 368
rect -209 -440 -175 -424
rect -81 352 -47 368
rect -81 -440 -47 -424
rect 47 352 81 368
rect 47 -440 81 -424
rect 175 352 209 368
rect 175 -440 209 -424
rect 303 352 337 368
rect 303 -440 337 -424
rect 431 352 465 368
rect 431 -440 465 -424
<< viali >>
rect -403 411 -365 445
rect -275 411 -237 445
rect -147 411 -109 445
rect -19 411 19 445
rect 109 411 147 445
rect 237 411 275 445
rect 365 411 403 445
rect -465 -424 -431 352
rect -337 -424 -303 352
rect -209 -424 -175 352
rect -81 -424 -47 352
rect 47 -424 81 352
rect 175 -424 209 352
rect 303 -424 337 352
rect 431 -424 465 352
<< metal1 >>
rect -415 445 -353 451
rect -415 411 -403 445
rect -365 411 -353 445
rect -415 405 -353 411
rect -287 445 -225 451
rect -287 411 -275 445
rect -237 411 -225 445
rect -287 405 -225 411
rect -159 445 -97 451
rect -159 411 -147 445
rect -109 411 -97 445
rect -159 405 -97 411
rect -31 445 31 451
rect -31 411 -19 445
rect 19 411 31 445
rect -31 405 31 411
rect 97 445 159 451
rect 97 411 109 445
rect 147 411 159 445
rect 97 405 159 411
rect 225 445 287 451
rect 225 411 237 445
rect 275 411 287 445
rect 225 405 287 411
rect 353 445 415 451
rect 353 411 365 445
rect 403 411 415 445
rect 353 405 415 411
rect -471 352 -425 364
rect -471 -424 -465 352
rect -431 -424 -425 352
rect -471 -436 -425 -424
rect -343 352 -297 364
rect -343 -424 -337 352
rect -303 -424 -297 352
rect -343 -436 -297 -424
rect -215 352 -169 364
rect -215 -424 -209 352
rect -175 -424 -169 352
rect -215 -436 -169 -424
rect -87 352 -41 364
rect -87 -424 -81 352
rect -47 -424 -41 352
rect -87 -436 -41 -424
rect 41 352 87 364
rect 41 -424 47 352
rect 81 -424 87 352
rect 41 -436 87 -424
rect 169 352 215 364
rect 169 -424 175 352
rect 209 -424 215 352
rect 169 -436 215 -424
rect 297 352 343 364
rect 297 -424 303 352
rect 337 -424 343 352
rect 297 -436 343 -424
rect 425 352 471 364
rect 425 -424 431 352
rect 465 -424 471 352
rect 425 -436 471 -424
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 4 l 0.35 m 1 nf 7 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
