magic
tech sky130A
magscale 1 2
timestamp 1711964565
<< error_p >>
rect -29 872 29 878
rect -29 838 -17 872
rect -29 832 29 838
rect -29 -838 29 -832
rect -29 -872 -17 -838
rect -29 -878 29 -872
<< pwell >>
rect -211 -1010 211 1010
<< nmos >>
rect -15 -800 15 800
<< ndiff >>
rect -73 788 -15 800
rect -73 -788 -61 788
rect -27 -788 -15 788
rect -73 -800 -15 -788
rect 15 788 73 800
rect 15 -788 27 788
rect 61 -788 73 788
rect 15 -800 73 -788
<< ndiffc >>
rect -61 -788 -27 788
rect 27 -788 61 788
<< psubdiff >>
rect -175 940 175 974
rect -175 878 -141 940
rect 141 878 175 940
rect -175 -940 -141 -878
rect 141 -940 175 -878
rect -175 -974 -79 -940
rect 79 -974 175 -940
<< psubdiffcont >>
rect -175 -878 -141 878
rect 141 -878 175 878
rect -79 -974 79 -940
<< poly >>
rect -33 872 33 888
rect -33 838 -17 872
rect 17 838 33 872
rect -33 822 33 838
rect -15 800 15 822
rect -15 -822 15 -800
rect -33 -838 33 -822
rect -33 -872 -17 -838
rect 17 -872 33 -838
rect -33 -888 33 -872
<< polycont >>
rect -17 838 17 872
rect -17 -872 17 -838
<< locali >>
rect -175 940 175 974
rect -175 878 -141 940
rect 141 878 175 940
rect -33 838 -17 872
rect 17 838 33 872
rect -61 788 -27 804
rect -61 -804 -27 -788
rect 27 788 61 804
rect 27 -804 61 -788
rect -33 -872 -17 -838
rect 17 -872 33 -838
rect -175 -940 -141 -878
rect 141 -940 175 -878
rect -175 -974 -79 -940
rect 79 -974 175 -940
<< viali >>
rect -17 838 17 872
rect -61 -788 -27 788
rect 27 -788 61 788
rect -17 -872 17 -838
<< metal1 >>
rect -29 872 29 878
rect -29 838 -17 872
rect 17 838 29 872
rect -29 832 29 838
rect -67 788 -21 800
rect -67 -788 -61 788
rect -27 -788 -21 788
rect -67 -800 -21 -788
rect 21 788 67 800
rect 21 -788 27 788
rect 61 -788 67 788
rect 21 -800 67 -788
rect -29 -838 29 -832
rect -29 -872 -17 -838
rect 17 -872 29 -838
rect -29 -878 29 -872
<< properties >>
string FIXED_BBOX -158 -957 158 957
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
