magic
tech sky130A
magscale 1 2
timestamp 1713906399
<< error_s >>
rect -5320 41455 -5310 41468
rect -5250 41455 -5240 41468
rect -5213 41380 -5206 41530
rect -5185 41408 -5178 41558
rect -5153 41380 -5131 41530
rect -5125 41408 -5095 41558
rect -5086 41380 -5067 41530
rect -5039 41408 -5035 41558
rect -5011 41380 -5007 41530
rect -4913 41380 -4906 41530
rect -4885 41408 -4878 41558
rect -4853 41380 -4831 41530
rect -4825 41408 -4795 41558
rect -4786 41380 -4767 41530
rect -4738 41408 -4735 41558
rect -4710 41380 -4707 41530
rect -4613 41380 -4606 41530
rect -4585 41408 -4578 41558
rect -4553 41380 -4531 41530
rect -4525 41408 -4495 41558
rect -4486 41380 -4467 41530
rect -5213 36290 -5206 36350
rect -5185 36262 -5178 36322
rect -5153 36290 -5131 36350
rect -5125 36262 -5095 36322
rect -5086 36290 -5067 36350
rect -5039 36262 -5035 36322
rect -5011 36290 -5007 36350
rect -4913 36290 -4906 36350
rect -4885 36262 -4878 36322
rect -4853 36290 -4831 36350
rect -4825 36262 -4795 36322
rect -4786 36290 -4767 36350
rect -4739 36262 -4735 36322
rect -4711 36290 -4707 36350
rect -4613 36290 -4606 36350
rect -4585 36262 -4578 36322
rect -4553 36290 -4531 36350
rect -4525 36262 -4495 36322
rect -4486 36290 -4467 36350
rect -4454 36262 -4435 36322
rect -4426 36290 -4407 36350
rect -4394 36262 -4375 36322
rect -4366 36290 -4347 36350
rect -4334 36262 -4315 36322
rect -4306 36290 -4287 36350
rect -4274 36262 -4255 36322
rect -4246 36290 -4227 36350
rect -4214 36262 -4195 36322
rect -4186 36290 -4167 36350
rect -4154 36262 -4135 36322
rect -4126 36290 -4107 36350
rect -4094 36262 -4075 36322
rect -4066 36290 -4047 36350
rect -4034 36262 -4015 36322
rect -4006 36290 -3987 36350
rect -3974 36262 -3950 36322
rect -3946 36290 -3916 36350
rect -3895 36262 -3888 36322
<< metal1 >>
rect 10980 48530 10990 48590
rect 11050 48568 11060 48590
rect 11050 48540 24074 48568
rect 11050 48530 11060 48540
rect -3925 48470 -3865 48480
rect -3925 48400 -3865 48410
rect -4005 48210 -3945 48220
rect -4005 48140 -3945 48150
rect -4075 47940 -4015 47950
rect -4075 47870 -4015 47880
rect -4135 47660 -4075 47670
rect -4135 47590 -4075 47600
rect -4195 47390 -4135 47400
rect -4195 47320 -4135 47330
rect -4255 47110 -4195 47120
rect -4255 47040 -4195 47050
rect -4315 46850 -4255 46860
rect -4315 46780 -4255 46790
rect -4375 46580 -4315 46590
rect -4375 46510 -4315 46520
rect -4435 46300 -4375 46310
rect -4435 46230 -4375 46240
rect -4495 46030 -4435 46040
rect -4495 45960 -4435 45970
rect -4555 45770 -4495 45780
rect -4555 45700 -4495 45710
rect -4615 45490 -4555 45500
rect -4615 45420 -4555 45430
rect -4675 45220 -4615 45230
rect -4675 45150 -4615 45160
rect -4735 44940 -4675 44950
rect -4735 44870 -4675 44880
rect -4795 44680 -4735 44690
rect -4795 44610 -4735 44620
rect -4855 44410 -4795 44420
rect -4855 44340 -4795 44350
rect -4915 44140 -4855 44150
rect -4915 44070 -4855 44080
rect -4975 43850 -4915 43860
rect -4975 43780 -4915 43790
rect -5035 43580 -4975 43590
rect -5035 43510 -4975 43520
rect -5095 43320 -5035 43330
rect -5095 43250 -5035 43260
rect -5155 43030 -5095 43040
rect -5155 42960 -5095 42970
rect -5215 42760 -5155 42770
rect -5215 42690 -5155 42700
rect -5275 42480 -5215 42490
rect -5275 42410 -5215 42420
rect -5245 41408 -5215 42410
rect -5185 41408 -5155 42690
rect -5125 41408 -5095 42960
rect -5065 41408 -5035 43250
rect -5005 41408 -4975 43510
rect -4945 41408 -4915 43780
rect -4885 41408 -4855 44070
rect -4825 41408 -4795 44340
rect -4765 41408 -4735 44610
rect -4705 41408 -4675 44870
rect -4645 41408 -4615 45150
rect -4585 41408 -4555 45420
rect -4525 41408 -4495 45700
rect -4465 41408 -4435 45960
rect -4405 41408 -4375 46230
rect -4345 41408 -4315 46510
rect -4285 41408 -4255 46780
rect -4225 41408 -4195 47040
rect -4165 41408 -4135 47320
rect -4105 41408 -4075 47590
rect -4045 41408 -4015 47870
rect -3980 41408 -3950 48140
rect -3895 41408 -3865 48400
rect 15080 42261 15090 42321
rect 15150 42305 15160 42321
rect 24046 42305 24074 48540
rect 15150 42277 24074 42305
rect 24152 48490 24212 48500
rect 24152 48420 24212 48430
rect 15150 42261 15160 42277
rect 15390 42180 15400 42240
rect 15460 42220 15470 42240
rect 16590 42220 16600 42240
rect 15460 42190 16600 42220
rect 15460 42180 15470 42190
rect 16590 42180 16600 42190
rect 16660 42180 16670 42240
rect 22750 42170 22760 42240
rect 22830 42220 22840 42240
rect 23190 42220 23200 42240
rect 22830 42190 23200 42220
rect 22830 42170 22840 42190
rect 23190 42180 23200 42190
rect 23260 42180 23270 42240
rect -2731 42067 -2721 42127
rect -2661 42110 -2651 42127
rect 1130 42110 1140 42130
rect -2661 42080 1140 42110
rect -2661 42067 -2651 42080
rect 1130 42070 1140 42080
rect 1200 42110 1210 42130
rect 14470 42110 14480 42130
rect 1200 42080 14480 42110
rect 1200 42070 1210 42080
rect 14470 42070 14480 42080
rect 14540 42070 14550 42130
rect 14970 42100 14980 42160
rect 15040 42150 15050 42160
rect 20280 42150 20290 42160
rect 15040 42120 20290 42150
rect 15040 42100 15050 42120
rect 20280 42100 20290 42120
rect 20345 42100 20355 42160
rect 15260 42030 15270 42090
rect 15330 42070 15340 42090
rect 15330 42040 24092 42070
rect 15330 42030 15340 42040
rect -1807 41964 -1797 42017
rect -1744 42000 -1734 42017
rect 2330 42000 2340 42030
rect -1744 41970 2340 42000
rect 2400 42000 2410 42030
rect 2400 41970 23770 42000
rect -1744 41964 -1734 41970
rect 23760 41940 23770 41970
rect 23830 41940 23840 42000
rect 23760 41930 23840 41940
rect -888 41860 -878 41912
rect -823 41901 -813 41912
rect 3357 41901 3367 41915
rect -823 41871 3367 41901
rect -823 41860 -813 41871
rect 3357 41855 3367 41871
rect 3427 41855 3437 41915
rect 14470 41870 14480 41930
rect 14540 41920 14550 41930
rect 14540 41910 23730 41920
rect 14540 41890 23660 41910
rect 14540 41870 14550 41890
rect 18430 41825 18440 41860
rect -3272 41790 -3262 41815
rect -3805 41760 -3262 41790
rect -3805 41408 -3775 41760
rect -3272 41755 -3262 41760
rect -3202 41790 -3192 41815
rect 15260 41790 15270 41810
rect -3202 41760 15270 41790
rect -3202 41755 -3192 41760
rect 15260 41750 15270 41760
rect 15330 41750 15340 41810
rect 15500 41800 18440 41825
rect 18500 41800 18510 41860
rect 23650 41850 23660 41890
rect 23720 41850 23730 41910
rect 15500 41795 18510 41800
rect 15380 41510 15390 41570
rect 15450 41510 15470 41570
rect 14750 41420 14760 41480
rect 14820 41465 14830 41480
rect 14820 41435 15410 41465
rect 14820 41420 14830 41435
rect 12910 41330 12920 41390
rect 12980 41375 12990 41390
rect 12980 41345 15350 41375
rect 12980 41330 12990 41345
rect 960 41240 970 41300
rect 1030 41285 1040 41300
rect 1030 41255 15290 41285
rect 1030 41240 1040 41255
rect 2790 41150 2800 41210
rect 2860 41195 2870 41210
rect 2860 41165 15230 41195
rect 2860 41150 2870 41165
rect 12000 41105 12010 41120
rect 185 41075 12010 41105
rect 185 36490 215 41075
rect 12000 41060 12010 41075
rect 12070 41060 12080 41120
rect 15080 41040 15090 41100
rect 15150 41040 15160 41100
rect 10150 41015 10160 41030
rect 245 40985 10160 41015
rect 245 36550 275 40985
rect 10150 40970 10160 40985
rect 10220 40970 10230 41030
rect 8310 40925 8320 40940
rect 305 40895 8320 40925
rect 305 36610 335 40895
rect 8310 40880 8320 40895
rect 8380 40880 8390 40940
rect 14970 40835 14980 40850
rect 365 40805 14980 40835
rect 365 36670 395 40805
rect 14970 40790 14980 40805
rect 15040 40790 15050 40850
rect 6450 40745 6460 40750
rect 425 40715 6460 40745
rect 425 36730 455 40715
rect 6450 40690 6460 40715
rect 6520 40690 6530 40750
rect 4620 40655 4630 40660
rect 485 40625 4630 40655
rect 485 36790 515 40625
rect 4620 40600 4630 40625
rect 4690 40600 4700 40660
rect 2320 40565 2330 40580
rect 595 40535 2330 40565
rect 595 39820 625 40535
rect 2320 40520 2330 40535
rect 2390 40520 2400 40580
rect 3350 40475 3360 40490
rect 545 39760 555 39820
rect 615 39760 625 39820
rect 655 40445 3360 40475
rect 655 39350 685 40445
rect 3350 40430 3360 40445
rect 3420 40430 3430 40490
rect 1140 40385 1150 40400
rect 605 39290 615 39350
rect 675 39290 685 39350
rect 715 40355 1150 40385
rect 715 38730 745 40355
rect 1140 40340 1150 40355
rect 1210 40340 1220 40400
rect 9250 40340 9260 40680
rect 9630 40340 9640 40680
rect 1530 40170 1540 40270
rect 1910 40170 1920 40270
rect 665 38670 675 38730
rect 735 38670 745 38730
rect 3400 38020 3410 38080
rect 3470 38020 3480 38080
rect 14830 38020 14860 38030
rect 3420 37670 3460 38020
rect 14800 37960 14810 38020
rect 14870 38005 14880 38020
rect 15120 38005 15150 41040
rect 14870 37975 15150 38005
rect 14870 37960 14880 37975
rect 3400 37610 3410 37670
rect 3470 37610 3480 37670
rect 1960 37330 2300 37510
rect 1950 36990 1960 37330
rect 2300 36990 2310 37330
rect 7400 36990 7410 37330
rect 7750 36990 7760 37330
rect 15200 36850 15230 41165
rect 10095 36840 15230 36850
rect 485 36780 10035 36790
rect 485 36760 9975 36780
rect 425 36720 9945 36730
rect 425 36700 9885 36720
rect 365 36660 9855 36670
rect 365 36640 9795 36660
rect 305 36600 9765 36610
rect 305 36580 9705 36600
rect 245 36540 9675 36550
rect 245 36520 9615 36540
rect 185 36480 9585 36490
rect 185 36460 9525 36480
rect 10155 36820 15230 36840
rect 15260 36790 15290 41255
rect 10095 36770 10155 36780
rect 10185 36780 15290 36790
rect 9975 36710 10035 36720
rect 10245 36760 15290 36780
rect 15320 36730 15350 41345
rect 10185 36710 10245 36720
rect 10275 36720 15350 36730
rect 9885 36650 9945 36660
rect 10335 36700 15350 36720
rect 15380 36670 15410 41435
rect 10275 36650 10335 36660
rect 10365 36660 15410 36670
rect 9795 36590 9855 36600
rect 10425 36640 15410 36660
rect 15440 36610 15470 41510
rect 10365 36590 10425 36600
rect 10455 36600 15470 36610
rect 9705 36530 9765 36540
rect 10515 36580 15470 36600
rect 15500 36550 15530 41795
rect 21190 41765 21200 41800
rect 10455 36530 10515 36540
rect 10545 36540 15530 36550
rect 9615 36470 9675 36480
rect 10605 36520 15530 36540
rect 15560 41740 21200 41765
rect 21260 41740 21270 41800
rect 15560 41735 21265 41740
rect 15560 36490 15590 41735
rect 17070 41590 17080 41680
rect 17450 41590 17460 41680
rect 22470 41530 22480 41680
rect 23040 41530 23050 41680
rect 23180 41480 23190 41540
rect 23250 41480 23260 41540
rect 23510 41480 23520 41540
rect 23580 41525 23590 41540
rect 23580 41480 23591 41525
rect 23630 41480 23640 41540
rect 23700 41480 23710 41540
rect 23210 41340 23240 41480
rect 23561 39695 23591 41480
rect 23650 40830 23680 41480
rect 23620 40770 23630 40830
rect 23690 40770 23700 40830
rect 15760 39330 15770 39390
rect 15830 39330 15840 39390
rect 15670 38440 15680 38500
rect 15740 38440 15750 38500
rect 15700 37880 15730 38440
rect 15670 37820 15680 37880
rect 15740 37820 15750 37880
rect 15790 37750 15820 39330
rect 15740 37690 15750 37750
rect 15810 37690 15820 37750
rect 10545 36470 10605 36480
rect 10635 36480 15590 36490
rect 9525 36410 9585 36420
rect 10695 36460 15590 36480
rect 10635 36410 10695 36420
rect -5245 36270 -5215 36322
rect -5185 36270 -5155 36322
rect -5125 36270 -5095 36322
rect -5065 36270 -5035 36322
rect -5005 36270 -4975 36322
rect -4945 36270 -4915 36322
rect -4885 36270 -4855 36322
rect -4825 36270 -4795 36322
rect -4765 36270 -4735 36322
rect -4705 36270 -4675 36322
rect -4645 36270 -4615 36322
rect -4585 36270 -4555 36322
rect -4525 36270 -4495 36322
rect -4465 36270 -4435 36322
rect -4405 36270 -4375 36322
rect -4345 36270 -4315 36322
rect -4285 36270 -4255 36322
rect -4225 36270 -4195 36322
rect -4165 36270 -4135 36322
rect -4105 36270 -4075 36322
rect -4045 36270 -4015 36322
rect -3980 36270 -3950 36322
rect -3895 36270 -3865 36322
rect -3805 36270 -3775 36322
rect 24062 36190 24092 42040
rect 24152 36190 24182 48420
rect 24232 48230 24292 48240
rect 24232 48160 24292 48170
rect 24237 36190 24267 48160
rect 24302 47960 24362 47970
rect 24302 47890 24362 47900
rect 24302 36190 24332 47890
rect 24362 47680 24422 47690
rect 24362 47610 24422 47620
rect 24362 36190 24392 47610
rect 24422 47410 24482 47420
rect 24422 47340 24482 47350
rect 24422 36190 24452 47340
rect 24482 47130 24542 47140
rect 24482 47060 24542 47070
rect 24482 36190 24512 47060
rect 24542 46870 24602 46880
rect 24542 46800 24602 46810
rect 24542 36190 24572 46800
rect 24602 46600 24662 46610
rect 24602 46530 24662 46540
rect 24602 36190 24632 46530
rect 24662 46320 24722 46330
rect 24662 46250 24722 46260
rect 24662 36190 24692 46250
rect 24722 46050 24782 46060
rect 24722 45980 24782 45990
rect 24722 36190 24752 45980
rect 24782 45790 24842 45800
rect 24782 45720 24842 45730
rect 24782 36190 24812 45720
rect 24842 45510 24902 45520
rect 24842 45440 24902 45450
rect 24842 36190 24872 45440
rect 24902 45240 24962 45250
rect 24902 45170 24962 45180
rect 24902 36190 24932 45170
rect 24962 44960 25022 44970
rect 24962 44890 25022 44900
rect 24962 36190 24992 44890
rect 25022 44700 25082 44710
rect 25022 44630 25082 44640
rect 25022 36190 25052 44630
rect 25082 44430 25142 44440
rect 25082 44360 25142 44370
rect 25082 36190 25112 44360
rect 25142 44160 25202 44170
rect 25142 44090 25202 44100
rect 25142 36190 25172 44090
rect 25202 43870 25262 43880
rect 25202 43800 25262 43810
rect 25202 36190 25232 43800
rect 25262 43600 25322 43610
rect 25262 43530 25322 43540
rect 25262 36190 25292 43530
rect 25322 43340 25382 43350
rect 25322 43270 25382 43280
rect 25322 36190 25352 43270
rect 25382 43050 25442 43060
rect 25382 42980 25442 42990
rect 25382 36190 25412 42980
rect 25442 42780 25502 42790
rect 25442 42710 25502 42720
rect 25442 36190 25472 42710
rect 25502 42500 25562 42510
rect 25502 42430 25562 42440
rect 25502 36190 25532 42430
rect 10610 33670 10620 33730
rect 10680 33670 10690 33730
rect 10520 33580 10530 33640
rect 10590 33580 10600 33640
rect 10430 33490 10440 33550
rect 10500 33490 10510 33550
rect 10340 33400 10350 33460
rect 10410 33400 10420 33460
rect 10250 33310 10260 33370
rect 10320 33310 10330 33370
rect 10160 33220 10170 33280
rect 10230 33220 10240 33280
rect 10070 33130 10080 33190
rect 10140 33130 10150 33190
rect 9980 33040 9990 33100
rect 10050 33040 10060 33100
rect 9890 32950 9900 33010
rect 9960 32950 9970 33010
rect 9800 32860 9810 32920
rect 9870 32860 9880 32920
rect 9710 32770 9720 32830
rect 9780 32770 9790 32830
rect 9620 32680 9630 32740
rect 9690 32680 9700 32740
rect 9530 32590 9540 32650
rect 9600 32590 9610 32650
<< via1 >>
rect 10990 48530 11050 48590
rect -3925 48410 -3865 48470
rect -4005 48150 -3945 48210
rect -4075 47880 -4015 47940
rect -4135 47600 -4075 47660
rect -4195 47330 -4135 47390
rect -4255 47050 -4195 47110
rect -4315 46790 -4255 46850
rect -4375 46520 -4315 46580
rect -4435 46240 -4375 46300
rect -4495 45970 -4435 46030
rect -4555 45710 -4495 45770
rect -4615 45430 -4555 45490
rect -4675 45160 -4615 45220
rect -4735 44880 -4675 44940
rect -4795 44620 -4735 44680
rect -4855 44350 -4795 44410
rect -4915 44080 -4855 44140
rect -4975 43790 -4915 43850
rect -5035 43520 -4975 43580
rect -5095 43260 -5035 43320
rect -5155 42970 -5095 43030
rect -5215 42700 -5155 42760
rect -5275 42420 -5215 42480
rect 15090 42261 15150 42321
rect 24152 48430 24212 48490
rect 15400 42180 15460 42240
rect 16600 42180 16660 42240
rect 22760 42170 22830 42240
rect 23200 42180 23260 42240
rect -2721 42067 -2661 42127
rect 1140 42070 1200 42130
rect 14480 42070 14540 42130
rect 14980 42100 15040 42160
rect 20290 42100 20345 42160
rect 15270 42030 15330 42090
rect -1797 41964 -1744 42017
rect 2340 41970 2400 42030
rect 23770 41940 23830 42000
rect -878 41860 -823 41912
rect 3367 41855 3427 41915
rect 14480 41870 14540 41930
rect -3262 41755 -3202 41815
rect 15270 41750 15330 41810
rect 18440 41800 18500 41860
rect 23660 41850 23720 41910
rect 15390 41510 15450 41570
rect 14760 41420 14820 41480
rect 12920 41330 12980 41390
rect 970 41240 1030 41300
rect 2800 41150 2860 41210
rect 12010 41060 12070 41120
rect 15090 41040 15150 41100
rect 10160 40970 10220 41030
rect 8320 40880 8380 40940
rect 14980 40790 15040 40850
rect 6460 40690 6520 40750
rect 4630 40600 4690 40660
rect 2330 40520 2390 40580
rect 555 39760 615 39820
rect 3360 40430 3420 40490
rect 615 39290 675 39350
rect 1150 40340 1210 40400
rect 9260 40340 9630 40680
rect 1540 40170 1910 40270
rect 675 38670 735 38730
rect 3410 38020 3470 38080
rect 14810 37960 14870 38020
rect 3410 37610 3470 37670
rect 1960 36990 2300 37330
rect 7410 36990 7750 37330
rect 9525 36420 9585 36480
rect 9615 36480 9675 36540
rect 9705 36540 9765 36600
rect 9795 36600 9855 36660
rect 9885 36660 9945 36720
rect 9975 36720 10035 36780
rect 10095 36780 10155 36840
rect 10185 36720 10245 36780
rect 10275 36660 10335 36720
rect 10365 36600 10425 36660
rect 10455 36540 10515 36600
rect 10545 36480 10605 36540
rect 21200 41740 21260 41800
rect 17080 41590 17450 41680
rect 22480 41530 23040 41680
rect 23190 41480 23250 41540
rect 23520 41480 23580 41540
rect 23640 41480 23700 41540
rect 23630 40770 23690 40830
rect 15770 39330 15830 39390
rect 15680 38440 15740 38500
rect 15680 37820 15740 37880
rect 15750 37690 15810 37750
rect 10635 36420 10695 36480
rect 24232 48170 24292 48230
rect 24302 47900 24362 47960
rect 24362 47620 24422 47680
rect 24422 47350 24482 47410
rect 24482 47070 24542 47130
rect 24542 46810 24602 46870
rect 24602 46540 24662 46600
rect 24662 46260 24722 46320
rect 24722 45990 24782 46050
rect 24782 45730 24842 45790
rect 24842 45450 24902 45510
rect 24902 45180 24962 45240
rect 24962 44900 25022 44960
rect 25022 44640 25082 44700
rect 25082 44370 25142 44430
rect 25142 44100 25202 44160
rect 25202 43810 25262 43870
rect 25262 43540 25322 43600
rect 25322 43280 25382 43340
rect 25382 42990 25442 43050
rect 25442 42720 25502 42780
rect 25502 42440 25562 42500
rect 10620 33670 10680 33730
rect 10530 33580 10590 33640
rect 10440 33490 10500 33550
rect 10350 33400 10410 33460
rect 10260 33310 10320 33370
rect 10170 33220 10230 33280
rect 10080 33130 10140 33190
rect 9990 33040 10050 33100
rect 9900 32950 9960 33010
rect 9810 32860 9870 32920
rect 9720 32770 9780 32830
rect 9630 32680 9690 32740
rect 9540 32590 9600 32650
<< metal2 >>
rect 10990 48590 11050 48600
rect 10990 48520 11050 48530
rect -3540 48480 -3480 48490
rect -3925 48470 -3865 48480
rect -3865 48420 -3540 48450
rect -3540 48410 -3480 48420
rect -3925 48400 -3865 48410
rect -2990 48260 -2940 48440
rect -1150 48280 -1100 48460
rect 410 48290 460 48470
rect 2250 48290 2300 48470
rect 4000 48290 4050 48470
rect 5750 48290 5800 48470
rect 7500 48290 7550 48470
rect 9240 48280 9290 48460
rect -4005 48210 -3945 48220
rect -3540 48200 -3480 48210
rect -3945 48160 -3540 48190
rect -4005 48140 -3945 48150
rect 10990 48192 11046 48520
rect 24152 48490 24212 48500
rect 23950 48480 24010 48490
rect 12740 48260 12790 48440
rect 14490 48240 14540 48420
rect 16240 48240 16290 48420
rect 17990 48290 18040 48470
rect 19730 48250 19780 48430
rect 21480 48270 21530 48450
rect 23230 48280 23280 48460
rect 24010 48440 24152 48470
rect 24152 48420 24212 48430
rect 23950 48410 24010 48420
rect 24232 48230 24292 48240
rect 23950 48210 24010 48220
rect 24010 48180 24232 48210
rect 24232 48160 24292 48170
rect 23950 48140 24010 48150
rect -3540 48130 -3480 48140
rect 24302 47960 24362 47970
rect -4075 47940 -4015 47950
rect -3540 47940 -3480 47950
rect -4015 47890 -3540 47920
rect -4075 47870 -4015 47880
rect -3540 47870 -3480 47880
rect 23950 47940 24010 47950
rect 24010 47910 24302 47940
rect 24302 47890 24362 47900
rect 23950 47870 24010 47880
rect 24362 47680 24422 47690
rect 23950 47670 24010 47680
rect -4135 47660 -4075 47670
rect -3540 47660 -3480 47670
rect -4075 47610 -3540 47640
rect -4135 47590 -4075 47600
rect 24010 47630 24362 47660
rect 24362 47610 24422 47620
rect 23950 47600 24010 47610
rect -3540 47590 -3480 47600
rect 24422 47410 24482 47420
rect -4195 47390 -4135 47400
rect -3550 47390 -3490 47400
rect -4135 47340 -3550 47370
rect -4195 47320 -4135 47330
rect -3550 47320 -3490 47330
rect 23950 47390 24010 47400
rect 24010 47360 24422 47390
rect 24422 47340 24482 47350
rect 23950 47320 24010 47330
rect 24482 47130 24542 47140
rect -3550 47120 -3490 47130
rect -4255 47110 -4195 47120
rect -4195 47060 -3550 47090
rect -3550 47050 -3490 47060
rect 23950 47110 24010 47120
rect 24010 47080 24482 47110
rect 24482 47060 24542 47070
rect -4255 47040 -4195 47050
rect 23950 47040 24010 47050
rect 24542 46870 24602 46880
rect -4315 46850 -4255 46860
rect -3540 46850 -3480 46860
rect -4255 46800 -3540 46830
rect -4315 46780 -4255 46790
rect -3540 46780 -3480 46790
rect 23950 46850 24010 46860
rect 24010 46820 24542 46850
rect 24542 46800 24602 46810
rect 23950 46780 24010 46790
rect 24602 46600 24662 46610
rect -4375 46580 -4315 46590
rect -3550 46580 -3490 46590
rect -4315 46530 -3550 46560
rect -4375 46510 -4315 46520
rect -3550 46510 -3490 46520
rect 23950 46580 24010 46590
rect 24010 46550 24602 46580
rect 24602 46530 24662 46540
rect 23950 46510 24010 46520
rect 24662 46320 24722 46330
rect -3540 46310 -3480 46320
rect -4435 46300 -4375 46310
rect -4375 46250 -3540 46280
rect -3540 46240 -3480 46250
rect 23950 46310 24010 46320
rect 24010 46270 24662 46300
rect 24662 46250 24722 46260
rect 23950 46240 24010 46250
rect -4435 46230 -4375 46240
rect 24722 46050 24782 46060
rect -3540 46040 -3480 46050
rect -4495 46030 -4435 46040
rect -4435 45980 -3540 46010
rect -3540 45970 -3480 45980
rect 23950 46030 24010 46040
rect 24010 46000 24722 46030
rect 24722 45980 24782 45990
rect -4495 45960 -4435 45970
rect 23950 45960 24010 45970
rect 24782 45790 24842 45800
rect -4555 45770 -4495 45780
rect 23950 45770 24010 45780
rect -3540 45760 -3480 45770
rect -4495 45720 -3540 45750
rect -4555 45700 -4495 45710
rect 24010 45740 24782 45770
rect 24782 45720 24842 45730
rect 23950 45700 24010 45710
rect -3540 45690 -3480 45700
rect 24842 45510 24902 45520
rect 23950 45500 24010 45510
rect -4615 45490 -4555 45500
rect -3540 45490 -3480 45500
rect -4555 45440 -3540 45470
rect -4615 45420 -4555 45430
rect 24010 45460 24842 45490
rect 24842 45440 24902 45450
rect 23950 45430 24010 45440
rect -3540 45420 -3480 45430
rect 24902 45240 24962 45250
rect 23950 45230 24010 45240
rect -4675 45220 -4615 45230
rect -3540 45210 -3480 45220
rect -4615 45170 -3540 45200
rect -4675 45150 -4615 45160
rect 24010 45190 24902 45220
rect 24902 45170 24962 45180
rect 23950 45160 24010 45170
rect -3540 45140 -3480 45150
rect 24962 44960 25022 44970
rect 23950 44950 24010 44960
rect -4735 44940 -4675 44950
rect -3540 44940 -3480 44950
rect -4675 44890 -3540 44920
rect -4735 44870 -4675 44880
rect 24010 44910 24962 44940
rect 24962 44890 25022 44900
rect 23950 44880 24010 44890
rect -3540 44870 -3480 44880
rect 25022 44700 25082 44710
rect 23950 44690 24010 44700
rect -4795 44680 -4735 44690
rect -3540 44670 -3480 44680
rect -4735 44630 -3540 44660
rect -4795 44610 -4735 44620
rect 24010 44650 25022 44680
rect 25022 44630 25082 44640
rect 23950 44620 24010 44630
rect -3540 44600 -3480 44610
rect 25082 44430 25142 44440
rect -4855 44410 -4795 44420
rect 23950 44410 24010 44420
rect -3540 44400 -3480 44410
rect -4795 44360 -3540 44390
rect -4855 44340 -4795 44350
rect 24010 44380 25082 44410
rect 25082 44360 25142 44370
rect 23950 44340 24010 44350
rect -3540 44330 -3480 44340
rect 25142 44160 25202 44170
rect -4915 44140 -4855 44150
rect 23950 44140 24010 44150
rect -3540 44130 -3480 44140
rect -4855 44090 -3540 44120
rect -4915 44070 -4855 44080
rect 24010 44110 25142 44140
rect 25142 44090 25202 44100
rect 23950 44070 24010 44080
rect -3540 44060 -3480 44070
rect 25202 43870 25262 43880
rect -3540 43860 -3480 43870
rect -4975 43850 -4915 43860
rect -4915 43800 -3540 43830
rect -3540 43790 -3480 43800
rect 23950 43860 24010 43870
rect 24010 43820 25202 43850
rect 25202 43800 25262 43810
rect 23950 43790 24010 43800
rect -4975 43780 -4915 43790
rect 25262 43600 25322 43610
rect -3540 43590 -3480 43600
rect -5035 43580 -4975 43590
rect -4975 43530 -3540 43560
rect 23960 43590 24020 43600
rect 23957 43550 23960 43580
rect -3540 43520 -3480 43530
rect 24020 43550 25262 43580
rect 25262 43530 25322 43540
rect 23960 43520 24020 43530
rect -5035 43510 -4975 43520
rect 25322 43340 25382 43350
rect 23950 43330 24010 43340
rect -5095 43320 -5035 43330
rect -3540 43320 -3480 43330
rect -5035 43270 -3540 43300
rect -5095 43250 -5035 43260
rect 24010 43290 25322 43320
rect 25322 43270 25382 43280
rect 23950 43260 24010 43270
rect -3540 43250 -3480 43260
rect -3540 43050 -3480 43060
rect 25382 43050 25442 43060
rect -5155 43030 -5095 43040
rect -5095 42990 -3540 43010
rect -5095 42980 -3480 42990
rect 23950 43040 24010 43050
rect 24010 43000 25382 43030
rect 25382 42980 25442 42990
rect 23950 42970 24010 42980
rect -5155 42960 -5095 42970
rect -3540 42780 -3480 42790
rect -5215 42760 -5155 42770
rect -5155 42720 -3540 42740
rect -5155 42710 -3480 42720
rect 23950 42780 24010 42790
rect 25442 42780 25502 42790
rect 24010 42730 25442 42760
rect 23950 42710 24010 42720
rect 25442 42710 25502 42720
rect -5215 42690 -5155 42700
rect 15696 42554 15724 42614
rect -5275 42480 -5215 42490
rect -3540 42470 -3480 42480
rect -5215 42430 -3540 42460
rect -5275 42410 -5215 42420
rect -3540 42400 -3480 42410
rect 2816 42354 2844 42534
rect 8336 42474 8364 42554
rect 10176 42494 10204 42534
rect 12016 42494 12044 42534
rect 14786 42526 15724 42554
rect 17536 42544 17564 42614
rect 16616 42516 17564 42544
rect 7440 42446 8364 42474
rect 9266 42466 10204 42494
rect 11106 42466 12044 42494
rect 6496 42414 6524 42434
rect 4656 42354 4684 42414
rect 5586 42386 6524 42414
rect 976 42258 1004 42346
rect 1906 42326 2844 42354
rect 3746 42326 4684 42354
rect 19376 42344 19404 42454
rect 22136 42354 22164 42534
rect 23940 42500 24000 42510
rect 25502 42500 25562 42510
rect 24000 42450 25502 42480
rect 23940 42430 24000 42440
rect 25502 42430 25562 42440
rect 15090 42321 15150 42331
rect 62 42230 1004 42258
rect 13856 42174 13884 42314
rect 18466 42316 19404 42344
rect 21226 42326 22164 42354
rect 15090 42251 15150 42261
rect 12946 42146 13884 42174
rect 14980 42160 15040 42170
rect -2721 42127 -2661 42137
rect -2721 42057 -2661 42067
rect 1140 42130 1200 42140
rect 14480 42130 14540 42140
rect 1140 42060 1200 42070
rect -1797 42017 -1744 42027
rect -1797 41954 -1744 41964
rect -878 41912 -823 41922
rect -3260 41825 -3204 41908
rect -878 41850 -823 41860
rect -3262 41815 -3202 41825
rect -5050 41780 -4990 41790
rect -3660 41780 -3580 41790
rect -4990 41700 -3660 41780
rect -3262 41745 -3202 41755
rect -5050 41690 -4990 41700
rect -3660 41690 -3580 41700
rect -4790 41620 -4730 41630
rect -3660 41620 -3580 41630
rect -4730 41540 -3660 41620
rect -4790 41530 -4730 41540
rect -3660 41530 -3580 41540
rect 980 41310 1010 41935
rect 970 41300 1030 41310
rect 970 41230 1030 41240
rect -100 40680 240 40690
rect 1160 40410 1190 42060
rect 2350 42040 2380 42045
rect 2340 42030 2400 42040
rect 2340 41960 2400 41970
rect 1540 40680 1910 40690
rect -100 40330 240 40340
rect 1150 40400 1210 40410
rect 1150 40330 1210 40340
rect 2350 40590 2380 41960
rect 3367 41915 3427 41925
rect 2820 41220 2850 41895
rect 3367 41845 3427 41855
rect 2800 41210 2860 41220
rect 2800 41140 2860 41150
rect 2330 40580 2390 40590
rect 2330 40510 2390 40520
rect 3380 40500 3410 41845
rect 4640 40670 4670 41920
rect 6480 40760 6510 41960
rect 8330 40950 8360 41940
rect 10170 41040 10200 41920
rect 12020 41130 12050 42110
rect 14980 42090 15040 42100
rect 14480 42060 14540 42070
rect 12940 41400 12970 41970
rect 14490 41940 14530 42060
rect 14480 41930 14540 41940
rect 14480 41860 14540 41870
rect 14780 41490 14810 42055
rect 14760 41480 14820 41490
rect 14760 41410 14820 41420
rect 12920 41390 12980 41400
rect 12920 41320 12980 41330
rect 12010 41120 12070 41130
rect 12010 41050 12070 41060
rect 10160 41030 10220 41040
rect 10160 40960 10220 40970
rect 8320 40940 8380 40950
rect 8320 40870 8380 40880
rect 15000 40860 15030 42090
rect 15110 41110 15140 42251
rect 15400 42240 15460 42250
rect 15400 42170 15460 42180
rect 16600 42240 16660 42250
rect 16600 42170 16660 42180
rect 22760 42240 22830 42250
rect 23200 42240 23260 42250
rect 23200 42170 23260 42180
rect 15270 42090 15330 42100
rect 15270 42020 15330 42030
rect 15280 41820 15310 42020
rect 15270 41810 15330 41820
rect 15270 41740 15330 41750
rect 15410 41580 15440 42170
rect 20290 42160 20345 42170
rect 22760 42160 22830 42170
rect 20290 42090 20345 42100
rect 18440 41860 18500 41870
rect 18440 41790 18500 41800
rect 21200 41800 21260 41890
rect 21200 41730 21260 41740
rect 17080 41680 17450 41690
rect 15390 41570 15450 41580
rect 15390 41500 15450 41510
rect 15090 41100 15150 41110
rect 15090 41030 15150 41040
rect 14980 40850 15040 40860
rect 14980 40780 15040 40790
rect 6460 40750 6520 40760
rect 6460 40680 6520 40690
rect 9260 40680 9630 40690
rect 4630 40660 4690 40670
rect 4630 40590 4690 40600
rect 3360 40490 3420 40500
rect 3360 40420 3420 40430
rect 1540 40270 1910 40340
rect 9260 40330 9630 40340
rect 17080 40680 17450 41590
rect 22480 41680 23040 41690
rect 23210 41550 23240 42170
rect 23770 42000 23830 42010
rect 23770 41930 23830 41940
rect 23660 41910 23720 41920
rect 23540 41550 23570 41875
rect 23660 41840 23720 41850
rect 23680 41550 23710 41840
rect 22480 41520 23040 41530
rect 23190 41540 23250 41550
rect 23190 41470 23250 41480
rect 23520 41540 23580 41550
rect 23520 41470 23580 41480
rect 23640 41540 23710 41550
rect 23700 41505 23710 41540
rect 23640 41470 23700 41480
rect 23780 41410 23810 41930
rect 23630 40830 23690 40840
rect 23630 40760 23690 40770
rect 17080 40330 17450 40340
rect 1540 40160 1910 40170
rect 555 39820 615 39830
rect 615 39780 960 39820
rect 555 39750 615 39760
rect 10360 39670 10420 39680
rect 10360 39600 10420 39610
rect 15770 39390 15830 39400
rect 615 39350 675 39360
rect 675 39310 960 39350
rect 15770 39320 15830 39330
rect 615 39280 675 39290
rect 9980 38910 10040 38920
rect 9980 38840 10040 38850
rect 14530 38750 15060 38850
rect 675 38730 735 38740
rect 735 38690 970 38730
rect 675 38660 735 38670
rect 3410 38080 3470 38090
rect 3290 38040 3410 38080
rect 3410 38010 3470 38020
rect 14810 38020 14870 38030
rect 14750 37970 14810 38000
rect 14810 37950 14870 37960
rect 15010 37920 15060 38750
rect 15680 38500 15740 38510
rect 15740 38451 15880 38491
rect 15680 38430 15740 38440
rect 14695 37890 14905 37918
rect 14695 37888 14920 37890
rect 14860 37880 14920 37888
rect 14695 37798 14805 37828
rect 14860 37810 14920 37820
rect 3345 37750 3486 37768
rect 3250 37738 3486 37750
rect 3250 37710 3390 37738
rect 14775 37735 14805 37798
rect 14860 37750 14920 37760
rect 14775 37705 14860 37735
rect 14860 37680 14920 37690
rect 3410 37670 3470 37680
rect 15010 37640 15630 37920
rect 15680 37880 15740 37890
rect 15680 37810 15740 37820
rect 15750 37750 15810 37760
rect 15750 37680 15810 37690
rect 3410 37600 3470 37610
rect 1960 37330 2300 37340
rect 1960 36980 2300 36990
rect 7410 37330 7750 37340
rect 7410 36980 7750 36990
rect 10095 36840 10155 36850
rect 9975 36780 10035 36790
rect 9885 36720 9945 36730
rect 9795 36660 9855 36670
rect 9705 36600 9765 36610
rect 9615 36540 9675 36550
rect 9525 36480 9585 36490
rect 9975 36710 10035 36720
rect 9885 36650 9945 36660
rect 9795 36590 9855 36600
rect 9705 36530 9765 36540
rect 9615 36470 9675 36480
rect 9525 36410 9585 36420
rect -100 34950 240 34960
rect -100 34600 240 34610
rect 9555 32660 9585 36410
rect 9645 32750 9675 36470
rect 9735 32840 9765 36530
rect 9825 32930 9855 36590
rect 9915 33020 9945 36650
rect 10005 33110 10035 36710
rect 10095 36770 10155 36780
rect 10185 36780 10245 36790
rect 10095 33200 10125 36770
rect 10185 36710 10245 36720
rect 10275 36720 10335 36730
rect 10185 33290 10215 36710
rect 10275 36650 10335 36660
rect 10365 36660 10425 36670
rect 10275 33380 10305 36650
rect 10365 36590 10425 36600
rect 10455 36600 10515 36610
rect 10365 33470 10395 36590
rect 10455 36530 10515 36540
rect 10545 36540 10605 36550
rect 10455 33560 10485 36530
rect 10545 36470 10605 36480
rect 10635 36480 10695 36490
rect 10545 33650 10575 36470
rect 10635 36410 10695 36420
rect 10635 33740 10665 36410
rect 19540 35030 19910 35040
rect 19540 34650 19910 34660
rect 10620 33730 10680 33740
rect 10620 33660 10680 33670
rect 10530 33640 10590 33650
rect 10530 33570 10590 33580
rect 10440 33550 10500 33560
rect 10440 33480 10500 33490
rect 10350 33460 10410 33470
rect 10350 33390 10410 33400
rect 10260 33370 10320 33380
rect 10260 33300 10320 33310
rect 10170 33280 10230 33290
rect 10170 33210 10230 33220
rect 10080 33190 10140 33200
rect 10080 33120 10140 33130
rect 9990 33100 10050 33110
rect 9990 33030 10050 33040
rect 9900 33010 9960 33020
rect 9900 32940 9960 32950
rect 9810 32920 9870 32930
rect 9810 32850 9870 32860
rect 9720 32830 9780 32840
rect 9720 32760 9780 32770
rect 9630 32740 9690 32750
rect 9630 32670 9690 32680
rect 9540 32650 9600 32660
rect 9540 32580 9600 32590
rect 18840 31560 19200 31570
rect 1090 31540 1430 31550
rect 1090 31190 1430 31200
rect 18840 31190 19200 31200
<< via2 >>
rect -3540 48420 -3480 48480
rect -3540 48140 -3480 48200
rect 23950 48420 24010 48480
rect 23950 48150 24010 48210
rect -3540 47880 -3480 47940
rect 23950 47880 24010 47940
rect -3540 47600 -3480 47660
rect 23950 47610 24010 47670
rect -3550 47330 -3490 47390
rect 23950 47330 24010 47390
rect -3550 47060 -3490 47120
rect 23950 47050 24010 47110
rect -3540 46790 -3480 46850
rect 23950 46790 24010 46850
rect -3550 46520 -3490 46580
rect 23950 46520 24010 46580
rect -3540 46250 -3480 46310
rect 23950 46250 24010 46310
rect -3540 45980 -3480 46040
rect 23950 45970 24010 46030
rect -3540 45700 -3480 45760
rect 23950 45710 24010 45770
rect -3540 45430 -3480 45490
rect 23950 45440 24010 45500
rect -3540 45150 -3480 45210
rect 23950 45170 24010 45230
rect -3540 44880 -3480 44940
rect 23950 44890 24010 44950
rect -3540 44610 -3480 44670
rect 23950 44630 24010 44690
rect -3540 44340 -3480 44400
rect 23950 44350 24010 44410
rect -3540 44070 -3480 44130
rect 23950 44080 24010 44140
rect -3540 43800 -3480 43860
rect 23950 43800 24010 43860
rect -3540 43530 -3480 43590
rect 23960 43530 24020 43590
rect -3540 43260 -3480 43320
rect 23950 43270 24010 43330
rect -3540 42990 -3480 43050
rect 23950 42980 24010 43040
rect -3540 42720 -3480 42780
rect 23950 42720 24010 42780
rect -3540 42410 -3480 42470
rect 23940 42440 24000 42500
rect -5050 41700 -4990 41780
rect -3660 41700 -3580 41780
rect -4790 41540 -4730 41620
rect -3660 41540 -3580 41620
rect -100 40340 240 40680
rect 1540 40340 1910 40680
rect 9260 40340 9630 40680
rect 22480 41530 23040 41680
rect 17080 40340 17450 40680
rect 10360 39610 10420 39670
rect 9980 38850 10040 38910
rect 14860 37820 14920 37880
rect 14860 37690 14920 37750
rect 15680 37820 15740 37880
rect 15750 37690 15810 37750
rect 1960 36990 2300 37330
rect 7410 36990 7750 37330
rect -100 34610 240 34950
rect 19540 34660 19910 35030
rect 1090 31200 1430 31540
rect 18840 31200 19200 31560
<< metal3 >>
rect -5310 41455 -5250 48700
rect -5050 41785 -4990 48700
rect -5060 41780 -4980 41785
rect -5060 41700 -5050 41780
rect -4990 41700 -4980 41780
rect -5060 41695 -4980 41700
rect -5320 41408 -5240 41455
rect -5050 41408 -4990 41695
rect -4790 41625 -4730 48700
rect -3550 48480 -3470 48485
rect -3550 48420 -3540 48480
rect -3480 48420 -3470 48480
rect -3550 48415 -3470 48420
rect 23940 48480 24020 48485
rect 23940 48420 23950 48480
rect 24010 48420 24020 48480
rect 23940 48415 24020 48420
rect 23940 48210 24020 48215
rect -3550 48200 -3470 48205
rect -3550 48140 -3540 48200
rect -3480 48140 -3470 48200
rect 23940 48150 23950 48210
rect 24010 48150 24020 48210
rect 23940 48145 24020 48150
rect -3550 48135 -3470 48140
rect -3550 47940 -3470 47945
rect -3550 47880 -3540 47940
rect -3480 47880 -3470 47940
rect -3550 47875 -3470 47880
rect 23940 47940 24020 47945
rect 23940 47880 23950 47940
rect 24010 47880 24020 47940
rect 23940 47875 24020 47880
rect 23940 47670 24020 47675
rect -3550 47660 -3470 47665
rect -3550 47600 -3540 47660
rect -3480 47600 -3470 47660
rect 23940 47610 23950 47670
rect 24010 47610 24020 47670
rect 23940 47605 24020 47610
rect -3550 47595 -3470 47600
rect -3560 47390 -3480 47395
rect -3560 47330 -3550 47390
rect -3490 47330 -3480 47390
rect -3560 47325 -3480 47330
rect 23940 47390 24020 47395
rect 23940 47330 23950 47390
rect 24010 47330 24020 47390
rect 23940 47325 24020 47330
rect -3560 47120 -3480 47125
rect -3560 47060 -3550 47120
rect -3490 47060 -3480 47120
rect -3560 47055 -3480 47060
rect 23940 47110 24020 47115
rect 23940 47050 23950 47110
rect 24010 47050 24020 47110
rect 23940 47045 24020 47050
rect -3550 46850 -3470 46855
rect -3550 46790 -3540 46850
rect -3480 46790 -3470 46850
rect -3550 46785 -3470 46790
rect 23940 46850 24020 46855
rect 23940 46790 23950 46850
rect 24010 46790 24020 46850
rect 23940 46785 24020 46790
rect -3560 46580 -3480 46585
rect -3560 46520 -3550 46580
rect -3490 46520 -3480 46580
rect -3560 46515 -3480 46520
rect 23940 46580 24020 46585
rect 23940 46520 23950 46580
rect 24010 46520 24020 46580
rect 23940 46515 24020 46520
rect -3550 46310 -3470 46315
rect -3550 46250 -3540 46310
rect -3480 46250 -3470 46310
rect -3550 46245 -3470 46250
rect 23940 46310 24020 46315
rect 23940 46250 23950 46310
rect 24010 46250 24020 46310
rect 23940 46245 24020 46250
rect -3550 46040 -3470 46045
rect -3550 45980 -3540 46040
rect -3480 45980 -3470 46040
rect -3550 45975 -3470 45980
rect 23940 46030 24020 46035
rect 23940 45970 23950 46030
rect 24010 45970 24020 46030
rect 23940 45965 24020 45970
rect 23940 45770 24020 45775
rect -3550 45760 -3470 45765
rect -3550 45700 -3540 45760
rect -3480 45700 -3470 45760
rect 23940 45710 23950 45770
rect 24010 45710 24020 45770
rect 23940 45705 24020 45710
rect -3550 45695 -3470 45700
rect 23940 45500 24020 45505
rect -3550 45490 -3470 45495
rect -3550 45430 -3540 45490
rect -3480 45430 -3470 45490
rect 23940 45440 23950 45500
rect 24010 45440 24020 45500
rect 23940 45435 24020 45440
rect -3550 45425 -3470 45430
rect 23940 45230 24020 45235
rect -3550 45210 -3470 45215
rect -3550 45150 -3540 45210
rect -3480 45150 -3470 45210
rect 23940 45170 23950 45230
rect 24010 45170 24020 45230
rect 23940 45165 24020 45170
rect -3550 45145 -3470 45150
rect 23940 44950 24020 44955
rect -3550 44940 -3470 44945
rect -3550 44880 -3540 44940
rect -3480 44880 -3470 44940
rect 23940 44890 23950 44950
rect 24010 44890 24020 44950
rect 23940 44885 24020 44890
rect -3550 44875 -3470 44880
rect 23940 44690 24020 44695
rect -3550 44670 -3470 44675
rect -3550 44610 -3540 44670
rect -3480 44610 -3470 44670
rect 23940 44630 23950 44690
rect 24010 44630 24020 44690
rect 23940 44625 24020 44630
rect -3550 44605 -3470 44610
rect 23940 44410 24020 44415
rect -3550 44400 -3470 44405
rect -3550 44340 -3540 44400
rect -3480 44340 -3470 44400
rect 23940 44350 23950 44410
rect 24010 44350 24020 44410
rect 23940 44345 24020 44350
rect -3550 44335 -3470 44340
rect 23940 44140 24020 44145
rect -3550 44130 -3470 44135
rect -3550 44070 -3540 44130
rect -3480 44070 -3470 44130
rect 23940 44080 23950 44140
rect 24010 44080 24020 44140
rect 23940 44075 24020 44080
rect -3550 44065 -3470 44070
rect -3550 43860 -3470 43865
rect -3550 43800 -3540 43860
rect -3480 43800 -3470 43860
rect -3550 43795 -3470 43800
rect 23940 43860 24020 43865
rect 23940 43800 23950 43860
rect 24010 43800 24020 43860
rect 23940 43795 24020 43800
rect -3550 43590 -3470 43595
rect -3550 43530 -3540 43590
rect -3480 43530 -3470 43590
rect -3550 43525 -3470 43530
rect 23950 43590 24030 43595
rect 23950 43530 23960 43590
rect 24020 43530 24030 43590
rect 23950 43525 24030 43530
rect 23940 43330 24020 43335
rect -3550 43320 -3470 43325
rect -3550 43260 -3540 43320
rect -3480 43260 -3470 43320
rect 23940 43270 23950 43330
rect 24010 43270 24020 43330
rect 23940 43265 24020 43270
rect -3550 43255 -3470 43260
rect -3550 43050 -3470 43055
rect -3550 42990 -3540 43050
rect -3480 42990 -3470 43050
rect -3550 42985 -3470 42990
rect 23940 43040 24020 43045
rect 23940 42980 23950 43040
rect 24010 42980 24020 43040
rect 23940 42975 24020 42980
rect -3550 42780 -3470 42785
rect -3550 42720 -3540 42780
rect -3480 42720 -3470 42780
rect -3550 42715 -3470 42720
rect 23940 42780 24020 42785
rect 23940 42720 23950 42780
rect 24010 42720 24020 42780
rect 23940 42715 24020 42720
rect 23930 42500 24010 42505
rect -3550 42470 -3470 42475
rect -3550 42410 -3540 42470
rect -3480 42410 -3470 42470
rect 23930 42440 23940 42500
rect 24000 42440 24010 42500
rect 23930 42435 24010 42440
rect -3550 42405 -3470 42410
rect 21970 41830 25340 41910
rect -3670 41780 -3570 41785
rect 21970 41780 22050 41830
rect -3670 41700 -3660 41780
rect -3580 41700 22050 41780
rect -3670 41695 -3570 41700
rect 22470 41680 23050 41685
rect -4800 41620 -4720 41625
rect -4800 41540 -4790 41620
rect -4730 41540 -4720 41620
rect -4800 41535 -4720 41540
rect -3670 41620 -3570 41625
rect -3670 41540 -3660 41620
rect -3580 41540 22060 41620
rect -3670 41535 -3570 41540
rect -4790 41408 -4730 41535
rect 21980 41310 22060 41540
rect 22470 41530 22480 41680
rect 23040 41530 23050 41680
rect 22470 41525 23050 41530
rect 21980 41230 25077 41310
rect -110 40680 250 40685
rect 1530 40680 1920 40685
rect 9250 40680 9640 40685
rect 17070 40680 17460 40685
rect -110 40340 -100 40680
rect 240 40340 1540 40680
rect 1910 40340 9260 40680
rect 9630 40340 17080 40680
rect 17450 40340 19170 40680
rect 19540 40340 22390 40680
rect -110 40335 250 40340
rect 1530 40335 1920 40340
rect 9250 40335 9640 40340
rect 17070 40335 17460 40340
rect 9670 39810 10690 40020
rect 9670 39460 10240 39810
rect 10340 39680 10440 39690
rect 10340 39610 10360 39680
rect 10430 39610 10440 39680
rect 10340 39590 10440 39610
rect 10570 39460 10690 39810
rect 9670 39060 10690 39460
rect 9670 38710 9840 39060
rect 9950 38920 10060 38930
rect 9950 38850 9970 38920
rect 10040 38850 10060 38920
rect 9950 38830 10060 38850
rect 10170 38710 10690 39060
rect 1950 37330 2310 37335
rect 7400 37330 7760 37335
rect 9670 37330 10690 38710
rect 14850 37880 14930 37885
rect 15670 37880 15750 37885
rect 14850 37820 14860 37880
rect 14920 37820 15680 37880
rect 15740 37820 15750 37880
rect 14850 37815 14930 37820
rect 15670 37815 15750 37820
rect 14850 37750 14930 37755
rect 15740 37750 15820 37755
rect 14850 37690 14860 37750
rect 14920 37690 15750 37750
rect 15810 37690 15820 37750
rect 14850 37685 14930 37690
rect 15740 37685 15820 37690
rect 550 36990 560 37330
rect 900 36990 1960 37330
rect 2300 36990 7410 37330
rect 7750 36990 22480 37330
rect 23040 36990 23050 37330
rect 1950 36985 2310 36990
rect 7400 36985 7760 36990
rect -5310 36170 -5250 36322
rect -5050 36240 -4990 36322
rect -4790 36240 -4730 36322
rect -110 34950 250 34955
rect -110 34610 -100 34950
rect 240 34610 250 34950
rect -110 34605 250 34610
rect 3170 32130 3990 32410
rect 3170 31880 3470 32130
rect 3690 31880 3990 32130
rect 1080 31540 1440 31550
rect 1080 31200 1090 31540
rect 1430 31200 1440 31540
rect 1080 30270 1440 31200
rect 3170 30470 3990 31880
rect 9670 30480 10690 36990
rect 25017 35840 25077 41230
rect 25277 36200 25337 41830
rect 25537 36130 25597 48690
rect 19530 35030 19920 35035
rect 19530 34660 19540 35030
rect 19910 34660 19920 35030
rect 19530 34655 19920 34660
rect 16310 32130 17130 32410
rect 16310 31880 16590 32130
rect 16820 31880 17130 32130
rect 16310 30480 17130 31880
rect 18830 31560 19210 31565
rect 18830 31200 18840 31560
rect 19200 31200 19210 31560
rect 18830 31195 19210 31200
rect 9670 30470 17130 30480
rect 3170 30270 17130 30470
rect 18850 30270 19210 31195
rect 1080 29910 19210 30270
rect 3170 29760 17130 29910
rect 3170 29750 12210 29760
rect 16310 29750 17130 29760
rect 8080 28870 12210 29750
<< via3 >>
rect 22480 41530 23040 41680
rect -100 40340 240 40680
rect 19170 40340 19540 40680
rect 10360 39670 10430 39680
rect 10360 39610 10420 39670
rect 10420 39610 10430 39670
rect 9970 38910 10040 38920
rect 9970 38850 9980 38910
rect 9980 38850 10040 38910
rect 560 36990 900 37330
rect 22480 36990 23040 37330
rect -100 34610 240 34950
rect 1090 31200 1430 31540
rect 19540 34660 19910 35030
<< metal4 >>
rect -92 47215 228 49050
rect 568 47290 888 49040
rect -100 41431 240 42870
rect 560 42141 900 42870
rect 559 41799 901 42141
rect -101 41089 241 41431
rect -100 40681 240 41089
rect -101 40680 241 40681
rect -101 40340 -100 40680
rect 240 40340 241 40680
rect -101 40339 241 40340
rect -100 34951 240 40339
rect 560 37331 900 41799
rect 22480 41681 23040 41720
rect 22479 41680 23041 41681
rect 22479 41530 22480 41680
rect 23040 41530 23041 41680
rect 22479 41529 23041 41530
rect 19169 40680 19541 40681
rect 19169 40340 19170 40680
rect 19540 40340 19541 40680
rect 19169 40339 19541 40340
rect 10359 39680 10431 39681
rect 10359 39610 10360 39680
rect 10430 39610 10431 39680
rect 10359 39609 10431 39610
rect 9969 38920 10041 38921
rect 9969 38850 9970 38920
rect 10040 38890 10041 38920
rect 10040 38850 10050 38890
rect 9969 38849 10050 38850
rect 559 37330 901 37331
rect 559 36990 560 37330
rect 900 36990 901 37330
rect 559 36989 901 36990
rect -101 34950 241 34951
rect -101 34610 -100 34950
rect 240 34610 241 34950
rect -101 34609 241 34610
rect -100 34580 240 34609
rect 560 32751 900 36989
rect 559 31541 901 32751
rect 3539 31979 3621 32061
rect 559 31540 1431 31541
rect 559 31200 1090 31540
rect 1430 31200 1431 31540
rect 559 31199 1431 31200
rect 3550 30100 3610 31979
rect 9990 30100 10050 38849
rect 3550 30040 10050 30100
rect 9990 29140 10050 30040
rect 8170 29080 10050 29140
rect 10370 30100 10430 39609
rect 19170 35031 19540 40339
rect 22480 37331 23040 41529
rect 22479 37330 23041 37331
rect 22479 36990 22480 37330
rect 23040 36990 23041 37330
rect 22479 36989 23041 36990
rect 19170 35030 19911 35031
rect 19170 34660 19540 35030
rect 19910 34660 19911 35030
rect 19539 34659 19911 34660
rect 16680 32051 16740 32065
rect 16669 31969 16751 32051
rect 16680 30100 16740 31969
rect 10370 30040 16740 30100
rect 10370 29140 10430 30040
rect 10370 29080 12117 29140
rect 8170 28860 8230 29080
rect 12057 28870 12117 29080
use break_before_make  break_before_make_0 ~/Desktop/SAR_ADC_12bit/break_before_make/layout
timestamp 1713906110
transform 1 0 -7051 0 1 29930
box 1725 6360 6167 11600
use DAC_and_SW  DAC_and_SW_0
timestamp 1713606823
transform -1 0 25087 0 1 4500
box -520 0 15040 31800
use DAC_and_SW  DAC_and_SW_1
timestamp 1713606823
transform 1 0 -4800 0 1 4500
box -520 0 15040 31800
use latched_comparator  latched_comparator_0 ~/Desktop/SAR_ADC_12bit/layout/../latched_comparator/layout
timestamp 1712061640
transform -1 0 8780 0 1 39170
box 5450 -1740 7860 1100
use offset_calibration  offset_calibration_0 ~/Desktop/SAR_ADC_12bit/layout/../offset_calibration/layout
timestamp 1712002773
transform 1 0 12181 0 1 38781
box 3610 -1900 11750 2900
use preamplifier  preamplifier_0 ~/Desktop/SAR_ADC_12bit/layout/../preamplifier/layout
timestamp 1711972782
transform -1 0 11136 0 1 30538
box -3630 6580 7680 9930
use state_machine  state_machine_0 ~/Desktop/SAR_ADC_12bit/layout/../state_machine/layout
timestamp 1713020991
transform 1 0 -4300 0 1 40495
box 480 1360 28477 8022
<< labels >>
rlabel metal3 -5310 48640 -5250 48700 1 VIN_P
port 16 n
rlabel metal3 -5050 48640 -4990 48700 1 VREF
port 17 n
rlabel metal3 -4790 48640 -4730 48700 1 VCM
port 18 n
rlabel metal3 25537 48630 25597 48690 1 VIN_N
port 19 n
rlabel metal4 -80 48760 200 49020 1 VDD
port 20 n
rlabel metal4 600 48770 880 49030 1 VSS
port 21 n
rlabel metal2 -2990 48260 -2940 48440 1 CLK_DATA
port 1 n
rlabel metal2 -1150 48280 -1100 48460 1 DATA[0]
port 2 n
rlabel metal2 410 48290 460 48470 1 DATA[1]
port 3 n
rlabel metal2 2250 48290 2300 48470 1 DATA[2]
port 4 n
rlabel metal2 4000 48290 4050 48470 1 DATA[3]
port 5 n
rlabel metal2 5750 48290 5800 48470 1 DATA[4]
port 6 n
rlabel metal2 7500 48290 7550 48470 1 DATA[5]
port 7 n
rlabel metal2 9240 48280 9290 48460 1 DEBUG_OUT
port 8 n
rlabel metal2 10990 48280 11040 48460 1 RST_Z
port 9 n
rlabel metal2 14490 48240 14540 48420 1 START
port 10 n
rlabel metal2 16240 48240 16290 48420 1 EN_OFFSET_CAL
port 11 n
rlabel metal2 17990 48290 18040 48470 1 DEBUG_MUX[0]
port 12 n
rlabel metal2 19730 48250 19780 48430 1 DEBUG_MUX[1]
port 13 n
rlabel metal2 21480 48270 21530 48450 1 DEBUG_MUX[2]
port 14 n
rlabel metal2 23230 48280 23280 48460 1 DEBUG_MUX[3]
port 15 n
rlabel metal2 12740 48260 12790 48440 1 CLK
port 22 n
rlabel metal2 8960 8890 8980 8960 1 C10_P_btm
rlabel metal2 11310 8870 11330 8940 1 C10_N_btm
rlabel metal2 9050 11080 9070 11180 1 C9_P_btm
rlabel metal2 11220 11090 11240 11190 1 C9_N_btm
rlabel metal2 9140 12890 9160 12980 1 C8_P_btm
rlabel metal2 11120 12900 11140 12990 1 C8_N_btm
rlabel metal2 9230 14000 9250 14120 1 C7_P_btm
rlabel metal2 11040 14030 11060 14150 1 C7_N_btm
rlabel metal2 9320 14730 9340 14810 1 C6_P_btm
rlabel metal2 10950 14740 10970 14820 1 C6_N_btm
rlabel metal2 9410 15120 9430 15200 1 C5_P_btm
rlabel metal2 10860 15100 10880 15180 1 C5_N_btm
rlabel metal2 9500 15830 9520 15910 1 C4_P_btm
rlabel metal2 10760 15830 10780 15910 1 C4_N_btm
rlabel metal2 9580 16300 9600 16360 1 C2_P_btm
rlabel metal2 10680 16230 10700 16290 1 C2_N_btm
rlabel metal2 9680 16590 9700 16660 1 C0_dummy_P_btm
rlabel metal2 10590 16590 10610 16660 1 C0_dummy_N_btm
rlabel metal2 9770 16960 9790 17020 1 C0_P_btm
rlabel metal2 10500 16970 10520 17030 1 C0_N_btm
rlabel metal2 9860 17320 9880 17380 1 C1_P_btm
rlabel metal2 10410 17330 10430 17390 1 C1_N_btm
rlabel metal2 9950 17690 9970 17750 1 C3_P_btm
rlabel metal2 10320 17700 10340 17760 1 C3_N_btm
rlabel metal4 8180 28890 8220 28910 1 VDAC_P
rlabel metal4 12070 28890 12110 28910 1 VDAC_N
rlabel metal2 3350 38050 3380 38070 1 VDAC_Pi
rlabel metal2 3340 37720 3370 37740 1 VDAC_Ni
rlabel metal2 930 38700 960 38720 1 EN_COMP
rlabel metal2 920 39320 950 39340 1 COMP_N
rlabel metal2 910 39790 940 39810 1 COMP_P
rlabel metal3 15640 37700 15660 37730 1 CAL_N
rlabel metal3 15640 37830 15660 37860 1 CAL_P
rlabel metal2 -3248 41854 -3224 41880 1 SMPL
rlabel metal2 -3744 48428 -3716 48444 1 SMPL_ON_P
rlabel metal2 24104 48446 24132 48462 1 SMPL_ON_N
rlabel metal2 1166 34386 1194 34402 1 EN_VIN_BSTR_P
rlabel metal2 19090 34368 19120 34400 1 EN_VIN_BSTR_N
<< end >>
