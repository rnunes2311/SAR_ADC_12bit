** sch_path: /Users/ricardonunes/Desktop/SAR_ADC_12bit/simulations/top_level_differential_sim.sch

* Skywater 130 nm PDK models
.lib /opt/pdk/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

* Models for standard digital cells
.include /opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

* C extraction spice netlist for CDAC
*.include /Users/ricardonunes/Desktop/SAR_ADC_12bit/simulations/../layout/subcells/CDAC/CDAC_mim_12bit_flat.spice

* Spice netlist for state machine generated by openlane
*.include /Users/ricardonunes/Desktop/SAR_ADC_12bit/simulations/../layout/subcells/state_machine/state_machine_openlane_generated.spice

* C or RC extraction of the SAR ADC
.include /Users/ricardonunes/Desktop/SAR_ADC_12bit/simulations/../layout/SAR_ADC_12bit_flat.spice

**.subckt top_level_differential_sim
V1 VDD VSS {VDD}
.save i(v1)
V2 net1 VSS {VCM}
.save i(v2)
V3 net2 VSS {VREF}
.save i(v3)
V4 VSS GND 0
V7 START VSS pulse(0 1.8 20n 1n 1n 100n 1u)
V8 RST_Z VSS pwl(0 0 10n 0 10.1n 1.8)
V5 net4 VSS pwl(0.000u 0.6 1u 0.6 1.000u 0.4000 2u 0.4000 2.001u 0.8000 3u 0.8000 3.001u 0.9599 4u 0.9599 4.001u 0.2401 5u 0.2401
+ 5.001u 0.0186 6u 0.0186 6.001u 1.1814 7u 1.1814)
x1 VDD VCM VSS VREF VIN_P VIN_N RST_Z CLK_DATA DATA[5] DATA[4] DATA[3] DATA[2] DATA[1] DATA[0] START EN_OFFSET_CAL CLK VREF_GND
+ SINGLE_ENDED SAR_ADC_12bit
R1 net1 VCM 500 m=1
V9 CLK VSS pulse(0 1.8 0 1n 1n 40n 50n)
V6 net5 VSS pwl(0.000u 0.6 1u 0.6 1.000u 0.8000 2u 0.8000 2.001u 0.4000 3u 0.4000 3.001u 0.2401 4u 0.2401 4.001u 0.9599 5u 0.9599
+ 5.001u 1.1814 6u 1.1814 6.001u 0.0186 7u 0.0186)
V10 net3 VSS {VREF_GND}
.save i(v10)
R6 net2 VREF 500 m=1
R7 net3 VREF_GND 500 m=1
R8 net4 VIN_P 500 m=1
R9 net5 VIN_N 500 m=1
V11 EN_OFFSET_CAL VSS pwl(0 0 3u 0 3.001u 1.8)
V12 SINGLE_ENDED VSS 0
**** begin user architecture code


* Supply, common mode and reference voltage
.param VDD = 1.8
.param VREF = 1.2
.param VREF_GND = 0
.param VCM = 0.6

.option temp = 27

*.save all

* Control signals
.save start rst_z clk en_offset_cal

* Input signals
.save vin_p vin_n

* Reference, supply
.save vref vref_gnd vcm vdd

* Output signals
.save clk_data data[5] data[4] data[3] data[2] data[1] data[0]

* Internal signals
.save x1.vdac_p x1.vdac_n x1.vdac_pi x1.vdac_ni x1.smpl x1.en_comp x1.comp_p x1.comp_n x1.cal_p x1.cal_n
.save x1.en_vin_bstr_p x1.en_vin_bstr_n
.save x1.c10_p_btm x1.c9_p_btm x1.c8_p_btm x1.c7_p_btm x1.c6_p_btm x1.c5_p_btm x1.c4_p_btm x1.c3_p_btm x1.c2_p_btm x1.c1_p_btm x1.c0_p_btm x1.C0_dummy_p_btm
.save x1.c10_n_btm x1.c9_n_btm x1.c8_n_btm x1.c7_n_btm x1.c6_n_btm x1.c5_n_btm x1.c4_n_btm x1.c3_n_btm x1.c2_n_btm x1.c1_n_btm x1.c0_n_btm x1.C0_dummy_n_btm

.option GMIN=1e-12 reltol=1e-5
.control
		set ngbehavior=hsa
          		set skywaterpdk
          		set ng_nomodcheck
          		set num_threads=4
          		option noinit
          		option klu
		tran 10n 7u
		write top_level_differential_sim.raw
.endc


**** end user architecture code
**.ends
.end
