* SPICE3 file created from SAR_ADC_12bit_flat.ext - technology: sky130A
* Changed subckt name from SAR_ADC_12bit_flat to SAR_ADC_12bit

.subckt SAR_ADC_12bit VDD VCM VSS VREF VIN_P VIN_N RST_Z CLK_DATA DATA[5] DATA[4] DATA[3] DATA[2] DATA[1] DATA[0] START
+ EN_OFFSET_CAL CLK VREF_GND SINGLE_ENDED
X0 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1 a_13076_44458# a_13259_45724# a_13296_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VDD a_2324_44458# a_949_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4 VSS a_12427_45724# a_10490_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X9 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=361.2627 ps=3.22652k w=10 l=10
X10 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X11 VDD a_2903_42308# a_3080_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X12 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X13 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X14 VDD a_12861_44030# a_17829_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VSS a_1209_43370# a_n1557_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X16 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X17 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X18 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X19 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X20 a_16237_45028# a_16147_45260# a_16019_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 a_2075_43172# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VDD a_n755_45592# a_1176_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X23 a_6756_44260# a_5937_45572# a_6453_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X24 a_n1533_42852# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X25 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X26 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X27 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X28 a_15868_43402# a_15681_43442# a_15781_43660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X29 a_8103_44636# a_8375_44464# a_8333_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X31 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X32 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X33 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X34 VSS a_16327_47482# a_16377_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X35 a_2437_43646# a_n443_46116# a_2437_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X36 a_5088_37509# VSS VDAC_Ni VDD sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X37 a_n2810_45028# a_n2840_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X38 a_2113_38308# VDAC_Ni a_2112_39137# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X39 VDD a_3626_43646# a_19647_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X40 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X41 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X42 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X43 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X44 VSS a_10334_44484# a_10440_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X45 a_1576_42282# a_1755_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X46 a_10933_46660# a_10554_47026# a_10861_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X47 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X48 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X49 a_16867_43762# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X50 a_14021_43940# a_13483_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X51 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X52 VREF a_21076_30879# C8_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X53 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X54 VSS a_n2946_37690# a_n3565_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X55 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X56 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X57 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X58 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X59 a_n913_45002# a_1307_43914# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X60 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X61 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X62 a_n2840_43370# a_n2661_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X63 a_3457_43396# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X64 a_1343_38525# a_1177_38525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X65 VSS a_9672_43914# a_2107_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X66 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X67 a_14180_46482# a_14035_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X68 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X69 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X70 VSS C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X71 a_n1059_45260# a_17499_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X72 VSS a_18989_43940# a_19006_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X73 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X74 a_20749_43396# a_12549_44172# a_743_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X75 a_n2104_42282# a_n1925_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X76 VSS a_10695_43548# a_10057_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X77 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X78 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X79 VDD a_3877_44458# a_2382_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X80 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X81 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X82 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X83 VSS a_n4334_39616# a_n4064_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X84 a_n1699_44726# a_n1917_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X85 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X86 VDD a_12883_44458# a_n2293_43922# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X87 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X88 a_9241_45822# a_5066_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X89 a_11909_44484# a_3232_43370# a_11827_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X90 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X91 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X92 a_835_46155# a_584_46384# a_376_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X93 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X94 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X95 a_5210_46155# a_5164_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X96 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X97 VDD a_n3690_39392# a_n3420_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X98 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X99 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X100 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X101 VDD a_167_45260# a_1609_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X102 VSS a_526_44458# a_3363_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X103 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X104 a_19268_43646# a_19319_43548# a_19095_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X105 VSS a_22959_44484# a_19237_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X106 VDAC_P C2_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X107 a_n2216_39072# a_n2312_39304# a_n2302_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X108 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X109 VDD a_1177_38525# a_1343_38525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X110 a_19987_42826# a_10193_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X111 a_6151_47436# a_14311_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X112 a_8145_46902# a_7927_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X113 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X114 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X115 a_14275_46494# a_13925_46122# a_14180_46482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X116 a_20512_43084# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X117 a_14539_43914# a_17701_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X118 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X119 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X120 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X121 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X122 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X123 a_6298_44484# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X124 a_644_44056# a_626_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X125 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X126 a_10949_43914# a_12429_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.28 ps=2.56 w=1 l=0.15
X127 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X128 VSS a_n2302_39866# a_n4209_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X129 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X130 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X131 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X132 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X133 VDD a_3699_46634# a_3686_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X134 VSS a_21811_47423# a_20916_46384# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X135 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X136 a_5691_45260# a_5111_44636# a_5837_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X137 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X138 a_18249_42858# a_18083_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X139 a_8035_47026# a_7411_46660# a_7927_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X140 VDD a_1307_43914# a_1241_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X141 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X142 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X143 VDD a_104_43370# a_n971_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X144 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X145 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X146 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X147 VSS a_n3565_39590# a_n3607_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X148 a_n1331_43914# a_n1549_44318# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X149 VDD a_n2833_47464# CLK_DATA VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X150 a_3363_44484# a_1823_45246# a_3232_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X151 VCM a_4958_30871# C9_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X152 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X153 VSS a_12281_43396# a_12563_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X154 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X155 VSS a_22400_42852# a_22780_40081# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X156 VSS a_18780_47178# a_13661_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X157 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X158 a_n4318_39768# a_n2840_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X159 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X160 DATA[5] a_11459_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X161 a_15004_44636# a_11691_44458# a_15146_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X162 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X163 VDD a_8049_45260# a_22959_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X164 a_7230_45938# a_6472_45840# a_6667_45809# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X165 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X166 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X167 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X168 a_8746_45002# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X169 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X170 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X171 a_n984_44318# a_n1899_43946# a_n1331_43914# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X172 a_n4064_39616# a_n4334_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X173 a_17124_42282# a_17303_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X174 a_16223_45938# a_15599_45572# a_16115_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X175 a_n809_44244# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X176 VSS a_3065_45002# a_2680_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X177 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X178 a_5193_42852# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X179 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X180 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X181 VDD a_6969_46634# a_6999_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X182 VDD a_10623_46897# a_10554_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X183 a_16137_43396# a_15781_43660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X184 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X185 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X186 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X187 VDD a_n2472_46634# a_n2442_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X188 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X189 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X190 VDD a_4185_45028# a_22959_45036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X191 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X192 a_15225_45822# a_15037_45618# a_15143_45578# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X193 VSS a_3537_45260# a_4640_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X194 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X195 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X196 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X197 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X198 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X199 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X200 VSS C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X201 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X202 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X203 a_n2012_43396# a_n2129_43609# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X204 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X205 VDD a_n13_43084# a_n1853_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X206 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X207 a_5068_46348# a_n1151_42308# a_5210_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X208 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X209 a_873_42968# a_685_42968# a_791_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X210 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X211 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X212 VDD a_22485_44484# a_20974_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X213 a_17730_32519# a_22591_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X214 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X215 a_n1021_46688# a_n1151_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X216 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X217 VSS a_11599_46634# a_11735_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X218 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X219 a_13163_45724# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.14075 ps=1.325 w=0.42 l=0.15
X220 C9_P_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X221 a_n2012_44484# a_n2129_44697# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X222 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X223 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X224 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X225 a_8487_44056# a_4223_44672# a_8415_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X226 a_13940_44484# a_13556_45296# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X227 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X228 VSS a_1414_42308# a_1525_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X229 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X230 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X231 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X232 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X233 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X234 a_16434_46660# a_16388_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X235 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X236 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X237 a_3315_47570# a_n1151_42308# a_2952_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X238 a_2680_45002# a_1823_45246# a_2903_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X239 a_1307_43914# a_2779_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X240 VSS a_n1630_35242# a_18194_35068# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X241 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X242 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X243 a_22731_47423# SMPL_ON_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X244 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X245 VDD a_1307_43914# a_3681_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X246 a_n863_45724# a_1667_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X247 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X248 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X249 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X250 a_22521_40599# COMP_P VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X251 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X252 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X253 VDD a_11459_47204# DATA[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X254 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X255 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X256 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X257 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X258 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X259 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=218.18214 ps=2.11206k w=0.55 l=0.59
X260 a_n4209_38216# a_n2302_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X261 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X262 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X263 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X264 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X265 a_10467_46802# a_11599_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X266 VDD a_13747_46662# a_19862_44208# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X267 a_n2946_39866# a_n2956_39768# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X268 a_n1013_45572# a_n1079_45724# a_n1099_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X269 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X270 VSS a_15279_43071# a_14579_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X271 DATA[3] a_7227_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X272 a_7584_44260# a_7542_44172# a_7281_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X273 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X274 VSS a_8049_45260# a_22959_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X275 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X276 a_n97_42460# a_19700_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X277 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X278 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X279 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X280 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X281 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X282 VDAC_P C2_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X283 VDD a_19647_42308# a_13258_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X284 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X285 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X286 a_3754_39466# a_7754_39300# VSS sky130_fd_pr__res_high_po_0p35 l=18
X287 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X288 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X289 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X290 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X291 VDD a_16751_45260# a_6171_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X292 VSS a_2952_47436# a_2747_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X293 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X294 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X295 a_18326_43940# a_18079_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X296 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X297 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X298 VDAC_N C0_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X299 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X300 a_9248_44260# a_8270_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X301 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X302 a_3503_45724# a_3775_45552# a_3733_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X303 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X304 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X305 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X306 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X307 a_n2017_45002# a_19987_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X308 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X309 a_288_46660# a_171_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X310 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X311 VDD a_196_42282# a_n3674_37592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X312 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X313 a_10037_46155# a_9804_47204# a_9823_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X314 a_20075_46420# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X315 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X316 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X317 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X318 a_n4064_39072# a_n4334_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X319 a_1149_42558# a_961_42354# a_1067_42314# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X320 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X321 VSS a_14513_46634# a_14447_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X322 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X323 a_13569_47204# a_13381_47204# a_13487_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X324 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X325 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X326 VDD a_14840_46494# a_15015_46420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X327 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X328 C6_P_btm a_n3565_39304# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=0.35
X329 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X330 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X331 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X332 a_14537_43396# a_14358_43442# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X333 VDD a_14955_47212# a_10227_46804# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X334 a_n3565_39590# a_n2946_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X335 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X336 VDD a_7754_40130# a_11206_38545# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X337 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X338 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X339 a_n901_43156# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X340 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X341 a_17668_45572# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X342 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X343 a_7309_43172# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X344 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X345 a_15493_43396# a_14955_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X346 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X347 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X348 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X349 VDD a_1138_42852# a_1337_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X350 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X351 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X352 a_1427_43646# a_1568_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X353 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X354 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X355 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X356 a_18184_42460# a_15743_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X357 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X358 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X359 VDD a_13351_46090# a_10903_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X360 VDD a_9290_44172# a_10949_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X361 a_8379_46155# a_8128_46384# a_7920_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X362 VSS a_3483_46348# a_17325_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X363 a_18310_42308# a_10193_42453# a_18220_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X364 VSS a_11823_42460# a_14358_43442# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X365 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X366 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X367 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X368 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X369 VDD a_n2288_47178# a_n2312_40392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X370 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X371 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X372 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X373 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X374 a_17719_45144# a_16375_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X375 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X376 VDD a_5891_43370# a_5147_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X377 a_22609_38406# a_22469_39537# CAL_N VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X378 a_7287_43370# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X379 a_11173_44260# a_2063_45854# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X380 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X381 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X382 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X383 a_11897_42308# a_11823_42460# a_11551_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X384 a_19466_46812# a_19778_44110# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X385 a_n3565_38502# a_n2946_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X386 a_9049_44484# a_8701_44490# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X387 VDD a_12861_44030# a_13759_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X388 VDD a_16588_47582# a_16763_47508# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X389 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X390 a_9396_43370# a_4883_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X391 C0_P_btm a_n784_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X392 a_n1736_42282# a_n1557_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X393 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X394 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X395 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X396 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X397 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X398 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X399 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X400 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X401 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X402 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X403 VDD a_14113_42308# a_16522_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X404 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X405 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X406 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X407 a_10651_43940# a_3090_45724# a_10555_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X408 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X409 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X410 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X411 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X412 VDD a_8667_46634# a_n237_47217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X413 a_7499_43078# a_10083_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X414 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X415 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X416 a_6123_31319# a_7227_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X417 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X418 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X419 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X420 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X421 VSS a_n755_45592# a_1145_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X422 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X423 C7_P_btm a_5534_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X424 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X425 VSS a_n4064_37984# a_n2302_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X426 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X427 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X428 VDD a_1239_39587# COMP_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X429 a_n3674_38680# a_n2840_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X430 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X431 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X432 a_3581_42558# a_3539_42460# a_3497_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X433 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X434 VSS a_5907_45546# a_5937_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X435 a_18783_43370# a_15743_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X436 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X437 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X438 VSS a_1799_45572# a_1983_46706# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X439 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X440 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X441 VDD a_22959_46660# a_21076_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X442 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X443 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X444 VDD a_1736_39043# a_1239_39043# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X445 a_13467_32519# a_21487_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X446 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X447 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X448 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X449 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X450 a_2864_46660# a_2747_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X451 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X452 a_8199_44636# a_10355_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X453 a_14403_45348# a_13259_45724# a_14309_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X454 a_556_44484# a_742_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X455 VSS a_15433_44458# a_15367_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X456 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X457 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X458 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X459 a_n1630_35242# a_564_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X460 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X461 a_n2840_43370# a_n2661_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X462 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X463 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X464 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X465 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X466 VSS a_13747_46662# a_13693_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X467 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X468 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X469 a_18245_44484# a_17767_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X470 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X471 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X472 a_13113_42826# a_12895_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X473 a_16855_43396# a_16409_43396# a_16759_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X474 a_19741_43940# a_19862_44208# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X475 a_n1079_45724# a_n755_45592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X476 VSS a_22365_46825# a_20202_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X477 a_19386_47436# a_19321_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X478 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X479 VSS a_526_44458# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X480 a_1176_45822# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X481 a_13887_32519# a_22223_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X482 a_n89_47570# a_n237_47217# a_n452_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X483 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X484 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=10.615 ps=76.96 w=3.75 l=15
X485 a_10341_43396# a_9803_43646# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X486 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X487 a_5111_42852# a_4905_42826# a_5193_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X488 VDD a_n4209_38502# a_n4334_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X489 a_5437_45600# a_n881_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X490 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X491 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X492 a_18953_45572# a_18909_45814# a_18787_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X493 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X494 a_n3607_39616# a_n3674_39768# a_n3690_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X495 VDD a_3429_45260# a_3316_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X496 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X497 VDD a_4791_45118# a_6165_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X498 a_4842_47570# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X499 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X500 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X501 a_1337_46116# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X502 a_n2661_42834# a_10809_44734# a_12189_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X503 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X504 VSS C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X505 a_11136_45572# a_11322_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X506 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X507 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X508 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X509 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X510 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X511 VREF_GND a_n3420_39072# C6_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X512 a_n3565_37414# a_n2946_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X513 VSS a_10249_46116# a_11186_47026# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X514 a_16655_46660# a_n743_46660# a_16292_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X515 a_n1991_46122# a_n2157_46122# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X516 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X517 VDD a_1576_42282# a_1606_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X518 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X519 VSS C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X520 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X521 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X522 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X523 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X524 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X525 a_2075_43172# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X526 a_5159_47243# a_n443_46116# a_4700_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X527 VSS a_5891_43370# a_8375_44464# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X528 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X529 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X530 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X531 VSS a_14539_43914# a_14485_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X532 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X533 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X534 VDD a_13076_44458# a_12883_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X535 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X536 VDD en_comp a_1177_38525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X537 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X538 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X539 C0_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X540 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X541 a_15297_45822# a_11823_42460# a_15225_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X542 a_8103_44636# a_8199_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X543 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X544 a_1423_45028# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X545 a_n1899_43946# a_n2065_43946# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X546 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X547 a_18479_47436# a_20075_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X548 a_2382_45260# a_3877_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X549 a_6765_43638# a_6547_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X550 a_n2293_43922# a_12741_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X551 a_945_42968# a_n1059_45260# a_873_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X552 a_n3565_38216# a_n2946_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X553 VDD a_n3690_39392# a_n3420_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X554 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X555 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X556 VDD a_3785_47178# a_3815_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X557 VDD a_14084_46812# a_14035_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X558 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X559 a_765_45546# a_12549_44172# a_17829_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X560 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X561 VDD a_20974_43370# a_20556_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X562 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X563 VSS a_15051_42282# a_11823_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X564 a_14275_46494# a_13759_46122# a_14180_46482# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X565 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X566 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X567 a_17517_44484# a_16979_44734# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X568 a_1609_45822# a_n443_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X569 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X570 VDD a_4915_47217# a_12891_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X571 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X572 a_20679_44626# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X573 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X574 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X575 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X576 a_13921_42308# a_13259_45724# a_13575_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X577 VSS a_1423_45028# a_9838_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X578 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X579 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X580 VCM a_n784_42308# C0_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X581 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X582 VSS a_11599_46634# a_13759_46122# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X583 a_14127_45572# a_11823_42460# a_14033_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X584 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X585 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X586 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X587 a_13569_43230# a_12379_42858# a_13460_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X588 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X589 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X590 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X591 a_5072_46660# a_4955_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X592 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X593 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X594 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X595 a_8037_42858# a_7871_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X596 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X597 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X598 VSS a_22591_46660# a_20820_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X599 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X600 a_3686_47026# a_2609_46660# a_3524_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X601 a_9672_43914# a_10057_43914# a_9801_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X602 VDD a_18429_43548# a_16823_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X603 VDD a_n2833_47464# CLK_DATA VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X604 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X605 a_17339_46660# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X606 VSS a_1606_42308# a_2351_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X607 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X608 a_16409_43396# a_16243_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X609 VDD a_n4209_37414# a_n4334_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X610 VSS a_9625_46129# a_10044_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X611 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X612 VSS a_n2302_39072# a_n4209_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X613 a_13468_44734# a_768_44030# a_13213_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X614 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X615 a_2124_47436# a_584_46384# a_2266_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X616 VDD a_n971_45724# a_2809_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X617 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X618 a_10809_44734# a_2063_45854# a_10809_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X619 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X620 a_7577_46660# a_7411_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X621 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X622 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X623 a_4921_42308# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X624 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X625 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X626 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X627 a_16023_47582# a_15507_47210# a_15928_47570# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X628 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X629 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X630 a_10193_42453# a_20712_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X631 a_12791_45546# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X632 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X633 a_6481_42558# a_n913_45002# a_1755_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X634 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X635 VSS a_n881_46662# a_n659_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X636 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X637 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X638 a_14955_43940# a_14537_43396# a_15037_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X639 VSS C2_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X640 a_n2956_38680# a_n2472_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X641 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X642 VREF_GND a_14097_32519# C4_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X643 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X644 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X645 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X646 VDD a_21188_45572# a_21363_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X647 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X648 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X649 a_15682_43940# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X650 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X651 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X652 a_18907_42674# a_18727_42674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X653 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X654 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X655 a_12545_42858# a_12379_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X656 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X657 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X658 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X659 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X660 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X661 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X662 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X663 C9_P_btm a_n4064_39616# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X664 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X665 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X666 a_15125_43396# a_15095_43370# a_15037_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X667 VREF a_20692_30879# C6_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=0.35
X668 a_13720_44458# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X669 a_20974_43370# a_22485_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X670 a_18548_42308# a_18494_42460# a_18057_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X671 a_2998_44172# a_584_46384# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X672 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X673 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X674 a_n875_44318# a_n2065_43946# a_n984_44318# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X675 w_11334_34010# a_18194_35068# EN_VIN_BSTR_N w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X676 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X677 a_n2293_42834# a_8049_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X678 VSS a_4743_44484# a_4791_45118# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X679 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X680 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X681 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X682 a_3626_43646# a_3232_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X683 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X684 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X685 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X686 VSS a_n2438_43548# a_n2433_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X687 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X688 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X689 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X690 a_n1076_43230# a_n2157_42858# a_n1423_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X691 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X692 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X693 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X694 VDD a_17973_43940# a_18079_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X695 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X696 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X697 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X698 VREF_GND a_17538_32519# C8_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X699 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X700 VDD a_22223_46124# a_20205_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X701 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X702 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X703 a_4704_46090# a_4883_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X704 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X705 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X706 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X707 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X708 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X709 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X710 a_17478_45572# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X711 a_5815_47464# a_6151_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X712 DATA[3] a_7227_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X713 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X714 a_22609_38406# a_22521_39511# CAL_N VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X715 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X716 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X717 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X718 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X719 VSS a_19864_35138# a_21589_35634# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X720 VSS a_n3420_39616# a_n2946_39866# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X721 VDAC_P C0_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X722 a_17034_45572# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X723 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X724 a_133_42852# a_n97_42460# a_n13_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X725 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X726 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X727 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X728 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X729 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X730 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X731 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X732 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X733 a_n1925_46634# a_8162_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X734 a_21350_47026# a_20273_46660# a_21188_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X735 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X736 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X737 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X738 VDD a_2713_42308# a_2903_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X739 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X740 a_n3674_39304# a_n2840_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X741 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X742 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X743 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X744 a_n4315_30879# a_n2302_40160# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X745 a_13565_43940# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X746 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X747 VDD a_1823_45246# a_2202_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X748 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X749 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X750 VSS a_n3690_38304# a_n3420_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X751 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X752 a_2211_45572# a_2063_45854# a_1848_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X753 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X754 VSS a_16112_44458# a_14673_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X755 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X756 VSS a_3316_45546# a_3260_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X757 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X758 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X759 VDD a_n443_46116# a_2896_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X760 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X761 a_21177_47436# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X762 VSS a_9290_44172# a_13943_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X763 a_n3674_37592# a_196_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X764 a_n310_47570# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X765 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X766 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X767 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X768 a_421_43172# a_n97_42460# a_n13_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X769 a_18780_47178# a_18597_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X770 VSS a_8791_42308# a_5934_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X771 VDD a_17339_46660# a_18051_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X772 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X773 VSS a_n2840_46090# a_n2956_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X774 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X775 a_n2661_43370# a_10907_45822# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X776 a_9396_43370# a_4883_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X777 VDD a_19333_46634# a_19123_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X778 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X779 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X780 a_5755_42852# a_n97_42460# a_5837_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X781 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X782 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X783 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X784 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X785 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X786 a_n4251_39392# a_n4318_39304# a_n4334_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X787 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X788 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X789 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X790 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X791 a_805_46414# a_472_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X792 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X793 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X794 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X795 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X796 VDD a_n1076_43230# a_n901_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X797 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X798 VDD a_4520_42826# a_4093_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X799 a_21845_43940# a_12549_44172# a_19692_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X800 a_15415_45028# a_15227_44166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X801 a_12469_46902# a_12251_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X802 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X803 a_19479_31679# a_22223_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X804 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X805 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X806 VSS a_22165_42308# a_22223_42860# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X807 a_7542_44172# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X808 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X809 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X810 a_3080_42308# a_2903_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X811 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X812 VDD a_10249_46116# a_11186_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X813 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X814 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X815 a_3905_42558# a_2382_45260# a_3823_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X816 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X817 a_12347_46660# a_11901_46660# a_12251_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X818 VSS a_16137_43396# a_16414_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X819 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X820 a_5066_45546# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X821 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X822 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X823 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X824 VSS C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X825 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X826 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X827 a_14581_44484# a_13249_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X828 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X829 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X830 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X831 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X832 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X833 a_2113_38308# a_1343_38525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X834 a_n473_42460# a_n755_45592# a_n327_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X835 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X836 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X837 VDD a_n1699_43638# a_n1809_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X838 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X839 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X840 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X841 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X842 a_13759_47204# a_13717_47436# a_13675_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X843 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X844 a_n3420_39616# a_n3690_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X845 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X846 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X847 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X848 C4_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X849 VDD a_9127_43156# a_5891_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X850 a_2779_44458# a_1423_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X851 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X852 a_n967_46494# a_n2157_46122# a_n1076_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X853 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X854 VDD a_19319_43548# a_19268_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.195 ps=1.39 w=1 l=0.15
X855 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X856 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X857 a_1123_46634# a_948_46660# a_1302_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X858 a_n755_45592# a_n809_44244# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X859 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X860 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X861 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X862 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X863 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X864 a_5807_45002# a_16763_47508# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X865 a_3726_37500# a_3754_38470# VDAC_Ni VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X866 a_6293_42852# a_5755_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X867 a_2952_47436# a_3160_47472# a_3094_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X868 a_8120_45572# a_8034_45724# a_n1925_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X869 a_11541_44484# a_11691_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X870 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X871 VSS a_10083_42826# a_7499_43078# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X872 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X873 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X874 VSS a_21589_35634# SMPL_ON_N VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X875 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X876 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X877 VDD a_n1630_35242# a_18194_35068# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X878 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X879 a_4880_45572# a_5066_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X880 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X881 VIN_P EN_VIN_BSTR_P C0_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X882 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X883 a_5257_43370# a_5907_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X884 COMP_P a_1239_39587# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X885 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X886 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X887 a_3497_42558# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X888 VSS a_1123_46634# a_584_46384# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X889 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X890 a_16223_45938# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X891 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X892 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X893 a_2711_45572# a_768_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X894 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X895 a_4883_46098# a_21363_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X896 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X897 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X898 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X899 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X900 VSS a_2553_47502# a_2487_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X901 VDD a_12469_46902# a_12359_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X902 a_6453_43914# a_6109_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X903 a_7765_42852# a_7227_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X904 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X905 a_18450_45144# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X906 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X907 a_17786_45822# a_15861_45028# a_17478_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X908 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X909 a_6765_43638# a_6547_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X910 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X911 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X912 a_12089_42308# a_11551_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X913 a_16547_43609# a_16414_43172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X914 a_n914_46116# a_n1991_46122# a_n1076_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X915 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X916 a_1343_38525# a_1177_38525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X917 VSS a_n4334_40480# a_n4064_40160# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X918 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X919 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X920 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X921 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X922 a_3221_46660# a_3177_46902# a_3055_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X923 a_6667_45809# a_6472_45840# a_6977_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X924 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X925 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X926 a_6643_43396# a_6197_43396# a_6547_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X927 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X928 a_n1190_43762# a_n2267_43396# a_n1352_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X929 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X930 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X931 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X932 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X933 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X934 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X935 a_5837_45348# a_5807_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X936 a_5565_43396# a_4905_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X937 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X938 a_1307_43914# a_2779_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X939 a_7418_45067# a_7229_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X940 a_1793_42852# a_742_44458# a_1709_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X941 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X942 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X943 VDD a_10227_46804# a_10083_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X944 a_11301_43218# a_10922_42852# a_11229_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X945 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X946 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X947 VSS C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X948 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X949 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X950 VSS a_13291_42460# a_13249_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X951 a_18341_45572# a_18175_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X952 a_19113_45348# a_19321_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X953 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X954 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X955 a_8696_44636# a_16855_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X956 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X957 a_12189_44484# a_8975_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X958 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X959 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X960 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X961 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X962 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X963 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X964 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X965 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X966 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X967 a_n1736_46482# a_n1853_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X968 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X969 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X970 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X971 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X972 a_n4064_37984# a_n4334_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X973 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X974 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X975 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X976 a_1239_47204# a_1209_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X977 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X978 a_1606_42308# a_1576_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X979 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X980 VDD VDAC_Ni a_6886_37412# VSS sky130_fd_pr__nfet_03v3_nvt ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X981 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X982 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X983 VDD a_n443_42852# a_6481_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X984 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X985 a_16795_42852# a_n97_42460# a_16877_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X986 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X987 a_18315_45260# a_18587_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X988 VSS a_768_44030# a_3600_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X989 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X990 VDD a_12005_46116# a_n1741_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X991 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X992 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X993 VDD a_4958_30871# a_17531_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X994 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X995 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X996 a_17973_43940# a_17737_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X997 a_18900_46660# a_18834_46812# a_18285_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X998 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X999 VSS a_22821_38993# a_22876_39857# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1000 a_6419_46155# a_5257_43370# a_6347_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1001 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1002 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1003 a_18597_46090# a_19431_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1004 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1005 a_3737_43940# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1006 VDD a_1823_45246# a_4419_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X1007 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1008 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1009 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1010 EN_VIN_BSTR_P VDD a_n1386_35608# VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.9
X1011 VDD a_4007_47204# DATA[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1012 VSS a_21496_47436# a_13507_46334# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1013 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1014 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1015 VSS a_10723_42308# a_5742_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1016 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1017 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1018 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1019 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1020 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1021 a_11823_42460# a_15051_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1022 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1023 VSS a_n4209_38216# a_n4251_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1024 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1025 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1026 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1027 a_12891_46348# a_4915_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1028 VSS a_20679_44626# a_20640_44752# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1029 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1030 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1031 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1032 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1033 a_21115_43940# a_20935_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1034 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1035 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1036 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1037 a_n1821_43396# a_n2267_43396# a_n1917_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1038 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1039 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1040 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1041 VDD a_10951_45334# a_10775_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1042 a_20850_46155# a_19692_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X1043 VDD a_13661_43548# a_18587_45118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1044 a_11649_44734# a_3232_43370# a_n2661_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.174 ps=1.39 w=1 l=0.15
X1045 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1046 a_17364_32525# a_22959_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1047 a_20820_30879# a_22591_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1048 VSS a_21359_45002# a_21101_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X1049 EN_VIN_BSTR_P VDD a_n83_35174# VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.9
X1050 a_18989_43940# a_18451_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1051 a_6197_43396# a_6031_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1052 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1053 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X1054 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1055 VDD a_12891_46348# a_13213_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1056 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1057 VREF_GND a_13467_32519# C1_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1058 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1059 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1060 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1061 VSS a_n4334_39392# a_n4064_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1062 a_8873_43396# a_5891_43370# a_8791_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1063 VDD a_584_46384# a_3540_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X1064 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1065 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1066 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1067 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1068 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1069 C9_P_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1070 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1071 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1072 C6_N_btm a_5742_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1073 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1074 a_10809_44484# a_10057_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1075 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1076 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1077 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1078 a_n4318_38216# a_n2472_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1079 VSS C0_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1080 a_6545_47178# a_6419_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X1081 a_6109_44484# a_5518_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1082 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1083 a_13258_32519# a_19647_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1084 VDD a_n901_46420# a_n443_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X1085 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1086 VDD a_11599_46634# a_18819_46122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1087 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1088 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1089 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1090 a_15682_43940# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1091 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X1092 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1093 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1094 a_n1435_47204# a_n1605_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1095 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1096 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1097 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1098 a_14113_42308# a_13575_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1099 VSS a_4646_46812# a_4651_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1100 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1101 VSS a_n2472_46090# a_n2956_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1102 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1103 a_4958_30871# a_17124_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1104 VSS a_22223_42860# a_22400_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1105 a_13381_47204# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1106 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1107 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1108 C0_P_btm a_n3565_37414# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1109 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1110 VDD a_1208_46090# a_472_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1111 VSS a_n2302_39072# a_n4209_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1112 VSS a_18479_47436# a_19452_47524# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1113 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1114 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1115 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1116 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1117 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1118 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1119 a_22545_38993# a_22459_39145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1120 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X1121 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1122 a_n443_46116# a_n901_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1123 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1124 a_20623_45572# a_20107_45572# a_20528_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1125 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1126 VSS a_n3565_39304# a_n3607_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1127 a_12281_43396# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1128 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1129 a_15486_42560# a_15764_42576# a_15720_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1130 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1131 C1_P_btm a_n4209_37414# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1132 VSS a_n1613_43370# a_8649_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1133 a_15765_45572# a_15599_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1134 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1135 VSS a_n2946_39866# a_n3565_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1136 VCM a_5932_42308# C3_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1137 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1138 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1139 a_n1613_43370# a_5815_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X1140 VSS a_14495_45572# a_n881_46662# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1141 a_10617_44484# a_10440_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1142 VDD a_5111_44636# a_8487_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1143 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1144 VSS a_1847_42826# a_2905_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1145 a_n2267_44484# a_n2433_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1146 a_20708_46348# a_15227_44166# a_20850_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1147 a_1115_44172# a_453_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1148 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1149 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1150 VSS COMP_P a_n1329_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X1151 VSS a_15861_45028# a_17023_45118# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1152 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1153 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1154 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1155 a_16292_46812# a_5807_45002# a_16434_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1156 a_n4064_39072# a_n4334_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X1157 a_17325_44484# a_15227_44166# a_16979_44734# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1158 a_5534_30871# a_12563_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1159 a_15803_42450# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1160 VSS a_3381_47502# a_3315_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1161 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1162 VDD a_9863_46634# a_2063_45854# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X1163 VDD a_n1838_35608# SMPL_ON_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1164 VIN_N EN_VIN_BSTR_N C3_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1165 VSS a_584_46384# a_3457_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1166 a_3863_42891# a_3681_42891# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1167 VDD a_n2840_43370# a_n4318_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1168 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1169 VDD a_9049_44484# a_9313_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X1170 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1171 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1172 a_11541_44484# a_11453_44696# a_n2661_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1173 VDD a_376_46348# a_171_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1174 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1175 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1176 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1177 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1178 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1179 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1180 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1181 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1182 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1183 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1184 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1185 VDD a_1431_47204# DATA[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1186 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1187 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1188 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1189 a_21589_35634# a_19864_35138# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1190 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1191 a_19553_46090# a_19335_46494# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1192 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1193 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1194 a_18727_42674# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1195 a_n1613_43370# a_5815_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X1196 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1197 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1198 VDD a_n2302_37984# a_n4209_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1199 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1200 a_n1925_42282# a_4185_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1201 VDD a_19164_43230# a_19339_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1202 VSS a_17591_47464# a_16327_47482# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1203 VSS a_n3690_38304# a_n3420_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1204 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1205 VSS a_4361_42308# a_21855_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1206 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1207 a_2479_44172# a_2905_42968# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X1208 VDD a_8103_44636# a_7640_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X1209 a_n1741_47186# a_12891_46348# a_12839_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1210 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1211 a_8192_45572# a_8162_45546# a_8120_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X1212 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1213 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1214 a_5009_45028# a_3090_45724# a_4927_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1215 a_12549_44172# a_20567_45036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1216 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1217 VSS a_n2840_42282# a_n3674_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1218 a_5129_47502# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1219 a_14840_46494# a_13759_46122# a_14493_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1220 VSS a_2324_44458# a_949_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1221 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1222 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1223 VSS a_n913_45002# a_2713_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1224 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1225 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1226 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1227 VDD a_n863_45724# a_1221_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X1228 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1229 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1230 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1231 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1232 a_2307_45899# a_n237_47217# a_1848_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1233 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1234 VDD a_n4209_39304# a_n4334_39392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X1235 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1236 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X1237 a_8601_46660# a_7411_46660# a_8492_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1238 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1239 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1240 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1241 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1242 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1243 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1244 a_n2946_39072# a_n2956_39304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1245 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1246 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1247 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1248 a_15861_45028# a_15595_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1249 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1250 VSS a_n1613_43370# a_3221_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1251 VSS a_1239_39587# COMP_P VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1252 a_1756_43548# a_768_44030# a_1987_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1253 a_3754_39134# a_7754_39300# VSS sky130_fd_pr__res_high_po_0p35 l=18
X1254 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1255 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1256 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1257 a_n4318_40392# a_n2840_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1258 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1259 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1260 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1261 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1262 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1263 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1264 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1265 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1266 VSS a_18143_47464# a_12861_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1267 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1268 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1269 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1270 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1271 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1272 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1273 a_19332_42282# a_19511_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1274 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1275 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1276 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1277 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1278 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1279 VSS a_17583_46090# a_13259_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X1280 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1281 VSS a_7754_38470# a_6886_37412# VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1282 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1283 a_20623_43914# a_19321_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1284 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1285 a_n3420_39616# a_n3690_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1286 VSS a_17499_43370# a_n1059_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1287 a_n2661_46634# a_13017_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1288 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1289 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1290 a_4185_45348# a_3065_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1291 VDD a_19321_45002# a_20567_45036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1292 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1293 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1294 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1295 VDD a_6545_47178# a_6575_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1296 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1297 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1298 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1299 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1300 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1301 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1302 VDD a_18285_46348# a_18051_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.16 ps=1.32 w=1 l=0.15
X1303 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1304 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1305 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1306 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1307 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1308 a_2864_46660# a_2747_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1309 VSS a_n809_44244# a_n755_45592# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1310 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1311 VDD a_1307_43914# a_2253_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1312 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1313 a_18374_44850# a_18248_44752# a_17970_44736# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1314 a_n913_45002# a_1307_43914# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1315 a_13351_46090# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X1316 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1317 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1318 a_18194_35068# a_n1630_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1319 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1320 a_13657_42308# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1321 a_3090_45724# a_19321_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X1322 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1323 VSS a_1239_39043# comp_n VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1324 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1325 a_375_42282# a_413_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1326 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1327 a_5700_37509# VSS VDAC_Pi VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1328 VSS a_10903_43370# a_10057_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1329 a_10334_44484# a_10157_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1330 a_2113_38308# a_2113_38308# a_2113_38308# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=3.02 ps=24.88 w=1 l=0.15
X1331 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1332 VSS a_22959_46124# a_20692_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1333 a_n3674_39768# a_n2472_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1334 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1335 a_584_46384# a_1123_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1336 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1337 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1338 VREF a_n4209_39304# C7_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1339 VSS a_20107_42308# a_7174_31319# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1340 VSS a_n2438_43548# a_n133_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1341 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1342 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1343 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1344 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1345 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1346 VDAC_N C1_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1347 a_n4209_39590# a_n2302_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1348 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1349 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1350 a_526_44458# a_3147_46376# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1351 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1352 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1353 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1354 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1355 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1356 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1357 a_20301_43646# a_19692_46634# a_20556_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1358 VDD a_n901_46420# a_n914_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1359 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1360 VSS a_1177_38525# a_1343_38525# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1361 a_n971_45724# a_104_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1362 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1363 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1364 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1365 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1366 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1367 a_20447_31679# a_22959_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1368 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1369 a_n4334_38304# a_n4318_38216# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1370 VSS a_13348_45260# a_13159_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1371 a_8685_42308# a_8515_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1372 VSS a_n881_46662# a_6517_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1373 a_768_44030# a_13487_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X1374 VDD a_14493_46090# a_14383_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1375 VSS a_6491_46660# a_6851_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1376 a_n327_42308# a_n357_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X1377 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1378 a_22485_44484# a_22315_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1379 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1380 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1381 VSS C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1382 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1383 a_8605_42826# a_8387_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1384 a_15673_47210# a_15507_47210# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1385 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1386 a_1709_42852# a_n863_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1387 VDD a_n1736_42282# a_n4318_37592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1388 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1389 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1390 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1391 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1392 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1393 VREF a_19721_31679# C2_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1394 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1395 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1396 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1397 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1398 VSS a_895_43940# a_2537_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X1399 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1400 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1401 a_13249_42308# a_10903_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1402 a_8945_43396# a_3537_45260# a_8873_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1403 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1404 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1405 a_17609_46634# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1406 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1407 VDD a_11599_46634# a_18175_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1408 a_601_46902# a_383_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1409 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1410 a_4640_45348# a_4574_45260# a_4558_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1411 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1412 a_n467_45028# a_n745_45366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1413 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1414 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1415 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1416 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1417 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1418 a_1208_46090# a_765_45546# a_1337_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1419 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1420 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1421 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1422 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1423 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1424 VSS a_n863_45724# a_2905_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1425 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1426 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1427 a_3820_44260# a_2382_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X1428 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1429 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1430 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1431 C5_P_btm a_n4064_38528# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1432 VSS a_16721_46634# a_16655_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1433 a_21588_30879# a_22223_47212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1434 a_16877_42852# a_16823_43084# a_16795_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1435 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1436 VSS a_17715_44484# a_17737_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1437 a_16241_47178# a_16023_47582# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1438 a_17665_42852# a_17595_43084# a_14539_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X1439 VSS a_n2438_43548# a_n2157_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1440 a_16759_43396# a_16409_43396# a_16664_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1441 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1442 a_22876_39857# a_22545_38993# a_22780_39857# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1443 a_12359_47026# a_11735_46660# a_12251_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1444 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1445 a_5883_43914# a_8333_44056# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X1446 VDD a_n3565_39590# a_n3690_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X1447 VDD a_4007_47204# DATA[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1448 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1449 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1450 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1451 a_1990_45572# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1452 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1453 a_5072_46660# a_4955_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1454 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1455 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1456 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1457 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1458 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1459 VDD a_3357_43084# a_22591_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1460 VSS a_3815_47204# a_4007_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X1461 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1462 a_1736_39587# a_1736_39043# a_2112_39137# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1463 a_15803_42450# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1464 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1465 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1466 a_20528_46660# a_20411_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1467 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1468 a_n3607_39392# a_n3674_39304# a_n3690_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X1469 a_21421_42336# a_16327_47482# a_21335_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1470 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1471 VDD a_n4064_39616# a_n2216_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X1472 a_n1838_35608# a_n1386_35608# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1473 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1474 a_6655_43762# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1475 a_14371_46494# a_13925_46122# a_14275_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1476 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1477 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1478 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1479 VDD a_3503_45724# a_3218_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X1480 VSS a_n901_43156# a_n443_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1481 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1482 VDD a_n2840_43914# a_n4318_39768# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1483 a_15037_43940# a_13556_45296# a_14955_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1484 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1485 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1486 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1487 VDD a_10467_46802# a_10428_46928# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1488 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1489 a_15060_45348# a_13661_43548# a_14976_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X1490 a_9895_44260# a_9290_44172# a_9801_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1491 VDD a_6171_42473# a_5379_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1492 a_5009_45028# a_5147_45002# a_5093_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1493 a_13904_45546# a_10903_43370# a_14127_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1494 a_3537_45260# a_7287_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1495 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1496 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1497 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1498 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1499 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1500 VDD a_8696_44636# a_17478_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X1501 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1502 a_19900_46494# a_18985_46122# a_19553_46090# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1503 a_3935_42891# a_3905_42865# a_3863_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1504 VSS a_n881_46662# a_11117_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1505 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1506 C3_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1507 VSS C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1508 VSS a_n4334_39616# a_n4064_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1509 DATA[0] a_327_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1510 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1511 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1512 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1513 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1514 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1515 DATA[2] a_4007_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1516 a_15682_46116# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1517 a_1057_46660# a_n133_46660# a_948_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1518 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1519 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1520 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1521 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1522 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1523 VSS a_2982_43646# a_21487_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1524 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1525 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1526 a_21363_45546# a_21188_45572# a_21542_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1527 a_18204_44850# a_17767_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1528 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1529 a_n443_42852# a_n901_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1530 VSS a_11823_42460# a_11322_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1531 a_n447_43370# a_n2497_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1532 VSS a_n4064_38528# a_n2302_38778# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X1533 a_17324_43396# a_16409_43396# a_16977_43638# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1534 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1535 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1536 a_15095_43370# a_15567_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X1537 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1538 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1539 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1540 a_10150_46912# a_10428_46928# a_10384_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1541 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1542 VSS a_n2472_42282# a_n4318_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1543 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1544 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1545 VDD a_n1630_35242# a_n1532_35090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1546 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1547 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1548 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1549 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1550 a_8492_46660# a_7577_46660# a_8145_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1551 a_5649_42852# a_5111_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1552 VDD a_18287_44626# a_18248_44752# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1553 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1554 a_20894_47436# a_20990_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X1555 a_19636_46660# a_19594_46812# a_19333_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X1556 a_10249_46116# a_9823_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X1557 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1558 a_739_46482# a_n743_46660# a_376_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1559 VSS a_10775_45002# a_10180_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X1560 a_2896_43646# a_2479_44172# a_2982_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X1561 a_10227_46804# a_14955_47212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1562 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1563 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1564 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1565 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1566 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1567 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1568 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1569 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1570 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1571 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1572 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1573 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1574 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1575 a_12791_45546# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1576 VSS a_5807_45002# a_11691_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1577 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1578 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1579 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1580 VSS a_2382_45260# a_2304_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X1581 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1582 a_n4315_30879# a_n2302_40160# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1583 VSS a_3357_43084# a_22591_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1584 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1585 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1586 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1587 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1588 a_6298_44484# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1589 a_949_44458# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1590 VDD a_n901_46420# a_n443_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1591 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1592 VDD a_2277_45546# a_2307_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1593 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1594 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1595 a_10053_45546# a_8746_45002# a_10306_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X1596 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1597 a_n2956_39768# a_n2840_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1598 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1599 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1600 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1601 VDD a_4361_42308# a_21855_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1602 VDD a_17591_47464# a_16327_47482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1603 VSS a_6945_45028# a_22223_46124# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1604 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1605 a_n3565_39590# a_n2946_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1606 VDD a_5257_43370# a_5263_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1607 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1608 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1609 a_18494_42460# a_18907_42674# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1610 VDAC_Ni VSS a_5088_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1611 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1612 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1613 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1614 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1615 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1616 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1617 a_n1151_42308# a_n1329_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1618 SMPL_ON_P a_n1838_35608# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1619 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1620 a_16763_47508# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1621 a_21259_43561# a_4190_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1622 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1623 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1624 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1625 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1626 a_8349_46414# a_8016_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1627 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1628 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1629 a_17970_44736# a_18287_44626# a_18245_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1630 VDD a_1431_47204# DATA[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1631 a_1123_46634# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1632 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1633 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1634 a_n237_47217# a_8667_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X1635 VSS C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1636 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1637 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1638 a_5837_42852# a_3537_45260# a_5755_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1639 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1640 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1641 VSS a_19692_46634# a_19636_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1642 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1643 a_8697_45572# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1644 a_1145_45348# a_n863_45724# a_626_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1645 VSS a_5934_30871# a_8515_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1646 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1647 VSS a_1239_47204# a_1431_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X1648 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1649 a_22705_38406# a_22521_40055# a_22609_38406# VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1650 a_11173_44260# a_10729_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X1651 VSS a_17591_47464# a_16327_47482# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1652 VDD a_n4334_38304# a_n4064_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1653 a_22165_42308# a_21887_42336# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1654 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1655 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1656 VDD a_8952_43230# a_9127_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1657 VSS a_n4064_37440# a_n2302_37690# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X1658 a_5244_44056# a_5147_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1659 VSS a_2127_44172# a_n2661_45010# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X1660 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1661 a_n3565_38502# a_n2946_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X1662 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1663 a_n2956_37592# a_n2472_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1664 VSS a_15493_43940# a_22959_43948# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1665 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1666 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1667 a_19339_43156# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1668 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1669 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1670 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1671 VDD a_n1177_44458# a_n1190_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1672 VDD a_n1920_47178# a_n2312_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1673 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1674 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1675 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1676 VDD a_16292_46812# a_15811_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1677 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1678 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1679 a_5164_46348# a_4927_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X1680 a_9482_43914# a_9838_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1681 a_20835_44721# a_20679_44626# a_20980_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1682 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1683 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1684 a_5837_42852# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1685 VSS a_5937_45572# a_8781_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1686 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1687 a_7221_43396# a_6031_43396# a_7112_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1688 a_10037_47542# a_n881_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X1689 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1690 C7_N_btm a_20820_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1691 VSS a_5937_45572# a_8560_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X1692 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1693 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1694 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1695 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1696 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1697 VSS a_15559_46634# a_13059_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X1698 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1699 a_5385_46902# a_5167_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1700 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1701 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1702 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1703 VDD a_21589_35634# SMPL_ON_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1704 VDD a_10334_44484# a_10440_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1705 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1706 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1707 a_19597_46482# a_19553_46090# a_19431_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1708 VDD a_n2302_37984# a_n4209_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1709 a_18051_46116# a_18189_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X1710 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1711 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1712 a_16414_43172# a_n1059_45260# a_16328_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X1713 a_15493_43940# a_14955_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1714 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1715 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1716 a_21297_46660# a_20107_46660# a_21188_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1717 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1718 a_11813_46116# a_11387_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X1719 VSS SMPL_ON_P a_n1605_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1720 VDD a_4699_43561# a_3539_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1721 VSS a_n3420_39072# a_n2946_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X1722 DATA[4] a_9067_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1723 a_5894_47026# a_4817_46660# a_5732_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1724 VDD a_n97_42460# a_16245_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1725 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1726 VDD a_13163_45724# a_11962_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1727 a_15433_44458# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1728 VDD a_16327_47482# a_20980_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1729 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1730 a_18114_32519# a_22223_45036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1731 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1732 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1733 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1734 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1735 a_n452_44636# a_n1151_42308# a_n310_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1736 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1737 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1738 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1739 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1740 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1741 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1742 VDD a_22959_43396# a_17364_32525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1743 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1744 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1745 VSS a_n357_42282# a_7573_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X1746 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1747 a_n4064_37984# a_n4334_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1748 VDD a_1307_43914# a_4149_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X1749 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1750 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1751 VDD a_9863_47436# a_9804_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1752 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1753 a_22821_38993# a_22400_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1754 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1755 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1756 a_3754_39134# a_7754_38968# VSS sky130_fd_pr__res_high_po_0p35 l=18
X1757 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1758 a_4649_43172# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1759 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1760 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1761 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1762 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1763 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1764 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1765 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1766 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1767 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1768 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1769 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1770 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1771 a_526_44458# a_3147_46376# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X1772 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1773 a_22465_38105# a_22775_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1774 VSS a_1848_45724# a_1799_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1775 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1776 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1777 a_20885_45572# a_20841_45814# a_20719_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1778 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1779 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1780 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1781 a_10554_47026# a_10428_46928# a_10150_46912# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1782 a_n746_45260# a_n1177_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1783 a_7_44811# a_n1151_42308# a_n452_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1784 VDD a_2324_44458# a_15682_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1785 VDD a_10355_46116# a_8199_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1786 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1787 a_4181_43396# a_4093_43548# a_n2661_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1788 a_21005_45260# a_21101_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X1789 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1790 a_n3565_37414# a_n2946_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X1791 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1792 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1793 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1794 VDD a_2437_43646# a_22223_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1795 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1796 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1797 a_3754_38802# a_7754_38968# VSS sky130_fd_pr__res_high_po_0p35 l=18
X1798 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1799 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1800 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1801 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1802 a_2075_43172# a_1307_43914# a_n913_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1803 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1804 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1805 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1806 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1807 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1808 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1809 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1810 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1811 comp_n a_1239_39043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1812 VSS a_17499_43370# a_n1059_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1813 VDD a_n2840_45002# a_n2810_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1814 VSS a_12861_44030# a_17339_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1815 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1816 a_10057_43914# a_10807_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1817 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1818 a_5343_44458# a_7963_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1819 a_n1423_42826# a_n1641_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1820 VDD a_11827_44484# a_22223_45036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1821 VDD a_n2472_43914# a_n3674_39768# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1822 a_526_44458# a_3147_46376# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X1823 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X1824 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1825 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1826 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1827 a_6945_45028# a_5937_45572# a_6945_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1828 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1829 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1830 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1831 VDD a_n3690_39616# a_n3420_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1832 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1833 a_20301_43646# a_13661_43548# a_743_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1834 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1835 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1836 a_n2216_39866# a_n2442_46660# a_n2302_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1837 VDD a_22000_46634# a_15227_44166# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1838 a_n3674_38216# a_n2104_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1839 VSS a_2889_44172# a_413_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1840 VSS a_n97_42460# a_n144_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1841 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1842 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1843 a_133_42852# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X1844 a_16321_45348# a_1307_43914# a_16019_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
X1845 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1846 VDD a_9290_44172# a_13070_42354# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X1847 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1848 VDD a_22465_38105# a_22521_39511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1849 a_n3420_39072# a_n3690_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X1850 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1851 a_n2860_38778# a_n2956_38680# a_n2946_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1852 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1853 a_22465_38105# a_22775_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1854 a_10555_44260# a_10729_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X1855 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1856 a_6517_45366# a_5937_45572# a_6431_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1857 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1858 a_14401_32519# a_22223_43948# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1859 VDD a_5111_44636# a_5837_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X1860 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1861 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1862 VSS a_9290_44172# a_13070_42354# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1863 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1864 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1865 VDD a_9290_44172# a_10586_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1866 a_16751_45260# a_8696_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1867 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1868 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1869 VSS a_5068_46348# a_4955_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1870 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1871 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1872 a_1736_39587# a_1736_39043# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X1873 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1874 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1875 a_n913_45002# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1876 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1877 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1878 VSS a_11599_46634# a_15507_47210# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1879 VSS a_768_44030# a_644_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1880 VDD a_n357_42282# a_16877_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1881 a_5193_43172# a_3905_42865# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1882 VSS a_18783_43370# a_18525_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X1883 a_12465_44636# a_5807_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1884 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1885 a_3540_43646# a_1414_42308# a_3626_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X1886 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1887 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1888 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1889 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1890 a_5421_42558# a_5379_42460# a_5337_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1891 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1892 VSS a_n3690_38528# a_n3420_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1893 a_21363_45546# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1894 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1895 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1896 VDD a_12861_44030# a_17609_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1897 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1898 a_n2956_38216# a_n2472_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1899 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1900 VCM a_4958_30871# C9_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1901 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1902 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1903 a_13885_46660# a_13607_46688# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1904 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1905 a_2232_45348# a_1609_45822# a_n2293_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X1906 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1907 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1908 a_5691_45260# a_6171_45002# a_5837_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1909 a_9801_44260# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1910 VCM a_3080_42308# C2_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1911 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1912 a_15743_43084# a_19339_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1913 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1914 VSS a_22591_43396# a_14209_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1915 a_327_44734# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X1916 VSS a_7499_43078# a_8746_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1917 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1918 VSS a_2437_43646# a_22223_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1919 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1920 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1921 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1922 a_6547_43396# a_6197_43396# a_6452_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1923 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1924 a_20556_43646# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1925 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1926 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1927 a_1987_43646# a_742_44458# a_1891_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1928 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1929 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1930 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1931 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1932 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1933 a_648_43396# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X1934 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1935 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1936 VDD CLK a_8953_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1937 VDD a_n23_47502# a_7_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1938 a_17609_46634# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X1939 a_3602_45348# a_3537_45260# a_3495_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X1940 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1941 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1942 VDD a_2982_43646# a_21487_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1943 a_13661_43548# a_18780_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1944 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1945 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1946 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1947 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1948 a_11323_42473# a_5742_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1949 a_9313_44734# a_3232_43370# a_9159_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1950 C6_P_btm a_5742_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1951 a_14383_46116# a_13759_46122# a_14275_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1952 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1953 a_2813_43396# a_2479_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1954 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1955 a_16721_46634# a_16388_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1956 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1957 VREF a_20820_30879# C7_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1958 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1959 VDD a_526_44458# a_9885_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1960 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1961 VDD a_15681_43442# a_15781_43660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X1962 a_6125_45348# a_3232_43370# a_5691_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1963 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1964 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1965 a_10907_45822# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X1966 a_14955_43396# a_9145_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1967 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1968 a_3429_45260# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1969 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1970 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1971 a_8128_46384# a_7903_47542# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1972 VDD a_15227_44166# a_17969_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X1973 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1974 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1975 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1976 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1977 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1978 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1979 VSS C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1980 a_n2860_37690# a_n2956_37592# a_n2946_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1981 DATA[0] a_327_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1982 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1983 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1984 VSS a_7287_43370# a_3537_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1985 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1986 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1987 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1988 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1989 C4_P_btm a_n3420_38528# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1990 a_15682_46116# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1991 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1992 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1993 a_18599_43230# a_18083_42858# a_18504_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1994 DATA[2] a_4007_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X1995 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1996 a_18057_42282# a_18494_42460# a_18214_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X1997 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1998 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1999 a_11117_47542# a_4915_47217# a_11031_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2000 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2001 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2002 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2003 VDD a_22400_42852# a_22521_40599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2004 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2005 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2006 a_7112_43396# a_6197_43396# a_6765_43638# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2007 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2008 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2009 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2010 a_584_46384# a_1123_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2011 VSS a_n3690_37440# a_n3420_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2012 VSS a_n901_43156# a_n443_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2013 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2014 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2015 a_19240_46482# a_19123_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2016 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2017 VCM a_5742_30871# C6_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2018 VSS a_10193_42453# a_10149_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2019 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2020 VDD a_10193_42453# a_10210_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X2021 a_564_42282# a_743_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2022 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2023 VSS a_2324_44458# a_15682_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2024 VSS a_n967_45348# a_n961_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2025 a_21195_42852# a_20922_43172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2026 VDD a_6575_47204# a_9067_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2027 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2028 a_22612_30879# a_22959_47212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2029 a_21188_46660# a_20273_46660# a_20841_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2030 a_13749_43396# a_13661_43548# a_13667_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X2031 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2032 VSS a_n2840_45546# a_n2810_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2033 a_13490_45394# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2034 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2035 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2036 a_n2840_43914# a_n2661_43922# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2037 a_n822_43940# a_n1899_43946# a_n984_44318# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2038 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2039 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2040 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2041 a_21613_42308# a_21335_42336# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X2042 a_14537_43396# a_13059_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2043 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2044 VDAC_Pi a_3754_38470# a_4338_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2045 a_7112_43396# a_6031_43396# a_6765_43638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2046 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2047 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2048 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2049 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2050 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2051 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2052 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2053 a_n4064_39616# a_n4334_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2054 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2055 a_n23_47502# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2056 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2057 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2058 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2059 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2060 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2061 a_14543_43071# a_5534_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2062 VDD a_7227_45028# a_7230_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2063 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2064 VDD a_19900_46494# a_20075_46420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2065 VSS a_16327_47482# a_19597_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2066 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2067 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2068 a_9823_46155# a_n743_46660# a_9751_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2069 a_18214_42558# a_16137_43396# a_18057_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2070 VDD a_22959_43948# a_17538_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2071 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2072 a_n3690_38304# a_n3674_38216# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2073 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2074 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2075 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2076 a_15009_46634# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X2077 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2078 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2079 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2080 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2081 VSS a_10227_46804# a_15521_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X2082 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2083 a_17591_47464# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2084 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2085 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2086 a_22485_44484# a_22315_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2087 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2088 a_n1644_44306# a_n1761_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2089 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2090 VDD a_n1329_42308# a_n1151_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2091 VDD RST_Z a_8530_39574# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2092 VSS a_13507_46334# a_18184_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2093 a_n630_44306# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2094 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2095 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2096 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2097 a_18783_43370# a_15743_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2098 VSS C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2099 a_n4064_38528# a_n4334_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2100 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2101 a_8325_42308# a_n913_45002# a_8337_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2102 VSS a_22521_40599# a_22469_40625# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2103 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2104 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2105 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X2106 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2107 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2108 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2109 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2110 a_21973_42336# a_20202_43084# a_21887_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2111 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2112 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2113 VSS a_n1613_43370# a_645_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2114 a_10341_42308# a_9803_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2115 VSS a_10807_43548# a_11173_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2116 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2117 VSS a_16327_47482# a_20885_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2118 a_n1920_47178# a_n1741_47186# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2119 a_9127_43156# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2120 VSS a_5257_43370# a_3905_42865# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2121 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2122 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2123 VSS a_n2946_39072# a_n3565_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2124 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2125 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2126 VDD a_n2472_45002# a_n2956_37592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2127 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2128 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2129 a_13259_45724# a_17583_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2130 VSS a_10586_45546# a_10544_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X2131 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2132 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2133 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2134 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2135 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2136 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2137 a_16751_45260# a_17023_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2138 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2139 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2140 VSS a_n4209_38502# a_n4251_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2141 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2142 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2143 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2144 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2145 VSS a_10083_42826# a_7499_43078# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2146 a_n2840_42826# a_n2661_42834# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2147 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2148 VSS a_7227_42308# a_6123_31319# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2149 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2150 a_1302_46660# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2151 a_5907_45546# a_6194_45824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X2152 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2153 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2154 a_n2302_37984# a_n2810_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2155 a_13059_46348# a_15559_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2156 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2157 COMP_P a_1239_39587# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2158 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2159 VREF_GND a_14209_32519# C5_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2160 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2161 a_3065_45002# a_3318_42354# a_3581_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X2162 a_16023_47582# a_15673_47210# a_15928_47570# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2163 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2164 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2165 VSS a_n881_46662# a_n935_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2166 VDD a_21487_43396# a_13467_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2167 C6_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2168 VDD a_n443_42852# a_997_45618# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2169 a_2553_47502# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2170 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2171 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2172 a_13635_43156# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2173 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2174 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2175 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2176 a_8568_45546# a_8199_44636# a_8791_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2177 a_4338_37500# a_3754_38470# VDAC_Pi VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2178 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2179 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2180 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2181 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2182 VDD a_564_42282# a_n1630_35242# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2183 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2184 a_n473_42460# a_n971_45724# a_n327_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X2185 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2186 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2187 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2188 a_16335_44484# a_13661_43548# a_16241_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X2189 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2190 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2191 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2192 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2193 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2194 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2195 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2196 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2197 VDD a_15861_45028# a_17023_45118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2198 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2199 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2200 a_5205_44734# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2201 a_7499_43078# a_10083_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=2.61 w=1 l=0.15
X2202 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2203 VSS a_1123_46634# a_1057_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2204 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2205 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2206 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2207 w_1575_34946# a_n1532_35090# EN_VIN_BSTR_P w_1575_34946# sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2208 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2209 a_5700_37509# VSS VDAC_Pi VDD sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2210 a_n4064_37440# a_n4334_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2211 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2212 VSS a_13259_45724# a_18315_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2213 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2214 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2215 VSS a_22223_43396# a_13887_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2216 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2217 a_n1453_44318# a_n1899_43946# a_n1549_44318# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2218 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2219 a_11682_45822# a_11322_45546# a_11525_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2220 VDD a_22591_45572# a_19963_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2221 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2222 a_18429_43548# a_18525_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X2223 a_5934_30871# a_8791_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2224 a_509_45822# a_n1099_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2225 a_4190_30871# a_19332_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2226 a_20980_44850# a_20766_44850# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X2227 a_3381_47502# a_2905_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2228 VDD a_3537_45260# a_4649_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2229 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2230 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2231 VDD a_1423_45028# a_9838_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2232 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2233 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2234 a_6682_46660# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2235 a_20273_45572# a_20107_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2236 VDD a_11963_45334# a_11787_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X2237 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2238 a_n755_45592# a_n809_44244# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2239 a_19256_45572# a_18175_45572# a_18909_45814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2240 VSS a_5937_45572# a_9159_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2241 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2242 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2243 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2244 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2245 VSS a_3699_46634# a_3633_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2246 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2247 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2248 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2249 VSS a_n2438_43548# a_n2157_46122# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2250 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2251 a_14226_46987# a_14180_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2252 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2253 a_n722_43218# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2254 a_n2840_45002# a_n2661_45010# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2255 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2256 VSS a_8953_45546# a_9241_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2257 a_12005_46436# a_2063_45854# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2258 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2259 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2260 a_9885_43396# a_8270_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2261 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2262 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2263 VSS a_n4209_37414# a_n4251_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2264 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2265 a_18817_42826# a_18599_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2266 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2267 VDD a_n3690_39616# a_n3420_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2268 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2269 EN_VIN_BSTR_P a_n1532_35090# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2270 VDAC_Pi VSS a_5700_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2271 VDD a_167_45260# a_1423_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2272 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2273 VSS a_4704_46090# a_1823_45246# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2274 a_16886_45144# a_8696_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X2275 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2276 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2277 VSS C0_dummy_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2278 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2279 a_11688_45572# a_11652_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X2280 a_8953_45002# CLK VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2281 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2282 a_4520_42826# a_1823_45246# a_4743_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2283 a_949_44458# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2284 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2285 a_n3420_39072# a_n3690_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2286 VDD a_n2104_42282# a_n3674_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2287 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2288 VDD RST_Z a_14311_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2289 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2290 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2291 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2292 a_19339_43156# a_19164_43230# a_19518_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2293 a_19721_31679# a_22959_45036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2294 a_458_43396# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X2295 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2296 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2297 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2298 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2299 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2300 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2301 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2302 a_11453_44696# a_17719_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X2303 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2304 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2305 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2306 a_22717_36887# a_22459_39145# a_22609_37990# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2307 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2308 VDD a_n3420_37984# a_n2860_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2309 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2310 a_13711_45394# a_12891_46348# a_13348_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2311 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2312 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2313 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2314 a_1138_42852# a_791_42968# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X2315 a_16664_43396# a_16547_43609# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2316 a_21259_43561# a_4190_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2317 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2318 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2319 a_10586_45546# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2320 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2321 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2322 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2323 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2324 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2325 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2326 VSS a_n3690_38528# a_n3420_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2327 VSS a_11599_46634# a_15599_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2328 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2329 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2330 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X2331 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2332 a_196_42282# a_375_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2333 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2334 VSS a_n881_46662# a_7989_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2335 a_7832_46660# a_7715_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2336 VDD a_n2109_45247# en_comp VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2337 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2338 a_3633_46660# a_2443_46660# a_3524_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2339 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2340 a_15928_47570# a_15811_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2341 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2342 a_2127_44172# a_2675_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2343 a_9885_43646# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X2344 VSS a_n2472_45546# a_n2956_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2345 a_n2472_43914# a_n2293_43922# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2346 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2347 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2348 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2349 VDD a_12991_46634# a_12978_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2350 VDD a_1667_45002# a_n863_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2351 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2352 a_n4209_39304# a_n2302_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2353 a_5837_45028# a_3232_43370# a_5691_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X2354 VDD a_21195_42852# a_21671_42860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2355 a_14084_46812# a_n1151_42308# a_14226_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2356 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2357 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2358 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2359 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2360 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2361 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2362 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2363 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2364 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2365 VSS a_n913_45002# a_4921_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2366 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2367 a_14209_32519# a_22591_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2368 a_12427_45724# a_12791_45546# a_12749_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2369 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2370 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2371 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2372 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2373 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2374 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2375 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2376 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2377 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2378 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2379 a_12553_44484# a_12465_44636# a_n2661_43922# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2380 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2381 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2382 a_5829_43940# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2383 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2384 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2385 a_16237_45028# a_n743_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2386 VDD a_22959_45036# a_19721_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2387 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2388 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2389 a_14761_44260# a_14673_44172# a_n2293_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2390 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2391 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2392 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2393 VSS a_n1613_43370# a_5429_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2394 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2395 VDD a_n452_45724# a_n1853_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2396 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2397 VSS a_21363_46634# a_21297_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2398 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2399 VDD a_584_46384# a_2998_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2400 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2401 VSS C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2402 VDD a_15959_42545# a_15890_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X2403 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2404 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2405 VSS a_4699_43561# a_3539_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2406 VSS a_10227_46804# a_13157_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2407 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2408 VSS a_n2946_39866# a_n3565_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2409 a_n4209_38502# a_n2302_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X2410 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2411 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2412 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2413 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2414 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2415 a_n144_43396# a_n971_45724# a_n447_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X2416 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2417 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2418 a_17538_32519# a_22959_43948# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2419 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2420 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2421 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2422 a_16680_45572# a_15599_45572# a_16333_45814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2423 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2424 VSS a_5937_45572# a_6101_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X2425 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2426 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2427 a_8387_43230# a_7871_42858# a_8292_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2428 a_15231_43396# a_9145_43396# a_15125_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X2429 a_9672_43914# a_8199_44636# a_9895_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2430 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2431 VDD a_22731_47423# a_13717_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2432 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2433 VDD a_9290_44172# a_13667_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X2434 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2435 a_n3420_37984# a_n3690_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2436 VDD a_17767_44458# a_17715_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X2437 VDD a_7845_44172# a_7542_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X2438 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2439 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2440 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2441 VDD a_10903_43370# a_13163_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.06615 ps=0.735 w=0.42 l=0.15
X2442 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2443 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2444 a_n2840_44458# a_n2661_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2445 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2446 VDD a_n863_45724# a_945_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X2447 a_22400_42852# a_22223_42860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2448 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2449 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2450 VDD a_12549_44172# a_10949_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.195 ps=1.39 w=1 l=0.15
X2451 a_4933_42558# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2452 VSS a_9482_43914# a_10157_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2453 a_19333_46634# a_19466_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X2454 a_13565_44260# a_12891_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2455 VSS a_n3690_37440# a_n3420_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2456 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2457 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2458 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2459 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2460 a_n2293_46098# a_5663_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X2461 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2462 VSS a_11453_44696# a_22959_47212# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2463 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2464 VSS a_12563_42308# a_5534_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2465 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2466 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2467 a_n2472_42826# a_n2293_42834# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2468 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2469 a_n13_43084# a_n443_42852# a_133_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2470 a_7920_46348# a_8128_46384# a_8062_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2471 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2472 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2473 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2474 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2475 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2476 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2477 a_2698_46116# a_2521_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X2478 a_15785_43172# a_15743_43084# a_15095_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X2479 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2480 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2481 a_8654_47026# a_7577_46660# a_8492_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2482 VDD a_21363_46634# a_21350_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2483 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2484 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2485 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2486 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2487 VDD a_n809_44244# a_n822_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2488 a_766_43646# a_626_44172# a_458_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X2489 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2490 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2491 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2492 a_n784_42308# a_n961_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2493 a_12895_43230# a_12379_42858# a_12800_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2494 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2495 VSS a_8191_45002# a_8137_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2496 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2497 a_15959_42545# a_15803_42450# a_16104_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X2498 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2499 VSS a_805_46414# a_739_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2500 a_11341_43940# a_3232_43370# a_11173_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.19825 ps=1.26 w=0.65 l=0.15
X2501 a_5210_46482# a_5164_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2502 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2503 VDD a_7705_45326# a_7735_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2504 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2505 a_13720_44458# a_13661_43548# a_13940_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2506 a_2162_46660# a_2107_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2507 VSS a_n4334_39392# a_n4064_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2508 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2509 a_n1423_42826# a_n1641_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2510 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2511 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2512 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2513 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2514 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2515 a_n2956_39304# a_n2840_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2516 VDD a_11415_45002# a_n2661_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2517 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2518 a_15037_43940# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X2519 VDD a_1606_42308# a_2351_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2520 a_2277_45546# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2521 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2522 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2523 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2524 VDD a_14180_45002# a_13017_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X2525 a_3232_43370# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2526 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2527 a_6903_46660# a_6755_46942# a_6540_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2528 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2529 VDD a_n2302_40160# a_n4315_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2530 a_22521_40055# en_comp VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2531 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2532 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2533 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2534 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2535 VSS C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2536 a_1576_42282# a_1755_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2537 VDD a_8199_44636# a_8191_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X2538 a_n4209_37414# a_n2302_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X2539 VSS a_21855_43396# a_13678_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2540 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2541 a_7573_43172# a_7499_43078# a_7227_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2542 VDD a_18989_43940# a_19006_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2543 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2544 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2545 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2546 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2547 VSS a_6540_46812# a_6491_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2548 VDD a_22223_45572# a_19479_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2549 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2550 VIN_N EN_VIN_BSTR_N C0_dummy_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2551 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2552 VSS a_2903_42308# a_3080_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2553 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2554 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2555 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2556 VSS a_n863_45724# a_n906_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X2557 a_3823_42558# a_3065_45002# a_3905_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2558 a_n2840_44458# a_n2661_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2559 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2560 VSS a_2779_44458# a_1307_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2561 VSS a_5263_45724# a_5204_45822# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X2562 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2563 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2564 VDD a_2124_47436# a_1209_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2565 VSS a_2957_45546# a_2905_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2566 a_12925_46660# a_11735_46660# a_12816_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2567 a_376_46348# a_n743_46660# a_518_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2568 a_11415_45002# a_4915_47217# a_14581_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2569 VDD a_7754_40130# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.5
X2570 a_n2104_42282# a_n1925_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2571 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2572 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2573 a_n2472_45002# a_n2293_45010# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2574 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2575 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2576 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2577 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2578 a_21398_44850# a_20679_44626# a_20835_44721# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2579 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2580 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2581 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2582 VDD a_22521_40599# a_22705_38406# VDD sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2583 VSS a_8685_43396# a_15231_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X2584 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2585 VDD a_16333_45814# a_16223_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2586 a_16241_44484# a_2711_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X2587 a_3905_42865# a_5257_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2588 a_13485_45572# a_12549_44172# a_13385_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X2589 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2590 C3_P_btm a_n4209_38216# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2591 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2592 VSS a_10623_46897# a_10554_47026# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2593 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2594 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2595 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2596 VSS a_22959_45572# a_20447_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2597 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2598 a_19120_35138# a_18194_35068# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2599 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2600 VDD a_19987_42826# a_n2017_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.135 ps=1.27 w=1 l=0.15
X2601 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2602 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2603 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2604 a_9028_43914# a_9482_43914# a_9420_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2605 a_1343_38525# a_1177_38525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2606 a_n2860_39072# a_n2956_39304# a_n2946_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X2607 VSS a_17973_43940# a_18079_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X2608 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2609 a_9290_44172# a_13635_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2610 a_3059_42968# a_742_44458# a_2987_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2611 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2612 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2613 a_18194_35068# a_n1630_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2614 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2615 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2616 a_n452_44636# a_n467_45028# a_n310_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2617 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2618 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2619 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2620 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2621 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2622 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2623 VDD a_768_44030# a_2711_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2624 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2625 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2626 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2627 VDAC_N C0_dummy_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2628 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2629 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2630 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2631 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2632 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2633 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2634 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2635 VDD a_12281_43396# a_12563_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2636 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2637 VDD a_12741_44636# a_22959_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2638 SMPL_ON_N a_21589_35634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2639 a_8333_44734# a_3537_45260# a_8238_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X2640 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2641 VSS a_1177_38525# a_1343_38525# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2642 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2643 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2644 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2645 VSS C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2646 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2647 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2648 a_17124_42282# a_17303_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2649 a_12156_46660# a_11813_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2650 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2651 VDD a_n447_43370# a_n2129_43609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2652 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2653 VDD a_10809_44734# a_22959_46124# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2654 VSS a_1115_44172# a_n2293_45010# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X2655 a_5013_44260# a_1307_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2656 a_3357_43084# a_5257_43370# a_5565_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2657 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2658 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2659 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2660 a_n967_43230# a_n2157_42858# a_n1076_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2661 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2662 a_1568_43370# a_1847_42826# a_1793_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2663 a_11682_45822# a_10586_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X2664 a_n2012_44484# a_n2129_44697# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2665 a_18315_45260# a_15227_44166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X2666 a_14543_43071# a_5534_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2667 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2668 a_16147_45260# a_17478_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2669 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2670 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2671 a_19963_31679# a_22591_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2672 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2673 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2674 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2675 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2676 a_n967_45348# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2677 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2678 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2679 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2680 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2681 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2682 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2683 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2684 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2685 VSS a_7276_45260# a_7227_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2686 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2687 a_1241_44260# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X2688 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2689 VDD a_11599_46634# a_20107_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2690 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2691 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2692 VDD a_n809_44244# a_n755_45592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2693 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2694 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2695 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2696 a_n4334_40480# a_n4318_40392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2697 VSS a_n815_47178# a_n785_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2698 a_3175_45822# a_3090_45724# a_2957_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2699 a_14621_43646# a_14579_43548# a_14537_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2700 VDD a_n1386_35608# a_n1838_35608# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2701 VDD a_n2946_37984# a_n3565_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2702 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2703 VREF a_20205_31679# C4_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2704 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2705 VSS a_15227_44166# a_18900_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X2706 a_n310_44811# a_n356_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2707 VDD a_16977_43638# a_16867_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2708 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2709 VDD a_15227_44166# a_17749_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X2710 a_3147_46376# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X2711 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2712 a_12638_46436# a_12594_46348# a_12379_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2713 VSS a_2324_44458# a_6298_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2714 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2715 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2716 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2717 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2718 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2719 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2720 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2721 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2722 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2723 a_21071_46482# a_15227_44166# a_20708_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2724 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2725 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2726 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2727 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2728 a_9127_43156# a_8952_43230# a_9306_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2729 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2730 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2731 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2732 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2733 VDD a_1343_38525# a_2684_37794# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2734 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2735 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2736 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2737 a_961_42354# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2738 a_n1059_45260# a_17499_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2739 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2740 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2741 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2742 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2743 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2744 VSS a_8349_46414# a_8283_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2745 VSS a_11787_45002# a_11652_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X2746 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2747 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2748 VSS a_12741_44636# a_22959_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2749 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2750 a_4223_44672# a_3537_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2751 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2752 a_n1532_35090# a_n1630_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2753 a_509_45822# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2754 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2755 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2756 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2757 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2758 a_16119_47582# a_15673_47210# a_16023_47582# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2759 a_6452_43396# a_6293_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2760 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2761 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2762 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2763 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2764 VSS CLK a_8953_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2765 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2766 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2767 a_6194_45824# a_6472_45840# a_6428_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2768 a_3754_38802# a_7754_38636# VSS sky130_fd_pr__res_high_po_0p35 l=18
X2769 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2770 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2771 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2772 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2773 VDD a_n881_46662# a_11031_47542# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2774 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2775 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2776 VSS a_1209_47178# a_1239_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2777 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2778 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2779 a_12429_44172# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X2780 a_15559_46634# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X2781 a_11229_43218# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2782 a_16020_45572# a_15903_45785# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2783 a_10149_42308# a_9290_44172# a_9803_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2784 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2785 C3_P_btm a_5932_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2786 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2787 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2788 a_10793_43218# a_10083_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2789 VSS a_20708_46348# a_20411_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2790 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2791 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2792 C9_N_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2793 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2794 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2795 a_13635_43156# a_13460_43230# a_13814_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2796 a_n863_45724# a_1667_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2797 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2798 VDAC_N C2_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2799 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2800 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2801 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2802 a_12379_46436# a_12594_46348# a_12638_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2803 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2804 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2805 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2806 a_1209_43370# a_1049_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X2807 a_2982_43646# a_3232_43370# a_2813_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2808 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2809 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2810 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2811 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2812 a_21542_45572# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2813 VSS a_19647_42308# a_13258_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2814 a_n443_46116# a_n901_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2815 a_18985_46122# a_18819_46122# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2816 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2817 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2818 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2819 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2820 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2821 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2822 a_12839_46116# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2823 VDD a_n2438_43548# a_2443_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2824 VDD a_9028_43914# a_8975_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X2825 VDD a_17124_42282# a_4958_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2826 VSS a_10053_45546# a_9625_46129# VSS sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X2827 VSS a_380_45546# a_n356_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X2828 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2829 VSS a_20193_45348# a_21973_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2830 VSS a_196_42282# a_n3674_37592# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2831 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2832 VSS C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2833 a_17639_46660# a_17609_46634# a_765_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2834 VDD a_5257_43370# a_5826_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X2835 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2836 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2837 a_9803_42558# a_n97_42460# a_9885_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2838 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2839 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2840 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2841 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2842 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2843 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2844 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2845 VSS a_10227_46804# a_10553_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X2846 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2847 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2848 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2849 VSS a_n913_45002# a_12281_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2850 VSS a_18597_46090# a_16375_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2851 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2852 a_12816_46660# a_11901_46660# a_12469_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2853 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2854 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2855 a_n3565_39590# a_n2946_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2856 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2857 a_20205_45028# a_18184_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2858 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2859 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2860 a_n3420_37984# a_n3690_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2861 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2862 VDD a_13259_45724# a_13667_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X2863 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2864 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2865 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2866 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2867 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2868 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2869 a_n1736_42282# a_n1557_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2870 a_13747_46662# a_19386_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2871 VSS a_4791_45118# a_6165_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X2872 a_261_44278# a_n863_45724# a_175_44278# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2873 a_8325_42308# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2874 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2875 SMPL_ON_P a_n1838_35608# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2876 a_10623_46897# a_10467_46802# a_10768_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X2877 a_2675_43914# a_2998_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2878 a_18695_43230# a_18249_42858# a_18599_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2879 a_17957_46116# a_765_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X2880 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2881 a_17613_45144# a_8696_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2882 a_n4318_39304# a_n2840_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2883 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2884 a_18799_45938# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2885 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2886 VSS a_19862_44208# a_20922_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X2887 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2888 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2889 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2890 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2891 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2892 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2893 a_6151_47436# a_14311_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2894 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2895 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2896 VSS a_5129_47502# a_5063_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2897 VSS a_167_45260# a_2521_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2898 a_16333_45814# a_16115_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2899 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2900 a_3733_45822# a_n755_45592# a_3638_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X2901 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2902 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2903 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2904 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2905 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2906 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2907 SMPL_ON_N a_21589_35634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2908 a_13163_45724# a_13527_45546# a_13485_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2909 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2910 a_8605_42826# a_8387_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2911 a_1337_46116# a_1176_45822# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2912 a_n4209_38216# a_n2302_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2913 a_n83_35174# a_n1532_35090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2914 VDD a_4419_46090# a_n1925_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2915 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2916 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2917 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2918 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2919 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2920 a_20712_42282# a_n357_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2921 a_1241_43940# a_1467_44172# a_1443_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2922 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2923 VDD a_n961_42308# a_n784_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2924 a_7227_42852# a_n97_42460# a_7309_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2925 a_9145_43396# a_8791_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2926 a_14976_45348# a_13059_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2927 a_9863_47436# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X2928 a_743_42282# a_19692_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2929 VSS a_12891_46348# a_12638_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2930 a_4915_47217# a_12991_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2931 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2932 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2933 VSS a_1239_39587# COMP_P VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2934 a_n3674_38680# a_n2840_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2935 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2936 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2937 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2938 VCM a_4958_30871# C9_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2939 VSS a_3539_42460# a_3065_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2940 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2941 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2942 a_17801_45144# a_17613_45144# a_17719_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X2943 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2944 VDD a_n4209_39590# a_n4334_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X2945 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2946 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2947 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2948 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2949 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2950 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2951 a_18787_45572# a_18341_45572# a_18691_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2952 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2953 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2954 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2955 a_10922_42852# a_10796_42968# a_10518_42984# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2956 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2957 a_3754_39964# a_7754_40130# VSS sky130_fd_pr__res_high_po_0p35 l=18
X2958 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2959 VDD a_n4334_40480# a_n4064_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2960 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2961 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2962 VDD a_526_44458# a_3232_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2963 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2964 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2965 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2966 a_n1630_35242# a_564_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2967 a_167_45260# a_2202_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2968 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2969 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2970 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2971 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2972 VDD a_11967_42832# a_20512_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2973 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2974 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2975 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2976 VDD a_16019_45002# a_15903_45785# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2977 a_2896_43646# a_n443_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2978 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2979 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2980 VSS a_9067_47204# DATA[4] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2981 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2982 a_12005_46116# a_10903_43370# a_12005_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2983 a_n2312_38680# a_n2104_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2984 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2985 a_14097_32519# a_22959_42860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2986 a_n2288_47178# a_n2109_47186# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2987 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2988 a_6999_46987# a_3877_44458# a_6540_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X2989 a_8199_44636# a_10355_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X2990 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2991 a_3429_45260# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X2992 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2993 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2994 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2995 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2996 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2997 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2998 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2999 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3000 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3001 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3002 C8_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3003 a_9293_42558# a_9223_42460# a_8953_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X3004 a_4338_37500# VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.589 ps=4.42 w=1.9 l=0.15
X3005 VDD a_n2302_40160# a_n4315_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3006 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3007 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3008 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3009 VDD a_n452_47436# a_n815_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3010 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3011 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3012 a_13807_45067# a_13556_45296# a_13348_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3013 a_14309_45348# a_2711_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X3014 a_1176_45822# a_997_45618# a_1260_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X3015 VDD a_13159_45002# a_n2661_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3016 VSS a_20269_44172# a_19319_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3017 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3018 a_16104_42674# a_15890_42674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X3019 a_2981_46116# a_2804_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3020 a_4185_45028# a_3877_44458# a_4185_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3021 a_n1655_43396# a_n1699_43638# a_n1821_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3022 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3023 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3024 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3025 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3026 a_22731_47423# SMPL_ON_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3027 a_n722_46482# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3028 VSS a_n443_42852# a_997_45618# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X3029 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3030 a_6945_45348# a_5205_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3031 a_4791_45118# a_4743_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X3032 a_21513_45002# a_21363_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3033 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3034 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3035 VSS a_1576_42282# a_1606_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3036 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3037 a_n1533_46116# a_n2157_46122# a_n1641_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3038 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3039 a_15227_44166# a_22000_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3040 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3041 VDAC_P C0_dummy_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3042 VSS en_comp a_1177_38525# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3043 a_n743_46660# a_n1021_46688# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3044 a_n4064_40160# a_n4334_40480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X3045 a_2075_43172# a_1307_43914# a_n913_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3046 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3047 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3048 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3049 VSS a_5205_44484# a_6756_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3050 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3051 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3052 comp_n a_1239_39043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3053 VDD a_19321_45002# a_3090_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X3054 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3055 VSS a_3483_46348# a_13829_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3056 VDD a_327_44734# a_375_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3057 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3058 VDD a_7754_40130# a_11206_38545# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3059 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3060 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3061 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3062 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3063 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3064 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3065 VDD a_526_44458# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3066 VDD a_5937_45572# a_6671_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3067 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3068 VDD a_n863_45724# a_458_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X3069 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3070 VDD a_n4334_38304# a_n4064_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X3071 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3072 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3073 VDD a_1756_43548# a_1467_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.28 ps=2.56 w=1 l=0.15
X3074 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3075 a_20269_44172# a_20365_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X3076 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3077 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3078 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3079 VDD a_4791_45118# a_5066_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3080 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3081 VDD a_14976_45028# a_15227_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3082 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3083 VSS a_13904_45546# a_12594_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X3084 VSS a_8953_45546# a_8568_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3085 VDAC_Pi a_3754_38470# a_4338_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3086 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3087 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3088 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3089 a_16112_44458# a_15227_44166# a_16335_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3090 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3091 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3092 VSS a_20974_43370# a_20749_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3093 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3094 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3095 a_n913_45002# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3096 VSS a_16327_47482# a_17021_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3097 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3098 a_16388_46812# a_17957_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1725 ps=1.345 w=1 l=0.15
X3099 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3100 a_n4318_37592# a_n1736_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3101 VSS a_20159_44458# a_19321_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X3102 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3103 VDD a_9672_43914# a_2107_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3104 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3105 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3106 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3107 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3108 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3109 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3110 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3111 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3112 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3113 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3114 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3115 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3116 VSS a_6151_47436# a_8189_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3117 VDD a_12549_44172# a_17609_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3118 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3119 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3120 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3121 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3122 VDD a_1239_39043# comp_n VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3123 a_6229_45572# a_6194_45824# a_5907_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3124 VDD a_19700_43370# a_n97_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3125 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3126 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3127 a_6851_47204# a_6491_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3128 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3129 a_8423_43396# a_n443_42852# a_8317_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X3130 VDD a_19615_44636# a_18579_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X3131 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3132 a_1755_42282# a_n913_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3133 a_18799_45938# a_18175_45572# a_18691_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3134 VDD a_7499_43078# a_8697_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X3135 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3136 a_n4209_39304# a_n2302_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X3137 VDD a_6765_43638# a_6655_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3138 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3139 VSS a_2324_44458# a_6298_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3140 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3141 a_n1741_47186# a_12005_46116# a_12379_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X3142 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3143 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3144 VDD a_22223_47212# a_21588_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3145 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3146 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3147 a_685_42968# a_n443_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3148 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3149 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3150 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3151 a_10467_46802# a_11599_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3152 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3153 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3154 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3155 a_17749_42852# a_17701_42308# a_17665_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3156 VDD a_n443_42852# a_15781_43660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X3157 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3158 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3159 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3160 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3161 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3162 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3163 a_18599_43230# a_18249_42858# a_18504_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3164 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3165 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3166 CLK_DATA a_n2833_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X3167 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3168 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3169 VDD a_7920_46348# a_7715_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3170 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3171 a_3537_45260# a_7287_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3172 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3173 a_2809_45028# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X3174 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3175 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3176 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3177 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3178 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3179 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3180 a_7832_46660# a_7715_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3181 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3182 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3183 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3184 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3185 VSS a_4905_42826# a_4520_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3186 a_3873_46454# a_n881_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X3187 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3188 VSS a_20202_43084# a_21421_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3189 a_6709_45028# a_6431_45366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3190 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3191 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3192 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3193 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3194 a_20623_43914# a_19321_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3195 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3196 a_20193_45348# a_18494_42460# a_20205_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3197 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3198 VSS a_9313_45822# a_11459_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X3199 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3200 a_n443_42852# a_n901_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3201 a_n4318_39768# a_n2840_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3202 VSS a_22469_40625# a_22717_36887# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3203 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3204 a_6428_45938# a_5907_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3205 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3206 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3207 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3208 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3209 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3210 a_n2104_46634# a_n1925_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3211 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3212 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3213 VSS a_7287_43370# a_3537_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3214 EN_VIN_BSTR_N VDD a_19120_35138# VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.9
X3215 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3216 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3217 a_2987_42968# a_1847_42826# a_2905_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3218 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3219 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3220 a_11031_47542# a_4915_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3221 VSS a_12991_46634# a_12925_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3222 VDAC_Ni a_7754_38636# VSS sky130_fd_pr__res_high_po_0p35 l=18
X3223 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3224 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3225 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3226 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3227 VDAC_N C2_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3228 VSS a_20894_47436# a_20843_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3229 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3230 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3231 a_10752_42852# a_10083_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3232 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3233 a_13076_44458# a_9482_43914# a_13468_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X3234 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3235 a_n1809_43762# a_n2433_43396# a_n1917_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3236 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3237 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3238 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3239 a_17970_44736# a_18248_44752# a_18204_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X3240 a_5663_43940# a_5883_43914# a_5841_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X3241 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3242 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3243 a_n2302_38778# a_n2312_38680# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3244 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3245 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3246 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3247 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3248 a_16588_47582# a_15507_47210# a_16241_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3249 VSS a_4099_45572# a_3483_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3250 VSS a_14539_43914# a_16112_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3251 a_16867_43762# a_16243_43396# a_16759_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3252 a_n745_45366# a_n746_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3253 a_10518_42984# a_10835_43094# a_10793_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X3254 C2_P_btm a_n3420_37984# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X3255 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3256 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3257 VIN_P EN_VIN_BSTR_P C5_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X3258 a_n37_45144# a_n443_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3259 VSS a_11341_43940# a_22223_43948# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3260 VSS a_8530_39574# a_3754_38470# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3261 a_18287_44626# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3262 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3263 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3264 a_20159_44458# a_20362_44736# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X3265 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3266 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3267 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3268 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3269 a_6969_46634# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3270 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3271 DATA[5] a_11459_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3272 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3273 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3274 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3275 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3276 a_18861_43218# a_18817_42826# a_18695_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3277 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3278 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3279 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3280 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3281 a_11322_45546# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3282 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3283 a_n3674_37592# a_196_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3284 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3285 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3286 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3287 a_n1809_43762# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3288 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3289 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3290 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3291 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3292 a_4419_46090# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X3293 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3294 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3295 VDD a_11189_46129# a_11133_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X3296 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3297 a_15959_42545# a_15764_42576# a_16269_42308# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X3298 VIN_P EN_VIN_BSTR_P a_n923_35174# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3299 VSS a_7640_43914# a_7584_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3300 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3301 VDD a_7227_47204# DATA[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X3302 a_n1076_46494# a_n1991_46122# a_n1423_46090# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3303 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3304 a_16375_45002# a_18597_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3305 a_4235_43370# a_3935_42891# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X3306 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3307 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3308 VDD a_n1699_44726# a_n1809_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3309 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3310 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3311 a_21177_47436# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X3312 a_7418_45394# a_7229_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3313 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3314 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3315 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3316 a_22000_46634# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3317 VDD a_7542_44172# a_7499_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3318 a_11309_47204# a_11031_47542# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3319 VDD a_1307_43914# a_3353_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3320 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3321 a_3905_42308# a_2382_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3322 a_8483_43230# a_8037_42858# a_8387_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3323 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3324 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3325 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3326 a_n2104_46634# a_n1925_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3327 a_7281_43914# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X3328 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3329 a_9028_43914# a_9290_44172# a_9248_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3330 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3331 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3332 a_453_43940# a_175_44278# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3333 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3334 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3335 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3336 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3337 VDD a_n2302_38778# a_n4209_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3338 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3339 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3340 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3341 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3342 a_15521_42308# a_15486_42560# a_15051_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3343 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3344 VDD a_4700_47436# a_3785_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3345 a_18909_45814# a_18691_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3346 a_11551_42558# a_n97_42460# a_11633_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3347 VSS a_11459_47204# DATA[5] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3348 VDD a_15227_44166# a_15415_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X3349 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3350 VSS a_16327_47482# a_20397_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X3351 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3352 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3353 VDD a_8270_45546# a_9165_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3354 a_n809_44244# a_n984_44318# a_n630_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3355 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3356 VDD a_948_46660# a_1123_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3357 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3358 a_20766_44850# a_20679_44626# a_20362_44736# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X3359 VDD a_15009_46634# a_14180_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3360 a_13385_45572# a_10903_43370# a_13297_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X3361 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3362 VDD a_13777_45326# a_13807_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3363 VSS a_n755_45592# a_n39_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3364 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3365 a_14976_45028# a_14797_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X3366 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3367 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3368 a_6886_37412# VDAC_Pi VDD VSS sky130_fd_pr__nfet_03v3_nvt ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X3369 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3370 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3371 a_6419_46482# a_6165_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X3372 a_n2302_37690# a_n2810_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3373 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3374 VSS a_768_44030# a_5244_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3375 VSS a_n2946_39072# a_n3565_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3376 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3377 a_20623_45572# a_20273_45572# a_20528_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3378 VDD a_8199_44636# a_8336_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X3379 VSS a_9396_43370# a_5111_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3380 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3381 a_743_42282# a_13661_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3382 a_n1190_44850# a_n2267_44484# a_n1352_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3383 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3384 a_20009_46494# a_18819_46122# a_19900_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3385 a_7309_42852# a_5891_43370# a_7227_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3386 a_n2312_39304# a_n1920_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3387 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3388 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3389 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3390 VSS a_n4064_40160# a_n2302_40160# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X3391 a_12991_43230# a_12545_42858# a_12895_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3392 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3393 a_22397_42558# a_n913_45002# a_17303_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3394 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3395 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3396 VSS a_3905_42865# a_5013_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3397 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3398 VSS C0_dummy_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3399 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3400 a_22765_42852# a_15743_43084# a_18184_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3401 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3402 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3403 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3404 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3405 COMP_P a_1239_39587# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3406 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3407 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3408 a_7705_45326# a_7229_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3409 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3410 a_3065_45002# a_1823_45246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X3411 VSS a_10405_44172# a_8016_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3412 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3413 a_742_44458# a_n443_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3414 VDD a_526_44458# a_3905_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3415 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3416 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3417 a_310_45028# a_n37_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X3418 VDD a_3232_43370# a_2982_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3419 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3420 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3421 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3422 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3423 VSS a_18184_42460# a_20256_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.11375 ps=1 w=0.65 l=0.15
X3424 a_19466_46812# a_13747_46662# a_19929_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3425 VDD a_16241_47178# a_16131_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3426 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3427 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3428 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3429 VSS a_768_44030# a_9028_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X3430 a_20850_46482# a_19692_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3431 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3432 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3433 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3434 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3435 a_12089_42308# a_11551_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3436 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3437 a_11173_43940# a_2063_45854# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3438 a_3457_43396# a_1414_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3439 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3440 a_8034_45724# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3441 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3442 VDD a_5907_46634# a_5894_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3443 a_22000_46634# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3444 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3445 a_5841_46660# a_4651_46660# a_5732_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3446 VSS a_3699_46348# a_3160_47472# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X3447 VSS a_22223_45036# a_18114_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3448 a_2437_43396# a_1568_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3449 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3450 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3451 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3452 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3453 a_2448_45028# a_2382_45260# a_n2293_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X3454 VDD a_n2104_46634# a_n2312_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3455 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3456 a_21167_46155# a_20916_46384# a_20708_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3457 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3458 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3459 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3460 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3461 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3462 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3463 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3464 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3465 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3466 a_5205_44484# a_5343_44458# a_5289_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3467 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3468 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3469 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3470 a_7499_43078# a_10083_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3471 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3472 VDD a_n2302_37690# a_n4209_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3473 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3474 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3475 a_948_46660# a_33_46660# a_601_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3476 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3477 VSS a_21005_45260# a_19778_44110# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3478 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3479 a_9241_46436# a_n237_47217# a_8049_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3480 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3481 a_15015_46420# a_14840_46494# a_15194_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3482 VSS a_13487_47204# a_768_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X3483 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3484 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3485 VDD a_20567_45036# a_12549_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3486 a_22717_37285# a_22459_39145# a_22609_38406# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3487 a_21398_44850# a_20640_44752# a_20835_44721# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X3488 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3489 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3490 a_5527_46155# a_5204_45822# a_5068_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3491 a_1823_45246# a_4704_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3492 a_1606_42308# a_1576_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3493 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3494 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3495 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3496 VSS a_4235_43370# a_4181_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3497 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3498 VSS a_18194_35068# a_19120_35138# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3499 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3500 VDD a_18783_43370# a_18525_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X3501 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3502 VCM a_5534_30871# C7_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X3503 a_n881_46662# a_14495_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X3504 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3505 a_n1821_44484# a_n2267_44484# a_n1917_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3506 a_21188_45572# a_20107_45572# a_20841_45814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3507 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3508 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3509 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3510 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3511 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3512 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3513 VSS a_8270_45546# a_8192_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X3514 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3515 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3516 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3517 a_5891_43370# a_9127_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3518 VDD a_n863_45724# a_3059_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3519 VDD a_17609_46634# a_765_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3520 VSS a_n755_45592# a_3503_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3521 a_19237_31679# a_22959_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3522 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3523 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3524 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3525 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3526 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3527 a_n4334_38528# a_n4318_38680# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3528 VSS C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3529 a_12156_46660# a_11813_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3530 a_n901_43156# a_n1076_43230# a_n722_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3531 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3532 a_n2810_45028# a_n2840_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3533 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3534 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3535 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3536 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3537 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3538 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3539 a_16333_45814# a_16115_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3540 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3541 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3542 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3543 a_n913_45002# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3544 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3545 a_16795_42852# a_n97_42460# a_16877_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3546 a_6905_45572# a_6151_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X3547 VDD a_21188_46660# a_21363_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3548 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3549 VDD a_5934_30871# a_8515_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3550 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3551 a_14180_45002# a_13059_46348# a_14403_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3552 a_16405_45348# a_16375_45002# a_16321_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3553 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3554 w_1575_34946# a_n923_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=10.615 ps=76.96 w=3.75 l=15
X3555 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3556 VREF a_19963_31679# C3_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X3557 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3558 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3559 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3560 VDD a_3422_30871# a_22315_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3561 a_2123_42473# a_n784_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3562 VSS a_n1613_43370# a_n1287_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3563 VSS a_22223_43948# a_14401_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3564 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3565 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3566 a_19518_43218# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3567 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3568 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3569 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3570 VSS a_20075_46420# a_20009_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3571 VSS a_16922_45042# a_16751_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3572 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3573 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3574 a_1049_43396# a_458_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3575 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3576 VDD a_3232_43370# a_11341_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.3925 ps=1.785 w=1 l=0.15
X3577 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3578 VDD a_526_44458# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3579 VDD a_n237_47217# a_8270_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3580 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3581 a_1848_45724# a_n237_47217# a_1990_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3582 VDD a_14539_43914# a_12465_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3583 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3584 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3585 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3586 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3587 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3588 VDD a_n881_46662# a_7903_47542# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3589 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3590 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3591 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3592 VDD a_n1423_46090# a_n1533_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3593 VDD a_5111_44636# a_5421_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3594 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3595 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3596 a_11778_45572# a_10193_42453# a_11688_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X3597 a_20623_46660# a_20107_46660# a_20528_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3598 a_6347_46155# a_6165_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3599 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3600 VDD a_21359_45002# a_21101_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X3601 a_4700_47436# a_n443_46116# a_4842_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3602 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3603 C4_P_btm a_n3565_38502# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X3604 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3605 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3606 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3607 VDD a_5755_42308# a_5932_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3608 a_14113_42308# a_13575_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3609 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3610 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3611 a_17333_42852# a_16795_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3612 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3613 a_10695_43548# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X3614 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3615 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3616 a_4958_30871# a_17124_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3617 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3618 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3619 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3620 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3621 VSS a_19339_43156# a_19273_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3622 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3623 a_8387_43230# a_8037_42858# a_8292_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3624 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3625 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3626 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3627 VSS a_16327_47482# a_18861_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3628 VDD a_n2840_44458# a_n4318_40392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3629 VDD a_15004_44636# a_14815_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3630 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3631 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3632 VSS a_1823_45246# a_3602_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3633 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3634 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3635 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3636 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3637 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3638 a_n4334_37440# a_n4318_37592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3639 VDD a_18780_47178# a_13661_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3640 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3641 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3642 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3643 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3644 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3645 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3646 a_2455_43940# a_895_43940# a_2253_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3647 a_13667_43396# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X3648 CAL_P a_22465_38105# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3649 a_2680_45002# a_3065_45002# a_2809_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3650 a_21381_43940# a_21115_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X3651 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3652 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3653 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3654 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3655 VSS a_22521_39511# a_22469_39537# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3656 a_15781_43660# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X3657 a_380_45546# a_765_45546# a_509_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3658 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3659 a_16019_45002# a_16147_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.160875 ps=1.145 w=0.65 l=0.15
X3660 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3661 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3662 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3663 a_5534_30871# a_12563_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3664 a_12741_44636# a_6755_46942# a_16789_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3665 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3666 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3667 VDD a_3537_45260# a_4558_45348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3668 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3669 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3670 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3671 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3672 VSS a_2324_44458# a_15682_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3673 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3674 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3675 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3676 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3677 VDD a_n473_42460# a_n1761_44111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X3678 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3679 VSS a_7754_38470# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X3680 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3681 a_12895_43230# a_12545_42858# a_12800_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3682 a_20836_43172# a_20193_45348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3683 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3684 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3685 VSS a_n2833_47464# CLK_DATA VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3686 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3687 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3688 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3689 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3690 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3691 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X3692 a_726_44056# a_626_44172# a_644_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3693 a_6655_43762# a_6031_43396# a_6547_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3694 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3695 VDD a_1123_46634# a_584_46384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3696 DATA[5] a_11459_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X3697 VDD a_3232_43370# a_3626_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3698 a_5343_44458# a_7963_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3699 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3700 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3701 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3702 a_2889_44172# a_1414_42308# a_3052_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3703 a_9313_44734# a_5883_43914# a_9241_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3704 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3705 a_3483_46348# a_4099_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3706 a_2809_45028# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3707 VDD a_6171_45002# a_11827_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3708 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3709 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3710 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3711 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3712 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3713 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3714 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3715 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3716 VDD a_9625_46129# a_9569_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X3717 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3718 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3719 a_15567_42826# a_15227_44166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3720 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3721 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X3722 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3723 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3724 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3725 a_2113_38308# a_2113_38308# a_2113_38308# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X3726 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3727 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3728 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3729 a_n2810_45572# a_n2840_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3730 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3731 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3732 a_7_45899# a_n443_46116# a_n452_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3733 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3734 VDD a_13259_45724# a_22397_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3735 a_5708_44484# a_3483_46348# a_5608_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X3736 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3737 a_5732_46660# a_4817_46660# a_5385_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3738 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3739 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3740 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3741 VDD a_13507_46334# a_22765_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3742 a_11823_42460# a_15051_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=2.61 w=1 l=0.15
X3743 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3744 VSS a_22521_40055# a_22459_39145# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3745 a_13678_32519# a_21855_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3746 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3747 a_5365_45348# a_5111_44636# a_4927_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3748 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3749 a_17021_43396# a_16977_43638# a_16855_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3750 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3751 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3752 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3753 VREF_GND a_n4064_39616# C9_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3754 VDD a_7227_47204# DATA[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3755 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3756 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3757 a_7989_47542# a_n237_47217# a_7903_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3758 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3759 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3760 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3761 a_19332_42282# a_19511_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3762 VSS a_6851_47204# a_7227_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X3763 a_13607_46688# a_6755_46942# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3764 EN_VIN_BSTR_N a_18194_35068# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3765 a_4880_45572# a_526_44458# a_4808_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X3766 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3767 a_20922_43172# a_10193_42453# a_20836_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X3768 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3769 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3770 a_12978_47026# a_11901_46660# a_12816_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3771 VDD a_13720_44458# a_12607_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X3772 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3773 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3774 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3775 VDD a_2952_47436# a_2747_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3776 a_5147_45002# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3777 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3778 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3779 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3780 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3781 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3782 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3783 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3784 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3785 VDD a_14513_46634# a_14543_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3786 VDD a_21259_43561# a_16922_45042# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3787 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3788 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3789 VDD a_n4334_38528# a_n4064_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3790 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3791 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3792 VSS a_11459_47204# DATA[5] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3793 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3794 C9_N_btm a_17730_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3795 VDD a_21137_46414# a_21167_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3796 a_3905_42558# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3797 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3798 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3799 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3800 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3801 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3802 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3803 VSS a_22959_47212# a_22612_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3804 VSS a_6755_46942# a_13556_45296# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3805 a_383_46660# a_33_46660# a_288_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3806 a_n4209_38216# a_n2302_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X3807 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3808 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3809 a_17061_44734# a_11691_44458# a_16979_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3810 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3811 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3812 a_4149_42891# a_2382_45260# a_3935_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X3813 DATA[3] a_7227_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3814 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3815 VDD a_n755_45592# a_3318_42354# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X3816 VDD a_n443_46116# a_1427_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3817 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3818 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3819 VDD a_5497_46414# a_5527_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3820 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3821 a_5937_45572# a_5907_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3822 a_11323_42473# a_5742_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3823 VSS a_4921_42308# a_5755_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3824 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3825 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3826 a_n3565_39304# a_n2946_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3827 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3828 a_21076_30879# a_22959_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3829 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3830 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3831 VDD a_n2302_38778# a_n4209_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3832 VSS a_n755_45592# a_3318_42354# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X3833 VDD a_17583_46090# a_13259_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3834 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3835 a_3699_46634# a_3524_46660# a_3878_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3836 VSS a_3600_43914# a_3499_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X3837 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3838 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3839 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3840 a_17595_43084# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X3841 a_5111_44636# a_9396_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3842 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3843 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3844 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3845 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3846 a_13829_44260# a_13059_46348# a_13483_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3847 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3848 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3849 a_18341_45572# a_18175_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3850 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3851 a_9290_44172# a_13635_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3852 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3853 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3854 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3855 a_12991_46634# a_12816_46660# a_13170_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3856 VSS a_2277_45546# a_2211_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3857 a_18429_43548# a_18525_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X3858 VSS a_6453_43914# a_n2661_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X3859 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3860 a_6773_42558# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3861 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3862 a_2253_44260# a_n443_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X3863 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3864 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3865 a_9885_42558# a_7499_43078# a_9803_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3866 a_16414_43172# a_16137_43396# a_16245_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X3867 a_3726_37500# a_6886_37412# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X3868 a_2304_45348# a_n863_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X3869 a_21811_47423# SINGLE_ENDED VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3870 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3871 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3872 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3873 a_13351_46090# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X3874 VSS C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3875 a_n4064_38528# a_n4334_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X3876 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3877 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3878 a_n1435_47204# a_n1605_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3879 a_n935_46688# a_n1151_42308# a_n1021_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3880 VSS a_12549_44172# a_17639_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X3881 a_6977_45572# a_6598_45938# a_6905_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X3882 a_11530_34132# EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3883 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3884 VSS a_n1177_43370# a_n1243_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3885 VSS a_n23_44458# a_n89_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3886 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3887 VDD a_13460_43230# a_13635_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3888 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3889 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3890 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3891 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3892 VSS a_n913_45002# a_n967_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3893 VDD a_11525_45546# a_11189_46129# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X3894 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3895 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3896 VDD a_n755_45592# a_626_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3897 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3898 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3899 a_n1287_44306# a_n1331_43914# a_n1453_44318# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3900 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3901 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3902 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3903 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3904 VDD a_10227_46804# a_10768_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X3905 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3906 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3907 a_895_43940# a_644_44056# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3908 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3909 a_11136_42852# a_10922_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X3910 a_n755_45592# a_n809_44244# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3911 a_n699_43396# a_n1177_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3912 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3913 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3914 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3915 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3916 VDD a_n4334_37440# a_n4064_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3917 VDD a_8568_45546# a_8162_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3918 a_11551_42558# a_n97_42460# a_11633_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3919 a_6293_42852# a_5755_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3920 a_n2840_42826# a_n2661_42834# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3921 a_14033_45572# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X3922 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3923 VSS a_n1736_42282# a_n4318_37592# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3924 a_16131_47204# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3925 a_5289_44734# a_4223_44672# a_5205_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3926 VDD a_10083_42826# a_7499_43078# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3927 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3928 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3929 VSS a_5147_45002# a_5708_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X3930 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3931 a_768_44030# a_13487_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3932 VDD a_11415_45002# a_22591_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3933 VIN_N EN_VIN_BSTR_N C8_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3934 VSS a_6886_37412# a_4338_37500# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X3935 VDD a_13259_45724# a_14309_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X3936 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3937 a_10053_45546# a_10490_45724# a_10210_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X3938 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3939 VDD a_19332_42282# a_4190_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3940 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3941 a_n4064_40160# a_n4334_40480# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3942 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3943 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3944 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3945 a_n998_43396# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3946 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3947 a_6671_43940# a_6109_44484# a_6453_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3948 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3949 a_3090_45724# a_18911_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1468 ps=1.34 w=1 l=0.15
X3950 VSS a_18287_44626# a_18248_44752# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3951 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3952 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3953 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3954 a_n1352_43396# a_n2433_43396# a_n1699_43638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3955 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3956 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3957 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3958 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3959 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3960 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3961 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3962 VSS C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3963 VDD a_n2302_37690# a_n4209_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3964 VDD a_n2946_37984# a_n3565_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3965 a_16131_47204# a_15507_47210# a_16023_47582# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3966 a_11750_44172# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X3967 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3968 VSS a_2779_44458# a_1307_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3969 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3970 a_n23_44458# a_n356_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3971 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3972 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3973 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3974 VIN_N EN_VIN_BSTR_N C1_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X3975 a_7845_44172# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X3976 VSS a_6123_31319# a_7963_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3977 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3978 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3979 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3980 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3981 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3982 a_8560_45348# a_8746_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X3983 a_5907_46634# a_5732_46660# a_6086_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3984 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3985 a_19095_43396# a_13661_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X3986 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3987 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3988 a_21363_46634# a_21188_46660# a_21542_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3989 VSS a_n4315_30879# a_n4251_40480# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X3990 VSS a_n4064_39616# a_n2302_39866# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X3991 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3992 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3993 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3994 a_14180_46482# a_14035_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3995 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3996 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3997 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3998 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3999 a_n4064_37440# a_n4334_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X4000 a_18315_45260# a_18587_45118# a_18545_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X4001 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4002 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4003 a_8349_46414# a_8016_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X4004 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4005 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4006 VSS a_3499_42826# a_3445_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4007 a_n1532_35090# a_n1630_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4008 a_2537_44260# a_2479_44172# a_2127_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X4009 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4010 VDD a_3815_47204# a_4007_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4011 a_9306_43218# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X4012 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4013 VDD a_6667_45809# a_6598_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X4014 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4015 a_7230_45938# a_6511_45714# a_6667_45809# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X4016 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4017 VDD a_2779_44458# a_1307_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X4018 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4019 a_8685_43396# a_8147_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X4020 VDD a_1343_38525# a_1736_39043# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4021 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4022 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4023 VSS VSS a_3726_37500# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.589 pd=4.42 as=0.3135 ps=2.23 w=1.9 l=0.15
X4024 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4025 a_8270_45546# a_n237_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4026 a_3992_43940# a_768_44030# a_3737_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X4027 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4028 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4029 a_15765_45572# a_15599_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4030 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4031 a_3815_47204# a_3785_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4032 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4033 a_2063_45854# a_9863_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4034 VDD a_19431_45546# a_19418_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4035 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4036 VSS a_14021_43940# a_22959_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4037 VSS a_11415_45002# a_22591_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4038 a_6755_46942# a_15015_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X4039 a_19328_44172# a_19478_44306# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X4040 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4041 VDD a_768_44030# a_726_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4042 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4043 VSS a_10227_46804# a_14537_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4044 a_21073_44484# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X4045 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4046 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4047 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4048 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X4049 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4050 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4051 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4052 VDD a_13059_46348# a_15297_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X4053 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4054 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4055 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4056 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4057 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4058 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4059 VSS a_12465_44636# a_22223_47212# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4060 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4061 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4062 a_19164_43230# a_18083_42858# a_18817_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4063 VDD a_n1352_43396# a_n1177_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4064 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4065 VSS a_n863_45724# a_1067_42314# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4066 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4067 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4068 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4069 a_383_46660# a_n133_46660# a_288_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4070 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4071 a_13814_43218# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X4072 VSS a_9127_43156# a_9061_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4073 a_3524_46660# a_2443_46660# a_3177_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4074 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4075 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4076 VDD a_9482_43914# a_10157_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4077 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4078 VSS a_12607_44458# a_12553_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4079 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4080 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4081 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4082 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4083 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4084 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4085 VSS a_17499_43370# a_17433_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4086 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4087 VSS a_10903_43370# a_11963_45334# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4088 C1_P_btm a_1606_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4089 VSS a_14815_43914# a_14761_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4090 a_13213_44734# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4091 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4092 VDD a_12427_45724# a_10490_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X4093 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4094 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4095 VDD a_n2302_39072# a_n4209_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4096 VSS a_11323_42473# a_10807_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4097 a_12513_46660# a_12469_46902# a_12347_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X4098 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4099 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4100 VDD a_1209_43370# a_n1557_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4101 a_18989_43940# a_18451_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4102 VSS a_8667_46634# a_8601_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4103 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4104 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4105 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4106 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4107 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4108 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4109 a_2889_44172# a_2998_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X4110 VSS a_7281_43914# a_7229_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X4111 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4112 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4113 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4114 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4115 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4116 VSS a_21195_42852# a_21671_42860# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4117 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4118 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4119 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4120 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4121 VSS a_n699_43396# a_4743_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X4122 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4123 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4124 a_n3565_39590# a_n2946_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X4125 VDD a_n443_46116# a_2437_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4126 a_n2956_38680# a_n2472_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4127 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4128 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4129 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4130 a_10553_43218# a_10518_42984# a_10083_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X4131 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4132 VSS a_13635_43156# a_13569_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4133 a_16789_44484# a_14537_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4134 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4135 a_18834_46812# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X4136 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4137 a_n1151_42308# a_n1329_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X4138 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4139 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4140 a_10405_44172# a_7499_43078# a_10555_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X4141 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4142 VSS a_n2833_47464# CLK_DATA VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X4143 VSS a_18315_45260# a_18189_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X4144 a_n1917_43396# a_n2433_43396# a_n2012_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4145 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4146 a_n1441_43940# a_n2065_43946# a_n1549_44318# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4147 VDD a_17499_43370# a_17486_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4148 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4149 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4150 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4151 VDD a_22223_42860# a_22400_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4152 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4153 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4154 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4155 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4156 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4157 VDD a_3524_46660# a_3699_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4158 a_n1059_45260# a_17499_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4159 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4160 a_10765_43646# a_10695_43548# a_10057_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X4161 a_15890_42674# a_15803_42450# a_15486_42560# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X4162 VDD a_12549_44172# a_20556_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4163 VSS a_12861_44030# a_17639_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X4164 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4165 VDD a_5815_47464# a_n1613_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4166 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4167 VCM a_4958_30871# C9_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4168 a_17433_43396# a_16243_43396# a_17324_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4169 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4170 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4171 a_11827_44484# a_3232_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4172 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4173 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4174 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4175 a_1847_42826# a_2351_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4176 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4177 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4178 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4179 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4180 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4181 VSS a_6151_47436# a_14955_47212# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4182 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4183 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4184 a_20205_31679# a_22223_46124# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4185 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4186 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4187 VSS a_15227_44166# a_15785_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4188 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4189 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4190 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4191 VDD a_8667_46634# a_8654_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4192 a_n452_45724# a_n443_46116# a_n310_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4193 VDD a_1239_47204# a_1431_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4194 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4195 a_700_44734# a_n746_45260# a_327_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X4196 a_19862_44208# a_13747_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4197 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4198 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4199 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4200 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4201 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4202 a_10775_45002# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X4203 a_1115_44172# a_453_43940# a_1443_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4204 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4205 a_3232_43370# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4206 VDD a_22959_44484# a_19237_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4207 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4208 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4209 a_n3690_38528# a_n3674_38680# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4210 a_484_44484# a_n863_45724# a_327_44734# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X4211 VDD a_14543_43071# a_13291_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4212 VSS a_12549_44172# a_21205_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X4213 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4214 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4215 a_20512_43084# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4216 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4217 a_20256_43172# a_20202_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.203125 ps=1.275 w=0.65 l=0.15
X4218 a_6761_42308# a_n913_45002# a_6773_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4219 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4220 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4221 a_n2840_42282# a_n2661_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4222 a_6298_44484# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4223 VDD a_19864_35138# a_21589_35634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4224 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4225 a_n2661_46098# a_1983_46706# a_2162_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4226 VDD a_8685_43396# a_14955_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X4227 VSS a_15368_46634# a_15312_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4228 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4229 a_5429_46660# a_5385_46902# a_5263_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X4230 VDD a_16855_45546# a_16842_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4231 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4232 a_1221_42558# a_1184_42692# a_1149_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X4233 VSS a_5815_47464# a_n1613_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4234 a_11315_46155# a_11133_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4235 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4236 a_16522_42674# a_15803_42450# a_15959_42545# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X4237 a_n923_35174# EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X4238 a_20885_46660# a_20841_46902# a_20719_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X4239 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4240 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4241 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4242 a_14456_42282# a_14635_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4243 a_20719_45572# a_20273_45572# a_20623_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4244 a_1756_43548# a_1307_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X4245 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4246 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4247 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4248 a_n2472_42826# a_n2293_42834# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4249 a_7276_45260# a_6709_45028# a_7418_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4250 VDD a_1823_45246# a_3232_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4251 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4252 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4253 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4254 VDD a_22400_42852# a_22521_40055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4255 a_n4315_30879# a_n2302_40160# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4256 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4257 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4258 VSS a_3422_30871# a_22315_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4259 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4260 VDD a_10341_42308# a_11554_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X4261 a_n2497_47436# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4262 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4263 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4264 a_3260_45572# a_3218_45724# a_2957_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X4265 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4266 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4267 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4268 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4269 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4270 a_11280_45822# a_2063_45854# a_10907_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X4271 a_603_45572# a_310_45028# a_509_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X4272 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4273 a_8746_45002# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4274 a_15002_46116# a_13925_46122# a_14840_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4275 a_2479_44172# a_2905_42968# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X4276 a_11064_45572# a_10903_43370# a_10907_45822# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X4277 a_n906_45572# a_n971_45724# a_n1013_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X4278 a_21205_44306# a_20935_43940# a_21115_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X4279 a_12861_44030# a_18143_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4280 VDD a_n2840_46090# a_n2956_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4281 DATA[3] a_7227_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X4282 VDD a_6945_45028# a_22223_46124# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4283 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4284 a_13556_45296# a_6755_46942# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4285 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4286 VSS C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4287 VCM a_7174_31319# C0_dummy_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4288 VDD a_8199_44636# a_9377_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X4289 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4290 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4291 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4292 a_n4334_39392# a_n4318_39304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4293 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X4294 a_12710_44260# a_10903_43370# a_12603_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X4295 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4296 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4297 a_13777_45326# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4298 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4299 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4300 a_16522_42674# a_15764_42576# a_15959_42545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X4301 a_14205_43396# a_13667_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X4302 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4303 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4304 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4305 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4306 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4307 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4308 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4309 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4310 a_6419_46155# a_5807_45002# a_6419_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4311 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4312 VDD a_5732_46660# a_5907_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4313 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4314 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4315 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4316 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4317 a_n2860_39866# a_n2956_39768# a_n2946_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X4318 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4319 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X4320 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4321 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4322 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4323 a_18533_44260# a_18326_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4324 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4325 VDD a_13556_45296# a_13857_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4326 a_5066_45546# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4327 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4328 w_1575_34946# a_n923_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X4329 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4330 a_n901_46420# a_n1076_46494# a_n722_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X4331 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4332 VSS a_11599_46634# a_18175_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4333 a_12861_44030# a_18143_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4334 VSS a_13635_43156# a_9290_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4335 VSS a_11599_46634# a_18819_46122# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4336 VDD a_n1630_35242# a_18194_35068# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4337 a_n3690_37440# a_n3674_37592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4338 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4339 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4340 VSS a_n3690_39616# a_n3420_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4341 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4342 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4343 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4344 a_n2442_46660# a_n2472_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4345 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4346 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4347 VSS a_n1435_47204# a_13487_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X4348 VDD a_3147_46376# a_526_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X4349 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4350 a_8317_43396# a_n755_45592# a_8229_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X4351 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4352 a_n3674_38216# a_n2104_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4353 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4354 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4355 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4356 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4357 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4358 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4359 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4360 a_n2312_40392# a_n2288_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4361 VSS a_22591_44484# a_17730_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4362 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4363 VDD a_21589_35634# SMPL_ON_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4364 VDD a_n1079_45724# a_n1099_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X4365 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4366 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4367 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4368 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4369 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4370 a_n914_42852# a_n1991_42858# a_n1076_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4371 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4372 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4373 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4374 a_n97_42460# a_19700_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4375 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4376 VDD a_n809_44244# a_n755_45592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X4377 a_3877_44458# a_3699_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X4378 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4379 a_n913_45002# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4380 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4381 a_15368_46634# a_15143_45578# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X4382 a_11206_38545# CAL_N a_4338_37500# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X4383 a_4905_42826# a_5379_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4384 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4385 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4386 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4387 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4388 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4389 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4390 VSS a_10467_46802# a_10428_46928# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4391 VSS a_3147_46376# a_526_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X4392 VDD a_n4334_40480# a_n4064_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4393 a_9313_45822# a_9049_44484# a_9159_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4394 a_21145_44484# a_20766_44850# a_21073_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X4395 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4396 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4397 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4398 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4399 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4400 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4401 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4402 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4403 VSS a_22521_40599# a_22717_37285# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X4404 VDD a_2324_44458# a_15682_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4405 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4406 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4407 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4408 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4409 VSS a_2680_45002# a_2274_45254# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X4410 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4411 a_10768_47026# a_10554_47026# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X4412 VSS C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4413 VSS a_21671_42860# a_3422_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4414 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4415 a_5837_45028# a_5807_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X4416 C0_dummy_P_btm a_7174_31319# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4417 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4418 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4419 a_n785_47204# a_n815_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4420 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4421 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4422 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4423 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4424 a_14537_43396# a_14358_43442# a_14621_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X4425 a_n1736_43218# a_n1853_43023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X4426 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4427 a_n3565_38216# a_n2946_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4428 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4429 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4430 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4431 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4432 a_16877_42852# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4433 a_6640_46482# a_5257_43370# a_6419_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4434 VDD a_3090_45724# a_17786_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X4435 a_15493_43396# a_14955_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X4436 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4437 a_9823_46482# a_9569_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X4438 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4439 VDD a_14021_43940# a_22959_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4440 VDD a_n3420_38528# a_n2860_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X4441 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4442 VSS a_10227_46804# a_12513_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4443 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4444 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4445 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4446 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4447 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4448 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4449 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4450 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4451 VDD a_3483_46348# a_17061_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4452 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4453 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4454 VSS a_17339_46660# a_19095_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4455 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4456 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4457 VSS a_n1532_35090# a_n83_35174# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X4458 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4459 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4460 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4461 a_3699_46348# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X4462 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4463 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4464 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4465 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4466 VSS a_10533_42308# a_10723_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4467 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4468 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4469 a_18214_42558# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X4470 VSS a_3537_45260# a_4223_44672# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4471 VSS a_n1630_35242# a_n1532_35090# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4472 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4473 VSS a_14537_43396# a_14180_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X4474 a_16501_45348# a_10193_42453# a_16405_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4475 VSS a_21259_43561# a_16922_45042# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4476 VSS a_15743_43084# a_15567_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4477 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4478 VDD a_22821_38993# a_22521_39511# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4479 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4480 VSS a_n2840_46634# a_n2956_39768# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4481 a_9049_44484# a_8701_44490# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X4482 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4483 VDD a_2382_45260# a_3737_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4484 VDD a_n967_45348# a_n961_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4485 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4486 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4487 a_19615_44636# a_12861_44030# a_19789_44512# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X4488 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4489 a_9863_46634# a_10150_46912# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X4490 VDD a_n881_46662# a_n745_45366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X4491 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4492 a_n2109_45247# a_n2017_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4493 VDD a_21496_47436# a_13507_46334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X4494 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4495 VSS a_n143_45144# a_n37_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4496 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4497 a_19418_45938# a_18341_45572# a_19256_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4498 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4499 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4500 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4501 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4502 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4503 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4504 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4505 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4506 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4507 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4508 VDD a_n2438_43548# a_n2433_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4509 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4510 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4511 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4512 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4513 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4514 VDD a_5907_45546# a_5937_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X4515 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4516 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4517 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4518 C5_P_btm a_n4209_38502# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X4519 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4520 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4521 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4522 VSS a_n452_44636# a_n2129_44697# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4523 a_n4318_38680# a_n2472_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4524 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4525 a_n2472_42282# a_n2293_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4526 a_5608_44484# a_5111_44636# a_5518_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X4527 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4528 VDD a_742_44458# a_700_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X4529 VDD a_n901_43156# a_n443_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X4530 VSS a_7287_43370# a_7221_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4531 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4532 VSS a_768_44030# a_13720_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4533 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4534 a_n89_44484# a_n467_45028# a_n452_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4535 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4536 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4537 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4538 a_2609_46660# a_2443_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4539 VDD a_9290_44172# a_9801_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X4540 VSS a_n1613_43370# a_6809_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4541 VDD a_327_47204# DATA[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4542 a_n4064_39616# a_n4334_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4543 a_556_44484# a_526_44458# a_484_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X4544 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4545 VDD a_n4334_39392# a_n4064_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4546 VDD a_2324_44458# a_15682_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4547 VSS a_4007_47204# DATA[2] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4548 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4549 a_2112_39137# a_1343_38525# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4550 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4551 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4552 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4553 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4554 VSS a_19328_44172# a_19279_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
X4555 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4556 VDD a_n3420_37440# a_n2860_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X4557 a_n3420_38528# a_n3690_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X4558 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4559 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X4560 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4561 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4562 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4563 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4564 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4565 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4566 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4567 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4568 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4569 a_13887_32519# a_22223_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4570 a_11387_46155# a_n1151_42308# a_11315_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4571 a_10341_43396# a_9803_43646# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4572 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4573 a_10554_47026# a_10467_46802# a_10150_46912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X4574 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4575 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4576 VSS a_16137_43396# a_18548_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X4577 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4578 C0_P_btm a_n3420_37440# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4579 VSS a_10227_46804# a_20885_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4580 VIN_P EN_VIN_BSTR_P C2_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X4581 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4582 a_n452_45724# a_n743_46660# a_n310_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4583 a_11682_45822# a_11652_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X4584 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4585 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4586 a_n443_42852# a_n901_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4587 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4588 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4589 VDD a_n2472_46090# a_n2956_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4590 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X4591 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4592 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4593 VSS a_13747_46662# a_14495_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X4594 VDD a_10809_44734# a_n2661_42834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4595 C0_dummy_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X4596 VDD a_11322_45546# a_11280_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X4597 VSS a_n1329_42308# a_n1151_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4598 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4599 VSS a_n4209_39590# a_n4251_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X4600 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4601 VDD a_n2302_39072# a_n4209_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4602 a_5649_42852# a_5111_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4603 VDD a_18479_47436# a_13747_46662# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X4604 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4605 a_3381_47502# a_2905_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X4606 VSS a_n746_45260# a_261_44278# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4607 VDAC_P C1_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4608 VSS a_n913_45002# a_8325_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4609 a_17486_43762# a_16409_43396# a_17324_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4610 a_11136_45572# a_3483_46348# a_11064_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X4611 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4612 VSS a_13249_42308# a_13904_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X4613 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4614 VSS a_1307_43914# a_2675_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4615 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4616 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4617 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4618 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4619 VSS a_n1532_35090# a_n923_35174# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X4620 VSS a_13259_45724# a_14797_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X4621 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4622 VSS a_2324_44458# a_949_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4623 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4624 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4625 a_3699_46634# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4626 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4627 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4628 VIN_N EN_VIN_BSTR_N C9_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X4629 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4630 a_20841_45814# a_20623_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4631 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4632 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4633 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4634 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4635 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4636 a_10341_42308# a_9803_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X4637 a_17639_46660# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4638 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4639 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4640 a_16327_47482# a_17591_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4641 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4642 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4643 VSS a_2324_44458# a_15682_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4644 a_20397_44484# a_20362_44736# a_20159_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X4645 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4646 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4647 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4648 a_1260_45572# a_n755_45592# a_1176_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X4649 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4650 a_12991_46634# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4651 a_n4064_39072# a_n4334_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X4652 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4653 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4654 a_518_46155# a_472_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4655 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4656 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4657 VDD a_20841_45814# a_20731_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4658 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4659 a_9751_46155# a_9569_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4660 a_1443_43940# a_1414_42308# a_1241_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4661 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=0.35
X4662 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4663 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4664 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4665 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4666 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4667 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4668 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4669 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4670 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4671 DATA[1] a_1431_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4672 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4673 VDD a_11823_42460# a_14033_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X4674 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4675 COMP_P a_1239_39587# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4676 VSS a_n2840_42826# a_n3674_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4677 VSS a_3537_45260# a_5365_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X4678 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4679 a_21589_35634# a_19864_35138# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4680 a_3065_45002# a_3318_42354# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X4681 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4682 C8_P_btm a_n3420_39616# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4683 a_n310_45899# a_n356_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4684 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4685 VDD a_22591_46660# a_20820_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4686 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4687 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4688 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4689 a_16327_47482# a_17591_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4690 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4691 a_n3420_37440# a_n3690_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X4692 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4693 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4694 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4695 a_8337_42558# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4696 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4697 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4698 VDD a_n1331_43914# a_n1441_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4699 VDD a_4646_46812# a_7411_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4700 VSS a_3877_44458# a_2382_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4701 w_11334_34010# a_18194_35068# EN_VIN_BSTR_N w_11334_34010# sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X4702 a_11186_47026# a_10428_46928# a_10623_46897# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X4703 a_20273_46660# a_20107_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4704 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4705 VDD a_10835_43094# a_10796_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4706 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4707 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4708 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4709 VSS a_12883_44458# a_12829_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4710 a_11341_43940# a_10729_43914# a_11257_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3925 pd=1.785 as=0.135 ps=1.27 w=1 l=0.15
X4711 VSS a_564_42282# a_n1630_35242# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4712 VSS a_5066_45546# a_9159_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4713 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4714 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4715 a_12549_44172# a_20567_45036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4716 VDD a_14456_42282# a_5342_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4717 VDD a_2063_45854# a_10809_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4718 VDD a_10227_46804# a_16104_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X4719 a_645_46660# a_601_46902# a_479_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X4720 VDD a_2127_44172# a_n2661_45010# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X4721 a_n2840_46090# a_n2661_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4722 a_5088_37509# VSS VDAC_Ni VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X4723 a_12861_44030# a_18143_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X4724 a_14513_46634# a_14180_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4725 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4726 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4727 VREF_GND a_17730_32519# C9_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4728 a_14635_42282# a_n913_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4729 a_21137_46414# a_19692_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4730 a_1609_45822# a_167_45260# a_1609_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4731 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4732 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4733 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4734 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4735 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4736 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4737 a_10544_45572# a_10490_45724# a_10053_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X4738 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4739 a_10555_44260# a_10949_43914# a_10405_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.13325 ps=1.06 w=0.65 l=0.15
X4740 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4741 C2_P_btm a_n3565_38216# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X4742 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X4743 a_8952_43230# a_7871_42858# a_8605_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4744 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4745 VSS a_1431_47204# DATA[1] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4746 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4747 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4748 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4749 VDD a_1736_39587# a_1239_39587# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4750 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4751 a_9377_42558# a_8685_42308# a_9293_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4752 a_3067_47026# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X4753 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4754 a_4190_30871# a_19332_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4755 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4756 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4757 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4758 a_15861_45028# a_15595_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X4759 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4760 VDD a_9067_47204# DATA[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4761 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4762 a_13720_44458# a_9482_43914# a_14112_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X4763 a_n1352_43396# a_n2267_43396# a_n1699_43638# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4764 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4765 a_16245_42852# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X4766 a_6469_45572# a_5907_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X4767 VSS a_n357_42282# a_6101_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4768 a_15194_46482# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X4769 a_15493_43940# a_14955_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4770 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4771 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4772 a_20692_30879# a_22959_46124# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4773 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4774 VSS a_n2302_37984# a_n4209_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4775 a_5497_46414# a_5164_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4776 VSS a_104_43370# a_n971_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4777 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4778 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4779 a_5907_46634# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4780 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4781 a_3177_46902# a_2959_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4782 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4783 VREF_GND a_13258_32519# C0_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4784 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4785 VDD a_4743_44484# a_4791_45118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4786 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4787 a_19700_43370# a_18579_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4788 a_12861_44030# a_18143_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X4789 a_21363_46634# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4790 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4791 VSS a_n443_42852# a_15940_43402# VSS sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X4792 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4793 a_12427_45724# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.14075 ps=1.325 w=0.42 l=0.15
X4794 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4795 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4796 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4797 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4798 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4799 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4800 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4801 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4802 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4803 VSS a_n3690_39616# a_n3420_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X4804 VDAC_N C3_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4805 a_5891_43370# a_9127_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4806 a_n1920_47178# a_n1741_47186# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X4807 a_10903_43370# a_13351_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4808 a_n955_45028# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4809 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4810 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4811 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4812 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4813 VDD a_n357_42282# a_7309_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4814 a_4185_45028# a_3065_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4815 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4816 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4817 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4818 VDD a_3147_46376# a_526_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4819 a_18596_45572# a_18479_45785# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4820 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4821 VSS a_22775_42308# a_22465_38105# VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4822 a_16137_43396# a_15781_43660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X4823 a_6575_47204# a_6545_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4824 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4825 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4826 a_4649_42852# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X4827 VSS a_n2472_46634# a_n2442_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4828 VSS a_2711_45572# a_20107_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4829 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4830 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4831 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4832 VSS a_n2104_42282# a_n3674_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4833 VIN_N EN_VIN_BSTR_N a_11530_34132# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X4834 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4835 VSS a_15015_46420# a_14949_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4836 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4837 VSS a_5691_45260# a_n2109_47186# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4838 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4839 a_17730_32519# a_22591_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4840 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4841 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4842 a_3600_43914# a_1307_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X4843 a_17583_46090# a_17715_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X4844 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4845 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4846 a_13925_46122# a_13759_46122# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4847 VDD a_n901_43156# a_n914_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4848 VDD a_1239_39043# comp_n VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4849 a_8191_45002# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4850 a_n310_44484# a_n356_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4851 a_21125_42558# a_18597_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4852 VDD a_22959_46124# a_20692_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4853 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4854 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4855 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4856 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4857 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4858 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4859 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4860 VSS a_14543_43071# a_13291_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4861 a_5932_42308# a_5755_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4862 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4863 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4864 VDD a_1307_43914# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4865 VSS a_3147_46376# a_526_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4866 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4867 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4868 VDD a_n2946_38778# a_n3565_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4869 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4870 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4871 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4872 VDD a_16112_44458# a_14673_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X4873 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4874 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4875 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4876 a_n1641_46494# a_n1991_46122# a_n1736_46482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4877 a_3175_45822# a_3316_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4878 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4879 VSS a_16763_47508# a_5807_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4880 VREF a_20447_31679# C5_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X4881 a_14226_46660# a_14180_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4882 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4883 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4884 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4885 VDD a_13348_45260# a_13159_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X4886 a_n4209_39590# a_n2302_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X4887 VDD a_6491_46660# a_6851_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4888 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4889 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4890 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4891 VDD a_22775_42308# a_22465_38105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4892 a_6511_45714# a_4646_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4893 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4894 a_3422_30871# a_21671_42860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4895 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4896 VDD a_2889_44172# a_413_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X4897 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4898 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4899 VSS a_16763_47508# a_16697_47582# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4900 VSS a_n443_42852# a_1755_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4901 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4902 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4903 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4904 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4905 a_10405_44172# a_10729_43914# a_10651_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4906 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4907 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4908 a_n2840_45546# a_n2661_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X4909 a_14401_32519# a_22223_43948# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4910 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4911 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4912 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4913 VREF a_21076_30879# C8_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4914 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4915 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4916 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4917 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4918 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4919 a_4558_45348# a_4574_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4920 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4921 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4922 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4923 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4924 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4925 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4926 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4927 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4928 a_5193_42852# a_3905_42865# a_5111_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4929 a_18143_47464# a_18479_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X4930 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4931 a_10533_42308# a_n913_45002# a_10545_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4932 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4933 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4934 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4935 VDD a_16721_46634# a_16751_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4936 a_18909_45814# a_18691_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4937 a_n2840_45002# a_n2661_45010# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X4938 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4939 a_948_46660# a_n133_46660# a_601_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4940 a_117_45144# a_n443_42852# a_45_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X4941 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4942 a_11415_45002# a_13249_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4943 a_3699_46348# a_3877_44458# a_3873_46454# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X4944 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4945 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4946 a_n4209_38502# a_n2302_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X4947 a_15681_43442# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4948 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4949 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4950 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=10
X4951 VDD a_n1059_45260# a_18727_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X4952 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4953 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4954 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4955 a_n4251_38304# a_n4318_38216# a_n4334_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X4956 VSS a_5013_44260# a_5663_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4957 a_9801_43940# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X4958 a_22521_39511# a_22545_38993# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X4959 VSS a_10193_42453# a_18797_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4960 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4961 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4962 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4963 a_19789_44512# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X4964 VDD a_18057_42282# a_n356_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X4965 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4966 a_2779_44458# a_1423_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X4967 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4968 a_13113_42826# a_12895_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4969 a_16197_42308# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X4970 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4971 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4972 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4973 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4974 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4975 VDD a_8034_45724# a_n1925_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X4976 VDD a_11691_44458# a_11649_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4977 a_15761_42308# a_15051_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X4978 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4979 a_n3690_39392# a_n3674_39304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4980 VSS a_1568_43370# a_1512_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4981 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4982 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4983 a_16680_45572# a_15765_45572# a_16333_45814# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4984 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4985 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4986 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4987 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4988 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4989 VDD a_5066_45546# a_5024_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X4990 VSS a_n809_44244# a_n875_44318# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4991 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4992 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4993 VDD a_n2946_37690# a_n3565_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4994 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4995 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4996 a_10518_42984# a_10796_42968# a_10752_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X4997 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4998 a_n2267_43396# a_n2433_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4999 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5000 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5001 a_8189_46660# a_8145_46902# a_8023_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X5002 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5003 VDD a_1123_46634# a_584_46384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X5004 VSS a_n4064_39072# a_n2302_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X5005 VDD a_13661_43548# a_14976_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X5006 a_11691_44458# a_5807_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5007 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5008 VSS a_5891_43370# a_5837_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5009 a_20062_46116# a_18985_46122# a_19900_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5010 a_20269_44172# a_20365_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X5011 VSS a_n2472_42826# a_n4318_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5012 a_18707_42852# a_18083_42858# a_18599_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5013 VSS a_7754_38470# a_7754_38470# VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X5014 VDD a_327_47204# DATA[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5015 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5016 a_n784_42308# a_n961_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5017 a_12638_46436# a_13059_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5018 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X5019 a_13157_43218# a_13113_42826# a_12991_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X5020 VSS a_4007_47204# DATA[2] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5021 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5022 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5023 VDD a_15015_46420# a_15002_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5024 VDD a_16327_47482# a_20159_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5025 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5026 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X5027 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5028 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5029 VSS a_n785_47204# a_327_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X5030 a_18834_46812# a_13661_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X5031 a_n2840_45546# a_n2661_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5032 VSS a_21177_47436# a_20990_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X5033 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5034 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5035 a_n3420_38528# a_n3690_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5036 VSS a_7499_43078# a_11816_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5037 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5038 a_6761_42308# a_3537_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5039 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5040 VSS C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5041 a_10623_46897# a_10428_46928# a_10933_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X5042 a_5263_45724# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X5043 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5044 VDD a_11823_42460# a_11322_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5045 VSS a_5111_44636# a_8018_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5046 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5047 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5048 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5049 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5050 a_3357_43084# a_4905_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5051 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5052 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5053 a_7903_47542# a_n237_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X5054 VSS a_8667_46634# a_n237_47217# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5055 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5056 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5057 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5058 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5059 a_n2472_46090# a_n2293_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5060 VREF a_19237_31679# C0_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X5061 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5062 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5063 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5064 VCM a_5742_30871# C6_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X5065 VDD a_n901_43156# a_n443_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5066 a_10249_46116# a_9823_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X5067 a_2684_37794# VDAC_Pi a_2113_38308# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X5068 VSS a_22959_46660# a_21076_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5069 VDD a_10775_45002# a_10180_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X5070 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5071 a_n4209_37414# a_n2302_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X5072 a_13467_32519# a_21487_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5073 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5074 a_8696_44636# a_16855_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X5075 a_6633_46155# a_5807_45002# a_6419_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X5076 a_n2661_42834# a_8975_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5077 a_n1243_43396# a_n2433_43396# a_n1352_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5078 a_7274_43762# a_6197_43396# a_7112_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5079 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5080 a_10922_42852# a_10835_43094# a_10518_42984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X5081 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5082 VDD a_5807_45002# a_11691_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5083 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5084 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5085 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5086 DATA[0] a_327_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5087 a_n1917_43396# a_n2267_43396# a_n2012_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5088 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5089 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5090 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5091 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5092 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5093 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5094 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5095 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5096 a_n4209_38502# a_n2302_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5097 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5098 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5099 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5100 VSS RST_Z a_14311_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5101 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5102 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5103 a_18285_46348# a_18834_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5104 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5105 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5106 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5107 a_16327_47482# a_17591_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X5108 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5109 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5110 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5111 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5112 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5113 VSS a_18443_44721# a_18374_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X5114 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5115 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5116 a_18597_46090# a_19431_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X5117 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5118 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5119 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5120 VSS a_8199_44636# a_10951_45334# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5121 a_7735_45067# a_6709_45028# a_7276_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X5122 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5123 a_1176_45572# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X5124 C8_P_btm a_5342_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5125 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5126 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5127 VSS a_n1838_35608# SMPL_ON_P VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5128 a_n3565_39304# a_n2946_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X5129 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5130 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5131 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=0.35
X5132 DATA[4] a_9067_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X5133 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5134 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5135 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5136 a_n1076_43230# a_n1991_42858# a_n1423_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5137 VSS a_n2109_45247# en_comp VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5138 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5139 DATA[1] a_1431_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X5140 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5141 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5142 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5143 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5144 a_13348_45260# a_13556_45296# a_13490_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5145 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5146 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5147 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5148 a_n2302_40160# a_n2312_40392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5149 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5150 VSS a_21356_42826# a_n357_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5151 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5152 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5153 VDD a_11453_44696# a_22959_47212# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X5154 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5155 VSS a_8696_44636# a_8701_44490# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5156 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5157 VSS a_15037_45618# a_15143_45578# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5158 a_3878_46660# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X5159 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5160 a_626_44172# a_n863_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5161 a_2277_45546# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X5162 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5163 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5164 a_18479_45785# a_19268_43646# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.3275 ps=1.655 w=1 l=0.15
X5165 a_16327_47482# a_17591_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X5166 a_20273_45572# a_20107_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5167 a_n3420_37440# a_n3690_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5168 VSS a_n443_42852# a_742_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5169 VSS a_n901_43156# a_n967_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X5170 a_10555_44260# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X5171 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5172 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5173 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5174 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5175 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5176 a_20820_30879# a_22591_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5177 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5178 a_17364_32525# a_22959_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5179 VSS a_13076_44458# a_12883_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X5180 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5181 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5182 a_685_42968# a_n443_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5183 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5184 a_11633_42558# a_9290_44172# a_11551_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5185 a_13170_46660# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X5186 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5187 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5188 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5189 a_20731_45938# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X5190 VDD a_4791_45118# a_6633_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X5191 a_19700_43370# a_18579_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5192 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5193 a_2382_45260# a_3877_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5194 VDD a_11599_46634# a_20107_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5195 a_16751_45260# a_17023_45118# a_16981_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5196 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5197 VSS a_13487_47204# a_768_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5198 a_11257_43940# a_10807_43548# a_11173_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5199 a_12829_44484# a_12741_44636# a_n2293_43922# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5200 VCM a_6123_31319# C4_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X5201 a_5342_30871# a_14456_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5202 VDD a_5937_45572# a_8034_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5203 VSS a_14084_46812# a_14035_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X5204 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5205 a_17639_46660# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X5206 a_10809_44734# a_10057_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5207 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5208 VDD a_11823_42460# a_14853_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5209 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5210 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5211 a_20749_43396# a_20974_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5212 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5213 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5214 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5215 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5216 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5217 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5218 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5219 a_19511_42282# a_n913_45002# a_21125_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5220 VDD a_11967_42832# a_16243_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5221 a_17517_44484# a_16979_44734# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X5222 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5223 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5224 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5225 a_1609_45572# a_n443_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5226 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5227 VSS a_1431_47204# DATA[1] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5228 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5229 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5230 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5231 a_20075_46420# a_19900_46494# a_20254_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5232 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5233 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5234 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5235 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5236 VDD a_10083_42826# a_7499_43078# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5237 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5238 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5239 a_n4209_37414# a_n2302_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5240 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5241 a_16020_45572# a_15903_45785# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X5242 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5243 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5244 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5245 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5246 a_20731_45938# a_20107_45572# a_20623_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5247 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5248 VDD a_n3420_39072# a_n2860_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X5249 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5250 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5251 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5252 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5253 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5254 a_16855_45546# a_16680_45572# a_17034_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5255 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5256 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5257 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5258 VSS a_22731_47423# a_13717_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5259 a_18114_32519# a_22223_45036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5260 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5261 VSS a_18429_43548# a_16823_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X5262 VSS a_n4334_38304# a_n4064_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5263 VSS a_8325_42308# a_8791_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5264 a_17339_46660# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5265 a_n2472_45546# a_n2293_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5266 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5267 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5268 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5269 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5270 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5271 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5272 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5273 VDD a_n4334_38528# a_n4064_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5274 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5275 VSS a_768_44030# a_13076_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X5276 VSS a_12861_44030# a_19692_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5277 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5278 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5279 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5280 VDD a_14495_45572# a_n881_46662# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5281 a_18596_45572# a_18479_45785# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X5282 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5283 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5284 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5285 a_n2472_45002# a_n2293_45010# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5286 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5287 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5288 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5289 a_3445_43172# a_3357_43084# a_n2293_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5290 a_5326_44056# a_5147_45002# a_5244_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5291 VSS a_22959_42860# a_14097_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5292 VDD a_n881_46662# a_6431_45366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X5293 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5294 a_13003_42852# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X5295 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5296 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5297 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5298 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5299 VSS a_9127_43156# a_5891_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5300 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5301 a_3503_45724# a_3775_45552# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5302 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5303 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5304 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5305 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5306 C6_N_btm a_14401_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X5307 a_3540_43646# a_584_46384# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5308 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5309 VSS a_n2302_37984# a_n4209_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5310 a_19929_45028# a_19778_44110# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5311 VDD a_167_45260# a_117_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5312 DATA[4] a_9067_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5313 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5314 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5315 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5316 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5317 a_3147_46376# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X5318 a_6086_46660# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X5319 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5320 a_n1533_46116# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X5321 VSS a_n3565_38216# a_n3607_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X5322 a_5337_42558# a_5267_42460# a_4905_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X5323 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X5324 a_21542_46660# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X5325 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5326 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5327 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5328 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5329 comp_n a_1239_39043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5330 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5331 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5332 a_10216_45572# a_10180_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X5333 a_3626_43646# a_3232_43370# a_3457_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5334 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5335 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5336 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5337 a_4699_43561# a_3080_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5338 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5339 a_1067_42314# a_1184_42692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5340 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5341 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5342 VDD a_21613_42308# a_22775_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5343 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5344 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5345 a_n4064_37984# a_n4334_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X5346 a_16269_42308# a_15890_42674# a_16197_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X5347 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5348 VDD a_5937_45572# a_6945_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5349 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5350 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5351 a_22545_38993# a_22459_39145# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5352 a_21356_42826# a_21381_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5353 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5354 VDD CLK a_8953_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5355 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5356 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5357 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5358 VDD a_2324_44458# a_949_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5359 a_n1549_44318# a_n2065_43946# a_n1644_44306# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5360 VSS a_19862_44208# a_19808_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5361 VSS a_n3690_39392# a_n3420_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5362 VDD a_1307_43914# a_16237_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5363 VDD a_5891_43370# a_8791_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5364 a_20256_43172# a_18494_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X5365 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X5366 VREF_GND a_13887_32519# C3_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X5367 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5368 a_n3420_39072# a_n3690_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X5369 a_7927_46660# a_7411_46660# a_7832_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5370 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5371 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5372 a_n2472_45546# a_n2293_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5373 VSS C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5374 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5375 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5376 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5377 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5378 C9_P_btm a_n4064_39616# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5379 a_4649_42852# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5380 a_17668_45572# a_n881_46662# a_17568_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X5381 VSS a_15493_43396# a_19478_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5382 a_16664_43396# a_16547_43609# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X5383 VDD a_6511_45714# a_6472_45840# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5384 a_6540_46812# a_3877_44458# a_6682_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5385 VDD a_5068_46348# a_4955_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X5386 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5387 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5388 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5389 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5390 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5391 a_9159_44484# a_5883_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X5392 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5393 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5394 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5395 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5396 VSS a_10341_43396# a_22591_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5397 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5398 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5399 VDD a_n4334_37440# a_n4064_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5400 VSS a_17124_42282# a_4958_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5401 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5402 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5403 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5404 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5405 C8_P_btm a_n3565_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5406 a_5267_42460# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X5407 a_n1545_46494# a_n1991_46122# a_n1641_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5408 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5409 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5410 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5411 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5412 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5413 a_1138_42852# a_791_42968# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X5414 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5415 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5416 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5417 a_n4318_40392# a_n2840_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5418 a_n1644_44306# a_n1761_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X5419 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5420 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5421 VDD a_7754_40130# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.5
X5422 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5423 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5424 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5425 a_5267_42460# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X5426 VDD a_1609_45822# a_n2293_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X5427 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5428 VREF_GND a_17364_32525# C7_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X5429 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X5430 a_2127_44172# a_2675_43914# a_2455_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5431 a_11787_45002# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X5432 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5433 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5434 VDD a_17499_43370# a_n1059_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5435 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5436 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5437 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5438 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5439 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5440 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5441 a_n2946_37984# a_n2956_38216# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5442 VSS a_19333_46634# a_19123_46287# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5443 a_3316_45546# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X5444 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5445 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5446 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5447 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5448 VSS a_13777_45326# a_13711_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5449 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5450 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5451 a_20712_42282# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5452 VSS C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5453 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5454 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5455 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5456 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5457 a_20573_43172# a_20512_43084# a_20256_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X5458 a_19479_31679# a_22223_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5459 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5460 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5461 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5462 a_n2293_46634# a_14673_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5463 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X5464 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5465 a_n1177_43370# a_n1352_43396# a_n998_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5466 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5467 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5468 VSS a_526_44458# a_5457_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X5469 a_33_46660# a_n133_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5470 VDD a_10903_43370# a_10849_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X5471 VDD a_7754_40130# a_7754_40130# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X5472 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5473 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5474 a_584_46384# a_1123_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5475 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5476 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5477 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5478 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X5479 a_8495_42852# a_7871_42858# a_8387_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5480 a_5495_43940# a_5244_44056# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X5481 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5482 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5483 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5484 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5485 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5486 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5487 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5488 a_16842_45938# a_15765_45572# a_16680_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5489 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5490 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5491 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5492 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5493 VDD a_2779_44458# a_1307_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5494 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5495 VSS a_n961_42308# a_n784_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5496 VDD a_167_45260# a_2521_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X5497 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5498 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5499 VSS a_13259_45724# a_17303_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5500 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5501 a_22780_40945# COMP_P a_22521_40599# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5502 a_17538_32519# a_22959_43948# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5503 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5504 VDD a_5937_45572# a_5829_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X5505 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5506 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5507 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5508 a_5742_30871# a_10723_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5509 a_9801_43940# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5510 a_21496_47436# a_4883_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5511 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5512 a_11816_44260# a_11750_44172# a_10729_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5513 VDD a_15051_42282# a_11823_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5514 a_2123_42473# a_n784_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5515 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5516 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5517 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5518 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5519 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5520 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5521 a_13565_43940# a_12891_46348# a_13483_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5522 VSS a_n1630_35242# a_18194_35068# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5523 a_7227_42852# a_n97_42460# a_7309_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X5524 VDD a_13747_46662# a_13607_46688# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X5525 a_n1655_44484# a_n1699_44726# a_n1821_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X5526 a_5257_43370# a_5907_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X5527 a_1667_45002# a_1823_45246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X5528 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5529 a_n2293_46098# a_5663_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X5530 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5531 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5532 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5533 a_13003_42852# a_12379_42858# a_12895_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5534 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5535 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5536 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5537 a_2711_45572# a_768_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5538 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5539 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5540 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X5541 a_4883_46098# a_21363_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X5542 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5543 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5544 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5545 DATA[0] a_327_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X5546 VSS a_16751_45260# a_6171_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X5547 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5548 a_16763_47508# a_16588_47582# a_16942_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5549 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5550 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5551 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5552 a_11750_44172# a_10903_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X5553 VDD a_20835_44721# a_20766_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X5554 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5555 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5556 VSS a_15861_45028# a_17668_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X5557 a_7845_44172# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X5558 a_15597_42852# a_15743_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5559 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5560 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5561 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5562 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5563 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5564 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5565 a_n4064_39072# a_n4334_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5566 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5567 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5568 VSS a_9223_42460# a_8953_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X5569 VDD a_11967_42832# a_18083_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5570 a_13487_47204# a_13381_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.16535 ps=1.82 w=0.65 l=0.15
X5571 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5572 C2_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X5573 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5574 a_13297_45572# a_13259_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1034 ps=1 w=0.42 l=0.15
X5575 a_n923_35174# a_n1532_35090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X5576 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5577 VDD a_n3565_38216# a_n3690_38304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X5578 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5579 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5580 C10_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5581 a_6101_43172# a_5891_43370# a_5755_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5582 VSS C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5583 a_11901_46660# a_11735_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5584 a_16979_44734# a_14539_43914# a_17061_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5585 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5586 VSS a_14955_47212# a_10227_46804# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5587 a_18443_44721# a_18248_44752# a_18753_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X5588 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5589 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5590 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5591 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5592 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X5593 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5594 VDD a_18909_45814# a_18799_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X5595 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5596 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5597 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5598 VDAC_N C2_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5599 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5600 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5601 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5602 a_1431_46436# a_1138_42852# a_1337_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X5603 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5604 VDD a_n4064_37984# a_n2216_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X5605 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5606 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5607 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5608 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5609 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5610 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5611 VDD a_22521_40599# a_22469_40625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X5612 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5613 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5614 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5615 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5616 VDD a_768_44030# a_5326_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X5617 a_18443_44721# a_18287_44626# a_18588_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X5618 VSS a_n4209_39304# a_n4251_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X5619 a_n357_42282# a_21356_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X5620 a_491_47026# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X5621 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5622 VSS a_n2288_47178# a_n2312_40392# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5623 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5624 VCM a_1606_42308# C1_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X5625 VDD a_20712_42282# a_10193_42453# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5626 VSS a_3483_46348# a_15301_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X5627 VSS a_13635_43156# a_9290_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X5628 a_n901_46420# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5629 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5630 a_5068_46348# a_5204_45822# a_5210_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5631 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5632 a_14033_45822# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5633 VSS a_6761_42308# a_7227_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5634 VSS a_11599_46634# a_20107_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5635 a_3537_45260# a_7287_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5636 w_1575_34946# EN_VIN_BSTR_P VDD w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X5637 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5638 VDD a_13661_43548# a_15595_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X5639 a_9803_42558# a_n97_42460# a_9885_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5640 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5641 VDD a_10227_46804# a_11136_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X5642 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5643 a_n1177_43370# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5644 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5645 VREF_GND a_n3420_39616# C8_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5646 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5647 VDD a_n2946_39072# a_n3565_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5648 a_601_46902# a_383_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X5649 VDAC_Ni a_3754_38470# a_3726_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X5650 a_5024_45822# a_n443_46116# a_4419_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X5651 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5652 a_17701_42308# a_17531_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5653 VSS a_12861_44030# a_13487_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X5654 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X5655 a_6598_45938# a_6472_45840# a_6194_45824# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X5656 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5657 a_4808_45572# a_1823_45246# a_4419_46090# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X5658 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5659 a_n3607_38304# a_n3674_38216# a_n3690_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X5660 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5661 a_n229_43646# a_n2497_47436# a_n447_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X5662 VSS a_6969_46634# a_6903_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5663 a_18214_42558# a_18184_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X5664 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5665 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5666 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5667 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5668 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5669 VSS a_4883_46098# a_10355_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X5670 VDD a_4646_46812# a_6031_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5671 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5672 a_491_47026# a_n133_46660# a_383_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5673 VDD a_16327_47482# a_18588_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X5674 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5675 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5676 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5677 VSS a_n1613_43370# a_n1655_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5678 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5679 VDAC_Ni VSS a_5088_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X5680 a_6812_45938# a_6598_45938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X5681 a_8147_43396# a_n443_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5682 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5683 a_12427_45724# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.1281 ps=1.03 w=0.42 l=0.15
X5684 C9_N_btm a_17730_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5685 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5686 VDD a_19594_46812# a_19551_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X5687 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5688 a_n4318_37592# a_n1736_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X5689 a_9290_44172# a_13635_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5690 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5691 VSS a_1736_39043# a_1239_39043# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5692 a_1414_42308# a_1067_42314# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X5693 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5694 VSS a_2698_46116# a_2804_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5695 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5696 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5697 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5698 VSS a_5649_42852# a_22223_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5699 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5700 VDD a_13259_45724# a_14797_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X5701 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5702 a_4817_46660# a_4651_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5703 a_n2288_47178# a_n2109_47186# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5704 a_8062_46155# a_8016_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X5705 VDD a_20623_43914# a_20365_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X5706 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5707 a_949_44458# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5708 a_13296_44484# a_12891_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X5709 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5710 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5711 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5712 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5713 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5714 a_11601_46155# a_11309_47204# a_11387_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X5715 a_10210_45822# a_8746_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X5716 a_18287_44626# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5717 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5718 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5719 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5720 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5721 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5722 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5723 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5724 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5725 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X5726 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5727 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5728 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5729 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5730 VSS a_11189_46129# a_11133_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X5731 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5732 a_n3565_38216# a_n2946_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X5733 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5734 a_6109_44484# a_5518_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5735 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5736 a_6431_45366# a_5937_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X5737 a_14021_43940# a_13483_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X5738 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5739 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5740 a_17499_43370# a_17324_43396# a_17678_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5741 a_3495_45348# a_3429_45260# a_3316_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X5742 VDD a_1115_44172# a_n2293_45010# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X5743 VDD a_19787_47423# a_19594_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5744 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5745 a_18707_42852# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X5746 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5747 a_1208_46090# a_n881_46662# a_1431_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X5748 a_n1809_44850# a_n2433_44484# a_n1917_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5749 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5750 a_5431_46482# a_n1151_42308# a_5068_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X5751 a_8667_46634# a_8492_46660# a_8846_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5752 a_19787_47423# START VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5753 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5754 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5755 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5756 a_n2302_39866# a_n2442_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5757 VSS a_n2438_43548# a_2443_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5758 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5759 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5760 a_18797_44260# a_13661_43548# a_18451_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5761 a_19551_46910# a_19692_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5762 VDD a_10341_43396# a_22591_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X5763 a_8697_45822# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X5764 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5765 VDD a_8953_45546# a_8049_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5766 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5767 a_12005_46116# a_2063_45854# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5768 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5769 VSS a_2123_42473# a_1184_42692# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5770 VSS a_12861_44030# a_18911_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.194 pd=1.95 as=0.1092 ps=1.36 w=0.42 l=0.15
X5771 a_1241_43940# a_584_46384# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X5772 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5773 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5774 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5775 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5776 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5777 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5778 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5779 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5780 a_16285_47570# a_16241_47178# a_16119_47582# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X5781 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5782 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5783 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5784 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5785 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5786 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5787 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5788 VSS a_961_42354# a_1067_42314# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5789 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X5790 a_10617_44484# a_10440_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X5791 a_1423_45028# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5792 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5793 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5794 C7_P_btm a_n4064_39072# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X5795 VDD a_4704_46090# a_1823_45246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5796 a_18479_47436# a_20075_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X5797 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5798 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5799 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5800 a_19987_42826# a_10193_42453# a_20573_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X5801 VDD a_9313_45822# a_11459_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X5802 VSS a_n3690_39392# a_n3420_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X5803 a_n1809_44850# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X5804 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5805 VSS a_3785_47178# a_3815_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5806 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5807 a_n3420_39072# a_n3690_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5808 VDD a_5891_43370# a_8375_44464# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5809 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5810 VSS a_9863_46634# a_2063_45854# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X5811 a_7920_46348# a_n1151_42308# a_8062_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5812 a_19721_31679# a_22959_45036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5813 a_19808_44306# a_19778_44110# a_19328_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5814 VDD a_10193_42453# a_11633_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5815 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5816 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5817 VDD a_15559_46634# a_13059_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5818 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5819 VSS a_n2840_43370# a_n4318_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5820 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5821 a_15037_43396# a_14205_43396# a_14955_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X5822 VDD a_11189_46129# a_11601_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X5823 a_5263_45724# a_5257_43370# a_5437_45600# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X5824 a_12495_44260# a_12429_44172# a_10949_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.2275 ps=2 w=0.65 l=0.15
X5825 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5826 a_6452_43396# a_6293_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X5827 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5828 VSS a_4915_47217# a_12891_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5829 a_14084_46812# a_13885_46660# a_14226_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5830 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5831 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5832 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5833 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5834 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5835 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5836 a_19478_44306# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X5837 a_7705_45326# a_7229_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X5838 a_1115_44172# a_1307_43914# a_1241_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X5839 a_8953_45002# CLK VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5840 a_16981_45144# a_16922_45042# a_16886_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X5841 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5842 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5843 a_4223_44672# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5844 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5845 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5846 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5847 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5848 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5849 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5850 a_7174_31319# a_20107_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5851 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5852 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5853 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5854 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5855 VDD a_10227_46804# a_15051_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5856 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5857 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5858 VDD a_n2302_39866# a_n4209_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5859 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5860 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5861 CLK_DATA a_n2833_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5862 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X5863 VSS a_8103_44636# a_7640_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X5864 a_15146_44811# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X5865 a_n4209_39304# a_n2302_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5866 a_n2833_47464# a_n2497_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X5867 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5868 a_2903_45348# a_n971_45724# a_2809_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X5869 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5870 VSS a_3537_45260# a_8103_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5871 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5872 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5873 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5874 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5875 VSS a_21137_46414# a_21071_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5876 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5877 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5878 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5879 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5880 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5881 VSS a_1414_42308# a_2889_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5882 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5883 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5884 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5885 VDD a_1848_45724# a_1799_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X5886 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5887 VSS a_n13_43084# a_n1853_43023# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X5888 a_18479_45785# a_19268_43646# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5889 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5890 VSS a_19279_43940# a_21398_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X5891 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5892 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5893 a_1736_39587# a_1343_38525# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X5894 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5895 VSS a_22485_44484# a_20974_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5896 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5897 VSS a_n3420_37984# a_n2946_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X5898 a_5841_44260# a_5495_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X5899 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5900 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5901 a_5275_47026# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X5902 C5_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X5903 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5904 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5905 a_n2661_45546# a_4093_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5906 VSS a_n2302_38778# a_n4209_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5907 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5908 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5909 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5910 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5911 VSS a_5497_46414# a_5431_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5912 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5913 VDD a_19339_43156# a_19326_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5914 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5915 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5916 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5917 VDD a_6123_31319# a_7963_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5918 a_8137_45348# a_8049_45260# a_n2293_42834# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5919 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5920 VDD a_17499_43370# a_n1059_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X5921 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5922 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5923 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5924 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5925 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5926 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5927 VDD a_12861_44030# a_17339_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5928 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5929 a_10849_43646# a_10807_43548# a_10765_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5930 VSS a_13507_46334# a_18997_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X5931 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5932 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5933 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5934 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5935 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5936 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5937 a_8560_45348# a_3483_46348# a_8488_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X5938 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5939 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5940 VDD a_n3690_38304# a_n3420_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5941 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5942 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5943 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5944 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5945 a_13249_42308# a_13070_42354# a_13333_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X5946 a_6969_46634# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X5947 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5948 a_n2216_37984# a_n2810_45572# a_n2302_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X5949 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5950 VSS a_22223_46124# a_20205_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5951 VSS a_n1613_43370# a_n1379_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5952 a_6194_45824# a_6511_45714# a_6469_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X5953 a_n229_43646# a_n97_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5954 a_17613_45144# a_8696_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5955 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5956 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5957 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5958 VSS a_13747_46662# a_19862_44208# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5959 a_22821_38993# a_22400_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5960 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5961 a_17303_42282# a_n913_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5962 a_8649_43218# a_8605_42826# a_8483_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X5963 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5964 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5965 VSS a_n901_46420# a_n967_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X5966 a_15004_44636# a_13556_45296# a_15146_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5967 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5968 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5969 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5970 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5971 a_11186_47026# a_10467_46802# a_10623_46897# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X5972 a_n1076_46494# a_n2157_46122# a_n1423_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X5973 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5974 VSS a_526_44458# a_4169_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X5975 a_3353_43940# a_2998_44172# a_2675_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5976 a_n23_45546# a_n356_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X5977 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5978 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5979 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5980 a_18326_43940# a_18079_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X5981 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5982 a_18194_35068# a_n1630_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5983 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5984 a_20922_43172# a_19862_44208# a_20753_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X5985 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5986 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5987 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5988 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5989 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5990 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5991 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5992 C5_P_btm a_5934_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X5993 a_10334_44484# a_10157_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X5994 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5995 a_n2017_45002# a_19987_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.208 ps=1.94 w=0.65 l=0.15
X5996 VSS a_742_44458# a_1756_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5997 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5998 a_n2956_38216# a_n2472_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5999 VDD a_10193_42453# a_13657_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6000 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6001 VDD a_8191_45002# a_n2293_42834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6002 a_13885_46660# a_13607_46688# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X6003 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6004 VSS RST_Z a_7754_39964# VSS sky130_fd_pr__nfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.15
X6005 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6006 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6007 VSS a_4223_44672# a_n2497_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6008 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6009 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6010 a_4699_43561# a_3080_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6011 a_19511_42282# a_18597_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6012 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6013 a_n3420_37984# a_n3690_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X6014 VSS a_19692_46634# a_743_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6015 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6016 VDD a_22591_43396# a_14209_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6017 a_n1991_46122# a_n2157_46122# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6018 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6019 VDD a_n4334_39392# a_n4064_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X6020 VDD a_7499_43078# a_8746_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6021 a_n971_45724# a_104_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X6022 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6023 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6024 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6025 a_20447_31679# a_22959_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6026 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6027 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6028 VDD a_15493_43940# a_22959_43948# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6029 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6030 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6031 VSS a_n2302_37690# a_n4209_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6032 a_n4334_39616# a_n4318_39768# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6033 VDD a_13527_45546# a_13163_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X6034 a_18147_46436# a_17339_46660# a_17957_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X6035 a_8336_45822# a_8270_45546# a_n1925_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X6036 a_n2956_39304# a_n2840_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X6037 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6038 VDD a_584_46384# a_766_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X6039 a_11361_45348# a_10907_45822# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6040 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6041 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6042 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6043 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6044 VDD a_11599_46634# a_11735_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6045 a_19431_45546# a_19256_45572# a_19610_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X6046 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6047 VSS a_9290_44172# a_12710_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.118125 pd=1.04 as=0.08775 ps=0.92 w=0.65 l=0.15
X6048 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6049 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6050 VDD a_11323_42473# a_10807_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6051 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6052 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6053 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6054 a_2266_47243# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X6055 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6056 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6057 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6058 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6059 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6060 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6061 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6062 a_2982_43646# a_2479_44172# a_2896_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6063 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6064 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6065 a_18280_46660# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6066 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6067 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6068 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6069 C1_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X6070 VDD a_8492_46660# a_8667_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6071 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6072 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X6073 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6074 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6075 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6076 VDD a_11967_42832# a_12379_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6077 VDD a_n1076_46494# a_n901_46420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6078 a_n4251_38528# a_n4318_38680# a_n4334_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X6079 a_4361_42308# a_3823_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6080 VDD a_n971_45724# a_3775_45552# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6081 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6082 VDD a_11599_46634# a_13759_46122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6083 VDAC_P C2_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6084 VDD a_21811_47423# a_20916_46384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6085 a_18985_46122# a_18819_46122# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6086 VDD a_5649_42852# a_22223_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6087 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6088 VSS a_5343_44458# a_8333_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6089 VDD a_7287_43370# a_3537_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6090 VSS a_3090_45724# a_10555_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X6091 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6092 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6093 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6094 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6095 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6096 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6097 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6098 a_20528_45572# a_19466_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X6099 a_13487_47204# a_13717_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6100 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6101 VREF_GND a_13678_32519# C2_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X6102 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6103 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6104 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6105 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6106 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6107 VDD a_20269_44172# a_19319_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X6108 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6109 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6110 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6111 a_5807_45002# a_16763_47508# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X6112 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6113 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6114 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6115 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6116 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6117 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6118 VSS a_16327_47482# a_16285_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6119 a_n23_44458# a_n356_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6120 VDD a_n1059_45260# a_8791_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X6121 a_1847_42826# a_2351_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6122 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X6123 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6124 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6125 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6126 VSS a_3503_45724# a_3218_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X6127 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6128 a_19553_46090# a_19335_46494# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X6129 VDD a_n2840_45546# a_n2810_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X6130 a_15037_45618# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6131 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6132 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6133 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6134 a_14537_43646# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X6135 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6136 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6137 VDD a_1307_43914# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6138 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6139 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6140 a_n1699_43638# a_n1917_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X6141 VDD a_9313_44734# a_22959_42860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6142 C6_P_btm a_n3420_39072# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X6143 VDD a_n2946_38778# a_n3565_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6144 a_6671_43940# a_5205_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6145 VSS a_5111_44636# a_4905_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X6146 a_2124_47436# a_2063_45854# a_2266_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X6147 a_n4064_37984# a_n4334_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6148 VSS a_9625_46129# a_9569_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X6149 VDD a_3483_46348# a_13565_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X6150 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6151 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6152 VDD a_19279_43940# a_21398_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X6153 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6154 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6155 a_6171_42473# a_5932_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6156 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6157 a_17568_45572# a_8696_44636# a_17478_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X6158 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6159 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6160 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6161 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6162 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6163 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6164 a_18588_44850# a_18374_44850# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X6165 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6166 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6167 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6168 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6169 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6170 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6171 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6172 a_22465_38105# a_22775_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X6173 a_18451_43940# a_18579_44172# a_18533_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6174 VSS a_5755_42308# a_5932_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X6175 a_2959_46660# a_2609_46660# a_2864_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6176 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6177 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6178 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6179 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6180 a_21359_45002# a_21513_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6181 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6182 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6183 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6184 a_7_47243# a_n746_45260# a_n452_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X6185 a_14493_46090# a_14275_46494# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X6186 a_19478_44306# a_15493_43396# a_19478_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X6187 a_7287_43370# a_7112_43396# a_7466_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X6188 a_15227_46910# a_3090_45724# a_15009_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X6189 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6190 VSS a_n1630_35242# a_n1532_35090# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6191 a_12251_46660# a_11901_46660# a_12156_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6192 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6193 a_8495_42852# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X6194 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6195 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6196 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6197 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6198 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6199 a_11633_42558# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X6200 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6201 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6202 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6203 a_n4251_37440# a_n4318_37592# a_n4334_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X6204 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6205 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6206 a_15279_43071# a_5342_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6207 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6208 VDD a_7276_45260# a_7227_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X6209 VSS a_2479_44172# a_2813_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X6210 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6211 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6212 VREF_GND a_14401_32519# C6_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X6213 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6214 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6215 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6216 VDD a_n815_47178# a_n785_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6217 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6218 VDD a_3877_44458# a_3699_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X6219 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6220 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6221 a_9313_45822# a_5937_45572# a_9241_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X6222 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6223 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6224 a_1239_47204# a_1209_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6225 a_20841_45814# a_20623_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X6226 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6227 VDD a_805_46414# a_835_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6228 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6229 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6230 a_6298_44484# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6231 a_961_42354# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6232 a_12379_46436# a_12005_46116# a_n1741_47186# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6233 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6234 a_4338_37500# a_3754_38470# VDAC_Pi VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X6235 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6236 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6237 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6238 VDD a_5257_43370# a_3905_42865# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6239 VSS C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6240 a_n1741_47186# a_12594_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6241 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6242 a_n2956_39768# a_n2840_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X6243 VSS a_n473_42460# a_n1761_44111# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X6244 a_13163_45724# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.1281 ps=1.03 w=0.42 l=0.15
X6245 a_10210_45822# a_10586_45546# a_10053_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6246 VDD a_10227_46804# a_9863_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6247 a_22465_38105# a_22775_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X6248 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6249 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6250 VSS a_4185_45028# a_22959_45036# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6251 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6252 VDD a_n2438_43548# a_n2065_43946# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6253 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6254 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6255 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6256 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6257 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6258 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6259 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X6260 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6261 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6262 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6263 a_5457_43172# a_5111_44636# a_5111_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X6264 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6265 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6266 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6267 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6268 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6269 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6270 a_10695_43548# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X6271 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6272 VDD a_11787_45002# a_11652_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X6273 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6274 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6275 VDD a_n2946_37690# a_n3565_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6276 a_13059_46348# a_15559_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6277 VDD a_n23_44458# a_7_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6278 a_12891_46348# a_4915_47217# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6279 a_8023_46660# a_7577_46660# a_7927_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6280 VSS a_10057_43914# a_9672_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6281 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6282 a_20637_44484# a_20159_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X6283 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6284 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6285 a_n237_47217# a_8667_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X6286 a_n143_45144# a_n755_45592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6287 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6288 a_4520_42826# a_4905_42826# a_4649_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X6289 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6290 VSS RST_Z a_8530_39574# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6291 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6292 VSS a_n971_45724# a_8423_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X6293 a_n1379_43218# a_n1423_42826# a_n1545_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X6294 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6295 VSS a_n2946_37984# a_n3565_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6296 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X6297 VSS a_3626_43646# a_19647_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6298 a_8697_45822# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X6299 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6300 VDD a_n4334_39616# a_n4064_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6301 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6302 a_n443_42852# a_n901_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6303 a_3094_47243# a_2905_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X6304 a_15051_42282# a_15486_42560# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X6305 VDD a_1209_47178# a_1239_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6306 a_11823_42460# a_15051_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6307 a_n1641_46494# a_n2157_46122# a_n1736_46482# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6308 VDD a_13661_43548# a_16241_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X6309 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6310 a_5167_46660# a_4817_46660# a_5072_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6311 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6312 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6313 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6314 VSS a_10835_43094# a_10796_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6315 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6316 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6317 VDD a_20708_46348# a_20411_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X6318 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6319 VSS a_16327_47482# a_18005_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X6320 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6321 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6322 VSS a_16292_46812# a_15811_47375# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X6323 a_9482_43914# a_9838_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6324 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6325 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X6326 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6327 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6328 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6329 a_20623_46660# a_20273_46660# a_20528_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6330 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6331 VDD a_12594_46348# a_n1741_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6332 a_18374_44850# a_18287_44626# a_17970_44736# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X6333 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6334 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6335 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6336 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6337 a_16750_47204# a_15673_47210# a_16588_47582# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6338 a_6545_47178# a_6419_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X6339 VDD a_22223_43396# a_13887_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6340 a_8783_44734# a_8696_44636# a_8701_44490# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6341 a_175_44278# a_n863_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X6342 VSS C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6343 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6344 VSS a_7754_38470# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X6345 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X6346 VSS a_n901_46420# a_n443_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X6347 VDD a_18479_47436# a_20935_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6348 a_3754_38470# a_7754_38470# VSS sky130_fd_pr__res_high_po_0p35 l=18
X6349 VSS a_5907_46634# a_5841_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X6350 a_5745_43940# a_5883_43914# a_5829_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6351 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6352 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6353 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6354 a_1110_47026# a_33_46660# a_948_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6355 a_16434_46987# a_16388_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X6356 VSS a_2324_44458# a_15682_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6357 VDD a_n2302_39866# a_n4209_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6358 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6359 a_20974_43370# a_22485_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6360 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6361 a_2998_44172# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6362 a_13381_47204# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6363 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6364 VDD a_4921_42308# a_5755_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6365 a_10991_42826# a_10835_43094# a_11136_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X6366 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6367 VSS a_n4334_38528# a_n4064_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6368 VDD a_6851_47204# a_7227_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X6369 a_3052_44056# a_2998_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X6370 a_n1699_43638# a_n1917_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X6371 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6372 CAL_N a_22465_38105# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X6373 a_3177_46902# a_2959_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X6374 a_9241_44734# a_5937_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6375 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6376 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6377 VSS a_1208_46090# a_472_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X6378 a_22365_46825# EN_OFFSET_CAL VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6379 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6380 VSS a_13163_45724# a_11962_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X6381 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6382 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6383 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6384 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6385 a_3055_46660# a_2609_46660# a_2959_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6386 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6387 a_19326_42852# a_18249_42858# a_19164_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6388 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6389 a_9885_43646# a_8270_45546# a_9803_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6390 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6391 a_n443_46116# a_n901_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6392 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6393 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6394 VDD a_18597_46090# a_16375_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6395 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6396 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6397 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6398 VSS a_22959_43396# a_17364_32525# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X6399 a_19431_45546# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6400 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6401 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6402 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6403 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6404 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6405 VDD a_n3690_38304# a_n3420_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X6406 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6407 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6408 a_n4064_39616# a_n4334_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X6409 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6410 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6411 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6412 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6413 VSS a_n1177_44458# a_n1243_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X6414 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6415 VSS a_n23_45546# a_n89_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X6416 VDD a_12816_46660# a_12991_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6417 a_7499_43940# a_7640_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6418 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6419 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X6420 a_2952_47436# a_n1151_42308# a_3094_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X6421 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6422 VSS a_n2302_38778# a_n4209_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6423 a_n452_47436# a_n746_45260# a_n310_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X6424 a_4235_43370# a_3935_42891# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X6425 a_5105_45348# a_4558_45348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6426 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6427 VSS a_n1838_35608# SMPL_ON_P VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6428 a_18051_46116# a_765_45546# a_17957_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X6429 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6430 a_n1441_43940# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X6431 a_15301_44260# a_15227_44166# a_14955_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X6432 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6433 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6434 VSS a_n3565_38502# a_n3607_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X6435 a_n746_45260# a_n1177_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X6436 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6437 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6438 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6439 a_n2840_43914# a_n2661_43922# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X6440 a_6809_43396# a_6765_43638# a_6643_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X6441 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6442 VSS a_376_46348# a_171_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X6443 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6444 VSS a_8199_44636# a_8701_44490# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6445 a_7499_43940# a_3090_45724# a_7281_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X6446 a_9165_43940# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6447 a_19443_46116# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X6448 VSS a_13059_46348# a_15143_45578# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X6449 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6450 a_453_43940# a_175_44278# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X6451 a_9885_42308# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6452 a_n3674_39304# a_n2840_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X6453 a_2959_46660# a_2443_46660# a_2864_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6454 a_14543_46987# a_13885_46660# a_14084_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X6455 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6456 VDD a_413_45260# a_22959_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6457 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6458 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6459 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6460 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6461 a_17969_45144# a_16375_45002# a_17896_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X6462 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6463 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6464 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6465 a_n4064_38528# a_n4334_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X6466 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6467 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6468 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6469 a_16292_46812# a_n743_46660# a_16434_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X6470 a_21188_46660# a_20107_46660# a_20841_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X6471 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6472 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6473 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6474 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6475 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6476 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6477 a_4365_46436# a_4185_45028# a_n1925_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6478 a_12251_46660# a_11735_46660# a_12156_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6479 a_n998_44484# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X6480 VDD a_n2472_45546# a_n2956_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X6481 a_7577_46660# a_7411_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6482 a_10835_43094# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6483 VDD a_3177_46902# a_3067_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X6484 a_14976_45028# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X6485 a_n3420_37984# a_n3690_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6486 VSS a_13661_43548# a_743_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6487 a_12638_46436# a_12891_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X6488 a_n1352_44484# a_n2433_44484# a_n1699_44726# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X6489 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6490 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6491 a_12839_46116# a_12891_46348# a_n1741_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6492 VSS a_3090_45724# a_4927_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6493 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6494 VSS a_22000_46634# a_15227_44166# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X6495 VSS a_n863_45724# a_791_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X6496 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6497 a_14209_32519# a_22591_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X6498 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6499 VSS a_n4334_37440# a_n4064_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6500 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6501 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6502 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6503 a_n2012_43396# a_n2129_43609# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X6504 VSS a_11823_42460# a_14635_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6505 a_n1613_43370# a_5815_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6506 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6507 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6508 a_n2661_43922# a_12465_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6509 C8_P_btm a_n3565_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6510 VSS a_4520_42826# a_4093_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X6511 a_19692_46634# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6512 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6513 a_5013_44260# a_3905_42865# a_5025_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6514 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6515 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6516 VSS C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6517 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6518 a_8018_44260# a_7499_43078# a_7911_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X6519 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6520 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6521 VDD a_11823_42460# a_14358_43442# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X6522 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6523 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6524 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6525 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6526 a_742_44458# a_n443_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6527 VDD a_10405_44172# a_8016_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X6528 a_20254_46482# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X6529 VIN_N EN_VIN_BSTR_N C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X6530 a_167_45260# a_2202_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X6531 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6532 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6533 VSS a_19332_42282# a_4190_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X6534 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6535 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6536 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6537 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6538 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6539 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6540 a_20356_42852# a_18184_42460# a_20256_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.175 ps=1.35 w=1 l=0.15
X6541 a_14840_46494# a_13925_46122# a_14493_46090# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6542 VSS a_1414_42308# a_3457_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X6543 a_19006_44850# a_18287_44626# a_18443_44721# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X6544 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6545 a_9420_43940# a_768_44030# a_9165_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X6546 VDD a_10903_43370# a_12005_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6547 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6548 a_n4209_38216# a_n2302_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6549 VSS a_13661_43548# a_15685_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X6550 VSS a_12861_44030# a_18280_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6551 C4_P_btm a_6123_31319# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X6552 a_13575_42558# a_n97_42460# a_13657_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X6553 VSS a_n2302_37690# a_n4209_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6554 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6555 VDAC_P C2_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6556 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6557 a_8667_46634# a_6151_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6558 a_n1533_42852# a_n2157_42858# a_n1641_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X6559 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6560 VDD a_n971_45724# a_n229_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X6561 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6562 a_n1613_43370# a_5815_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6563 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6564 a_21335_42336# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X6565 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6566 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6567 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6568 VSS a_n3565_37414# a_n3607_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X6569 a_n2946_38778# a_n2956_38680# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6570 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6571 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6572 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6573 VSS a_9127_43156# a_5891_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X6574 VSS a_13351_46090# a_10903_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X6575 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6576 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6577 a_743_42282# a_12549_44172# a_20749_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X6578 a_14309_45028# a_2711_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X6579 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6580 VSS a_413_45260# a_22959_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6581 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6582 VDD a_3877_44458# a_4185_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6583 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6584 a_13105_45348# a_13017_45260# a_n2661_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6585 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6586 a_8229_43396# a_7499_43078# a_8147_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X6587 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6588 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6589 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6590 VSS a_6545_47178# a_6575_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6591 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6592 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6593 a_19551_46910# a_19466_46812# a_19333_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X6594 a_6945_45028# a_5205_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6595 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6596 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6597 a_18280_46660# a_12549_44172# a_17609_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X6598 VSS a_18285_46348# a_18243_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X6599 a_3726_37500# a_3754_38470# VDAC_Ni VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X6600 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6601 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6602 a_n4064_37440# a_n4334_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X6603 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6604 a_20708_46348# a_20916_46384# a_20850_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X6605 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6606 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6607 a_5167_46660# a_4651_46660# a_5072_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6608 VDD a_n1352_44484# a_n1177_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6609 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6610 a_15685_45394# a_15415_45028# a_15595_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X6611 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6612 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6613 VDD a_10193_42453# a_18214_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X6614 a_21350_45938# a_20273_45572# a_21188_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6615 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6616 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6617 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6618 comp_n a_1239_39043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6619 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6620 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6621 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6622 a_7765_42852# a_7227_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X6623 VSS a_526_44458# a_10149_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X6624 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6625 a_7639_45394# a_n1151_42308# a_7276_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X6626 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6627 a_501_45348# a_413_45260# a_375_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6628 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6629 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6630 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6631 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6632 a_16547_43609# a_16414_43172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X6633 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6634 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6635 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6636 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6637 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X6638 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6639 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6640 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6641 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6642 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6643 a_5891_43370# a_9127_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6644 a_n3565_38502# a_n2946_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6645 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6646 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6647 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6648 a_13857_44734# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6649 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6650 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6651 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6652 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6653 a_n2661_46098# a_2107_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X6654 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6655 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6656 VSS a_16327_47482# a_18953_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6657 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6658 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6659 VSS a_742_44458# a_1568_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6660 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6661 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6662 a_19273_43230# a_18083_42858# a_19164_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6663 a_6123_31319# a_7227_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X6664 a_768_44030# a_13487_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X6665 a_12293_43646# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X6666 a_584_46384# a_1123_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6667 VDD a_2711_45572# a_4099_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6668 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6669 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6670 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6671 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6672 C8_N_btm a_5342_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X6673 a_10306_45572# a_10193_42453# a_10216_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X6674 a_n1917_44484# a_n2433_44484# a_n2012_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6675 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6676 a_8035_47026# a_6151_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X6677 a_18545_45144# a_13259_45724# a_18450_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X6678 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6679 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6680 VDD a_21855_43396# a_13678_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6681 a_16977_43638# a_16759_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X6682 a_n1423_46090# a_n1641_46494# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X6683 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6684 VDD a_22223_43948# a_14401_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6685 VDD a_6540_46812# a_6491_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X6686 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6687 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6688 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6689 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6690 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6691 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6692 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6693 VDD a_n863_45724# a_n1099_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X6694 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6695 a_n2946_37690# a_n2956_37592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6696 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6697 C10_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X6698 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6699 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6700 a_5111_42852# a_4905_42826# a_5193_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6701 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6702 VDD a_5263_45724# a_5204_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X6703 a_n467_45028# a_n745_45366# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X6704 VDD a_15095_43370# a_14955_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X6705 VSS a_n4334_38304# a_n4064_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X6706 VSS a_765_45546# a_1208_46090# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6707 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6708 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X6709 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6710 VDD a_2957_45546# a_2905_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6711 a_8855_44734# a_4791_45118# a_8783_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6712 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6713 a_11963_45334# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X6714 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6715 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6716 a_n2661_44458# a_11453_44696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.182 ps=1.92 w=0.7 l=0.15
X6717 VDD a_4915_47217# a_11415_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6718 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6719 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6720 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6721 a_3600_43914# a_3537_45260# a_3820_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6722 a_n1741_47186# a_12005_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6723 a_1848_45724# a_2063_45854# a_1990_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X6724 a_21588_30879# a_22223_47212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6725 a_14537_46482# a_14493_46090# a_14371_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X6726 a_16241_44734# a_2711_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X6727 a_3905_42865# a_5257_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6728 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6729 a_10425_46660# a_9863_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X6730 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6731 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6732 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6733 a_19365_45572# a_18175_45572# a_19256_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6734 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6735 a_21811_47423# SINGLE_ENDED VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6736 VDD a_22959_45572# a_20447_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6737 a_3090_45724# a_18911_45144# a_19113_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6738 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6739 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6740 a_13777_45326# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6741 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6742 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6743 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6744 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6745 VCM a_5934_30871# C5_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X6746 a_n3690_39616# a_n3674_39768# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6747 a_17333_42852# a_16795_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6748 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X6749 DATA[2] a_4007_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6750 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6751 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6752 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6753 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6754 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6755 a_11525_45546# a_11962_45724# a_11682_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X6756 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6757 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6758 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6759 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6760 a_17595_43084# a_13259_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X6761 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6762 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6763 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6764 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6765 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6766 a_n13_43084# a_n755_45592# a_133_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X6767 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6768 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6769 a_n1838_35608# a_n1386_35608# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6770 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6771 a_n3565_37414# a_n2946_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6772 a_n2840_42282# a_n2661_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X6773 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6774 a_20193_45348# a_18184_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6775 a_1756_43548# a_768_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6776 a_20719_46660# a_20273_46660# a_20623_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6777 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6778 a_n2302_39072# a_n2312_39304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6779 VSS a_n1613_43370# a_n1379_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6780 a_n2472_43914# a_n2293_43922# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X6781 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6782 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6783 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6784 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6785 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6786 a_14456_42282# a_14635_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X6787 VSS a_2711_45572# a_4099_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6788 VDD a_20075_46420# a_20062_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6789 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6790 a_4927_45028# a_5147_45002# a_5105_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X6791 a_21381_43940# a_21115_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X6792 VSS C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6793 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6794 VSS a_10227_46804# a_10185_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X6795 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6796 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6797 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6798 a_4169_42308# a_1823_45246# a_3823_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X6799 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6800 a_n3607_38528# a_n3674_38680# a_n3690_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X6801 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6802 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6803 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6804 a_4704_46090# a_4883_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X6805 VDD a_20894_47436# a_20843_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X6806 CLK_DATA a_n2833_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X6807 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6808 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6809 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6810 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6811 VSS a_n913_45002# a_6761_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6812 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6813 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6814 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6815 VDD a_15051_42282# a_11823_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6816 VDD a_12465_44636# a_22223_47212# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6817 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6818 VDD a_20193_45348# a_20753_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6819 VSS C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6820 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6821 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6822 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6823 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6824 VDD a_5257_43370# a_3357_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6825 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6826 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X6827 VSS a_14113_42308# a_16522_42674# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X6828 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6829 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6830 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6831 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6832 a_13460_43230# a_12379_42858# a_13113_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X6833 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6834 a_19240_46482# a_19123_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X6835 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6836 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6837 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6838 a_22609_37990# a_22521_39511# CAL_P VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X6839 a_5829_43940# a_5495_43940# a_5745_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6840 VSS C1_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6841 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6842 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6843 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6844 VSS a_21487_43396# a_13467_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X6845 a_10227_46804# a_14955_47212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6846 VDD a_7287_43370# a_7274_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6847 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6848 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6849 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6850 a_14955_43940# a_14537_43396# a_15037_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6851 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6852 VDD a_12861_44030# a_18911_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1468 pd=1.34 as=0.1092 ps=1.36 w=0.42 l=0.15
X6853 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6854 a_15953_42852# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6855 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6856 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6857 a_9114_42852# a_8037_42858# a_8952_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6858 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6859 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6860 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6861 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6862 a_n4315_30879# a_n2302_40160# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X6863 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6864 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6865 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6866 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6867 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6868 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6869 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X6870 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6871 VSS a_8199_44636# a_8953_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X6872 VSS a_n901_46420# a_n443_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6873 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6874 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6875 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6876 VDD a_15227_44166# a_18285_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X6877 a_16375_45002# a_18597_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6878 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6879 a_15279_43071# a_5342_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6880 a_18780_47178# a_18597_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X6881 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6882 VDD a_2324_44458# a_6298_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6883 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6884 a_10193_42453# a_20712_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X6885 a_5205_44484# a_5111_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6886 a_19335_46494# a_18985_46122# a_19240_46482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6887 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6888 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6889 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6890 VSS a_685_42968# a_791_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6891 a_4842_47243# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X6892 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6893 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6894 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6895 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6896 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6897 C8_N_btm a_21076_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6898 VSS a_22591_45572# a_19963_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X6899 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6900 VSS a_11322_45546# a_12016_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X6901 a_20753_42852# a_10193_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X6902 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6903 a_n1059_45260# a_17499_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6904 a_509_45572# a_n1099_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X6905 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6906 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6907 SMPL_ON_P a_n1838_35608# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6908 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6909 DATA[5] a_11459_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6910 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6911 a_n1532_35090# a_n1630_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6912 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6913 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6914 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6915 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6916 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6917 a_n1991_42858# a_n2157_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6918 a_16789_45572# a_15599_45572# a_16680_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6919 a_20362_44736# a_20640_44752# a_20596_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X6920 a_13622_42852# a_12545_42858# a_13460_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6921 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6922 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6923 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6924 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6925 a_8701_44490# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6926 a_n3607_37440# a_n3674_37592# a_n3690_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X6927 VSS a_n746_45260# a_556_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X6928 a_15143_45578# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6929 a_10775_45002# a_10951_45334# a_10903_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X6930 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6931 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6932 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6933 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6934 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6935 VSS a_7227_47204# DATA[3] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X6936 VDD a_6151_47436# a_14955_47212# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6937 a_15673_47210# a_15507_47210# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6938 a_19120_35138# VDD EN_VIN_BSTR_N VSS sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.9
X6939 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6940 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6941 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6942 a_20679_44626# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6943 VDD a_n2946_39072# a_n3565_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6944 VDD a_10991_42826# a_10922_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X6945 a_5815_47464# a_6151_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X6946 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X6947 a_n2956_37592# a_n2472_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X6948 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6949 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6950 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6951 a_13667_43396# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X6952 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6953 VSS a_n1920_47178# a_n2312_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X6954 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6955 VDD a_n4064_40160# a_n2216_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X6956 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6957 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6958 a_5164_46348# a_4927_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X6959 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6960 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6961 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6962 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6963 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6964 a_949_44458# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6965 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6966 a_15940_43402# a_12549_44172# a_15868_43402# VSS sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6967 VDD a_4646_46812# a_4651_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6968 a_1427_43646# a_1049_43396# a_1209_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X6969 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6970 a_19164_43230# a_18249_42858# a_18817_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6971 a_2982_43646# a_3232_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X6972 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6973 VDD a_12861_44030# a_21845_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6974 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6975 a_648_43396# a_526_44458# a_548_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X6976 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6977 VDD a_3600_43914# a_3499_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X6978 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6979 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6980 a_16409_43396# a_16243_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6981 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6982 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6983 VSS a_2063_45854# a_11136_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X6984 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6985 VSS a_21589_35634# SMPL_ON_N VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6986 VSS a_1823_45246# a_2202_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6987 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6988 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6989 VDD a_n3420_39616# a_n2860_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X6990 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6991 a_10903_45394# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X6992 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6993 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6994 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6995 a_9290_44172# a_13635_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6996 VSS a_n971_45724# a_3775_45552# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6997 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6998 a_18243_46436# a_18189_46348# a_18147_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
X6999 a_4700_47436# a_4915_47217# a_4842_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X7000 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7001 VDD a_6453_43914# a_n2661_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7002 VSS a_n2438_43548# a_n2433_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7003 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7004 VDD a_10053_45546# a_9625_46129# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X7005 VDD a_12861_44030# a_19615_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X7006 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7007 VDD a_13113_42826# a_13003_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X7008 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7009 VDD a_380_45546# a_n356_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X7010 a_11813_46116# a_11387_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X7011 a_2253_43940# a_n443_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X7012 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7013 a_765_45546# a_17609_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7014 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7015 a_3503_45724# a_1823_45246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X7016 VDD a_9625_46129# a_10037_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X7017 VDD a_3699_46348# a_3160_47472# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X7018 a_18997_42308# a_18727_42674# a_18907_42674# VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X7019 a_5755_42852# a_n97_42460# a_5837_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7020 VDD a_22223_45036# a_18114_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7021 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7022 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7023 EN_VIN_BSTR_P a_n1532_35090# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X7024 VDAC_Pi VSS a_5700_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X7025 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7026 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7027 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7028 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7029 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7030 a_12281_43396# a_n913_45002# a_12293_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7031 VDD a_10533_42308# a_10723_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7032 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7033 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7034 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7035 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7036 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7037 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7038 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7039 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7040 VSS a_9863_47436# a_9804_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X7041 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7042 VDD a_8791_42308# a_5934_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7043 a_11387_46482# a_11133_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X7044 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7045 VDD a_21005_45260# a_19778_44110# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X7046 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7047 a_8049_45260# a_n237_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7048 VDD a_13487_47204# a_768_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7049 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7050 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7051 VSS a_n3420_38528# a_n2946_38778# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X7052 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7053 VDD a_4646_46812# a_7871_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7054 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X7055 a_895_43940# a_644_44056# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X7056 C3_P_btm a_n4064_37984# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X7057 a_19256_45572# a_18341_45572# a_18909_45814# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7058 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7059 VSS a_2713_42308# a_2903_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7060 a_3067_47026# a_2443_46660# a_2959_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X7061 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7062 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7063 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7064 a_9863_47436# a_2063_45854# a_10037_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X7065 a_15037_45618# a_13259_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7066 a_10991_42826# a_10796_42968# a_11301_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X7067 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7068 a_3726_37500# CAL_P a_11206_38545# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X7069 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7070 a_2127_44172# a_1307_43914# a_2253_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X7071 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7072 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7073 a_1823_45246# a_4704_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7074 VDD a_n2438_43548# a_n2433_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7075 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7076 a_17678_43396# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X7077 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7078 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7079 a_3080_42308# a_2903_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7080 VDD a_10903_43370# a_12427_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.06615 ps=0.735 w=0.42 l=0.15
X7081 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7082 a_n452_47436# a_n237_47217# a_n310_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X7083 a_18057_42282# a_n1059_45260# a_18310_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X7084 VSS a_n452_45724# a_n1853_46287# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X7085 a_n3674_39768# a_n2472_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7086 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7087 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7088 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7089 a_8846_46660# a_6151_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X7090 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7091 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7092 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7093 a_1307_43914# a_2779_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7094 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7095 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7096 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=10
X7097 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7098 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7099 a_22365_46825# EN_OFFSET_CAL VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7100 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7101 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7102 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7103 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7104 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7105 a_n2472_42282# a_n2293_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X7106 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7107 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7108 a_n89_45572# a_n743_46660# a_n452_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7109 VSS a_n2840_45002# a_n2810_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7110 a_15928_47570# a_15811_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X7111 a_518_46482# a_472_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X7112 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7113 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7114 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7115 a_n3420_39616# a_n3690_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X7116 a_15463_44811# a_11691_44458# a_15004_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X7117 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7118 a_20556_43646# a_19692_46634# a_20301_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7119 VSS a_17767_44458# a_17715_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X7120 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7121 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7122 a_9061_43230# a_7871_42858# a_8952_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X7123 a_14309_45028# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X7124 a_16237_45028# a_16375_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7125 a_8791_43396# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X7126 VDD a_n4209_38216# a_n4334_38304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X7127 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7128 VDD a_n1423_42826# a_n1533_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X7129 a_1568_43370# a_n863_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7130 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7131 a_22780_39857# a_22465_38105# a_22521_39511# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X7132 a_n1379_46482# a_n1423_46090# a_n1545_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X7133 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7134 a_13575_42558# a_n97_42460# a_13657_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7135 a_6667_45809# a_6511_45714# a_6812_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X7136 a_3754_39964# a_7754_39964# VSS sky130_fd_pr__res_high_po_0p35 l=18
X7137 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7138 a_16115_45572# a_15765_45572# a_16020_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7139 VDD a_18911_45144# a_3090_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.165 ps=1.33 w=1 l=0.15
X7140 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7141 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7142 VSS a_9290_44172# a_10586_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7143 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7144 VDD a_3499_42826# a_n2293_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7145 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7146 a_2725_42558# a_n755_45592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7147 a_18504_43218# a_17333_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X7148 a_2253_43940# a_2479_44172# a_2455_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7149 a_16979_44734# a_14539_43914# a_17061_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X7150 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7151 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7152 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7153 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7154 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7155 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7156 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7157 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7158 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7159 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7160 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7161 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7162 VSS a_1307_43914# a_3681_42891# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X7163 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7164 VSS a_626_44172# a_648_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X7165 VSS a_n3420_37440# a_n2946_37690# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X7166 a_n3420_38528# a_n3690_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X7167 a_21356_42826# a_21381_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7168 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7169 a_1343_38525# a_1177_38525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7170 a_n310_47243# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X7171 a_5025_43940# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7172 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7173 a_16877_43172# a_16823_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7174 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X7175 a_20841_46902# a_20623_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X7176 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7177 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7178 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7179 VSS a_6171_45002# a_6125_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X7180 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7181 VSS a_17595_43084# a_14539_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X7182 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7183 a_5883_43914# a_8333_44056# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X7184 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7185 a_21137_46414# a_19692_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X7186 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7187 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7188 a_20766_44850# a_20640_44752# a_20362_44736# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X7189 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7190 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7191 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7192 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7193 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7194 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7195 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7196 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7197 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7198 a_805_46414# a_472_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X7199 a_1176_45822# a_997_45618# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X7200 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7201 VDAC_N C1_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7202 a_21887_42336# a_20202_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7203 VSS a_11967_42832# a_18083_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7204 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X7205 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7206 DATA[2] a_4007_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X7207 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7208 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7209 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7210 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7211 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7212 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7213 VDD a_1823_45246# a_3316_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X7214 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7215 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7216 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7217 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7218 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7219 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7220 a_21513_45002# a_21363_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X7221 a_8704_45028# a_5937_45572# a_8191_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X7222 a_3232_43370# a_1823_45246# a_3363_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7223 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7224 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7225 a_22780_40081# en_comp a_22521_40055# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7226 a_13333_42558# a_13291_42460# a_13249_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7227 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7228 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7229 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7230 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7231 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7232 a_13661_43548# a_18780_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7233 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7234 VSS a_n2840_43914# a_n4318_39768# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7235 a_15037_44260# a_13556_45296# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7236 a_5497_46414# a_5164_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X7237 a_12749_45572# a_12549_44172# a_12649_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X7238 VSS a_22223_45572# a_19479_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7239 w_1575_34946# a_n923_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X7240 VDD a_n2438_43548# a_n133_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7241 VDD a_14815_43914# a_n2293_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7242 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7243 VDD a_n984_44318# a_n809_44244# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X7244 a_n1545_43230# a_n1991_42858# a_n1641_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7245 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7246 VDD a_22521_39511# a_22469_39537# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7247 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7248 a_11530_34132# a_18194_35068# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X7249 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7250 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7251 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7252 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7253 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7254 a_8128_46384# a_7903_47542# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X7255 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7256 VDD a_7281_43914# a_7229_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7257 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7258 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7259 VDD a_13507_46334# a_18907_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X7260 CLK_DATA a_n2833_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7261 VDD a_13904_45546# a_12594_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X7262 a_479_46660# a_33_46660# a_383_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7263 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7264 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7265 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7266 VSS a_6667_45809# a_6598_45938# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X7267 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7268 a_8568_45546# a_8953_45546# a_8697_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X7269 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7270 VREF a_19479_31679# C1_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X7271 VDD a_n881_46662# a_n1021_46688# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X7272 VDD a_2324_44458# a_15682_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7273 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7274 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7275 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7276 a_17767_44458# a_17970_44736# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X7277 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7278 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7279 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7280 VSS a_22400_42852# a_22780_40945# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7281 VDD a_n755_45592# a_133_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X7282 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7283 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7284 a_10867_43940# a_7499_43078# a_10405_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
X7285 VDD a_10723_42308# a_5742_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7286 a_16241_44734# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X7287 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7288 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7289 a_11823_42460# a_15051_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7290 a_20556_43646# a_20974_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7291 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7292 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7293 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7294 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7295 a_n3420_37440# a_n3690_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X7296 a_4574_45260# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X7297 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7298 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7299 a_13483_43940# a_13249_42308# a_13565_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7300 a_18194_35068# a_n1630_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7301 VDD a_20159_44458# a_19321_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X7302 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7303 a_n1352_44484# a_n2267_44484# a_n1699_44726# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7304 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7305 a_2583_47243# a_584_46384# a_2124_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X7306 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7307 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7308 a_22612_30879# a_22959_47212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X7309 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7310 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7311 VDD a_8349_46414# a_8379_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7312 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7313 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7314 a_n2216_40160# a_n2312_40392# a_n2302_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X7315 VSS a_14456_42282# a_5342_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7316 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7317 VSS a_768_44030# a_2711_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7318 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7319 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7320 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7321 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7322 a_n984_44318# a_n2065_43946# a_n1331_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X7323 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7324 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7325 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7326 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7327 a_5093_45028# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X7328 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7329 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7330 a_11608_46482# a_n1151_42308# a_11387_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7331 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7332 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7333 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7334 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7335 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7336 VDD a_15227_44166# a_15597_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7337 a_19862_44208# a_13747_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7338 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7339 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7340 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7341 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7342 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7343 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7344 a_19335_46494# a_18819_46122# a_19240_46482# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X7345 VDD a_2324_44458# a_6298_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7346 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7347 VSS a_1736_39587# a_1239_39587# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7348 a_n4318_38216# a_n2472_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7349 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X7350 a_8953_45546# a_8685_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7351 a_18249_42858# a_18083_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7352 a_12816_46660# a_11735_46660# a_12469_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X7353 a_19268_43646# a_13661_43548# a_19177_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.1525 ps=1.305 w=1 l=0.15
X7354 a_20256_42852# a_20202_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3125 ps=1.625 w=1 l=0.15
X7355 a_13258_32519# a_19647_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7356 VDD a_16680_45572# a_16855_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X7357 VSS a_n447_43370# a_n2129_43609# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X7358 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7359 a_20528_45572# a_19466_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X7360 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7361 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7362 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7363 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7364 a_11525_45546# a_10586_45546# a_11778_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X7365 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7366 VREF a_n3565_39590# C8_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7367 a_3537_45260# a_7287_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7368 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7369 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7370 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7371 VDD a_2711_45572# a_20107_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7372 a_16147_45260# a_17478_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X7373 a_n2109_45247# a_n2017_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7374 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7375 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7376 a_19963_31679# a_22591_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X7377 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7378 a_19610_45572# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X7379 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7380 a_5837_43172# a_3537_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7381 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7382 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7383 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7384 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7385 a_n143_45144# a_n755_45592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7386 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7387 a_n310_45572# a_n356_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X7388 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7389 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7390 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7391 VDD a_18143_47464# a_12861_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X7392 VDD a_22959_47212# a_22612_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7393 a_15015_46420# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7394 a_20596_44850# a_20159_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7395 VSS a_7227_47204# DATA[3] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7396 VSS a_7227_45028# a_7230_45938# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X7397 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7398 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7399 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7400 a_2957_45546# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X7401 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7402 VSS a_14579_43548# a_14537_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7403 VDD a_n2946_39866# a_n3565_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X7404 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7405 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X7406 VSS a_5111_44636# a_8333_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X7407 VDD a_7287_43370# a_3537_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7408 VDD a_11599_46634# a_15507_47210# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7409 VDD a_6151_47436# a_6812_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X7410 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7411 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7412 VDD COMP_P a_n1329_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X7413 VDD a_20679_44626# a_20640_44752# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7414 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7415 a_n3565_39304# a_n2946_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7416 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7417 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7418 VSS a_19321_45002# a_20567_45036# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7419 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7420 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7421 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7422 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7423 VSS a_n2472_45002# a_n2956_37592# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7424 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7425 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7426 VSS C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7427 a_10903_43370# a_13351_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7428 a_14513_46634# a_14180_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X7429 a_10949_43914# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X7430 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7431 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7432 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7433 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7434 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7435 a_10149_43396# a_5111_44636# a_9803_43646# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7436 VSS a_19431_45546# a_19365_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X7437 a_13943_43396# a_11823_42460# a_13837_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X7438 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7439 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7440 VSS a_16922_45042# a_17719_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X7441 a_16112_44458# a_14539_43914# a_16241_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X7442 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7443 C8_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X7444 VDD a_4099_45572# a_3483_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7445 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7446 a_6197_43396# a_6031_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7447 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7448 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7449 VSS a_18143_47464# a_12861_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X7450 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7451 a_7309_42852# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X7452 a_n2840_46634# a_n2661_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X7453 a_380_45546# a_n357_42282# a_603_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7454 a_18533_43940# a_18326_43940# a_18451_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7455 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7456 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7457 a_5932_42308# a_5755_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X7458 VDD a_n863_45724# a_2448_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X7459 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7460 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7461 a_16328_43172# a_n97_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7462 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7463 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7464 VSS a_n2946_38778# a_n3565_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7465 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7466 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7467 a_17583_46090# a_17715_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X7468 VDD a_13635_43156# a_9290_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7469 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7470 VDD a_n755_45592# a_8147_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X7471 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7472 VSS a_10991_42826# a_10922_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X7473 VDD a_15433_44458# a_15463_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7474 a_n2267_43396# a_n2433_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7475 a_19615_44636# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X7476 a_5732_46660# a_4651_46660# a_5385_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X7477 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X7478 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7479 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7480 a_n2840_46090# a_n2661_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X7481 VDD a_5129_47502# a_5159_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7482 a_n967_45348# a_n913_45002# a_n955_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7483 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7484 a_19006_44850# a_18248_44752# a_18443_44721# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X7485 a_n4209_39590# a_n2302_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X7486 VDD a_18817_42826# a_18707_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X7487 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7488 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7489 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7490 a_15559_46634# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X7491 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7492 a_9803_43646# a_8953_45546# a_9885_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X7493 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7494 VDD a_n2840_42282# a_n3674_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X7495 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7496 VDD a_3232_43370# a_9313_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X7497 a_13460_43230# a_12545_42858# a_13113_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7498 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7499 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7500 a_20362_44736# a_20679_44626# a_20637_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X7501 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7502 a_2713_42308# a_n913_45002# a_2725_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7503 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7504 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7505 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7506 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7507 a_768_44030# a_13487_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7508 a_16241_47178# a_16023_47582# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X7509 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7510 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7511 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7512 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7513 a_14955_43396# a_14205_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X7514 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7515 VSS C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7516 VSS a_n913_45002# a_10533_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7517 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7518 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7519 a_7466_43396# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X7520 a_n4064_40160# a_n4334_40480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7521 VDD a_6151_47436# a_5907_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X7522 a_16697_47582# a_15507_47210# a_16588_47582# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X7523 a_n2267_44484# a_n2433_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7524 a_15682_43940# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7525 VDD a_1239_39587# COMP_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7526 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7527 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7528 a_13693_46688# a_6755_46942# a_13607_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7529 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7530 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7531 VDAC_Ni a_3754_38470# a_3726_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X7532 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X7533 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X7534 VDD a_19778_44110# a_19741_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7535 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7536 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7537 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7538 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7539 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7540 a_2609_46660# a_2443_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7541 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7542 a_5708_44484# a_5257_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X7543 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7544 VSS a_n2472_43914# a_n3674_39768# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7545 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7546 a_18143_47464# a_18479_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X7547 a_5263_46660# a_4817_46660# a_5167_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7548 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7549 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7550 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7551 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7552 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7553 a_12016_45572# a_11962_45724# a_11525_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X7554 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7555 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7556 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7557 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7558 VSS a_18057_42282# a_n356_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X7559 VDD a_21671_42860# a_3422_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7560 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7561 C9_N_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7562 VDD a_8746_45002# a_8704_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X7563 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7564 a_3411_47243# a_3160_47472# a_2952_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X7565 a_n2840_46634# a_n2661_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7566 VSS a_7705_45326# a_7639_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X7567 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7568 a_n3420_39616# a_n3690_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7569 a_133_43172# a_n357_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X7570 VDD a_9396_43370# a_5111_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X7571 VSS a_167_45260# a_1423_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7572 a_743_42282# a_13661_43548# a_20301_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7573 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7574 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7575 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7576 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7577 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7578 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7579 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7580 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7581 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7582 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7583 VDD a_20512_43084# a_19987_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X7584 VSS a_n2946_37690# a_n3565_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7585 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7586 a_1891_43646# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.14825 ps=1.34 w=0.42 l=0.15
X7587 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7588 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7589 VSS a_526_44458# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7590 VSS a_n357_42282# a_17141_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X7591 a_n4318_39304# a_n2840_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7592 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7593 VIN_P EN_VIN_BSTR_P C8_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X7594 a_14485_44260# a_5807_45002# a_12465_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7595 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7596 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7597 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7598 VSS a_n1059_45260# a_8945_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X7599 a_11453_44696# a_17719_45144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X7600 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7601 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7602 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7603 a_10545_42558# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7604 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7605 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7606 a_17701_42308# a_17531_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7607 a_8292_43218# a_7765_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X7608 a_13657_42558# a_11823_42460# a_13575_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7609 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7610 a_16751_46987# a_5807_45002# a_16292_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X7611 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7612 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7613 a_10586_45546# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7614 a_n1243_44484# a_n2433_44484# a_n1352_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X7615 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7616 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7617 VDD a_3537_45260# a_4223_44672# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7618 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7619 VSS a_16855_45546# a_16789_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X7620 a_3626_43646# a_1414_42308# a_3540_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7621 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7622 VSS a_n2946_37984# a_n3565_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7623 a_45_45144# a_n143_45144# a_n37_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7624 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7625 VDD a_20107_42308# a_7174_31319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7626 a_3815_47204# a_3785_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7627 a_15567_42826# a_15743_43084# a_15953_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7628 VSS a_10341_42308# a_11554_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X7629 a_n1917_44484# a_n2267_44484# a_n2012_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7630 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7631 VCM a_5342_30871# C8_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7632 a_n83_35174# VDD EN_VIN_BSTR_P VSS sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.9
X7633 a_6755_46942# a_15015_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X7634 a_n3420_38528# a_n3690_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7635 VSS a_4791_45118# a_6640_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X7636 a_2437_43646# a_1568_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7637 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7638 VDAC_Pi a_7754_39632# VSS sky130_fd_pr__res_high_po_0p35 l=18
X7639 a_n4209_39590# a_n2302_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7640 a_9823_46155# a_9804_47204# a_9823_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X7641 a_1990_45899# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X7642 a_15743_43084# a_19339_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X7643 VDD a_5385_46902# a_5275_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X7644 a_5129_47502# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X7645 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7646 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7647 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7648 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7649 VDAC_P C1_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7650 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7651 VDD a_1177_38525# a_1343_38525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7652 a_9145_43396# a_8791_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7653 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7654 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7655 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7656 VIN_P EN_VIN_BSTR_P C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7657 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7658 VDD a_20841_46902# a_20731_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X7659 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7660 a_7276_45260# a_n1151_42308# a_7418_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X7661 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7662 VDD a_n785_47204# a_327_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X7663 a_8103_44636# a_8375_44464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7664 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7665 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7666 a_4915_47217# a_12991_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X7667 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7668 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7669 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7670 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7671 VDD a_8199_44636# a_8855_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X7672 VDD a_12549_44172# a_21115_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X7673 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7674 VDD a_2553_47502# a_2583_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7675 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7676 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7677 a_n327_42558# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X7678 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7679 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7680 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7681 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7682 a_19864_35138# VDD EN_VIN_BSTR_N VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.9
X7683 a_12800_43218# a_12089_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X7684 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7685 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7686 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7687 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7688 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7689 VSS a_20623_43914# a_20365_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X7690 VSS a_n743_46660# a_16501_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X7691 VSS a_22959_45036# a_19721_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7692 VDD a_7754_40130# a_11206_38545# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X7693 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7694 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7695 a_n4318_38680# a_n2472_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7696 VSS a_11967_42832# a_16243_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7697 a_7754_40130# RST_Z VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X7698 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7699 a_13483_43940# a_13249_42308# a_13565_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X7700 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7701 a_3363_44484# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7702 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7703 a_13249_42558# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X7704 a_18504_43218# a_17333_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X7705 VDD a_4235_43370# a_n2661_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7706 a_n4209_38502# a_n2302_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7707 a_n39_42308# a_n97_42460# a_n473_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7708 a_10210_45822# a_10180_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X7709 VSS a_11967_42832# a_20512_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7710 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7711 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7712 VSS a_n443_46116# a_2813_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7713 VSS a_4646_46812# a_7411_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7714 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7715 a_20273_46660# a_20107_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7716 VDD a_11341_43940# a_22223_43948# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7717 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X7718 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7719 a_n2312_38680# a_n2104_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7720 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7721 VDD a_12791_45546# a_12427_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X7722 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7723 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7724 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7725 a_19237_31679# a_22959_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7726 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7727 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7728 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7729 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7730 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7731 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7732 VDD a_19328_44172# a_19279_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X7733 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7734 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7735 VDD SMPL_ON_P a_n1605_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7736 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7737 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7738 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7739 VSS a_11967_42832# a_12379_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7740 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7741 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7742 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7743 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7744 VDD a_18315_45260# a_18189_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X7745 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7746 VSS a_15227_44166# a_17719_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X7747 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7748 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7749 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7750 a_10951_45334# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X7751 VSS C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7752 VDD a_2123_42473# a_1184_42692# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7753 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7754 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7755 a_4791_45118# a_4743_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X7756 a_21195_42852# a_20922_43172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X7757 a_4156_43218# a_3905_42865# a_3935_42891# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7758 a_n3420_37440# a_n3690_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7759 a_15227_44166# a_22000_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7760 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7761 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7762 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7763 a_n1899_43946# a_n2065_43946# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7764 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7765 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7766 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7767 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7768 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7769 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7770 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7771 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7772 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7773 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7774 a_n743_46660# a_n1021_46688# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X7775 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7776 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7777 VDD a_17591_47464# a_16327_47482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X7778 a_n2293_45546# a_2274_45254# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X7779 a_11633_42308# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7780 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7781 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7782 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7783 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7784 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7785 a_15682_46116# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7786 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7787 a_20205_31679# a_22223_46124# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7788 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7789 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X7790 a_n2472_46634# a_n2293_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X7791 a_2698_46116# a_2521_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X7792 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7793 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7794 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7795 VDD a_10193_42453# a_11682_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X7796 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7797 a_22705_37990# a_22521_40055# a_22609_37990# VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X7798 VDD a_n3565_38502# a_n3690_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X7799 a_5342_30871# a_14456_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7800 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7801 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7802 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7803 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7804 VDD a_8325_42308# a_8791_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7805 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7806 a_548_43396# a_n863_45724# a_458_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X7807 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7808 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7809 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7810 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7811 VDD a_n4334_39616# a_n4064_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X7812 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7813 VSS a_1756_43548# a_1467_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.182 ps=1.86 w=0.65 l=0.15
X7814 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7815 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7816 VDD a_17517_44484# a_22591_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7817 VSS a_n913_45002# a_19511_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7818 a_288_46660# a_171_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X7819 a_15312_46660# a_14976_45028# a_15009_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X7820 a_n2472_46090# a_n2293_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X7821 VSS a_22959_43948# a_17538_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7822 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7823 C9_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X7824 a_20894_47436# a_20990_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7825 VDD a_n2438_43548# a_n2157_46122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7826 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7827 VDD a_n4064_38528# a_n2216_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X7828 a_8037_42858# a_7871_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7829 a_n1736_43218# a_n1853_43023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X7830 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7831 a_n4209_37414# a_n2302_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7832 a_13527_45546# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7833 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7834 VDD a_n2472_42282# a_n4318_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X7835 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7836 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7837 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7838 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7839 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7840 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7841 a_n2661_43370# a_11415_45002# a_11361_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7842 VDD a_n2840_42826# a_n3674_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X7843 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7844 VSS a_1343_38525# a_2113_38308# VSS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X7845 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7846 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7847 VDD a_22165_42308# a_22223_42860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7848 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7849 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7850 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X7851 VSS a_14180_45002# a_13017_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X7852 a_15681_43442# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7853 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7854 C8_N_btm a_21076_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7855 VSS a_n2302_40160# a_n4315_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7856 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7857 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7858 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7859 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7860 a_8488_45348# a_8199_44636# a_8191_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X7861 a_16588_47582# a_15673_47210# a_16241_47178# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7862 a_18220_42308# a_18184_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X7863 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7864 a_n1423_46090# a_n1641_46494# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X7865 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7866 VSS a_n4334_38528# a_n4064_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X7867 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7868 VDD a_18143_47464# a_12861_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7869 a_17609_46634# a_12549_44172# a_18280_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7870 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7871 a_16115_45572# a_15599_45572# a_16020_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X7872 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7873 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7874 VSS a_19700_43370# a_n97_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7875 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7876 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7877 VSS a_2124_47436# a_1209_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X7878 VSS C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7879 VREF_GND a_17730_32519# C9_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7880 VDD a_6755_46942# a_12741_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7881 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7882 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7883 VSS a_19615_44636# a_18579_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X7884 a_15595_45028# a_15415_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X7885 a_12545_42858# a_12379_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7886 a_8791_45572# a_7499_43078# a_8697_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X7887 a_16942_47570# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X7888 a_14853_42852# a_n913_45002# a_14635_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7889 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7890 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7891 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7892 VSS a_4958_30871# a_17531_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X7893 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7894 a_8333_44056# a_4223_44672# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7895 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7896 a_6511_45714# a_4646_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7897 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7898 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7899 VDD a_10949_43914# a_10867_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X7900 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7901 a_17973_43940# a_17737_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7902 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7903 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7904 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7905 a_18494_42460# a_18907_42674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X7906 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7907 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7908 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7909 a_17061_44734# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X7910 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7911 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7912 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7913 a_n2472_46634# a_n2293_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7914 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7915 C2_P_btm a_3080_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X7916 VSS a_5267_42460# a_4905_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X7917 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7918 VSS a_n2438_43548# a_n2065_43946# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7919 VDD a_7754_40130# a_3754_38470# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X7920 VDD a_n357_42282# a_5837_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X7921 a_9159_45572# a_5937_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X7922 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7923 a_3483_46348# a_4099_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7924 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7925 VDD a_n3565_37414# a_n3690_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X7926 a_8238_44734# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X7927 VSS a_17517_44484# a_22591_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7928 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7929 VSS a_21613_42308# a_22775_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X7930 VDD a_3381_47502# a_3411_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7931 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7932 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7933 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7934 a_10150_46912# a_10467_46802# a_10425_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X7935 a_526_44458# a_3147_46376# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7936 a_n2810_45572# a_n2840_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7937 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7938 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7939 a_13675_47204# a_n1435_47204# a_13569_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X7940 a_22165_42308# a_21887_42336# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X7941 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7942 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7943 VDD a_n4064_37440# a_n2216_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X7944 VSS a_11827_44484# a_22223_45036# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7945 a_5518_44484# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X7946 a_5891_43370# a_9127_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7947 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7948 a_n3565_38502# a_n2946_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X7949 VDD a_22521_40055# a_22459_39145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7950 a_13678_32519# a_21855_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7951 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7952 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7953 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7954 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7955 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7956 VDD a_8605_42826# a_8495_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X7957 a_n2312_40392# a_n2288_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7958 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7959 a_7499_43078# a_10083_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7960 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7961 SMPL_ON_N a_21589_35634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7962 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7963 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7964 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7965 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7966 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7967 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7968 VDD a_20193_45348# a_21887_42336# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X7969 a_13076_44458# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X7970 w_1575_34946# a_n1532_35090# EN_VIN_BSTR_P w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X7971 a_18691_45572# a_18341_45572# a_18596_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7972 VSS a_n4334_37440# a_n4064_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X7973 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7974 a_3600_43914# a_1307_43914# a_3992_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X7975 a_4743_43172# a_3537_45260# a_4649_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X7976 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7977 VSS C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7978 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7979 a_11387_46155# a_11309_47204# a_11387_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X7980 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7981 a_n755_45592# a_n809_44244# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7982 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7983 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7984 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7985 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7986 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7987 a_15682_43940# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7988 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7989 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7990 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7991 a_22609_37990# a_22469_39537# CAL_P VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X7992 a_n1177_44458# a_n1352_44484# a_n998_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X7993 a_11554_42852# a_10835_43094# a_10991_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X7994 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7995 VSS a_9313_44734# a_22959_42860# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7996 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7997 VDD a_2680_45002# a_2274_45254# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X7998 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7999 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8000 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X8001 VSS C1_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8002 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8003 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X8004 VDD a_n1177_43370# a_n1190_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X8005 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8006 w_1575_34946# a_n923_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X8007 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8008 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8009 VDD a_6755_46942# a_13556_45296# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8010 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8011 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8012 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8013 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8014 VDD a_n971_45724# a_8147_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X8015 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8016 a_n785_47204# a_n815_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8017 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8018 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8019 a_n4251_40480# a_n4318_40392# a_n4334_40480# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X8020 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X8021 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8022 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8023 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8024 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8025 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8026 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X8027 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8028 a_19900_46494# a_18819_46122# a_19553_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X8029 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X8030 VSS a_n1386_35608# a_n1838_35608# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8031 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8032 a_12561_45572# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1034 ps=1 w=0.42 l=0.15
X8033 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8034 a_10083_42826# a_10518_42984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X8035 a_12359_47026# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X8036 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8037 VSS a_10355_46116# a_8199_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8038 a_3422_30871# a_21671_42860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X8039 a_5937_45572# a_5907_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8040 VDD a_16327_47482# a_17767_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X8041 a_21005_45260# a_21101_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X8042 a_12649_45572# a_10903_43370# a_12561_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X8043 VSS a_19321_45002# a_19113_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8044 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8045 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8046 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8047 a_5111_44636# a_9396_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8048 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8049 a_21297_45572# a_20107_45572# a_21188_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X8050 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8051 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8052 a_12469_46902# a_12251_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X8053 a_376_46348# a_584_46384# a_518_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X8054 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8055 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8056 a_15146_44484# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X8057 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8058 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8059 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8060 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8061 VIN_P EN_VIN_BSTR_P C6_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X8062 VSS C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8063 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8064 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8065 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8066 VDD a_n971_45724# a_n327_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X8067 a_n3565_37414# a_n2946_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X8068 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8069 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8070 a_14180_45002# a_14537_43396# a_14309_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X8071 VDD a_10193_42453# a_16237_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X8072 a_18681_44484# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X8073 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8074 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8075 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8076 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8077 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8078 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8079 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8080 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8081 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8082 a_17829_46910# a_12549_44172# a_765_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1525 ps=1.305 w=1 l=0.15
X8083 VSS a_15009_46634# a_14180_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X8084 a_2304_45348# a_2274_45254# a_2232_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X8085 a_6598_45938# a_6511_45714# a_6194_45824# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X8086 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8087 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8088 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8089 a_n3565_38216# a_n2946_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8090 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8091 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8092 a_5745_43940# a_5013_44260# a_5663_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8093 VDD a_10193_42453# a_18533_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X8094 a_5742_30871# a_10723_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8095 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8096 a_19478_44056# a_3090_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X8097 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8098 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8099 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8100 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8101 VSS a_15051_42282# a_11823_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8102 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8103 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8104 a_8192_45572# a_8199_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X8105 a_10185_46660# a_10150_46912# a_9863_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X8106 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8107 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8108 a_10835_43094# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8109 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8110 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8111 a_15890_42674# a_15764_42576# a_15486_42560# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X8112 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8113 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8114 a_n699_43396# a_n1177_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X8115 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8116 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8117 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8118 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8119 a_14033_45822# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X8120 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X8121 a_6101_44260# a_1307_43914# a_5663_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X8122 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8123 a_7927_46660# a_7577_46660# a_7832_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X8124 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8125 a_16721_46634# a_16388_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X8126 a_5826_44734# a_5147_45002# a_5518_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X8127 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8128 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8129 a_21496_47436# a_4883_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X8130 VDD a_16763_47508# a_16750_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X8131 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8132 VDD a_n746_45260# a_175_44278# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X8133 a_n443_46116# a_n901_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8134 a_2813_43396# a_3232_43370# a_2982_43646# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X8135 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8136 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8137 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8138 a_6171_42473# a_5932_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X8139 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8140 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8141 VDD a_601_46902# a_491_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X8142 VSS a_4646_46812# a_6031_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8143 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8144 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8145 VSS a_13059_46348# a_12638_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X8146 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X8147 VDD a_1123_46634# a_1110_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X8148 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8149 a_8292_43218# a_7765_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X8150 a_11787_45002# a_11963_45334# a_11915_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X8151 VSS a_584_46384# a_2998_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8152 VDD a_n2472_42826# a_n4318_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X8153 a_1667_45002# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X8154 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8155 VDD a_n3690_38528# a_n3420_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8156 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8157 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8158 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8159 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8160 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8161 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8162 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8163 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8164 a_20731_47026# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X8165 a_8062_46482# a_8016_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X8166 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8167 a_n2216_38778# a_n2312_38680# a_n2302_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X8168 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8169 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8170 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8171 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8172 a_13925_46122# a_13759_46122# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8173 VSS a_11599_46634# a_20107_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8174 VSS CLK a_8953_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X8175 a_5385_46902# a_5167_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X8176 VDD a_7499_43078# a_10729_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X8177 a_9803_43646# a_8953_45546# a_9885_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8178 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8179 VSS a_n2104_46634# a_n2312_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X8180 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8181 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8182 a_n1177_44458# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X8183 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8184 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8185 VDD a_5111_44636# a_7542_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X8186 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8187 VDD a_19256_45572# a_19431_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X8188 VDD a_6761_42308# a_7227_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X8189 a_7911_44260# a_7845_44172# a_7542_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X8190 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8191 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8192 a_n1641_43230# a_n2157_42858# a_n1736_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X8193 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8194 VDD a_19553_46090# a_19443_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X8195 a_5205_44484# a_5343_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8196 a_22400_42852# a_22223_42860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8197 a_12603_44260# a_12549_44172# a_12495_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.12675 ps=1.04 w=0.65 l=0.15
X8198 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8199 VSS a_18194_35068# a_11530_34132# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X8200 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8201 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8202 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8203 a_3638_45822# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X8204 VSS C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8205 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8206 a_17324_43396# a_16243_43396# a_16977_43638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X8207 a_5275_47026# a_4651_46660# a_5167_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X8208 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8209 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8210 a_19452_47524# a_19386_47436# a_13747_46662# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8211 a_11915_45394# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X8212 VSS a_327_47204# DATA[0] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X8213 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8214 a_14447_46660# a_n1151_42308# a_14084_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X8215 SMPL_ON_P a_n1838_35608# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8216 a_12800_43218# a_12089_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X8217 VSS a_n1613_43370# a_n1655_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8218 a_20731_47026# a_20107_46660# a_20623_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X8219 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8220 a_n1532_35090# a_n1630_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8221 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8222 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8223 VSS a_20712_42282# a_10193_42453# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X8224 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8225 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8226 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8227 VSS a_n443_42852# a_421_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X8228 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8229 a_15720_42674# a_15051_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X8230 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8231 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8232 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8233 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8234 VDD a_11599_46634# a_15599_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8235 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8236 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8237 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8238 a_n659_45366# a_n746_45260# a_n745_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X8239 a_14493_46090# a_14275_46494# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X8240 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8241 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8242 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8243 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8244 a_15682_46116# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X8245 a_n881_46662# a_14495_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X8246 a_8685_43396# a_8147_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X8247 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8248 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8249 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8250 C7_P_btm a_n4209_39304# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X8251 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8252 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8253 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8254 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8255 a_11554_42852# a_10796_42968# a_10991_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X8256 a_765_45546# a_17609_46634# a_17639_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8257 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X8258 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8259 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8260 SMPL_ON_N a_21589_35634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8261 VDD a_15803_42450# a_15764_42576# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8262 a_2063_45854# a_9863_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8263 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8264 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8265 a_19386_47436# a_19321_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X8266 a_8492_46660# a_7411_46660# a_8145_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X8267 a_1337_46436# a_1176_45822# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X8268 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8269 VSS a_4419_46090# a_4365_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8270 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8271 a_n1549_44318# a_n1899_43946# a_n1644_44306# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X8272 VDD a_9067_47204# DATA[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8273 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8274 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8275 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8276 VDAC_P C3_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8277 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8278 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8279 VSS a_6575_47204# a_9067_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X8280 a_n1331_43914# a_n1549_44318# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X8281 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8282 VDD a_3537_45260# a_5093_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X8283 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8284 a_20835_44721# a_20640_44752# a_21145_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X8285 VSS a_11189_46129# a_11608_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X8286 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8287 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8288 a_n327_42558# a_n97_42460# a_n473_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X8289 a_8147_43396# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X8290 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8291 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8292 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8293 VDD a_n3690_37440# a_n3420_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8294 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8295 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8296 a_8685_42308# a_8515_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8297 VDD a_17324_43396# a_17499_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X8298 a_19431_46494# a_18985_46122# a_19335_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X8299 VDD a_12607_44458# a_n2661_43922# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8300 a_1414_42308# a_1067_42314# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X8301 VDD a_10193_42453# a_9885_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X8302 VDD a_21356_42826# a_n357_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X8303 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8304 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8305 a_n2216_37690# a_n2810_45028# a_n2302_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X8306 VDD a_4883_46098# a_10355_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X8307 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8308 a_16977_43638# a_16759_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X8309 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8310 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8311 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8312 VSS a_n4334_40480# a_n4064_40160# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8313 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8314 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8315 a_1049_43396# a_458_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8316 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8317 VDD a_n443_42852# a_742_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8318 a_10555_43940# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X8319 VSS a_22775_42308# a_22465_38105# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8320 VSS a_n237_47217# a_8270_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8321 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8322 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8323 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8324 a_21613_42308# a_21335_42336# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X8325 a_8145_46902# a_7927_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X8326 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8327 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8328 VSS a_16019_45002# a_15903_45785# VSS sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X8329 VCM a_5342_30871# C8_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8330 VDD a_n23_45546# a_7_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X8331 VDD a_2698_46116# a_2804_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8332 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8333 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8334 a_20935_43940# a_18479_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8335 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8336 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8337 a_2713_42308# a_n755_45592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8338 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8339 VSS C2_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8340 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8341 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8342 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8343 VDD a_n699_43396# a_4743_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X8344 DATA[1] a_1431_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8345 a_17591_47464# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X8346 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8347 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8348 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8349 a_9223_42460# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X8350 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8351 a_12741_44636# a_14537_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8352 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8353 VDD a_20202_43084# a_21335_42336# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X8354 a_564_42282# a_743_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X8355 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8356 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8357 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8358 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8359 a_2684_37794# a_1736_39587# a_1736_39043# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X8360 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8361 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8362 VSS a_n2302_40160# a_n4315_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8363 a_15367_44484# a_13556_45296# a_15004_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X8364 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8365 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8366 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8367 VSS a_n452_47436# a_n815_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X8368 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8369 VDD a_2063_45854# a_9863_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X8370 VSS a_6511_45714# a_6472_45840# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8371 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8372 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8373 a_9223_42460# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X8374 VSS a_19987_42826# a_n2017_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.08775 ps=0.92 w=0.65 l=0.15
X8375 VSS a_13159_45002# a_13105_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8376 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8377 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8378 a_2981_46116# a_2804_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X8379 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8380 a_21188_45572# a_20273_45572# a_20841_45814# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X8381 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8382 a_20692_30879# a_22959_46124# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X8383 a_9028_43914# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X8384 VDD a_17715_44484# a_17737_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8385 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8386 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8387 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8388 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8389 VSS a_n2840_44458# a_n4318_40392# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X8390 VSS a_15004_44636# a_14815_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X8391 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8392 a_16759_43396# a_16243_43396# a_16664_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X8393 a_4574_45260# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X8394 a_17829_46910# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X8395 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8396 a_n4064_38528# a_n4334_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8397 VSS a_n443_46116# a_4880_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X8398 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8399 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8400 VDD a_1799_45572# a_1983_46706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X8401 VDD a_21363_45546# a_21350_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X8402 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8403 a_n4064_40160# a_n4334_40480# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X8404 VDD a_22775_42308# a_22465_38105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8405 VDAC_P C5_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8406 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8407 a_13259_45724# a_17583_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8408 C1_P_btm a_n4064_37440# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X8409 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8410 VIN_P EN_VIN_BSTR_P C4_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X8411 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8412 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8413 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8414 VSS a_327_44734# a_501_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8415 a_6575_47204# a_6545_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8416 VSS a_765_45546# a_380_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X8417 a_104_43370# a_n699_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X8418 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8419 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8420 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8421 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8422 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8423 a_n2293_42282# a_3357_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8424 VDD a_22959_42860# a_14097_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8425 a_3935_42891# a_2382_45260# a_3935_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X8426 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8427 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8428 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8429 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8430 VSS a_6171_42473# a_5379_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X8431 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8432 VDD a_9127_43156# a_5891_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8433 VDD a_n863_45724# a_327_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X8434 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8435 VDD a_8145_46902# a_8035_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X8436 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X8437 a_17141_43172# a_n1059_45260# a_16795_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X8438 VSS a_9067_47204# DATA[4] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X8439 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8440 VSS a_10193_42453# a_11897_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X8441 a_15433_44458# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X8442 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8443 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8444 VSS a_4791_45118# a_5066_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8445 VDD a_5691_45260# a_n2109_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X8446 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8447 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X8448 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8449 a_15486_42560# a_15803_42450# a_15761_42308# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X8450 a_18753_44484# a_18374_44850# a_18681_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X8451 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8452 a_n1641_43230# a_n1991_42858# a_n1736_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X8453 VDD a_1983_46706# a_n2661_46098# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8454 a_15227_46910# a_15368_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8455 a_6682_46987# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X8456 a_n1079_45724# a_n755_45592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X8457 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8458 a_12429_44172# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.118125 ps=1.04 w=0.42 l=0.15
X8459 a_1568_43370# a_1847_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8460 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X8461 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8462 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X8463 VDD a_7227_42308# a_6123_31319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8464 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8465 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8466 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8467 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8468 VSS a_1123_46634# a_584_46384# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8469 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8470 a_8952_43230# a_8037_42858# a_8605_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X8471 a_3457_43396# a_3232_43370# a_3626_43646# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X8472 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8473 a_7174_31319# a_20107_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8474 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8475 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8476 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8477 VSS a_167_45260# a_n37_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X8478 a_13490_45067# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X8479 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8480 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8481 VSS a_6171_45002# a_11909_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8482 VSS a_n2302_39866# a_n4209_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8483 a_4181_44734# a_3090_45724# a_n2497_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X8484 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8485 a_16388_46812# a_17957_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.112125 ps=0.995 w=0.65 l=0.15
X8486 VDD a_3218_45724# a_3175_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X8487 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8488 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8489 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8490 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8491 a_33_46660# a_n133_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8492 a_8283_46482# a_n1151_42308# a_7920_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X8493 VSS a_n809_44244# a_n755_45592# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8494 VDD a_15279_43071# a_14579_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8495 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8496 a_8953_45002# CLK VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8497 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8498 VDD a_16763_47508# a_5807_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8499 VDD a_310_45028# a_509_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8500 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8501 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8502 a_n23_47502# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X8503 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8504 a_3935_43218# a_3681_42891# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X8505 VDD a_10903_43370# a_10907_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X8506 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8507 a_n1099_45572# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X8508 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8509 a_14949_46494# a_13759_46122# a_14840_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X8510 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8511 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8512 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8513 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8514 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8515 VSS a_1239_39043# comp_n VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8516 VSS C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8517 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8518 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8519 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8520 VDD a_n4315_30879# a_n4334_40480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X8521 a_6851_47204# a_6491_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8522 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8523 a_13556_45296# a_6755_46942# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8524 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8525 VSS a_15227_44166# a_14539_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X8526 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8527 a_19987_42826# a_18494_42460# a_20356_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X8528 a_n4209_39304# a_n2302_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X8529 a_n2833_47464# a_n2497_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X8530 a_3524_46660# a_2609_46660# a_3177_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X8531 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8532 VREF a_n3565_39590# C8_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X8533 VSS a_6151_47436# a_6229_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X8534 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8535 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8536 VSS a_22223_47212# a_21588_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X8537 a_18533_43940# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X8538 a_14205_43396# a_13667_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X8539 a_n4064_37440# a_n4334_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8540 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8541 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8542 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8543 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8544 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8545 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X8546 a_16377_45572# a_16333_45814# a_16211_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X8547 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8548 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8549 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8550 a_10044_46482# a_n743_46660# a_9823_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X8551 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8552 a_19113_45348# a_18911_45144# a_3090_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8553 VSS a_13720_44458# a_12607_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X8554 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8555 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8556 a_n2860_37984# a_n2956_38216# a_n2946_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X8557 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8558 a_5934_30871# a_8791_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X8559 a_5837_43396# a_5111_44636# a_5147_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8560 a_2266_47570# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X8561 a_10861_46660# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X8562 VSS a_7920_46348# a_7715_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X8563 a_14383_46116# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X8564 a_2905_42968# a_742_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8565 a_2809_45348# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X8566 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8567 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8568 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8569 a_6540_46812# a_6755_46942# a_6682_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X8570 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8571 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8572 a_6709_45028# a_6431_45366# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X8573 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8574 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8575 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8576 a_8953_45002# CLK VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8577 VSS a_18494_42460# a_20193_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8578 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8579 C7_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X8580 a_n1991_42858# a_n2157_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8581 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8582 a_13249_42308# a_13070_42354# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X8583 a_n2442_46660# a_n2472_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8584 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8585 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X8586 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X8587 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8588 a_13348_45260# a_12891_46348# a_13490_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X8589 VREF_GND a_n4064_39616# C9_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8590 a_17061_44484# a_11691_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X8591 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8592 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8593 VDAC_N C6_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8594 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X8595 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8596 VDD a_18443_44721# a_18374_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X8597 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8598 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8599 VDD a_n3565_39304# a_n3690_39392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X8600 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X8601 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8602 a_1512_43396# a_n443_46116# a_1209_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X8603 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8604 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8605 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8606 VSS a_15803_42450# a_15764_42576# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8607 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8608 VDD a_22591_44484# a_17730_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8609 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8610 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8611 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8612 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8613 EN_VIN_BSTR_N a_18194_35068# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X8614 a_11901_46660# a_11735_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8615 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8616 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8617 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8618 a_21076_30879# a_22959_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8619 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8620 a_3877_44458# a_3699_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X8621 VDD a_n4064_39072# a_n2216_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X8622 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8623 a_11691_44458# a_5807_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8624 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8625 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8626 a_2813_43396# a_n443_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X8627 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8628 a_15368_46634# a_15143_45578# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X8629 VSS a_9028_43914# a_8975_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X8630 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8631 C8_N_btm a_17538_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8632 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8633 a_5093_45028# a_4558_45348# a_5009_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8634 VSS a_10193_42453# a_13921_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X8635 a_15597_42852# a_15567_42826# a_15095_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X8636 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X8637 VDD a_13059_46348# a_12839_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8638 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8639 a_3823_42558# a_3065_45002# a_3905_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X8640 VDD a_526_44458# a_5193_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X8641 a_2553_47502# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X8642 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8643 VSS a_1667_45002# a_n863_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X8644 a_1307_43914# a_2779_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8645 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8646 VDD a_n3690_38528# a_n3420_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X8647 a_16855_45546# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X8648 a_5495_43940# a_5244_44056# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X8649 VDD a_21177_47436# a_20990_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X8650 VDAC_N C4_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8651 VDD a_22365_46825# a_20202_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X8652 VSS a_19787_47423# a_19594_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X8653 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8654 VDD a_5815_47464# a_n1613_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X8655 a_n1736_46482# a_n1853_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X8656 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8657 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8658 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8659 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8660 a_5063_47570# a_4915_47217# a_4700_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X8661 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8662 VDD a_11459_47204# DATA[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X8663 a_11322_45546# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8664 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8665 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8666 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8667 a_19787_47423# START VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X8668 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8669 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8670 VDD a_9127_43156# a_9114_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X8671 a_n4251_39616# a_n4318_39768# a_n4334_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X8672 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8673 a_3754_39466# a_7754_39632# VSS sky130_fd_pr__res_high_po_0p35 l=18
X8674 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X8675 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8676 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8677 a_10384_47026# a_9863_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X8678 VSS a_11525_45546# a_11189_46129# VSS sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X8679 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8680 a_10729_43914# a_11750_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8681 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X8682 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8683 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8684 a_4921_42308# a_n913_45002# a_4933_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X8685 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8686 VSS a_8568_45546# a_8162_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X8687 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8688 a_20528_46660# a_20411_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X8689 VSS a_n23_47502# a_n89_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X8690 a_13657_42558# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X8691 VSS a_4223_44672# a_5205_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8692 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8693 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X8694 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8695 a_791_42968# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8696 a_13837_43396# a_13259_45724# a_13749_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X8697 a_19177_43646# a_17339_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X8698 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8699 a_196_42282# a_375_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X8700 a_18005_44484# a_17970_44736# a_17767_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X8701 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8702 VSS a_327_47204# DATA[0] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8703 a_11309_47204# a_11031_47542# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X8704 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8705 VDAC_P C4_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8706 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8707 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8708 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8709 VSS a_4646_46812# a_7871_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8710 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8711 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8712 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8713 VSS a_5815_47464# a_n1613_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X8714 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8715 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8716 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8717 a_18691_45572# a_18175_45572# a_18596_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X8718 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8719 a_n23_45546# a_n356_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X8720 VDAC_N C2_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8721 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8722 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8723 VDD a_n1630_35242# a_n1532_35090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8724 a_9885_42558# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X8725 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8726 VSS a_4700_47436# a_3785_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X8727 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8728 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8729 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8730 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8731 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8732 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8733 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X8734 a_4361_42308# a_3823_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X8735 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8736 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8737 VDD a_n2438_43548# a_n2157_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8738 VDD a_n2840_46634# a_n2956_39768# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X8739 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8740 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8741 VDD a_13635_43156# a_13622_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X8742 a_4817_46660# a_4651_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8743 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8744 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8745 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8746 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8747 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8748 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8749 VSS a_1307_43914# a_4156_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X8750 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X8751 a_8415_44056# a_5343_44458# a_8333_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8752 a_n1699_44726# a_n1917_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X8753 VDD a_n2946_39866# a_n3565_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8754 a_1525_44260# a_1467_44172# a_1115_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X8755 a_14976_45028# a_14797_45144# a_15060_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X8756 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8757 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8758 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X8759 VSS a_15959_42545# a_15890_42674# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X8760 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X8761 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8762 VDD a_n1838_35608# SMPL_ON_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8763 a_n3565_39304# a_n2946_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X8764 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8765 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8766 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8767 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8768 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8769 VDD a_22469_40625# a_22705_37990# VDD sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X8770 a_n2312_39304# a_n1920_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X8771 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8772 VDAC_P C6_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8773 VIN_N EN_VIN_BSTR_N C7_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X8774 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8775 VDD a_1736_39587# a_1736_39043# VDD sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X8776 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8777 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8778 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8779 VDD a_n3690_37440# a_n3420_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X8780 VDAC_N C5_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8781 VDD a_n452_44636# a_n2129_44697# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X8782 VSS a_21363_45546# a_21297_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X8783 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8784 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8785 VDD a_7112_43396# a_7287_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X8786 a_19443_46116# a_18819_46122# a_19335_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X8787 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8788 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8789 VDD a_5111_44636# a_5518_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X8790 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8791 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8792 VDD EN_VIN_BSTR_N w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X8793 a_310_45028# a_n37_45144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X8794 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8795 a_17719_45144# a_17613_45144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X8796 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8797 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8798 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8799 VDD a_12563_42308# a_5534_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8800 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8801 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8802 a_17499_43370# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X8803 a_n357_42282# a_21356_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8804 VSS a_13747_46662# a_19466_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8805 a_14112_44734# a_768_44030# a_13857_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X8806 VSS a_n2946_38778# a_n3565_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8807 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8808 VDD a_3483_46348# a_15037_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X8809 VDD a_13635_43156# a_9290_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X8810 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X8811 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8812 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X8813 VDD a_13487_47204# a_768_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8814 a_14097_32519# a_22959_42860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8815 a_8270_45546# a_n237_47217# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8816 a_3094_47570# a_2905_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X8817 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8818 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X8819 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8820 VSS a_3232_43370# a_11541_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X8821 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8822 VSS C0_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8823 a_8781_46436# a_8199_44636# a_8034_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8824 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8825 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8826 a_10533_42308# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8827 DATA[4] a_9067_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8828 a_20841_46902# a_20623_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X8829 a_13527_45546# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8830 VDAC_N C7_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8831 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8832 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8833 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8834 a_17896_45144# a_16922_45042# a_17801_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X8835 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8836 VDAC_P C8_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8837 DATA[1] a_1431_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8838 a_18817_42826# a_18599_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X8839 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8840 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8841 VDAC_N C9_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8842 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8843 VSS C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8844 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8845 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X8846 a_104_43370# a_n699_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X8847 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8848 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8849 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8850 VDAC_N VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8851 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8852 a_16211_45572# a_15765_45572# a_16115_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X8853 VSS a_20835_44721# a_20766_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X8854 a_19741_43940# a_19478_44306# a_19328_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8855 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8856 VDAC_P VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8857 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8858 VDD a_4223_44672# a_4181_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X8859 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8860 VDD a_13747_46662# a_14495_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X8861 VSS VSS sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8862 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8863 a_2487_47570# a_2063_45854# a_2124_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X8864 VSS a_10809_44734# a_22959_46124# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X8865 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8866 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8867 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8868 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8869 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8870 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8871 VDAC_N C8_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8872 VDAC_N C10_N_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8873 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8874 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8875 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8876 VDAC_P C9_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8877 VDAC_P C10_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8878 VSS a_7754_38470# a_6886_37412# VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X8879 VSS a_20567_45036# a_12549_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X8880 a_18451_43940# a_18579_44172# a_18533_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X8881 a_21359_45002# a_21513_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8882 a_13904_45546# a_13249_42308# a_14033_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X8883 VDAC_P C7_P_btm sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8884 VSS a_13661_43548# a_18587_45118# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X8885 a_6547_43396# a_6031_43396# a_6452_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
C0 VDD CLK 0.49309f
C1 a_3877_44458# a_5263_46660# 0.004328f
C2 a_4646_46812# a_5894_47026# 2.49e-19
C3 a_13661_43548# a_15227_44166# 0.805606f
C4 a_5807_45002# a_19333_46634# 5.26e-20
C5 a_13747_46662# a_18834_46812# 0.00381f
C6 a_12891_46348# a_12925_46660# 4.23e-19
C7 a_6151_47436# a_3483_46348# 2.14e-20
C8 a_n443_46116# a_4704_46090# 0.017894f
C9 C10_N_btm VIN_N 3.66034f
C10 a_18479_47436# a_11415_45002# 0.033153f
C11 a_10227_46804# a_20820_30879# 3.25e-20
C12 a_5907_46634# a_5732_46660# 0.233657f
C13 a_4817_46660# a_5275_47026# 0.031068f
C14 a_n2661_46634# a_12991_46634# 2.4e-19
C15 C9_N_btm VREF 7.369471f
C16 RST_Z EN_OFFSET_CAL 0.044122f
C17 a_n1151_42308# a_7920_46348# 0.085186f
C18 a_2063_45854# a_8953_45546# 5.65e-19
C19 a_4791_45118# a_5068_46348# 0.003762f
C20 C8_N_btm VREF_GND 2.58605f
C21 C7_N_btm VCM 1.58335f
C22 a_13507_46334# a_18280_46660# 0.004063f
C23 a_11453_44696# a_21363_46634# 0.027075f
C24 a_7_47243# a_765_45546# 1.52e-21
C25 a_14579_43548# a_16795_42852# 4.68e-21
C26 a_n97_42460# a_14635_42282# 0.077798f
C27 a_13678_32519# a_17364_32525# 0.050075f
C28 a_22223_43396# a_14209_32519# 0.001768f
C29 a_10341_43396# a_14543_43071# 6.95e-20
C30 a_15095_43370# a_5342_30871# 0.238762f
C31 a_19721_31679# EN_VIN_BSTR_N 0.005343f
C32 a_18114_32519# a_18194_35068# 6.3e-20
C33 a_14955_43396# a_15279_43071# 4.47e-19
C34 a_17023_45118# VDD 0.086861f
C35 a_13887_32519# a_22591_43396# 0.006001f
C36 a_10951_45334# a_8975_43940# 2.96e-20
C37 a_9482_43914# a_5883_43914# 0.003705f
C38 a_375_42282# a_742_44458# 1.19e-20
C39 a_2711_45572# a_17973_43940# 0.011171f
C40 a_18175_45572# a_18588_44850# 1.76e-20
C41 a_3090_45724# a_12545_42858# 0.002446f
C42 a_768_44030# a_1184_42692# 6.5e-19
C43 a_13259_45724# a_13565_43940# 3.63e-19
C44 a_1307_43914# a_2779_44458# 0.332183f
C45 a_n2661_45010# a_n89_44484# 1.47e-19
C46 a_9290_44172# a_13667_43396# 0.136018f
C47 a_8199_44636# a_10341_43396# 2.94e-19
C48 a_4185_45028# a_15781_43660# 4.43e-21
C49 a_12861_44030# a_15764_42576# 1.78e-19
C50 a_526_44458# a_766_43646# 1.14e-19
C51 a_n1925_42282# a_4905_42826# 8.84e-21
C52 SMPL_ON_P a_n4334_40480# 1.83e-19
C53 a_6945_45028# a_6197_43396# 4.56e-21
C54 a_10227_46804# a_11323_42473# 4.75e-21
C55 a_n881_46662# a_2957_45546# 2.67e-20
C56 a_20107_46660# a_20719_46660# 3.82e-19
C57 a_5807_45002# a_20062_46116# 1.96e-20
C58 a_15227_44166# a_4185_45028# 3.86e-20
C59 a_8145_46902# a_6945_45028# 3.44e-20
C60 a_n743_46660# a_11315_46155# 1.84e-19
C61 a_6755_46942# a_17715_44484# 2.63e-19
C62 a_768_44030# a_n2293_45546# 3.42e-20
C63 a_10768_47026# a_9290_44172# 3.45e-19
C64 a_15743_43084# a_15959_42545# 0.00371f
C65 a_16137_43396# a_17124_42282# 6.71e-20
C66 a_4361_42308# a_8791_42308# 0.009181f
C67 a_1847_42826# a_2351_42308# 0.120686f
C68 a_10341_43396# a_19511_42282# 1.05e-21
C69 a_5342_30871# a_14097_32519# 0.028503f
C70 a_9127_43156# a_n784_42308# 1.7e-20
C71 a_2905_42968# a_1755_42282# 2.89e-20
C72 a_743_42282# a_9885_42558# 0.006242f
C73 a_14209_32519# a_5934_30871# 0.004208f
C74 a_n630_44306# VDD 1.8e-19
C75 a_n2017_45002# a_21381_43940# 3.18e-20
C76 a_13259_45724# a_5534_30871# 0.032063f
C77 a_16019_45002# a_15493_43940# 3.46e-19
C78 a_3090_45724# a_19332_42282# 1.58e-19
C79 a_15004_44636# a_15146_44484# 0.007833f
C80 a_16979_44734# a_17061_44734# 0.171361f
C81 a_14539_43914# a_17517_44484# 6.45e-19
C82 a_n443_42852# a_n901_43156# 0.367747f
C83 a_n357_42282# a_1847_42826# 0.037548f
C84 a_526_44458# a_8292_43218# 0.02177f
C85 a_7903_47542# DATA[4] 2.01e-19
C86 a_9482_43914# a_12495_44260# 0.002157f
C87 a_5147_45002# a_5745_43940# 0.007407f
C88 a_5111_44636# a_5326_44056# 2.81e-20
C89 a_13717_47436# VDD 0.314317f
C90 a_6575_47204# DATA[3] 0.055018f
C91 a_3232_43370# a_3737_43940# 6.52e-19
C92 a_n1435_47204# RST_Z 0.179508f
C93 a_18114_32519# a_22591_44484# 0.018563f
C94 a_2437_43646# a_n97_42460# 0.201806f
C95 a_n881_46662# a_9482_43914# 1.52e-20
C96 a_17715_44484# a_8049_45260# 0.03139f
C97 a_12005_46116# a_12379_46436# 0.038694f
C98 a_10903_43370# a_12638_46436# 0.006548f
C99 a_n2293_46098# a_3218_45724# 0.007233f
C100 SMPL_ON_P a_n2661_44458# 0.002144f
C101 a_n2293_46634# a_n659_45366# 6.05e-19
C102 a_n2661_46098# a_2437_43646# 0.025093f
C103 a_6945_45028# a_5066_45546# 0.018752f
C104 a_n2497_47436# a_n1917_44484# 0.011319f
C105 a_n1076_46494# a_n1099_45572# 3.72e-20
C106 a_376_46348# a_380_45546# 0.011689f
C107 a_1176_45822# a_n2293_45546# 2.19e-20
C108 a_11415_45002# a_n443_42852# 1.47e-20
C109 a_n2312_38680# en_comp 5.01e-19
C110 a_n2438_43548# a_n913_45002# 6.79e-21
C111 a_12861_44030# a_13711_45394# 6.53e-20
C112 a_11189_46129# a_11315_46155# 0.005516f
C113 a_9290_44172# a_11601_46155# 8.23e-19
C114 a_805_46414# a_n863_45724# 8.12e-20
C115 a_2202_46116# a_n2661_45546# 6.86e-21
C116 a_5807_45002# a_5147_45002# 0.035651f
C117 a_6755_46942# a_15861_45028# 0.033041f
C118 a_14209_32519# a_11530_34132# 0.004282f
C119 a_19268_43646# VDD 0.237793f
C120 COMP_P a_4958_30871# 0.02709f
C121 a_15743_43084# RST_Z 2.97e-19
C122 a_6761_42308# a_8791_42308# 6.62e-21
C123 a_6123_31319# a_8325_42308# 6.08e-19
C124 a_7227_42308# a_8685_42308# 7.46e-20
C125 a_4190_30871# C2_P_btm 9.13e-20
C126 a_5343_44458# a_7287_43370# 2.75e-19
C127 a_16922_45042# a_16243_43396# 6.03e-22
C128 a_n913_45002# a_18083_42858# 6.19e-20
C129 a_n2017_45002# a_18249_42858# 0.545311f
C130 a_n1059_45260# a_17333_42852# 0.270324f
C131 a_13259_45724# a_19647_42308# 1.03e-19
C132 a_3422_30871# a_19862_44208# 0.030442f
C133 a_5883_43914# a_6031_43396# 0.001063f
C134 a_2998_44172# a_1525_44260# 4.65e-22
C135 a_21076_30879# a_22469_39537# 8.69e-20
C136 a_5111_44636# a_10083_42826# 0.005394f
C137 a_n443_42852# a_10533_42308# 1.11e-21
C138 a_9313_44734# a_20974_43370# 1.96e-19
C139 a_14035_46660# VDD 0.363878f
C140 a_6298_44484# a_6765_43638# 0.001141f
C141 a_n2956_39304# a_n2946_38778# 0.004064f
C142 a_n2956_38680# a_n3420_38528# 0.233147f
C143 a_n357_42282# a_15486_42560# 1.89e-20
C144 a_3232_43370# a_8387_43230# 1.01e-22
C145 a_13885_46660# RST_Z 2.35e-19
C146 a_1414_42308# a_n2661_42282# 1.17e-20
C147 a_8049_45260# a_15861_45028# 0.001507f
C148 a_5164_46348# a_3065_45002# 1.51e-21
C149 a_4704_46090# a_3537_45260# 4.91e-19
C150 a_4419_46090# a_4574_45260# 3.99e-20
C151 a_15227_44166# a_18587_45118# 0.040339f
C152 a_18834_46812# a_18911_45144# 1.88e-21
C153 a_n2442_46660# a_n2661_42834# 7.66e-20
C154 a_17583_46090# a_3357_43084# 1.42e-21
C155 a_n443_46116# a_2253_44260# 0.0014f
C156 a_n2438_43548# a_556_44484# 0.011144f
C157 a_12741_44636# a_16019_45002# 5.77e-19
C158 a_8016_46348# a_413_45260# 1.13e-21
C159 a_3483_46348# a_5111_44636# 0.340106f
C160 a_10903_43370# a_n2017_45002# 0.029479f
C161 a_4185_45028# a_4558_45348# 0.059418f
C162 a_2711_45572# a_3175_45822# 7.71e-19
C163 a_n237_47217# a_4883_46098# 0.181672f
C164 a_n4334_39392# a_n4064_38528# 7.84e-19
C165 a_n4209_39304# a_n2302_38778# 0.001019f
C166 a_1736_39587# a_2684_37794# 0.565517f
C167 a_5932_42308# C6_P_btm 3.73e-19
C168 a_6851_47204# a_n1435_47204# 2.24e-19
C169 a_9067_47204# a_11031_47542# 6.46e-21
C170 a_6151_47436# a_13487_47204# 0.038134f
C171 a_6575_47204# a_9313_45822# 0.017088f
C172 a_n3690_39392# a_n3420_38528# 7.84e-19
C173 a_n2946_39072# a_n3565_38502# 9.15e-19
C174 a_n2302_39072# a_n4209_38502# 9.15e-19
C175 a_n3420_39072# a_n3690_38528# 0.017537f
C176 a_n4064_39072# a_n4334_38528# 0.00115f
C177 a_n3565_39304# a_n2946_38778# 9.15e-19
C178 a_1736_39043# comp_n 0.005064f
C179 a_n4064_39616# a_n3565_38216# 0.028071f
C180 a_n3420_39616# a_n3420_37984# 0.047086f
C181 a_1755_42282# VDD 0.215277f
C182 a_n2109_47186# a_n2312_39304# 0.06316f
C183 a_n1920_47178# a_n2312_40392# 7.09e-19
C184 a_n3565_39590# a_n4064_37984# 0.031327f
C185 a_4915_47217# a_11599_46634# 0.015066f
C186 a_1606_42308# RST_Z 1.44945f
C187 a_19237_31679# a_13678_32519# 0.052466f
C188 a_20512_43084# a_14209_32519# 0.006512f
C189 en_comp a_7174_31319# 5.65154f
C190 a_n1099_45572# VDD 0.89411f
C191 a_n913_45002# a_22775_42308# 7.44e-19
C192 a_22485_44484# a_22591_43396# 0.025074f
C193 a_20205_31679# VIN_N 0.028894f
C194 a_14401_32519# a_17538_32519# 0.052152f
C195 a_13483_43940# a_9145_43396# 0.002944f
C196 a_9313_44734# a_18599_43230# 0.008115f
C197 a_18341_45572# a_19418_45938# 1.46e-19
C198 a_18479_45785# a_18787_45572# 0.004823f
C199 a_6598_45938# a_1423_45028# 2.06e-21
C200 a_2711_45572# a_5105_45348# 1.42e-19
C201 a_768_44030# a_2896_43646# 0.005068f
C202 a_12549_44172# a_2982_43646# 5e-19
C203 a_5937_45572# a_n2661_43922# 0.048264f
C204 a_8953_45546# a_n2661_42834# 0.019463f
C205 a_8199_44636# a_n2293_43922# 6.69e-20
C206 a_n881_46662# a_6031_43396# 1.13e-19
C207 a_n1613_43370# a_6293_42852# 0.004944f
C208 a_n2497_47436# a_n1853_43023# 4.11e-19
C209 a_584_46384# a_743_42282# 3.35e-20
C210 a_n2438_43548# a_n4318_39304# 9.42e-19
C211 a_8746_45002# a_10775_45002# 2.04e-20
C212 a_2324_44458# a_7640_43914# 3.17e-20
C213 a_10490_45724# a_8953_45002# 4.57e-19
C214 a_13163_45724# a_6171_45002# 1.51e-20
C215 a_13259_45724# a_11691_44458# 0.337184f
C216 a_10193_42453# a_10951_45334# 1.8e-20
C217 a_11530_34132# a_19120_35138# 0.480251f
C218 EN_VIN_BSTR_N a_18194_35068# 0.340036f
C219 a_n3565_37414# VCM 0.03748f
C220 VDAC_P VDD 5.19214f
C221 a_12861_44030# a_19692_46634# 0.097215f
C222 a_8912_37509# RST_Z 0.082942f
C223 a_4883_46098# a_8270_45546# 0.278829f
C224 a_15811_47375# a_16292_46812# 0.080078f
C225 a_16327_47482# a_14976_45028# 1.2e-20
C226 a_n2438_43548# a_2107_46812# 0.111283f
C227 a_n133_46660# a_948_46660# 0.102355f
C228 a_n2312_38680# a_n935_46688# 7.7e-20
C229 a_n743_46660# a_1983_46706# 0.001758f
C230 a_n4064_37440# VIN_P 0.078489f
C231 a_n881_46662# a_7715_46873# 0.02091f
C232 a_6151_47436# a_14513_46634# 3.62e-20
C233 a_n1613_43370# a_7577_46660# 3.27e-20
C234 a_n1151_42308# a_14447_46660# 0.003689f
C235 a_2952_47436# a_765_45546# 0.004287f
C236 a_n3420_37440# VREF 9.37e-19
C237 a_n2661_46634# a_n2661_46098# 0.066513f
C238 a_171_46873# a_1123_46634# 1.13e-20
C239 a_33_46660# a_383_46660# 0.20669f
C240 a_11599_46634# a_18834_46812# 0.012948f
C241 a_10227_46804# a_12816_46660# 0.253017f
C242 a_648_43396# a_685_42968# 5.58e-19
C243 a_n2661_42282# a_n3674_38680# 0.00768f
C244 a_10951_45334# VDD 0.226705f
C245 a_15095_43370# a_743_42282# 2.85e-19
C246 a_10341_43396# a_21259_43561# 0.00679f
C247 a_16243_43396# a_15743_43084# 0.600668f
C248 a_16759_43396# a_17324_43396# 7.99e-20
C249 a_16409_43396# a_18525_43370# 1.15e-20
C250 a_11967_42832# a_14113_42308# 0.003103f
C251 a_n97_42460# a_14543_43071# 7.94e-21
C252 a_2982_43646# a_5111_42852# 2.74e-20
C253 a_3626_43646# a_3935_42891# 0.002569f
C254 a_3539_42460# a_3681_42891# 4.58e-21
C255 a_4646_46812# a_9127_43156# 4.29e-21
C256 a_13017_45260# a_13105_45348# 2.63e-19
C257 a_n443_42852# a_n984_44318# 1.59e-20
C258 a_n357_42282# a_5244_44056# 2.74e-21
C259 a_n755_45592# a_3905_42865# 4.59e-20
C260 a_n2840_45002# a_n4318_40392# 4.48e-19
C261 a_2437_43646# a_742_44458# 0.081793f
C262 a_19692_46634# a_19700_43370# 4.58e-19
C263 a_n2442_46660# a_n2293_42282# 5.92e-20
C264 a_6171_45002# a_16501_45348# 2.67e-19
C265 a_n2293_46098# a_6293_42852# 0.001583f
C266 a_3218_45724# a_2675_43914# 6.54e-21
C267 a_18175_45572# a_18443_44721# 9.32e-21
C268 a_18341_45572# a_18248_44752# 3.18e-20
C269 a_18479_45785# a_18287_44626# 0.024431f
C270 a_n2956_38216# a_n4318_39768# 0.045702f
C271 a_7499_43078# a_11967_42832# 5.46e-21
C272 a_413_45260# a_22223_45036# 2.66e-19
C273 a_n2661_45010# a_n2840_44458# 3.06e-19
C274 a_8199_44636# a_n97_42460# 0.003284f
C275 a_1423_45028# a_2809_45028# 8.35e-21
C276 a_13059_46348# a_14537_43646# 0.003923f
C277 a_n443_46116# a_2713_42308# 1.17e-19
C278 a_n971_45724# a_8515_42308# 3.09e-19
C279 a_16327_47482# a_18051_46116# 2.01e-20
C280 a_n2109_47186# a_6511_45714# 5.45e-21
C281 a_n1741_47186# a_6194_45824# 3.64e-21
C282 a_2063_45854# a_1609_45822# 0.035351f
C283 a_n443_46116# a_2957_45546# 0.020365f
C284 a_n881_46662# a_5210_46482# 0.002203f
C285 a_12991_46634# a_765_45546# 1.31e-19
C286 a_n1613_43370# a_5431_46482# 6.82e-22
C287 a_4883_46098# a_12638_46436# 0.009375f
C288 a_17591_47464# a_16375_45002# 4.87e-19
C289 a_19321_45002# a_6945_45028# 0.042647f
C290 a_2107_46812# a_11133_46155# 7.92e-20
C291 a_13747_46662# a_10809_44734# 0.045104f
C292 a_n971_45724# a_2711_45572# 0.214535f
C293 a_15559_46634# a_16388_46812# 2.85e-19
C294 a_13507_46334# a_14371_46494# 0.001286f
C295 a_n743_46660# a_14275_46494# 0.006268f
C296 a_14401_32519# a_22465_38105# 8.57e-20
C297 a_3422_30871# C7_P_btm 2.94e-19
C298 a_18249_42858# a_19164_43230# 0.118759f
C299 a_3626_43646# a_15890_42674# 0.003304f
C300 a_n97_42460# a_19511_42282# 7.78e-21
C301 a_8037_42858# a_8483_43230# 2.28e-19
C302 a_526_44458# a_3681_42891# 0.002914f
C303 a_n1925_42282# a_2905_42968# 1.42e-20
C304 a_13259_45724# a_4190_30871# 0.271537f
C305 a_n2442_46660# a_n3565_39590# 0.134948f
C306 a_375_42282# a_n984_44318# 1.76e-20
C307 a_18114_32519# a_9313_44734# 1.28e-20
C308 a_n913_45002# a_12429_44172# 1.57e-21
C309 a_n1059_45260# a_13483_43940# 1.59e-20
C310 a_n2661_44458# a_8333_44734# 9.44e-20
C311 a_11691_44458# a_n2661_43922# 0.038882f
C312 a_1307_43914# a_644_44056# 1.94e-20
C313 a_3065_45002# a_3499_42826# 3.27e-19
C314 a_n2956_39768# a_n2946_39866# 0.14868f
C315 a_n443_42852# a_9885_43646# 0.001927f
C316 a_4883_46098# a_n2017_45002# 1.86e-19
C317 a_10903_43370# a_13759_46122# 8.61e-19
C318 a_1208_46090# a_1337_46436# 0.010132f
C319 a_n743_46660# a_15765_45572# 0.026376f
C320 a_7411_46660# a_8568_45546# 0.001217f
C321 a_13507_46334# a_n913_45002# 0.023897f
C322 a_17591_47464# a_413_45260# 4.35e-19
C323 a_12005_46116# a_13351_46090# 1.07e-19
C324 a_584_46384# a_626_44172# 0.450256f
C325 a_n2293_46634# a_8696_44636# 3.28e-20
C326 a_13661_43548# a_16377_45572# 1.08e-20
C327 a_22365_46825# a_8049_45260# 0.001257f
C328 a_17829_46910# a_13259_45724# 8.1e-20
C329 a_17339_46660# a_18243_46436# 0.001467f
C330 a_2905_45572# a_1307_43914# 1.08e-21
C331 a_9823_46155# a_2324_44458# 1.64e-20
C332 a_n784_42308# a_1755_42282# 0.073102f
C333 a_n1243_43396# VDD 4.56e-20
C334 a_n1630_35242# a_961_42354# 3.02e-19
C335 a_1067_42314# a_1184_42692# 0.147283f
C336 a_n863_45724# a_564_42282# 1.21e-19
C337 a_18287_44626# a_14021_43940# 2.78e-20
C338 a_9313_44734# a_17737_43940# 1.96e-20
C339 a_7499_43078# a_9114_42852# 2.49e-19
C340 a_1307_43914# a_10765_43646# 8.56e-19
C341 a_n2661_43922# a_8333_44056# 7.64e-20
C342 a_n2661_42834# a_9028_43914# 0.009687f
C343 a_22485_44484# a_22591_44484# 0.15878f
C344 a_19721_31679# a_14401_32519# 0.053967f
C345 a_5883_43914# a_6671_43940# 0.051304f
C346 a_n755_45592# a_n961_42308# 2.27e-20
C347 a_n357_42282# a_n473_42460# 0.179066f
C348 a_n2017_45002# a_5649_42852# 0.03149f
C349 a_n913_45002# a_21855_43396# 3.57e-20
C350 a_3090_45724# a_14797_45144# 9.53e-19
C351 a_14976_45028# a_14537_43396# 0.087031f
C352 a_n2497_47436# a_n1899_43946# 0.040963f
C353 a_11415_45002# a_2437_43646# 0.01065f
C354 a_12465_44636# a_9313_44734# 2.57e-20
C355 a_13259_45724# a_n443_42852# 0.022577f
C356 a_n2661_45546# a_n1079_45724# 0.008911f
C357 a_n2472_45546# a_n2293_45546# 0.171197f
C358 a_7411_46660# a_n2661_43370# 5.29e-21
C359 a_3483_46348# a_16147_45260# 6.65e-20
C360 a_20885_46660# a_3357_43084# 5.68e-19
C361 a_12741_44636# a_20719_45572# 3.43e-19
C362 a_12861_44030# a_13296_44484# 1.28e-19
C363 a_12549_44172# a_14539_43914# 0.110516f
C364 a_n2293_46634# a_n1177_44458# 1.56e-19
C365 a_2324_44458# a_10306_45572# 7.74e-19
C366 a_n2438_43548# a_n2661_44458# 0.136664f
C367 a_6945_45028# a_6977_45572# 0.001758f
C368 a_n784_42308# VDAC_P 0.005839f
C369 a_n452_47436# a_n971_45724# 0.330438f
C370 a_n1741_47186# a_n785_47204# 0.026399f
C371 a_n2109_47186# a_1209_47178# 0.226908f
C372 a_n815_47178# a_n746_45260# 0.001861f
C373 COMP_P a_22780_40945# 3.32e-19
C374 a_5934_30871# VDAC_Pi 1.75e-19
C375 a_9313_44734# a_13887_32519# 0.191376f
C376 a_19478_44306# a_19319_43548# 0.005956f
C377 a_3065_45002# a_3318_42354# 0.146272f
C378 en_comp a_5932_42308# 0.233106f
C379 a_11967_42832# a_15781_43660# 0.026392f
C380 a_n1059_45260# a_6123_31319# 0.001842f
C381 a_n913_45002# a_7227_42308# 0.052824f
C382 a_n2017_45002# a_7963_42308# 0.003883f
C383 a_17517_44484# a_17324_43396# 7.13e-22
C384 a_1241_43940# a_1443_43940# 0.092725f
C385 a_11341_43940# a_11173_43940# 1.36e-19
C386 a_19328_44172# a_19478_44056# 0.003538f
C387 a_n1925_42282# VDD 0.728242f
C388 a_10334_44484# a_10083_42826# 5.56e-20
C389 a_20708_46348# a_20567_45036# 5.99e-19
C390 a_n443_42852# a_n467_45028# 0.007314f
C391 a_3316_45546# a_3065_45002# 0.141454f
C392 a_3218_45724# a_3429_45260# 0.001528f
C393 a_n357_42282# a_5111_44636# 0.033023f
C394 a_584_46384# a_2813_43396# 0.00985f
C395 a_15227_44166# a_11967_42832# 0.132673f
C396 a_n1613_43370# a_7499_43940# 0.001731f
C397 a_n881_46662# a_6671_43940# 1.87e-19
C398 a_18189_46348# a_11691_44458# 6.35e-20
C399 a_16375_45002# a_16019_45002# 0.032313f
C400 a_768_44030# a_1443_43940# 0.003817f
C401 a_22612_30879# a_15493_43940# 1.68e-20
C402 a_n3420_39072# VIN_P 0.031754f
C403 a_12891_46348# a_13569_47204# 9.78e-20
C404 a_6575_47204# a_6540_46812# 1.87e-19
C405 a_4915_47217# a_7411_46660# 4.06e-20
C406 a_n881_46662# a_13747_46662# 0.550574f
C407 a_n310_47243# a_n2661_46634# 2.6e-19
C408 a_n4334_38528# VDD 0.385889f
C409 a_n4209_39304# VCM 0.05604f
C410 a_n3565_39304# VREF 0.098117f
C411 a_n2312_39304# a_n1925_46634# 0.071018f
C412 a_3726_37500# a_5088_37509# 0.189392f
C413 a_n3420_37984# C2_P_btm 0.03058f
C414 a_n4064_37984# C4_P_btm 0.001746f
C415 a_n1435_47204# a_4651_46660# 5.31e-20
C416 a_2063_45854# a_10249_46116# 0.078073f
C417 a_n1151_42308# a_10150_46912# 8.58e-20
C418 a_2982_43646# a_16977_43638# 3.11e-21
C419 a_3626_43646# a_16547_43609# 3.44e-21
C420 a_8685_43396# a_8423_43396# 2.34e-19
C421 a_18079_43940# a_18249_42858# 7.49e-20
C422 a_18326_43940# a_17333_42852# 7.02e-19
C423 a_18451_43940# a_18083_42858# 2.66e-22
C424 a_15493_43396# a_17595_43084# 1.05e-20
C425 a_n2293_43922# a_4921_42308# 1.79e-19
C426 a_11341_43940# a_13460_43230# 2.23e-21
C427 a_14401_32519# a_22591_43396# 0.01561f
C428 a_20974_43370# a_13887_32519# 0.033282f
C429 a_5891_43370# a_8791_42308# 7.71e-19
C430 a_19418_45938# VDD 4.6e-19
C431 a_n356_44636# a_13070_42354# 1.4e-19
C432 a_8270_45546# a_8685_43396# 0.006203f
C433 a_2711_45572# a_9313_44734# 0.036278f
C434 a_3537_45260# a_9482_43914# 3.66e-21
C435 a_7276_45260# a_6709_45028# 0.215102f
C436 w_11334_34010# a_14097_32519# 5.84e-19
C437 a_1138_42852# a_1241_43940# 0.006402f
C438 a_6469_45572# a_5883_43914# 3.18e-21
C439 a_n443_42852# a_n2661_43922# 0.045456f
C440 a_10193_42453# a_18248_44752# 0.004992f
C441 a_6598_45938# a_6109_44484# 6.27e-20
C442 a_16147_45260# a_17719_45144# 0.049848f
C443 a_13507_46334# a_20922_43172# 2.68e-20
C444 a_n2442_46660# a_n1423_42826# 4.46e-21
C445 a_3090_45724# a_7287_43370# 0.005365f
C446 a_18341_45572# a_16922_45042# 3.38e-20
C447 a_2324_44458# a_10729_43914# 2.83e-21
C448 a_8696_44636# a_16237_45028# 3.7e-19
C449 a_6431_45366# a_8191_45002# 8.63e-21
C450 a_6171_45002# a_8953_45002# 0.034987f
C451 a_3232_43370# a_10775_45002# 1.54e-20
C452 a_11823_42460# a_13076_44458# 1.17e-19
C453 a_3483_46348# a_13565_44260# 3.95e-19
C454 w_1575_34946# a_6123_31319# 0.002297f
C455 a_6755_46942# a_11901_46660# 0.587021f
C456 a_10249_46116# a_12469_46902# 8.44e-20
C457 a_n881_46662# a_4419_46090# 0.045203f
C458 a_n1613_43370# a_4704_46090# 4.05e-20
C459 a_12465_44636# a_12594_46348# 9.31e-21
C460 a_4883_46098# a_13759_46122# 0.044004f
C461 a_16327_47482# a_19900_46494# 0.216811f
C462 a_4791_45118# a_5431_46482# 0.001192f
C463 a_n2661_46098# a_765_45546# 0.0407f
C464 a_22612_30879# a_12741_44636# 1.68e-20
C465 a_21588_30879# a_22959_46660# 0.001846f
C466 a_13507_46334# a_14493_46090# 0.001974f
C467 a_10227_46804# a_18819_46122# 2.52e-20
C468 a_15811_47375# a_6945_45028# 0.037131f
C469 a_18597_46090# a_17583_46090# 4.74e-20
C470 a_11599_46634# a_10809_44734# 0.06157f
C471 a_768_44030# a_1138_42852# 0.021091f
C472 a_n2661_46634# a_11415_45002# 0.494836f
C473 a_n1435_47204# a_n1379_46482# 7.65e-21
C474 a_20916_46384# a_21076_30879# 9.97e-20
C475 a_10341_43396# a_13291_42460# 7.32e-20
C476 a_14021_43940# a_17124_42282# 4.98e-21
C477 a_4361_42308# a_21356_42826# 0.017293f
C478 a_13467_32519# a_21195_42852# 0.034759f
C479 a_20623_43914# a_13258_32519# 1.97e-21
C480 a_3080_42308# a_1755_42282# 0.047244f
C481 a_5649_42852# a_19164_43230# 5.64e-21
C482 a_18248_44752# VDD 0.251171f
C483 a_n97_42460# a_4921_42308# 3.35e-20
C484 a_10057_43914# CLK 1.02e-19
C485 a_1823_45246# a_5111_42852# 5.16e-20
C486 a_n443_42852# a_n447_43370# 0.002103f
C487 a_14537_43396# a_15433_44458# 0.018743f
C488 a_14797_45144# a_14815_43914# 3.57e-20
C489 a_n2661_43370# a_n2012_44484# 8.13e-19
C490 a_5807_45002# a_14113_42308# 1.48e-22
C491 a_13661_43548# a_13657_42558# 3.59e-20
C492 a_13249_42308# a_13829_44260# 7.14e-19
C493 a_13904_45546# a_14021_43940# 1.09e-21
C494 a_n863_45724# a_n1557_42282# 0.034373f
C495 a_4646_46812# a_1755_42282# 1.48e-21
C496 a_8696_44636# a_9672_43914# 4.19e-20
C497 a_n2661_45546# a_2982_43646# 0.007559f
C498 a_375_42282# a_n2661_43922# 0.024229f
C499 a_n755_45592# a_4093_43548# 1.18e-21
C500 a_n357_42282# a_4235_43370# 0.005266f
C501 a_3090_45724# a_13157_43218# 7.17e-19
C502 w_1575_34946# EN_VIN_BSTR_P 3.99222f
C503 a_n1925_46634# a_6511_45714# 0.028817f
C504 a_12549_44172# a_12427_45724# 0.152925f
C505 a_12891_46348# a_11823_42460# 0.033376f
C506 a_765_45546# a_17957_46116# 0.133328f
C507 a_6755_46942# a_15194_46482# 0.002244f
C508 a_1208_46090# a_1823_45246# 0.006027f
C509 a_n746_45260# a_n2661_45010# 0.400342f
C510 a_12465_44636# a_15037_45618# 2.95e-21
C511 a_5807_45002# a_7499_43078# 6.76e-20
C512 a_11901_46660# a_8049_45260# 8.89e-20
C513 a_n2293_46098# a_4704_46090# 2.86e-20
C514 a_1176_45822# a_1138_42852# 0.41217f
C515 a_11415_45002# a_8199_44636# 4.09e-20
C516 a_n881_46662# a_6469_45572# 3.11e-19
C517 a_n1613_43370# a_6905_45572# 8.54e-19
C518 a_n743_46660# a_6194_45824# 0.002138f
C519 a_1799_45572# a_n443_42852# 4.66e-20
C520 a_13507_46334# a_15903_45785# 7.77e-20
C521 a_2553_47502# a_2437_43646# 0.004656f
C522 a_12861_44030# a_18175_45572# 0.031037f
C523 a_n2497_47436# en_comp 4.47e-20
C524 a_472_46348# a_167_45260# 0.001848f
C525 a_13059_46348# a_6945_45028# 3.04e-19
C526 a_18285_46348# a_17715_44484# 2.97e-20
C527 a_19123_46287# a_17583_46090# 1.17e-20
C528 a_17829_46910# a_18189_46348# 4.65e-19
C529 a_17538_32519# a_11530_34132# 0.002953f
C530 a_12089_42308# a_12563_42308# 0.03299f
C531 a_12379_42858# a_13070_42354# 6.78e-21
C532 a_3080_42308# VDAC_P 0.009704f
C533 a_3737_43940# VDD 0.18423f
C534 a_13887_32519# a_22397_42558# 0.002537f
C535 a_5649_42852# a_21973_42336# 0.001208f
C536 a_7499_43078# a_10518_42984# 0.03265f
C537 a_20193_45348# a_20623_43914# 0.048456f
C538 a_16241_44734# a_16241_44484# 6.96e-20
C539 a_14673_44172# a_16335_44484# 6.01e-19
C540 a_11117_47542# DATA[5] 3.92e-19
C541 a_18479_45785# a_19268_43646# 0.12682f
C542 a_8953_45546# a_9885_42558# 0.024699f
C543 a_8199_44636# a_10533_42308# 4.26e-20
C544 a_22223_45036# a_22223_43948# 6.3e-19
C545 a_11827_44484# a_15493_43940# 0.010315f
C546 a_20202_43084# a_19647_42308# 6.58e-21
C547 a_3232_43370# a_3539_42460# 1.57e-22
C548 a_3537_45260# a_6031_43396# 0.034593f
C549 a_n699_43396# a_n2661_42282# 4.19e-21
C550 a_13759_47204# RST_Z 9.49e-19
C551 a_2711_45572# a_18599_43230# 4e-19
C552 a_9804_47204# CLK 5.1e-19
C553 a_n1925_42282# a_n784_42308# 0.235613f
C554 a_13259_45724# a_14635_42282# 3.09e-19
C555 a_9313_44734# a_22485_44484# 2.92e-21
C556 a_1307_43914# a_104_43370# 7.32e-21
C557 a_n2017_45002# a_8685_43396# 2.66e-19
C558 a_12594_46348# a_2711_45572# 0.009529f
C559 a_11453_44696# a_18450_45144# 3.07e-19
C560 a_6540_46812# a_5205_44484# 1.12e-21
C561 a_3483_46348# a_9049_44484# 0.117501f
C562 a_11813_46116# a_3357_43084# 1.83e-20
C563 a_15227_44166# a_20273_45572# 2.83e-19
C564 a_17829_46910# a_17478_45572# 2.26e-21
C565 a_10428_46928# a_413_45260# 1.23e-20
C566 a_5263_46660# a_5111_44636# 5.58e-20
C567 a_5257_43370# a_4558_45348# 2.74e-21
C568 a_8387_43230# VDD 0.200672f
C569 a_9803_42558# a_7174_31319# 4.88e-21
C570 a_6123_31319# a_n4315_30879# 7.4e-21
C571 a_5342_30871# C5_P_btm 9.85e-20
C572 a_5534_30871# C3_P_btm 7.69e-20
C573 a_15764_42576# a_17124_42282# 1e-19
C574 a_14113_42308# a_16197_42308# 0.002157f
C575 a_15959_42545# a_16104_42674# 0.057222f
C576 a_15803_42450# a_16522_42674# 0.089677f
C577 a_22485_44484# a_20974_43370# 0.101193f
C578 a_20512_43084# a_17538_32519# 5.55e-20
C579 a_18114_32519# a_13887_32519# 0.054996f
C580 a_n2017_45002# a_15953_42852# 9.63e-19
C581 a_n1059_45260# a_15597_42852# 0.056846f
C582 a_n913_45002# a_14853_42852# 7.37e-19
C583 a_5244_44056# a_5025_43940# 6.46e-21
C584 a_2698_46116# VDD 0.195879f
C585 a_16979_44734# a_16409_43396# 6.95e-19
C586 a_14539_43914# a_16977_43638# 0.013865f
C587 a_14673_44172# a_3626_43646# 4.56e-21
C588 a_22591_44484# a_14401_32519# 0.001482f
C589 a_19479_31679# a_14097_32519# 0.05096f
C590 a_n2497_47436# a_n1699_43638# 0.038204f
C591 SMPL_ON_P a_n2840_43370# 8.96e-19
C592 a_12861_44030# a_13829_44260# 3.01e-20
C593 a_11652_45724# a_11962_45724# 0.002072f
C594 a_2711_45572# a_15037_45618# 0.005856f
C595 a_10490_45724# a_12791_45546# 8.97e-21
C596 a_12741_44636# a_11827_44484# 0.305294f
C597 a_11415_45002# a_19113_45348# 0.012208f
C598 a_13259_45724# a_2437_43646# 3.14e-20
C599 a_18597_46090# a_20365_43914# 4.85e-21
C600 a_13507_46334# a_18451_43940# 2.1e-20
C601 a_2324_44458# a_1423_45028# 0.154419f
C602 a_11322_45546# a_11823_42460# 0.133185f
C603 a_3483_46348# a_13105_45348# 4.98e-19
C604 a_18479_47436# a_20935_43940# 0.207572f
C605 a_11453_44696# a_12429_44172# 2.89e-21
C606 a_10227_46804# a_11341_43940# 0.057378f
C607 a_4185_45028# a_n2661_43370# 0.053994f
C608 a_5937_45572# a_5837_45028# 0.043505f
C609 a_7920_46348# a_n2293_42834# 4.35e-20
C610 a_526_44458# a_3232_43370# 0.461444f
C611 a_n3565_38502# a_n4064_37440# 0.028296f
C612 a_n4064_38528# a_n3565_37414# 0.029213f
C613 a_n3420_38528# a_n3420_37440# 0.051118f
C614 a_2553_47502# a_n2661_46634# 3.46e-20
C615 a_4883_46098# a_22731_47423# 9.43e-21
C616 a_4915_47217# a_13661_43548# 3.51e-19
C617 a_9313_45822# a_12891_46348# 2.26e-20
C618 a_11459_47204# a_11309_47204# 0.183357f
C619 a_4958_30871# C6_N_btm 0.005441f
C620 a_7174_31319# C7_P_btm 9.97e-20
C621 a_11599_46634# a_n881_46662# 0.100714f
C622 a_n4064_40160# a_n1532_35090# 6.3e-20
C623 a_n785_47204# a_n743_46660# 7.46e-20
C624 a_n23_47502# a_n2438_43548# 3.57e-20
C625 a_n237_47217# a_n133_46660# 6.22e-19
C626 a_13507_46334# a_11453_44696# 0.060476f
C627 a_21811_47423# a_22223_47212# 0.031065f
C628 a_n1741_47186# a_2107_46812# 2.24e-19
C629 a_n746_45260# a_171_46873# 0.120194f
C630 a_n971_45724# a_33_46660# 5.37e-19
C631 a_1209_47178# a_n1925_46634# 3.96e-20
C632 a_16522_42674# VDD 0.077608f
C633 a_7542_44172# a_7871_42858# 6.14e-20
C634 a_15037_43940# a_15095_43370# 1.6e-19
C635 a_13527_45546# VDD 0.1902f
C636 a_20935_43940# a_4190_30871# 6.17e-21
C637 a_21115_43940# a_21259_43561# 1.55e-19
C638 a_20623_43914# a_20301_43646# 0.002259f
C639 a_1568_43370# a_1512_43396# 5.16e-20
C640 a_4905_42826# a_3539_42460# 4.19e-20
C641 a_n97_42460# a_6452_43396# 5.26e-20
C642 a_14021_43940# a_19268_43646# 0.007741f
C643 a_10180_45724# CLK 0.095799f
C644 a_3422_30871# a_21671_42860# 0.199876f
C645 a_n2293_43922# a_13291_42460# 5.94e-19
C646 a_19862_44208# a_21487_43396# 0.00184f
C647 a_20365_43914# a_743_42282# 0.001315f
C648 SMPL_ON_N a_13678_32519# 0.029315f
C649 a_6229_45572# a_n2661_43370# 4.04e-19
C650 a_13507_46334# a_17364_32525# 3.3e-20
C651 a_16223_45938# a_1307_43914# 2.89e-19
C652 a_4185_45028# a_2998_44172# 0.001414f
C653 a_n2472_45002# a_n2293_45010# 0.177252f
C654 a_n2661_45010# a_n2109_45247# 0.025907f
C655 a_n2840_45002# a_n2017_45002# 1.31e-20
C656 a_n2293_46634# a_14205_43396# 0.0055f
C657 a_17339_46660# a_11341_43940# 0.023304f
C658 a_3090_45724# a_9420_43940# 0.00133f
C659 a_10193_42453# a_16922_45042# 0.035103f
C660 a_n357_42282# a_10334_44484# 9.23e-21
C661 a_12549_44172# a_17324_43396# 6.76e-20
C662 a_3483_46348# a_3905_42865# 3.18e-20
C663 a_18819_46122# a_18579_44172# 8.68e-21
C664 a_2063_45854# a_5937_45572# 0.012248f
C665 a_n1151_42308# a_6419_46155# 0.028969f
C666 a_4700_47436# a_5068_46348# 1.09e-20
C667 a_n1435_47204# a_n1076_46494# 2.92e-21
C668 a_n2497_47436# a_2324_44458# 0.796031f
C669 a_5807_45002# a_15227_44166# 0.042586f
C670 a_13661_43548# a_18834_46812# 0.1407f
C671 a_12891_46348# a_12513_46660# 3.56e-19
C672 a_n443_46116# a_4419_46090# 0.20069f
C673 a_4791_45118# a_4704_46090# 0.001482f
C674 C9_N_btm VIN_N 1.82823f
C675 DATA[0] DATA[1] 1.62e-19
C676 a_18479_47436# a_20202_43084# 0.040227f
C677 a_4817_46660# a_5072_46660# 0.06121f
C678 a_5167_46660# a_5732_46660# 7.99e-20
C679 a_4955_46873# a_5275_47026# 7.88e-19
C680 a_n2661_46634# a_12251_46660# 0.001121f
C681 C8_N_btm VREF 3.6701f
C682 C6_N_btm VCM 0.877241f
C683 C7_N_btm VREF_GND 1.61142f
C684 a_13507_46334# a_17639_46660# 0.005147f
C685 a_11453_44696# a_20623_46660# 0.029618f
C686 VDD EN_OFFSET_CAL 0.489629f
C687 a_14579_43548# a_16414_43172# 1.1e-20
C688 a_n97_42460# a_13291_42460# 0.419357f
C689 a_2982_43646# a_3863_42891# 5.25e-19
C690 a_21855_43396# a_17364_32525# 7.4e-20
C691 a_14205_43396# a_5342_30871# 1.54e-19
C692 a_10341_43396# a_13460_43230# 3.71e-20
C693 a_12281_43396# a_12545_42858# 0.029151f
C694 a_18114_32519# EN_VIN_BSTR_N 0.187697f
C695 a_4361_42308# a_20749_43396# 3.4e-19
C696 a_15095_43370# a_15279_43071# 0.105784f
C697 a_16922_45042# VDD 1.54713f
C698 a_5649_42852# a_14209_32519# 4.85e-19
C699 a_22223_43396# a_22591_43396# 7.52e-19
C700 a_2382_45260# a_n356_44636# 2.62e-19
C701 a_2711_45572# a_17737_43940# 0.005447f
C702 a_2437_43646# a_n2661_43922# 0.033401f
C703 a_20202_43084# a_4190_30871# 4.66e-19
C704 a_3090_45724# a_12089_42308# 0.002716f
C705 a_768_44030# a_1576_42282# 6.84e-23
C706 a_1307_43914# a_949_44458# 0.028157f
C707 a_327_44734# a_7_44811# 9.51e-20
C708 a_9290_44172# a_10695_43548# 0.011352f
C709 a_8199_44636# a_9885_43646# 0.007796f
C710 a_12861_44030# a_15486_42560# 1.58e-19
C711 a_526_44458# a_4905_42826# 0.202895f
C712 a_n1925_42282# a_3080_42308# 0.897997f
C713 a_10775_45002# a_8975_43940# 4.88e-21
C714 SMPL_ON_P a_n4315_30879# 3.70932f
C715 a_10227_46804# a_10723_42308# 6.28e-21
C716 a_n881_46662# a_1848_45724# 8.39e-20
C717 a_19123_46287# a_20885_46660# 5.98e-21
C718 a_12465_44636# a_2711_45572# 0.027219f
C719 a_19321_45002# a_20009_46494# 1.68e-19
C720 a_13747_46662# a_19443_46116# 1.58e-20
C721 a_11459_47204# a_10490_45724# 3.69e-22
C722 a_n1435_47204# a_10193_42453# 9.87e-21
C723 a_2107_46812# a_10586_45546# 1.85e-19
C724 a_n2661_46634# a_13259_45724# 0.009129f
C725 a_4651_46660# a_526_44458# 6.28e-21
C726 a_7577_46660# a_6945_45028# 0.001401f
C727 a_16137_43396# a_16522_42674# 0.001223f
C728 a_15743_43084# a_15803_42450# 1.96e-19
C729 a_1847_42826# a_2123_42473# 0.004599f
C730 a_4361_42308# a_8685_42308# 0.014949f
C731 a_18083_42858# a_19273_43230# 2.56e-19
C732 a_18249_42858# a_17749_42852# 4.27e-20
C733 a_8387_43230# a_n784_42308# 2.3e-21
C734 a_743_42282# a_9377_42558# 0.00119f
C735 a_n875_44318# VDD 4.97e-20
C736 a_3537_45260# a_6671_43940# 0.00223f
C737 a_18114_32519# a_22485_44484# 0.020813f
C738 a_13259_45724# a_14543_43071# 2.13e-20
C739 a_1307_43914# a_11341_43940# 2.31482f
C740 a_1138_42852# a_1067_42314# 3.59e-19
C741 a_14539_43914# a_17061_44734# 0.020462f
C742 a_9241_44734# a_9313_44734# 5.24e-19
C743 a_16112_44458# a_17517_44484# 1.99e-21
C744 a_13249_42308# a_13837_43396# 8.11e-20
C745 a_n755_45592# a_685_42968# 2.82e-19
C746 a_n357_42282# a_791_42968# 0.009083f
C747 a_n443_42852# a_n1641_43230# 8.55e-20
C748 a_526_44458# a_7573_43172# 0.001584f
C749 a_7227_47204# DATA[4] 1.74e-19
C750 a_9482_43914# a_11816_44260# 0.003029f
C751 a_13059_46348# a_14456_42282# 0.001136f
C752 a_4185_45028# COMP_P 3.46e-20
C753 a_n863_45724# a_3935_42891# 4.1e-20
C754 a_10193_42453# a_15743_43084# 0.027326f
C755 a_13381_47204# RST_Z 2.25e-20
C756 a_7903_47542# DATA[3] 0.01066f
C757 a_n1435_47204# VDD 0.267875f
C758 a_1823_45246# a_n2661_45546# 0.181403f
C759 a_5807_45002# a_4558_45348# 9.02e-19
C760 a_6755_46942# a_8696_44636# 0.04097f
C761 a_n2293_46634# a_n967_45348# 0.007362f
C762 a_17583_46090# a_8049_45260# 5.45e-20
C763 a_12005_46116# a_12005_46436# 0.009374f
C764 a_10903_43370# a_12379_46436# 2.66e-19
C765 a_n2293_46098# a_2957_45546# 0.00827f
C766 SMPL_ON_P a_n4318_40392# 0.039594f
C767 a_12359_47026# a_11823_42460# 5.24e-20
C768 a_22612_30879# a_413_45260# 0.11791f
C769 a_1799_45572# a_2437_43646# 0.002971f
C770 a_n2497_47436# a_n1699_44726# 0.012807f
C771 a_n901_46420# a_n1099_45572# 0.002063f
C772 a_768_44030# a_7229_43940# 0.042486f
C773 a_15227_44166# a_15143_45578# 0.010748f
C774 a_n2312_38680# a_n2956_37592# 0.048307f
C775 a_2063_45854# a_11691_44458# 4.35e-20
C776 a_n2438_43548# a_n1059_45260# 3.13e-20
C777 a_9290_44172# a_11315_46155# 0.001284f
C778 a_472_46348# a_n863_45724# 1.63e-20
C779 a_15743_43084# VDD 0.572249f
C780 a_14097_32519# a_13258_32519# 0.051815f
C781 a_13887_32519# EN_VIN_BSTR_N 0.031746f
C782 a_6761_42308# a_8685_42308# 3.39e-20
C783 a_7227_42308# a_8325_42308# 4.47e-20
C784 a_4190_30871# C3_P_btm 1.1e-19
C785 a_18579_44172# a_11341_43940# 0.030765f
C786 a_5343_44458# a_6547_43396# 3.36e-21
C787 a_n1059_45260# a_18083_42858# 0.021784f
C788 a_n913_45002# a_17701_42308# 1.16e-19
C789 a_n2017_45002# a_17333_42852# 0.314084f
C790 a_10193_42453# a_1606_42308# 1.31e-19
C791 a_13259_45724# a_19511_42282# 7.13e-20
C792 a_21398_44850# a_19862_44208# 9.39e-19
C793 a_4223_44672# a_8147_43396# 0.001199f
C794 a_2479_44172# a_3499_42826# 0.004494f
C795 a_895_43940# a_2537_44260# 7.13e-20
C796 a_21076_30879# a_22821_38993# 1.66e-19
C797 a_5111_44636# a_8952_43230# 1.01e-19
C798 a_11691_44458# a_14955_43396# 6.92e-19
C799 a_9313_44734# a_14401_32519# 0.00363f
C800 a_13885_46660# VDD 0.499249f
C801 a_n357_42282# a_15051_42282# 3.44e-19
C802 a_n2956_39304# a_n3420_38528# 0.001161f
C803 a_n2956_38680# a_n3690_38528# 0.015398f
C804 a_6298_44484# a_6197_43396# 0.002222f
C805 a_21137_46414# a_21188_45572# 1.5e-20
C806 a_6945_45028# a_21363_45546# 2.51e-20
C807 a_3483_46348# a_5147_45002# 0.363215f
C808 a_18189_46348# a_2437_43646# 3.03e-20
C809 a_8049_45260# a_8696_44636# 0.005215f
C810 a_11415_45002# a_16751_45260# 0.009485f
C811 a_4419_46090# a_3537_45260# 0.003458f
C812 a_4185_45028# a_4574_45260# 0.006766f
C813 a_15227_44166# a_18315_45260# 0.272047f
C814 a_n2956_39768# a_n2293_43922# 6.42e-20
C815 a_n2661_46634# a_n2661_43922# 1.58e-19
C816 a_15682_46116# a_3357_43084# 3.34e-20
C817 a_n1151_42308# a_n2661_42282# 1.58e-19
C818 a_n755_45592# a_7499_43078# 0.157526f
C819 a_n2438_43548# a_484_44484# 7.2e-20
C820 a_12741_44636# a_15595_45028# 3.6e-19
C821 a_1823_45246# a_5205_44484# 4.61e-19
C822 a_13507_46334# a_19237_31679# 6.88e-20
C823 a_1736_39587# a_1177_38525# 0.001279f
C824 a_n4209_39304# a_n4064_38528# 0.029379f
C825 a_n4209_39590# a_n2302_37984# 7.57e-20
C826 a_5932_42308# C7_P_btm 0.003981f
C827 a_6491_46660# a_n1435_47204# 7.35e-19
C828 a_9067_47204# a_9863_47436# 0.007473f
C829 a_6151_47436# a_12861_44030# 0.39397f
C830 a_7903_47542# a_9313_45822# 3.57e-20
C831 a_n3690_39392# a_n3690_38528# 0.050585f
C832 a_1239_39043# comp_n 0.38743f
C833 a_n3420_39072# a_n3565_38502# 0.034254f
C834 a_n4064_39072# a_n4209_38502# 0.030674f
C835 a_n3565_39304# a_n3420_38528# 0.028052f
C836 a_n4064_39616# a_n4334_38304# 8e-19
C837 a_1606_42308# VDD 0.631207f
C838 a_n2109_47186# a_n2312_40392# 0.005539f
C839 a_n2288_47178# a_n2312_39304# 0.01565f
C840 a_12429_44172# a_9145_43396# 1.63e-19
C841 en_comp a_20712_42282# 4.59e-20
C842 a_380_45546# VDD 0.154763f
C843 a_n913_45002# a_21613_42308# 0.259761f
C844 a_22485_44484# a_13887_32519# 5.15e-23
C845 a_20512_43084# a_22591_43396# 5.83e-19
C846 a_10807_43548# a_10695_43548# 0.159782f
C847 a_20193_45348# a_14097_32519# 4.63e-20
C848 a_14401_32519# a_20974_43370# 0.118041f
C849 a_9313_44734# a_18817_42826# 0.003505f
C850 a_17478_45572# a_2437_43646# 1.42e-21
C851 a_18175_45572# a_18787_45572# 3.82e-19
C852 a_16147_45260# a_18953_45572# 2.59e-20
C853 a_10227_46804# a_10341_43396# 0.188948f
C854 a_6667_45809# a_1423_45028# 8.66e-22
C855 a_768_44030# a_1987_43646# 3.01e-19
C856 a_12791_45546# a_6171_45002# 9.74e-21
C857 a_8199_44636# a_n2661_43922# 0.04879f
C858 a_5937_45572# a_n2661_42834# 0.043505f
C859 a_n1613_43370# a_6031_43396# 0.308901f
C860 a_n2497_47436# a_n2157_42858# 1.22e-19
C861 a_n2438_43548# a_n2840_43370# 0.00955f
C862 a_5066_45546# a_6298_44484# 7.32e-21
C863 a_526_44458# a_8975_43940# 3.81e-21
C864 a_10193_42453# a_10775_45002# 1.13e-21
C865 a_2324_44458# a_6109_44484# 0.101116f
C866 a_8746_45002# a_8953_45002# 0.257529f
C867 a_10180_45724# a_10951_45334# 6.34e-19
C868 a_10586_45546# a_n2661_44458# 9.07e-20
C869 a_16375_45002# a_11827_44484# 2.06e-19
C870 a_11530_34132# a_18194_35068# 0.4004f
C871 a_n3565_37414# VREF_GND 0.0061f
C872 a_8912_37509# VDD 18.3523f
C873 a_13717_47436# a_19692_46634# 3.9e-20
C874 a_12861_44030# a_19466_46812# 0.004139f
C875 a_16327_47482# a_3090_45724# 1.00134f
C876 a_15811_47375# a_15559_46634# 0.018669f
C877 a_n743_46660# a_2107_46812# 0.72755f
C878 a_n2438_43548# a_948_46660# 0.054839f
C879 a_n133_46660# a_1123_46634# 0.043619f
C880 a_n1925_46634# a_288_46660# 0.003365f
C881 VDAC_N RST_Z 0.154233f
C882 a_6151_47436# a_14180_46812# 6.21e-19
C883 a_n1613_43370# a_7715_46873# 8.67e-20
C884 a_2553_47502# a_765_45546# 0.003113f
C885 a_n1151_42308# a_14226_46660# 2.85e-20
C886 a_n881_46662# a_7411_46660# 0.025876f
C887 a_n2661_46634# a_1799_45572# 0.0082f
C888 a_n2956_39768# a_n2661_46098# 1.22e-20
C889 a_171_46873# a_383_46660# 3.12e-19
C890 a_33_46660# a_601_46902# 0.17072f
C891 a_15507_47210# a_16292_46812# 3.28e-19
C892 a_11599_46634# a_17609_46634# 5.91e-20
C893 a_10227_46804# a_12991_46634# 0.349162f
C894 a_10775_45002# VDD 0.148349f
C895 a_n2661_42282# a_n2840_42282# 0.173771f
C896 a_14205_43396# a_743_42282# 2.22e-20
C897 a_10341_43396# a_19177_43646# 2.93e-19
C898 a_2675_43914# a_2713_42308# 8.11e-22
C899 a_n3674_39768# a_n1630_35242# 1.64e-19
C900 a_16243_43396# a_18783_43370# 2.36e-21
C901 a_16137_43396# a_15743_43084# 0.029757f
C902 a_16977_43638# a_17324_43396# 0.051162f
C903 a_16409_43396# a_18429_43548# 1.76e-19
C904 a_n97_42460# a_13460_43230# 1.61e-19
C905 a_2982_43646# a_4520_42826# 3.49e-20
C906 a_3626_43646# a_3681_42891# 0.001623f
C907 a_n2840_45002# a_n2840_44458# 0.025171f
C908 a_18597_46090# a_22400_42852# 2.28e-21
C909 a_4646_46812# a_8387_43230# 4.44e-20
C910 a_3483_46348# a_4093_43548# 4.56e-21
C911 a_n443_42852# a_n809_44244# 1.06e-19
C912 a_n357_42282# a_3905_42865# 0.059842f
C913 a_17339_46660# a_10341_43396# 0.023552f
C914 a_n755_45592# a_3600_43914# 7.02e-21
C915 a_6171_45002# a_16405_45348# 2.48e-19
C916 a_n2293_46098# a_6031_43396# 1.36e-21
C917 a_1423_45028# a_2448_45028# 6.07e-21
C918 a_18479_45785# a_18248_44752# 0.002693f
C919 a_18175_45572# a_18287_44626# 2.34e-19
C920 a_n971_45724# a_5934_30871# 7.07e-19
C921 a_19692_46634# a_19268_43646# 5.49e-20
C922 a_11453_44696# a_10586_45546# 0.005294f
C923 a_2124_47436# a_2277_45546# 5.88e-21
C924 a_n443_46116# a_1848_45724# 0.041711f
C925 a_2063_45854# a_n443_42852# 8.99e-20
C926 a_584_46384# a_1609_45822# 1.57e-20
C927 a_n881_46662# a_4365_46436# 5.52e-19
C928 a_14084_46812# a_14226_46660# 0.007833f
C929 a_12251_46660# a_765_45546# 0.001931f
C930 a_4883_46098# a_12379_46436# 0.007631f
C931 a_2107_46812# a_11189_46129# 1.06e-20
C932 a_13661_43548# a_10809_44734# 0.043589f
C933 a_19452_47524# a_6945_45028# 4.72e-19
C934 a_15559_46634# a_13059_46348# 0.167936f
C935 a_n743_46660# a_14493_46090# 0.007037f
C936 a_11599_46634# a_19443_46116# 0.026712f
C937 a_13507_46334# a_14180_46482# 0.001677f
C938 a_4190_30871# a_19326_42852# 1.16e-19
C939 a_3422_30871# C8_P_btm 4.06e-19
C940 a_18817_42826# a_18599_43230# 0.209641f
C941 a_18083_42858# a_19987_42826# 6.28e-21
C942 a_18249_42858# a_19339_43156# 0.042415f
C943 a_17333_42852# a_19164_43230# 3.85e-20
C944 a_3626_43646# a_15959_42545# 0.005102f
C945 a_5111_42852# a_5193_42852# 0.171361f
C946 a_8037_42858# a_8292_43218# 0.064178f
C947 a_2382_45260# a_3820_44260# 0.001415f
C948 a_526_44458# a_2905_42968# 0.007721f
C949 a_4185_45028# a_4743_43172# 5.73e-19
C950 a_n443_42852# a_14955_43396# 0.076467f
C951 a_5343_44458# a_n356_44636# 5.46e-20
C952 a_n2661_44458# a_8238_44734# 5.96e-19
C953 a_n2442_46660# a_n4334_39616# 6.16e-20
C954 a_n2017_45002# a_13483_43940# 1.15e-21
C955 a_n913_45002# a_11750_44172# 9.36e-22
C956 a_11691_44458# a_n2661_42834# 0.018854f
C957 a_1307_43914# a_175_44278# 8.72e-21
C958 a_7229_43940# a_7845_44172# 1.1e-20
C959 a_n2956_39768# a_n3420_39616# 0.233256f
C960 a_2324_44458# a_15567_42826# 7.25e-19
C961 a_9569_46155# a_2324_44458# 5.17e-20
C962 a_472_46348# a_1431_46436# 6.01e-19
C963 a_n743_46660# a_15903_45785# 2.48e-19
C964 a_7411_46660# a_8162_45546# 4.69e-20
C965 a_4791_45118# a_9482_43914# 6.76e-20
C966 a_765_45546# a_13259_45724# 0.036082f
C967 a_17339_46660# a_18147_46436# 0.002157f
C968 a_13507_46334# a_n1059_45260# 3.96e-20
C969 a_16588_47582# a_413_45260# 8.28e-20
C970 a_10903_43370# a_13351_46090# 0.181897f
C971 a_12005_46116# a_12594_46348# 0.065075f
C972 a_584_46384# a_501_45348# 1.78e-19
C973 a_13747_46662# a_16842_45938# 3.67e-19
C974 a_13661_43548# a_16211_45572# 6.84e-20
C975 a_2747_46873# a_2437_43646# 0.003933f
C976 a_6755_46942# a_7227_45028# 2.07e-20
C977 a_6969_46634# a_6598_45938# 6.03e-19
C978 a_22959_42860# a_13258_32519# 7.81e-21
C979 a_564_42282# a_961_42354# 0.003943f
C980 a_n784_42308# a_1606_42308# 15.027599f
C981 COMP_P a_n39_42308# 5.96e-21
C982 a_3539_42460# VDD 0.363092f
C983 a_21195_42852# a_21335_42336# 8.75e-20
C984 a_n1630_35242# a_1184_42692# 0.003096f
C985 a_1067_42314# a_1576_42282# 0.017282f
C986 a_3626_43646# RST_Z 4.03e-19
C987 a_20512_43084# a_22591_44484# 2.48e-20
C988 a_n913_45002# a_4361_42308# 0.250497f
C989 a_18248_44752# a_14021_43940# 1.74e-20
C990 a_n2293_42834# a_8147_43396# 7.84e-19
C991 a_9313_44734# a_15682_43940# 1.54e-19
C992 a_7499_43078# a_10793_43218# 3.95e-19
C993 a_n755_45592# a_n1329_42308# 2.67e-21
C994 a_1307_43914# a_10341_43396# 2.19e-19
C995 a_14539_43914# a_15301_44260# 6.38e-21
C996 a_n2661_42834# a_8333_44056# 0.007771f
C997 a_18114_32519# a_14401_32519# 0.087478f
C998 a_5883_43914# a_5829_43940# 0.009634f
C999 a_n357_42282# a_n961_42308# 7.65e-19
C1000 a_8049_45260# a_7227_45028# 3.6e-19
C1001 a_12594_46348# a_14033_45822# 0.001526f
C1002 a_15227_44166# a_13017_45260# 5.47e-20
C1003 a_3090_45724# a_14537_43396# 0.530123f
C1004 a_n2497_47436# a_n1761_44111# 0.045728f
C1005 a_8953_45546# a_8696_44636# 0.022578f
C1006 a_20202_43084# a_2437_43646# 0.129143f
C1007 a_11415_45002# a_21513_45002# 0.050445f
C1008 a_526_44458# a_10193_42453# 1.72e-19
C1009 a_5257_43370# a_n2661_43370# 0.027779f
C1010 a_n2472_45546# a_n2956_38216# 0.157892f
C1011 a_n2661_45546# a_n2293_45546# 0.077901f
C1012 a_n1613_43370# a_n1809_44850# 0.012196f
C1013 a_20719_46660# a_3357_43084# 0.001371f
C1014 a_4915_47217# a_11967_42832# 1.34e-21
C1015 a_12891_46348# a_14539_43914# 3.29e-20
C1016 a_12549_44172# a_16112_44458# 1.91e-20
C1017 a_2324_44458# a_10216_45572# 9.53e-19
C1018 a_n2438_43548# a_n4318_40392# 0.001259f
C1019 a_n743_46660# a_n2661_44458# 8.9e-21
C1020 a_6945_45028# a_6905_45572# 7.62e-19
C1021 a_10227_46804# a_n2293_43922# 1.57e-19
C1022 a_22400_42852# a_22705_37990# 1.13e-20
C1023 a_5742_30871# a_n4209_38216# 4.02e-21
C1024 COMP_P a_22469_40625# 0.120018f
C1025 a_n815_47178# a_n971_45724# 0.013837f
C1026 a_n1741_47186# a_n23_47502# 0.007866f
C1027 a_n2109_47186# a_327_47204# 0.041762f
C1028 SMPL_ON_P a_n237_47217# 4.88e-23
C1029 a_n1920_47178# a_n785_47204# 1.29e-19
C1030 a_9313_44734# a_22223_43396# 1.02e-20
C1031 a_2382_45260# a_3823_42558# 0.058499f
C1032 a_3065_45002# a_2903_42308# 2.87e-19
C1033 a_11967_42832# a_15681_43442# 1.86e-19
C1034 a_18579_44172# a_10341_43396# 0.023217f
C1035 a_n913_45002# a_6761_42308# 0.350952f
C1036 a_n1059_45260# a_7227_42308# 1.26e-19
C1037 a_n2017_45002# a_6123_31319# 0.007053f
C1038 a_17517_44484# a_17499_43370# 1.98e-19
C1039 a_11341_43940# a_10867_43940# 3.41e-19
C1040 a_15493_43396# a_19319_43548# 0.120111f
C1041 a_526_44458# VDD 2.35177f
C1042 a_10157_44484# a_10083_42826# 1.72e-19
C1043 a_13259_45724# a_16751_45260# 1.84e-20
C1044 a_3483_46348# a_10157_44484# 2.51e-21
C1045 a_4185_45028# a_5883_43914# 4.3e-21
C1046 a_10227_46804# a_n97_42460# 0.18445f
C1047 a_5164_46348# a_5518_44484# 7.19e-19
C1048 a_3503_45724# a_2382_45260# 3.72e-20
C1049 a_3218_45724# a_3065_45002# 0.002508f
C1050 a_n357_42282# a_5147_45002# 1.06e-21
C1051 a_3316_45546# a_2680_45002# 0.050127f
C1052 a_4791_45118# a_6031_43396# 4.86e-20
C1053 a_n443_46116# a_1512_43396# 0.010064f
C1054 a_584_46384# a_2437_43396# 8.66e-20
C1055 a_n1613_43370# a_6671_43940# 0.03314f
C1056 a_8791_45572# a_8696_44636# 1.87e-19
C1057 a_10907_45822# a_12649_45572# 4.44e-21
C1058 a_17715_44484# a_11691_44458# 0.036149f
C1059 a_11189_46129# a_n2661_44458# 2.93e-21
C1060 a_15682_46116# a_16237_45028# 3.39e-20
C1061 a_18189_46348# a_19113_45348# 2.31e-19
C1062 a_768_44030# a_1241_43940# 0.003504f
C1063 a_21588_30879# a_15493_43940# 1.53e-20
C1064 a_n4064_37440# VDAC_P 3.73e-19
C1065 a_4915_47217# a_5257_43370# 8.75e-20
C1066 a_n881_46662# a_13661_43548# 3.79e-20
C1067 a_2747_46873# a_n2661_46634# 0.019513f
C1068 a_n4209_38502# VDD 0.811731f
C1069 a_n4209_39304# VREF_GND 0.02097f
C1070 a_n237_47217# a_8035_47026# 1.8e-20
C1071 a_n2312_39304# a_n2312_38680# 0.082563f
C1072 a_3726_37500# a_4338_37500# 0.212154f
C1073 a_11453_44696# a_n743_46660# 0.004481f
C1074 a_n4064_37984# C5_P_btm 1.01e-19
C1075 a_n3420_37984# C3_P_btm 0.001771f
C1076 a_n1435_47204# a_4646_46812# 4.92e-20
C1077 a_2063_45854# a_10554_47026# 0.002948f
C1078 a_n1151_42308# a_9863_46634# 2.6e-19
C1079 a_4791_45118# a_7715_46873# 1.8e-19
C1080 a_3626_43646# a_16243_43396# 5.34e-20
C1081 a_2982_43646# a_16409_43396# 5.61e-21
C1082 a_8685_43396# a_8317_43396# 2.29e-19
C1083 a_18079_43940# a_17333_42852# 1.33e-20
C1084 a_18326_43940# a_18083_42858# 1e-20
C1085 a_9396_43370# a_10341_43396# 5.02e-19
C1086 a_11341_43940# a_13635_43156# 3.77e-20
C1087 a_20974_43370# a_22223_43396# 0.04256f
C1088 a_14401_32519# a_13887_32519# 0.07508f
C1089 a_5891_43370# a_8685_42308# 0.048111f
C1090 a_21845_43940# a_13678_32519# 1.2e-19
C1091 a_17668_45572# VDD 9.68e-19
C1092 a_n356_44636# a_12563_42308# 2.77e-19
C1093 a_7276_45260# a_7229_43940# 0.322065f
C1094 a_5205_44484# a_6709_45028# 0.095031f
C1095 a_n443_42852# a_n2661_42834# 0.076984f
C1096 a_10193_42453# a_17970_44736# 9.16e-19
C1097 a_6511_45714# a_7640_43914# 3.14e-19
C1098 a_16375_45002# a_18005_44484# 8.14e-20
C1099 a_16147_45260# a_17613_45144# 0.028566f
C1100 a_13507_46334# a_19987_42826# 6.44e-20
C1101 a_768_44030# a_5755_42852# 2.35e-21
C1102 a_3090_45724# a_6547_43396# 0.003527f
C1103 a_18479_45785# a_16922_45042# 0.02321f
C1104 a_15861_45028# a_11691_44458# 2.17e-19
C1105 a_3232_43370# a_8953_45002# 0.012103f
C1106 a_6171_45002# a_8191_45002# 0.024424f
C1107 a_17339_46660# a_n97_42460# 0.001432f
C1108 a_11823_42460# a_12883_44458# 0.026633f
C1109 a_n1613_43370# a_10796_42968# 1.91e-20
C1110 a_14955_47212# a_10809_44734# 9.82e-20
C1111 a_15507_47210# a_6945_45028# 0.04755f
C1112 a_2063_45854# a_6633_46155# 4.03e-21
C1113 a_6755_46942# a_11813_46116# 0.028837f
C1114 a_10249_46116# a_11901_46660# 3.57e-19
C1115 a_n881_46662# a_4185_45028# 0.001491f
C1116 a_n1613_43370# a_4419_46090# 2.2e-19
C1117 a_16327_47482# a_20075_46420# 0.270434f
C1118 a_n443_46116# a_4365_46436# 1.01e-19
C1119 a_4791_45118# a_5210_46482# 1.81e-19
C1120 a_21588_30879# a_12741_44636# 0.001298f
C1121 a_1799_45572# a_765_45546# 0.225248f
C1122 a_22612_30879# a_20820_30879# 0.061094f
C1123 a_4883_46098# a_13351_46090# 0.006426f
C1124 a_13507_46334# a_13925_46122# 0.003355f
C1125 a_18143_47464# a_18189_46348# 1.76e-19
C1126 a_11453_44696# a_11189_46129# 2.99e-20
C1127 a_18597_46090# a_15682_46116# 1.97e-20
C1128 a_8035_47026# a_8270_45546# 7.91e-21
C1129 a_n1435_47204# a_n1545_46494# 4.84e-20
C1130 a_21487_43396# a_21671_42860# 3.61e-19
C1131 a_4361_42308# a_20922_43172# 0.00325f
C1132 a_13467_32519# a_21356_42826# 0.001409f
C1133 a_15095_43370# a_15785_43172# 0.002407f
C1134 a_20269_44172# a_20107_42308# 3.94e-19
C1135 a_20365_43914# a_13258_32519# 6.32e-21
C1136 a_19862_44208# a_20712_42282# 3.07e-21
C1137 a_4699_43561# a_1755_42282# 2.85e-21
C1138 a_n1557_42282# a_961_42354# 1.02e-20
C1139 a_3080_42308# a_1606_42308# 4.87174f
C1140 a_3539_42460# a_n784_42308# 2.97e-20
C1141 a_5649_42852# a_19339_43156# 2.62e-21
C1142 a_17970_44736# VDD 0.27753f
C1143 a_10440_44484# CLK 0.013272f
C1144 a_1823_45246# a_4520_42826# 0.053569f
C1145 a_n443_42852# a_n1352_43396# 2.4e-19
C1146 a_14537_43396# a_14815_43914# 0.015948f
C1147 a_1307_43914# a_n2293_43922# 0.022859f
C1148 a_n2312_39304# a_7174_31319# 4.73e-21
C1149 a_13249_42308# a_13565_44260# 0.002149f
C1150 SMPL_ON_N a_22775_42308# 9.64e-21
C1151 a_8696_44636# a_9028_43914# 4.56e-21
C1152 a_375_42282# a_n2661_42834# 0.035547f
C1153 a_n357_42282# a_4093_43548# 0.002194f
C1154 a_3090_45724# a_12991_43230# 0.001405f
C1155 w_1575_34946# a_n923_35174# 37.7438f
C1156 a_n1925_46634# a_6472_45840# 9.08e-19
C1157 a_768_44030# a_11652_45724# 4.54e-22
C1158 a_12549_44172# a_11962_45724# 0.034917f
C1159 a_12891_46348# a_12427_45724# 1.55e-19
C1160 a_17339_46660# a_17957_46116# 0.098952f
C1161 a_6755_46942# a_14949_46494# 5.41e-19
C1162 a_765_45546# a_18189_46348# 0.013467f
C1163 a_805_46414# a_1823_45246# 6.82e-20
C1164 a_472_46348# a_2202_46116# 3.26e-20
C1165 a_n971_45724# a_n2661_45010# 0.017233f
C1166 SMPL_ON_P a_n2017_45002# 1.46e-21
C1167 a_3524_46660# a_3503_45724# 8.08e-21
C1168 a_5807_45002# a_8568_45546# 7.37e-22
C1169 a_11813_46116# a_8049_45260# 0.00127f
C1170 a_n2293_46098# a_4419_46090# 0.051687f
C1171 a_1208_46090# a_1138_42852# 0.043831f
C1172 a_10227_46804# a_16020_45572# 3.37e-19
C1173 a_13507_46334# a_15599_45572# 4.46e-20
C1174 a_2063_45854# a_2437_43646# 0.392331f
C1175 a_12861_44030# a_16147_45260# 3.97e-19
C1176 a_n2497_47436# a_n2956_37592# 1.14e-20
C1177 a_376_46348# a_167_45260# 1.16e-21
C1178 a_14543_46987# a_10809_44734# 4.31e-19
C1179 a_n743_46660# a_5907_45546# 0.002962f
C1180 a_13678_32519# a_21973_42336# 3.77e-19
C1181 a_5649_42852# a_22465_38105# 7.91e-21
C1182 a_14401_32519# EN_VIN_BSTR_N 0.772414f
C1183 a_12379_42858# a_12563_42308# 2.54e-20
C1184 a_12089_42308# a_11633_42558# 0.003531f
C1185 a_3353_43940# VDD 0.005542f
C1186 a_22959_43396# a_22775_42308# 2.94e-20
C1187 a_7499_43078# a_10083_42826# 0.375624f
C1188 a_9290_44172# a_8685_42308# 1.4e-21
C1189 a_20193_45348# a_20365_43914# 0.025746f
C1190 a_16922_45042# a_14021_43940# 0.11663f
C1191 a_14673_44172# a_16241_44484# 9.76e-19
C1192 a_17517_44484# a_18204_44850# 6.24e-19
C1193 a_18479_45785# a_15743_43084# 0.001697f
C1194 a_n443_42852# a_n2293_42282# 4.9e-19
C1195 a_8953_45546# a_9377_42558# 0.007183f
C1196 a_11827_44484# a_22223_43948# 0.003019f
C1197 a_21359_45002# a_15493_43940# 8.21e-21
C1198 a_22223_45036# a_11341_43940# 7.11e-20
C1199 a_20202_43084# a_19511_42282# 0.082529f
C1200 a_375_42282# a_n1352_43396# 9.86e-21
C1201 a_13759_47204# VDD 0.004261f
C1202 a_3232_43370# a_3626_43646# 0.204337f
C1203 a_4223_44672# a_n2661_42282# 0.064384f
C1204 a_n356_44636# a_453_43940# 0.02089f
C1205 a_2711_45572# a_18817_42826# 0.001093f
C1206 a_9313_44734# a_20512_43084# 0.028182f
C1207 a_1307_43914# a_n97_42460# 0.23336f
C1208 a_13259_45724# a_13291_42460# 0.089962f
C1209 a_n1925_42282# a_196_42282# 2.11e-19
C1210 a_526_44458# a_n784_42308# 0.011818f
C1211 a_n2293_46634# a_2809_45028# 4.98e-19
C1212 a_5204_45822# a_4880_45572# 0.046074f
C1213 a_765_45546# a_17478_45572# 0.00712f
C1214 a_12005_46116# a_2711_45572# 6.25e-20
C1215 a_n1533_46116# a_n2293_45546# 2.26e-19
C1216 a_768_44030# a_13490_45067# 2.87e-19
C1217 a_3483_46348# a_7499_43078# 0.207714f
C1218 a_11735_46660# a_3357_43084# 5.8e-20
C1219 a_15227_44166# a_20107_45572# 1.29e-19
C1220 a_13059_46348# a_14033_45572# 2.71e-20
C1221 a_10150_46912# a_413_45260# 9.34e-21
C1222 a_5807_45002# a_n2661_43370# 0.018021f
C1223 a_8605_42826# VDD 0.204898f
C1224 a_9223_42460# a_7174_31319# 4.88e-21
C1225 a_5342_30871# C6_P_btm 0.012f
C1226 a_5534_30871# C4_P_btm 8.01e-20
C1227 a_14113_42308# a_15761_42308# 9.35e-19
C1228 a_15051_42282# a_15521_42308# 0.007399f
C1229 a_n4318_37592# a_n4064_38528# 0.020352f
C1230 a_15764_42576# a_16522_42674# 0.05936f
C1231 a_15803_42450# a_16104_42674# 9.73e-19
C1232 a_5111_44636# a_8495_42852# 2.05e-20
C1233 a_13249_42308# a_15051_42282# 4.99e-21
C1234 a_22485_44484# a_14401_32519# 0.01705f
C1235 a_20512_43084# a_20974_43370# 0.020132f
C1236 a_15682_43940# a_17737_43940# 1.13e-19
C1237 a_18114_32519# a_22223_43396# 4.85e-19
C1238 a_11823_42460# a_15890_42674# 1.45e-19
C1239 a_5891_43370# a_9803_43646# 0.011447f
C1240 a_n2017_45002# a_15597_42852# 0.004498f
C1241 a_n1059_45260# a_14853_42852# 0.003368f
C1242 a_n913_45002# a_13622_42852# 4.2e-19
C1243 a_3905_42865# a_5025_43940# 4.14e-19
C1244 a_2521_46116# VDD 0.163553f
C1245 a_18579_44172# a_n97_42460# 0.005302f
C1246 a_14539_43914# a_16409_43396# 0.031761f
C1247 a_375_42282# a_n2293_42282# 5.08e-19
C1248 a_19479_31679# a_22400_42852# 3.1e-20
C1249 a_n2497_47436# a_n2267_43396# 0.222725f
C1250 a_10490_45724# a_11823_42460# 0.022778f
C1251 a_2711_45572# a_14033_45822# 7.91e-19
C1252 a_3090_45724# a_n356_44636# 5.97e-22
C1253 a_12741_44636# a_21359_45002# 4.18e-19
C1254 a_11415_45002# a_22959_45036# 0.001254f
C1255 a_11525_45546# a_11962_45724# 0.095856f
C1256 a_11322_45546# a_12427_45724# 0.010517f
C1257 a_n2293_46634# a_n1899_43946# 5.11e-21
C1258 a_768_44030# a_7845_44172# 0.004571f
C1259 a_18479_47436# a_20623_43914# 0.012705f
C1260 a_11453_44696# a_11750_44172# 1.03e-20
C1261 a_15227_44166# a_18374_44850# 4.22e-19
C1262 a_3483_46348# a_11915_45394# 0.002345f
C1263 a_3699_46348# a_n2661_43370# 5.24e-21
C1264 a_5937_45572# a_5093_45028# 9.15e-20
C1265 a_n2109_47186# a_1983_46706# 9.03e-20
C1266 a_n1741_47186# a_948_46660# 1.63e-20
C1267 a_n971_45724# a_171_46873# 0.002898f
C1268 a_n785_47204# a_n1021_46688# 0.001633f
C1269 a_327_47204# a_n1925_46634# 1.53e-19
C1270 a_n4209_38502# a_n2302_37690# 4.92e-19
C1271 a_n3565_38502# a_n2946_37690# 4.07e-19
C1272 a_2684_37794# a_3754_38470# 5.6e-20
C1273 a_n4064_38528# a_n4334_37440# 1.78e-19
C1274 a_2063_45854# a_n2661_46634# 1.75382f
C1275 a_4915_47217# a_5807_45002# 0.766023f
C1276 a_9313_45822# a_11309_47204# 0.027145f
C1277 a_n1435_47204# a_9804_47204# 1.58e-19
C1278 a_7754_40130# a_7754_39964# 0.301877f
C1279 a_4958_30871# C5_N_btm 1.35e-19
C1280 a_7174_31319# C8_P_btm 7.53e-20
C1281 a_n3420_39072# VDAC_P 2.6e-19
C1282 a_14955_47212# a_n881_46662# 0.008266f
C1283 a_n23_47502# a_n743_46660# 1.99e-20
C1284 a_n237_47217# a_n2438_43548# 0.02231f
C1285 a_n746_45260# a_n133_46660# 0.042075f
C1286 a_21177_47436# a_11453_44696# 3.75e-20
C1287 a_4883_46098# a_22223_47212# 1.16e-19
C1288 a_21811_47423# a_12465_44636# 0.00101f
C1289 a_16104_42674# VDD 0.134357f
C1290 a_15493_43396# a_19095_43396# 1.29e-19
C1291 a_7542_44172# a_7227_42852# 2.27e-20
C1292 a_9313_44734# a_16245_42852# 2.19e-19
C1293 a_13163_45724# VDD 0.322298f
C1294 a_20365_43914# a_20301_43646# 0.001115f
C1295 a_20623_43914# a_4190_30871# 6.24e-20
C1296 a_15493_43940# a_16823_43084# 6.79e-20
C1297 a_19862_44208# a_20556_43646# 0.009839f
C1298 a_10193_42453# DATA[5] 4.15e-19
C1299 a_4905_42826# a_3626_43646# 1.99e-19
C1300 a_3080_42308# a_3539_42460# 0.037567f
C1301 a_1568_43370# a_648_43396# 4.6e-20
C1302 a_n97_42460# a_9396_43370# 1.44e-20
C1303 a_14021_43940# a_15743_43084# 0.045789f
C1304 a_10053_45546# CLK 0.001305f
C1305 a_3422_30871# a_21195_42852# 0.289298f
C1306 a_20269_44172# a_743_42282# 7.1e-21
C1307 a_10809_44734# a_11967_42832# 7.41e-21
C1308 a_n2661_45010# a_n2293_45010# 0.400159f
C1309 a_n2293_46634# a_14358_43442# 0.008808f
C1310 a_3090_45724# a_9165_43940# 0.006052f
C1311 a_8049_45260# a_9159_44484# 1.3e-21
C1312 a_10193_42453# a_16501_45348# 0.009694f
C1313 a_13661_43548# a_14621_43646# 1.53e-19
C1314 a_12549_44172# a_17499_43370# 1.62e-19
C1315 a_4646_46812# a_3539_42460# 1.05e-20
C1316 a_n1151_42308# a_6165_46155# 0.055317f
C1317 a_2063_45854# a_8199_44636# 0.037924f
C1318 a_n1435_47204# a_n901_46420# 4.38e-21
C1319 a_12465_44636# a_22000_46634# 0.001537f
C1320 a_4651_46660# a_5275_47026# 9.73e-19
C1321 a_3877_44458# a_3878_46660# 8.89e-19
C1322 a_2107_46812# a_6086_46660# 2.62e-19
C1323 a_13661_43548# a_17609_46634# 0.002022f
C1324 a_12891_46348# a_12347_46660# 4.22e-19
C1325 a_n443_46116# a_4185_45028# 6.94e-20
C1326 a_4700_47436# a_4704_46090# 1.44e-19
C1327 a_4791_45118# a_4419_46090# 4.81e-19
C1328 C8_N_btm VIN_N 0.907642f
C1329 a_4955_46873# a_5072_46660# 0.17431f
C1330 a_5385_46902# a_5732_46660# 0.051162f
C1331 a_4817_46660# a_6540_46812# 2.48e-19
C1332 VDD DATA[5] 0.504354f
C1333 a_n2661_46634# a_12469_46902# 0.001353f
C1334 a_10227_46804# a_11415_45002# 0.139042f
C1335 C5_N_btm VCM 0.719982f
C1336 C6_N_btm VREF_GND 0.836236f
C1337 a_11453_44696# a_20841_46902# 0.0185f
C1338 a_2747_46873# a_765_45546# 0.040029f
C1339 C7_N_btm VREF 1.818f
C1340 a_n2661_42282# a_5742_30871# 3.56e-20
C1341 a_5649_42852# a_22591_43396# 2.81e-19
C1342 a_14358_43442# a_5342_30871# 2.31e-19
C1343 a_12281_43396# a_12089_42308# 0.210903f
C1344 a_10341_43396# a_13635_43156# 2.32e-19
C1345 a_14579_43548# a_15567_42826# 4.33e-19
C1346 a_15095_43370# a_5534_30871# 1.69e-19
C1347 a_4361_42308# a_17364_32525# 4.28e-20
C1348 a_13678_32519# a_14209_32519# 0.048492f
C1349 a_22223_43396# a_13887_32519# 0.154411f
C1350 a_9290_44172# a_9803_43646# 0.010228f
C1351 a_2711_45572# a_15682_43940# 0.038198f
C1352 a_n2312_39304# a_5932_42308# 4.36e-21
C1353 a_n913_45002# a_5891_43370# 0.255618f
C1354 a_2437_43646# a_n2661_42834# 0.033942f
C1355 a_20202_43084# a_21259_43561# 1.84e-19
C1356 a_3090_45724# a_12379_42858# 0.00513f
C1357 a_1307_43914# a_742_44458# 0.355379f
C1358 a_327_44734# a_n310_44811# 1.25e-19
C1359 a_8016_46348# a_10341_43396# 0.00203f
C1360 a_12861_44030# a_15051_42282# 4e-21
C1361 a_n1925_42282# a_4699_43561# 5.23e-20
C1362 a_526_44458# a_3080_42308# 0.041925f
C1363 a_10775_45002# a_10057_43914# 0.010331f
C1364 a_12741_44636# a_16823_43084# 0.00226f
C1365 a_10227_46804# a_10533_42308# 0.001306f
C1366 a_8953_45002# a_8975_43940# 0.001233f
C1367 a_6945_45028# a_6031_43396# 3.75e-20
C1368 a_6755_46942# a_15682_46116# 0.116442f
C1369 a_6969_46634# a_2324_44458# 7e-22
C1370 a_6151_47436# a_13904_45546# 3.01e-22
C1371 a_n1613_43370# a_1848_45724# 6.13e-21
C1372 a_20107_46660# a_19636_46660# 3.64e-21
C1373 a_19123_46287# a_20719_46660# 8.64e-21
C1374 a_19321_45002# a_19597_46482# 5.66e-19
C1375 a_3090_45724# a_5204_45822# 2.88e-19
C1376 a_15227_44166# a_3483_46348# 0.595533f
C1377 a_17339_46660# a_11415_45002# 0.025523f
C1378 a_n881_46662# a_997_45618# 1.94e-19
C1379 a_3877_44458# a_n1925_42282# 0.034241f
C1380 a_7715_46873# a_6945_45028# 0.001653f
C1381 a_4646_46812# a_526_44458# 0.020719f
C1382 a_n743_46660# a_14180_46482# 0.002131f
C1383 a_13887_32519# a_5934_30871# 2.14e-19
C1384 a_15743_43084# a_15764_42576# 0.006278f
C1385 a_1847_42826# a_1755_42282# 2.18e-19
C1386 a_2075_43172# a_1606_42308# 4.06e-19
C1387 a_5534_30871# a_14097_32519# 0.041746f
C1388 a_4361_42308# a_8325_42308# 0.020707f
C1389 a_17333_42852# a_17749_42852# 0.002387f
C1390 a_18249_42858# a_17665_42852# 3.34e-20
C1391 a_8605_42826# a_n784_42308# 4.32e-21
C1392 a_743_42282# a_9293_42558# 9.79e-19
C1393 a_16664_43396# a_14113_42308# 2.4e-20
C1394 a_n1287_44306# VDD 1.78e-19
C1395 a_3537_45260# a_5829_43940# 3.27e-20
C1396 a_18114_32519# a_20512_43084# 5.22e-19
C1397 a_13259_45724# a_13460_43230# 0.015281f
C1398 a_15415_45028# a_15493_43940# 1.94e-21
C1399 a_13249_42308# a_13749_43396# 3.84e-19
C1400 a_14539_43914# a_16241_44734# 0.006538f
C1401 a_n2293_42834# a_n2661_42282# 0.026231f
C1402 a_n357_42282# a_685_42968# 0.004355f
C1403 a_n443_42852# a_n1423_42826# 1.28e-19
C1404 a_n755_45592# a_421_43172# 1.37e-20
C1405 a_526_44458# a_7309_43172# 0.003264f
C1406 a_9482_43914# a_11173_44260# 0.043729f
C1407 a_13059_46348# a_13575_42558# 3.09e-21
C1408 a_6151_47436# CLK 0.036587f
C1409 a_n863_45724# a_3681_42891# 4.05e-19
C1410 a_10193_42453# a_18783_43370# 0.007846f
C1411 a_7227_47204# DATA[3] 0.357377f
C1412 a_13381_47204# VDD 0.130765f
C1413 a_6109_44484# a_5708_44484# 0.002689f
C1414 a_376_46348# a_n863_45724# 1.69e-21
C1415 SMPL_ON_P a_n2840_44458# 8.99e-19
C1416 a_6755_46942# a_16680_45572# 9.94e-21
C1417 a_n2442_46660# a_n967_45348# 1.82e-19
C1418 a_n2293_46634# en_comp 0.00109f
C1419 a_n1021_46688# a_n913_45002# 2.23e-21
C1420 a_n2312_38680# a_n2810_45028# 0.044149f
C1421 a_15682_46116# a_8049_45260# 0.015666f
C1422 a_n2293_46098# a_1848_45724# 0.006569f
C1423 a_1138_42852# a_n2661_45546# 0.023338f
C1424 a_21588_30879# a_413_45260# 0.041669f
C1425 a_n2497_47436# a_n2267_44484# 0.025633f
C1426 a_n1853_46287# a_n755_45592# 0.021472f
C1427 a_n1641_46494# a_n1099_45572# 0.0023f
C1428 a_n2438_43548# a_n2017_45002# 0.29197f
C1429 a_12861_44030# a_13105_45348# 3.05e-19
C1430 a_18783_43370# VDD 0.289099f
C1431 a_22400_42852# a_13258_32519# 0.039664f
C1432 a_13887_32519# a_11530_34132# 0.005035f
C1433 a_6761_42308# a_8325_42308# 5.55e-19
C1434 a_5934_30871# a_8515_42308# 0.222946f
C1435 a_4190_30871# C4_P_btm 1.36e-19
C1436 a_19279_43940# a_15493_43940# 0.019758f
C1437 a_5343_44458# a_6765_43638# 9.35e-22
C1438 en_comp a_5342_30871# 0.032532f
C1439 a_n913_45002# a_17595_43084# 1.88e-20
C1440 a_n1059_45260# a_17701_42308# 0.073596f
C1441 a_n2017_45002# a_18083_42858# 0.03192f
C1442 a_20980_44850# a_19862_44208# 1.48e-19
C1443 a_4223_44672# a_7112_43396# 3.59e-20
C1444 a_5111_44636# a_9127_43156# 4.76e-19
C1445 a_11691_44458# a_15095_43370# 1.02e-20
C1446 a_22223_45036# a_10341_43396# 2.09e-19
C1447 a_9313_44734# a_21381_43940# 0.028978f
C1448 a_n357_42282# a_14113_42308# 5.29e-20
C1449 a_n2956_38680# a_n3565_38502# 0.302523f
C1450 a_3232_43370# a_8037_42858# 2.1e-22
C1451 a_6298_44484# a_6293_42852# 2.36e-20
C1452 a_12741_44636# a_15415_45028# 1.4e-19
C1453 a_21137_46414# a_21363_45546# 0.001589f
C1454 a_6945_45028# a_20623_45572# 5.77e-19
C1455 a_3483_46348# a_4558_45348# 0.068916f
C1456 a_17715_44484# a_2437_43646# 3.38e-20
C1457 a_8049_45260# a_16680_45572# 0.005473f
C1458 a_11415_45002# a_1307_43914# 0.001965f
C1459 a_4185_45028# a_3537_45260# 1.06643f
C1460 a_15227_44166# a_17719_45144# 0.187414f
C1461 a_19692_46634# a_16922_45042# 0.055961f
C1462 a_n2956_39768# a_n2661_43922# 1.22e-20
C1463 a_n2661_46634# a_n2661_42834# 1.68e-20
C1464 a_2324_44458# a_3357_43084# 0.216574f
C1465 a_9290_44172# a_n913_45002# 0.632534f
C1466 a_5257_43370# a_5883_43914# 0.019234f
C1467 a_2107_46812# a_5891_43370# 1.37e-20
C1468 a_n357_42282# a_7499_43078# 0.259858f
C1469 a_n881_46662# a_11967_42832# 9.73e-21
C1470 a_n3565_39590# a_n3420_37984# 0.031465f
C1471 a_n971_45724# a_4883_46098# 0.031452f
C1472 a_4915_47217# a_14311_47204# 0.001913f
C1473 a_14113_42308# CAL_N 0.001678f
C1474 a_1239_39587# a_1177_38525# 3.88e-21
C1475 a_n4209_39590# a_n4064_37984# 0.032388f
C1476 a_5932_42308# C8_P_btm 1.4e-19
C1477 a_6545_47178# a_n1435_47204# 9.45e-19
C1478 a_6151_47436# a_13717_47436# 0.17202f
C1479 a_1239_39043# a_1736_39043# 0.08488f
C1480 a_n3565_39304# a_n3690_38528# 6.38e-20
C1481 a_n3420_39072# a_n4334_38528# 0.008604f
C1482 a_n3690_39392# a_n3565_38502# 6.38e-20
C1483 a_n2302_39072# a_n2216_39072# 0.011479f
C1484 a_n4064_39616# a_n4209_38216# 0.027937f
C1485 a_n3420_39616# a_n3565_38216# 0.028042f
C1486 a_1221_42558# VDD 2.13e-19
C1487 a_n2288_47178# a_n2312_40392# 0.153632f
C1488 a_n2497_47436# a_n2312_39304# 0.061823f
C1489 a_5934_30871# EN_VIN_BSTR_N 0.073476f
C1490 a_20193_45348# a_22400_42852# 0.05078f
C1491 a_21381_43940# a_20974_43370# 0.02221f
C1492 a_10807_43548# a_9803_43646# 3.09e-19
C1493 a_5883_43914# a_9114_42852# 8.7e-21
C1494 a_1307_43914# a_10533_42308# 1.27e-21
C1495 a_n913_45002# a_21887_42336# 0.060677f
C1496 a_17730_32519# a_13678_32519# 0.054146f
C1497 a_20512_43084# a_13887_32519# 8.15e-19
C1498 a_n356_44636# a_945_42968# 2.2e-19
C1499 a_10949_43914# a_10695_43548# 2.27e-19
C1500 a_20692_30879# EN_OFFSET_CAL 0.004501f
C1501 en_comp a_20107_42308# 4.59e-20
C1502 a_n452_45724# VDD 0.112977f
C1503 a_9313_44734# a_18249_42858# 0.007699f
C1504 a_11415_45002# a_18579_44172# 2.58e-23
C1505 a_16147_45260# a_18787_45572# 4.04e-20
C1506 a_18479_45785# a_17668_45572# 1.16e-19
C1507 a_3877_44458# a_3737_43940# 1.04e-19
C1508 a_6511_45714# a_1423_45028# 4.54e-21
C1509 a_n755_45592# a_n2661_43370# 0.036276f
C1510 a_768_44030# a_1891_43646# 5.62e-19
C1511 a_11823_42460# a_6171_45002# 0.123118f
C1512 a_8199_44636# a_n2661_42834# 0.032396f
C1513 a_8953_45546# a_9159_44484# 0.004058f
C1514 a_526_44458# a_10057_43914# 3.21e-19
C1515 a_10180_45724# a_10775_45002# 0.073185f
C1516 a_10903_43370# a_9313_44734# 0.030402f
C1517 a_2324_44458# a_5826_44734# 9.11e-19
C1518 a_10193_42453# a_8953_45002# 0.001294f
C1519 a_8746_45002# a_8191_45002# 7.28e-19
C1520 a_12741_44636# a_19279_43940# 6.8e-19
C1521 a_n971_45724# a_5649_42852# 7.13e-21
C1522 a_11530_34132# EN_VIN_BSTR_N 1.02927f
C1523 a_n4209_37414# VCM 0.03628f
C1524 a_13717_47436# a_19466_46812# 2.28e-20
C1525 VDAC_N VDD 4.62327f
C1526 a_15811_47375# a_15368_46634# 2.18e-19
C1527 a_n743_46660# a_948_46660# 0.038448f
C1528 a_n2438_43548# a_1123_46634# 0.075317f
C1529 a_n133_46660# a_383_46660# 0.105995f
C1530 a_6886_37412# RST_Z 0.031637f
C1531 a_n3420_37440# VIN_P 0.143165f
C1532 a_6151_47436# a_14035_46660# 6.85e-19
C1533 a_4915_47217# a_14226_46987# 8.89e-19
C1534 a_n3565_37414# VREF 0.046045f
C1535 a_2063_45854# a_765_45546# 1.71006f
C1536 a_n881_46662# a_5257_43370# 0.447042f
C1537 a_n1613_43370# a_7411_46660# 1.61e-20
C1538 a_n2840_46634# a_n2661_46098# 3.35e-19
C1539 a_n1925_46634# a_1983_46706# 0.007111f
C1540 a_171_46873# a_601_46902# 2.33e-20
C1541 a_15507_47210# a_15559_46634# 0.011624f
C1542 a_11599_46634# a_16292_46812# 7.78e-19
C1543 a_10227_46804# a_12251_46660# 0.188053f
C1544 a_15682_43940# a_16877_42852# 2.72e-20
C1545 a_8953_45002# VDD 1.24336f
C1546 a_14358_43442# a_743_42282# 1.97e-20
C1547 a_9145_43396# a_4361_42308# 1.15e-19
C1548 a_10341_43396# a_17678_43396# 2.66e-19
C1549 a_2479_44172# a_2903_42308# 2.23e-20
C1550 a_n4318_39768# a_n1630_35242# 1.81e-19
C1551 a_16409_43396# a_17324_43396# 0.118759f
C1552 a_16243_43396# a_18525_43370# 4.59e-21
C1553 a_9313_44734# a_21125_42558# 2.22e-19
C1554 a_n97_42460# a_13635_43156# 0.001861f
C1555 a_1138_42852# a_1427_43646# 7.47e-20
C1556 a_18175_45572# a_18248_44752# 8.43e-19
C1557 a_4646_46812# a_8605_42826# 9.01e-21
C1558 a_11823_42460# a_14673_44172# 7.39e-20
C1559 a_n755_45592# a_2998_44172# 5.92e-21
C1560 a_6171_45002# a_16321_45348# 3.7e-19
C1561 a_2711_45572# a_20512_43084# 7.39e-20
C1562 a_n2810_45572# a_n3674_39768# 0.023119f
C1563 a_19692_46634# a_15743_43084# 5.26e-19
C1564 a_16327_47482# a_19431_46494# 1.79e-19
C1565 a_n2109_47186# a_6194_45824# 1.26e-19
C1566 a_584_46384# a_n443_42852# 1.36389f
C1567 a_3785_47178# a_3503_45724# 9.09e-22
C1568 a_10467_46802# a_11415_45002# 7.12e-22
C1569 a_n881_46662# a_1337_46116# 0.043447f
C1570 a_4883_46098# a_12005_46436# 1.01e-19
C1571 a_2107_46812# a_9290_44172# 0.091636f
C1572 a_5807_45002# a_10809_44734# 0.065594f
C1573 a_13747_46662# a_6945_45028# 0.035381f
C1574 a_n2293_46634# a_2324_44458# 0.021161f
C1575 a_3877_44458# a_2698_46116# 6.32e-21
C1576 a_13717_47436# a_20205_31679# 2.49e-20
C1577 a_15368_46634# a_13059_46348# 0.101997f
C1578 a_15559_46634# a_15227_46910# 7.75e-19
C1579 a_14976_45028# a_16388_46812# 4.43e-20
C1580 a_n443_46116# a_997_45618# 0.080297f
C1581 a_n743_46660# a_13925_46122# 0.041274f
C1582 a_11599_46634# a_20254_46482# 3.41e-19
C1583 a_10227_46804# a_13259_45724# 0.335001f
C1584 a_13507_46334# a_12638_46436# 0.001374f
C1585 a_4190_30871# a_14097_32519# 0.031855f
C1586 a_3422_30871# C9_P_btm 0.003737f
C1587 a_18249_42858# a_18599_43230# 0.210876f
C1588 a_18083_42858# a_19164_43230# 0.101963f
C1589 a_17333_42852# a_19339_43156# 4.42e-21
C1590 a_3626_43646# a_15803_42450# 0.006237f
C1591 a_2982_43646# a_15890_42674# 9.89e-20
C1592 a_5111_42852# a_4649_42852# 1.58e-19
C1593 a_7765_42852# a_8292_43218# 0.157652f
C1594 a_7229_43940# a_7542_44172# 0.086946f
C1595 a_2382_45260# a_3499_42826# 0.040227f
C1596 a_n443_42852# a_15095_43370# 0.006819f
C1597 a_n357_42282# a_15781_43660# 6.97e-20
C1598 a_n2956_39768# a_n3690_39616# 0.015398f
C1599 a_10193_42453# a_3626_43646# 0.13905f
C1600 a_n2661_44458# a_5891_43370# 0.013115f
C1601 a_3357_43084# a_19862_44208# 9.13e-21
C1602 a_526_44458# a_2075_43172# 0.227071f
C1603 a_n1925_42282# a_1847_42826# 2.13e-20
C1604 a_n2312_38680# a_n2302_40160# 4.94e-19
C1605 a_n2442_46660# a_n4209_39590# 0.095025f
C1606 a_n699_43396# a_n23_44458# 2.43e-20
C1607 a_626_44172# a_n1899_43946# 2.19e-20
C1608 a_n2017_45002# a_12429_44172# 3.24e-21
C1609 a_n913_45002# a_10807_43548# 0.023237f
C1610 a_n1059_45260# a_11750_44172# 1.48e-21
C1611 a_11691_44458# a_11649_44734# 4.78e-19
C1612 a_16763_47508# a_413_45260# 3.7e-19
C1613 a_9625_46129# a_2324_44458# 0.002476f
C1614 a_472_46348# a_1337_46436# 9.76e-19
C1615 a_n743_46660# a_15599_45572# 0.022482f
C1616 a_4915_47217# a_13017_45260# 0.002063f
C1617 a_17339_46660# a_13259_45724# 0.038367f
C1618 a_13507_46334# a_n2017_45002# 5.63e-19
C1619 a_18597_46090# en_comp 3.29e-20
C1620 a_10903_43370# a_12594_46348# 0.169312f
C1621 a_11387_46155# a_13351_46090# 5.76e-21
C1622 a_584_46384# a_375_42282# 0.480677f
C1623 a_3090_45724# a_3503_45724# 0.006081f
C1624 a_16388_46812# a_18051_46116# 3.66e-19
C1625 a_12549_44172# a_18596_45572# 1.55e-20
C1626 a_9313_45822# a_6171_45002# 1.31e-19
C1627 a_2487_47570# a_2437_43646# 0.001086f
C1628 a_15227_44166# a_n357_42282# 0.023198f
C1629 a_6755_46942# a_6598_45938# 2.16e-20
C1630 a_6969_46634# a_6667_45809# 1.42e-19
C1631 a_n971_45724# a_3602_45348# 0.003621f
C1632 a_22223_42860# a_13258_32519# 1.75e-20
C1633 a_564_42282# a_1184_42692# 0.00104f
C1634 a_n3674_37592# a_961_42354# 1.74e-21
C1635 a_12800_43218# a_12563_42308# 5.38e-19
C1636 COMP_P a_n327_42308# 3.18e-21
C1637 a_3626_43646# VDD 0.340378f
C1638 a_11136_42852# a_5742_30871# 6.68e-19
C1639 a_n1630_35242# a_1576_42282# 1.99e-20
C1640 a_21356_42826# a_21335_42336# 0.00235f
C1641 a_n2661_42834# a_8018_44260# 2.37e-19
C1642 a_20447_31679# a_17364_32525# 0.054026f
C1643 en_comp a_743_42282# 1.86e-20
C1644 a_n1059_45260# a_4361_42308# 0.033614f
C1645 a_n913_45002# a_13467_32519# 0.024166f
C1646 a_17970_44736# a_14021_43940# 2.51e-21
C1647 a_6298_44484# a_7499_43940# 3.16e-19
C1648 a_5275_47026# VDD 0.135766f
C1649 a_n2293_42834# a_7112_43396# 6.84e-20
C1650 a_9313_44734# a_14955_43940# 1.56e-20
C1651 a_20512_43084# a_22485_44484# 0.004999f
C1652 a_n357_42282# a_n1329_42308# 7.05e-20
C1653 a_n2956_38216# a_n1630_35242# 4.4e-19
C1654 a_n755_45592# COMP_P 1.75e-21
C1655 a_7499_43078# a_10553_43218# 1.15e-19
C1656 a_14539_43914# a_15037_44260# 8.96e-19
C1657 a_4223_44672# a_9801_43940# 3.24e-20
C1658 a_5883_43914# a_5745_43940# 0.007922f
C1659 a_8049_45260# a_6598_45938# 2.14e-19
C1660 a_5807_45002# a_5883_43914# 0.002403f
C1661 a_n2497_47436# a_n2065_43946# 0.036632f
C1662 a_5937_45572# a_8696_44636# 0.041815f
C1663 a_20202_43084# a_21513_45002# 0.13666f
C1664 a_11415_45002# a_20885_45572# 4.28e-19
C1665 a_22365_46825# a_2437_43646# 0.001459f
C1666 a_526_44458# a_10180_45724# 4e-22
C1667 a_n2661_45546# a_n2956_38216# 0.15505f
C1668 a_n2438_43548# a_n2840_44458# 0.00955f
C1669 a_n2810_45572# a_n2293_45546# 4.68e-19
C1670 a_n1613_43370# a_n2012_44484# 2.46e-19
C1671 a_12549_44172# a_15004_44636# 3.69e-20
C1672 a_768_44030# a_13720_44458# 0.178939f
C1673 a_2324_44458# a_9159_45572# 0.003342f
C1674 a_10809_44734# a_15143_45578# 1.76e-21
C1675 a_10227_46804# a_n2661_43922# 0.041913f
C1676 a_4883_46098# a_9313_44734# 0.015767f
C1677 a_n815_47178# a_n452_47436# 0.107449f
C1678 a_n1605_47204# a_n971_45724# 3.64e-19
C1679 a_n1741_47186# a_n237_47217# 0.083957f
C1680 a_n2109_47186# a_n785_47204# 0.43597f
C1681 SMPL_ON_P a_n746_45260# 9.03e-22
C1682 a_6123_31319# VDAC_Pi 1.96e-19
C1683 a_n784_42308# VDAC_N 0.010209f
C1684 a_1606_42308# a_n4064_37440# 0.002946f
C1685 COMP_P a_22521_40599# 0.204681f
C1686 a_5111_44636# a_1755_42282# 2.47e-19
C1687 a_3065_45002# a_2713_42308# 3.6e-19
C1688 a_2382_45260# a_3318_42354# 0.028613f
C1689 a_n2017_45002# a_7227_42308# 0.005025f
C1690 a_n1059_45260# a_6761_42308# 6.76e-21
C1691 a_n913_45002# a_6773_42558# 0.003807f
C1692 a_9313_44734# a_5649_42852# 0.028023f
C1693 a_11341_43940# a_10651_43940# 7.77e-20
C1694 a_19328_44172# a_19319_43548# 0.033025f
C1695 a_18451_43940# a_18533_43940# 0.171361f
C1696 a_2981_46116# VDD 0.111597f
C1697 a_20193_45348# a_22223_42860# 0.017179f
C1698 a_8975_43940# a_8037_42858# 2.54e-20
C1699 a_18819_46122# a_11827_44484# 1.7e-21
C1700 a_13259_45724# a_1307_43914# 0.023098f
C1701 a_3483_46348# a_9838_44484# 0.014242f
C1702 a_n443_42852# a_n659_45366# 1.08e-19
C1703 a_19900_46494# a_18494_42460# 0.001134f
C1704 a_5164_46348# a_5343_44458# 3.87e-20
C1705 a_3316_45546# a_2382_45260# 0.052075f
C1706 a_2957_45546# a_3065_45002# 4.26e-19
C1707 a_n1151_42308# a_7287_43370# 2.15e-20
C1708 a_3090_45724# a_20679_44626# 5.62e-22
C1709 a_10907_45822# a_12561_45572# 4.22e-21
C1710 a_9290_44172# a_n2661_44458# 0.027487f
C1711 a_17583_46090# a_11691_44458# 3.92e-21
C1712 a_n971_45724# a_8685_43396# 0.079658f
C1713 a_n3420_37984# C4_P_btm 1.42e-19
C1714 a_n4064_37984# C6_P_btm 1.01e-19
C1715 a_n3565_38216# C2_P_btm 0.040789f
C1716 a_n3565_39304# VIN_P 0.039159f
C1717 a_n4209_39304# VREF 0.195875f
C1718 a_12549_44172# a_768_44030# 0.490163f
C1719 a_n443_46116# a_5257_43370# 4.89e-19
C1720 a_n881_46662# a_5807_45002# 0.243322f
C1721 a_2112_39137# VDD 0.284849f
C1722 a_n1741_47186# a_8270_45546# 1.71e-19
C1723 a_n237_47217# a_7832_46660# 0.008175f
C1724 a_n2312_40392# a_n2312_38680# 0.052461f
C1725 a_n2312_39304# a_n2104_46634# 0.018871f
C1726 a_n1435_47204# a_3877_44458# 5.83e-20
C1727 a_2063_45854# a_10623_46897# 0.009821f
C1728 a_n1151_42308# a_8492_46660# 1.89e-20
C1729 a_2982_43646# a_16547_43609# 9.82e-21
C1730 a_3626_43646# a_16137_43396# 0.003078f
C1731 a_8685_43396# a_8229_43396# 1.2e-19
C1732 a_18079_43940# a_18083_42858# 7.22e-20
C1733 a_14539_43914# a_15890_42674# 3.49e-22
C1734 a_8791_43396# a_10341_43396# 1.01e-19
C1735 a_14401_32519# a_22223_43396# 0.006786f
C1736 a_5891_43370# a_8325_42308# 0.053347f
C1737 a_20447_31679# a_21589_35634# 3.86e-20
C1738 a_n97_42460# a_17678_43396# 2.62e-19
C1739 a_17538_32519# a_13678_32519# 0.051187f
C1740 a_20974_43370# a_5649_42852# 0.186094f
C1741 a_n2293_46098# a_5829_43940# 0.05512f
C1742 a_5205_44484# a_7229_43940# 0.006973f
C1743 a_6511_45714# a_6109_44484# 1.17e-19
C1744 a_13507_46334# a_19164_43230# 1.15e-20
C1745 a_n2442_46660# a_n1853_43023# 2.67e-21
C1746 a_768_44030# a_5111_42852# 3.09e-21
C1747 a_3090_45724# a_6765_43638# 0.002105f
C1748 a_16147_45260# a_17023_45118# 0.040001f
C1749 a_18175_45572# a_16922_45042# 5.86e-20
C1750 a_13259_45724# a_18579_44172# 5.71e-20
C1751 a_2324_44458# a_9672_43914# 1.42e-19
C1752 a_8696_44636# a_11691_44458# 0.141053f
C1753 a_3232_43370# a_8191_45002# 0.045343f
C1754 a_6171_45002# a_7705_45326# 0.009164f
C1755 a_6431_45366# a_6709_45028# 0.112564f
C1756 a_526_44458# a_5013_44260# 3.48e-20
C1757 a_11962_45724# a_13076_44458# 1.5e-19
C1758 a_11823_42460# a_12607_44458# 0.01822f
C1759 a_n1613_43370# a_10835_43094# 7.12e-22
C1760 a_11599_46634# a_6945_45028# 0.04727f
C1761 a_2063_45854# a_6347_46155# 2.92e-21
C1762 a_6755_46942# a_11735_46660# 0.61229f
C1763 a_10249_46116# a_11813_46116# 0.001399f
C1764 a_n743_46660# a_16655_46660# 0.004413f
C1765 a_n881_46662# a_3699_46348# 0.203393f
C1766 a_n1613_43370# a_4185_45028# 1.83e-19
C1767 a_16327_47482# a_19335_46494# 0.155998f
C1768 a_14311_47204# a_10809_44734# 3.31e-20
C1769 a_n1741_47186# a_12638_46436# 0.016323f
C1770 a_n443_46116# a_1337_46116# 0.002343f
C1771 a_20916_46384# a_12741_44636# 0.023496f
C1772 a_21588_30879# a_20820_30879# 0.084472f
C1773 a_12465_44636# a_10903_43370# 0.003556f
C1774 a_4883_46098# a_12594_46348# 0.022174f
C1775 a_13507_46334# a_13759_46122# 0.004601f
C1776 a_10227_46804# a_18189_46348# 2.07e-20
C1777 a_11453_44696# a_9290_44172# 0.064153f
C1778 a_5111_42852# a_5755_42852# 1.15e-19
C1779 a_13467_32519# a_20922_43172# 5.27e-19
C1780 a_21487_43396# a_21195_42852# 0.01192f
C1781 a_4361_42308# a_19987_42826# 1.33e-19
C1782 a_15095_43370# a_14635_42282# 0.001265f
C1783 a_20269_44172# a_13258_32519# 1.75e-21
C1784 a_20623_43914# a_19511_42282# 1.33e-21
C1785 a_15493_43940# a_19332_42282# 2.75e-21
C1786 a_4235_43370# a_1755_42282# 6.88e-21
C1787 a_n1557_42282# a_1184_42692# 1.23e-19
C1788 a_5649_42852# a_18599_43230# 9.69e-21
C1789 a_17767_44458# VDD 0.348803f
C1790 a_19862_44208# a_20107_42308# 2.1e-21
C1791 a_10334_44484# CLK 0.012484f
C1792 a_9145_43396# a_13622_42852# 5.7e-20
C1793 a_1823_45246# a_3935_42891# 0.002482f
C1794 a_n443_42852# a_n1177_43370# 1.95e-19
C1795 a_1307_43914# a_n2661_43922# 0.023892f
C1796 a_14976_45348# a_14539_43914# 4.77e-20
C1797 a_15037_45618# a_14955_43940# 3.52e-21
C1798 a_n2312_40392# a_7174_31319# 6.67e-21
C1799 a_2711_45572# a_21381_43940# 4.03e-21
C1800 a_9482_43914# a_15463_44811# 0.005265f
C1801 a_413_45260# a_19279_43940# 1.83e-21
C1802 a_2324_44458# a_743_42282# 8.04e-21
C1803 a_20447_31679# a_19237_31679# 0.051563f
C1804 a_n755_45592# a_1568_43370# 7.31e-20
C1805 a_3090_45724# a_12800_43218# 0.002125f
C1806 w_1575_34946# a_n1532_35090# 0.796778f
C1807 a_12891_46348# a_11962_45724# 0.001251f
C1808 a_12549_44172# a_11652_45724# 6.46e-20
C1809 a_17339_46660# a_18189_46348# 0.170772f
C1810 a_8270_45546# a_10586_45546# 3.82e-21
C1811 a_765_45546# a_17715_44484# 0.117636f
C1812 a_472_46348# a_1823_45246# 0.001742f
C1813 a_n2497_47436# a_n2810_45028# 9.88e-21
C1814 a_3699_46634# a_3503_45724# 6.06e-21
C1815 a_n2661_46634# a_3775_45552# 1.47e-21
C1816 a_768_44030# a_11525_45546# 1.76e-21
C1817 a_11735_46660# a_8049_45260# 8.52e-20
C1818 a_n2293_46098# a_4185_45028# 0.06423f
C1819 a_1208_46090# a_1176_45822# 0.141891f
C1820 a_805_46414# a_1138_42852# 2.41e-19
C1821 a_n881_46662# a_15143_45578# 0.069805f
C1822 a_4883_46098# a_15037_45618# 7.22e-21
C1823 a_10227_46804# a_17478_45572# 8.9e-22
C1824 a_584_46384# a_2437_43646# 0.302508f
C1825 a_14226_46987# a_10809_44734# 4.26e-19
C1826 a_n743_46660# a_5263_45724# 7.27e-19
C1827 a_13678_32519# a_22465_38105# 0.034429f
C1828 a_14401_32519# a_11530_34132# 0.004736f
C1829 a_n2293_42282# a_4921_42308# 2.29e-20
C1830 a_3052_44056# VDD 0.001151f
C1831 a_3080_42308# VDAC_N 0.007198f
C1832 a_14209_32519# a_22775_42308# 1.21e-19
C1833 a_12089_42308# a_11551_42558# 0.109508f
C1834 a_9049_44484# a_9127_43156# 1.35e-22
C1835 a_7499_43078# a_8952_43230# 0.054554f
C1836 a_9290_44172# a_8325_42308# 1.58e-20
C1837 a_20193_45348# a_20269_44172# 0.002705f
C1838 a_18479_45785# a_18783_43370# 2.61e-19
C1839 a_10037_47542# DATA[4] 1.79e-19
C1840 a_8199_44636# a_9885_42558# 0.009365f
C1841 a_8953_45546# a_9293_42558# 0.007436f
C1842 a_11827_44484# a_11341_43940# 0.231114f
C1843 a_13675_47204# VDD 0.004094f
C1844 a_3232_43370# a_3540_43646# 0.00217f
C1845 a_2711_45572# a_18249_42858# 0.001642f
C1846 a_n2661_44458# a_10807_43548# 1.72e-19
C1847 a_n356_44636# a_1414_42308# 0.179164f
C1848 a_n1925_42282# a_n473_42460# 1.12e-19
C1849 a_5937_45572# a_7227_45028# 0.064518f
C1850 a_5204_45822# a_4808_45572# 7.79e-20
C1851 a_5257_43370# a_3537_45260# 0.001934f
C1852 a_17339_46660# a_17478_45572# 2.92e-22
C1853 a_765_45546# a_15861_45028# 0.004302f
C1854 a_11901_46660# a_2437_43646# 9.19e-20
C1855 a_2324_44458# a_2277_45546# 8.22e-19
C1856 a_10903_43370# a_2711_45572# 0.213719f
C1857 a_3483_46348# a_8568_45546# 0.137016f
C1858 a_19466_46812# a_19418_45938# 2.93e-19
C1859 a_9863_46634# a_413_45260# 1.44e-20
C1860 a_n1151_42308# a_n23_44458# 0.101137f
C1861 a_2107_46812# a_2304_45348# 9.3e-21
C1862 a_1606_42308# a_n3420_39072# 0.001872f
C1863 a_8037_42858# VDD 0.344922f
C1864 a_8791_42308# a_7174_31319# 9.76e-21
C1865 a_5342_30871# C7_P_btm 5.39e-19
C1866 a_5534_30871# C5_P_btm 8.45e-20
C1867 a_14113_42308# a_15521_42308# 0.002088f
C1868 a_15764_42576# a_16104_42674# 0.029366f
C1869 a_1307_43914# a_3445_43172# 1.01e-21
C1870 a_13249_42308# a_14113_42308# 2.26e-19
C1871 a_20512_43084# a_14401_32519# 5.21e-19
C1872 a_11823_42460# a_15959_42545# 9.34e-20
C1873 a_5891_43370# a_9145_43396# 0.049186f
C1874 a_9313_44734# a_8685_43396# 0.124273f
C1875 a_n356_44636# a_12281_43396# 2.72e-19
C1876 a_10193_42453# a_13921_42308# 0.002387f
C1877 a_n1059_45260# a_13622_42852# 1.72e-19
C1878 a_167_45260# VDD 1.41955f
C1879 a_14539_43914# a_16547_43609# 0.01221f
C1880 a_16979_44734# a_16243_43396# 3.15e-20
C1881 a_19721_31679# a_13678_32519# 0.051384f
C1882 a_n2661_43922# a_9396_43370# 9.06e-21
C1883 a_2998_44172# a_5326_44056# 9.84e-20
C1884 a_n2497_47436# a_n2129_43609# 0.216536f
C1885 a_10490_45724# a_12427_45724# 0.108721f
C1886 a_8746_45002# a_11823_42460# 2.13e-21
C1887 a_7499_43078# a_13249_42308# 1.99e-20
C1888 a_2711_45572# a_12016_45572# 2.58e-19
C1889 a_12741_44636# a_21101_45002# 7.11e-19
C1890 a_12465_44636# a_14955_43940# 6.55e-20
C1891 a_10809_44734# a_13017_45260# 1.77e-20
C1892 a_11322_45546# a_11962_45724# 0.270736f
C1893 a_11525_45546# a_11652_45724# 0.138143f
C1894 a_n443_42852# a_8696_44636# 8.12e-20
C1895 a_n1925_42282# a_5111_44636# 5.66e-21
C1896 a_n2293_46634# a_n1761_44111# 4.77e-21
C1897 a_11415_45002# a_22223_45036# 0.011148f
C1898 a_768_44030# a_7542_44172# 0.005732f
C1899 a_18597_46090# a_19862_44208# 0.536021f
C1900 a_15227_44166# a_18443_44721# 0.002052f
C1901 a_3483_46348# a_n2661_43370# 0.953959f
C1902 a_5937_45572# a_5009_45028# 6.92e-20
C1903 a_n4315_30879# a_n1532_35090# 2.87e-19
C1904 a_n2109_47186# a_2107_46812# 0.032545f
C1905 a_n1741_47186# a_1123_46634# 9.86e-20
C1906 a_n785_47204# a_n1925_46634# 2.12e-19
C1907 a_n3565_38502# a_n3420_37440# 0.034147f
C1908 a_n4209_38502# a_n4064_37440# 0.028279f
C1909 a_n4064_38528# a_n4209_37414# 0.027936f
C1910 a_n3420_38528# a_n3565_37414# 0.029229f
C1911 a_584_46384# a_n2661_46634# 0.034039f
C1912 a_11031_47542# a_11309_47204# 0.110775f
C1913 a_9313_45822# a_11117_47542# 6.66e-19
C1914 a_n1435_47204# a_8128_46384# 9.08e-20
C1915 a_4958_30871# C4_N_btm 1.18e-19
C1916 a_7174_31319# C9_P_btm 9.33e-20
C1917 a_n746_45260# a_n2438_43548# 0.031949f
C1918 a_n237_47217# a_n743_46660# 0.192378f
C1919 a_n971_45724# a_n133_46660# 0.011188f
C1920 a_20990_47178# a_11453_44696# 1.3e-19
C1921 a_4883_46098# a_12465_44636# 0.024607f
C1922 a_14311_47204# a_n881_46662# 0.037789f
C1923 a_3754_39964# VDAC_Pi 0.296508f
C1924 a_9049_44484# CLK 7.29e-22
C1925 a_n2661_42282# a_n13_43084# 5.65e-21
C1926 a_20269_44172# a_20301_43646# 4.32e-19
C1927 a_20365_43914# a_4190_30871# 1.62e-20
C1928 a_19862_44208# a_743_42282# 4.04e-19
C1929 a_12791_45546# VDD 0.205486f
C1930 a_4699_43561# a_3539_42460# 0.109444f
C1931 a_3080_42308# a_3626_43646# 0.092602f
C1932 a_1049_43396# a_648_43396# 5.57e-19
C1933 a_1209_43370# a_1512_43396# 0.001377f
C1934 a_1568_43370# a_548_43396# 1.89e-20
C1935 a_n97_42460# a_8791_43396# 6.57e-22
C1936 a_14021_43940# a_18783_43370# 0.006778f
C1937 a_11823_42460# RST_Z 1.21e-19
C1938 a_n2956_37592# a_n2302_37984# 0.005102f
C1939 a_3422_30871# a_21356_42826# 0.024863f
C1940 a_22612_30879# a_10341_43396# 1.26e-21
C1941 a_16020_45572# a_16019_45002# 6.19e-19
C1942 a_15861_45028# a_16751_45260# 0.044248f
C1943 a_3483_46348# a_2998_44172# 2.54e-20
C1944 a_n2661_45010# a_n2472_45002# 0.065751f
C1945 a_n2840_45002# a_n2293_45010# 2.81e-19
C1946 a_19479_31679# en_comp 1.32e-19
C1947 a_n2293_46634# a_14579_43548# 0.035629f
C1948 a_8034_45724# a_n2661_43922# 6.46e-21
C1949 a_13507_46334# a_14209_32519# 0.008866f
C1950 a_10193_42453# a_16405_45348# 0.001843f
C1951 a_13661_43548# a_14537_43646# 1.89e-19
C1952 a_12549_44172# a_16759_43396# 1.5e-19
C1953 a_4646_46812# a_3626_43646# 4.2e-20
C1954 a_n755_45592# a_5883_43914# 1.16e-19
C1955 a_n743_46660# a_8270_45546# 0.274248f
C1956 a_n1151_42308# a_5497_46414# 0.089064f
C1957 a_n1435_47204# a_n1641_46494# 2.5e-20
C1958 a_12465_44636# a_21188_46660# 3.64e-21
C1959 a_4651_46660# a_5072_46660# 0.083408f
C1960 a_4646_46812# a_5275_47026# 8.49e-19
C1961 a_3877_44458# a_3633_46660# 2.14e-19
C1962 a_2107_46812# a_5841_46660# 1.55e-19
C1963 a_n1925_46634# a_8601_46660# 6.89e-21
C1964 a_5807_45002# a_17609_46634# 2.45e-19
C1965 a_13747_46662# a_15559_46634# 1.73e-20
C1966 a_12891_46348# a_12978_47026# 1.98e-19
C1967 a_4915_47217# a_3483_46348# 1.09e-19
C1968 a_4791_45118# a_4185_45028# 0.064362f
C1969 C7_N_btm VIN_N 1.52449f
C1970 a_18479_47436# a_20885_46660# 6.01e-19
C1971 a_4817_46660# a_5732_46660# 0.118759f
C1972 a_n2661_46634# a_11901_46660# 0.030789f
C1973 C5_N_btm VREF_GND 0.676559f
C1974 C4_N_btm VCM 0.716447f
C1975 a_10227_46804# a_20202_43084# 0.022898f
C1976 a_11453_44696# a_20273_46660# 0.545219f
C1977 VDD DATA[4] 0.326957f
C1978 C6_N_btm VREF 1.41944f
C1979 a_5649_42852# a_13887_32519# 0.004879f
C1980 a_4361_42308# a_22959_43396# 1.39e-19
C1981 a_14579_43548# a_5342_30871# 0.041574f
C1982 a_12281_43396# a_12379_42858# 0.036584f
C1983 a_14205_43396# a_5534_30871# 1.04e-19
C1984 a_15095_43370# a_14543_43071# 1.43e-19
C1985 a_21855_43396# a_14209_32519# 2.74e-19
C1986 a_13467_32519# a_17364_32525# 0.050014f
C1987 a_9290_44172# a_9145_43396# 0.103991f
C1988 a_6171_45002# a_14539_43914# 3.43e-19
C1989 a_n2312_40392# a_5932_42308# 6.05e-21
C1990 a_n1059_45260# a_5891_43370# 0.186322f
C1991 a_3090_45724# a_10341_42308# 0.002812f
C1992 a_8016_46348# a_9885_43646# 0.001881f
C1993 a_12861_44030# a_14113_42308# 1.46e-20
C1994 a_3357_43084# a_5708_44484# 0.005179f
C1995 a_327_44734# a_n23_44458# 0.141544f
C1996 a_8953_45002# a_10057_43914# 0.001204f
C1997 a_526_44458# a_4699_43561# 1.19e-19
C1998 a_n1925_42282# a_4235_43370# 0.199349f
C1999 a_3877_44458# a_526_44458# 0.017621f
C2000 a_6755_46942# a_2324_44458# 0.155169f
C2001 a_4915_47217# a_14495_45572# 0.001776f
C2002 a_6151_47436# a_13527_45546# 4.69e-21
C2003 a_19551_46910# a_19636_46660# 1.48e-19
C2004 a_7411_46660# a_6945_45028# 0.004283f
C2005 a_5807_45002# a_19443_46116# 0.003665f
C2006 a_13747_46662# a_20009_46494# 9.03e-20
C2007 a_3090_45724# a_5164_46348# 1.94e-19
C2008 a_11459_47204# a_10193_42453# 3.13e-19
C2009 a_9313_45822# a_8746_45002# 5.46e-20
C2010 a_4883_46098# a_2711_45572# 0.041245f
C2011 a_768_44030# a_n2661_45546# 0.07332f
C2012 a_4791_45118# a_6229_45572# 1.28e-19
C2013 a_n1613_43370# a_997_45618# 1.47e-20
C2014 a_n881_46662# a_n755_45592# 0.077214f
C2015 a_15743_43084# a_15486_42560# 6.65e-19
C2016 a_1847_42826# a_1606_42308# 0.025123f
C2017 a_5649_42852# a_8515_42308# 5.44e-20
C2018 a_18083_42858# a_17749_42852# 3.87e-19
C2019 a_17333_42852# a_17665_42852# 0.001922f
C2020 a_8037_42858# a_n784_42308# 6.19e-21
C2021 a_743_42282# a_9803_42558# 0.010183f
C2022 a_n1453_44318# VDD 3.29e-19
C2023 a_3537_45260# a_5745_43940# 1.23e-19
C2024 a_n1059_45260# a_18533_43940# 5.26e-21
C2025 a_2711_45572# a_5649_42852# 1.3e-19
C2026 a_13259_45724# a_13635_43156# 0.017822f
C2027 a_14539_43914# a_14673_44172# 0.205935f
C2028 a_16112_44458# a_16241_44734# 0.062574f
C2029 a_n755_45592# a_133_43172# 0.002433f
C2030 a_n443_42852# a_n1991_42858# 1.6e-19
C2031 a_n357_42282# a_421_43172# 2.38e-19
C2032 a_526_44458# a_6101_43172# 6.27e-21
C2033 a_9482_43914# a_10555_44260# 0.088693f
C2034 a_n863_45724# a_2905_42968# 0.269475f
C2035 a_10193_42453# a_18525_43370# 2.7e-19
C2036 a_18479_45785# a_3626_43646# 4.26e-20
C2037 a_6851_47204# DATA[3] 0.146601f
C2038 a_11459_47204# VDD 0.34771f
C2039 a_n998_44484# a_n2661_43922# 3.71e-19
C2040 a_6109_44484# a_5608_44484# 4.33e-19
C2041 a_5826_44734# a_5708_44484# 1.98e-20
C2042 a_11189_46129# a_12638_46436# 1.22e-19
C2043 a_n2293_46098# a_997_45618# 0.003758f
C2044 a_n1076_46494# a_n863_45724# 1.04e-19
C2045 a_n901_46420# a_n452_45724# 0.004896f
C2046 a_6755_46942# a_16855_45546# 3.44e-19
C2047 a_15227_44166# a_13249_42308# 2.89e-20
C2048 a_n2442_46660# en_comp 0.02478f
C2049 a_n2293_46634# a_n2956_37592# 4.76e-19
C2050 a_n1021_46688# a_n1059_45260# 3.15e-21
C2051 a_n1925_46634# a_n913_45002# 1.36e-21
C2052 a_2324_44458# a_8049_45260# 0.054166f
C2053 a_20916_46384# a_413_45260# 6.71e-20
C2054 a_1176_45822# a_n2661_45546# 0.004027f
C2055 a_5807_45002# a_3537_45260# 0.005102f
C2056 a_n2956_38680# a_n1925_42282# 4.34e-20
C2057 a_n2497_47436# a_n2129_44697# 0.019202f
C2058 a_768_44030# a_5205_44484# 0.033081f
C2059 a_9804_47204# a_8953_45002# 0.003283f
C2060 a_n2438_43548# a_n2109_45247# 0.007532f
C2061 a_18525_43370# VDD 0.263553f
C2062 a_5379_42460# a_5742_30871# 7.37e-20
C2063 a_4190_30871# C5_P_btm 1.71e-19
C2064 a_7963_42308# a_8515_42308# 8.26e-20
C2065 a_n2956_39304# a_n3565_38502# 0.001812f
C2066 a_20820_30879# a_22469_39537# 7.31e-20
C2067 a_5343_44458# a_6197_43396# 1.12e-20
C2068 a_n913_45002# a_16795_42852# 7.33e-21
C2069 a_n1059_45260# a_17595_43084# 0.049f
C2070 a_n2017_45002# a_17701_42308# 0.132871f
C2071 a_10057_43914# a_3626_43646# 2.08e-20
C2072 a_4223_44672# a_7287_43370# 2.11e-19
C2073 a_2127_44172# a_2537_44260# 0.007617f
C2074 a_21076_30879# a_22521_39511# 6.56e-20
C2075 a_5111_44636# a_8387_43230# 0.001241f
C2076 a_11827_44484# a_10341_43396# 3.05e-19
C2077 a_7542_44172# a_7845_44172# 0.137004f
C2078 a_6298_44484# a_6031_43396# 0.001377f
C2079 a_7715_46873# a_6298_44484# 3.13e-20
C2080 a_12741_44636# a_14797_45144# 1.29e-20
C2081 a_20075_46420# a_20528_45572# 5.63e-19
C2082 a_6165_46155# a_413_45260# 9.78e-21
C2083 a_11813_46116# a_11691_44458# 1.05e-21
C2084 a_6945_45028# a_20841_45814# 4.67e-19
C2085 a_17583_46090# a_2437_43646# 9.89e-22
C2086 a_13507_46334# a_17730_32519# 1.98e-20
C2087 a_8049_45260# a_16855_45546# 0.004398f
C2088 a_11415_45002# a_16019_45002# 0.007819f
C2089 a_3699_46348# a_3537_45260# 3.5e-21
C2090 a_19466_46812# a_16922_45042# 0.030378f
C2091 a_3483_46348# a_4574_45260# 0.022358f
C2092 a_15227_44166# a_17613_45144# 0.048772f
C2093 a_n2956_39768# a_n2661_42834# 7.06e-20
C2094 a_12549_44172# a_17517_44484# 0.019389f
C2095 a_14840_46494# a_3357_43084# 2.67e-21
C2096 a_9290_44172# a_n1059_45260# 0.092471f
C2097 a_3090_45724# a_18494_42460# 1.58e-20
C2098 a_4185_45028# a_3429_45260# 0.004974f
C2099 COMP_P VIN_N 0.001768f
C2100 a_n4209_39304# a_n3420_38528# 0.029412f
C2101 a_1606_42308# C10_N_btm 1.34e-19
C2102 a_5932_42308# C9_P_btm 9.33e-20
C2103 a_2063_45854# a_10227_46804# 0.186188f
C2104 a_6151_47436# a_n1435_47204# 0.061966f
C2105 a_6575_47204# a_9067_47204# 0.210614f
C2106 a_4915_47217# a_13487_47204# 0.013601f
C2107 a_n3565_39304# a_n3565_38502# 0.041674f
C2108 a_n3420_39072# a_n4209_38502# 0.032647f
C2109 a_n4064_39072# a_n2216_39072# 0.005565f
C2110 a_n3420_39616# a_n4334_38304# 4.87e-19
C2111 a_n4064_40160# a_n3607_38304# 5.58e-20
C2112 a_1149_42558# VDD 4.29e-19
C2113 a_4958_30871# a_8530_39574# 1.39e-19
C2114 a_5934_30871# a_11530_34132# 8.66e-19
C2115 a_n2833_47464# a_n2312_39304# 0.009425f
C2116 a_n2497_47436# a_n2312_40392# 0.194574f
C2117 a_20193_45348# a_20836_43172# 9.63e-20
C2118 a_14021_43940# a_3626_43646# 1.24e-20
C2119 a_21381_43940# a_14401_32519# 4.91e-20
C2120 a_10807_43548# a_9145_43396# 0.290878f
C2121 a_n2293_43922# a_12895_43230# 0.001356f
C2122 a_3422_30871# a_20749_43396# 1.42e-19
C2123 a_19237_31679# a_13467_32519# 0.052472f
C2124 a_n1761_44111# a_743_42282# 1.3e-19
C2125 a_20512_43084# a_22223_43396# 0.001484f
C2126 a_n356_44636# a_873_42968# 2.03e-19
C2127 a_n2293_42834# a_5379_42460# 1.97e-21
C2128 a_10729_43914# a_10695_43548# 0.00999f
C2129 a_20205_31679# EN_OFFSET_CAL 0.002855f
C2130 en_comp a_13258_32519# 0.007613f
C2131 a_n863_45724# VDD 1.89058f
C2132 a_n913_45002# a_21335_42336# 0.062808f
C2133 a_9313_44734# a_17333_42852# 0.010555f
C2134 a_18175_45572# a_17668_45572# 1.93e-20
C2135 a_18691_45572# a_18799_45938# 0.057222f
C2136 a_18479_45785# a_17568_45572# 5.46e-20
C2137 a_6472_45840# a_1423_45028# 3.3e-21
C2138 a_n2293_46634# a_n2267_43396# 7.31e-22
C2139 a_n357_42282# a_n2661_43370# 0.034578f
C2140 a_7499_43078# a_11787_45002# 4.1e-20
C2141 a_12427_45724# a_6171_45002# 8.61e-21
C2142 a_11823_42460# a_3232_43370# 0.002063f
C2143 a_8016_46348# a_n2661_43922# 0.02895f
C2144 a_5937_45572# a_9159_44484# 0.040512f
C2145 a_12465_44636# a_8685_43396# 5.48e-20
C2146 a_10227_46804# a_14955_43396# 0.035123f
C2147 a_2324_44458# a_5289_44734# 0.001168f
C2148 a_10180_45724# a_8953_45002# 0.107499f
C2149 a_12861_44030# a_15781_43660# 0.025765f
C2150 a_5066_45546# a_5343_44458# 1.18e-21
C2151 a_n1613_43370# a_5257_43370# 0.025984f
C2152 a_n4209_37414# VREF_GND 0.00198f
C2153 a_6886_37412# VDD 0.235486f
C2154 a_n743_46660# a_1123_46634# 0.054493f
C2155 a_n2438_43548# a_383_46660# 0.0336f
C2156 a_n133_46660# a_601_46902# 0.053479f
C2157 a_6151_47436# a_13885_46660# 0.001762f
C2158 a_4915_47217# a_14513_46634# 2.71e-19
C2159 a_12861_44030# a_15227_44166# 0.810382f
C2160 a_13717_47436# a_19333_46634# 1.58e-20
C2161 a_584_46384# a_765_45546# 0.086068f
C2162 a_n881_46662# a_5429_46660# 3.91e-20
C2163 a_5700_37509# RST_Z 0.051902f
C2164 a_n1925_46634# a_2107_46812# 1.12874f
C2165 a_171_46873# a_33_46660# 0.207108f
C2166 a_15811_47375# a_14976_45028# 2.33e-19
C2167 a_11599_46634# a_15559_46634# 0.028826f
C2168 a_10227_46804# a_12469_46902# 0.181535f
C2169 a_3905_42865# a_1755_42282# 5.4e-20
C2170 a_n3674_39768# a_n3674_37592# 0.024722f
C2171 a_15682_43940# a_16245_42852# 6.93e-20
C2172 a_8191_45002# VDD 0.39677f
C2173 a_3539_42460# a_1847_42826# 1.09e-20
C2174 a_14579_43548# a_743_42282# 3.98e-19
C2175 a_10341_43396# a_17433_43396# 1.6e-19
C2176 a_16409_43396# a_17499_43370# 0.042737f
C2177 a_16977_43638# a_16759_43396# 0.209641f
C2178 a_16243_43396# a_18429_43548# 6.92e-21
C2179 a_16137_43396# a_18525_43370# 2.8e-19
C2180 a_16547_43609# a_17324_43396# 5.47e-21
C2181 a_n97_42460# a_12895_43230# 1.91e-20
C2182 a_2982_43646# a_3681_42891# 0.006879f
C2183 a_1138_42852# a_n1557_42282# 0.009215f
C2184 a_18175_45572# a_17970_44736# 2.35e-20
C2185 a_21542_45572# a_19721_31679# 3.76e-20
C2186 a_4646_46812# a_8037_42858# 0.001539f
C2187 en_comp a_20193_45348# 6.75e-20
C2188 a_n2956_39768# a_n2293_42282# 5.23e-20
C2189 a_11787_45002# a_11915_45394# 0.004764f
C2190 a_11963_45334# a_n2661_43370# 2.8e-19
C2191 a_1307_43914# a_5837_45028# 1.79e-20
C2192 a_6171_45002# a_14309_45028# 0.00276f
C2193 a_n357_42282# a_2998_44172# 4.93e-20
C2194 a_n2810_45572# a_n4318_39768# 0.023737f
C2195 a_19692_46634# a_18783_43370# 1.14e-20
C2196 a_16327_47482# a_19240_46482# 2.52e-19
C2197 a_n2109_47186# a_5907_45546# 8.91e-19
C2198 a_n1151_42308# a_n356_45724# 4.29e-20
C2199 a_1431_47204# a_1609_45822# 9.46e-22
C2200 a_584_46384# a_509_45822# 3.94e-19
C2201 a_4955_46873# a_1823_45246# 0.001178f
C2202 a_5257_43370# a_n2293_46098# 0.049293f
C2203 a_n881_46662# a_835_46155# 2.99e-19
C2204 a_11901_46660# a_765_45546# 0.007273f
C2205 a_4883_46098# a_10037_46155# 4.58e-19
C2206 a_19321_45002# a_19900_46494# 0.002634f
C2207 a_20916_46384# a_18985_46122# 5.23e-20
C2208 a_2107_46812# a_10355_46116# 7.69e-19
C2209 a_13661_43548# a_6945_45028# 0.015293f
C2210 a_12156_46660# a_12347_46660# 4.61e-19
C2211 a_15368_46634# a_15227_46910# 0.050747f
C2212 a_n443_46116# a_n755_45592# 0.651643f
C2213 a_3090_45724# a_16388_46812# 1.08e-19
C2214 a_14976_45028# a_13059_46348# 0.209989f
C2215 a_n743_46660# a_13759_46122# 0.01783f
C2216 a_11599_46634# a_20009_46494# 2.17e-19
C2217 a_17591_47464# a_13259_45724# 3.28e-20
C2218 a_10227_46804# a_14383_46116# 0.01306f
C2219 a_13507_46334# a_12379_46436# 0.001281f
C2220 a_3422_30871# C10_P_btm 0.002966f
C2221 a_21381_43940# a_21421_42336# 1.07e-19
C2222 a_18249_42858# a_18817_42826# 0.16939f
C2223 a_18083_42858# a_19339_43156# 0.042271f
C2224 a_17333_42852# a_18599_43230# 3.68e-19
C2225 a_8685_43396# a_8515_42308# 5.84e-21
C2226 a_3626_43646# a_15764_42576# 0.002707f
C2227 a_2982_43646# a_15959_42545# 2.23e-19
C2228 a_7765_42852# a_7573_43172# 1.97e-19
C2229 a_4520_42826# a_4649_42852# 0.062574f
C2230 a_7871_42858# a_8292_43218# 0.086377f
C2231 a_1307_43914# a_n809_44244# 5.87e-21
C2232 a_7229_43940# a_7281_43914# 0.164835f
C2233 a_n443_42852# a_14205_43396# 0.118229f
C2234 a_n357_42282# a_15681_43442# 3.86e-20
C2235 a_n2956_39768# a_n3565_39590# 0.302561f
C2236 a_n2661_44458# a_8375_44464# 0.003111f
C2237 a_11827_44484# a_n2293_43922# 0.028646f
C2238 a_526_44458# a_1847_42826# 0.154735f
C2239 a_n2312_38680# a_n4064_40160# 8.3e-19
C2240 a_n2442_46660# a_n2216_40160# 0.001258f
C2241 a_n699_43396# a_n356_44636# 0.044884f
C2242 a_626_44172# a_n1761_44111# 3.66e-23
C2243 a_n913_45002# a_10949_43914# 0.001202f
C2244 a_n2017_45002# a_11750_44172# 1.48e-22
C2245 a_n1059_45260# a_10807_43548# 0.031771f
C2246 a_16023_47582# a_413_45260# 1.6e-19
C2247 a_8953_45546# a_2324_44458# 0.047906f
C2248 a_5257_43370# a_7230_45938# 6.16e-21
C2249 a_3483_46348# a_10809_44734# 0.02965f
C2250 a_n2293_46098# a_1337_46116# 0.002811f
C2251 a_3090_45724# a_3316_45546# 0.04556f
C2252 a_n2661_46634# a_8696_44636# 2.14e-19
C2253 a_5807_45002# a_16842_45938# 1.8e-19
C2254 a_9313_45822# a_3232_43370# 1.83e-20
C2255 a_2266_47570# a_2437_43646# 0.001239f
C2256 a_2063_45854# a_1307_43914# 0.005774f
C2257 a_6755_46942# a_6667_45809# 1.38e-20
C2258 a_6969_46634# a_6511_45714# 7.16e-20
C2259 a_n2109_47186# a_6125_45348# 3.53e-19
C2260 a_n971_45724# a_3495_45348# 0.005013f
C2261 a_10903_43370# a_12005_46116# 0.277468f
C2262 SMPL_ON_N a_20447_31679# 0.029368f
C2263 a_22165_42308# a_13258_32519# 0.004531f
C2264 a_n3674_37592# a_1184_42692# 1.16e-19
C2265 a_n1630_35242# a_1067_42314# 4.97e-19
C2266 a_3540_43646# VDD 0.209044f
C2267 a_11136_42852# a_11323_42473# 8.95e-19
C2268 a_2982_43646# RST_Z 0.015013f
C2269 a_n2661_42834# a_7911_44260# 4.06e-19
C2270 a_22315_44484# a_19237_31679# 4.46e-20
C2271 a_n2017_45002# a_4361_42308# 0.004087f
C2272 a_6298_44484# a_6671_43940# 4.34e-19
C2273 a_5072_46660# VDD 0.081835f
C2274 a_n2293_42834# a_7287_43370# 7.97e-19
C2275 a_9313_44734# a_13483_43940# 1.18e-20
C2276 a_n863_45724# a_n784_42308# 0.358682f
C2277 a_n357_42282# COMP_P 3.45e-20
C2278 a_14539_43914# a_14761_44260# 3.61e-19
C2279 a_11827_44484# a_n97_42460# 4.56e-20
C2280 a_1307_43914# a_14955_43396# 5.43e-20
C2281 a_8049_45260# a_6667_45809# 2.79e-19
C2282 a_n2661_45546# a_n2472_45546# 0.040937f
C2283 a_15368_46634# a_9482_43914# 3.52e-20
C2284 a_8199_44636# a_8696_44636# 0.265919f
C2285 a_11415_45002# a_20719_45572# 7.75e-19
C2286 a_5066_45546# a_4880_45572# 0.04794f
C2287 a_10903_43370# a_14033_45822# 0.040019f
C2288 a_n2840_45546# a_n2293_45546# 2.81e-19
C2289 a_n2810_45572# a_n2956_38216# 6.20057f
C2290 a_14976_45028# a_13556_45296# 0.003018f
C2291 a_12549_44172# a_13720_44458# 7.87e-20
C2292 a_768_44030# a_13076_44458# 0.132449f
C2293 a_n2293_46634# a_n2267_44484# 2.41e-19
C2294 a_10227_46804# a_n2661_42834# 0.024624f
C2295 a_n1605_47204# a_n452_47436# 3.88e-21
C2296 SMPL_ON_P a_n971_45724# 2.75e-21
C2297 a_n1741_47186# a_n746_45260# 0.032595f
C2298 a_n2109_47186# a_n23_47502# 0.043455f
C2299 a_n2288_47178# a_n785_47204# 6.98e-20
C2300 a_22400_42852# a_22705_38406# 2.84e-20
C2301 a_5934_30871# a_7754_40130# 0.007046f
C2302 a_22775_42308# a_22465_38105# 0.330766f
C2303 a_21613_42308# a_21973_42336# 0.001645f
C2304 a_7309_42852# VDD 0.177437f
C2305 a_n1630_35242# a_3726_37500# 0.001279f
C2306 a_6123_31319# a_7754_39964# 5.24e-20
C2307 COMP_P CAL_N 0.008927f
C2308 a_5111_44636# a_1606_42308# 1.35e-20
C2309 a_2382_45260# a_2903_42308# 1.98e-20
C2310 a_n2017_45002# a_6761_42308# 0.006728f
C2311 a_20692_30879# VDAC_N 4.47e-19
C2312 a_9313_44734# a_13678_32519# 0.097255f
C2313 a_n913_45002# a_6481_42558# 0.005099f
C2314 a_n2661_42282# a_104_43370# 5.48e-21
C2315 a_18326_43940# a_18533_43940# 0.001502f
C2316 a_19328_44172# a_19808_44306# 0.001696f
C2317 a_18451_43940# a_19319_43548# 1.99e-20
C2318 a_20193_45348# a_22165_42308# 0.252856f
C2319 a_13259_45724# a_16019_45002# 1.86e-19
C2320 a_3483_46348# a_5883_43914# 5.92e-19
C2321 a_13507_46334# a_17538_32519# 8.21e-20
C2322 a_20708_46348# a_19778_44110# 4.6e-21
C2323 a_19900_46494# a_18184_42460# 4.45e-21
C2324 a_20075_46420# a_18494_42460# 2.66e-19
C2325 a_5068_46348# a_5343_44458# 1.11e-21
C2326 a_3218_45724# a_2382_45260# 5.5e-20
C2327 a_2957_45546# a_2680_45002# 4.36e-19
C2328 a_3316_45546# a_2274_45254# 8.04e-21
C2329 a_2107_46812# a_10949_43914# 8.95e-21
C2330 a_6511_45714# a_3357_43084# 1.21e-20
C2331 a_15227_44166# a_17325_44484# 0.001944f
C2332 a_n443_42852# a_n967_45348# 3.13e-19
C2333 a_n755_45592# a_3537_45260# 0.025346f
C2334 a_15682_46116# a_11691_44458# 1.87e-21
C2335 a_n3420_37984# C5_P_btm 1.22e-19
C2336 a_n3565_38216# C3_P_btm 0.001023f
C2337 a_n4064_37984# C7_P_btm 4.26e-20
C2338 a_n3420_37440# VDAC_P 4.18e-19
C2339 VDAC_Pi a_n923_35174# 0.001372f
C2340 a_12891_46348# a_768_44030# 0.193145f
C2341 a_4791_45118# a_5257_43370# 0.36404f
C2342 a_n1613_43370# a_5807_45002# 0.086053f
C2343 a_n2216_39072# VDD 0.00419f
C2344 a_n971_45724# a_8035_47026# 8.58e-19
C2345 a_n2312_39304# a_n2293_46634# 0.021162f
C2346 a_2063_45854# a_10467_46802# 0.036614f
C2347 a_n1151_42308# a_8667_46634# 1.5e-19
C2348 a_2982_43646# a_16243_43396# 7.65e-20
C2349 a_8685_43396# a_7466_43396# 3.33e-20
C2350 a_14539_43914# a_15959_42545# 3.47e-21
C2351 a_n356_44636# a_11551_42558# 1.46e-19
C2352 a_19721_31679# a_22775_42308# 3.9e-21
C2353 a_10555_44260# a_10796_42968# 6.32e-21
C2354 a_15493_43396# a_15567_42826# 4.1e-20
C2355 a_5891_43370# a_8337_42558# 4.22e-21
C2356 a_20447_31679# a_19864_35138# 1.11e-20
C2357 a_17973_43940# a_18083_42858# 5.46e-19
C2358 a_n97_42460# a_17433_43396# 1.55e-19
C2359 a_20974_43370# a_13678_32519# 0.020999f
C2360 a_14401_32519# a_5649_42852# 3.64e-19
C2361 a_3090_45724# a_6197_43396# 0.010809f
C2362 a_n2293_46098# a_5745_43940# 0.019006f
C2363 a_11823_42460# a_8975_43940# 7.95e-20
C2364 a_526_44458# a_5244_44056# 4.69e-21
C2365 a_n1925_42282# a_3905_42865# 0.023709f
C2366 a_n967_45348# a_375_42282# 0.001506f
C2367 a_6472_45840# a_6109_44484# 7.09e-20
C2368 a_13507_46334# a_19339_43156# 4.77e-21
C2369 a_16147_45260# a_16922_45042# 0.016249f
C2370 a_13259_45724# a_18245_44484# 1.46e-19
C2371 a_2324_44458# a_9028_43914# 4.61e-20
C2372 a_16115_45572# a_16237_45028# 4.93e-20
C2373 a_3232_43370# a_7705_45326# 0.02181f
C2374 a_6171_45002# a_6709_45028# 0.021915f
C2375 a_6431_45366# a_7229_43940# 1.72e-19
C2376 a_10193_42453# a_16979_44734# 0.016398f
C2377 a_12427_45724# a_12607_44458# 3.74e-21
C2378 a_n2956_39768# a_n1423_42826# 3.32e-21
C2379 a_n2442_46660# a_n2157_42858# 5.35e-21
C2380 a_4883_46098# a_12005_46116# 0.012933f
C2381 a_13507_46334# a_13351_46090# 0.214666f
C2382 a_14955_47212# a_6945_45028# 0.013254f
C2383 a_2063_45854# a_8034_45724# 0.034258f
C2384 a_10249_46116# a_11735_46660# 7.95e-19
C2385 a_6755_46942# a_11186_47026# 0.014167f
C2386 a_n743_46660# a_16434_46660# 6.95e-19
C2387 a_n881_46662# a_3483_46348# 0.5947f
C2388 a_n1613_43370# a_3699_46348# 2.1e-19
C2389 a_16327_47482# a_19553_46090# 0.172776f
C2390 a_n1741_47186# a_12379_46436# 0.067348f
C2391 a_5807_45002# a_n2293_46098# 2.61e-20
C2392 a_20916_46384# a_20820_30879# 4.91e-20
C2393 a_10227_46804# a_17715_44484# 1.63e-20
C2394 a_13487_47204# a_10809_44734# 1.49e-19
C2395 a_22612_30879# a_11415_45002# 1.26e-21
C2396 a_21588_30879# a_22591_46660# 5.88e-20
C2397 a_6151_47436# a_526_44458# 3.76e-20
C2398 a_12281_43396# a_12800_43218# 9.09e-21
C2399 a_16979_44734# VDD 0.256327f
C2400 a_13467_32519# a_19987_42826# 5.32e-19
C2401 a_4361_42308# a_19164_43230# 1.97e-20
C2402 a_15095_43370# a_13291_42460# 6.1e-21
C2403 a_14205_43396# a_14635_42282# 6.79e-20
C2404 a_4093_43548# a_1755_42282# 1.31e-21
C2405 a_5649_42852# a_18817_42826# 1.52e-20
C2406 a_19862_44208# a_13258_32519# 3.59e-19
C2407 a_1568_43370# a_2351_42308# 3.07e-21
C2408 a_10157_44484# CLK 0.002339f
C2409 a_1823_45246# a_3681_42891# 2.81e-20
C2410 a_12741_44636# a_12089_42308# 6.17e-22
C2411 a_n2956_38216# a_n1557_42282# 1.25e-20
C2412 a_1307_43914# a_n2661_42834# 3.43601f
C2413 a_2711_45572# a_19741_43940# 0.005487f
C2414 a_n863_45724# a_3080_42308# 0.001926f
C2415 a_1423_45028# a_3363_44484# 8.49e-19
C2416 a_13556_45296# a_15433_44458# 0.1084f
C2417 a_9482_43914# a_15146_44811# 0.006879f
C2418 a_n2293_42834# a_n23_44458# 8.19e-21
C2419 a_n913_45002# a_3422_30871# 0.145467f
C2420 a_13507_46334# a_22465_38105# 9.82e-20
C2421 a_n755_45592# a_1049_43396# 8.22e-21
C2422 a_n357_42282# a_1568_43370# 0.036942f
C2423 a_n2293_46634# a_9223_42460# 1.9e-20
C2424 w_1575_34946# a_n1386_35608# 0.005843f
C2425 a_n1925_46634# a_5907_45546# 6.84e-21
C2426 a_8270_45546# a_8379_46155# 8.95e-21
C2427 a_17339_46660# a_17715_44484# 0.018672f
C2428 a_765_45546# a_17583_46090# 0.067337f
C2429 a_376_46348# a_1823_45246# 9.94e-21
C2430 SMPL_ON_P a_n2293_45010# 4.92e-20
C2431 a_n2661_46634# a_7227_45028# 3.38e-20
C2432 a_768_44030# a_11322_45546# 6.14e-20
C2433 a_12549_44172# a_11525_45546# 7.96e-19
C2434 a_n2293_46098# a_3699_46348# 3.53e-20
C2435 a_472_46348# a_1138_42852# 0.028956f
C2436 a_805_46414# a_1176_45822# 0.024739f
C2437 a_10227_46804# a_15861_45028# 0.002162f
C2438 a_17591_47464# a_17478_45572# 1.31e-20
C2439 a_2124_47436# a_2437_43646# 0.025048f
C2440 a_n881_46662# a_14495_45572# 0.170589f
C2441 a_3090_45724# a_5066_45546# 1.9e-19
C2442 a_14513_46634# a_10809_44734# 0.002278f
C2443 a_n743_46660# a_4099_45572# 1.05e-19
C2444 a_13678_32519# a_22397_42558# 0.001628f
C2445 a_10341_42308# a_11633_42558# 2.57e-19
C2446 a_2455_43940# VDD 0.144352f
C2447 a_3080_42308# a_6886_37412# 6.84e-19
C2448 a_14209_32519# a_21613_42308# 9.39e-21
C2449 a_12089_42308# a_5742_30871# 1.26e-19
C2450 a_22591_43396# a_22775_42308# 1.54e-19
C2451 a_7499_43078# a_9127_43156# 0.08498f
C2452 a_5111_44636# a_3539_42460# 2.98e-20
C2453 a_17061_44734# a_17517_44484# 0.004238f
C2454 a_9804_47204# DATA[4] 0.015379f
C2455 a_8953_45546# a_9803_42558# 0.031932f
C2456 a_8199_44636# a_9377_42558# 0.001018f
C2457 a_4185_45028# a_14456_42282# 1.64e-19
C2458 a_21359_45002# a_11341_43940# 1.28e-20
C2459 a_11827_44484# a_21115_43940# 0.005833f
C2460 a_20193_45348# a_19862_44208# 0.041264f
C2461 a_13569_47204# VDD 0.00491f
C2462 a_3232_43370# a_2982_43646# 0.416054f
C2463 a_n2661_44458# a_10949_43914# 1.28e-19
C2464 a_n356_44636# a_1467_44172# 0.061333f
C2465 a_13259_45724# a_13814_43218# 5.53e-19
C2466 a_n1925_42282# a_n961_42308# 2.27e-19
C2467 a_2711_45572# a_17333_42852# 2.07e-20
C2468 a_2107_46812# a_2232_45348# 1.12e-19
C2469 a_8199_44636# a_7227_45028# 3.82e-20
C2470 a_5937_45572# a_6598_45938# 2.01e-19
C2471 a_5204_45822# a_5024_45822# 1.6e-19
C2472 a_5732_46660# a_6171_45002# 1.44e-19
C2473 a_4646_46812# a_8191_45002# 7.69e-21
C2474 a_765_45546# a_8696_44636# 0.001141f
C2475 a_17339_46660# a_15861_45028# 5.36e-22
C2476 a_11813_46116# a_2437_43646# 7.51e-20
C2477 a_13507_46334# a_19721_31679# 8.21e-20
C2478 a_11387_46155# a_2711_45572# 4.02e-20
C2479 a_8049_45260# a_12839_46116# 0.004724f
C2480 a_12891_46348# a_13490_45067# 0.00125f
C2481 a_584_46384# a_700_44734# 5.41e-19
C2482 a_3483_46348# a_8162_45546# 0.009853f
C2483 a_9313_45822# a_8975_43940# 3.56e-20
C2484 a_n1151_42308# a_n356_44636# 0.093166f
C2485 a_7765_42852# VDD 0.333322f
C2486 a_8685_42308# a_7174_31319# 4.88e-21
C2487 a_n3674_38216# a_n4064_38528# 0.020875f
C2488 a_5342_30871# C8_P_btm 0.093874f
C2489 a_5534_30871# C6_P_btm 0.01116f
C2490 a_n4318_37592# a_n3420_38528# 0.024768f
C2491 a_14113_42308# a_17124_42282# 4.43e-19
C2492 a_1307_43914# a_n2293_42282# 0.004191f
C2493 a_13249_42308# a_13657_42558# 0.002219f
C2494 a_20512_43084# a_21381_43940# 0.019564f
C2495 a_11823_42460# a_15803_42450# 8.2e-20
C2496 a_5891_43370# a_8423_43396# 7.18e-21
C2497 a_10193_42453# a_13657_42308# 5.7e-19
C2498 a_16979_44734# a_16137_43396# 8.54e-22
C2499 a_14539_43914# a_16243_43396# 0.029808f
C2500 a_16112_44458# a_16547_43609# 1.97e-19
C2501 a_18114_32519# a_13678_32519# 0.055126f
C2502 a_n2661_43922# a_8791_43396# 3e-20
C2503 a_n2661_42834# a_9396_43370# 8.6e-21
C2504 a_2202_46116# VDD 0.20904f
C2505 a_2998_44172# a_5025_43940# 5.5e-20
C2506 a_3600_43914# a_3992_43940# 0.016359f
C2507 a_11453_44696# a_10949_43914# 7.02e-20
C2508 a_n2497_47436# a_n2433_43396# 0.173242f
C2509 a_17715_44484# a_1307_43914# 3.38e-21
C2510 a_10490_45724# a_11962_45724# 0.114064f
C2511 a_10193_42453# a_11823_42460# 0.235429f
C2512 a_2711_45572# a_11778_45572# 8.22e-19
C2513 a_12741_44636# a_21005_45260# 0.001247f
C2514 a_12465_44636# a_13483_43940# 3.64e-19
C2515 a_10809_44734# a_11963_45334# 4.58e-19
C2516 a_11322_45546# a_11652_45724# 0.26844f
C2517 a_526_44458# a_5111_44636# 0.338508f
C2518 a_n1925_42282# a_5147_45002# 9.69e-37
C2519 a_8270_45546# a_5891_43370# 0.052984f
C2520 a_n2293_46634# a_n2065_43946# 2.74e-19
C2521 a_11415_45002# a_11827_44484# 0.169126f
C2522 a_768_44030# a_7281_43914# 0.006034f
C2523 a_n1613_43370# a_n822_43940# 2.39e-19
C2524 a_16327_47482# a_15493_43940# 0.04211f
C2525 a_15227_44166# a_18287_44626# 5.33e-20
C2526 a_3483_46348# a_11361_45348# 5.71e-19
C2527 a_3147_46376# a_n2661_43370# 9.13e-21
C2528 a_7227_45028# a_8192_45572# 7.21e-20
C2529 a_n4315_30879# a_n1386_35608# 1.11e-19
C2530 a_n2109_47186# a_948_46660# 5.02e-20
C2531 a_n1741_47186# a_383_46660# 4.76e-20
C2532 a_n23_47502# a_n1925_46634# 4.04e-20
C2533 a_13507_46334# a_22223_47212# 0.001502f
C2534 a_21496_47436# a_12465_44636# 2.84e-19
C2535 a_4883_46098# a_21811_47423# 0.054014f
C2536 a_7174_31319# C10_P_btm 1.34e-19
C2537 a_n3565_38502# a_n3690_37440# 4.13e-19
C2538 a_n4209_38502# a_n2946_37690# 3.29e-19
C2539 a_n3420_38528# a_n4334_37440# 1.39e-19
C2540 a_2684_37794# VDAC_Ni 0.004723f
C2541 a_2124_47436# a_n2661_46634# 1.6e-20
C2542 a_4791_45118# a_5807_45002# 0.129041f
C2543 a_6151_47436# a_13759_47204# 0.00136f
C2544 a_11031_47542# a_11117_47542# 0.006584f
C2545 a_9313_45822# a_10037_47542# 0.00168f
C2546 a_13487_47204# a_n881_46662# 0.108977f
C2547 a_4958_30871# C3_N_btm 1.05e-19
C2548 a_n3565_39304# VDAC_P 4.47e-19
C2549 a_n746_45260# a_n743_46660# 0.068305f
C2550 a_n971_45724# a_n2438_43548# 0.038673f
C2551 a_20894_47436# a_11453_44696# 7.99e-20
C2552 a_7499_43078# CLK 9.27e-21
C2553 a_n2661_42282# a_n1076_43230# 2.25e-20
C2554 a_9313_44734# a_15597_42852# 4.48e-19
C2555 a_n2810_45028# a_n2302_37984# 0.003394f
C2556 a_20269_44172# a_4190_30871# 4.64e-20
C2557 a_11341_43940# a_16823_43084# 2.12e-19
C2558 a_15493_43396# a_20556_43646# 1.31e-20
C2559 a_11823_42460# VDD 4.44574f
C2560 a_4235_43370# a_3539_42460# 0.005553f
C2561 a_4699_43561# a_3626_43646# 5.64e-20
C2562 a_4905_42826# a_2982_43646# 1.34e-19
C2563 a_n97_42460# a_8147_43396# 8.39e-22
C2564 a_14021_43940# a_18525_43370# 0.007346f
C2565 a_19478_44306# a_743_42282# 1.05e-20
C2566 a_n2956_37592# a_n4064_37984# 0.012393f
C2567 a_3422_30871# a_20922_43172# 0.045027f
C2568 a_21398_44850# a_21356_42826# 1.64e-20
C2569 a_8696_44636# a_16751_45260# 0.265287f
C2570 a_15861_45028# a_1307_43914# 0.067929f
C2571 a_n2840_45002# a_n2472_45002# 7.52e-19
C2572 a_n2293_46634# a_13667_43396# 0.011502f
C2573 SMPL_ON_N a_13467_32519# 0.029246f
C2574 a_8034_45724# a_n2661_42834# 5.76e-21
C2575 a_10193_42453# a_16321_45348# 9.06e-20
C2576 a_12549_44172# a_16977_43638# 3.73e-20
C2577 a_1823_45246# a_5663_43940# 5.36e-19
C2578 a_17715_44484# a_18579_44172# 2.18e-19
C2579 a_13507_46334# a_22591_43396# 0.011335f
C2580 a_3877_44458# a_3626_43646# 1.07e-19
C2581 a_n357_42282# a_5883_43914# 1.93e-19
C2582 a_n1151_42308# a_5204_45822# 0.487224f
C2583 a_2063_45854# a_8016_46348# 8.48e-19
C2584 a_n1435_47204# a_n1423_46090# 2.49e-19
C2585 a_12465_44636# a_21363_46634# 5.44e-20
C2586 a_16327_47482# a_12741_44636# 0.074082f
C2587 a_4651_46660# a_6540_46812# 7.72e-21
C2588 a_4646_46812# a_5072_46660# 0.013764f
C2589 a_13661_43548# a_15559_46634# 8.86e-22
C2590 a_13747_46662# a_15368_46634# 0.110984f
C2591 a_5807_45002# a_16292_46812# 0.202526f
C2592 a_n443_46116# a_3483_46348# 0.009289f
C2593 a_n881_46662# a_14513_46634# 0.017832f
C2594 C6_N_btm VIN_N 0.391905f
C2595 a_4883_46098# a_22000_46634# 0.004514f
C2596 a_18479_47436# a_20719_46660# 8e-19
C2597 a_5385_46902# a_5167_46660# 0.209641f
C2598 a_4817_46660# a_5907_46634# 0.042415f
C2599 a_n1741_47186# a_13351_46090# 7.57e-20
C2600 a_13507_46334# a_20731_47026# 8.28e-19
C2601 C4_N_btm VREF_GND 0.671882f
C2602 C3_N_btm VCM 0.716273f
C2603 a_10227_46804# a_22365_46825# 2.64e-20
C2604 VDD DATA[3] 0.309692f
C2605 a_11453_44696# a_20411_46873# 0.020751f
C2606 C5_N_btm VREF 0.987144f
C2607 a_19321_45002# a_3090_45724# 0.163821f
C2608 a_n2661_46634# a_11813_46116# 0.162517f
C2609 a_5649_42852# a_22223_43396# 0.165664f
C2610 a_13678_32519# a_13887_32519# 10.751599f
C2611 a_4361_42308# a_14209_32519# 8.23e-20
C2612 a_12281_43396# a_10341_42308# 2.53e-20
C2613 a_14358_43442# a_5534_30871# 0.002889f
C2614 a_14205_43396# a_14543_43071# 9.94e-20
C2615 a_15095_43370# a_13460_43230# 5.97e-21
C2616 a_14579_43548# a_15279_43071# 0.108607f
C2617 a_768_44030# a_564_42282# 4.13e-22
C2618 a_6171_45002# a_16112_44458# 5.94e-20
C2619 a_2711_45572# a_13483_43940# 1.84e-21
C2620 a_19431_45546# a_17517_44484# 1.08e-20
C2621 a_n2017_45002# a_5891_43370# 0.065487f
C2622 a_3090_45724# a_10922_42852# 0.002693f
C2623 a_4646_46812# a_7309_42852# 1.16e-20
C2624 a_4883_46098# a_5934_30871# 0.005052f
C2625 a_327_44734# a_n356_44636# 0.085841f
C2626 a_14403_45348# a_14309_45028# 1.26e-19
C2627 a_8953_45002# a_10440_44484# 1.69e-19
C2628 a_n1925_42282# a_4093_43548# 0.018682f
C2629 a_526_44458# a_4235_43370# 0.032501f
C2630 w_1575_34946# a_2113_38308# 6.01e-20
C2631 a_n743_46660# a_12379_46436# 1.32e-19
C2632 a_6755_46942# a_14840_46494# 0.021842f
C2633 a_8270_45546# a_9290_44172# 0.433963f
C2634 a_4915_47217# a_13249_42308# 0.161597f
C2635 a_6151_47436# a_13163_45724# 1.73e-21
C2636 a_21188_46660# a_22000_46634# 2.08e-19
C2637 a_20623_46660# a_20731_47026# 0.057222f
C2638 a_19123_46287# a_19636_46660# 1.03e-19
C2639 a_5257_43370# a_6945_45028# 6.65e-21
C2640 a_2107_46812# a_10044_46482# 2.82e-19
C2641 a_2063_45854# a_11682_45822# 3.96e-19
C2642 a_n1613_43370# a_n755_45592# 0.052236f
C2643 a_n881_46662# a_n357_42282# 7.4e-19
C2644 a_15743_43084# a_15051_42282# 5.67e-19
C2645 a_n1644_44306# VDD 0.082968f
C2646 a_5649_42852# a_5934_30871# 0.058776f
C2647 a_13887_32519# a_6123_31319# 1.56e-19
C2648 a_4361_42308# a_4169_42308# 7.22e-19
C2649 a_17333_42852# a_16877_42852# 0.003649f
C2650 a_17701_42308# a_17749_42852# 0.004244f
C2651 a_18083_42858# a_17665_42852# 2.63e-19
C2652 a_743_42282# a_9223_42460# 0.010592f
C2653 a_n863_45724# a_2075_43172# 2.8e-19
C2654 a_13259_45724# a_12895_43230# 6.21e-19
C2655 a_15415_45028# a_11341_43940# 7.47e-21
C2656 a_14537_43396# a_15493_43940# 8.79e-19
C2657 a_16112_44458# a_14673_44172# 0.077293f
C2658 a_6151_47436# DATA[5] 0.19492f
C2659 a_n443_42852# a_n1853_43023# 0.141267f
C2660 a_n357_42282# a_133_43172# 0.001058f
C2661 a_9482_43914# a_9895_44260# 0.005015f
C2662 a_10193_42453# a_18429_43548# 0.002926f
C2663 a_11823_42460# a_16137_43396# 6.91e-20
C2664 a_6491_46660# DATA[3] 0.011549f
C2665 a_9313_45822# VDD 0.5747f
C2666 a_n998_44484# a_n2661_42834# 2.81e-19
C2667 a_n1243_44484# a_n2661_43922# 2.55e-19
C2668 a_5147_45002# a_3737_43940# 2.51e-20
C2669 a_11189_46129# a_12379_46436# 1.91e-20
C2670 a_n2293_46098# a_n755_45592# 0.086057f
C2671 a_n901_46420# a_n863_45724# 0.00998f
C2672 a_n1991_46122# a_n1099_45572# 5.38e-19
C2673 a_6755_46942# a_16115_45572# 0.004389f
C2674 a_765_45546# a_7227_45028# 2.27e-20
C2675 a_n2442_46660# a_n2956_37592# 0.049818f
C2676 a_14840_46494# a_8049_45260# 0.002948f
C2677 a_n2497_47436# a_n2433_44484# 0.027254f
C2678 a_1208_46090# a_n2661_45546# 4.43e-20
C2679 a_n2293_46634# a_n2810_45028# 0.004774f
C2680 a_n2956_39304# a_n1925_42282# 5.53e-20
C2681 a_n1076_46494# a_n1079_45724# 8.64e-19
C2682 a_376_46348# a_n2293_45546# 1.03e-21
C2683 a_n2438_43548# a_n2293_45010# 0.033143f
C2684 a_7963_42308# a_5934_30871# 0.002785f
C2685 a_6123_31319# a_8515_42308# 8.12e-20
C2686 a_18429_43548# VDD 0.163446f
C2687 a_5267_42460# a_5742_30871# 1.46e-20
C2688 a_20256_43172# a_20107_42308# 1.36e-19
C2689 a_22400_42852# a_19511_42282# 2.86e-21
C2690 a_1606_42308# a_15051_42282# 1.09e-19
C2691 a_4190_30871# C6_P_btm 0.005085f
C2692 a_13678_32519# EN_VIN_BSTR_N 0.031779f
C2693 a_n2956_38680# a_n4209_38502# 0.235751f
C2694 a_20835_44721# a_15493_43940# 7.97e-20
C2695 a_19279_43940# a_11341_43940# 0.003029f
C2696 a_18579_44172# a_20623_43914# 1.89e-20
C2697 a_5343_44458# a_6293_42852# 1.91e-20
C2698 a_20820_30879# a_22821_38993# 1.52e-19
C2699 a_n1059_45260# a_16795_42852# 0.182174f
C2700 a_n2017_45002# a_17595_43084# 0.016123f
C2701 a_11823_42460# a_n784_42308# 5.93e-20
C2702 a_n2661_42834# a_10867_43940# 6.15e-20
C2703 a_4223_44672# a_6547_43396# 3.73e-19
C2704 a_2127_44172# a_2253_44260# 0.013015f
C2705 en_comp a_5534_30871# 0.021896f
C2706 a_21359_45002# a_10341_43396# 7.35e-21
C2707 a_375_42282# a_n1853_43023# 2.99e-20
C2708 a_1414_42308# a_3499_42826# 0.023314f
C2709 a_12741_44636# a_14537_43396# 0.094691f
C2710 a_21137_46414# a_20841_45814# 2.76e-19
C2711 a_20708_46348# a_20623_45572# 9.36e-19
C2712 a_6945_45028# a_20273_45572# 2.17e-19
C2713 a_15682_46116# a_2437_43646# 4.97e-20
C2714 a_8049_45260# a_16115_45572# 0.004258f
C2715 a_11415_45002# a_15595_45028# 0.003773f
C2716 a_3483_46348# a_3537_45260# 0.605469f
C2717 a_13661_43548# a_15463_44811# 1.29e-19
C2718 a_1823_45246# a_3232_43370# 0.344002f
C2719 a_3090_45724# a_18184_42460# 2.47e-20
C2720 a_9290_44172# a_n2017_45002# 0.089856f
C2721 a_15227_44166# a_17023_45118# 2.94e-19
C2722 a_4185_45028# a_3065_45002# 0.060303f
C2723 a_15015_46420# a_3357_43084# 6.88e-21
C2724 a_3699_46348# a_3429_45260# 7.23e-21
C2725 a_5932_42308# C10_P_btm 1.34e-19
C2726 a_n3565_39590# a_n3565_38216# 0.031123f
C2727 a_6123_31319# EN_VIN_BSTR_N 0.050716f
C2728 a_n4209_39590# a_n3420_37984# 0.032713f
C2729 a_1606_42308# C9_N_btm 9.33e-20
C2730 a_5815_47464# a_n1435_47204# 0.001005f
C2731 a_4915_47217# a_12861_44030# 0.025257f
C2732 a_6151_47436# a_13381_47204# 0.014822f
C2733 a_n4064_39072# a_n2860_39072# 0.003765f
C2734 a_n3420_39616# a_n4209_38216# 0.027924f
C2735 a_n4064_40160# a_n4251_38304# 0.001069f
C2736 a_961_42354# VDD 0.091526f
C2737 a_n2833_47464# a_n2312_40392# 0.064992f
C2738 a_4958_30871# a_7754_38470# 9.47e-20
C2739 a_20193_45348# a_20573_43172# 1.16e-20
C2740 a_n2661_45546# CLK_DATA 1.81e-19
C2741 a_3422_30871# a_17364_32525# 0.007014f
C2742 a_n1079_45724# VDD 0.172275f
C2743 a_n2293_42834# a_5267_42460# 5.73e-21
C2744 a_22485_44484# a_13678_32519# 3.76e-22
C2745 a_20512_43084# a_5649_42852# 0.141324f
C2746 a_9313_44734# a_18083_42858# 0.05022f
C2747 a_n913_45002# a_7174_31319# 0.02792f
C2748 en_comp a_19647_42308# 4.59e-20
C2749 a_10405_44172# a_10695_43548# 1.89e-19
C2750 a_n2312_38680# a_n4318_39304# 0.023234f
C2751 a_8270_45546# a_10807_43548# 9.25e-21
C2752 a_19431_45546# a_19256_45572# 0.233657f
C2753 a_18909_45814# a_18799_45938# 0.097745f
C2754 a_16147_45260# a_17668_45572# 5.57e-19
C2755 a_18691_45572# a_18596_45572# 0.049827f
C2756 a_n2293_46634# a_n2129_43609# 4.29e-21
C2757 a_7499_43078# a_10951_45334# 0.008335f
C2758 a_768_44030# a_n1557_42282# 1.25e-19
C2759 a_11962_45724# a_6171_45002# 8.2e-19
C2760 a_13259_45724# a_11827_44484# 0.062801f
C2761 a_8199_44636# a_9159_44484# 4.07e-19
C2762 a_8016_46348# a_n2661_42834# 0.041785f
C2763 a_10227_46804# a_15095_43370# 0.264777f
C2764 a_310_45028# a_n2661_43370# 0.027265f
C2765 a_2324_44458# a_5205_44734# 5.38e-19
C2766 a_10053_45546# a_8953_45002# 0.009534f
C2767 a_12861_44030# a_15681_43442# 0.137136f
C2768 a_2124_47436# a_765_45546# 0.003536f
C2769 a_n881_46662# a_5263_46660# 2.48e-19
C2770 a_n1613_43370# a_5429_46660# 0.001925f
C2771 VDAC_N C10_N_btm 0.24639p
C2772 a_n743_46660# a_383_46660# 0.035839f
C2773 a_n2438_43548# a_601_46902# 0.043115f
C2774 a_n133_46660# a_33_46660# 0.580914f
C2775 a_n3565_37414# VIN_P 0.029764f
C2776 a_4915_47217# a_14180_46812# 0.017902f
C2777 a_13717_47436# a_15227_44166# 2.25e-20
C2778 a_12861_44030# a_18834_46812# 4.27e-19
C2779 a_n1925_46634# a_948_46660# 0.006613f
C2780 a_5088_37509# RST_Z 0.059771f
C2781 a_n2661_46634# a_1110_47026# 1.44e-19
C2782 a_n4209_37414# VREF 0.056254f
C2783 a_15811_47375# a_3090_45724# 1.43e-19
C2784 a_11599_46634# a_15368_46634# 0.320705f
C2785 a_10227_46804# a_11901_46660# 0.055248f
C2786 a_5700_37509# VDD 1.0734f
C2787 a_1414_42308# a_3318_42354# 0.001376f
C2788 a_9313_44734# a_22775_42308# 0.011571f
C2789 a_11967_42832# a_14456_42282# 4.2e-20
C2790 a_n4318_39768# a_n3674_37592# 0.024842f
C2791 a_7705_45326# VDD 0.211554f
C2792 a_19319_43548# a_19987_42826# 8.72e-20
C2793 a_3626_43646# a_1847_42826# 3.62e-21
C2794 a_n1441_43940# COMP_P 2.51e-20
C2795 a_10341_43396# a_16823_43084# 0.044262f
C2796 a_16243_43396# a_17324_43396# 0.102355f
C2797 a_16409_43396# a_16759_43396# 0.20669f
C2798 a_16547_43609# a_17499_43370# 1.26e-20
C2799 a_16137_43396# a_18429_43548# 9.56e-19
C2800 a_2982_43646# a_2905_42968# 3.17e-20
C2801 a_n97_42460# a_13113_42826# 4.45e-21
C2802 a_16147_45260# a_17970_44736# 2.03e-19
C2803 a_18175_45572# a_17767_44458# 6.65e-20
C2804 a_4646_46812# a_7765_42852# 0.122773f
C2805 a_3090_45724# a_15868_43402# 2.14e-21
C2806 a_n443_42852# a_n1899_43946# 2.87e-20
C2807 a_11787_45002# a_n2661_43370# 0.00108f
C2808 a_1823_45246# a_4905_42826# 0.110836f
C2809 a_n357_42282# a_2889_44172# 4.18e-22
C2810 a_6171_45002# a_13807_45067# 1.73e-19
C2811 a_n2840_45546# a_n4318_39768# 7.96e-20
C2812 a_n443_46116# a_2351_42308# 2.33e-20
C2813 a_14976_45028# a_15227_46910# 0.060892f
C2814 a_3090_45724# a_13059_46348# 0.167043f
C2815 a_15009_46634# a_16388_46812# 3.35e-20
C2816 a_16327_47482# a_16375_45002# 0.032962f
C2817 a_n743_46660# a_13351_46090# 0.008315f
C2818 a_n2109_47186# a_5263_45724# 9.21e-19
C2819 a_n881_46662# a_518_46155# 3.47e-19
C2820 a_11813_46116# a_765_45546# 0.003083f
C2821 a_4883_46098# a_9751_46155# 3.69e-19
C2822 a_19321_45002# a_20075_46420# 9.9e-20
C2823 a_20916_46384# a_18819_46122# 7.33e-21
C2824 a_19594_46812# a_19335_46494# 2.8e-19
C2825 a_2107_46812# a_9823_46155# 0.002289f
C2826 a_13747_46662# a_20708_46348# 2.93e-21
C2827 a_5807_45002# a_6945_45028# 0.057813f
C2828 a_3877_44458# a_167_45260# 5.06e-20
C2829 a_n443_46116# a_n357_42282# 0.153614f
C2830 a_4791_45118# a_n755_45592# 0.001705f
C2831 a_4651_46660# a_1823_45246# 0.001115f
C2832 a_10227_46804# a_15194_46482# 0.002224f
C2833 a_13507_46334# a_12005_46436# 7.68e-21
C2834 a_18083_42858# a_18599_43230# 0.113784f
C2835 a_17333_42852# a_18817_42826# 1.28e-19
C2836 a_8685_43396# a_5934_30871# 4.81e-19
C2837 a_7466_43396# a_6123_31319# 4.05e-20
C2838 a_3626_43646# a_15486_42560# 0.005343f
C2839 a_2982_43646# a_15803_42450# 4.86e-19
C2840 a_743_42282# a_20256_43172# 0.00713f
C2841 a_11691_44458# a_10617_44484# 1.65e-20
C2842 a_7229_43940# a_6453_43914# 0.001044f
C2843 a_5205_44484# a_7542_44172# 3.34e-20
C2844 a_n443_42852# a_14358_43442# 0.037176f
C2845 a_10193_42453# a_2982_43646# 0.231527f
C2846 a_11827_44484# a_n2661_43922# 0.32722f
C2847 a_526_44458# a_791_42968# 7.15e-19
C2848 a_n1925_42282# a_685_42968# 1.12e-20
C2849 a_n2661_44458# a_7640_43914# 0.005176f
C2850 a_626_44172# a_n2065_43946# 1.31e-21
C2851 a_375_42282# a_n1899_43946# 8.99e-21
C2852 a_n2312_38680# a_n4334_40480# 3.37e-19
C2853 a_n2017_45002# a_10807_43548# 0.0319f
C2854 a_16327_47482# a_413_45260# 2.72e-19
C2855 a_5937_45572# a_2324_44458# 0.407894f
C2856 a_5257_43370# a_6812_45938# 3.92e-20
C2857 a_n2293_46098# a_835_46155# 2.73e-19
C2858 a_3090_45724# a_3218_45724# 0.100752f
C2859 a_13059_46348# a_15002_46116# 1.85e-19
C2860 a_12549_44172# a_19431_45546# 1.86e-19
C2861 a_6969_46634# a_6472_45840# 2.28e-19
C2862 a_6755_46942# a_6511_45714# 2.73e-20
C2863 a_n1151_42308# a_14180_45002# 1.97e-20
C2864 a_584_46384# a_1307_43914# 0.314947f
C2865 a_6151_47436# a_8953_45002# 4.09e-20
C2866 a_n2109_47186# a_5837_45348# 8.23e-19
C2867 a_n971_45724# a_2903_45348# 0.004883f
C2868 a_21671_42860# a_13258_32519# 6.52e-20
C2869 a_5649_42852# a_7754_40130# 6.15e-19
C2870 a_564_42282# a_1067_42314# 1.81e-19
C2871 a_n327_42558# a_1184_42692# 1.76e-19
C2872 a_n784_42308# a_961_42354# 0.038477f
C2873 a_2982_43646# VDD 1.40372f
C2874 a_4646_46812# DATA[3] 0.001949f
C2875 a_n2293_43922# a_n2661_42282# 0.133253f
C2876 a_n2661_42834# a_7584_44260# 1.21e-19
C2877 a_3422_30871# a_19237_31679# 1.04e-19
C2878 a_n913_45002# a_21487_43396# 7.6e-21
C2879 a_n2017_45002# a_13467_32519# 2.68e-20
C2880 a_n356_44636# a_15493_43940# 9.87e-21
C2881 a_6540_46812# VDD 0.084698f
C2882 a_n2293_42834# a_6547_43396# 3.28e-20
C2883 a_9313_44734# a_12429_44172# 9.29e-21
C2884 a_19963_31679# a_17364_32525# 0.053794f
C2885 a_20447_31679# a_14209_32519# 0.051502f
C2886 en_comp a_4190_30871# 0.086973f
C2887 a_n863_45724# a_196_42282# 1.25e-19
C2888 a_n357_42282# a_n4318_37592# 4.71e-21
C2889 a_15415_45028# a_10341_43396# 3.51e-21
C2890 a_1423_45028# a_9803_43646# 3.46e-20
C2891 a_16979_44734# a_14021_43940# 3.43e-21
C2892 a_4223_44672# a_9165_43940# 1.39e-19
C2893 a_1307_43914# a_15095_43370# 1.5e-20
C2894 a_n2956_38216# a_n3674_37592# 0.025763f
C2895 a_13507_46334# a_9313_44734# 0.145766f
C2896 a_8049_45260# a_6511_45714# 0.001936f
C2897 a_7577_46660# a_8560_45348# 3.58e-21
C2898 a_n2312_38680# a_n2661_44458# 1.97e-21
C2899 a_14084_46812# a_14180_45002# 1.82e-22
C2900 a_n2810_45572# a_n2472_45546# 0.002308f
C2901 a_11415_45002# a_21350_45938# 8.06e-20
C2902 a_n2840_45546# a_n2956_38216# 0.019918f
C2903 a_10903_43370# a_12016_45572# 3.71e-20
C2904 a_14976_45028# a_9482_43914# 6.03e-19
C2905 a_3090_45724# a_13556_45296# 0.032207f
C2906 a_12549_44172# a_13076_44458# 5.14e-20
C2907 a_12891_46348# a_13720_44458# 8.1e-19
C2908 a_n2293_46634# a_n2129_44697# 5.68e-19
C2909 a_768_44030# a_12883_44458# 6.59e-19
C2910 a_6945_45028# a_15143_45578# 1.11e-21
C2911 a_n1741_47186# a_n971_45724# 0.157081f
C2912 a_n1605_47204# a_n815_47178# 2.38e-19
C2913 a_n2109_47186# a_n237_47217# 0.730469f
C2914 a_n2497_47436# a_n785_47204# 4.85e-19
C2915 SMPL_ON_P a_n452_47436# 3.73e-21
C2916 a_22400_42852# a_22609_38406# 1.37e-20
C2917 a_1606_42308# a_n3420_37440# 0.001369f
C2918 a_21887_42336# a_21973_42336# 0.006584f
C2919 a_21613_42308# a_22465_38105# 0.026117f
C2920 a_5837_42852# VDD 0.1774f
C2921 COMP_P a_11206_38545# 0.002821f
C2922 a_3905_42865# a_3539_42460# 0.022817f
C2923 a_n23_44458# a_n13_43084# 7.92e-19
C2924 a_2382_45260# a_2713_42308# 1.18e-20
C2925 a_19279_43940# a_10341_43396# 9.98e-20
C2926 a_n2017_45002# a_6773_42558# 0.001353f
C2927 a_9313_44734# a_21855_43396# 2.95e-19
C2928 a_n913_45002# a_5932_42308# 0.220872f
C2929 a_n2661_42282# a_n97_42460# 0.025699f
C2930 a_5883_43914# a_8952_43230# 3.2e-19
C2931 a_9838_44484# a_9127_43156# 8.54e-21
C2932 a_13259_45724# a_15595_45028# 2.25e-19
C2933 a_18189_46348# a_11827_44484# 1.03e-19
C2934 a_3483_46348# a_8701_44490# 1.31e-20
C2935 a_n755_45592# a_3429_45260# 2.78e-19
C2936 a_n23_45546# a_n37_45144# 0.001445f
C2937 a_n2293_46634# a_15493_43396# 4.09e-19
C2938 a_13507_46334# a_20974_43370# 0.017855f
C2939 a_19900_46494# a_19778_44110# 9.85e-21
C2940 a_20075_46420# a_18184_42460# 1.99e-20
C2941 a_2957_45546# a_2382_45260# 2.8e-21
C2942 a_n357_42282# a_3537_45260# 0.200175f
C2943 a_13059_46348# a_14815_43914# 0.004368f
C2944 a_3090_45724# a_20362_44736# 1.21e-21
C2945 a_5204_45822# a_4223_44672# 5.85e-20
C2946 a_2324_44458# a_11691_44458# 0.045025f
C2947 a_16375_45002# a_14537_43396# 3.44e-20
C2948 a_12549_44172# a_15301_44260# 4.3e-19
C2949 a_n3420_37984# C6_P_btm 1.22e-19
C2950 a_n3565_38216# C4_P_btm 9.91e-21
C2951 a_12891_46348# a_12549_44172# 0.309821f
C2952 a_6491_46660# a_6540_46812# 0.079263f
C2953 a_4791_45118# a_5429_46660# 6.03e-19
C2954 a_n2860_39072# VDD 0.004184f
C2955 a_n971_45724# a_7832_46660# 0.013782f
C2956 a_n2312_40392# a_n2293_46634# 4.37e-19
C2957 a_n2312_39304# a_n2442_46660# 0.15211f
C2958 a_2063_45854# a_10428_46928# 0.04306f
C2959 a_n1151_42308# a_7927_46660# 5.63e-20
C2960 a_7754_39964# a_n923_35174# 3.06e-20
C2961 a_n4209_39304# VIN_P 0.049722f
C2962 a_19963_31679# a_21589_35634# 1.55e-20
C2963 a_2982_43646# a_16137_43396# 5.37e-19
C2964 a_n356_44636# a_5742_30871# 0.120133f
C2965 a_14539_43914# a_15803_42450# 1.18e-22
C2966 a_11341_43940# a_12545_42858# 1.16e-20
C2967 a_8685_43396# a_7221_43396# 7.37e-21
C2968 a_n97_42460# a_16823_43084# 0.205258f
C2969 a_14401_32519# a_13678_32519# 0.050672f
C2970 a_21381_43940# a_5649_42852# 1.8e-20
C2971 a_20974_43370# a_21855_43396# 0.029556f
C2972 a_18597_46090# a_21195_42852# 0.01512f
C2973 a_526_44458# a_3905_42865# 0.321601f
C2974 a_n913_45002# a_1423_45028# 1.35e-22
C2975 a_12594_46348# a_12429_44172# 5.47e-22
C2976 a_6194_45824# a_6109_44484# 1.36e-19
C2977 a_n1925_42282# a_3600_43914# 2.11e-19
C2978 a_5111_44636# a_8953_45002# 3.17e-19
C2979 a_13507_46334# a_18599_43230# 0.00421f
C2980 a_6171_45002# a_7229_43940# 0.010208f
C2981 a_3232_43370# a_6709_45028# 0.086072f
C2982 a_16333_45814# a_16237_45028# 5.69e-20
C2983 a_16855_45546# a_11691_44458# 5.15e-22
C2984 a_13259_45724# a_18005_44484# 3.54e-19
C2985 a_3090_45724# a_6293_42852# 0.003062f
C2986 a_16147_45260# a_16501_45348# 9.04e-19
C2987 a_10193_42453# a_14539_43914# 0.278963f
C2988 a_11962_45724# a_12607_44458# 5.74e-21
C2989 a_n1613_43370# a_10083_42826# 1.52e-19
C2990 a_768_44030# a_3935_42891# 2.15e-21
C2991 a_13507_46334# a_12594_46348# 3.5e-19
C2992 a_4883_46098# a_10903_43370# 0.025531f
C2993 a_11599_46634# a_20708_46348# 1.58e-20
C2994 a_10467_46802# a_11901_46660# 0.001328f
C2995 a_10249_46116# a_11186_47026# 0.172467f
C2996 a_n881_46662# a_3147_46376# 0.073958f
C2997 a_n1613_43370# a_3483_46348# 0.029573f
C2998 a_16327_47482# a_18985_46122# 0.051538f
C2999 a_14311_47204# a_6945_45028# 0.008982f
C3000 a_n1741_47186# a_12005_46436# 5.93e-20
C3001 a_n443_46116# a_518_46155# 0.001648f
C3002 a_1110_47026# a_765_45546# 2.11e-20
C3003 a_10227_46804# a_17583_46090# 8.3e-22
C3004 a_17591_47464# a_17715_44484# 0.001482f
C3005 a_12861_44030# a_10809_44734# 0.156561f
C3006 a_7832_46660# a_8023_46660# 4.61e-19
C3007 a_21588_30879# a_11415_45002# 2.68e-19
C3008 a_n237_47217# a_8062_46155# 1.73e-19
C3009 a_5649_42852# a_18249_42858# 2.71e-20
C3010 a_14539_43914# VDD 0.873589f
C3011 a_4520_42826# a_5111_42852# 0.047152f
C3012 a_4361_42308# a_19339_43156# 3.07e-21
C3013 a_14358_43442# a_14635_42282# 9.06e-19
C3014 a_14205_43396# a_13291_42460# 6.79e-20
C3015 a_15493_43940# a_18727_42674# 1.18e-21
C3016 a_11341_43940# a_19332_42282# 5.32e-21
C3017 a_1756_43548# a_1755_42282# 1.07e-19
C3018 a_2982_43646# a_n784_42308# 0.026817f
C3019 a_n3674_39768# a_n4064_39072# 2.52e-21
C3020 a_19862_44208# a_19647_42308# 1.12e-20
C3021 a_17715_44484# a_17678_43396# 5.41e-20
C3022 a_19963_31679# a_19237_31679# 0.05162f
C3023 a_20447_31679# a_17730_32519# 0.051365f
C3024 a_5807_45002# a_14456_42282# 3.82e-19
C3025 a_13661_43548# a_13575_42558# 1.71e-20
C3026 a_9482_43914# a_15433_44458# 0.20244f
C3027 a_13556_45296# a_14815_43914# 0.378519f
C3028 a_n2293_42834# a_n356_44636# 0.027771f
C3029 a_n1059_45260# a_3422_30871# 7.02e-20
C3030 a_10903_43370# a_5649_42852# 9.98e-20
C3031 a_n357_42282# a_1049_43396# 0.001179f
C3032 a_11823_42460# a_14021_43940# 0.034191f
C3033 a_3090_45724# a_11554_42852# 0.001994f
C3034 a_13507_46334# a_15037_45618# 1.52e-20
C3035 a_8270_45546# a_8062_46155# 8.57e-21
C3036 a_17339_46660# a_17583_46090# 0.004328f
C3037 a_765_45546# a_15682_46116# 0.005634f
C3038 SMPL_ON_P a_n2472_45002# 1.75e-19
C3039 a_n2497_47436# a_n913_45002# 0.019337f
C3040 a_2959_46660# a_3316_45546# 5.39e-21
C3041 a_n2661_46634# a_6598_45938# 2.77e-21
C3042 a_12549_44172# a_11322_45546# 0.001723f
C3043 a_n2293_46098# a_3483_46348# 0.044283f
C3044 a_805_46414# a_1208_46090# 0.002746f
C3045 a_472_46348# a_1176_45822# 0.146555f
C3046 a_376_46348# a_1138_42852# 3.05e-21
C3047 a_1431_47204# a_2437_43646# 0.001971f
C3048 a_n881_46662# a_13249_42308# 9.77e-19
C3049 a_14180_46812# a_10809_44734# 0.012862f
C3050 a_3877_44458# a_n863_45724# 4.38e-21
C3051 a_10227_46804# a_8696_44636# 0.089585f
C3052 a_2253_43940# VDD 0.156797f
C3053 a_13467_32519# a_21973_42336# 0.00115f
C3054 a_10341_42308# a_11551_42558# 1.68e-19
C3055 a_12089_42308# a_11323_42473# 2.1e-19
C3056 a_20749_43396# a_20712_42282# 1.09e-20
C3057 a_13887_32519# a_22775_42308# 0.006279f
C3058 a_22591_43396# a_21613_42308# 2.05e-21
C3059 a_7499_43078# a_8387_43230# 0.008868f
C3060 a_5111_44636# a_3626_43646# 1.57e-19
C3061 a_742_44458# a_n2661_42282# 8.96e-21
C3062 a_n1925_42282# a_n1329_42308# 5.81e-19
C3063 a_8953_45546# a_9223_42460# 0.166987f
C3064 a_8016_46348# a_9885_42558# 5.79e-20
C3065 a_8128_46384# DATA[4] 6.38e-19
C3066 a_4185_45028# a_13575_42558# 8.71e-20
C3067 a_11827_44484# a_20935_43940# 0.003973f
C3068 a_3232_43370# a_2896_43646# 1.75e-19
C3069 a_n699_43396# a_3499_42826# 1.7e-19
C3070 a_n356_44636# a_1115_44172# 0.006316f
C3071 a_n2661_44458# a_10729_43914# 1.94e-19
C3072 a_13259_45724# a_13569_43230# 1.73e-19
C3073 a_2711_45572# a_18083_42858# 4.96e-19
C3074 a_2107_46812# a_1423_45028# 0.022467f
C3075 a_11133_46155# a_2711_45572# 1.16e-20
C3076 a_5937_45572# a_6667_45809# 0.002606f
C3077 a_4646_46812# a_7705_45326# 0.003014f
C3078 a_5732_46660# a_3232_43370# 2.77e-21
C3079 a_5907_46634# a_6171_45002# 1.1e-20
C3080 a_11415_45002# a_10907_45822# 0.050963f
C3081 a_17339_46660# a_8696_44636# 6.71e-19
C3082 a_n881_46662# a_17613_45144# 0.001826f
C3083 a_11735_46660# a_2437_43646# 6.77e-20
C3084 a_13507_46334# a_18114_32519# 0.001272f
C3085 a_2324_44458# a_n443_42852# 2.42e-19
C3086 a_n1379_46482# a_n2293_45546# 1.3e-20
C3087 a_8049_45260# a_11601_46155# 6.51e-19
C3088 a_8667_46634# a_413_45260# 2.03e-20
C3089 a_n1151_42308# a_n1655_44484# 1.11e-19
C3090 w_1575_34946# a_3422_30871# 1.88476f
C3091 a_7871_42858# VDD 0.395222f
C3092 a_8325_42308# a_7174_31319# 4.88e-21
C3093 a_5342_30871# C9_P_btm 5.28e-19
C3094 a_5534_30871# C7_P_btm 0.060228f
C3095 a_14113_42308# a_16522_42674# 0.183181f
C3096 a_13249_42308# a_13333_42558# 0.004402f
C3097 en_comp a_14635_42282# 4.34e-21
C3098 a_11823_42460# a_15764_42576# 4.46e-19
C3099 a_5891_43370# a_8317_43396# 5.61e-21
C3100 a_10193_42453# a_11897_42308# 0.00383f
C3101 a_n1059_45260# a_18504_43218# 2.15e-20
C3102 a_472_46348# DATA[0] 3.54e-20
C3103 a_19279_43940# a_n97_42460# 1.72e-21
C3104 a_14539_43914# a_16137_43396# 0.004691f
C3105 a_n2661_42834# a_8791_43396# 4.78e-20
C3106 a_n2661_43922# a_8147_43396# 2.31e-21
C3107 a_1823_45246# VDD 1.7584f
C3108 a_2998_44172# a_3992_43940# 5.62e-19
C3109 a_3600_43914# a_3737_43940# 0.126609f
C3110 a_n2956_38216# a_n2302_39072# 3.61e-19
C3111 a_18479_47436# a_19862_44208# 0.138185f
C3112 a_11453_44696# a_10729_43914# 5.66e-20
C3113 a_n2497_47436# a_n4318_39304# 3.31e-20
C3114 a_4791_45118# a_5326_44056# 1.55e-19
C3115 a_15682_46116# a_16751_45260# 3.1e-20
C3116 a_10490_45724# a_11652_45724# 0.044431f
C3117 a_8746_45002# a_11962_45724# 1.72e-21
C3118 a_10180_45724# a_11823_42460# 1.16e-20
C3119 a_2711_45572# a_11688_45572# 7.53e-19
C3120 a_12741_44636# a_20567_45036# 0.007778f
C3121 a_12465_44636# a_12429_44172# 0.003194f
C3122 a_10809_44734# a_11787_45002# 0.007368f
C3123 a_n1925_42282# a_4558_45348# 0.001226f
C3124 a_8270_45546# a_8375_44464# 1.34e-20
C3125 a_11415_45002# a_21359_45002# 0.015551f
C3126 a_20202_43084# a_11827_44484# 0.032881f
C3127 a_768_44030# a_6453_43914# 0.006009f
C3128 a_15227_44166# a_18248_44752# 0.001323f
C3129 a_3483_46348# a_8704_45028# 7.47e-19
C3130 a_2804_46116# a_n2661_43370# 1.16e-20
C3131 a_7227_45028# a_8120_45572# 1.01e-19
C3132 a_11322_45546# a_11525_45546# 0.055031f
C3133 a_18597_46090# a_15493_43396# 1.64e-21
C3134 a_n4315_30879# a_n1838_35608# 2.23e-19
C3135 a_n2109_47186# a_1123_46634# 3.71e-19
C3136 a_n746_45260# a_n1021_46688# 8.61e-21
C3137 a_n237_47217# a_n1925_46634# 0.079348f
C3138 a_13507_46334# a_12465_44636# 0.029101f
C3139 a_n3565_38502# a_n3565_37414# 0.030671f
C3140 a_n4209_38502# a_n3420_37440# 0.033073f
C3141 a_n3420_38528# a_n4209_37414# 0.027951f
C3142 a_1431_47204# a_n2661_46634# 0.001833f
C3143 a_6151_47436# a_13675_47204# 0.002433f
C3144 a_21496_47436# a_21811_47423# 3.73e-19
C3145 a_9313_45822# a_9804_47204# 0.171044f
C3146 a_12861_44030# a_n881_46662# 0.135351f
C3147 a_4958_30871# C2_N_btm 9.53e-20
C3148 a_19787_47423# a_11453_44696# 1.96e-19
C3149 a_n971_45724# a_n743_46660# 0.122713f
C3150 a_n452_47436# a_n2438_43548# 3.48e-19
C3151 a_n2661_42282# a_n901_43156# 5.27e-20
C3152 a_9313_44734# a_14853_42852# 4.55e-21
C3153 a_n2810_45028# a_n4064_37984# 0.002525f
C3154 a_15493_43396# a_743_42282# 1.59e-19
C3155 a_12427_45724# VDD 0.33808f
C3156 a_458_43396# a_648_43396# 0.045837f
C3157 a_4235_43370# a_3626_43646# 1.4e-19
C3158 a_4093_43548# a_3539_42460# 0.001457f
C3159 a_3080_42308# a_2982_43646# 0.095684f
C3160 a_n97_42460# a_7112_43396# 0.002373f
C3161 a_14021_43940# a_18429_43548# 0.00816f
C3162 a_19862_44208# a_4190_30871# 0.023868f
C3163 a_n2956_37592# a_n2946_37984# 0.004313f
C3164 a_4223_44672# a_3823_42558# 7.52e-22
C3165 a_3422_30871# a_19987_42826# 0.006447f
C3166 a_3316_45546# a_n699_43396# 1.1e-20
C3167 a_n755_45592# a_8103_44636# 4.46e-21
C3168 a_16680_45572# a_16751_45260# 9.83e-19
C3169 a_15861_45028# a_16019_45002# 0.04712f
C3170 a_8696_44636# a_1307_43914# 0.030679f
C3171 a_n2840_45002# a_n2661_45010# 0.189331f
C3172 a_n2293_46634# a_10695_43548# 0.007256f
C3173 a_3090_45724# a_7499_43940# 0.025901f
C3174 a_12549_44172# a_16409_43396# 3.09e-19
C3175 a_1823_45246# a_5495_43940# 0.001058f
C3176 a_13507_46334# a_13887_32519# 0.08088f
C3177 a_19900_46494# a_20159_44458# 7.47e-21
C3178 a_20075_46420# a_20362_44736# 4.79e-20
C3179 a_4646_46812# a_2982_43646# 2.9e-20
C3180 a_10227_46804# a_20885_46660# 0.001925f
C3181 VDD DATA[2] 0.3216f
C3182 a_2063_45854# a_7920_46348# 3.54e-19
C3183 a_n1151_42308# a_5164_46348# 0.110485f
C3184 a_12465_44636# a_20623_46660# 4.37e-20
C3185 a_18597_46090# a_18900_46660# 0.00136f
C3186 a_4646_46812# a_6540_46812# 0.029952f
C3187 a_4651_46660# a_5732_46660# 0.102355f
C3188 a_3877_44458# a_5072_46660# 0.021873f
C3189 a_n1925_46634# a_8270_45546# 0.109762f
C3190 a_5807_45002# a_15559_46634# 0.006621f
C3191 a_16131_47204# a_16292_46812# 2.31e-19
C3192 a_13661_43548# a_15368_46634# 3.74e-20
C3193 a_4791_45118# a_3483_46348# 0.088998f
C3194 a_n443_46116# a_3147_46376# 0.002662f
C3195 a_4007_47204# a_4185_45028# 7.03e-19
C3196 a_n1435_47204# a_n1991_46122# 1.76e-20
C3197 a_n881_46662# a_14180_46812# 0.028137f
C3198 C5_N_btm VIN_N 0.502041f
C3199 a_21811_47423# a_21363_46634# 0.010128f
C3200 a_4883_46098# a_21188_46660# 0.012559f
C3201 a_4817_46660# a_5167_46660# 0.218775f
C3202 a_n1741_47186# a_12594_46348# 0.150956f
C3203 a_11453_44696# a_20107_46660# 0.050203f
C3204 a_13507_46334# a_20528_46660# 0.00277f
C3205 C3_N_btm VREF_GND 0.67174f
C3206 C2_N_btm VCM 0.716172f
C3207 C4_N_btm VREF 0.98728f
C3208 a_13747_46662# a_14976_45028# 0.016638f
C3209 a_n2661_46634# a_11735_46660# 0.044956f
C3210 a_n237_47217# a_10355_46116# 1.06e-20
C3211 a_14579_43548# a_5534_30871# 0.030066f
C3212 a_14358_43442# a_14543_43071# 0.001166f
C3213 a_9028_43914# a_9223_42460# 3.81e-21
C3214 a_13467_32519# a_14209_32519# 0.048306f
C3215 a_13678_32519# a_22223_43396# 0.004894f
C3216 a_21855_43396# a_13887_32519# 3.59e-19
C3217 a_20556_43646# a_20749_43396# 0.018955f
C3218 a_n2661_43370# CLK 0.011991f
C3219 a_4905_42826# a_5193_42852# 0.016389f
C3220 a_4361_42308# a_22591_43396# 2.7e-19
C3221 a_10341_43396# a_12545_42858# 8.88e-20
C3222 a_14309_45028# VDD 0.189806f
C3223 a_6171_45002# a_15004_44636# 4.14e-20
C3224 a_2711_45572# a_12429_44172# 3.56e-22
C3225 a_3090_45724# a_10991_42826# 0.004747f
C3226 a_1423_45028# a_n2661_44458# 0.164701f
C3227 a_n1059_45260# a_7640_43914# 6.31e-21
C3228 a_4646_46812# a_5837_42852# 1.26e-20
C3229 a_10903_43370# a_8685_43396# 0.031035f
C3230 a_413_45260# a_n356_44636# 5.61e-19
C3231 a_n37_45144# a_n23_44458# 4.88e-19
C3232 a_14309_45348# a_14309_45028# 6.96e-20
C3233 a_9482_43914# a_5343_44458# 2.61e-20
C3234 a_526_44458# a_4093_43548# 0.107158f
C3235 a_6755_46942# a_15015_46420# 0.133517f
C3236 a_8270_45546# a_10355_46116# 2.83e-19
C3237 a_4915_47217# a_13904_45546# 0.013453f
C3238 a_n881_46662# a_310_45028# 7.88e-19
C3239 a_20841_46902# a_20731_47026# 0.097745f
C3240 a_21363_46634# a_22000_46634# 0.017308f
C3241 a_20623_46660# a_20528_46660# 0.049827f
C3242 a_19123_46287# a_18900_46660# 0.001018f
C3243 a_2107_46812# a_9823_46482# 2.17e-19
C3244 a_13507_46334# a_2711_45572# 9.2e-19
C3245 a_n1613_43370# a_n357_42282# 0.030838f
C3246 a_3090_45724# a_4704_46090# 4.99e-19
C3247 a_2063_45854# a_11280_45822# 0.009384f
C3248 a_15743_43084# a_14113_42308# 5.99e-20
C3249 a_n3674_39768# VDD 0.398971f
C3250 a_13678_32519# a_5934_30871# 2.14e-19
C3251 a_4361_42308# a_3905_42308# 3.53e-19
C3252 a_17701_42308# a_17665_42852# 0.002723f
C3253 a_17595_43084# a_17749_42852# 0.010303f
C3254 a_17333_42852# a_16245_42852# 1.21e-20
C3255 a_5649_42852# a_7963_42308# 5.44e-20
C3256 a_743_42282# a_8791_42308# 0.008346f
C3257 a_7871_42858# a_n784_42308# 4.17e-21
C3258 a_10341_43396# a_19332_42282# 2.01e-21
C3259 a_4915_47217# CLK 0.198293f
C3260 a_n863_45724# a_1847_42826# 0.216819f
C3261 a_n2661_45546# a_4520_42826# 2.03e-19
C3262 a_13259_45724# a_13113_42826# 1.98e-19
C3263 a_14797_45144# a_11341_43940# 1.37e-20
C3264 a_15004_44636# a_14673_44172# 0.039287f
C3265 a_20447_31679# a_17538_32519# 0.051306f
C3266 a_n443_42852# a_n2157_42858# 8.79e-20
C3267 a_526_44458# a_5457_43172# 7.33e-19
C3268 a_6151_47436# DATA[4] 2.92e-19
C3269 a_9482_43914# a_9801_44260# 0.003952f
C3270 a_1823_45246# a_n784_42308# 6e-20
C3271 a_11823_42460# a_13943_43396# 0.006456f
C3272 a_10193_42453# a_17324_43396# 9.84e-20
C3273 a_18479_45785# a_2982_43646# 2.74e-20
C3274 a_6545_47178# DATA[3] 0.178561f
C3275 a_11031_47542# VDD 0.214104f
C3276 a_n1243_44484# a_n2661_42834# 1.91e-19
C3277 a_n2293_46098# a_n357_42282# 0.014918f
C3278 a_n1853_46287# a_n1099_45572# 0.067343f
C3279 a_765_45546# a_6598_45938# 2.98e-21
C3280 a_6755_46942# a_16333_45814# 0.001253f
C3281 a_2063_45854# a_11827_44484# 8.5e-20
C3282 a_15015_46420# a_8049_45260# 0.002448f
C3283 a_12594_46348# a_10586_45546# 8.27e-20
C3284 a_n2497_47436# a_n2661_44458# 0.138848f
C3285 a_805_46414# a_n2661_45546# 7.52e-20
C3286 a_768_44030# a_6171_45002# 0.027851f
C3287 a_n2293_46634# a_n745_45366# 0.006631f
C3288 a_n2442_46660# a_n2810_45028# 0.045466f
C3289 a_8128_46384# a_8191_45002# 2.38e-19
C3290 a_n2438_43548# a_n2472_45002# 0.023014f
C3291 a_n901_46420# a_n1079_45724# 1.93e-20
C3292 a_n1076_46494# a_n2293_45546# 7.13e-22
C3293 a_6123_31319# a_5934_30871# 15.8951f
C3294 a_17324_43396# VDD 0.274722f
C3295 a_3823_42558# a_5742_30871# 1.54e-20
C3296 a_4190_30871# C7_P_btm 2.94e-19
C3297 a_13678_32519# a_11530_34132# 0.002459f
C3298 a_3537_45260# a_8952_43230# 3.58e-20
C3299 a_11827_44484# a_14955_43396# 5.17e-21
C3300 a_20679_44626# a_15493_43940# 1.03e-19
C3301 a_19279_43940# a_21115_43940# 1.52e-19
C3302 a_18579_44172# a_20365_43914# 1.9e-19
C3303 a_5343_44458# a_6031_43396# 9.7e-21
C3304 a_n1059_45260# a_16414_43172# 0.094309f
C3305 a_n2017_45002# a_16795_42852# 6.5e-19
C3306 a_n2661_42834# a_10651_43940# 5.65e-20
C3307 a_21076_30879# a_22459_39145# 3.89e-20
C3308 a_5111_44636# a_8037_42858# 2.31e-19
C3309 a_n913_45002# a_15567_42826# 6.93e-20
C3310 a_7499_43078# a_1606_42308# 5.24e-20
C3311 a_375_42282# a_n2157_42858# 2.28e-21
C3312 a_1414_42308# a_2537_44260# 4.33e-19
C3313 a_7281_43914# a_7542_44172# 0.060549f
C3314 a_n23_44458# a_104_43370# 1.77e-20
C3315 a_15227_44166# EN_OFFSET_CAL 2.2e-20
C3316 a_21137_46414# a_20273_45572# 0.002347f
C3317 a_5204_45822# a_413_45260# 4.29e-21
C3318 a_20708_46348# a_20841_45814# 1.63e-19
C3319 a_6945_45028# a_20107_45572# 1.37e-19
C3320 a_2324_44458# a_2437_43646# 0.011046f
C3321 a_7715_46873# a_5343_44458# 2.03e-20
C3322 a_8049_45260# a_16333_45814# 0.002964f
C3323 a_8034_45724# a_8696_44636# 9.58e-21
C3324 a_11415_45002# a_15415_45028# 0.0035f
C3325 a_17609_46634# a_17613_45144# 4.03e-21
C3326 a_3147_46376# a_3537_45260# 1.82e-19
C3327 a_13507_46334# a_22485_44484# 0.008777f
C3328 a_13747_46662# a_15433_44458# 1.47e-21
C3329 a_n2293_46634# a_3363_44484# 0.001146f
C3330 a_3090_45724# a_19778_44110# 9.48e-19
C3331 a_8199_44636# en_comp 4.34e-21
C3332 a_15227_44166# a_16922_45042# 0.533576f
C3333 a_3483_46348# a_3429_45260# 4.53e-19
C3334 a_3699_46348# a_3065_45002# 3.29e-21
C3335 a_14275_46494# a_3357_43084# 4.55e-22
C3336 a_768_44030# a_14673_44172# 2.39e-20
C3337 a_6123_31319# a_11530_34132# 0.001062f
C3338 a_n4334_39392# a_n4334_38528# 0.050585f
C3339 a_n4209_39304# a_n3565_38502# 0.029672f
C3340 a_1606_42308# C8_N_btm 6.73e-20
C3341 a_5129_47502# a_n1435_47204# 4.12e-19
C3342 a_7227_47204# a_9067_47204# 3.76e-21
C3343 a_7903_47542# a_6575_47204# 0.046223f
C3344 a_6151_47436# a_11459_47204# 0.034818f
C3345 a_4915_47217# a_13717_47436# 4.05e-19
C3346 a_n3565_39304# a_n4209_38502# 5.79402f
C3347 a_n2946_39072# a_n2860_39072# 0.011479f
C3348 a_n3420_39072# a_n2216_39072# 7.08e-20
C3349 a_5934_30871# EN_VIN_BSTR_P 0.075302f
C3350 a_n1741_47186# a_12465_44636# 4.19e-22
C3351 a_1184_42692# VDD 0.813074f
C3352 a_14021_43940# a_2982_43646# 0.00345f
C3353 a_10729_43914# a_9145_43396# 2.31e-20
C3354 a_n2293_43922# a_12545_42858# 0.022686f
C3355 a_14955_43940# a_8685_43396# 2.16e-19
C3356 a_n2293_45546# VDD 2.06545f
C3357 a_n2293_42834# a_3823_42558# 2.98e-20
C3358 a_17730_32519# a_13467_32519# 0.054292f
C3359 a_20512_43084# a_13678_32519# 0.059475f
C3360 a_9313_44734# a_17701_42308# 0.008094f
C3361 a_20447_31679# a_22465_38105# 4.46e-19
C3362 a_n913_45002# a_20712_42282# 0.003267f
C3363 a_n1059_45260# a_7174_31319# 5.53e-20
C3364 en_comp a_19511_42282# 2.68e-20
C3365 a_12861_44030# a_14621_43646# 1.73e-20
C3366 a_7499_43078# a_10775_45002# 0.00194f
C3367 a_9049_44484# a_8953_45002# 0.031391f
C3368 a_11415_45002# a_19279_43940# 0.003698f
C3369 a_17786_45822# a_17668_45572# 1.98e-20
C3370 a_18341_45572# a_18799_45938# 0.027606f
C3371 a_18691_45572# a_19256_45572# 7.99e-20
C3372 a_n971_45724# a_4361_42308# 6.67e-20
C3373 a_5907_45546# a_1423_45028# 3.15e-20
C3374 a_11652_45724# a_6171_45002# 0.072138f
C3375 a_5937_45572# a_5708_44484# 5.12e-19
C3376 a_10227_46804# a_14205_43396# 0.422372f
C3377 a_526_44458# a_10157_44484# 4.13e-20
C3378 a_n1099_45572# a_n2661_43370# 2.12e-19
C3379 a_2324_44458# a_4181_44734# 3.09e-19
C3380 a_4883_46098# a_8685_43396# 0.011038f
C3381 a_6755_46942# a_15493_43396# 8.69e-20
C3382 a_1431_47204# a_765_45546# 0.00505f
C3383 a_n1613_43370# a_5263_46660# 7.38e-19
C3384 VDAC_N C9_N_btm 0.123386p
C3385 a_11599_46634# a_14976_45028# 0.020184f
C3386 a_n743_46660# a_601_46902# 0.022066f
C3387 a_n2438_43548# a_33_46660# 0.588568f
C3388 a_n133_46660# a_171_46873# 0.163873f
C3389 a_4915_47217# a_14035_46660# 0.075669f
C3390 a_12861_44030# a_17609_46634# 0.183853f
C3391 a_n1925_46634# a_1123_46634# 0.018809f
C3392 a_4338_37500# RST_Z 0.01719f
C3393 a_15811_47375# a_15009_46634# 2.23e-19
C3394 a_10227_46804# a_11813_46116# 0.094518f
C3395 a_5088_37509# VDD 1.15925f
C3396 a_9313_44734# a_21613_42308# 0.001498f
C3397 a_1414_42308# a_2903_42308# 1.7e-19
C3398 a_6709_45028# VDD 0.390566f
C3399 a_19319_43548# a_19164_43230# 7.09e-19
C3400 a_18326_43940# a_18504_43218# 2.4e-20
C3401 a_15781_43660# a_15743_43084# 0.050751f
C3402 a_8685_43396# a_5649_42852# 2.05e-20
C3403 a_10341_43396# a_17021_43396# 4.33e-19
C3404 a_n97_42460# a_12545_42858# 3.58e-19
C3405 a_16547_43609# a_16759_43396# 9.49e-19
C3406 a_16137_43396# a_17324_43396# 1.29e-20
C3407 a_16243_43396# a_17499_43370# 0.043633f
C3408 a_16409_43396# a_16977_43638# 0.17072f
C3409 a_10907_45822# a_n2661_43922# 2.58e-19
C3410 a_16147_45260# a_17767_44458# 1.74e-19
C3411 a_8049_45260# a_15493_43396# 6.61e-22
C3412 a_4646_46812# a_7871_42858# 0.26422f
C3413 a_15227_44166# a_15743_43084# 0.513622f
C3414 a_3218_45724# a_1414_42308# 3.53e-21
C3415 a_n443_42852# a_n1761_44111# 0.007283f
C3416 a_20447_31679# a_19721_31679# 0.070259f
C3417 a_10951_45334# a_n2661_43370# 0.004229f
C3418 a_1307_43914# a_5009_45028# 2.65e-20
C3419 a_1823_45246# a_3080_42308# 0.049986f
C3420 a_n357_42282# a_2675_43914# 1.8e-19
C3421 a_n755_45592# a_895_43940# 8.1e-20
C3422 a_6171_45002# a_13490_45067# 3.54e-19
C3423 a_16327_47482# a_20753_42852# 0.00568f
C3424 w_1575_34946# a_7174_31319# 0.001988f
C3425 a_15009_46634# a_13059_46348# 0.054389f
C3426 a_3090_45724# a_15227_46910# 0.010657f
C3427 a_n743_46660# a_12594_46348# 0.0427f
C3428 a_n2109_47186# a_4099_45572# 8.98e-22
C3429 a_n1151_42308# a_3316_45546# 5.6e-21
C3430 a_n443_46116# a_310_45028# 0.06667f
C3431 a_n881_46662# a_3873_46454# 0.003191f
C3432 a_11735_46660# a_765_45546# 0.006002f
C3433 a_4883_46098# a_11608_46482# 5.79e-19
C3434 a_19321_45002# a_19335_46494# 0.006071f
C3435 a_19594_46812# a_19553_46090# 8.61e-19
C3436 a_13747_46662# a_19900_46494# 0.001247f
C3437 a_16131_47204# a_6945_45028# 0.003013f
C3438 a_n2661_46634# a_2324_44458# 0.0278f
C3439 a_n1741_47186# a_2711_45572# 6.27e-20
C3440 a_2107_46812# a_9569_46155# 0.018199f
C3441 a_4791_45118# a_n357_42282# 0.020355f
C3442 a_4646_46812# a_1823_45246# 8.67e-19
C3443 a_11599_46634# a_18051_46116# 0.03664f
C3444 a_10227_46804# a_14949_46494# 6.03e-19
C3445 a_n97_42460# a_19332_42282# 2.35e-20
C3446 a_14401_32519# a_22775_42308# 3.78e-20
C3447 a_17333_42852# a_18249_42858# 0.311255f
C3448 a_18083_42858# a_18817_42826# 0.0532f
C3449 a_3626_43646# a_15051_42282# 0.009723f
C3450 a_2982_43646# a_15764_42576# 3.1e-19
C3451 a_7227_42852# a_7573_43172# 0.013377f
C3452 a_3935_42891# a_4149_42891# 0.005572f
C3453 a_n1352_44484# a_n1243_44484# 0.007416f
C3454 a_n1177_44458# a_n998_44484# 0.007399f
C3455 a_n452_44636# a_7_44811# 6.64e-19
C3456 a_5205_44484# a_7281_43914# 0.008497f
C3457 a_13259_45724# a_16823_43084# 0.017563f
C3458 a_n443_42852# a_14579_43548# 0.04846f
C3459 a_949_44458# a_n23_44458# 3.38e-20
C3460 a_11827_44484# a_n2661_42834# 0.046936f
C3461 a_526_44458# a_685_42968# 1.6e-19
C3462 a_n2956_39768# a_n4209_39590# 0.334714f
C3463 a_12741_44636# a_12800_43218# 3.89e-21
C3464 a_12607_44458# a_15004_44636# 1.81e-20
C3465 a_n2661_44458# a_6109_44484# 0.004386f
C3466 a_375_42282# a_n1761_44111# 1.36e-19
C3467 a_n2312_38680# a_n4315_30879# 0.024522f
C3468 a_n2442_46660# a_n2302_40160# 0.017419f
C3469 a_n1059_45260# a_10729_43914# 5.14e-23
C3470 a_n913_45002# a_10405_44172# 2.38e-20
C3471 SMPL_ON_N a_19963_31679# 0.029334f
C3472 a_16241_47178# a_413_45260# 8.41e-20
C3473 a_11189_46129# a_12594_46348# 0.001927f
C3474 a_8199_44636# a_2324_44458# 0.412215f
C3475 a_n1076_46494# a_n914_46116# 0.006453f
C3476 a_n743_46660# a_15037_45618# 3.95e-20
C3477 a_n1151_42308# a_13777_45326# 2.49e-21
C3478 a_3483_46348# a_6945_45028# 0.002307f
C3479 a_n2293_46098# a_518_46155# 3.23e-19
C3480 a_3090_45724# a_2957_45546# 0.167712f
C3481 a_11387_46155# a_10903_43370# 7.72e-19
C3482 a_n971_45724# a_2809_45348# 0.00154f
C3483 a_6755_46942# a_6472_45840# 1.91e-20
C3484 a_21195_42852# a_13258_32519# 1.05e-19
C3485 a_22165_42308# a_19511_42282# 1.52e-19
C3486 a_n784_42308# a_1184_42692# 0.026118f
C3487 a_564_42282# a_n1630_35242# 0.156633f
C3488 a_196_42282# a_961_42354# 1.2e-21
C3489 a_19987_42826# a_7174_31319# 6.85e-20
C3490 a_2896_43646# VDD 0.208317f
C3491 a_3877_44458# DATA[3] 1.85e-20
C3492 a_n2661_42834# a_6756_44260# 1.06e-19
C3493 a_8696_44636# a_13635_43156# 2.2e-22
C3494 a_n2810_45572# a_n1630_35242# 5.26e-19
C3495 a_5732_46660# VDD 0.277366f
C3496 a_9313_44734# a_11750_44172# 2.81e-21
C3497 a_3422_30871# a_22959_44484# 2.88e-19
C3498 a_22315_44484# a_17730_32519# 0.001043f
C3499 a_1423_45028# a_9145_43396# 3.76e-21
C3500 a_14539_43914# a_14021_43940# 0.043922f
C3501 a_5518_44484# a_5829_43940# 1.88e-20
C3502 a_n357_42282# a_n1736_42282# 2.32e-20
C3503 a_1307_43914# a_14205_43396# 1.03e-20
C3504 a_12741_44636# a_20528_45572# 0.006514f
C3505 a_11599_46634# a_15433_44458# 1.57e-21
C3506 a_10586_45546# a_2711_45572# 0.295169f
C3507 a_10809_44734# a_13904_45546# 9.68e-22
C3508 a_8034_45724# a_7227_45028# 2.26e-19
C3509 a_8049_45260# a_6472_45840# 4.08e-19
C3510 a_n2312_38680# a_n4318_40392# 0.023897f
C3511 a_n2810_45572# a_n2661_45546# 0.006676f
C3512 a_n2840_45546# a_n2472_45546# 7.52e-19
C3513 a_8016_46348# a_8696_44636# 0.031525f
C3514 a_20202_43084# a_21350_45938# 1.43e-19
C3515 a_11415_45002# a_19610_45572# 5.19e-19
C3516 a_5066_45546# a_5024_45822# 3.47e-19
C3517 a_5807_45002# a_6298_44484# 1.01e-19
C3518 a_10903_43370# a_11778_45572# 3.1e-20
C3519 a_n2293_46634# a_n2433_44484# 7.85e-20
C3520 a_3090_45724# a_9482_43914# 0.029795f
C3521 a_3483_46348# a_14127_45572# 1.22e-19
C3522 a_16721_46634# a_413_45260# 6.74e-22
C3523 a_526_44458# a_7499_43078# 0.2203f
C3524 a_12891_46348# a_13076_44458# 0.182315f
C3525 a_768_44030# a_12607_44458# 0.215512f
C3526 a_12549_44172# a_12883_44458# 7.5e-19
C3527 a_n1741_47186# a_n452_47436# 0.013149f
C3528 a_n1920_47178# a_n971_45724# 1.39e-20
C3529 a_n2109_47186# a_n746_45260# 0.295988f
C3530 SMPL_ON_P a_n815_47178# 0.002605f
C3531 a_n2833_47464# a_n785_47204# 5.95e-22
C3532 a_5742_30871# a_1177_38525# 1.05e-19
C3533 a_21613_42308# a_22397_42558# 0.001996f
C3534 a_21887_42336# a_22465_38105# 7.29e-21
C3535 a_7174_31319# a_n4315_30879# 6.67e-21
C3536 a_5193_42852# VDD 0.187605f
C3537 a_6123_31319# a_7754_40130# 6.87e-20
C3538 COMP_P VDAC_P 0.003408f
C3539 a_18451_43940# a_18797_44260# 0.013377f
C3540 a_3905_42865# a_3626_43646# 0.036343f
C3541 a_10809_44734# CLK 0.002918f
C3542 a_n2956_38216# a_n2860_37690# 8.73e-19
C3543 a_17061_44734# a_16409_43396# 1.3e-20
C3544 a_n1059_45260# a_5932_42308# 8.52e-19
C3545 a_n913_45002# a_6171_42473# 0.034189f
C3546 a_n2017_45002# a_6481_42558# 0.001353f
C3547 a_17973_43940# a_18533_43940# 5.23e-19
C3548 a_n914_46116# VDD 7.75e-19
C3549 a_20193_45348# a_21195_42852# 1.43e-20
C3550 a_5883_43914# a_9127_43156# 3.96e-19
C3551 a_9313_44734# a_4361_42308# 0.082952f
C3552 a_13259_45724# a_15415_45028# 1.67e-19
C3553 a_n1925_42282# a_n2661_43370# 0.027962f
C3554 a_17715_44484# a_11827_44484# 0.037803f
C3555 a_n755_45592# a_3065_45002# 0.027852f
C3556 a_n23_45546# a_n143_45144# 0.004979f
C3557 a_n356_45724# a_n37_45144# 0.001109f
C3558 a_3503_45724# a_413_45260# 7.76e-19
C3559 a_13507_46334# a_14401_32519# 0.001279f
C3560 a_20075_46420# a_19778_44110# 1.42e-20
C3561 a_3483_46348# a_8103_44636# 0.00166f
C3562 a_6194_45824# a_3357_43084# 0.004141f
C3563 a_10193_42453# a_18799_45938# 3.31e-21
C3564 a_14840_46494# a_11691_44458# 2.41e-21
C3565 a_5164_46348# a_4223_44672# 2.5e-21
C3566 a_4704_46090# a_4743_44484# 4.57e-21
C3567 a_12549_44172# a_15037_44260# 4.91e-19
C3568 a_n2312_39304# a_n2472_46634# 0.016291f
C3569 a_n2312_40392# a_n2442_46660# 5.91846f
C3570 a_n4209_38216# C3_P_btm 0.041776f
C3571 a_n3565_38216# C5_P_btm 1.11e-20
C3572 a_n3420_37984# C7_P_btm 2.68e-20
C3573 a_6491_46660# a_5732_46660# 6.78e-19
C3574 a_6545_47178# a_6540_46812# 0.013617f
C3575 a_4791_45118# a_5263_46660# 0.001102f
C3576 comp_n VDD 0.504719f
C3577 a_12465_44636# a_n743_46660# 0.026136f
C3578 a_2063_45854# a_10150_46912# 0.008885f
C3579 a_n1151_42308# a_8145_46902# 3.91e-20
C3580 a_18799_45938# VDD 0.132317f
C3581 a_19963_31679# a_19864_35138# 1.38e-21
C3582 a_20974_43370# a_4361_42308# 0.122936f
C3583 a_17538_32519# a_13467_32519# 0.051209f
C3584 a_n2293_43922# a_5379_42460# 0.4571f
C3585 a_n356_44636# a_11323_42473# 1.17e-19
C3586 a_20835_44721# a_20753_42852# 5.18e-21
C3587 a_20447_31679# a_18194_35068# 9.11e-20
C3588 a_17737_43940# a_17701_42308# 1.13e-19
C3589 a_n97_42460# a_17021_43396# 4.28e-19
C3590 a_14401_32519# a_21855_43396# 0.00125f
C3591 a_21381_43940# a_13678_32519# 5.1e-21
C3592 a_n2293_46098# a_5025_43940# 0.002209f
C3593 a_11962_45724# a_8975_43940# 3.26e-21
C3594 a_19692_46634# a_2982_43646# 0.003269f
C3595 a_15861_45028# a_11827_44484# 1.34e-19
C3596 a_n1059_45260# a_1423_45028# 8.02e-22
C3597 a_n1925_42282# a_2998_44172# 0.02835f
C3598 a_526_44458# a_3600_43914# 9.66e-19
C3599 a_5111_44636# a_8191_45002# 1.43e-20
C3600 a_10903_43370# a_13483_43940# 1.22e-19
C3601 a_2437_43646# a_2448_45028# 4.11e-19
C3602 a_13507_46334# a_18817_42826# 0.001318f
C3603 a_10193_42453# a_16112_44458# 1.55e-19
C3604 a_6431_45366# a_5205_44484# 0.018787f
C3605 a_6171_45002# a_7276_45260# 0.00899f
C3606 a_3232_43370# a_7229_43940# 0.180766f
C3607 a_16115_45572# a_11691_44458# 1.01e-20
C3608 a_3090_45724# a_6031_43396# 0.00482f
C3609 a_16147_45260# a_16405_45348# 0.001516f
C3610 a_n1613_43370# a_8952_43230# 0.213002f
C3611 a_768_44030# a_3681_42891# 1.91e-20
C3612 a_n2956_39768# a_n1853_43023# 1.99e-21
C3613 w_1575_34946# a_5932_42308# 0.0018f
C3614 a_4883_46098# a_11387_46155# 0.010865f
C3615 a_11599_46634# a_19900_46494# 0.055271f
C3616 a_10467_46802# a_11813_46116# 2.89e-19
C3617 a_10249_46116# a_10768_47026# 0.027091f
C3618 a_6755_46942# a_8846_46660# 8.14e-19
C3619 a_10428_46928# a_11901_46660# 0.004685f
C3620 a_n881_46662# a_2804_46116# 0.050669f
C3621 a_n1613_43370# a_3147_46376# 0.004069f
C3622 a_13507_46334# a_12005_46116# 2.73e-19
C3623 a_16327_47482# a_18819_46122# 0.324239f
C3624 a_n1151_42308# a_5066_45546# 0.5423f
C3625 a_19594_46812# a_12741_44636# 6.75e-20
C3626 a_13487_47204# a_6945_45028# 0.015556f
C3627 a_13717_47436# a_10809_44734# 0.004969f
C3628 a_20916_46384# a_11415_45002# 7.86e-20
C3629 a_17591_47464# a_17583_46090# 6.37e-19
C3630 a_10227_46804# a_15682_46116# 0.001531f
C3631 a_5649_42852# a_17333_42852# 1.49e-20
C3632 a_19478_44306# a_19647_42308# 2.55e-20
C3633 a_16112_44458# VDD 0.182397f
C3634 a_4361_42308# a_18599_43230# 9.24e-21
C3635 a_14579_43548# a_14635_42282# 0.124652f
C3636 a_1568_43370# a_1755_42282# 7.17e-19
C3637 a_3080_42308# a_1184_42692# 1.44e-20
C3638 a_1756_43548# a_1606_42308# 3.46e-19
C3639 a_n4318_39768# a_n4064_39072# 2.48e-21
C3640 a_n1557_42282# a_n1630_35242# 0.865968f
C3641 a_19862_44208# a_19511_42282# 1.12e-19
C3642 a_n443_42852# a_n2267_43396# 9.52e-20
C3643 a_12549_44172# a_15890_42674# 5.15e-21
C3644 a_2711_45572# a_19478_44056# 4.36e-19
C3645 a_n863_45724# a_4235_43370# 1.09e-20
C3646 a_13777_45326# a_13857_44734# 8.93e-19
C3647 a_9482_43914# a_14815_43914# 0.024524f
C3648 a_n2017_45002# a_3422_30871# 2.49e-20
C3649 a_n357_42282# a_1209_43370# 1.52e-19
C3650 a_n755_45592# a_458_43396# 0.001112f
C3651 a_3090_45724# a_11301_43218# 0.001286f
C3652 a_n1925_46634# a_4099_45572# 2.99e-20
C3653 a_n743_46660# a_2711_45572# 0.525746f
C3654 a_768_44030# a_8746_45002# 0.001081f
C3655 a_12549_44172# a_10490_45724# 0.00731f
C3656 a_765_45546# a_2324_44458# 5.17e-20
C3657 a_17339_46660# a_15682_46116# 2.86e-19
C3658 SMPL_ON_P a_n2661_45010# 0.006065f
C3659 a_n2497_47436# a_n1059_45260# 0.073215f
C3660 a_16327_47482# a_16223_45938# 0.016725f
C3661 a_2609_46660# a_3503_45724# 2.66e-19
C3662 a_2959_46660# a_3218_45724# 1.15e-19
C3663 a_n2661_46634# a_6667_45809# 5.79e-21
C3664 a_12891_46348# a_11322_45546# 1.18e-20
C3665 a_11309_47204# a_11525_45546# 0.004008f
C3666 a_376_46348# a_1176_45822# 0.001135f
C3667 a_n2293_46098# a_3147_46376# 1.09e-19
C3668 a_472_46348# a_1208_46090# 0.088629f
C3669 a_1239_47204# a_2437_43646# 4.55e-19
C3670 a_n881_46662# a_13904_45546# 9.09e-19
C3671 a_14513_46634# a_6945_45028# 3.51e-20
C3672 a_14035_46660# a_10809_44734# 0.00805f
C3673 a_10227_46804# a_16680_45572# 2.11e-19
C3674 a_n2293_42282# a_3581_42558# 0.001341f
C3675 a_1443_43940# VDD 0.144342f
C3676 a_13467_32519# a_22465_38105# 0.076379f
C3677 a_10341_42308# a_5742_30871# 0.031841f
C3678 a_13887_32519# a_21613_42308# 0.00157f
C3679 a_7499_43078# a_8605_42826# 0.026478f
C3680 a_n1925_42282# COMP_P 0.071512f
C3681 a_8199_44636# a_9803_42558# 0.036259f
C3682 a_8953_45546# a_8791_42308# 0.006945f
C3683 a_4185_45028# a_13070_42354# 8.35e-20
C3684 a_21101_45002# a_21115_43940# 3.47e-20
C3685 a_11827_44484# a_20623_43914# 0.004538f
C3686 a_15928_47570# VDD 0.08228f
C3687 a_12549_44172# START 8.3e-19
C3688 a_8128_46384# DATA[3] 1.73e-19
C3689 a_20193_45348# a_15493_43396# 3.33e-21
C3690 a_768_44030# RST_Z 0.05505f
C3691 a_n356_44636# a_644_44056# 2.5e-19
C3692 a_n2661_44458# a_10405_44172# 1.99e-20
C3693 a_11691_44458# a_19478_44306# 3.14e-20
C3694 a_18494_42460# a_15493_43940# 0.02195f
C3695 a_n881_46662# CLK 0.023376f
C3696 a_n357_42282# a_3059_42968# 7.39e-19
C3697 a_2711_45572# a_17701_42308# 5.54e-20
C3698 a_11189_46129# a_2711_45572# 0.011492f
C3699 a_5937_45572# a_6511_45714# 9.66e-19
C3700 a_8199_44636# a_6667_45809# 4.59e-21
C3701 a_4646_46812# a_6709_45028# 0.031325f
C3702 a_5732_46660# a_5691_45260# 9.85e-21
C3703 a_5907_46634# a_3232_43370# 1.41e-20
C3704 a_n971_45724# a_5891_43370# 0.084717f
C3705 a_17339_46660# a_16680_45572# 2.93e-21
C3706 a_n1545_46494# a_n2293_45546# 8.21e-20
C3707 a_8049_45260# a_11315_46155# 1.74e-19
C3708 a_n237_47217# a_7640_43914# 4.56e-21
C3709 a_4419_46090# a_4880_45572# 0.032829f
C3710 a_n881_46662# a_17023_45118# 2.61e-20
C3711 a_15227_44166# a_17668_45572# 2.59e-20
C3712 a_7927_46660# a_413_45260# 1.45e-20
C3713 a_n1151_42308# a_n1821_44484# 1.76e-19
C3714 a_5342_30871# C10_P_btm 2.16e-19
C3715 a_7227_42852# VDD 0.254613f
C3716 a_n3674_38216# a_n3420_38528# 0.152701f
C3717 a_5932_42308# a_n4315_30879# 6.05e-21
C3718 a_n4318_38216# a_n4064_38528# 0.057645f
C3719 a_5534_30871# C8_P_btm 5.29e-19
C3720 a_n4318_37592# a_n3565_38502# 3.09e-20
C3721 a_19721_31679# a_13467_32519# 0.051394f
C3722 a_13249_42308# a_13249_42558# 0.003175f
C3723 en_comp a_13291_42460# 4.34e-21
C3724 a_1138_42852# VDD 0.397518f
C3725 a_11823_42460# a_15486_42560# 0.003207f
C3726 a_5891_43370# a_8229_43396# 1.73e-20
C3727 a_10193_42453# a_11633_42308# 0.003739f
C3728 a_n1059_45260# a_17141_43172# 0.001223f
C3729 a_n2017_45002# a_18504_43218# 0.016191f
C3730 a_3422_30871# a_21845_43940# 4.36e-19
C3731 a_16112_44458# a_16137_43396# 2.27e-19
C3732 a_n2661_43922# a_7112_43396# 3.6e-21
C3733 a_n2661_42834# a_8147_43396# 1.43e-20
C3734 a_2998_44172# a_3737_43940# 0.003753f
C3735 a_15682_46116# a_1307_43914# 0.001505f
C3736 a_10193_42453# a_11962_45724# 0.044438f
C3737 a_2711_45572# a_11136_45572# 0.002612f
C3738 a_8746_45002# a_11652_45724# 2.41e-21
C3739 a_10809_44734# a_10951_45334# 0.015679f
C3740 a_10490_45724# a_11525_45546# 0.06936f
C3741 a_526_44458# a_4558_45348# 7.28e-20
C3742 a_12741_44636# a_18494_42460# 0.114105f
C3743 a_11415_45002# a_21101_45002# 0.018873f
C3744 a_768_44030# a_5663_43940# 0.011502f
C3745 a_20202_43084# a_21359_45002# 0.008822f
C3746 a_n1613_43370# a_n1441_43940# 0.012196f
C3747 a_16327_47482# a_11341_43940# 0.063063f
C3748 a_8270_45546# a_7640_43914# 2.57e-20
C3749 a_15227_44166# a_17970_44736# 0.002254f
C3750 a_3483_46348# a_7735_45067# 2.41e-19
C3751 a_2698_46116# a_n2661_43370# 1.36e-20
C3752 a_n1925_42282# a_4574_45260# 3.52e-19
C3753 a_n2109_47186# a_383_46660# 2.96e-20
C3754 a_n1741_47186# a_33_46660# 4.45e-20
C3755 a_n971_45724# a_n1021_46688# 0.002801f
C3756 a_n746_45260# a_n1925_46634# 0.036469f
C3757 a_21177_47436# a_12465_44636# 2.23e-19
C3758 a_19386_47436# a_11453_44696# 1.38e-19
C3759 a_2113_38308# VDAC_Pi 0.170908f
C3760 a_n3565_38502# a_n4334_37440# 4.13e-19
C3761 a_n4209_38502# a_n3690_37440# 3.34e-19
C3762 a_n4209_39304# VDAC_P 4.55e-19
C3763 a_1239_47204# a_n2661_46634# 0.002062f
C3764 a_6151_47436# a_13569_47204# 0.004336f
C3765 a_21496_47436# a_4883_46098# 0.257837f
C3766 a_13507_46334# a_21811_47423# 4.35e-19
C3767 a_9863_47436# a_10037_47542# 0.006584f
C3768 a_9313_45822# a_8128_46384# 0.013269f
C3769 a_13717_47436# a_n881_46662# 0.039579f
C3770 a_4958_30871# C1_N_btm 9.46e-20
C3771 a_n815_47178# a_n2438_43548# 1.87e-19
C3772 a_n452_47436# a_n743_46660# 6.22e-21
C3773 a_19478_44306# a_4190_30871# 2.22e-20
C3774 a_5663_43940# a_5755_42852# 0.001147f
C3775 a_n2661_42282# a_n1641_43230# 1.25e-20
C3776 a_20512_43084# a_18083_42858# 1.67e-21
C3777 a_5883_43914# a_1755_42282# 2.89e-20
C3778 a_11962_45724# VDD 0.210594f
C3779 a_4699_43561# a_2982_43646# 1.91e-20
C3780 a_4093_43548# a_3626_43646# 0.011002f
C3781 a_458_43396# a_548_43396# 0.008441f
C3782 a_n97_42460# a_7287_43370# 0.004081f
C3783 a_14021_43940# a_17324_43396# 0.009103f
C3784 a_19862_44208# a_21259_43561# 8.37e-19
C3785 a_n2956_37592# a_n3420_37984# 0.001223f
C3786 a_n699_43396# a_2903_42308# 1.29e-19
C3787 a_3422_30871# a_19164_43230# 5.64e-20
C3788 a_9049_44484# DATA[4] 1.59e-19
C3789 a_15493_43396# a_20301_43646# 2.14e-19
C3790 a_17737_43940# a_4361_42308# 1.14e-20
C3791 a_12549_44172# a_16547_43609# 4.68e-19
C3792 a_3218_45724# a_n699_43396# 1.28e-20
C3793 a_16855_45546# a_16751_45260# 4.68e-19
C3794 a_15861_45028# a_15595_45028# 0.072432f
C3795 a_8696_44636# a_16019_45002# 2.28e-19
C3796 a_3090_45724# a_6671_43940# 0.00493f
C3797 a_3357_43084# a_n913_45002# 2.04e-19
C3798 a_18597_46090# a_20749_43396# 0.005121f
C3799 a_1823_45246# a_5013_44260# 0.001797f
C3800 a_13507_46334# a_22223_43396# 0.006729f
C3801 a_20075_46420# a_20159_44458# 1.46e-19
C3802 a_n2293_46634# a_9803_43646# 0.01299f
C3803 C2_N_btm VREF_GND 0.671742f
C3804 C1_N_btm VCM 0.716121f
C3805 VDD DATA[1] 0.321585f
C3806 C4_N_btm VIN_N 0.50261f
C3807 C3_N_btm VREF 0.984942f
C3808 a_13507_46334# a_22000_46634# 0.183978f
C3809 a_20990_47178# a_20731_47026# 6.38e-19
C3810 a_21496_47436# a_21188_46660# 2.45e-19
C3811 a_10227_46804# a_20719_46660# 3.17e-19
C3812 a_n1741_47186# a_12005_46116# 0.174477f
C3813 a_2063_45854# a_6419_46155# 1.49e-19
C3814 a_3160_47472# a_5164_46348# 9.48e-21
C3815 a_n1151_42308# a_5068_46348# 0.089946f
C3816 a_12465_44636# a_20841_46902# 3.04e-20
C3817 a_18597_46090# a_18280_46660# 3.97e-19
C3818 a_3877_44458# a_6540_46812# 0.244975f
C3819 a_4646_46812# a_5732_46660# 0.050752f
C3820 a_4651_46660# a_5907_46634# 0.043482f
C3821 a_n1925_46634# a_8189_46660# 1.2e-19
C3822 a_5807_45002# a_15368_46634# 0.029781f
C3823 a_12891_46348# a_12359_47026# 0.002172f
C3824 a_3785_47178# a_4419_46090# 2.07e-20
C3825 a_n443_46116# a_2804_46116# 0.018109f
C3826 a_n1435_47204# a_n1853_46287# 2.54e-20
C3827 a_n881_46662# a_14035_46660# 9.06e-20
C3828 a_4883_46098# a_21363_46634# 0.066909f
C3829 a_11453_44696# a_19551_46910# 0.047386f
C3830 a_13661_43548# a_14976_45028# 0.162789f
C3831 a_13747_46662# a_3090_45724# 0.139869f
C3832 a_n2661_46634# a_11186_47026# 0.002094f
C3833 a_n237_47217# a_9823_46155# 4.34e-20
C3834 a_2107_46812# a_6969_46634# 2.09e-19
C3835 a_4955_46873# a_5167_46660# 0.003269f
C3836 a_4817_46660# a_5385_46902# 0.170485f
C3837 a_14579_43548# a_14543_43071# 0.032593f
C3838 a_14205_43396# a_13635_43156# 0.002342f
C3839 a_21855_43396# a_22223_43396# 7.52e-19
C3840 a_743_42282# a_20749_43396# 0.09037f
C3841 a_11361_45348# CLK 3.72e-20
C3842 a_4905_42826# a_4649_42852# 0.006342f
C3843 a_13678_32519# a_5649_42852# 0.506367f
C3844 a_13467_32519# a_22591_43396# 4.5e-22
C3845 a_4361_42308# a_13887_32519# 2.22e-19
C3846 a_13807_45067# VDD 2.18e-20
C3847 a_6171_45002# a_13720_44458# 3.19e-20
C3848 a_n967_45348# a_n998_44484# 0.001023f
C3849 a_20447_31679# a_9313_44734# 1.21e-20
C3850 a_3090_45724# a_10796_42968# 0.004117f
C3851 a_n37_45144# a_n356_44636# 4.09e-19
C3852 a_n143_45144# a_n23_44458# 0.001215f
C3853 a_2324_44458# a_6452_43396# 1.62e-20
C3854 a_8953_45002# a_10157_44484# 0.002321f
C3855 a_n1925_42282# a_1568_43370# 1.62e-21
C3856 a_526_44458# a_1756_43548# 0.01292f
C3857 a_22612_30879# a_14097_32519# 0.059759f
C3858 a_2107_46812# a_9241_46436# 2.55e-19
C3859 a_n743_46660# a_10037_46155# 3.34e-19
C3860 a_6755_46942# a_14275_46494# 1.11e-19
C3861 a_10623_46897# a_2324_44458# 1.46e-20
C3862 a_8270_45546# a_9823_46155# 3.17e-19
C3863 a_n881_46662# a_n1099_45572# 0.088565f
C3864 a_n1613_43370# a_310_45028# 1.46e-20
C3865 a_21363_46634# a_21188_46660# 0.233657f
C3866 a_18285_46348# a_18900_46660# 0.004259f
C3867 a_20273_46660# a_20731_47026# 0.027606f
C3868 a_19123_46287# a_18280_46660# 8.18e-20
C3869 a_5807_45002# a_19597_46482# 1.86e-20
C3870 a_6151_47436# a_11823_42460# 4.56e-21
C3871 a_9313_45822# a_10053_45546# 4.44e-20
C3872 a_3090_45724# a_4419_46090# 0.001764f
C3873 a_2063_45854# a_10907_45822# 0.22153f
C3874 a_15781_43660# a_16104_42674# 4.99e-20
C3875 a_3080_42308# comp_n 2.82e-19
C3876 a_n4318_39768# VDD 0.469044f
C3877 a_17595_43084# a_17665_42852# 0.011552f
C3878 a_5649_42852# a_6123_31319# 0.062309f
C3879 a_4361_42308# a_8515_42308# 0.007572f
C3880 a_743_42282# a_8685_42308# 0.039566f
C3881 a_1138_42852# a_n784_42308# 3.74e-20
C3882 a_n863_45724# a_791_42968# 0.338631f
C3883 a_n2661_45546# a_3935_42891# 1.6e-19
C3884 a_13259_45724# a_12545_42858# 3.09e-19
C3885 a_14537_43396# a_11341_43940# 0.032289f
C3886 a_13720_44458# a_14673_44172# 2.95e-20
C3887 a_n2293_42834# a_3499_42826# 0.029158f
C3888 a_2711_45572# a_4361_42308# 0.031943f
C3889 a_526_44458# a_5193_43172# 3.3e-19
C3890 a_11823_42460# a_13837_43396# 0.001813f
C3891 a_10193_42453# a_17499_43370# 0.009503f
C3892 a_8696_44636# a_8791_43396# 3.5e-20
C3893 a_6151_47436# DATA[3] 0.041263f
C3894 a_9863_47436# VDD 0.207794f
C3895 a_5891_43370# a_9313_44734# 0.028253f
C3896 a_9482_43914# a_9248_44260# 5.36e-21
C3897 a_11813_46116# a_11682_45822# 2.39e-19
C3898 a_n2956_39768# en_comp 0.003442f
C3899 a_n2312_38680# a_n2017_45002# 8.38e-22
C3900 a_14275_46494# a_8049_45260# 0.001971f
C3901 a_11387_46155# a_11608_46482# 0.007833f
C3902 a_n2293_46098# a_310_45028# 0.017313f
C3903 a_n2157_46122# a_n1099_45572# 1.52e-19
C3904 a_12549_44172# a_6171_45002# 0.029809f
C3905 a_472_46348# a_n2661_45546# 2.09e-20
C3906 a_19594_46812# a_413_45260# 4.71e-20
C3907 a_768_44030# a_3232_43370# 0.224083f
C3908 a_6755_46942# a_15765_45572# 0.026052f
C3909 a_2107_46812# a_3357_43084# 0.033995f
C3910 a_n2293_46634# a_n913_45002# 0.024406f
C3911 a_n2438_43548# a_n2661_45010# 0.220364f
C3912 a_15368_46634# a_15143_45578# 0.105334f
C3913 a_n901_46420# a_n2293_45546# 1.79e-20
C3914 a_6761_42308# a_8515_42308# 1.96e-20
C3915 a_7227_42308# a_5934_30871# 5.66e-20
C3916 a_17499_43370# VDD 0.453381f
C3917 a_3318_42354# a_5742_30871# 1.46e-20
C3918 a_6123_31319# a_7963_42308# 0.192155f
C3919 a_4190_30871# C8_P_btm 4.06e-19
C3920 a_3232_43370# a_5755_42852# 5.23e-21
C3921 a_n357_42282# a_14456_42282# 7.69e-20
C3922 a_20835_44721# a_11341_43940# 6.34e-20
C3923 a_20766_44850# a_21115_43940# 4.08e-19
C3924 a_20640_44752# a_15493_43940# 7.7e-20
C3925 a_18579_44172# a_20269_44172# 7.35e-20
C3926 a_19279_43940# a_20935_43940# 2.95e-19
C3927 a_20820_30879# a_22521_39511# 5.7e-20
C3928 a_n2017_45002# a_16414_43172# 2.51e-19
C3929 a_13259_45724# a_19332_42282# 1.03e-19
C3930 a_n2661_42834# a_10555_43940# 8.1e-20
C3931 a_21076_30879# a_22521_40055# 2.11e-20
C3932 a_4223_44672# a_6197_43396# 1.94e-19
C3933 a_5111_44636# a_7765_42852# 3.95e-20
C3934 a_n443_42852# a_9223_42460# 1.18e-20
C3935 a_n913_45002# a_5342_30871# 0.122483f
C3936 a_n1059_45260# a_15567_42826# 0.048229f
C3937 a_6453_43914# a_7542_44172# 2.4e-20
C3938 a_1414_42308# a_2253_44260# 0.001444f
C3939 a_12978_47026# VDD 7.19e-19
C3940 a_n23_44458# a_n97_42460# 4.48e-19
C3941 a_n356_44636# a_104_43370# 0.001131f
C3942 a_11691_44458# a_13667_43396# 3.82e-21
C3943 a_21137_46414# a_20107_45572# 0.002164f
C3944 a_20708_46348# a_20273_45572# 4.47e-20
C3945 a_14840_46494# a_2437_43646# 1.19e-36
C3946 a_3316_45546# a_3260_45572# 4.85e-19
C3947 a_11415_45002# a_14797_45144# 0.021281f
C3948 a_12741_44636# a_13777_45326# 4.48e-20
C3949 a_13507_46334# a_20512_43084# 0.497215f
C3950 a_4185_45028# a_2382_45260# 0.008734f
C3951 a_3090_45724# a_18911_45144# 0.190188f
C3952 a_3483_46348# a_3065_45002# 0.001025f
C3953 a_3147_46376# a_3429_45260# 1.69e-19
C3954 a_12549_44172# a_14673_44172# 0.024138f
C3955 a_8049_45260# a_15765_45572# 0.012841f
C3956 a_13661_43548# a_15433_44458# 0.038412f
C3957 a_5257_43370# a_5518_44484# 0.095452f
C3958 a_n3565_39590# a_n4209_38216# 0.0313f
C3959 a_n4209_39304# a_n4334_38528# 6.38e-20
C3960 a_n4334_39392# a_n4209_38502# 6.38e-20
C3961 a_n4209_39590# a_n3565_38216# 0.03183f
C3962 a_1606_42308# C7_N_btm 0.00238f
C3963 a_n1151_42308# a_15811_47375# 1.38e-21
C3964 a_4915_47217# a_n1435_47204# 0.038318f
C3965 a_7227_47204# a_6575_47204# 0.028925f
C3966 a_6151_47436# a_9313_45822# 0.032544f
C3967 a_5934_30871# a_n923_35174# 0.009397f
C3968 a_1576_42282# VDD 0.26017f
C3969 a_n4064_40160# a_n4064_37984# 0.067467f
C3970 a_n3420_39072# a_n2860_39072# 0.003211f
C3971 a_20512_43084# a_21855_43396# 0.013929f
C3972 a_9313_44734# a_17595_43084# 0.006038f
C3973 a_21205_44306# a_21381_43940# 8.17e-20
C3974 a_10405_44172# a_9145_43396# 1.63e-19
C3975 a_n913_45002# a_20107_42308# 3.57e-19
C3976 a_n2293_43922# a_12089_42308# 0.183316f
C3977 a_13483_43940# a_8685_43396# 2.97e-20
C3978 a_n2956_38216# VDD 0.484692f
C3979 a_3422_30871# a_14209_32519# 0.031148f
C3980 a_n2293_42834# a_3318_42354# 4.09e-21
C3981 a_n2017_45002# a_7174_31319# 2.34e-19
C3982 a_12861_44030# a_14537_43646# 1.95e-20
C3983 a_n443_42852# a_117_45144# 6.39e-19
C3984 a_20202_43084# a_19279_43940# 0.020761f
C3985 a_11415_45002# a_20766_44850# 0.001727f
C3986 a_18341_45572# a_18596_45572# 0.056391f
C3987 a_18909_45814# a_19256_45572# 0.051162f
C3988 a_5263_45724# a_1423_45028# 5.02e-21
C3989 a_5066_45546# a_4223_44672# 2.22e-20
C3990 a_9290_44172# a_9313_44734# 0.140741f
C3991 a_768_44030# a_4905_42826# 4.03e-20
C3992 a_11652_45724# a_3232_43370# 0.009948f
C3993 a_n1613_43370# a_n998_43396# 0.001965f
C3994 a_10227_46804# a_14358_43442# 0.019948f
C3995 a_526_44458# a_9838_44484# 1.68e-22
C3996 a_380_45546# a_n2661_43370# 4.07e-20
C3997 a_16327_47482# a_10341_43396# 0.159266f
C3998 a_11525_45546# a_6171_45002# 9.43e-19
C3999 a_1239_47204# a_765_45546# 9.93e-19
C4000 a_n1613_43370# a_5894_47026# 5.16e-19
C4001 EN_VIN_BSTR_P a_n83_35174# 0.652984f
C4002 VDAC_N C8_N_btm 61.723f
C4003 a_11599_46634# a_3090_45724# 0.133107f
C4004 a_n2293_46634# a_2107_46812# 3.61e-19
C4005 a_n743_46660# a_33_46660# 0.025563f
C4006 a_n2438_43548# a_171_46873# 0.029723f
C4007 a_n4209_37414# VIN_P 0.029528f
C4008 a_4915_47217# a_13885_46660# 0.179458f
C4009 a_n1151_42308# a_13059_46348# 0.003065f
C4010 a_12861_44030# a_16292_46812# 0.059827f
C4011 a_n1925_46634# a_383_46660# 0.009919f
C4012 a_3726_37500# RST_Z 1.60318f
C4013 a_n2661_46634# a_491_47026# 0.003523f
C4014 a_15811_47375# a_14084_46812# 7.3e-20
C4015 a_10227_46804# a_11735_46660# 0.54163f
C4016 a_4338_37500# VDD 0.525635f
C4017 a_9313_44734# a_21887_42336# 0.001765f
C4018 a_7229_43940# VDD 0.821851f
C4019 a_19319_43548# a_19339_43156# 0.006943f
C4020 a_2982_43646# a_1847_42826# 4.13e-21
C4021 a_15681_43442# a_15743_43084# 0.001131f
C4022 a_10341_43396# a_16855_43396# 8.56e-19
C4023 a_n97_42460# a_12089_42308# 4.02e-19
C4024 a_16547_43609# a_16977_43638# 6.72e-20
C4025 a_16137_43396# a_17499_43370# 1.55e-19
C4026 a_16243_43396# a_16759_43396# 0.106647f
C4027 a_10907_45822# a_n2661_42834# 7.86e-20
C4028 a_n863_45724# a_3905_42865# 1.11e-19
C4029 a_4646_46812# a_7227_42852# 0.032378f
C4030 a_n1613_43370# a_8495_42852# 0.012196f
C4031 a_10775_45002# a_n2661_43370# 0.009126f
C4032 a_n443_42852# a_n2065_43946# 5.59e-21
C4033 a_2957_45546# a_1414_42308# 9.39e-21
C4034 a_16147_45260# a_16979_44734# 6.23e-20
C4035 a_20447_31679# a_18114_32519# 0.051474f
C4036 a_n443_46116# a_1755_42282# 3.6e-20
C4037 a_16327_47482# a_20356_42852# 7.6e-21
C4038 a_3357_43084# a_n2661_44458# 0.027126f
C4039 a_22959_45572# a_19721_31679# 0.005929f
C4040 a_n357_42282# a_895_43940# 0.008143f
C4041 a_n755_45592# a_2479_44172# 1.32e-20
C4042 a_1823_45246# a_4699_43561# 0.003517f
C4043 a_11823_42460# a_12829_44484# 2.31e-19
C4044 a_3877_44458# a_1823_45246# 0.231164f
C4045 a_14084_46812# a_13059_46348# 5.17e-19
C4046 a_15009_46634# a_15227_46910# 0.08213f
C4047 a_2905_45572# a_3503_45724# 0.001385f
C4048 a_n1151_42308# a_3218_45724# 5.24e-20
C4049 a_3160_47472# a_3316_45546# 0.003495f
C4050 a_n443_46116# a_n1099_45572# 0.368941f
C4051 a_11186_47026# a_765_45546# 5.79e-19
C4052 a_19321_45002# a_19553_46090# 0.008717f
C4053 a_19594_46812# a_18985_46122# 9.08e-20
C4054 a_n743_46660# a_12005_46116# 0.024033f
C4055 a_13747_46662# a_20075_46420# 1.64e-20
C4056 a_16942_47570# a_6945_45028# 1.33e-19
C4057 a_5807_45002# a_20708_46348# 1.89e-19
C4058 a_n881_46662# a_n1925_42282# 0.041426f
C4059 a_15559_46634# a_14513_46634# 2.81e-20
C4060 a_2107_46812# a_9625_46129# 0.184645f
C4061 a_11599_46634# a_15002_46116# 4.2e-19
C4062 a_10227_46804# a_14537_46482# 0.001903f
C4063 a_4883_46098# a_11387_46482# 2.91e-19
C4064 a_18204_44850# VDD 4.6e-19
C4065 a_17517_44484# RST_Z 0.004664f
C4066 a_20974_43370# a_21887_42336# 8.61e-21
C4067 a_18083_42858# a_18249_42858# 0.699797f
C4068 a_2982_43646# a_15486_42560# 9.69e-20
C4069 a_3626_43646# a_14113_42308# 0.077829f
C4070 a_7227_42852# a_7309_43172# 0.003935f
C4071 a_3935_42891# a_3863_42891# 6.64e-19
C4072 a_n452_44636# a_n310_44811# 0.005572f
C4073 a_5205_44484# a_6453_43914# 7.72e-19
C4074 a_7229_43940# a_5495_43940# 6.48e-21
C4075 a_n443_42852# a_13667_43396# 0.035517f
C4076 a_949_44458# a_n356_44636# 0.009584f
C4077 a_11827_44484# a_11649_44734# 5.76e-21
C4078 a_526_44458# a_421_43172# 3.36e-20
C4079 a_12883_44458# a_13076_44458# 0.142643f
C4080 a_12607_44458# a_13720_44458# 0.122704f
C4081 a_n2442_46660# a_n4064_40160# 0.006941f
C4082 a_n1059_45260# a_10405_44172# 2.46e-20
C4083 a_413_45260# a_3499_42826# 4.69e-19
C4084 a_n2661_44458# a_5826_44734# 6.36e-19
C4085 a_375_42282# a_n2065_43946# 2.58e-21
C4086 a_7499_43078# a_3626_43646# 0.002457f
C4087 a_6545_47178# a_6709_45028# 1.46e-20
C4088 a_10227_46804# en_comp 2.31e-20
C4089 a_9290_44172# a_12594_46348# 1.22e-21
C4090 a_n237_47217# a_1423_45028# 5.23e-20
C4091 a_376_46348# a_518_46482# 0.007833f
C4092 a_15673_47210# a_413_45260# 2.52e-19
C4093 a_11189_46129# a_12005_46116# 0.00104f
C4094 a_11133_46155# a_10903_43370# 2.09e-20
C4095 a_2107_46812# a_9159_45572# 6.31e-20
C4096 a_3090_45724# a_1848_45724# 3.59e-19
C4097 a_16388_46812# a_16375_45002# 0.039999f
C4098 a_n971_45724# a_2304_45348# 0.00123f
C4099 a_18597_46090# a_n913_45002# 0.126328f
C4100 a_11453_44696# a_3357_43084# 0.020072f
C4101 a_21356_42826# a_13258_32519# 6.82e-21
C4102 COMP_P a_1606_42308# 2.6775f
C4103 a_n4318_38680# a_n2860_38778# 1.77e-20
C4104 a_196_42282# a_1184_42692# 2.75e-19
C4105 a_n784_42308# a_1576_42282# 0.038241f
C4106 a_n473_42460# a_961_42354# 2.64e-21
C4107 a_n3674_37592# a_n1630_35242# 0.096752f
C4108 a_19164_43230# a_7174_31319# 3.33e-21
C4109 a_10752_42852# a_5742_30871# 5.4e-20
C4110 a_n2661_42834# a_n2661_42282# 0.019795f
C4111 a_3877_44458# DATA[2] 0.001477f
C4112 a_5907_46634# VDD 0.341121f
C4113 a_9313_44734# a_10807_43548# 0.033005f
C4114 a_22315_44484# a_22591_44484# 0.001038f
C4115 a_3422_30871# a_17730_32519# 0.004485f
C4116 a_n2293_42834# a_6197_43396# 1.31e-19
C4117 a_n913_45002# a_743_42282# 0.25834f
C4118 a_7499_43078# a_8649_43218# 5.01e-19
C4119 a_14537_43396# a_10341_43396# 0.013753f
C4120 a_1307_43914# a_14358_43442# 1.45e-20
C4121 a_20447_31679# a_13887_32519# 0.051465f
C4122 a_19963_31679# a_14209_32519# 0.051256f
C4123 a_10809_44734# a_13527_45546# 3.56e-21
C4124 a_8049_45260# a_6194_45824# 4.11e-20
C4125 a_768_44030# a_8975_43940# 0.124155f
C4126 a_n2840_45546# a_n2661_45546# 0.175179f
C4127 a_11415_45002# a_19365_45572# 1.55e-19
C4128 a_7411_46660# a_8560_45348# 2.42e-21
C4129 a_8270_45546# a_1423_45028# 0.023554f
C4130 a_10903_43370# a_11688_45572# 2.55e-20
C4131 a_n2293_46634# a_n2661_44458# 0.029279f
C4132 a_13607_46688# a_13777_45326# 2.78e-21
C4133 a_3483_46348# a_14033_45572# 0.003201f
C4134 a_16388_46812# a_413_45260# 4.56e-20
C4135 a_12549_44172# a_12607_44458# 0.033279f
C4136 a_12891_46348# a_12883_44458# 0.018059f
C4137 a_5807_45002# a_5518_44484# 7.14e-20
C4138 a_10227_46804# a_10617_44484# 0.006757f
C4139 a_n2497_47436# a_n237_47217# 4.7e-20
C4140 SMPL_ON_P a_n1605_47204# 0.194856f
C4141 a_n1741_47186# a_n815_47178# 0.031488f
C4142 a_n2109_47186# a_n971_45724# 1.21934f
C4143 a_21613_42308# a_21421_42336# 5.76e-19
C4144 a_4649_42852# VDD 0.194775f
C4145 a_18451_43940# a_18533_44260# 0.003935f
C4146 a_20835_44721# a_10341_43396# 2.07e-20
C4147 a_3600_43914# a_3626_43646# 3.68e-19
C4148 a_3537_45260# a_1755_42282# 0.002095f
C4149 a_n1059_45260# a_6171_42473# 2.78e-20
C4150 a_n2017_45002# a_5932_42308# 0.005049f
C4151 a_n913_45002# a_5755_42308# 0.036226f
C4152 a_10809_44734# EN_OFFSET_CAL 0.035912f
C4153 a_20193_45348# a_21356_42826# 1.21e-20
C4154 a_5883_43914# a_8387_43230# 2.5e-20
C4155 a_9313_44734# a_13467_32519# 0.057668f
C4156 a_5841_44260# a_n97_42460# 6.63e-22
C4157 a_17973_43940# a_19319_43548# 2.01e-22
C4158 a_6511_45714# a_2437_43646# 2.64e-21
C4159 a_16327_47482# a_n97_42460# 0.113034f
C4160 a_13259_45724# a_14797_45144# 0.092924f
C4161 a_526_44458# a_n2661_43370# 0.054473f
C4162 a_5066_45546# a_n2293_42834# 3.17e-20
C4163 a_17583_46090# a_11827_44484# 6.39e-21
C4164 a_n356_45724# a_n143_45144# 3.1e-21
C4165 a_n357_42282# a_3065_45002# 0.023226f
C4166 a_3316_45546# a_413_45260# 0.110075f
C4167 a_n755_45592# a_2680_45002# 5.6e-20
C4168 a_n743_46660# a_15682_43940# 0.001683f
C4169 a_13507_46334# a_21381_43940# 5.15e-20
C4170 a_19335_46494# a_19778_44110# 4.32e-19
C4171 a_3483_46348# a_6298_44484# 0.017162f
C4172 a_2107_46812# a_9672_43914# 0.079349f
C4173 a_5907_45546# a_3357_43084# 0.023698f
C4174 a_15015_46420# a_11691_44458# 4.75e-21
C4175 a_5068_46348# a_4223_44672# 1.13e-20
C4176 a_4419_46090# a_4743_44484# 8.99e-21
C4177 a_4185_45028# a_5343_44458# 5.81e-20
C4178 a_n1013_45572# a_n967_45348# 2.46e-19
C4179 a_12549_44172# a_14761_44260# 1.08e-19
C4180 a_19321_45002# a_15493_43940# 0.050579f
C4181 a_n2312_39304# a_n2661_46634# 0.105298f
C4182 a_n2312_40392# a_n2472_46634# 3.86e-20
C4183 a_n4209_38216# C4_P_btm 0.001041f
C4184 a_n3565_38216# C6_P_btm 1.26e-20
C4185 a_8530_39574# CAL_N 0.644218f
C4186 a_6545_47178# a_5732_46660# 1.97e-20
C4187 a_6151_47436# a_6540_46812# 0.043688f
C4188 a_6491_46660# a_5907_46634# 0.002903f
C4189 a_11309_47204# a_12891_46348# 9.04e-21
C4190 a_1736_39043# VDD 2.8939f
C4191 a_2063_45854# a_9863_46634# 0.10786f
C4192 a_n1151_42308# a_7577_46660# 0.001579f
C4193 a_18596_45572# VDD 0.077608f
C4194 a_20974_43370# a_13467_32519# 0.017399f
C4195 a_14401_32519# a_4361_42308# 8.07e-20
C4196 a_n2293_43922# a_5267_42460# 4.38e-20
C4197 a_n356_44636# a_10723_42308# 2.77e-19
C4198 a_14539_43914# a_15486_42560# 4.81e-21
C4199 a_11341_43940# a_12379_42858# 2.86e-20
C4200 a_10555_44260# a_10083_42826# 9.41e-22
C4201 a_20447_31679# EN_VIN_BSTR_N 0.002888f
C4202 a_17737_43940# a_17595_43084# 8.42e-21
C4203 a_n2661_42282# a_n2293_42282# 1.04835f
C4204 a_5891_43370# a_8515_42308# 1.03e-19
C4205 a_n97_42460# a_16855_43396# 8.47e-19
C4206 a_16147_45260# a_16321_45348# 0.002641f
C4207 a_18597_46090# a_20922_43172# 0.021228f
C4208 a_11652_45724# a_8975_43940# 1.25e-20
C4209 a_8696_44636# a_11827_44484# 0.039f
C4210 a_3357_43084# a_6125_45348# 0.001261f
C4211 a_2063_45854# a_11136_42852# 2.55e-20
C4212 a_2711_45572# a_5891_43370# 8.73e-21
C4213 a_526_44458# a_2998_44172# 0.028337f
C4214 a_15227_44166# a_3626_43646# 1.37e-19
C4215 a_n913_45002# a_626_44172# 7.19e-20
C4216 a_10903_43370# a_12429_44172# 0.116356f
C4217 a_13507_46334# a_18249_42858# 5.85e-19
C4218 a_6171_45002# a_5205_44484# 0.0168f
C4219 a_5691_45260# a_7229_43940# 2.13e-20
C4220 a_3232_43370# a_7276_45260# 0.027376f
C4221 a_16333_45814# a_11691_44458# 3.71e-21
C4222 a_n1613_43370# a_9127_43156# 0.267842f
C4223 a_768_44030# a_2905_42968# 4.25e-19
C4224 a_n2956_39768# a_n2157_42858# 3.98e-21
C4225 a_11599_46634# a_20075_46420# 0.021805f
C4226 a_2063_45854# a_5527_46155# 8.53e-21
C4227 a_10428_46928# a_11813_46116# 1.23e-19
C4228 a_10467_46802# a_11735_46660# 0.096658f
C4229 a_10554_47026# a_10768_47026# 0.097745f
C4230 a_10623_46897# a_11186_47026# 0.049827f
C4231 a_6755_46942# a_8601_46660# 5.59e-19
C4232 a_n881_46662# a_2698_46116# 0.058407f
C4233 a_12465_44636# a_9290_44172# 7.82e-20
C4234 a_13507_46334# a_10903_43370# 0.016027f
C4235 a_16327_47482# a_17957_46116# 6.07e-20
C4236 a_n1151_42308# a_5431_46482# 0.004507f
C4237 a_3160_47472# a_5066_45546# 1.83e-20
C4238 a_491_47026# a_765_45546# 1.57e-19
C4239 a_19321_45002# a_12741_44636# 0.113088f
C4240 a_21588_30879# a_22365_46825# 5.32e-19
C4241 a_12861_44030# a_6945_45028# 0.108969f
C4242 a_n1435_47204# a_10809_44734# 9.93e-19
C4243 a_20916_46384# a_20202_43084# 0.181561f
C4244 a_n443_46116# a_n1925_42282# 0.001452f
C4245 a_10227_46804# a_2324_44458# 0.051051f
C4246 a_4883_46098# a_11133_46155# 0.007956f
C4247 a_5649_42852# a_18083_42858# 4.21e-20
C4248 a_4190_30871# a_21195_42852# 1.06e-20
C4249 a_15493_43940# a_17531_42308# 1.35e-21
C4250 a_n1557_42282# a_564_42282# 0.003471f
C4251 a_15004_44636# VDD 0.090175f
C4252 a_3935_42891# a_4520_42826# 0.017436f
C4253 a_4361_42308# a_18817_42826# 1.3e-20
C4254 a_14579_43548# a_13291_42460# 0.007999f
C4255 a_11341_43940# a_18727_42674# 3.06e-21
C4256 a_1568_43370# a_1606_42308# 0.007194f
C4257 a_3080_42308# a_1576_42282# 1.7e-20
C4258 a_n3674_39768# a_n3420_39072# 2.58e-20
C4259 a_17715_44484# a_16823_43084# 4.72e-20
C4260 a_n443_42852# a_n2129_43609# 1.4e-19
C4261 a_1823_45246# a_1847_42826# 1.28e-20
C4262 a_12549_44172# a_15959_42545# 2.73e-19
C4263 a_2711_45572# a_18533_43940# 0.004398f
C4264 a_n863_45724# a_4093_43548# 9.16e-21
C4265 a_13556_45296# a_13857_44734# 0.01375f
C4266 a_9482_43914# a_14112_44734# 0.004038f
C4267 a_19963_31679# a_17730_32519# 0.054244f
C4268 a_n357_42282# a_458_43396# 0.016095f
C4269 a_n755_45592# a_n229_43646# 0.049717f
C4270 a_626_44172# a_556_44484# 0.00387f
C4271 a_n2810_45572# a_n1557_42282# 1.35e-20
C4272 a_3090_45724# a_11229_43218# 7.17e-19
C4273 a_2107_46812# a_2277_45546# 4.99e-20
C4274 a_n2438_43548# a_1260_45572# 0.001032f
C4275 a_768_44030# a_10193_42453# 0.030504f
C4276 a_n2497_47436# a_n2017_45002# 0.125552f
C4277 SMPL_ON_P a_n2840_45002# 7.52e-19
C4278 a_16327_47482# a_16020_45572# 0.001041f
C4279 a_2959_46660# a_2957_45546# 1.67e-20
C4280 a_2443_46660# a_3503_45724# 3.68e-20
C4281 a_n2661_46634# a_6511_45714# 1.3e-20
C4282 a_5807_45002# a_6428_45938# 3.09e-19
C4283 a_11309_47204# a_11322_45546# 2.89e-19
C4284 a_376_46348# a_1208_46090# 5.21e-19
C4285 a_n2293_46098# a_2804_46116# 1.46e-20
C4286 a_472_46348# a_805_46414# 0.360492f
C4287 a_n881_46662# a_13527_45546# 1.35e-19
C4288 a_1209_47178# a_2437_43646# 0.025116f
C4289 a_16388_46812# a_18985_46122# 5.62e-21
C4290 a_14180_46812# a_6945_45028# 4.2e-20
C4291 a_13885_46660# a_10809_44734# 0.026009f
C4292 a_288_46660# a_n443_42852# 2.55e-21
C4293 a_n2293_42282# a_3497_42558# 0.001879f
C4294 a_1241_43940# VDD 0.162129f
C4295 a_13467_32519# a_22397_42558# 5.38e-19
C4296 a_4361_42308# a_21421_42336# 6.95e-19
C4297 a_10922_42852# a_5742_30871# 7.65e-19
C4298 a_12089_42308# a_10533_42308# 8.19e-21
C4299 a_10341_42308# a_11323_42473# 1.11e-19
C4300 a_n2661_44458# a_9672_43914# 4.07e-20
C4301 a_7499_43078# a_8037_42858# 0.160087f
C4302 a_5111_44636# a_2982_43646# 1.32e-19
C4303 a_15433_44458# a_11967_42832# 7e-22
C4304 a_9313_44734# a_22315_44484# 2.17e-21
C4305 a_n1925_42282# a_n4318_37592# 0.024213f
C4306 a_8953_45546# a_8685_42308# 0.250058f
C4307 a_8199_44636# a_9223_42460# 0.065156f
C4308 a_4185_45028# a_12563_42308# 1.64e-19
C4309 a_21101_45002# a_20935_43940# 0.001207f
C4310 a_11827_44484# a_20365_43914# 0.0059f
C4311 a_768_44030# VDD 1.53454f
C4312 a_4574_45260# a_3539_42460# 5.02e-22
C4313 a_11691_44458# a_15493_43396# 1.33e-19
C4314 a_n913_45002# a_2813_43396# 5.93e-20
C4315 a_n356_44636# a_175_44278# 6.51e-20
C4316 a_14537_43396# a_n97_42460# 1.86e-20
C4317 a_18184_42460# a_15493_43940# 0.022388f
C4318 a_n357_42282# a_2987_42968# 4.17e-19
C4319 a_2711_45572# a_17595_43084# 2.52e-20
C4320 a_12549_44172# RST_Z 9.94e-19
C4321 a_11453_44696# a_16237_45028# 0.008411f
C4322 a_9290_44172# a_2711_45572# 0.030631f
C4323 a_8199_44636# a_6511_45714# 1.7e-19
C4324 a_5937_45572# a_6472_45840# 0.001997f
C4325 a_4646_46812# a_7229_43940# 0.104864f
C4326 a_n971_45724# a_8375_44464# 0.007671f
C4327 a_n237_47217# a_6109_44484# 4.56e-21
C4328 a_4419_46090# a_4808_45572# 0.004093f
C4329 a_3483_46348# a_5437_45600# 9.84e-20
C4330 a_n881_46662# a_16922_45042# 4.59e-20
C4331 a_8145_46902# a_413_45260# 2.46e-21
C4332 a_5755_42852# VDD 0.179985f
C4333 a_n784_42308# a_1736_39043# 1.49e-20
C4334 a_n3674_38216# a_n3690_38528# 4.64e-19
C4335 a_n1630_35242# a_n2302_39072# 5.02e-20
C4336 a_5534_30871# C9_P_btm 7.29e-20
C4337 a_n4318_37592# a_n4334_38528# 7.61e-20
C4338 a_15890_42674# a_15720_42674# 2.6e-19
C4339 a_14113_42308# a_13921_42308# 2.46e-19
C4340 a_18114_32519# a_13467_32519# 0.055508f
C4341 a_13249_42308# a_14456_42282# 1.37e-19
C4342 a_5111_44636# a_5837_42852# 7.13e-19
C4343 a_1176_45822# VDD 0.781481f
C4344 a_11823_42460# a_15051_42282# 0.367924f
C4345 a_n356_44636# a_10341_43396# 1.27e-20
C4346 a_10193_42453# a_10149_42308# 0.002618f
C4347 a_22315_44484# a_20974_43370# 1.76e-21
C4348 a_3422_30871# a_17538_32519# 0.005569f
C4349 a_20193_45348# a_20749_43396# 0.003298f
C4350 a_21076_30879# VCM 0.097317f
C4351 a_2998_44172# a_3353_43940# 3.09e-19
C4352 a_n2661_42834# a_7112_43396# 3.36e-20
C4353 a_n2661_43922# a_7287_43370# 2.05e-21
C4354 a_n1151_42308# a_7499_43940# 4.39e-20
C4355 a_15682_46116# a_16019_45002# 5.53e-19
C4356 a_10809_44734# a_10775_45002# 0.022389f
C4357 a_2324_44458# a_1307_43914# 0.129761f
C4358 a_10193_42453# a_11652_45724# 0.197229f
C4359 a_2711_45572# a_11064_45572# 2.3e-19
C4360 a_18900_46660# a_11691_44458# 6.04e-20
C4361 a_10490_45724# a_11322_45546# 0.246478f
C4362 a_8746_45002# a_11525_45546# 3.44e-21
C4363 a_11415_45002# a_21005_45260# 0.01592f
C4364 a_12741_44636# a_18184_42460# 0.041879f
C4365 a_768_44030# a_5495_43940# 0.017815f
C4366 a_20202_43084# a_21101_45002# 4.9e-19
C4367 a_n1613_43370# a_n630_44306# 0.003389f
C4368 a_16327_47482# a_21115_43940# 2.26e-21
C4369 a_15227_44166# a_17767_44458# 0.023473f
C4370 a_3483_46348# a_7418_45067# 3.85e-19
C4371 a_n1925_42282# a_3537_45260# 0.055426f
C4372 a_526_44458# a_4574_45260# 6.77e-19
C4373 a_6511_45714# a_8192_45572# 1.94e-20
C4374 a_n1741_47186# a_171_46873# 3.56e-20
C4375 a_n971_45724# a_n1925_46634# 0.163523f
C4376 a_20990_47178# a_12465_44636# 3.04e-19
C4377 a_18597_46090# a_11453_44696# 0.022871f
C4378 a_n3565_38502# a_n4209_37414# 0.029366f
C4379 a_n4209_38502# a_n3565_37414# 0.030019f
C4380 a_1209_47178# a_n2661_46634# 0.001337f
C4381 a_13507_46334# a_4883_46098# 4.09671f
C4382 a_9863_47436# a_9804_47204# 0.109361f
C4383 a_n1435_47204# a_n881_46662# 0.068194f
C4384 a_4958_30871# C0_N_btm 9.29e-20
C4385 a_n815_47178# a_n743_46660# 0.001755f
C4386 a_5495_43940# a_5755_42852# 8.96e-22
C4387 a_n2661_42282# a_n1423_42826# 2.27e-20
C4388 a_9313_44734# a_18695_43230# 5.53e-19
C4389 a_n2810_45028# a_n3420_37984# 5.66e-21
C4390 a_11652_45724# VDD 0.155048f
C4391 a_4235_43370# a_2982_43646# 7.35e-20
C4392 a_n97_42460# a_6547_43396# 8.98e-20
C4393 a_14021_43940# a_17499_43370# 0.011011f
C4394 a_n2956_37592# a_n3690_38304# 1.91e-20
C4395 a_3422_30871# a_19339_43156# 1.85e-21
C4396 a_15682_43940# a_4361_42308# 1.15e-20
C4397 a_15493_43396# a_4190_30871# 6e-19
C4398 a_12549_44172# a_16243_43396# 0.001317f
C4399 a_13059_46348# a_15493_43940# 1.93e-19
C4400 a_n357_42282# a_6298_44484# 3.34e-19
C4401 a_2957_45546# a_n699_43396# 2.21e-19
C4402 a_19900_46494# a_11967_42832# 2.43e-21
C4403 a_8696_44636# a_15595_45028# 1.68e-20
C4404 a_13507_46334# a_5649_42852# 0.136078f
C4405 a_1823_45246# a_5244_44056# 5.63e-19
C4406 a_3090_45724# a_5829_43940# 0.003937f
C4407 a_2277_45546# a_n2661_44458# 1.47e-21
C4408 a_3357_43084# a_n1059_45260# 0.003773f
C4409 a_21188_45572# a_413_45260# 2.54e-21
C4410 a_n443_42852# a_n2129_44697# 8.3e-20
C4411 a_n2293_46634# a_9145_43396# 0.238561f
C4412 a_21496_47436# a_21363_46634# 4.81e-20
C4413 a_13507_46334# a_21188_46660# 0.03408f
C4414 a_20894_47436# a_20731_47026# 2.28e-19
C4415 C1_N_btm VREF_GND 0.673422f
C4416 C0_N_btm VCM 0.717064f
C4417 a_n1741_47186# a_10903_43370# 0.066687f
C4418 a_2063_45854# a_6165_46155# 8.02e-20
C4419 a_n237_47217# a_9569_46155# 6.37e-20
C4420 START SINGLE_ENDED 0.002177f
C4421 VDD DATA[0] 1.05526f
C4422 a_12465_44636# a_20273_46660# 3.92e-21
C4423 a_3877_44458# a_5732_46660# 0.040487f
C4424 a_4646_46812# a_5907_46634# 0.037052f
C4425 a_4651_46660# a_5167_46660# 0.102946f
C4426 a_n1925_46634# a_8023_46660# 2.21e-19
C4427 a_n443_46116# a_2698_46116# 0.012019f
C4428 a_n1151_42308# a_4704_46090# 0.001193f
C4429 a_4007_47204# a_3483_46348# 1.93e-19
C4430 a_3785_47178# a_4185_45028# 2.07e-20
C4431 a_n881_46662# a_13885_46660# 2.09e-19
C4432 C3_N_btm VIN_N 0.455045f
C4433 a_4883_46098# a_20623_46660# 3.47e-20
C4434 a_16327_47482# a_11415_45002# 0.94171f
C4435 a_11453_44696# a_19123_46287# 0.021733f
C4436 C2_N_btm VREF 0.987884f
C4437 a_n1435_47204# a_n2157_46122# 1.63e-20
C4438 a_6151_47436# a_1823_45246# 3.85e-20
C4439 a_13747_46662# a_15009_46634# 6.01e-21
C4440 a_5807_45002# a_14976_45028# 0.026261f
C4441 a_13661_43548# a_3090_45724# 0.177565f
C4442 a_n2661_46634# a_10768_47026# 0.002208f
C4443 a_2107_46812# a_6755_46942# 0.002513f
C4444 a_9145_43396# a_5342_30871# 0.002082f
C4445 a_14358_43442# a_13635_43156# 8.12e-19
C4446 a_14579_43548# a_13460_43230# 1.97e-19
C4447 a_9028_43914# a_8685_42308# 1.61e-21
C4448 a_3080_42308# a_4649_42852# 5.53e-20
C4449 a_3539_42460# a_4743_43172# 8.63e-20
C4450 a_20512_43084# a_21613_42308# 2.76e-20
C4451 a_4361_42308# a_22223_43396# 9.86e-19
C4452 a_21855_43396# a_5649_42852# 0.057783f
C4453 a_13467_32519# a_13887_32519# 0.058303f
C4454 a_10341_43396# a_12379_42858# 2.27e-19
C4455 a_13490_45067# VDD 6.34e-20
C4456 a_375_42282# a_n2129_44697# 1.85e-20
C4457 a_6171_45002# a_13076_44458# 2.44e-20
C4458 a_n443_42852# a_15493_43396# 0.025952f
C4459 a_18341_45572# a_17517_44484# 1.28e-20
C4460 a_3090_45724# a_10835_43094# 0.008534f
C4461 a_768_44030# a_n784_42308# 3.1e-20
C4462 a_8953_45546# a_9803_43646# 0.091141f
C4463 a_n467_45028# a_n23_44458# 0.038286f
C4464 a_n143_45144# a_n356_44636# 4.67e-19
C4465 a_8953_45002# a_9838_44484# 0.013986f
C4466 a_626_44172# a_n2661_44458# 0.031248f
C4467 a_526_44458# a_1568_43370# 0.220609f
C4468 a_21588_30879# a_14097_32519# 0.056136f
C4469 a_22612_30879# a_22400_42852# 2.55e-19
C4470 a_2107_46812# a_8049_45260# 0.029889f
C4471 a_n743_46660# a_9751_46155# 3.19e-19
C4472 a_6755_46942# a_14493_46090# 1.15e-20
C4473 a_4915_47217# a_13163_45724# 1.03e-19
C4474 a_n881_46662# a_380_45546# 0.001604f
C4475 a_n1613_43370# a_n1099_45572# 0.025553f
C4476 a_18285_46348# a_18280_46660# 0.089884f
C4477 a_20273_46660# a_20528_46660# 0.056391f
C4478 a_20623_46660# a_21188_46660# 7.99e-20
C4479 a_19321_45002# a_16375_45002# 8.59e-21
C4480 a_5807_45002# a_18051_46116# 0.006001f
C4481 a_13747_46662# a_19431_46494# 1.74e-19
C4482 a_8846_46660# a_5937_45572# 2.62e-19
C4483 a_8270_45546# a_9569_46155# 1.61e-19
C4484 a_15368_46634# a_3483_46348# 1.42e-21
C4485 a_13059_46348# a_12741_44636# 0.02008f
C4486 a_3090_45724# a_4185_45028# 0.770164f
C4487 a_9313_45822# a_9049_44484# 0.119007f
C4488 a_3080_42308# a_1736_39043# 1.41e-19
C4489 a_16759_43396# a_15803_42450# 8.82e-20
C4490 a_791_42968# a_961_42354# 0.003403f
C4491 a_1847_42826# a_1184_42692# 0.001067f
C4492 a_18599_43230# a_18695_43230# 0.013793f
C4493 a_7845_44172# VDD 0.11772f
C4494 a_4361_42308# a_5934_30871# 0.092304f
C4495 a_5649_42852# a_7227_42308# 1.31e-19
C4496 a_743_42282# a_8325_42308# 0.02734f
C4497 a_13678_32519# a_6123_31319# 0.00363f
C4498 a_10341_43396# a_18727_42674# 1.72e-20
C4499 a_10193_42453# a_16759_43396# 5.51e-19
C4500 a_3537_45260# a_3737_43940# 0.012872f
C4501 a_n23_44458# a_n2661_43922# 0.007348f
C4502 a_n356_44636# a_n2293_43922# 0.025509f
C4503 a_n863_45724# a_685_42968# 0.052365f
C4504 a_20447_31679# a_14401_32519# 0.054145f
C4505 a_18114_32519# a_22315_44484# 0.017551f
C4506 a_4915_47217# DATA[5] 0.121371f
C4507 a_2711_45572# a_13467_32519# 2.9e-19
C4508 a_526_44458# a_4743_43172# 0.00549f
C4509 a_19963_31679# a_17538_32519# 0.051095f
C4510 a_5815_47464# DATA[3] 0.00149f
C4511 a_9067_47204# VDD 0.47483f
C4512 a_8375_44464# a_9313_44734# 8.59e-20
C4513 a_11823_42460# a_13749_43396# 1.72e-20
C4514 a_13556_45296# a_15493_43940# 2.77e-19
C4515 a_14976_45028# a_15143_45578# 0.005582f
C4516 a_15368_46634# a_14495_45572# 3.5e-20
C4517 a_765_45546# a_6511_45714# 5.27e-21
C4518 a_11735_46660# a_11682_45822# 1.59e-20
C4519 a_n2956_39768# a_n2956_37592# 0.047483f
C4520 a_n1925_46634# a_n2293_45010# 3.1e-20
C4521 a_2324_44458# a_8034_45724# 1.84e-19
C4522 a_14493_46090# a_8049_45260# 0.001687f
C4523 a_n2293_46098# a_n1099_45572# 0.069723f
C4524 a_n1853_46287# a_n452_45724# 0.080546f
C4525 a_12891_46348# a_6171_45002# 0.040434f
C4526 a_376_46348# a_n2661_45546# 4.24e-21
C4527 a_19321_45002# a_413_45260# 2.02e-19
C4528 a_768_44030# a_5691_45260# 4.31e-21
C4529 a_12549_44172# a_3232_43370# 3.99e-21
C4530 a_6755_46942# a_15903_45785# 0.192397f
C4531 a_n2293_46634# a_n1059_45260# 0.051525f
C4532 a_n2104_46634# a_n2017_45002# 7.56e-20
C4533 a_n2438_43548# a_n2840_45002# 0.002993f
C4534 a_n743_46660# a_n2661_45010# 8.45e-21
C4535 a_n1641_46494# a_n2293_45546# 1.27e-19
C4536 a_n1423_46090# a_n1079_45724# 1.85e-19
C4537 a_10903_43370# a_10586_45546# 0.238199f
C4538 a_6761_42308# a_5934_30871# 1.73e-20
C4539 a_13467_32519# EN_VIN_BSTR_N 0.031982f
C4540 a_16759_43396# VDD 0.191873f
C4541 a_2903_42308# a_5742_30871# 2.87e-20
C4542 a_4190_30871# C9_P_btm 0.002182f
C4543 a_3232_43370# a_5111_42852# 1.6e-21
C4544 a_3537_45260# a_8387_43230# 3.75e-19
C4545 a_n357_42282# a_13575_42558# 3.32e-21
C4546 a_n913_45002# a_15279_43071# 2.22e-19
C4547 a_n2956_39304# a_n2216_39072# 8.63e-19
C4548 a_n2956_38680# a_n2860_39072# 8.73e-19
C4549 a_11827_44484# a_14205_43396# 5.23e-22
C4550 a_20679_44626# a_11341_43940# 4.56e-20
C4551 a_20766_44850# a_20935_43940# 0.003556f
C4552 a_19279_43940# a_20623_43914# 1.14e-19
C4553 a_20835_44721# a_21115_43940# 3.62e-19
C4554 a_13259_45724# a_18907_42674# 4.44e-20
C4555 a_n2661_42834# a_9801_43940# 4.77e-19
C4556 a_18579_44172# a_19862_44208# 0.091151f
C4557 a_4223_44672# a_6293_42852# 2.53e-19
C4558 a_453_43940# a_1241_44260# 5.21e-19
C4559 a_5111_44636# a_7871_42858# 2.52e-19
C4560 a_5663_43940# a_7542_44172# 7.37e-21
C4561 a_1414_42308# a_1525_44260# 2.45e-19
C4562 a_n356_44636# a_n97_42460# 1.46232f
C4563 a_9313_44734# a_19319_43548# 1.9e-20
C4564 a_n2017_45002# a_15567_42826# 0.002448f
C4565 a_n1059_45260# a_5342_30871# 0.030512f
C4566 a_19900_46494# a_20273_45572# 9.45e-19
C4567 a_20708_46348# a_20107_45572# 0.007797f
C4568 a_5068_46348# a_413_45260# 2.65e-21
C4569 a_15015_46420# a_2437_43646# 1.91e-20
C4570 a_8953_45546# a_n913_45002# 0.052161f
C4571 a_3218_45724# a_3260_45572# 0.010055f
C4572 a_10586_45546# a_12016_45572# 6.73e-20
C4573 a_11415_45002# a_14537_43396# 0.04406f
C4574 a_12741_44636# a_13556_45296# 0.046411f
C4575 a_1823_45246# a_5111_44636# 0.002758f
C4576 a_584_46384# a_n2661_42282# 3.54e-21
C4577 a_3090_45724# a_18587_45118# 0.039584f
C4578 a_13925_46122# a_3357_43084# 1.09e-20
C4579 a_3147_46376# a_3065_45002# 2.49e-20
C4580 a_3699_46348# a_2382_45260# 2.18e-21
C4581 a_768_44030# a_13940_44484# 0.003215f
C4582 a_8049_45260# a_15903_45785# 0.003516f
C4583 a_13661_43548# a_14815_43914# 0.060575f
C4584 a_5257_43370# a_5343_44458# 0.063407f
C4585 a_n4315_30879# a_n2302_37984# 6.48e-20
C4586 a_1067_42314# VDD 0.128996f
C4587 a_n1741_47186# a_4883_46098# 0.031761f
C4588 a_n1630_35242# RST_Z 0.001585f
C4589 a_6123_31319# EN_VIN_BSTR_P 0.052187f
C4590 a_n4209_39304# a_n4209_38502# 0.042459f
C4591 a_1606_42308# C6_N_btm 2.33e-19
C4592 a_5934_30871# a_n1532_35090# 1.62e-19
C4593 a_n4064_40160# a_n2946_37984# 2.04e-20
C4594 a_7174_31319# VDAC_Pi 2.22e-19
C4595 a_n3565_39304# a_n2216_39072# 0.003034f
C4596 a_6151_47436# a_11031_47542# 0.03901f
C4597 a_6851_47204# a_6575_47204# 0.027563f
C4598 a_4915_47217# a_13381_47204# 0.045103f
C4599 a_7227_47204# a_7903_47542# 0.002513f
C4600 a_n443_46116# a_n1435_47204# 8.31e-19
C4601 a_22315_44484# a_13887_32519# 2.2e-22
C4602 a_9313_44734# a_16795_42852# 0.008194f
C4603 a_18184_42460# a_22765_42852# 0.012194f
C4604 a_9672_43914# a_9145_43396# 1.12e-19
C4605 a_n913_45002# a_13258_32519# 0.025596f
C4606 a_19963_31679# a_22465_38105# 3.53e-19
C4607 a_n2472_45546# VDD 0.290266f
C4608 a_20512_43084# a_4361_42308# 0.02826f
C4609 a_n2293_43922# a_12379_42858# 0.030458f
C4610 a_12429_44172# a_8685_43396# 2.43e-20
C4611 a_n2293_42834# a_2903_42308# 1.2e-20
C4612 a_n443_42852# a_45_45144# 2.99e-19
C4613 a_n452_45724# a_n2661_43370# 2.54e-20
C4614 a_8568_45546# a_8953_45002# 0.001119f
C4615 a_7499_43078# a_8191_45002# 0.002543f
C4616 a_11415_45002# a_20835_44721# 0.002797f
C4617 a_18479_45785# a_18596_45572# 0.183223f
C4618 a_18175_45572# a_18799_45938# 9.73e-19
C4619 a_18341_45572# a_19256_45572# 0.116691f
C4620 a_4099_45572# a_1423_45028# 2.06e-20
C4621 a_n2442_46660# a_n4318_39304# 0.023691f
C4622 a_8049_45260# a_n2661_44458# 5.47e-19
C4623 a_768_44030# a_3080_42308# 1.6e-19
C4624 a_n1613_43370# a_n1243_43396# 2.95e-19
C4625 a_10227_46804# a_14579_43548# 0.118896f
C4626 w_11334_34010# a_17364_32525# 0.016546f
C4627 a_12741_44636# a_20362_44736# 0.00339f
C4628 a_11322_45546# a_6171_45002# 0.069025f
C4629 a_11525_45546# a_3232_43370# 7.67e-19
C4630 a_526_44458# a_5883_43914# 0.0033f
C4631 w_1575_34946# a_5342_30871# 0.002142f
C4632 a_n2661_46634# a_288_46660# 0.002871f
C4633 a_1209_47178# a_765_45546# 0.003605f
C4634 a_n1613_43370# a_3878_46660# 0.002879f
C4635 a_n923_35174# a_n83_35174# 0.480251f
C4636 a_11453_44696# a_6755_46942# 0.026496f
C4637 VDAC_N C7_N_btm 30.844f
C4638 a_11599_46634# a_15009_46634# 6.85e-19
C4639 a_14955_47212# a_3090_45724# 0.009113f
C4640 a_n2438_43548# a_n133_46660# 0.848709f
C4641 a_n743_46660# a_171_46873# 0.075858f
C4642 a_768_44030# a_4646_46812# 0.047094f
C4643 a_n1925_46634# a_601_46902# 0.004874f
C4644 a_n1021_46688# a_33_46660# 1.18e-19
C4645 a_10227_46804# a_11186_47026# 0.018916f
C4646 a_3726_37500# VDD 0.341303f
C4647 a_13717_47436# a_16292_46812# 1.08e-20
C4648 a_12861_44030# a_15559_46634# 0.066578f
C4649 a_4905_42826# a_5111_42852# 0.105155f
C4650 a_n97_42460# a_12379_42858# 5.61e-19
C4651 a_11967_42832# a_12563_42308# 1.15e-20
C4652 a_7276_45260# VDD 0.093163f
C4653 a_2896_43646# a_1847_42826# 9.63e-20
C4654 a_9313_44734# a_21335_42336# 0.002222f
C4655 a_10341_43396# a_17486_43762# 1.07e-19
C4656 a_9145_43396# a_743_42282# 1.59e-19
C4657 a_16137_43396# a_16759_43396# 2.32e-19
C4658 a_16547_43609# a_16409_43396# 0.206231f
C4659 a_16243_43396# a_16977_43638# 0.053479f
C4660 a_4646_46812# a_5755_42852# 5.33e-19
C4661 a_15227_44166# a_18525_43370# 2.71e-21
C4662 a_3090_45724# a_15037_43396# 1.16e-20
C4663 a_n1613_43370# a_9306_43218# 0.001965f
C4664 a_8953_45002# a_n2661_43370# 0.034058f
C4665 a_10544_45572# a_9313_44734# 5.83e-20
C4666 a_16147_45260# a_14539_43914# 4.45e-20
C4667 a_n443_46116# a_1606_42308# 3.46e-19
C4668 a_4791_45118# a_1755_42282# 0.002644f
C4669 a_16327_47482# a_20256_42852# 8.08e-21
C4670 a_19963_31679# a_19721_31679# 9.01086f
C4671 a_n913_45002# a_20193_45348# 0.224918f
C4672 a_6171_45002# a_15060_45348# 2.19e-19
C4673 a_n357_42282# a_2479_44172# 0.008172f
C4674 a_10193_42453# a_17517_44484# 4.26e-19
C4675 a_1823_45246# a_4235_43370# 0.029154f
C4676 a_11823_42460# a_12553_44484# 1.28e-19
C4677 a_2107_46812# a_8953_45546# 0.007676f
C4678 a_13607_46688# a_13059_46348# 9.43e-19
C4679 a_2905_45572# a_3316_45546# 0.004332f
C4680 a_327_47204# a_n443_42852# 3.15e-21
C4681 a_n443_46116# a_380_45546# 0.073277f
C4682 a_11453_44696# a_8049_45260# 0.032046f
C4683 a_16327_47482# a_13259_45724# 0.584328f
C4684 a_19321_45002# a_18985_46122# 0.019556f
C4685 a_19594_46812# a_18819_46122# 1.63e-19
C4686 a_n743_46660# a_10903_43370# 0.080542f
C4687 a_13747_46662# a_19335_46494# 0.005102f
C4688 a_16697_47582# a_6945_45028# 1.16e-19
C4689 a_5807_45002# a_19900_46494# 0.00115f
C4690 a_n2109_47186# a_2711_45572# 0.032969f
C4691 a_n237_47217# a_1990_45899# 8.97e-19
C4692 a_3067_47026# a_3147_46376# 2.75e-19
C4693 a_3524_46660# a_3699_46348# 4.06e-19
C4694 a_n881_46662# a_526_44458# 0.060324f
C4695 a_10227_46804# a_12839_46116# 8.43e-21
C4696 a_4883_46098# a_10586_45546# 0.006953f
C4697 a_n1613_43370# a_n1925_42282# 1.08e-19
C4698 a_15559_46634# a_14180_46812# 0.001017f
C4699 a_n97_42460# a_18727_42674# 3.76e-20
C4700 a_17517_44484# VDD 2.99662f
C4701 a_4190_30871# a_18707_42852# 0.006254f
C4702 a_18083_42858# a_17333_42852# 0.284837f
C4703 a_17701_42308# a_18249_42858# 2.98e-20
C4704 a_2982_43646# a_15051_42282# 6.3e-19
C4705 SMPL_ON_P EN_VIN_BSTR_P 1.58e-19
C4706 a_n443_42852# a_10695_43548# 0.042055f
C4707 a_n2442_46660# a_n4334_40480# 3.24e-19
C4708 a_21363_45546# a_15493_43940# 1.34e-22
C4709 a_742_44458# a_n356_44636# 0.207503f
C4710 a_526_44458# a_133_43172# 3.34e-20
C4711 a_12607_44458# a_13076_44458# 0.200168f
C4712 a_n2017_45002# a_10405_44172# 1.01e-20
C4713 a_413_45260# a_2537_44260# 1.26e-19
C4714 a_3232_43370# a_7542_44172# 1.17e-20
C4715 a_n2661_44458# a_5289_44734# 5.74e-19
C4716 a_n2293_46098# a_n1925_42282# 0.020467f
C4717 a_6151_47436# a_6709_45028# 6.61e-22
C4718 a_n971_45724# a_2232_45348# 2.25e-19
C4719 a_8016_46348# a_2324_44458# 0.048711f
C4720 a_15811_47375# a_413_45260# 2.19e-19
C4721 a_11189_46129# a_10903_43370# 0.151119f
C4722 a_9290_44172# a_12005_46116# 1.48e-19
C4723 a_16388_46812# a_18243_46436# 0.004535f
C4724 a_12549_44172# a_18341_45572# 2.55e-20
C4725 a_n881_46662# a_17668_45572# 0.005485f
C4726 a_19987_42826# a_20107_42308# 0.001063f
C4727 a_20922_43172# a_13258_32519# 7.84e-20
C4728 a_n473_42460# a_1184_42692# 1.41e-19
C4729 a_n784_42308# a_1067_42314# 0.064066f
C4730 a_n327_42558# a_n1630_35242# 0.053474f
C4731 a_n3674_37592# a_564_42282# 1.04e-19
C4732 a_11554_42852# a_5742_30871# 3.85e-19
C4733 a_4223_44672# a_7499_43940# 0.030206f
C4734 a_n2661_42834# a_6101_44260# 2.26e-19
C4735 a_6171_45002# a_16409_43396# 6.7e-20
C4736 a_19479_31679# a_17364_32525# 0.05375f
C4737 a_5167_46660# VDD 0.203378f
C4738 a_n2293_42834# a_6293_42852# 0.008221f
C4739 a_9313_44734# a_10949_43914# 3.03e-20
C4740 a_3422_30871# a_22591_44484# 8.92e-19
C4741 a_n1059_45260# a_743_42282# 0.198704f
C4742 a_7499_43078# a_7309_42852# 0.011818f
C4743 a_n2810_45572# a_n3674_37592# 0.025877f
C4744 a_15004_44636# a_14021_43940# 7.55e-21
C4745 a_14797_45144# a_14955_43396# 4.74e-21
C4746 a_22315_44484# a_22485_44484# 0.109468f
C4747 a_12891_46348# a_12607_44458# 0.067773f
C4748 a_5807_45002# a_5343_44458# 4.88e-20
C4749 a_10809_44734# a_13163_45724# 4.78e-21
C4750 a_8062_46155# a_2711_45572# 1.41e-19
C4751 a_768_44030# a_10057_43914# 0.041949f
C4752 a_n2840_45546# a_n2810_45572# 0.162234f
C4753 a_11415_45002# a_20731_45938# 0.001207f
C4754 a_7577_46660# a_n2293_42834# 1.2e-20
C4755 a_10903_43370# a_11136_45572# 0.002788f
C4756 a_n2442_46660# a_n2661_44458# 2.17e-20
C4757 a_14976_45028# a_13017_45260# 2.91e-20
C4758 a_13059_46348# a_413_45260# 1.63e-20
C4759 a_2324_44458# a_11682_45822# 1.62e-20
C4760 COMP_P VDAC_N 0.003716f
C4761 a_n1741_47186# a_n1605_47204# 0.011722f
C4762 a_n2109_47186# a_n452_47436# 0.039314f
C4763 a_n2497_47436# a_n746_45260# 0.046973f
C4764 a_n1920_47178# a_n815_47178# 6.26e-20
C4765 a_14097_32519# a_22469_39537# 1.25e-20
C4766 a_5932_42308# VDAC_Pi 2.52e-19
C4767 a_4149_42891# VDD 0.001563f
C4768 a_22223_46124# EN_OFFSET_CAL 0.011048f
C4769 a_518_46482# VDD 3.14e-19
C4770 a_18326_43940# a_18533_44260# 6.08e-19
C4771 a_3905_42865# a_2982_43646# 0.006358f
C4772 a_6945_45028# CLK 0.027466f
C4773 a_20679_44626# a_10341_43396# 1.82e-20
C4774 a_n2956_38216# a_n4064_37440# 0.001421f
C4775 a_3600_43914# a_3540_43646# 1.75e-19
C4776 a_2998_44172# a_3626_43646# 1.65e-19
C4777 a_3537_45260# a_1606_42308# 3.89e-20
C4778 a_n1059_45260# a_5755_42308# 1.66e-19
C4779 a_n2017_45002# a_6171_42473# 0.003106f
C4780 a_n913_45002# a_5421_42558# 0.006411f
C4781 a_20193_45348# a_20922_43172# 7.72e-19
C4782 a_8701_44490# a_8387_43230# 1.48e-20
C4783 a_1414_42308# a_1512_43396# 8.62e-19
C4784 a_n2661_42282# a_n1177_43370# 1.78e-22
C4785 a_4185_45028# a_4743_44484# 0.007252f
C4786 a_3483_46348# a_5518_44484# 0.081879f
C4787 a_10907_45822# a_8696_44636# 0.001403f
C4788 a_n2661_45546# a_3232_43370# 0.038743f
C4789 a_4646_46812# a_7845_44172# 0.002985f
C4790 a_6472_45840# a_2437_43646# 3.74e-21
C4791 a_13259_45724# a_14537_43396# 0.083218f
C4792 a_15682_46116# a_11827_44484# 6.61e-22
C4793 a_n755_45592# a_2382_45260# 5.27e-19
C4794 a_1848_45724# a_1667_45002# 1.61e-19
C4795 a_3218_45724# a_413_45260# 0.016434f
C4796 a_4419_46090# a_n699_43396# 1.59e-20
C4797 a_8953_45546# a_n2661_44458# 0.019448f
C4798 a_13904_45546# a_14127_45572# 0.011458f
C4799 a_n443_42852# a_n745_45366# 4.76e-19
C4800 a_3090_45724# a_11967_42832# 0.12811f
C4801 a_19553_46090# a_19778_44110# 4.76e-20
C4802 a_2107_46812# a_9028_43914# 0.110155f
C4803 a_768_44030# a_14021_43940# 1.82e-19
C4804 a_12549_44172# a_14485_44260# 2.93e-20
C4805 a_14275_46494# a_11691_44458# 1.05e-20
C4806 a_n2312_40392# a_n2661_46634# 1.45e-20
C4807 a_n2312_39304# a_n2956_39768# 5.91067f
C4808 a_n4209_38216# C5_P_btm 1.11e-20
C4809 a_n3565_38216# C7_P_btm 1.43e-20
C4810 a_7754_38470# CAL_N 3.08e-19
C4811 a_8530_39574# a_11206_38545# 0.046219f
C4812 a_6151_47436# a_5732_46660# 0.002133f
C4813 a_n881_46662# a_13759_47204# 2.74e-19
C4814 a_1239_39043# VDD 0.507578f
C4815 a_n971_45724# a_6999_46987# 0.005614f
C4816 a_n1151_42308# a_7715_46873# 0.09029f
C4817 a_n237_47217# a_6969_46634# 1.13e-19
C4818 a_2063_45854# a_8492_46660# 0.005635f
C4819 a_4883_46098# a_n743_46660# 5.6639f
C4820 a_19256_45572# VDD 0.27151f
C4821 a_21381_43940# a_4361_42308# 0.195418f
C4822 a_14401_32519# a_13467_32519# 0.050489f
C4823 a_n2293_43922# a_3823_42558# 4.58e-20
C4824 a_n356_44636# a_10533_42308# 1.57e-19
C4825 a_14539_43914# a_15051_42282# 1.16e-20
C4826 a_11341_43940# a_10341_42308# 3.2e-20
C4827 a_5891_43370# a_5934_30871# 0.027588f
C4828 a_5244_44056# a_5193_42852# 3.06e-21
C4829 a_19963_31679# a_18194_35068# 1.2e-19
C4830 a_19479_31679# a_21589_35634# 7.02e-21
C4831 a_3232_43370# a_5205_44484# 0.217288f
C4832 a_768_44030# a_2075_43172# 0.00187f
C4833 a_n2956_38680# a_n3674_39768# 0.023133f
C4834 a_15765_45572# a_11691_44458# 3.92e-20
C4835 a_11525_45546# a_8975_43940# 1.35e-20
C4836 a_2711_45572# a_8375_44464# 1.54e-21
C4837 a_526_44458# a_2889_44172# 2.55e-20
C4838 a_6171_45002# a_6431_45366# 0.017465f
C4839 a_n1059_45260# a_626_44172# 2.24e-19
C4840 a_10903_43370# a_11750_44172# 0.135933f
C4841 a_3483_46348# a_9895_44260# 1.07e-19
C4842 a_n1613_43370# a_8387_43230# 0.163582f
C4843 a_11599_46634# a_19335_46494# 0.030852f
C4844 a_n237_47217# a_9241_46436# 2.14e-19
C4845 a_2063_45854# a_5210_46155# 1.39e-19
C4846 a_10428_46928# a_11735_46660# 0.001328f
C4847 a_10467_46802# a_11186_47026# 0.082642f
C4848 a_10623_46897# a_10768_47026# 0.057222f
C4849 a_n881_46662# a_2521_46116# 0.050613f
C4850 a_n1613_43370# a_2698_46116# 2.5e-20
C4851 a_16327_47482# a_18189_46348# 0.029513f
C4852 a_n1151_42308# a_5210_46482# 7.81e-19
C4853 a_288_46660# a_765_45546# 1.47e-21
C4854 a_5257_43370# a_3090_45724# 0.020885f
C4855 a_13381_47204# a_10809_44734# 1.08e-19
C4856 a_13717_47436# a_6945_45028# 0.038878f
C4857 a_4791_45118# a_n1925_42282# 1.87e-19
C4858 a_n443_46116# a_526_44458# 0.366438f
C4859 a_16588_47582# a_15682_46116# 0.00115f
C4860 a_10227_46804# a_14840_46494# 0.275527f
C4861 a_4883_46098# a_11189_46129# 0.008441f
C4862 a_n3674_39768# a_n3690_39392# 3.4e-19
C4863 a_n4318_39768# a_n3420_39072# 2.16e-21
C4864 a_15493_43396# a_19511_42282# 1.63e-19
C4865 a_5649_42852# a_17701_42308# 4.59e-20
C4866 a_21259_43561# a_21195_42852# 7.25e-20
C4867 a_4190_30871# a_21356_42826# 0.011885f
C4868 a_15493_43940# a_17303_42282# 7.91e-22
C4869 a_n1557_42282# a_n3674_37592# 0.022251f
C4870 a_13720_44458# VDD 0.202097f
C4871 a_4361_42308# a_18249_42858# 1.62e-19
C4872 a_19095_43396# a_18599_43230# 3.23e-19
C4873 a_n97_42460# a_3823_42558# 4.7e-21
C4874 a_743_42282# a_19987_42826# 0.009731f
C4875 a_19479_31679# a_19237_31679# 9.049419f
C4876 a_10903_43370# a_4361_42308# 0.00974f
C4877 a_22591_45572# a_17730_32519# 7.45e-20
C4878 a_12549_44172# a_15803_42450# 1.19e-21
C4879 a_2711_45572# a_19319_43548# 0.225335f
C4880 a_n863_45724# a_1756_43548# 9.82e-20
C4881 a_9482_43914# a_13857_44734# 0.011887f
C4882 a_19963_31679# a_22591_44484# 8.88e-20
C4883 a_n357_42282# a_n229_43646# 0.00541f
C4884 a_n2661_45546# a_4905_42826# 9.27e-20
C4885 a_13507_46334# a_18997_42308# 6.67e-19
C4886 a_3524_46660# a_n755_45592# 5.56e-20
C4887 a_4651_46660# a_n2661_45546# 2.36e-20
C4888 a_12549_44172# a_10193_42453# 0.116594f
C4889 a_768_44030# a_10180_45724# 7.51e-20
C4890 a_765_45546# a_15015_46420# 4.38e-20
C4891 a_11309_47204# a_10490_45724# 2.94e-20
C4892 a_n2497_47436# a_n2109_45247# 0.001006f
C4893 a_16327_47482# a_17478_45572# 0.012405f
C4894 a_n1925_46634# a_2711_45572# 0.030736f
C4895 a_n2661_46634# a_6472_45840# 1.74e-20
C4896 a_n2293_46098# a_2698_46116# 6.74e-20
C4897 a_n901_46420# a_1176_45822# 1.16e-19
C4898 a_n237_47217# a_3357_43084# 0.022871f
C4899 a_21076_30879# a_4185_45028# 2.52e-19
C4900 a_n881_46662# a_13163_45724# 2.21e-20
C4901 a_327_47204# a_2437_43646# 2.63e-19
C4902 a_14035_46660# a_6945_45028# 4.05e-19
C4903 a_16388_46812# a_18819_46122# 1.15e-19
C4904 a_10227_46804# a_16115_45572# 7.83e-19
C4905 a_13678_32519# a_22775_42308# 0.024479f
C4906 a_5649_42852# a_21613_42308# 0.02466f
C4907 a_10835_43094# a_11633_42558# 3.72e-19
C4908 a_726_44056# VDD 0.001151f
C4909 a_13467_32519# a_21421_42336# 6.18e-19
C4910 a_4361_42308# a_21125_42558# 2.86e-19
C4911 a_10991_42826# a_5742_30871# 0.002659f
C4912 a_10796_42968# a_11551_42558# 8.41e-19
C4913 a_10341_42308# a_10723_42308# 0.024028f
C4914 a_3080_42308# a_3726_37500# 0.004001f
C4915 a_17364_32525# a_13258_32519# 0.053358f
C4916 a_n2661_44458# a_9028_43914# 4.82e-21
C4917 a_7499_43078# a_7765_42852# 0.008252f
C4918 a_14815_43914# a_11967_42832# 5.37e-21
C4919 a_14673_44172# a_16241_44734# 0.002281f
C4920 a_9313_44734# a_3422_30871# 0.043499f
C4921 a_n881_46662# DATA[5] 0.082222f
C4922 a_9290_44172# a_5934_30871# 4.13e-20
C4923 a_8953_45546# a_8325_42308# 0.002755f
C4924 a_8199_44636# a_8791_42308# 6.71e-19
C4925 a_8016_46348# a_9803_42558# 1.11e-20
C4926 a_7989_47542# DATA[4] 1.37e-19
C4927 a_21005_45260# a_20935_43940# 4.06e-20
C4928 a_11827_44484# a_20269_44172# 0.002504f
C4929 a_12549_44172# VDD 3.08339f
C4930 a_3537_45260# a_3539_42460# 0.264936f
C4931 a_18494_42460# a_11341_43940# 0.025825f
C4932 a_19778_44110# a_15493_43940# 0.033844f
C4933 a_n1925_42282# a_n1736_42282# 0.029727f
C4934 a_n357_42282# a_1793_42852# 5.15e-19
C4935 a_12891_46348# RST_Z 9.63e-21
C4936 a_10355_46116# a_2711_45572# 3.59e-20
C4937 a_5937_45572# a_6194_45824# 0.002515f
C4938 a_8199_44636# a_6472_45840# 0.001875f
C4939 a_4646_46812# a_7276_45260# 0.016809f
C4940 a_5167_46660# a_5691_45260# 7.13e-20
C4941 a_8049_45260# a_14180_46482# 9.26e-19
C4942 a_n971_45724# a_7640_43914# 5.53e-20
C4943 a_4419_46090# a_5024_45822# 8.88e-19
C4944 a_19466_46812# a_18799_45938# 2.72e-19
C4945 a_6755_46942# a_n1059_45260# 1.35e-20
C4946 a_17609_46634# a_17668_45572# 1.45e-20
C4947 a_7577_46660# a_413_45260# 3.89e-21
C4948 a_5111_42852# VDD 0.178652f
C4949 a_5534_30871# C10_P_btm 1.08e-19
C4950 a_n1630_35242# a_n4064_39072# 1.85e-20
C4951 a_n4318_38216# a_n3420_38528# 0.31769f
C4952 a_n3674_38680# a_n4064_38528# 0.557806f
C4953 COMP_P a_2112_39137# 1.26e-21
C4954 a_14113_42308# a_13657_42308# 6.05e-20
C4955 a_n4318_37592# a_n4209_38502# 1.31e-19
C4956 a_1606_42308# a_1343_38525# 1.72e-20
C4957 a_n2661_43922# a_6547_43396# 6.85e-21
C4958 a_n2661_42834# a_7287_43370# 1.79e-19
C4959 a_5111_44636# a_5193_42852# 0.018763f
C4960 a_13249_42308# a_13575_42558# 0.088907f
C4961 a_1208_46090# VDD 0.178097f
C4962 a_20193_45348# a_17364_32525# 1.2e-19
C4963 a_11823_42460# a_14113_42308# 0.103699f
C4964 a_n2810_45572# a_n2302_39072# 2.61e-19
C4965 a_10193_42453# a_9885_42308# 2.33e-20
C4966 a_n1059_45260# a_16328_43172# 0.009298f
C4967 a_n901_46420# DATA[0] 2.21e-19
C4968 a_3422_30871# a_20974_43370# 0.020902f
C4969 a_22315_44484# a_14401_32519# 0.002016f
C4970 a_21076_30879# VREF_GND 0.041931f
C4971 a_2889_44172# a_3353_43940# 6.46e-21
C4972 a_2998_44172# a_3052_44056# 3.81e-19
C4973 a_15682_46116# a_15595_45028# 1.03e-20
C4974 a_10809_44734# a_8953_45002# 0.001885f
C4975 a_2711_45572# a_10544_45572# 2.65e-19
C4976 a_15227_44166# a_16979_44734# 0.181002f
C4977 a_3090_45724# a_18989_43940# 0.095784f
C4978 a_12465_44636# a_10949_43914# 3.08e-19
C4979 a_10193_42453# a_11525_45546# 0.0979f
C4980 a_7499_43078# a_11823_42460# 0.002874f
C4981 a_8746_45002# a_11322_45546# 3.97e-21
C4982 a_11415_45002# a_20567_45036# 0.011165f
C4983 a_12741_44636# a_19778_44110# 0.070586f
C4984 a_768_44030# a_5013_44260# 0.064017f
C4985 a_20202_43084# a_21005_45260# 1.88e-19
C4986 a_n1613_43370# a_n875_44318# 7.2e-19
C4987 a_16327_47482# a_20935_43940# 0.004638f
C4988 a_3483_46348# a_10903_45394# 0.002881f
C4989 a_167_45260# a_n2661_43370# 0.055202f
C4990 a_526_44458# a_3537_45260# 0.938783f
C4991 a_5937_45572# a_6517_45366# 2.26e-19
C4992 a_15720_42674# RST_Z 6.53e-21
C4993 a_n4209_38502# a_n4334_37440# 3.34e-19
C4994 a_2684_37794# a_3754_38802# 9.44e-20
C4995 a_4958_30871# C0_dummy_N_btm 1.65e-20
C4996 a_n2109_47186# a_33_46660# 6.32e-20
C4997 a_n815_47178# a_n1021_46688# 0.003455f
C4998 a_20894_47436# a_12465_44636# 2.12e-19
C4999 a_n237_47217# a_n2293_46634# 0.003267f
C5000 a_327_47204# a_n2661_46634# 0.004931f
C5001 a_n1151_42308# a_13747_46662# 0.050569f
C5002 a_6151_47436# a_15928_47570# 2.62e-20
C5003 a_21177_47436# a_4883_46098# 5.42e-19
C5004 a_18780_47178# a_11453_44696# 2.2e-19
C5005 a_9067_47204# a_9804_47204# 0.001602f
C5006 a_13381_47204# a_n881_46662# 0.025748f
C5007 a_n1435_47204# a_n1613_43370# 2.68e-19
C5008 a_13507_46334# a_21496_47436# 0.167302f
C5009 a_n1741_47186# a_n133_46660# 4.48e-20
C5010 SMPL_ON_P a_n2438_43548# 0.003035f
C5011 a_n2661_42282# a_n1991_42858# 7.14e-21
C5012 a_5495_43940# a_5111_42852# 5.29e-20
C5013 a_9313_44734# a_18504_43218# 0.002026f
C5014 a_15037_43940# a_9145_43396# 3.15e-19
C5015 a_4093_43548# a_2982_43646# 1.2e-20
C5016 a_n229_43646# a_n144_43396# 1.48e-19
C5017 a_n97_42460# a_6765_43638# 2.79e-19
C5018 a_14021_43940# a_16759_43396# 0.007414f
C5019 a_n2956_37592# a_n3565_38216# 0.074137f
C5020 a_11525_45546# VDD 0.133093f
C5021 a_n2293_43922# a_12800_43218# 0.011493f
C5022 a_3422_30871# a_18599_43230# 6.68e-21
C5023 a_19328_44172# a_4190_30871# 4.64e-22
C5024 a_12549_44172# a_16137_43396# 0.003438f
C5025 a_18479_47436# a_20749_43396# 4.66e-19
C5026 a_13661_43548# a_12281_43396# 1.07e-19
C5027 a_17339_46660# a_19478_44306# 9.54e-21
C5028 a_20075_46420# a_11967_42832# 1.89e-21
C5029 a_19335_46494# a_19615_44636# 2.3e-20
C5030 a_16115_45572# a_1307_43914# 0.001401f
C5031 a_8696_44636# a_15415_45028# 4.71e-20
C5032 a_13259_45724# a_n356_44636# 0.026337f
C5033 a_13507_46334# a_13678_32519# 0.037522f
C5034 a_4883_46098# a_4361_42308# 9.17e-20
C5035 a_1823_45246# a_3905_42865# 0.218008f
C5036 a_3090_45724# a_5745_43940# 0.003797f
C5037 a_n755_45592# a_5343_44458# 0.349527f
C5038 a_1609_45822# a_n2661_44458# 2.15e-19
C5039 a_3357_43084# a_n2017_45002# 3.91e-19
C5040 a_3218_45724# a_2779_44458# 3.4e-20
C5041 a_11453_44696# a_18285_46348# 0.236771f
C5042 a_13507_46334# a_21363_46634# 0.029223f
C5043 a_21177_47436# a_21188_46660# 5.06e-21
C5044 C0_N_btm VREF_GND 0.350401f
C5045 C0_dummy_N_btm VCM 0.311452f
C5046 VDD CLK_DATA 0.422202f
C5047 a_n1741_47186# a_11387_46155# 4.53e-19
C5048 a_n237_47217# a_9625_46129# 2.69e-19
C5049 a_2063_45854# a_5497_46414# 1.5e-19
C5050 a_12465_44636# a_20411_46873# 2.37e-20
C5051 RST_Z SINGLE_ENDED 0.0318f
C5052 a_3877_44458# a_5907_46634# 0.073504f
C5053 a_4646_46812# a_5167_46660# 0.033486f
C5054 a_4651_46660# a_5385_46902# 0.053479f
C5055 a_n1151_42308# a_4419_46090# 2.82e-19
C5056 a_n443_46116# a_2521_46116# 0.00999f
C5057 a_3785_47178# a_3699_46348# 4.8e-20
C5058 a_3815_47204# a_3483_46348# 2.65e-20
C5059 a_11309_47204# a_12156_46660# 4.26e-19
C5060 C2_N_btm VIN_N 0.502408f
C5061 a_4883_46098# a_20841_46902# 7.76e-20
C5062 a_16327_47482# a_20202_43084# 0.475502f
C5063 C1_N_btm VREF 0.98698f
C5064 a_13747_46662# a_14084_46812# 0.038349f
C5065 a_5807_45002# a_3090_45724# 0.032418f
C5066 a_n2293_46634# a_8270_45546# 0.030248f
C5067 a_2107_46812# a_10249_46116# 4.12e-19
C5068 a_4955_46873# a_4817_46660# 0.318259f
C5069 a_18479_47436# a_18280_46660# 4.42e-20
C5070 a_13667_43396# a_13460_43230# 8.37e-20
C5071 a_14579_43548# a_13635_43156# 0.003436f
C5072 a_4699_43561# a_4649_42852# 1.98e-20
C5073 a_3080_42308# a_4149_42891# 0.001517f
C5074 a_3539_42460# a_4649_43172# 0.001762f
C5075 a_n97_42460# a_12800_43218# 4.03e-19
C5076 a_19237_31679# a_13258_32519# 0.055803f
C5077 a_20512_43084# a_21887_42336# 1.58e-19
C5078 a_21855_43396# a_13678_32519# 0.17881f
C5079 a_4361_42308# a_5649_42852# 0.064476f
C5080 a_4190_30871# a_20749_43396# 0.018962f
C5081 a_10341_43396# a_10341_42308# 9.26e-19
C5082 a_12281_43396# a_10835_43094# 3.18e-20
C5083 a_4185_45028# a_12281_43396# 1.62e-19
C5084 a_9482_43914# a_4223_44672# 3.83e-21
C5085 a_3232_43370# a_13076_44458# 4.99e-21
C5086 a_18479_45785# a_17517_44484# 0.023114f
C5087 a_3090_45724# a_10518_42984# 0.004978f
C5088 a_8953_45546# a_9145_43396# 0.019849f
C5089 a_n467_45028# a_n356_44636# 0.052527f
C5090 a_2324_44458# a_8791_43396# 3.85e-21
C5091 a_8953_45002# a_5883_43914# 0.008516f
C5092 a_526_44458# a_1049_43396# 0.121121f
C5093 a_21588_30879# a_22400_42852# 2.09e-19
C5094 w_1575_34946# a_n4064_37984# 3.17e-19
C5095 a_2107_46812# a_8781_46436# 2.53e-19
C5096 a_6755_46942# a_13925_46122# 4.42e-19
C5097 a_10428_46928# a_2324_44458# 7.92e-21
C5098 a_20107_46660# a_20731_47026# 9.73e-19
C5099 a_20411_46873# a_20528_46660# 0.170785f
C5100 a_20841_46902# a_21188_46660# 0.051162f
C5101 a_20273_46660# a_22000_46634# 2.02e-19
C5102 a_18285_46348# a_17639_46660# 0.003315f
C5103 a_13747_46662# a_19240_46482# 0.012097f
C5104 a_8270_45546# a_9625_46129# 0.001176f
C5105 a_8846_46660# a_8199_44636# 6.28e-20
C5106 a_9863_47436# a_10053_45546# 3.03e-20
C5107 a_n881_46662# a_n452_45724# 0.005284f
C5108 a_14976_45028# a_3483_46348# 3.99e-20
C5109 a_n237_47217# a_9159_45572# 3.1e-20
C5110 a_5649_42852# a_6761_42308# 9.04e-20
C5111 a_13467_32519# a_5934_30871# 0.003932f
C5112 a_743_42282# a_8337_42558# 4.14e-19
C5113 a_5111_42852# a_n784_42308# 3.45e-21
C5114 a_3080_42308# a_1239_39043# 1.03e-19
C5115 a_16977_43638# a_15803_42450# 9.29e-20
C5116 a_4361_42308# a_7963_42308# 0.007925f
C5117 a_791_42968# a_1184_42692# 8.46e-19
C5118 a_1847_42826# a_1576_42282# 2.07e-19
C5119 a_8292_43218# a_8483_43230# 4.61e-19
C5120 a_16795_42852# a_16877_42852# 0.171361f
C5121 a_18599_43230# a_18504_43218# 0.049827f
C5122 a_18817_42826# a_18695_43230# 3.16e-19
C5123 a_7542_44172# VDD 0.412456f
C5124 a_10341_43396# a_18057_42282# 5.97e-21
C5125 a_5815_47464# DATA[2] 9.97e-21
C5126 a_10193_42453# a_16977_43638# 7.87e-19
C5127 a_n356_44636# a_n2661_43922# 0.041936f
C5128 a_n23_44458# a_n2661_42834# 0.001339f
C5129 a_7640_43914# a_9313_44734# 0.001487f
C5130 a_n863_45724# a_421_43172# 0.00331f
C5131 a_13259_45724# a_12379_42858# 0.001312f
C5132 a_3065_45002# a_3992_43940# 0.002689f
C5133 a_13720_44458# a_13940_44484# 0.009965f
C5134 a_18114_32519# a_3422_30871# 0.001438f
C5135 a_5129_47502# DATA[3] 4.21e-20
C5136 a_6575_47204# VDD 1.32036f
C5137 a_9482_43914# a_15493_43940# 1.42e-19
C5138 a_13777_45326# a_11341_43940# 3.2e-21
C5139 a_4915_47217# DATA[4] 0.069022f
C5140 a_526_44458# a_4649_43172# 0.005678f
C5141 a_n1991_46122# a_n1079_45724# 0.001345f
C5142 a_765_45546# a_6472_45840# 1.39e-20
C5143 a_3090_45724# a_15143_45578# 0.016572f
C5144 a_8270_45546# a_9159_45572# 8.13e-20
C5145 a_15368_46634# a_13249_42308# 4.76e-21
C5146 a_768_44030# a_4927_45028# 4.62e-21
C5147 a_22612_30879# en_comp 5.56e-19
C5148 a_13925_46122# a_8049_45260# 0.009027f
C5149 a_n2293_46098# a_380_45546# 0.007518f
C5150 a_n1853_46287# a_n863_45724# 0.019522f
C5151 a_n1076_46494# a_n2661_45546# 1.51e-20
C5152 a_12891_46348# a_3232_43370# 8.12e-21
C5153 a_6755_46942# a_15599_45572# 0.024601f
C5154 a_15227_44166# a_11823_42460# 1.79e-19
C5155 a_11309_47204# a_6171_45002# 3.85e-20
C5156 a_n2293_46634# a_n2017_45002# 0.039556f
C5157 a_n2956_39768# a_n2810_45028# 0.04304f
C5158 a_1983_46706# a_2437_43646# 0.01301f
C5159 a_n1423_46090# a_n2293_45546# 0.001036f
C5160 a_11387_46155# a_10586_45546# 7.66e-19
C5161 a_13467_32519# a_11530_34132# 0.002259f
C5162 a_4190_30871# C10_P_btm 0.446355f
C5163 a_16977_43638# VDD 0.206333f
C5164 a_2713_42308# a_5742_30871# 1.69e-20
C5165 a_6761_42308# a_7963_42308# 9.72e-20
C5166 a_7227_42308# a_6123_31319# 0.189956f
C5167 a_3537_45260# a_8605_42826# 2.91e-20
C5168 a_15559_46634# CLK 2.96e-21
C5169 a_n357_42282# a_13070_42354# 1.72e-20
C5170 a_n913_45002# a_5534_30871# 0.274894f
C5171 a_n1059_45260# a_15279_43071# 0.021145f
C5172 a_n2956_39304# a_n2860_39072# 0.001353f
C5173 a_18494_42460# a_10341_43396# 0.030934f
C5174 a_20159_44458# a_15493_43940# 7.59e-20
C5175 a_20835_44721# a_20935_43940# 4.15e-19
C5176 a_20640_44752# a_11341_43940# 4.18e-22
C5177 a_20679_44626# a_21115_43940# 0.003825f
C5178 a_19279_43940# a_20365_43914# 0.003068f
C5179 a_20820_30879# a_22459_39145# 3.4e-20
C5180 a_13259_45724# a_18727_42674# 8.73e-20
C5181 a_17517_44484# a_14021_43940# 6.77e-21
C5182 a_4223_44672# a_6031_43396# 1.22e-19
C5183 a_21076_30879# a_22469_40625# 6.02e-20
C5184 a_5111_44636# a_7227_42852# 1.22e-20
C5185 a_1414_42308# a_1241_44260# 9.75e-20
C5186 a_18579_44172# a_19478_44306# 0.040429f
C5187 a_n2017_45002# a_5342_30871# 0.038471f
C5188 a_n443_42852# a_8685_42308# 6.23e-22
C5189 a_19900_46494# a_20107_45572# 1.7e-19
C5190 a_20075_46420# a_20273_45572# 1.19e-20
C5191 a_8953_45546# a_n1059_45260# 0.318691f
C5192 a_3503_45724# a_3733_45822# 0.004937f
C5193 a_2957_45546# a_3260_45572# 0.001377f
C5194 a_10586_45546# a_11778_45572# 0.006085f
C5195 a_12741_44636# a_9482_43914# 0.101234f
C5196 a_11415_45002# a_14180_45002# 0.025987f
C5197 a_1823_45246# a_5147_45002# 0.001658f
C5198 a_3090_45724# a_18315_45260# 0.061731f
C5199 a_13759_46122# a_3357_43084# 1.98e-20
C5200 a_3147_46376# a_2680_45002# 3.68e-20
C5201 a_3483_46348# a_2382_45260# 1.72e-21
C5202 a_768_44030# a_13296_44484# 0.001019f
C5203 a_8049_45260# a_15599_45572# 0.003996f
C5204 a_5257_43370# a_4743_44484# 7.16e-21
C5205 a_n4315_30879# a_n4064_37984# 0.034375f
C5206 a_n1630_35242# VDD 3.16282f
C5207 a_6123_31319# a_n923_35174# 0.008058f
C5208 a_n4209_39590# a_n4209_38216# 0.031951f
C5209 a_1606_42308# C5_N_btm 1.89e-19
C5210 a_n1151_42308# a_11599_46634# 0.116147f
C5211 a_n4064_40160# a_n3420_37984# 0.053114f
C5212 a_n3565_39304# a_n2860_39072# 0.001021f
C5213 a_n4064_39072# a_n3607_39392# 4.68e-19
C5214 a_6151_47436# a_9863_47436# 0.030884f
C5215 a_4915_47217# a_11459_47204# 0.03966f
C5216 a_6491_46660# a_6575_47204# 0.029984f
C5217 a_4791_45118# a_n1435_47204# 5.92e-19
C5218 a_3422_30871# a_13887_32519# 0.031713f
C5219 a_9313_44734# a_16414_43172# 0.007521f
C5220 a_18494_42460# a_20356_42852# 0.014237f
C5221 a_18184_42460# a_20753_42852# 0.029113f
C5222 a_n913_45002# a_19647_42308# 3.13e-19
C5223 a_n1059_45260# a_13258_32519# 4.14e-21
C5224 a_n2661_45546# VDD 0.733118f
C5225 a_20512_43084# a_13467_32519# 0.021245f
C5226 a_n2661_43922# a_12379_42858# 2.39e-19
C5227 a_n2293_43922# a_10341_42308# 1.51e-20
C5228 a_n2661_42834# a_12089_42308# 1.12e-20
C5229 a_1307_43914# a_9223_42460# 3.82e-21
C5230 a_6511_45714# a_1307_43914# 9.73e-22
C5231 a_n863_45724# a_n2661_43370# 0.076347f
C5232 a_10903_43370# a_5891_43370# 1.39e-19
C5233 a_8568_45546# a_8191_45002# 9.41e-20
C5234 a_7499_43078# a_7705_45326# 2.7e-19
C5235 a_11415_45002# a_20679_44626# 0.007381f
C5236 a_8270_45546# a_9672_43914# 0.003127f
C5237 a_18175_45572# a_18596_45572# 0.086708f
C5238 a_18341_45572# a_19431_45546# 0.041762f
C5239 a_18909_45814# a_18691_45572# 0.209641f
C5240 a_18479_45785# a_19256_45572# 0.044595f
C5241 a_768_44030# a_4699_43561# 4.91e-20
C5242 a_18051_46116# a_17719_45144# 1.04e-20
C5243 a_10490_45724# a_6171_45002# 3.24e-19
C5244 a_10227_46804# a_13667_43396# 0.007746f
C5245 a_6755_46942# a_18326_43940# 1.01e-19
C5246 a_12741_44636# a_20159_44458# 0.006194f
C5247 a_3483_46348# a_15433_44458# 4.08e-20
C5248 a_11322_45546# a_3232_43370# 4.14e-19
C5249 a_n1925_46634# a_33_46660# 0.0095f
C5250 a_n1021_46688# a_171_46873# 1.98e-19
C5251 a_327_47204# a_765_45546# 8.96e-19
C5252 a_n1613_43370# a_3633_46660# 6.03e-19
C5253 a_n1532_35090# a_n83_35174# 0.558402f
C5254 a_n923_35174# EN_VIN_BSTR_P 1.02927f
C5255 VDAC_N C6_N_btm 15.440799f
C5256 a_14955_47212# a_15009_46634# 0.001517f
C5257 a_n743_46660# a_n133_46660# 0.205551f
C5258 a_n2661_46634# a_1983_46706# 0.005467f
C5259 a_n2293_46634# a_1123_46634# 6.6e-21
C5260 a_768_44030# a_3877_44458# 0.012394f
C5261 a_10227_46804# a_10768_47026# 0.012196f
C5262 a_n3607_37440# VDD 2.79e-20
C5263 a_12861_44030# a_15368_46634# 0.066698f
C5264 a_13717_47436# a_15559_46634# 2.06e-21
C5265 a_n1151_42308# a_13693_46688# 2.97e-19
C5266 a_4905_42826# a_4520_42826# 0.147708f
C5267 a_n97_42460# a_10341_42308# 0.005646f
C5268 a_5205_44484# VDD 0.508148f
C5269 a_18533_43940# a_18249_42858# 1.68e-20
C5270 a_895_43940# a_1755_42282# 3.72e-21
C5271 a_9313_44734# a_7174_31319# 1.37e-19
C5272 a_10341_43396# a_15940_43402# 4.63e-19
C5273 a_8685_43396# a_4361_42308# 1.36e-19
C5274 a_16137_43396# a_16977_43638# 6.31e-20
C5275 a_16243_43396# a_16409_43396# 0.575934f
C5276 a_2711_45572# a_3422_30871# 1.83e-19
C5277 a_n1613_43370# a_9061_43230# 2.95e-19
C5278 a_8191_45002# a_n2661_43370# 0.013381f
C5279 a_n356_45724# a_n809_44244# 3.24e-21
C5280 a_16147_45260# a_16112_44458# 7.04e-19
C5281 a_n863_45724# a_2998_44172# 2.34e-19
C5282 a_22591_45572# a_19721_31679# 0.001292f
C5283 a_16327_47482# a_19326_42852# 2.94e-19
C5284 a_4791_45118# a_1606_42308# 3.68e-20
C5285 a_8270_45546# a_743_42282# 9.44e-21
C5286 a_19963_31679# a_18114_32519# 0.051445f
C5287 a_n913_45002# a_11691_44458# 2.08e-20
C5288 a_n2293_46098# a_3539_42460# 4.77e-19
C5289 a_n357_42282# a_2127_44172# 0.00145f
C5290 a_6171_45002# a_14976_45348# 1.2e-19
C5291 a_n755_45592# a_453_43940# 0.003942f
C5292 a_10193_42453# a_17061_44734# 0.012286f
C5293 a_1823_45246# a_4093_43548# 0.17443f
C5294 a_2107_46812# a_5937_45572# 0.027091f
C5295 a_3785_47178# a_n755_45592# 8.67e-21
C5296 a_12816_46660# a_13059_46348# 3.67e-19
C5297 a_2905_45572# a_3218_45724# 0.021505f
C5298 a_n237_47217# a_2277_45546# 0.104529f
C5299 a_n1151_42308# a_1848_45724# 7.61e-21
C5300 a_327_47204# a_509_45822# 1.76e-20
C5301 SMPL_ON_N a_8049_45260# 1.15e-19
C5302 a_19321_45002# a_18819_46122# 0.018323f
C5303 a_n743_46660# a_11387_46155# 0.007599f
C5304 a_13747_46662# a_19553_46090# 3.31e-20
C5305 a_16285_47570# a_6945_45028# 1.12e-19
C5306 a_5807_45002# a_20075_46420# 4.74e-19
C5307 a_3699_46634# a_3699_46348# 0.005275f
C5308 a_3524_46660# a_3483_46348# 6.03e-20
C5309 a_n443_46116# a_n452_45724# 0.188857f
C5310 a_11599_46634# a_19240_46482# 0.016662f
C5311 a_n1613_43370# a_526_44458# 0.826565f
C5312 a_15368_46634# a_14180_46812# 4.62e-20
C5313 a_n881_46662# a_2981_46116# 0.026038f
C5314 a_n97_42460# a_18057_42282# 2.69e-20
C5315 a_9396_43370# a_9223_42460# 4.27e-20
C5316 a_17061_44734# VDD 0.17647f
C5317 a_17701_42308# a_17333_42852# 0.061051f
C5318 a_17595_43084# a_18249_42858# 2.35e-19
C5319 a_3422_30871# EN_VIN_BSTR_N 0.182769f
C5320 a_5755_42852# a_6101_43172# 0.013377f
C5321 a_2982_43646# a_14113_42308# 2.12e-19
C5322 a_n2956_39768# a_n2302_40160# 3.63e-19
C5323 a_n1699_44726# a_n1243_44484# 4.2e-19
C5324 a_5205_44484# a_5495_43940# 4.22e-20
C5325 SMPL_ON_P a_n923_35174# 2.32e-19
C5326 a_n2442_46660# a_n4315_30879# 0.361271f
C5327 a_20623_45572# a_15493_43940# 1.03e-21
C5328 w_11334_34010# a_19864_35138# 0.005843f
C5329 a_n1352_44484# a_n23_44458# 2.56e-20
C5330 a_n452_44636# a_n356_44636# 0.318214f
C5331 a_11827_44484# a_10617_44484# 1.33e-19
C5332 a_n967_45348# a_n2661_42282# 2.72e-19
C5333 a_n443_42852# a_9803_43646# 0.102893f
C5334 a_n1059_45260# a_9028_43914# 0.002455f
C5335 a_n913_45002# a_8333_44056# 3.9e-21
C5336 a_413_45260# a_2253_44260# 1.2e-19
C5337 a_3232_43370# a_7281_43914# 0.001158f
C5338 a_6171_45002# a_6453_43914# 1.38e-19
C5339 a_n2661_44458# a_5205_44734# 2.45e-19
C5340 a_7499_43078# a_2982_43646# 6.36e-19
C5341 a_12607_44458# a_12883_44458# 0.11453f
C5342 a_n2293_46098# a_526_44458# 0.053029f
C5343 a_16388_46812# a_18147_46436# 0.004345f
C5344 a_22959_47212# a_2437_43646# 4.39e-19
C5345 a_n971_45724# a_1423_45028# 0.021147f
C5346 a_7920_46348# a_2324_44458# 6.6e-21
C5347 a_n1423_46090# a_n914_46116# 2.6e-19
C5348 a_n1151_42308# a_13348_45260# 3.18e-22
C5349 a_3090_45724# a_n755_45592# 0.051041f
C5350 a_4883_46098# a_20447_31679# 0.003751f
C5351 a_9290_44172# a_10903_43370# 0.340316f
C5352 a_11189_46129# a_11387_46155# 0.320331f
C5353 a_15507_47210# a_413_45260# 3.64e-19
C5354 a_18597_46090# a_n2017_45002# 2.49e-21
C5355 SMPL_ON_N a_19479_31679# 0.029207f
C5356 a_n881_46662# a_17568_45572# 0.001221f
C5357 a_12549_44172# a_18479_45785# 0.105486f
C5358 a_19987_42826# a_13258_32519# 2.93e-19
C5359 a_n4318_38680# a_n4064_38528# 0.047936f
C5360 a_18599_43230# a_7174_31319# 2.71e-21
C5361 a_n784_42308# a_n1630_35242# 0.063076f
C5362 a_11301_43218# a_5742_30871# 1.38e-19
C5363 a_1427_43646# VDD 0.19291f
C5364 a_14797_45144# a_15095_43370# 1.1e-20
C5365 a_14537_43396# a_14955_43396# 0.027267f
C5366 a_4223_44672# a_6671_43940# 0.03251f
C5367 a_n2293_43922# a_3499_42826# 8.88e-21
C5368 a_n2661_42834# a_5841_44260# 5.31e-20
C5369 a_19963_31679# a_13887_32519# 0.051213f
C5370 a_5385_46902# VDD 0.203316f
C5371 a_18494_42460# a_n97_42460# 2.68e-19
C5372 a_n2293_42834# a_6031_43396# 1.5e-19
C5373 a_9313_44734# a_10729_43914# 0.001217f
C5374 a_n2017_45002# a_743_42282# 7.84646f
C5375 a_13720_44458# a_14021_43940# 8.41e-19
C5376 a_n913_45002# a_4190_30871# 0.061913f
C5377 a_3422_30871# a_22485_44484# 0.003365f
C5378 a_22315_44484# a_20512_43084# 0.004063f
C5379 a_12741_44636# a_20623_45572# 5.76e-19
C5380 a_4883_46098# a_5891_43370# 0.003161f
C5381 a_8034_45724# a_6511_45714# 0.001344f
C5382 a_768_44030# a_10440_44484# 0.002332f
C5383 a_12891_46348# a_8975_43940# 6.34e-21
C5384 a_20202_43084# a_20731_45938# 4.22e-19
C5385 a_11415_45002# a_20528_45572# 0.002765f
C5386 a_10809_44734# a_12791_45546# 3.56e-21
C5387 a_n2442_46660# a_n4318_40392# 0.023735f
C5388 a_3090_45724# a_13017_45260# 2.74e-21
C5389 a_5934_30871# a_2113_38308# 6.72e-20
C5390 a_n1630_35242# a_n2302_37690# 1.59e-19
C5391 a_21335_42336# a_21421_42336# 0.006584f
C5392 COMP_P a_6886_37412# 0.00104f
C5393 a_n1741_47186# SMPL_ON_P 0.178214f
C5394 a_n2497_47436# a_n971_45724# 0.229429f
C5395 a_n2109_47186# a_n815_47178# 0.160027f
C5396 a_n1920_47178# a_n1605_47204# 0.08571f
C5397 a_22400_42852# a_22469_39537# 0.019601f
C5398 a_3863_42891# VDD 8.63e-19
C5399 a_3065_45002# a_1755_42282# 4.51e-19
C5400 a_n913_45002# a_5337_42558# 0.006397f
C5401 a_n1533_46116# VDD 0.143145f
C5402 a_n2956_38216# a_n2946_37690# 0.004064f
C5403 a_11967_42832# a_12281_43396# 0.027232f
C5404 a_n2017_45002# a_5755_42308# 0.004115f
C5405 a_20193_45348# a_19987_42826# 0.008117f
C5406 a_5891_43370# a_5649_42852# 6.09e-19
C5407 a_9313_44734# a_21487_43396# 1.21e-19
C5408 a_1467_44172# a_1512_43396# 2.14e-20
C5409 a_3499_42826# a_n97_42460# 0.019497f
C5410 a_n2661_42282# a_n1917_43396# 4.78e-21
C5411 a_3483_46348# a_5343_44458# 0.046505f
C5412 a_4646_46812# a_7542_44172# 0.012612f
C5413 a_13259_45724# a_14180_45002# 0.04353f
C5414 a_2324_44458# a_11827_44484# 0.03555f
C5415 a_2957_45546# a_413_45260# 0.012841f
C5416 a_n755_45592# a_2274_45254# 1.63e-19
C5417 a_n357_42282# a_2382_45260# 0.025504f
C5418 a_5937_45572# a_n2661_44458# 0.061693f
C5419 a_4419_46090# a_4223_44672# 1.94e-20
C5420 a_4185_45028# a_n699_43396# 0.027874f
C5421 a_13904_45546# a_14033_45572# 0.010132f
C5422 a_n443_42852# a_n913_45002# 0.796158f
C5423 a_3090_45724# a_19006_44850# 0.001921f
C5424 a_18985_46122# a_19778_44110# 3.49e-19
C5425 a_4791_45118# a_3539_42460# 6.9e-19
C5426 a_19692_46634# a_17517_44484# 0.023737f
C5427 a_19321_45002# a_11341_43940# 0.009893f
C5428 a_13747_46662# a_15493_43940# 0.049242f
C5429 a_12549_44172# a_14021_43940# 0.150377f
C5430 a_n4209_38216# C6_P_btm 1.26e-20
C5431 a_n3565_38216# C8_P_btm 1.65e-20
C5432 a_8530_39574# VDAC_P 0.064895f
C5433 a_7754_38470# a_11206_38545# 7.39e-19
C5434 a_n3607_39392# VDD 2.79e-20
C5435 a_n2312_39304# a_n2840_46634# 0.018018f
C5436 a_n2312_40392# a_n2956_39768# 0.056063f
C5437 a_n1151_42308# a_7411_46660# 2.81e-19
C5438 a_4915_47217# a_5072_46660# 1.11e-19
C5439 a_5815_47464# a_5732_46660# 0.002408f
C5440 a_6151_47436# a_5907_46634# 9.7e-19
C5441 a_11117_47542# a_11309_47204# 5.76e-19
C5442 a_n881_46662# a_13675_47204# 0.001593f
C5443 a_n971_45724# a_6682_46987# 0.006879f
C5444 a_n237_47217# a_6755_46942# 0.073038f
C5445 a_2063_45854# a_8667_46634# 0.00593f
C5446 a_6575_47204# a_4646_46812# 1.71e-19
C5447 a_3905_42865# a_5193_42852# 0.001894f
C5448 a_2982_43646# a_15781_43660# 1.65e-20
C5449 a_19431_45546# VDD 0.342308f
C5450 a_18909_45814# START 2.56e-21
C5451 a_20974_43370# a_21487_43396# 0.03755f
C5452 a_21381_43940# a_13467_32519# 0.002377f
C5453 a_n2293_43922# a_3318_42354# 4.38e-20
C5454 a_5891_43370# a_7963_42308# 0.036306f
C5455 a_15682_43940# a_16795_42852# 7.6e-20
C5456 a_19963_31679# EN_VIN_BSTR_N 0.004167f
C5457 a_19479_31679# a_19864_35138# 6.24e-22
C5458 a_2711_45572# a_7640_43914# 3.03e-20
C5459 a_5691_45260# a_5205_44484# 9.01e-20
C5460 a_8049_45260# a_22959_44484# 5.34e-19
C5461 a_3537_45260# a_8953_45002# 2.96e-19
C5462 a_18597_46090# a_19164_43230# 2.45e-21
C5463 a_768_44030# a_1847_42826# 4.92e-19
C5464 a_n2956_39304# a_n3674_39768# 0.02324f
C5465 a_n2956_38680# a_n4318_39768# 0.023254f
C5466 a_15903_45785# a_11691_44458# 4.76e-21
C5467 a_16855_45546# a_11827_44484# 7.23e-23
C5468 a_18479_47436# a_20922_43172# 9.43e-20
C5469 a_n443_42852# a_556_44484# 4.78e-20
C5470 a_11322_45546# a_8975_43940# 2.88e-19
C5471 a_3503_45724# a_n2661_43922# 5.64e-21
C5472 a_526_44458# a_2675_43914# 0.03283f
C5473 a_5111_44636# a_7229_43940# 4.19e-21
C5474 a_3232_43370# a_6431_45366# 0.005731f
C5475 a_15227_44166# a_2982_43646# 8.62e-20
C5476 a_n2017_45002# a_626_44172# 1.24e-20
C5477 a_10903_43370# a_10807_43548# 0.193971f
C5478 a_n913_45002# a_375_42282# 0.01541f
C5479 a_13507_46334# a_18083_42858# 1.81e-19
C5480 a_n1613_43370# a_8605_42826# 0.159791f
C5481 a_4185_45028# a_22959_43948# 0.014665f
C5482 a_3483_46348# a_9801_44260# 0.002837f
C5483 a_11599_46634# a_19553_46090# 0.021903f
C5484 a_n237_47217# a_8049_45260# 0.109887f
C5485 a_6755_46942# a_8270_45546# 0.045608f
C5486 a_10428_46928# a_11186_47026# 0.055625f
C5487 a_10467_46802# a_10768_47026# 9.73e-19
C5488 a_10249_46116# a_10384_47026# 5.86e-19
C5489 a_n881_46662# a_167_45260# 0.108232f
C5490 a_n1613_43370# a_2521_46116# 8.1e-20
C5491 a_16327_47482# a_17715_44484# 0.03083f
C5492 a_16763_47508# a_15682_46116# 0.001945f
C5493 a_13747_46662# a_12741_44636# 0.099721f
C5494 a_4791_45118# a_526_44458# 0.042209f
C5495 a_n443_46116# a_2981_46116# 0.017561f
C5496 a_1983_46706# a_765_45546# 9.01e-19
C5497 a_19594_46812# a_11415_45002# 2.74e-20
C5498 a_n1435_47204# a_6945_45028# 0.030745f
C5499 a_10227_46804# a_15015_46420# 0.287571f
C5500 a_4883_46098# a_9290_44172# 0.055265f
C5501 a_19328_44172# a_19511_42282# 2.58e-21
C5502 a_5649_42852# a_17595_43084# 9.42e-21
C5503 a_4190_30871# a_20922_43172# 8.66e-20
C5504 a_21259_43561# a_21356_42826# 3.61e-19
C5505 a_11341_43940# a_17531_42308# 2.85e-21
C5506 a_15493_43940# a_4958_30871# 4.56e-21
C5507 a_13076_44458# VDD 0.180665f
C5508 a_4361_42308# a_17333_42852# 3.75e-20
C5509 a_1209_43370# a_1606_42308# 1.26e-20
C5510 a_n1557_42282# a_n327_42558# 0.001953f
C5511 a_3080_42308# a_n1630_35242# 0.032975f
C5512 a_743_42282# a_19164_43230# 5.07e-20
C5513 a_14209_32519# a_5342_30871# 0.028644f
C5514 a_n2661_45546# a_3080_42308# 0.155045f
C5515 a_11691_44458# a_n2661_44458# 0.021716f
C5516 a_6171_45002# a_14673_44172# 6.91e-20
C5517 a_19479_31679# a_22959_44484# 0.001721f
C5518 SMPL_ON_N a_13258_32519# 0.030848f
C5519 a_9290_44172# a_5649_42852# 3.77e-19
C5520 a_12549_44172# a_15764_42576# 7.49e-20
C5521 a_n863_45724# a_1568_43370# 0.202455f
C5522 a_9482_43914# a_13468_44734# 0.00165f
C5523 a_11823_42460# a_12603_44260# 2.91e-20
C5524 a_1423_45028# a_9313_44734# 0.241551f
C5525 a_3090_45724# a_10793_43218# 9.54e-20
C5526 a_1138_42852# a_791_42968# 0.100783f
C5527 a_13507_46334# a_22775_42308# 0.022177f
C5528 a_3699_46634# a_n755_45592# 3.16e-20
C5529 a_2107_46812# a_n443_42852# 1.15e-19
C5530 a_4646_46812# a_n2661_45546# 7e-20
C5531 a_12891_46348# a_10193_42453# 1.13e-20
C5532 a_n2497_47436# a_n2293_45010# 0.233882f
C5533 a_16327_47482# a_15861_45028# 0.030602f
C5534 a_2609_46660# a_2957_45546# 7.62e-19
C5535 a_n2661_46634# a_6194_45824# 1.76e-20
C5536 a_8270_45546# a_8049_45260# 0.321896f
C5537 a_n2293_46098# a_2521_46116# 1.28e-20
C5538 a_376_46348# a_472_46348# 0.318161f
C5539 a_16388_46812# a_17957_46116# 0.140894f
C5540 a_13885_46660# a_6945_45028# 7.75e-21
C5541 a_12925_46660# a_10809_44734# 7.99e-21
C5542 a_10227_46804# a_16333_45814# 3.14e-19
C5543 a_5649_42852# a_21887_42336# 0.017243f
C5544 a_13678_32519# a_21613_42308# 0.024855f
C5545 a_13887_32519# a_7174_31319# 0.003259f
C5546 a_13467_32519# a_21125_42558# 1.91e-19
C5547 a_4361_42308# a_18997_42308# 1.34e-19
C5548 a_10796_42968# a_5742_30871# 0.003276f
C5549 a_10835_43094# a_11551_42558# 4.09e-19
C5550 a_10341_42308# a_10533_42308# 0.035479f
C5551 a_10922_42852# a_10723_42308# 0.001007f
C5552 a_10991_42826# a_11323_42473# 1.78e-19
C5553 a_10555_44260# CLK 9.69e-20
C5554 a_n356_44636# a_n809_44244# 0.00336f
C5555 a_n2661_44458# a_8333_44056# 4.4e-20
C5556 a_7499_43078# a_7871_42858# 0.146369f
C5557 a_742_44458# a_3499_42826# 4.13e-19
C5558 a_16147_45260# a_17499_43370# 5.95e-20
C5559 a_8199_44636# a_8685_42308# 0.114007f
C5560 a_8953_45546# a_8337_42558# 1.56e-19
C5561 a_n881_46662# DATA[4] 0.087677f
C5562 a_12891_46348# VDD 1.01428f
C5563 a_3537_45260# a_3626_43646# 0.002395f
C5564 a_7989_47542# DATA[3] 2.61e-19
C5565 a_11691_44458# a_18451_43940# 0.001358f
C5566 a_18911_45144# a_15493_43940# 2.89e-20
C5567 a_18184_42460# a_11341_43940# 0.029749f
C5568 a_11827_44484# a_19862_44208# 0.015537f
C5569 a_4185_45028# a_11551_42558# 8.71e-20
C5570 a_n1925_42282# a_n3674_38216# 0.004354f
C5571 a_n357_42282# a_1709_42852# 5.74e-19
C5572 a_2711_45572# a_16414_43172# 3.78e-19
C5573 a_11453_44696# a_11691_44458# 0.035893f
C5574 a_9823_46155# a_2711_45572# 5.98e-20
C5575 a_n2956_38680# a_n2956_38216# 0.10753f
C5576 a_5937_45572# a_5907_45546# 0.104991f
C5577 a_6419_46155# a_6598_45938# 1.5e-19
C5578 a_4646_46812# a_5205_44484# 0.094488f
C5579 a_5385_46902# a_5691_45260# 3.11e-22
C5580 a_5275_47026# a_3537_45260# 7.68e-22
C5581 a_1123_46634# a_626_44172# 7.29e-21
C5582 a_768_44030# a_13490_45394# 1.56e-19
C5583 a_3483_46348# a_4880_45572# 4.49e-19
C5584 a_19692_46634# a_19256_45572# 2.88e-19
C5585 a_19466_46812# a_18596_45572# 7.53e-21
C5586 a_5732_46660# a_5147_45002# 5.29e-20
C5587 a_n1151_42308# a_n2012_44484# 9.03e-20
C5588 a_7715_46873# a_413_45260# 5.62e-20
C5589 a_6755_46942# a_n2017_45002# 1.28e-20
C5590 a_4520_42826# VDD 0.142755f
C5591 a_n3674_38216# a_n4334_38528# 2.59e-19
C5592 a_5742_30871# a_4958_30871# 0.032374f
C5593 a_8515_42308# a_7174_31319# 4.88e-21
C5594 a_n3674_38680# a_n2946_38778# 4.03e-21
C5595 a_15959_42545# a_15890_42674# 0.209641f
C5596 a_n2661_43922# a_6765_43638# 4.58e-22
C5597 a_n2661_42834# a_6547_43396# 2.31e-19
C5598 a_5147_45002# a_5193_42852# 4.91e-21
C5599 a_13249_42308# a_13070_42354# 0.141799f
C5600 a_2711_45572# a_7174_31319# 0.008877f
C5601 a_805_46414# VDD 0.154663f
C5602 a_20512_43084# a_19319_43548# 1.25e-19
C5603 a_21076_30879# VREF 0.417978f
C5604 a_11823_42460# a_13657_42558# 0.009593f
C5605 a_14539_43914# a_15781_43660# 1.8e-20
C5606 a_n913_45002# a_14635_42282# 0.332583f
C5607 a_n1059_45260# a_15785_43172# 3.54e-19
C5608 a_3422_30871# a_14401_32519# 0.096501f
C5609 a_2998_44172# a_2455_43940# 1.95e-19
C5610 a_2889_44172# a_3052_44056# 0.004767f
C5611 a_2675_43914# a_3353_43940# 0.011812f
C5612 a_n356_44636# a_14955_43396# 5.49e-21
C5613 a_5891_43370# a_8685_43396# 0.145735f
C5614 a_2324_44458# a_15595_45028# 0.04743f
C5615 a_2711_45572# a_10306_45572# 7.5e-19
C5616 a_8746_45002# a_10490_45724# 0.116339f
C5617 a_526_44458# a_3429_45260# 0.010386f
C5618 a_n1925_42282# a_3065_45002# 0.04956f
C5619 a_15227_44166# a_14539_43914# 0.520312f
C5620 a_3090_45724# a_18374_44850# 3.45e-19
C5621 a_10227_46804# a_15493_43396# 0.003705f
C5622 a_10193_42453# a_11322_45546# 0.024616f
C5623 a_12741_44636# a_18911_45144# 0.013476f
C5624 a_n1613_43370# a_n1287_44306# 0.003155f
C5625 a_16327_47482# a_20623_43914# 0.009946f
C5626 a_11415_45002# a_18494_42460# 0.006745f
C5627 a_768_44030# a_5244_44056# 0.167173f
C5628 a_3483_46348# a_8560_45348# 0.021507f
C5629 a_4883_46098# a_10807_43548# 2.5e-20
C5630 a_15890_42674# RST_Z 1.6e-20
C5631 a_n2109_47186# a_171_46873# 7.56e-20
C5632 a_n815_47178# a_n1925_46634# 9.48e-20
C5633 a_19787_47423# a_12465_44636# 2.07e-19
C5634 a_n4209_38502# a_n4209_37414# 0.028607f
C5635 a_n785_47204# a_n2661_46634# 0.006981f
C5636 a_n746_45260# a_n2293_46634# 0.048005f
C5637 a_4915_47217# a_13569_47204# 4.96e-19
C5638 a_6151_47436# a_768_44030# 0.096889f
C5639 a_20990_47178# a_4883_46098# 2.39e-20
C5640 a_18479_47436# a_11453_44696# 0.018416f
C5641 a_6575_47204# a_9804_47204# 3.95e-20
C5642 a_9067_47204# a_8128_46384# 4.87e-19
C5643 a_11459_47204# a_n881_46662# 0.0707f
C5644 a_4958_30871# C0_dummy_P_btm 1.65e-20
C5645 a_5742_30871# VCM 0.211981f
C5646 a_15720_42674# VDD 4.6e-19
C5647 a_n1741_47186# a_n2438_43548# 6.62e-19
C5648 a_7174_31319# EN_VIN_BSTR_N 0.051994f
C5649 a_n2661_42282# a_n1853_43023# 4.23e-20
C5650 a_5013_44260# a_5111_42852# 2.02e-21
C5651 a_9313_44734# a_17141_43172# 1.4e-19
C5652 a_n2810_45028# a_n3565_38216# 0.349341f
C5653 a_18079_43940# a_743_42282# 3.93e-21
C5654 a_13565_43940# a_9145_43396# 0.001581f
C5655 a_1756_43548# a_2982_43646# 7.54e-20
C5656 a_11322_45546# VDD 0.370908f
C5657 a_3422_30871# a_18817_42826# 1.01e-20
C5658 a_15493_43396# a_19177_43646# 0.001461f
C5659 a_18451_43940# a_4190_30871# 3.13e-19
C5660 a_n97_42460# a_6197_43396# 0.003645f
C5661 a_14021_43940# a_16977_43638# 0.005856f
C5662 a_4791_45118# a_8605_42826# 1.13e-21
C5663 a_19321_45002# a_10341_43396# 1.67e-19
C5664 a_13661_43548# a_12293_43646# 8.56e-20
C5665 a_13059_46348# a_11341_43940# 0.025185f
C5666 a_19335_46494# a_11967_42832# 4.62e-21
C5667 a_8696_44636# a_14797_45144# 7.63e-21
C5668 a_16333_45814# a_1307_43914# 6.14e-21
C5669 a_15861_45028# a_14537_43396# 2.27e-20
C5670 a_13507_46334# a_21855_43396# 0.003121f
C5671 a_3090_45724# a_5326_44056# 2.02e-19
C5672 a_n357_42282# a_5343_44458# 0.022768f
C5673 a_n443_42852# a_n2661_44458# 0.045408f
C5674 a_15765_45572# a_16751_45260# 8.52e-20
C5675 a_1823_45246# a_3600_43914# 0.016141f
C5676 a_17339_46660# a_15493_43396# 0.075223f
C5677 a_11823_42460# a_n2661_43370# 0.006541f
C5678 a_2957_45546# a_2779_44458# 6.96e-19
C5679 a_n2293_46634# a_8317_43396# 3.08e-19
C5680 a_11453_44696# a_17829_46910# 0.013408f
C5681 a_21177_47436# a_21363_46634# 2.52e-20
C5682 a_13507_46334# a_20623_46660# 0.005302f
C5683 C0_dummy_P_btm VCM 0.311452f
C5684 a_11599_46634# a_12741_44636# 0.183316f
C5685 a_2063_45854# a_5204_45822# 0.174206f
C5686 a_n237_47217# a_8953_45546# 0.090521f
C5687 RST_Z START 0.033428f
C5688 a_12549_44172# a_19692_46634# 0.491923f
C5689 VDD SINGLE_ENDED 0.210835f
C5690 a_12465_44636# a_20107_46660# 2.35e-20
C5691 a_3877_44458# a_5167_46660# 0.032716f
C5692 a_4646_46812# a_5385_46902# 0.042888f
C5693 a_4651_46660# a_4817_46660# 0.57393f
C5694 a_n1925_46634# a_6903_46660# 7.98e-20
C5695 a_n1151_42308# a_4185_45028# 7.97e-20
C5696 a_n443_46116# a_167_45260# 0.794635f
C5697 a_3785_47178# a_3483_46348# 2.62e-20
C5698 C1_N_btm VIN_N 0.39234f
C5699 a_4883_46098# a_20273_46660# 2.98e-19
C5700 C0_N_btm VREF 0.443884f
C5701 a_13747_46662# a_13607_46688# 0.168294f
C5702 a_5807_45002# a_15009_46634# 0.006271f
C5703 a_n1741_47186# a_11133_46155# 1.23e-20
C5704 a_13667_43396# a_13635_43156# 0.006368f
C5705 a_8333_44056# a_8325_42308# 1.23e-22
C5706 a_9145_43396# a_5534_30871# 2.86e-19
C5707 a_3080_42308# a_3863_42891# 9.93e-20
C5708 a_4190_30871# a_17364_32525# 1.46e-20
C5709 a_20512_43084# a_21335_42336# 1.26e-21
C5710 a_3422_30871# a_21421_42336# 5.28e-19
C5711 a_4361_42308# a_13678_32519# 0.048617f
C5712 a_13467_32519# a_5649_42852# 0.042596f
C5713 a_21259_43561# a_20749_43396# 7.22e-19
C5714 a_6171_45002# a_12607_44458# 5.85e-20
C5715 a_3232_43370# a_12883_44458# 1.44e-20
C5716 a_18175_45572# a_17517_44484# 1.07e-20
C5717 a_3090_45724# a_10083_42826# 0.005497f
C5718 a_9290_44172# a_8685_43396# 0.207262f
C5719 a_8199_44636# a_9803_43646# 0.009804f
C5720 a_8953_45002# a_8701_44490# 0.005993f
C5721 a_8191_45002# a_5883_43914# 4.94e-22
C5722 a_375_42282# a_n2661_44458# 0.025194f
C5723 a_526_44458# a_1209_43370# 0.057216f
C5724 a_12861_44030# a_13070_42354# 2.94e-20
C5725 a_6755_46942# a_13759_46122# 9.15e-19
C5726 a_20273_46660# a_21188_46660# 0.118759f
C5727 a_20107_46660# a_20528_46660# 0.083408f
C5728 a_13747_46662# a_16375_45002# 0.021583f
C5729 a_5807_45002# a_19431_46494# 1.86e-20
C5730 a_4915_47217# a_11823_42460# 0.016758f
C5731 a_6151_47436# a_11652_45724# 9.87e-21
C5732 a_8270_45546# a_8953_45546# 1.06716f
C5733 a_n881_46662# a_n863_45724# 0.023273f
C5734 a_n1613_43370# a_n452_45724# 6.53e-20
C5735 a_11453_44696# a_n443_42852# 4.16e-20
C5736 a_3090_45724# a_3483_46348# 0.060766f
C5737 a_9313_45822# a_8568_45546# 0.002981f
C5738 a_743_42282# a_4169_42308# 4.3e-19
C5739 a_13887_32519# a_5932_42308# 0.003117f
C5740 a_4520_42826# a_n784_42308# 4.32e-21
C5741 a_16409_43396# a_15803_42450# 9.67e-20
C5742 a_4361_42308# a_6123_31319# 0.065399f
C5743 a_16243_43396# a_15890_42674# 1.41e-20
C5744 a_7281_43914# VDD 0.198809f
C5745 a_18249_42858# a_18695_43230# 2.28e-19
C5746 a_5129_47502# DATA[2] 8.34e-20
C5747 a_10193_42453# a_16409_43396# 2.72e-19
C5748 a_n356_44636# a_n2661_42834# 0.024765f
C5749 a_n1655_44484# a_n2661_43922# 6.56e-19
C5750 a_n863_45724# a_133_43172# 7.15e-19
C5751 SMPL_ON_N a_22609_37990# 2.01e-20
C5752 a_3065_45002# a_3737_43940# 0.005754f
C5753 a_12607_44458# a_14673_44172# 2.97e-21
C5754 a_18114_32519# a_21398_44850# 4.06e-20
C5755 a_1307_43914# a_15493_43396# 2.1e-19
C5756 a_19963_31679# a_14401_32519# 0.053905f
C5757 a_4915_47217# DATA[3] 0.07179f
C5758 a_7903_47542# VDD 0.202868f
C5759 a_11823_42460# a_15681_43442# 6.78e-20
C5760 a_13556_45296# a_11341_43940# 0.001133f
C5761 a_10951_45334# a_10555_44260# 5.79e-20
C5762 a_9823_46155# a_10037_46155# 0.005572f
C5763 a_n1853_46287# a_n1079_45724# 0.02186f
C5764 a_n1991_46122# a_n2293_45546# 1.19e-19
C5765 a_765_45546# a_6194_45824# 9.06e-22
C5766 a_15368_46634# a_13904_45546# 8.27e-21
C5767 a_8270_45546# a_8791_45572# 9.56e-20
C5768 a_768_44030# a_5111_44636# 0.154519f
C5769 a_21588_30879# en_comp 4.44e-19
C5770 a_9313_45822# a_n2661_43370# 8.9e-20
C5771 a_13759_46122# a_8049_45260# 0.002564f
C5772 a_11133_46155# a_10586_45546# 0.006738f
C5773 a_n901_46420# a_n2661_45546# 1.05e-19
C5774 a_13747_46662# a_413_45260# 3.67e-20
C5775 a_11309_47204# a_3232_43370# 9.11e-20
C5776 a_n2293_46634# a_n2109_45247# 0.016559f
C5777 a_n2661_46634# a_n913_45002# 8.11e-21
C5778 a_n2442_46660# a_n2017_45002# 1.18e-21
C5779 a_n881_46662# a_8191_45002# 2.82e-21
C5780 a_2107_46812# a_2437_43646# 0.185914f
C5781 a_n2293_46098# a_n452_45724# 0.007729f
C5782 a_16409_43396# VDD 0.250832f
C5783 a_6761_42308# a_6123_31319# 0.187371f
C5784 a_1606_42308# a_14456_42282# 3.31e-20
C5785 a_3232_43370# a_3935_42891# 2.51e-20
C5786 a_3537_45260# a_8037_42858# 0.010068f
C5787 a_15368_46634# CLK 5.78e-20
C5788 a_n357_42282# a_12563_42308# 9.02e-20
C5789 a_n913_45002# a_14543_43071# 0.036401f
C5790 a_n1059_45260# a_5534_30871# 0.025423f
C5791 a_n2017_45002# a_15279_43071# 0.002198f
C5792 a_11691_44458# a_9145_43396# 4.24e-19
C5793 a_11827_44484# a_14579_43548# 9.5e-23
C5794 a_18184_42460# a_10341_43396# 0.034231f
C5795 a_20835_44721# a_20623_43914# 2.27e-19
C5796 a_20640_44752# a_21115_43940# 7.54e-19
C5797 a_19279_43940# a_20269_44172# 0.002186f
C5798 a_20679_44626# a_20935_43940# 7.96e-20
C5799 a_20820_30879# a_22521_40055# 1.31e-20
C5800 a_13259_45724# a_18057_42282# 4.22e-19
C5801 a_19615_44636# a_15493_43940# 4.39e-21
C5802 a_14673_44172# a_14761_44260# 1.45e-19
C5803 a_n2661_42834# a_9165_43940# 3.03e-20
C5804 a_n699_43396# a_648_43396# 3.48e-19
C5805 a_453_43940# a_261_44278# 5.76e-19
C5806 a_18579_44172# a_15493_43396# 0.070538f
C5807 a_21076_30879# a_22521_40599# 7.82e-20
C5808 a_5663_43940# a_6453_43914# 0.017005f
C5809 a_1115_44172# a_1525_44260# 0.007617f
C5810 a_5495_43940# a_7281_43914# 1.28e-20
C5811 a_12359_47026# VDD 0.142103f
C5812 a_n443_42852# a_8325_42308# 0.001008f
C5813 a_5111_44636# a_5755_42852# 0.002818f
C5814 a_20075_46420# a_20107_45572# 0.001614f
C5815 a_13351_46090# a_3357_43084# 3.73e-21
C5816 a_8199_44636# a_n913_45002# 0.018004f
C5817 a_5937_45572# a_n1059_45260# 2.49e-20
C5818 a_8953_45546# a_n2017_45002# 0.080521f
C5819 a_3503_45724# a_3638_45822# 0.008535f
C5820 a_10586_45546# a_11688_45572# 7.93e-19
C5821 a_12741_44636# a_13348_45260# 5.41e-21
C5822 a_1823_45246# a_4558_45348# 1.95e-19
C5823 a_4419_46090# a_413_45260# 7.46e-21
C5824 a_15227_44166# a_14309_45028# 8.19e-20
C5825 a_3090_45724# a_17719_45144# 0.001738f
C5826 a_2804_46116# a_2680_45002# 1.03e-20
C5827 a_3147_46376# a_2382_45260# 1.77e-20
C5828 a_768_44030# a_12829_44484# 3.4e-20
C5829 a_11415_45002# a_13777_45326# 0.021087f
C5830 a_8049_45260# a_15297_45822# 1.34e-19
C5831 a_13661_43548# a_13857_44734# 0.012574f
C5832 a_n2109_47186# a_4883_46098# 0.029241f
C5833 a_6123_31319# a_n1532_35090# 1.38e-19
C5834 a_1343_38525# a_2112_39137# 0.22564f
C5835 a_n4209_39304# a_n2216_39072# 0.001412f
C5836 a_564_42282# VDD 0.293756f
C5837 a_1606_42308# C4_N_btm 3.05e-19
C5838 a_n1741_47186# a_13507_46334# 8.99e-20
C5839 a_5932_42308# EN_VIN_BSTR_N 0.066129f
C5840 a_n4064_40160# a_n3690_38304# 3.42e-19
C5841 a_n4064_39072# a_n4251_39392# 4.37e-19
C5842 a_6491_46660# a_7903_47542# 5.79e-21
C5843 a_4915_47217# a_9313_45822# 0.366722f
C5844 a_6151_47436# a_9067_47204# 3.94e-19
C5845 a_6545_47178# a_6575_47204# 0.11927f
C5846 a_6851_47204# a_7227_47204# 0.241208f
C5847 a_4700_47436# a_n1435_47204# 2.1e-19
C5848 a_3422_30871# a_22223_43396# 2.47e-20
C5849 a_n356_44636# a_n2293_42282# 1.10197f
C5850 a_18184_42460# a_20356_42852# 0.008384f
C5851 a_18494_42460# a_20256_42852# 0.001548f
C5852 a_n913_45002# a_19511_42282# 0.120073f
C5853 a_n1059_45260# a_19647_42308# 2.95e-20
C5854 a_n2810_45572# VDD 0.557886f
C5855 a_20512_43084# a_19095_43396# 1.93e-19
C5856 a_n2293_43922# a_10922_42852# 1.19e-20
C5857 a_9313_44734# a_15567_42826# 0.01457f
C5858 a_10807_43548# a_8685_43396# 0.029811f
C5859 a_526_44458# a_8103_44636# 3.01e-21
C5860 a_17715_44484# a_n356_44636# 1.89e-21
C5861 a_8162_45546# a_8191_45002# 0.003007f
C5862 a_9049_44484# a_7229_43940# 4.55e-21
C5863 a_12741_44636# a_19615_44636# 0.001298f
C5864 a_11415_45002# a_20640_44752# 0.0058f
C5865 a_20202_43084# a_20679_44626# 0.035147f
C5866 a_8270_45546# a_9028_43914# 0.233359f
C5867 a_18175_45572# a_19256_45572# 0.102355f
C5868 a_18341_45572# a_18691_45572# 0.206455f
C5869 a_18479_45785# a_19431_45546# 0.009466f
C5870 a_16147_45260# a_18596_45572# 9.29e-20
C5871 w_11334_34010# a_14209_32519# 7.84e-19
C5872 a_5164_46348# a_n2661_43922# 8.9e-20
C5873 a_8746_45002# a_6171_45002# 0.069475f
C5874 a_10490_45724# a_3232_43370# 9.93e-20
C5875 a_n1613_43370# a_3626_43646# 1.21e-19
C5876 a_10227_46804# a_10695_43548# 2.31e-19
C5877 a_6755_46942# a_18079_43940# 2.17e-19
C5878 a_13259_45724# a_18494_42460# 1.69e-19
C5879 a_3483_46348# a_14815_43914# 0.036548f
C5880 a_n1079_45724# a_n2661_43370# 2.43e-20
C5881 a_2711_45572# a_1423_45028# 6.59e-21
C5882 w_1575_34946# a_5534_30871# 0.001804f
C5883 a_n1386_35608# a_n83_35174# 0.081924f
C5884 a_n1532_35090# EN_VIN_BSTR_P 0.340449f
C5885 VDAC_N C5_N_btm 7.72452f
C5886 a_n4251_37440# VDD 3.95e-19
C5887 a_n1925_46634# a_171_46873# 0.027689f
C5888 a_n785_47204# a_765_45546# 1.18e-19
C5889 a_12861_44030# a_14976_45028# 0.007077f
C5890 a_n1613_43370# a_5275_47026# 0.039193f
C5891 a_11599_46634# a_13607_46688# 3.8e-19
C5892 a_n743_46660# a_n2438_43548# 0.426835f
C5893 a_n2661_46634# a_2107_46812# 0.00917f
C5894 a_n1021_46688# a_n133_46660# 1.36e-19
C5895 a_13717_47436# a_15368_46634# 3.91e-20
C5896 a_3080_42308# a_4520_42826# 4.7e-19
C5897 a_n97_42460# a_10922_42852# 3.12e-20
C5898 a_19319_43548# a_18249_42858# 7.61e-19
C5899 a_2479_44172# a_1755_42282# 6.04e-21
C5900 a_11967_42832# a_11551_42558# 6.75e-19
C5901 a_9313_44734# a_20712_42282# 6.9e-20
C5902 a_3422_30871# a_5934_30871# 0.02193f
C5903 a_10341_43396# a_15868_43402# 7.33e-20
C5904 a_6431_45366# VDD 0.203167f
C5905 a_16137_43396# a_16409_43396# 0.011989f
C5906 a_16243_43396# a_16547_43609# 0.165289f
C5907 a_n1151_42308# a_n39_42308# 9.43e-20
C5908 a_n755_45592# a_1414_42308# 0.013035f
C5909 a_n2661_45546# a_5013_44260# 1.73e-19
C5910 a_2437_43646# a_n2661_44458# 0.036499f
C5911 a_15227_44166# a_17324_43396# 0.010717f
C5912 a_3090_45724# a_16664_43396# 1.05e-21
C5913 a_13059_46348# a_10341_43396# 0.014853f
C5914 a_n1613_43370# a_8649_43218# 0.001903f
C5915 a_7705_45326# a_n2661_43370# 0.00431f
C5916 a_n863_45724# a_2889_44172# 4.42e-22
C5917 a_3357_43084# a_19721_31679# 5.18e-19
C5918 a_n1059_45260# a_11691_44458# 4.15e-20
C5919 a_n2017_45002# a_20193_45348# 1.2e-20
C5920 a_6171_45002# a_14403_45348# 3.44e-19
C5921 a_n357_42282# a_453_43940# 0.027908f
C5922 a_10193_42453# a_16241_44734# 8.94e-19
C5923 a_1823_45246# a_1756_43548# 5.06e-21
C5924 a_2107_46812# a_8199_44636# 0.022874f
C5925 a_n1151_42308# a_997_45618# 9.32e-22
C5926 a_14976_45028# a_14180_46812# 1.12e-19
C5927 a_12991_46634# a_13059_46348# 0.003295f
C5928 a_13607_46688# a_13693_46688# 0.006584f
C5929 a_14084_46812# a_14543_46987# 6.64e-19
C5930 a_3090_45724# a_14513_46634# 6.29e-19
C5931 a_n743_46660# a_11133_46155# 0.006423f
C5932 a_n237_47217# a_1609_45822# 0.141985f
C5933 a_584_46384# a_n356_45724# 0.00412f
C5934 a_2063_45854# a_3503_45724# 0.002656f
C5935 a_2905_45572# a_2957_45546# 0.137248f
C5936 a_13747_46662# a_18985_46122# 0.035795f
C5937 a_5807_45002# a_19335_46494# 0.005114f
C5938 a_13759_47204# a_6945_45028# 7.25e-19
C5939 a_3699_46634# a_3483_46348# 3.01e-19
C5940 a_11599_46634# a_16375_45002# 0.407484f
C5941 a_15368_46634# a_14035_46660# 5.28e-22
C5942 a_15559_46634# a_13885_46660# 8.64e-20
C5943 a_12861_44030# a_18051_46116# 2.97e-19
C5944 a_n881_46662# a_1431_46436# 5.43e-19
C5945 a_n443_46116# a_n863_45724# 0.055503f
C5946 a_16241_44734# VDD 0.189894f
C5947 a_4190_30871# a_19273_43230# 5.82e-21
C5948 a_17595_43084# a_17333_42852# 0.057438f
C5949 a_17701_42308# a_18083_42858# 2.35e-19
C5950 a_3422_30871# a_11530_34132# 0.127528f
C5951 a_5755_42852# a_5837_43172# 0.003935f
C5952 a_n97_42460# a_17531_42308# 1.1e-21
C5953 a_21381_43940# a_21335_42336# 0.002309f
C5954 a_n2956_39768# a_n4064_40160# 0.002282f
C5955 a_n2267_44484# a_n1243_44484# 2.36e-20
C5956 a_5205_44484# a_5013_44260# 4e-20
C5957 w_11334_34010# a_19120_35138# 0.001523f
C5958 SMPL_ON_P a_n1532_35090# 4.33e-19
C5959 a_n1352_44484# a_n356_44636# 0.003615f
C5960 a_5111_44636# a_7845_44172# 0.063408f
C5961 en_comp a_n2661_42282# 0.103098f
C5962 a_n443_42852# a_9145_43396# 2.32123f
C5963 a_3232_43370# a_6453_43914# 0.001417f
C5964 a_6171_45002# a_5663_43940# 7.76e-21
C5965 a_n2661_44458# a_4181_44734# 5.47e-19
C5966 a_6545_47178# a_5205_44484# 1.89e-20
C5967 a_16388_46812# a_13259_45724# 0.030634f
C5968 a_11453_44696# a_2437_43646# 0.189184f
C5969 a_6419_46155# a_2324_44458# 2.12e-20
C5970 a_11189_46129# a_11133_46155# 0.203074f
C5971 a_5257_43370# a_5024_45822# 1.25e-19
C5972 a_3090_45724# a_n357_42282# 0.002409f
C5973 a_9290_44172# a_11387_46155# 0.008277f
C5974 a_n746_45260# a_626_44172# 0.011647f
C5975 a_n1991_46122# a_n914_46116# 1.46e-19
C5976 a_11599_46634# a_413_45260# 3.55e-19
C5977 a_12549_44172# a_18175_45572# 1.35e-20
C5978 a_196_42282# a_n1630_35242# 0.032791f
C5979 a_11229_43218# a_5742_30871# 8.46e-20
C5980 a_20922_43172# a_19511_42282# 2.35e-19
C5981 a_n784_42308# a_564_42282# 0.003938f
C5982 a_n327_42558# a_n3674_37592# 3.94e-19
C5983 a_n4318_38680# a_n2946_38778# 3.13e-20
C5984 a_18817_42826# a_7174_31319# 8.9e-21
C5985 a_n1557_42282# VDD 0.355513f
C5986 a_n913_45002# a_21259_43561# 1.9e-20
C5987 a_n1059_45260# a_4190_30871# 0.133926f
C5988 a_14537_43396# a_15095_43370# 0.019641f
C5989 a_1307_43914# a_10695_43548# 6.81e-19
C5990 a_20692_30879# a_n1630_35242# 2.27e-19
C5991 a_4223_44672# a_5829_43940# 0.037008f
C5992 a_n2661_43922# a_3499_42826# 0.001904f
C5993 a_n2661_42834# a_3820_44260# 5.39e-19
C5994 a_6171_45002# a_16243_43396# 1.07e-19
C5995 a_20447_31679# a_13678_32519# 0.051589f
C5996 a_4817_46660# VDD 0.370615f
C5997 a_18184_42460# a_n97_42460# 4.22e-19
C5998 a_9313_44734# a_10405_44172# 0.009407f
C5999 en_comp a_16823_43084# 6.51e-22
C6000 a_19479_31679# a_14209_32519# 0.051176f
C6001 a_3422_30871# a_20512_43084# 0.125955f
C6002 a_2324_44458# a_10907_45822# 0.025622f
C6003 w_11334_34010# a_17730_32519# 0.027505f
C6004 a_12861_44030# a_15433_44458# 0.002244f
C6005 a_20731_47026# a_3357_43084# 0.00277f
C6006 a_6945_45028# a_13163_45724# 3.09e-21
C6007 a_8034_45724# a_6472_45840# 1.02e-19
C6008 a_768_44030# a_10334_44484# 0.001784f
C6009 a_11133_46155# a_11136_45572# 5.62e-20
C6010 a_11309_47204# a_8975_43940# 4.06e-22
C6011 a_11415_45002# a_21188_45572# 0.009324f
C6012 a_10809_44734# a_11823_42460# 0.215753f
C6013 a_7715_46873# a_7639_45394# 2.05e-20
C6014 a_n1630_35242# a_n4064_37440# 2.18e-20
C6015 a_n1920_47178# SMPL_ON_P 0.007059f
C6016 a_n2109_47186# a_n1605_47204# 0.041602f
C6017 a_n2288_47178# a_n815_47178# 6.95e-21
C6018 a_22400_42852# a_22821_38993# 0.136515f
C6019 a_5742_30871# a_n4064_38528# 0.005505f
C6020 a_21613_42308# a_22775_42308# 0.225363f
C6021 a_1606_42308# a_8530_39574# 0.006802f
C6022 a_3065_45002# a_1606_42308# 1.43e-20
C6023 a_n913_45002# a_4921_42308# 0.169235f
C6024 a_n722_46482# VDD 1.22e-19
C6025 a_n2810_45572# a_n2302_37690# 5.35e-19
C6026 a_11827_44484# a_21671_42860# 3.44e-21
C6027 a_n2956_38216# a_n3420_37440# 0.001161f
C6028 a_2998_44172# a_2982_43646# 7.48e-19
C6029 a_16241_44734# a_16137_43396# 7.77e-20
C6030 a_n2017_45002# a_5421_42558# 0.001147f
C6031 a_5883_43914# a_7765_42852# 2.76e-21
C6032 a_8701_44490# a_8037_42858# 1.63e-21
C6033 a_20193_45348# a_19164_43230# 3.76e-21
C6034 a_6945_45028# DATA[5] 0.047689f
C6035 a_13925_46122# a_11691_44458# 3.94e-21
C6036 a_3483_46348# a_4743_44484# 6.71e-19
C6037 a_n755_45592# a_1667_45002# 0.002f
C6038 a_4646_46812# a_7281_43914# 0.021965f
C6039 a_13059_46348# a_n2293_43922# 5.13e-21
C6040 a_1848_45724# a_413_45260# 2.84e-21
C6041 a_8199_44636# a_n2661_44458# 0.069807f
C6042 a_4185_45028# a_4223_44672# 0.031094f
C6043 a_3699_46348# a_n699_43396# 1.2e-21
C6044 a_n443_42852# a_n1059_45260# 0.130036f
C6045 a_18819_46122# a_19778_44110# 5.3e-21
C6046 a_13259_45724# a_13777_45326# 0.043567f
C6047 a_18985_46122# a_18911_45144# 7.42e-22
C6048 a_n863_45724# a_3537_45260# 1.54e-20
C6049 a_n2661_45546# a_4927_45028# 0.001509f
C6050 a_4791_45118# a_3626_43646# 0.006599f
C6051 a_13661_43548# a_15493_43940# 1.28948f
C6052 a_12891_46348# a_14021_43940# 3.26e-20
C6053 a_768_44030# a_13565_44260# 7.87e-20
C6054 a_12549_44172# a_13829_44260# 4.49e-19
C6055 a_10193_42453# a_18691_45572# 6.6e-21
C6056 a_19466_46812# a_17517_44484# 1.01e-19
C6057 w_1575_34946# a_4190_30871# 0.004947f
C6058 a_n2312_40392# a_n2840_46634# 3.22e-21
C6059 a_4883_46098# a_n1925_46634# 0.030451f
C6060 a_13507_46334# a_n743_46660# 0.024694f
C6061 a_n4209_38216# C7_P_btm 1.43e-20
C6062 a_n3565_38216# C9_P_btm 1.91e-20
C6063 a_8530_39574# a_8912_37509# 0.426772f
C6064 a_7754_38470# VDAC_P 0.063714f
C6065 a_n1151_42308# a_5257_43370# 0.058425f
C6066 a_4915_47217# a_6540_46812# 1.17e-20
C6067 a_n443_46116# a_5072_46660# 3.53e-19
C6068 a_5815_47464# a_5907_46634# 0.004583f
C6069 a_4791_45118# a_5275_47026# 0.004467f
C6070 a_6491_46660# a_4817_46660# 1.23e-19
C6071 a_n881_46662# a_13569_47204# 0.001167f
C6072 a_n4251_39392# VDD 3.95e-19
C6073 a_n971_45724# a_6969_46634# 0.235123f
C6074 a_2063_45854# a_7927_46660# 0.004156f
C6075 a_n237_47217# a_10249_46116# 2.78e-20
C6076 a_6575_47204# a_3877_44458# 6.28e-20
C6077 a_n4064_39616# VCM 0.068103f
C6078 a_11453_44696# a_n2661_46634# 0.032889f
C6079 a_n4064_37440# a_n3607_37440# 7.1e-19
C6080 a_15682_43940# a_16414_43172# 3.58e-19
C6081 a_3499_42826# a_3445_43172# 2.31e-19
C6082 a_3905_42865# a_4649_42852# 0.04156f
C6083 a_18691_45572# VDD 0.191893f
C6084 a_18341_45572# START 7.1e-21
C6085 a_14401_32519# a_21487_43396# 6.94e-19
C6086 a_n2293_43922# a_2903_42308# 8.6e-20
C6087 a_5891_43370# a_6123_31319# 0.028865f
C6088 a_11341_43940# a_10991_42826# 2.93e-19
C6089 a_20974_43370# a_20556_43646# 0.076332f
C6090 en_comp a_22469_39537# 0.001226f
C6091 a_2711_45572# a_6109_44484# 3.03e-20
C6092 a_2324_44458# a_n2661_42282# 0.001316f
C6093 a_8049_45260# a_17730_32519# 3.56e-20
C6094 a_3537_45260# a_8191_45002# 0.00226f
C6095 a_768_44030# a_791_42968# 1.22e-19
C6096 a_n357_42282# a_14815_43914# 1.18e-20
C6097 a_10490_45724# a_8975_43940# 7.33e-22
C6098 a_n2956_39304# a_n4318_39768# 0.023377f
C6099 a_15599_45572# a_11691_44458# 1.35e-20
C6100 a_9290_44172# a_13483_43940# 0.005971f
C6101 a_n443_42852# a_484_44484# 3.87e-19
C6102 a_3503_45724# a_n2661_42834# 2.21e-21
C6103 a_3316_45546# a_n2661_43922# 3.15e-20
C6104 a_526_44458# a_895_43940# 0.018069f
C6105 a_n1925_42282# a_2479_44172# 3.15e-21
C6106 a_3232_43370# a_6171_45002# 0.314056f
C6107 a_4927_45028# a_5205_44484# 9.25e-21
C6108 a_5147_45002# a_7229_43940# 1.65e-22
C6109 a_5691_45260# a_6431_45366# 0.005044f
C6110 a_10903_43370# a_10949_43914# 0.451961f
C6111 a_n1059_45260# a_375_42282# 0.0165f
C6112 a_n1613_43370# a_8037_42858# 0.047354f
C6113 a_4185_45028# a_15493_43940# 0.039364f
C6114 a_13507_46334# a_17701_42308# 7.88e-21
C6115 a_11599_46634# a_18985_46122# 0.570252f
C6116 a_n237_47217# a_8781_46436# 5.45e-19
C6117 a_10554_47026# a_10384_47026# 2.6e-19
C6118 a_10428_46928# a_10768_47026# 0.027606f
C6119 a_6755_46942# a_8189_46660# 0.002345f
C6120 a_10249_46116# a_8270_45546# 1.06e-19
C6121 a_n1613_43370# a_167_45260# 1.05e-19
C6122 a_11453_44696# a_8199_44636# 3.39e-19
C6123 a_16327_47482# a_17583_46090# 1.09e-19
C6124 a_16023_47582# a_15682_46116# 0.001021f
C6125 a_13661_43548# a_12741_44636# 0.13948f
C6126 a_n881_46662# a_2202_46116# 0.051959f
C6127 a_n1741_47186# a_10586_45546# 3.67e-20
C6128 a_4700_47436# a_526_44458# 1.71e-21
C6129 a_4007_47204# a_n1925_42282# 8.11e-20
C6130 a_2107_46812# a_765_45546# 0.001701f
C6131 a_19321_45002# a_11415_45002# 0.065361f
C6132 a_13717_47436# a_20708_46348# 5.9e-22
C6133 a_13381_47204# a_6945_45028# 0.006113f
C6134 a_12861_44030# a_19900_46494# 4.29e-21
C6135 a_10227_46804# a_14275_46494# 0.18614f
C6136 a_4883_46098# a_10355_46116# 0.23167f
C6137 a_5649_42852# a_16795_42852# 4.02e-21
C6138 a_4190_30871# a_19987_42826# 3.95e-19
C6139 a_12883_44458# VDD 0.263743f
C6140 a_3422_30871# a_7754_40130# 4.49e-20
C6141 a_19095_43396# a_18249_42858# 6.34e-19
C6142 a_4361_42308# a_18083_42858# 2.01e-19
C6143 a_n1557_42282# a_n784_42308# 0.058812f
C6144 a_9145_43396# a_14635_42282# 3.74e-20
C6145 a_743_42282# a_19339_43156# 2.4e-20
C6146 a_n755_45592# a_n1190_43762# 2.34e-20
C6147 a_375_42282# a_484_44484# 8.95e-19
C6148 a_n2661_45546# a_4699_43561# 0.013733f
C6149 a_526_44458# a_10149_43396# 0.003062f
C6150 a_1307_43914# a_3363_44484# 5.2e-19
C6151 a_3357_43084# a_22591_44484# 7.11e-20
C6152 a_19479_31679# a_17730_32519# 0.052745f
C6153 a_12549_44172# a_15486_42560# 1.17e-21
C6154 a_n863_45724# a_1049_43396# 1.03e-19
C6155 a_9482_43914# a_13213_44734# 0.003145f
C6156 a_13556_45296# a_n2293_43922# 1.07e-20
C6157 a_3090_45724# a_10553_43218# 8.81e-20
C6158 a_11823_42460# a_12495_44260# 9.96e-20
C6159 a_n2312_38680# a_5934_30871# 4.54e-21
C6160 a_1138_42852# a_685_42968# 6.59e-20
C6161 a_13507_46334# a_21613_42308# 0.035917f
C6162 a_22591_45572# a_22485_44484# 1.77e-19
C6163 a_10227_46804# a_15765_45572# 4.04e-19
C6164 a_948_46660# a_n443_42852# 2.59e-20
C6165 a_2959_46660# a_n755_45592# 2.79e-21
C6166 a_1123_46634# a_1609_45822# 8.43e-20
C6167 a_n743_46660# a_603_45572# 1.47e-19
C6168 a_3877_44458# a_n2661_45546# 0.026409f
C6169 a_11309_47204# a_10193_42453# 0.006435f
C6170 a_n881_46662# a_11823_42460# 0.036994f
C6171 a_16327_47482# a_8696_44636# 0.087584f
C6172 a_2443_46660# a_2957_45546# 3.36e-19
C6173 a_n2661_46634# a_5907_45546# 7.09e-21
C6174 a_8189_46660# a_8049_45260# 2.51e-20
C6175 a_8270_45546# a_8781_46436# 2.13e-19
C6176 a_768_44030# a_9049_44484# 0.006069f
C6177 a_n2293_46098# a_167_45260# 0.086636f
C6178 a_n1076_46494# a_472_46348# 0.001137f
C6179 a_12741_44636# a_4185_45028# 1.08e-20
C6180 a_n971_45724# a_3357_43084# 0.565799f
C6181 a_n2293_46634# a_3175_45822# 1.98e-19
C6182 a_16388_46812# a_18189_46348# 0.0042f
C6183 a_12513_46660# a_10809_44734# 5.68e-19
C6184 a_1799_45572# a_3316_45546# 2.21e-21
C6185 a_21855_43396# a_21613_42308# 2.52e-21
C6186 a_13678_32519# a_21887_42336# 0.012293f
C6187 a_14209_32519# a_13258_32519# 0.051594f
C6188 a_n2293_42282# a_3823_42558# 3.04e-21
C6189 a_5649_42852# a_21335_42336# 6.37e-20
C6190 a_10835_43094# a_5742_30871# 0.011953f
C6191 a_10796_42968# a_11323_42473# 8.05e-20
C6192 a_10341_42308# a_10545_42558# 0.002951f
C6193 a_1793_42852# a_1755_42282# 3.44e-19
C6194 a_3065_45002# a_3539_42460# 0.300764f
C6195 a_15861_45028# a_17486_43762# 5.8e-21
C6196 a_7499_43078# a_7227_42852# 0.126148f
C6197 a_2711_45572# a_15567_42826# 6.6e-20
C6198 a_n1925_42282# a_n2104_42282# 0.166917f
C6199 a_11827_44484# a_19478_44306# 0.002282f
C6200 a_14581_44484# a_14673_44172# 7.47e-20
C6201 a_8199_44636# a_8325_42308# 0.004591f
C6202 a_20567_45036# a_20623_43914# 4.97e-21
C6203 a_11309_47204# VDD 0.358104f
C6204 a_3537_45260# a_3540_43646# 2.04e-20
C6205 a_4185_45028# a_5742_30871# 0.062132f
C6206 a_18587_45118# a_15493_43940# 4.11e-22
C6207 a_19778_44110# a_11341_43940# 0.004296f
C6208 a_18184_42460# a_21115_43940# 1.01e-21
C6209 a_21359_45002# a_19862_44208# 0.001254f
C6210 a_n357_42282# a_945_42968# 4.86e-19
C6211 a_n913_45002# a_6452_43396# 1.57e-20
C6212 a_n881_46662# DATA[3] 0.001196f
C6213 a_16388_46812# a_17478_45572# 5.42e-21
C6214 a_13059_46348# a_16020_45572# 2.07e-20
C6215 a_15227_44166# a_18799_45938# 7.44e-21
C6216 a_n2956_39304# a_n2956_38216# 0.05012f
C6217 a_5204_45822# a_3775_45552# 9.09e-22
C6218 a_6419_46155# a_6667_45809# 6.84e-19
C6219 a_5937_45572# a_5263_45724# 0.002746f
C6220 a_4817_46660# a_5691_45260# 8.09e-19
C6221 a_3877_44458# a_5205_44484# 5.39e-21
C6222 a_4915_47217# a_14539_43914# 1.6e-19
C6223 a_7411_46660# a_413_45260# 2.01e-20
C6224 a_9569_46155# a_2711_45572# 6.07e-20
C6225 a_12891_46348# a_13711_45394# 0.003687f
C6226 a_3483_46348# a_4808_45572# 3.56e-19
C6227 a_765_45546# a_15903_45785# 2.27e-20
C6228 a_19692_46634# a_19431_45546# 5.98e-20
C6229 a_19466_46812# a_19256_45572# 0.041135f
C6230 a_n2956_38680# a_n2472_45546# 4.48e-19
C6231 a_5167_46660# a_5111_44636# 1.66e-20
C6232 a_4646_46812# a_6431_45366# 8.39e-19
C6233 a_584_46384# a_n356_44636# 0.268036f
C6234 a_3935_42891# VDD 0.096403f
C6235 a_n3674_38216# a_n4209_38502# 4.47e-20
C6236 a_5934_30871# a_7174_31319# 0.473128f
C6237 a_15803_42450# a_15890_42674# 0.07009f
C6238 a_15764_42576# a_15720_42674# 1.46e-19
C6239 a_n3674_38680# a_n3420_38528# 0.07337f
C6240 a_n3674_37592# a_n4064_39072# 0.019349f
C6241 a_n2293_43922# a_6293_42852# 9.77e-21
C6242 a_n2661_42834# a_6765_43638# 4.91e-21
C6243 a_n2661_43922# a_6197_43396# 1.61e-20
C6244 a_21076_30879# VIN_N 0.068195f
C6245 a_13249_42308# a_12563_42308# 1.64e-19
C6246 a_2711_45572# a_20712_42282# 4.18e-19
C6247 a_472_46348# VDD 0.706547f
C6248 a_20820_30879# VCM 0.05604f
C6249 a_11750_44172# a_12429_44172# 1.03e-20
C6250 a_3537_45260# a_7309_42852# 4.49e-19
C6251 a_11823_42460# a_13333_42558# 0.003508f
C6252 a_14539_43914# a_15681_43442# 4.94e-20
C6253 a_10193_42453# a_15890_42674# 8.41e-20
C6254 a_n913_45002# a_13291_42460# 0.070562f
C6255 a_n1059_45260# a_14635_42282# 0.063373f
C6256 a_20980_44850# a_20974_43370# 4.87e-21
C6257 a_3422_30871# a_21381_43940# 0.006676f
C6258 a_2998_44172# a_2253_43940# 2.08e-19
C6259 a_2675_43914# a_3052_44056# 7.61e-19
C6260 a_n2956_38216# a_n3565_39304# 0.02162f
C6261 a_20193_45348# a_14209_32519# 5.6e-19
C6262 a_n443_46116# a_2455_43940# 0.010179f
C6263 w_11334_34010# a_17538_32519# 0.036508f
C6264 a_2324_44458# a_15415_45028# 0.03757f
C6265 a_2711_45572# a_10216_45572# 9.36e-19
C6266 a_10193_42453# a_10490_45724# 0.062365f
C6267 a_526_44458# a_3065_45002# 0.138202f
C6268 a_1823_45246# a_n2661_43370# 0.112095f
C6269 a_4185_45028# a_n2293_42834# 0.022725f
C6270 a_3090_45724# a_18443_44721# 3.2e-20
C6271 a_15227_44166# a_16112_44458# 0.073746f
C6272 a_765_45546# a_n2661_44458# 1.25e-21
C6273 a_12741_44636# a_18587_45118# 0.005591f
C6274 a_n1613_43370# a_n1453_44318# 9.54e-19
C6275 a_5937_45572# a_5837_45348# 2.99e-19
C6276 a_3483_46348# a_8488_45348# 0.003238f
C6277 a_11415_45002# a_18184_42460# 0.006818f
C6278 a_768_44030# a_3905_42865# 0.011432f
C6279 a_20202_43084# a_18494_42460# 0.166633f
C6280 a_4883_46098# a_10949_43914# 3.15e-21
C6281 a_16327_47482# a_20365_43914# 0.007136f
C6282 a_15959_42545# RST_Z 3.5e-20
C6283 a_n2497_47436# a_33_46660# 6.33e-21
C6284 a_22465_38105# a_22705_37990# 1.35e-19
C6285 a_n971_45724# a_n2293_46634# 0.090091f
C6286 a_n23_47502# a_n2661_46634# 5.47e-19
C6287 a_n1151_42308# a_5807_45002# 1.52318f
C6288 a_6151_47436# a_12549_44172# 0.214024f
C6289 a_19386_47436# a_12465_44636# 2.39e-19
C6290 a_6575_47204# a_8128_46384# 0.105633f
C6291 a_9313_45822# a_n881_46662# 1.00227f
C6292 a_5742_30871# VREF_GND 0.191352f
C6293 a_4958_30871# C0_P_btm 9.29e-20
C6294 a_15890_42674# VDD 0.203548f
C6295 a_18143_47464# a_11453_44696# 0.001066f
C6296 a_21177_47436# a_13507_46334# 0.329096f
C6297 a_n1920_47178# a_n2438_43548# 1.47e-19
C6298 a_n2109_47186# a_n133_46660# 2.86e-20
C6299 a_n1741_47186# a_n743_46660# 0.017496f
C6300 a_7174_31319# a_11530_34132# 0.001307f
C6301 a_n2661_42282# a_n2157_42858# 4.07e-20
C6302 a_9313_44734# a_16877_43172# 5.07e-19
C6303 a_5244_44056# a_5111_42852# 9.76e-21
C6304 a_742_44458# a_2903_42308# 0.0077f
C6305 a_10490_45724# VDD 0.162001f
C6306 a_n97_42460# a_6293_42852# 0.018467f
C6307 a_1568_43370# a_2982_43646# 0.002246f
C6308 a_n2956_37592# a_n4209_38216# 0.104159f
C6309 a_3422_30871# a_18249_42858# 1.45e-20
C6310 a_12429_44172# a_4361_42308# 1.84e-21
C6311 a_14021_43940# a_16409_43396# 0.025204f
C6312 a_2063_45854# a_10341_42308# 6.99e-21
C6313 a_8696_44636# a_14537_43396# 0.024289f
C6314 a_3090_45724# a_5025_43940# 4.03e-19
C6315 a_n357_42282# a_4743_44484# 5.15e-21
C6316 a_15765_45572# a_1307_43914# 9.23e-20
C6317 a_15903_45785# a_16751_45260# 2.12e-20
C6318 a_13507_46334# a_4361_42308# 0.040714f
C6319 a_1823_45246# a_2998_44172# 0.062531f
C6320 a_5066_45546# a_n2661_43922# 4.26e-20
C6321 a_n755_45592# a_n699_43396# 0.185444f
C6322 a_n2293_46634# a_8229_43396# 2.24e-19
C6323 VDD START 0.114358f
C6324 a_13507_46334# a_20841_46902# 0.005806f
C6325 C0_P_btm VCM 0.717283f
C6326 a_n971_45724# a_9625_46129# 2.11e-20
C6327 a_2063_45854# a_5164_46348# 0.022664f
C6328 a_n237_47217# a_5937_45572# 0.08715f
C6329 a_12549_44172# a_19466_46812# 1.6e-19
C6330 a_11453_44696# a_765_45546# 0.010973f
C6331 a_3877_44458# a_5385_46902# 0.021989f
C6332 a_4646_46812# a_4817_46660# 0.588038f
C6333 a_4651_46660# a_4955_46873# 0.140348f
C6334 a_n1925_46634# a_6682_46660# 1.03e-19
C6335 a_2905_45572# a_4419_46090# 1.32e-19
C6336 C0_N_btm VIN_N 0.529671f
C6337 a_n443_46116# a_2202_46116# 7.93e-21
C6338 a_13747_46662# a_12816_46660# 2.17e-21
C6339 a_5807_45002# a_14084_46812# 0.006112f
C6340 a_n2661_46634# a_10384_47026# 1.14e-19
C6341 a_n1741_47186# a_11189_46129# 4.54e-19
C6342 a_16327_47482# a_20885_46660# 8.54e-21
C6343 a_4883_46098# a_20411_46873# 0.012008f
C6344 a_15095_43370# a_12379_42858# 1.62e-21
C6345 a_10903_45394# CLK 0.001362f
C6346 a_17730_32519# a_13258_32519# 0.05785f
C6347 a_3422_30871# a_21125_42558# 2.49e-20
C6348 a_4361_42308# a_21855_43396# 0.167446f
C6349 a_13467_32519# a_13678_32519# 10.9526f
C6350 a_10341_43396# a_10991_42826# 7.08e-20
C6351 a_3232_43370# a_12607_44458# 1.04e-20
C6352 a_16147_45260# a_17517_44484# 8.68e-20
C6353 a_3090_45724# a_8952_43230# 1.36e-19
C6354 a_8199_44636# a_9145_43396# 0.020485f
C6355 a_6171_45002# a_8975_43940# 0.175346f
C6356 a_526_44458# a_458_43396# 0.085782f
C6357 w_1575_34946# a_n3420_37984# 3.98e-19
C6358 a_9863_46634# a_2324_44458# 2.26e-21
C6359 a_n881_46662# a_n1079_45724# 0.002262f
C6360 a_13059_46348# a_11415_45002# 0.225168f
C6361 a_20107_46660# a_22000_46634# 3.29e-20
C6362 a_20841_46902# a_20623_46660# 0.209641f
C6363 a_20273_46660# a_21363_46634# 0.042415f
C6364 a_n743_46660# a_10586_45546# 0.018104f
C6365 a_6755_46942# a_13351_46090# 3.38e-19
C6366 a_13661_43548# a_16375_45002# 0.003429f
C6367 a_5807_45002# a_19240_46482# 0.002625f
C6368 a_8270_45546# a_5937_45572# 0.29626f
C6369 a_n1613_43370# a_n863_45724# 0.027265f
C6370 a_765_45546# a_17639_46660# 0.094916f
C6371 a_17339_46660# a_18280_46660# 0.002515f
C6372 a_3090_45724# a_3147_46376# 0.010392f
C6373 a_9067_47204# a_9049_44484# 3.2e-20
C6374 a_19321_45002# a_13259_45724# 5.11e-20
C6375 a_6453_43914# VDD 0.194953f
C6376 a_743_42282# a_3905_42308# 3.67e-19
C6377 a_16547_43609# a_15803_42450# 1.5e-20
C6378 a_16243_43396# a_15959_42545# 6.33e-20
C6379 a_16409_43396# a_15764_42576# 6.83e-20
C6380 a_4361_42308# a_7227_42308# 0.01047f
C6381 a_16137_43396# a_15890_42674# 2.67e-21
C6382 a_13467_32519# a_6123_31319# 2.49e-19
C6383 a_10341_43396# a_17303_42282# 1.21e-20
C6384 a_16414_43172# a_16245_42852# 0.08213f
C6385 a_18249_42858# a_18504_43218# 0.05936f
C6386 a_791_42968# a_1067_42314# 2.04e-19
C6387 a_4915_47217# DATA[2] 9.44e-19
C6388 a_n1821_44484# a_n2661_43922# 0.001334f
C6389 a_n1655_44484# a_n2661_42834# 5.04e-19
C6390 a_10775_45002# a_10555_44260# 2.44e-20
C6391 a_2382_45260# a_3992_43940# 4.5e-19
C6392 a_13076_44458# a_13296_44484# 0.009965f
C6393 a_12607_44458# a_14581_44484# 3.05e-21
C6394 a_19479_31679# a_17538_32519# 0.051112f
C6395 a_n443_46116# DATA[3] 1.57e-20
C6396 a_n2661_43370# a_n3674_39768# 0.144159f
C6397 a_7227_47204# VDD 0.430714f
C6398 a_8375_44464# a_8783_44734# 5.23e-21
C6399 a_700_44734# a_556_44484# 6.84e-19
C6400 a_9482_43914# a_11341_43940# 0.037822f
C6401 a_9823_46155# a_9751_46155# 6.64e-19
C6402 a_n1853_46287# a_n2293_45546# 8.68e-20
C6403 a_765_45546# a_5907_45546# 6.13e-21
C6404 a_768_44030# a_5147_45002# 0.191082f
C6405 a_n2312_38680# a_n2661_45010# 1.97e-21
C6406 a_11453_44696# a_16751_45260# 0.002984f
C6407 a_11189_46129# a_10586_45546# 0.028266f
C6408 a_n2157_46122# a_n1079_45724# 0.006548f
C6409 a_n1641_46494# a_n2661_45546# 7.41e-20
C6410 a_3090_45724# a_13249_42308# 0.032019f
C6411 a_13661_43548# a_413_45260# 2.4e-20
C6412 a_n2293_46634# a_n2293_45010# 0.036081f
C6413 a_n1613_43370# a_8191_45002# 2.41e-21
C6414 a_n881_46662# a_7705_45326# 3.83e-20
C6415 a_948_46660# a_2437_43646# 2.21e-20
C6416 a_4915_47217# a_14309_45028# 0.004859f
C6417 a_n2293_46098# a_n863_45724# 0.003336f
C6418 a_13351_46090# a_8049_45260# 0.002917f
C6419 a_16547_43609# VDD 0.31275f
C6420 a_6761_42308# a_7227_42308# 0.173849f
C6421 a_5932_42308# a_5934_30871# 1.37963f
C6422 a_1606_42308# a_13575_42558# 1.77e-20
C6423 a_3232_43370# a_3681_42891# 0.005411f
C6424 a_3537_45260# a_7765_42852# 2.41e-19
C6425 a_n913_45002# a_13460_43230# 0.04239f
C6426 a_n1059_45260# a_14543_43071# 0.002239f
C6427 a_n2017_45002# a_5534_30871# 0.025363f
C6428 a_19778_44110# a_10341_43396# 1.31e-19
C6429 a_13259_45724# a_17531_42308# 0.009212f
C6430 a_20159_44458# a_11341_43940# 6.61e-20
C6431 a_20679_44626# a_20623_43914# 0.009865f
C6432 a_20640_44752# a_20935_43940# 4.13e-20
C6433 a_14976_45028# CLK 4.29e-20
C6434 a_11967_42832# a_15493_43940# 0.299734f
C6435 a_n2661_42834# a_8487_44056# 1.89e-21
C6436 a_19279_43940# a_19862_44208# 0.012567f
C6437 a_n699_43396# a_548_43396# 2.06e-19
C6438 a_18579_44172# a_19328_44172# 0.053539f
C6439 a_1115_44172# a_1241_44260# 0.013015f
C6440 a_5495_43940# a_6453_43914# 5.83e-20
C6441 a_n1761_44111# a_n2661_42282# 5.46e-20
C6442 a_12156_46660# VDD 0.082428f
C6443 a_19692_46634# SINGLE_ENDED 4.63e-20
C6444 a_5111_44636# a_5111_42852# 0.148196f
C6445 a_n755_45592# a_5024_45822# 1.65e-20
C6446 a_5257_43370# a_4223_44672# 0.016657f
C6447 a_n2293_46634# a_9313_44734# 0.022598f
C6448 a_13925_46122# a_2437_43646# 1.99e-20
C6449 a_12594_46348# a_3357_43084# 9.87e-21
C6450 a_8199_44636# a_n1059_45260# 0.019728f
C6451 a_5937_45572# a_n2017_45002# 2.08e-20
C6452 a_3503_45724# a_3775_45552# 0.13675f
C6453 a_10586_45546# a_11136_45572# 0.006861f
C6454 a_12741_44636# a_13159_45002# 7.19e-20
C6455 a_4185_45028# a_413_45260# 0.191095f
C6456 a_n1151_42308# a_n822_43940# 3.16e-20
C6457 a_3090_45724# a_17613_45144# 1.41e-19
C6458 a_2698_46116# a_2680_45002# 2.37e-20
C6459 a_2804_46116# a_2382_45260# 1.18e-21
C6460 a_1823_45246# a_4574_45260# 3.32e-19
C6461 a_12891_46348# a_13296_44484# 3.98e-19
C6462 a_12549_44172# a_12829_44484# 3.48e-20
C6463 a_11415_45002# a_13556_45296# 0.16025f
C6464 a_8049_45260# a_15225_45822# 7.33e-20
C6465 a_n4315_30879# a_n3420_37984# 0.034791f
C6466 a_n1151_42308# a_14311_47204# 0.003307f
C6467 a_7174_31319# a_7754_40130# 0.005009f
C6468 a_n3674_37592# VDD 0.357168f
C6469 a_1606_42308# C3_N_btm 5.68e-19
C6470 a_5932_42308# a_11530_34132# 0.001408f
C6471 a_n4064_40160# a_n3565_38216# 0.02828f
C6472 a_n4064_39616# a_n4064_38528# 0.05063f
C6473 a_n3420_39072# a_n3607_39392# 8.36e-19
C6474 a_n4064_39072# a_n2302_39072# 0.250408f
C6475 a_6545_47178# a_7903_47542# 1.49e-19
C6476 a_4915_47217# a_11031_47542# 0.125943f
C6477 a_6491_46660# a_7227_47204# 0.001647f
C6478 a_6151_47436# a_6575_47204# 0.047329f
C6479 a_4007_47204# a_n1435_47204# 0.001005f
C6480 a_18184_42460# a_20256_42852# 0.01674f
C6481 a_2253_43940# a_1568_43370# 3.94e-19
C6482 a_19319_43548# a_19741_43940# 0.048788f
C6483 a_n1059_45260# a_19511_42282# 3.28e-19
C6484 a_n2017_45002# a_19647_42308# 1.94e-19
C6485 a_n2840_45546# VDD 0.302566f
C6486 a_20512_43084# a_21487_43396# 0.003816f
C6487 a_3422_30871# a_5649_42852# 0.291966f
C6488 a_n2293_43922# a_10991_42826# 2.64e-20
C6489 a_9313_44734# a_5342_30871# 0.026413f
C6490 a_1307_43914# a_8685_42308# 1.98e-21
C6491 a_10949_43914# a_8685_43396# 4.56e-21
C6492 a_18579_44172# a_20749_43396# 5.9e-20
C6493 a_19479_31679# a_22465_38105# 2.87e-19
C6494 a_20447_31679# a_22775_42308# 4.98e-21
C6495 en_comp a_19332_42282# 4.59e-20
C6496 a_526_44458# a_6298_44484# 8.53e-21
C6497 a_8049_45260# a_19721_31679# 7.57e-19
C6498 a_7499_43078# a_7229_43940# 9.29e-21
C6499 a_12741_44636# a_11967_42832# 0.004783f
C6500 a_11415_45002# a_20362_44736# 0.001672f
C6501 a_20202_43084# a_20640_44752# 0.027593f
C6502 a_8270_45546# a_8333_44056# 0.001906f
C6503 a_18341_45572# a_18909_45814# 0.170692f
C6504 a_18479_45785# a_18691_45572# 0.036486f
C6505 a_18175_45572# a_19431_45546# 0.043567f
C6506 a_16147_45260# a_19256_45572# 2.79e-20
C6507 a_n2956_39768# a_n4318_39304# 0.02353f
C6508 a_768_44030# a_4093_43548# 1.82e-19
C6509 a_16375_45002# a_18587_45118# 2.59e-20
C6510 a_10193_42453# a_6171_45002# 0.411891f
C6511 a_8746_45002# a_3232_43370# 0.439467f
C6512 a_6755_46942# a_17973_43940# 6e-19
C6513 a_n971_45724# a_743_42282# 2.96e-19
C6514 a_10227_46804# a_9803_43646# 0.003261f
C6515 a_3483_46348# a_14112_44734# 2.1e-20
C6516 a_13259_45724# a_18184_42460# 0.001266f
C6517 a_n2293_45546# a_n2661_43370# 0.131199f
C6518 a_n23_47502# a_765_45546# 1.93e-20
C6519 a_n881_46662# a_6540_46812# 3.2e-19
C6520 a_12861_44030# a_3090_45724# 0.496275f
C6521 a_13717_47436# a_14976_45028# 2.92e-20
C6522 a_n1613_43370# a_5072_46660# 0.012366f
C6523 a_n1532_35090# a_n923_35174# 0.400297f
C6524 a_n1386_35608# EN_VIN_BSTR_P 0.573134f
C6525 VDAC_N C4_N_btm 3.92765f
C6526 a_11599_46634# a_12816_46660# 6.65e-20
C6527 a_n2661_46634# a_948_46660# 0.008972f
C6528 a_14311_47204# a_14084_46812# 2.83e-19
C6529 a_n2216_37690# VDD 0.003946f
C6530 a_n1021_46688# a_n2438_43548# 0.053225f
C6531 a_n1925_46634# a_n133_46660# 0.053144f
C6532 a_4699_43561# a_4520_42826# 1.02e-19
C6533 a_3080_42308# a_3935_42891# 0.017131f
C6534 a_n97_42460# a_10991_42826# 6.43e-20
C6535 a_10341_43396# a_15231_43396# 1.63e-19
C6536 a_14579_43548# a_16823_43084# 3.51e-21
C6537 a_6171_45002# VDD 0.441339f
C6538 a_16137_43396# a_16547_43609# 0.151161f
C6539 a_9313_44734# a_20107_42308# 8.02e-20
C6540 a_584_46384# a_3823_42558# 3.7e-20
C6541 a_n1151_42308# a_n327_42308# 1.59e-19
C6542 a_n357_42282# a_1414_42308# 0.027118f
C6543 a_15227_44166# a_17499_43370# 0.021724f
C6544 a_n1613_43370# a_7309_42852# 8.11e-20
C6545 a_13249_42308# a_14815_43914# 4.82e-21
C6546 a_6709_45028# a_n2661_43370# 0.041021f
C6547 a_8191_45002# a_8704_45028# 8.88e-19
C6548 a_n863_45724# a_2675_43914# 2e-20
C6549 a_3357_43084# a_18114_32519# 8.45e-21
C6550 a_19479_31679# a_19721_31679# 9.039419f
C6551 a_16327_47482# a_22400_42852# 1.22e-21
C6552 a_n2017_45002# a_11691_44458# 4.56e-21
C6553 a_6171_45002# a_14309_45348# 3.25e-19
C6554 a_2107_46812# a_8349_46414# 0.003223f
C6555 a_n1151_42308# a_n755_45592# 0.03818f
C6556 a_6151_47436# a_n2661_45546# 1.33e-19
C6557 a_15009_46634# a_14513_46634# 0.001266f
C6558 a_3090_45724# a_14180_46812# 0.001631f
C6559 a_14084_46812# a_14226_46987# 0.005572f
C6560 a_14976_45028# a_14035_46660# 7.08e-22
C6561 a_n743_46660# a_11189_46129# 0.039903f
C6562 a_n971_45724# a_2277_45546# 1.64e-20
C6563 a_n237_47217# a_n443_42852# 5.8e-21
C6564 a_2063_45854# a_3316_45546# 0.00135f
C6565 a_2905_45572# a_1848_45724# 5.22e-19
C6566 a_19321_45002# a_18189_46348# 8.52e-20
C6567 a_5807_45002# a_19553_46090# 0.00287f
C6568 a_13747_46662# a_18819_46122# 0.039742f
C6569 a_13661_43548# a_18985_46122# 0.006378f
C6570 a_13675_47204# a_6945_45028# 6.96e-19
C6571 a_10227_46804# a_14371_46494# 1.79e-19
C6572 a_4883_46098# a_10044_46482# 5.79e-19
C6573 a_15368_46634# a_13885_46660# 5.26e-20
C6574 a_n881_46662# a_1337_46436# 4.92e-19
C6575 a_2959_46660# a_3483_46348# 5.18e-19
C6576 a_2864_46660# a_2698_46116# 4.69e-19
C6577 a_17538_32519# a_13258_32519# 0.054578f
C6578 a_14673_44172# VDD 0.381917f
C6579 a_4190_30871# a_18861_43218# 9.99e-19
C6580 a_16795_42852# a_17333_42852# 0.108694f
C6581 a_17595_43084# a_18083_42858# 0.046381f
C6582 a_n97_42460# a_17303_42282# 2.32e-20
C6583 a_3626_43646# a_14456_42282# 0.005342f
C6584 a_8975_43940# a_12607_44458# 0.004748f
C6585 w_11334_34010# a_18194_35068# 0.796644f
C6586 SMPL_ON_P a_n1386_35608# 0.012082f
C6587 a_n2956_39768# a_n4334_40480# 4.08e-19
C6588 a_20623_45572# a_11341_43940# 1.76e-21
C6589 a_n1177_44458# a_n356_44636# 1.98e-19
C6590 a_5205_44484# a_5244_44056# 1.29e-20
C6591 a_5111_44636# a_7542_44172# 0.039468f
C6592 a_n2956_37592# a_n2661_42282# 1.91e-20
C6593 a_1823_45246# a_4743_43172# 1.5e-19
C6594 a_n357_42282# a_12281_43396# 0.022975f
C6595 a_n443_42852# a_8423_43396# 0.007509f
C6596 a_n2017_45002# a_8333_44056# 1.11e-21
C6597 a_3232_43370# a_5663_43940# 0.090892f
C6598 a_n2661_44458# a_700_44734# 5e-19
C6599 a_14955_47212# a_413_45260# 2.11e-19
C6600 a_6151_47436# a_5205_44484# 0.010575f
C6601 a_4791_45118# a_8191_45002# 5e-20
C6602 a_13059_46348# a_13259_45724# 0.812126f
C6603 a_12465_44636# a_3357_43084# 1.30897f
C6604 SMPL_ON_N a_2437_43646# 2.94e-19
C6605 a_9290_44172# a_11133_46155# 0.051331f
C6606 a_6165_46155# a_2324_44458# 4.51e-19
C6607 a_n1076_46494# a_n967_46494# 0.007416f
C6608 a_n901_46420# a_n722_46482# 0.007399f
C6609 a_n1641_46494# a_n1533_46116# 0.057222f
C6610 a_6969_46634# a_2711_45572# 5.57e-20
C6611 a_10227_46804# a_n913_45002# 0.344574f
C6612 a_13507_46334# a_20447_31679# 8.21e-20
C6613 a_12549_44172# a_16147_45260# 9.2e-20
C6614 a_13747_46662# a_16223_45938# 0.02646f
C6615 a_8270_45546# a_n443_42852# 0.063811f
C6616 a_n1853_46287# a_n914_46116# 3.05e-19
C6617 a_18249_42858# a_7174_31319# 1.28e-20
C6618 a_n473_42460# a_n1630_35242# 0.049561f
C6619 a_19987_42826# a_19511_42282# 1.28e-19
C6620 a_196_42282# a_564_42282# 7.52e-19
C6621 a_n784_42308# a_n3674_37592# 0.254719f
C6622 a_n4318_38680# a_n3420_38528# 0.001905f
C6623 a_766_43646# VDD 0.009527f
C6624 a_n2017_45002# a_4190_30871# 0.025499f
C6625 a_9482_43914# a_10341_43396# 7.76e-20
C6626 a_14537_43396# a_14205_43396# 0.080783f
C6627 a_20205_31679# a_n1630_35242# 1.48e-19
C6628 a_4223_44672# a_5745_43940# 0.040431f
C6629 a_n2661_42834# a_3499_42826# 0.009315f
C6630 a_n2661_43922# a_2537_44260# 1.23e-19
C6631 a_1307_43914# a_9803_43646# 9.06e-20
C6632 a_18989_43940# a_15493_43940# 0.025737f
C6633 a_4955_46873# VDD 0.467566f
C6634 a_n2293_42834# a_648_43396# 6.38e-19
C6635 a_9313_44734# a_9672_43914# 1.48e-19
C6636 a_n2293_45010# a_743_42282# 1.96e-21
C6637 a_10903_43370# a_7174_31319# 4.88e-21
C6638 a_3422_30871# a_21145_44484# 6.39e-20
C6639 a_20193_45348# a_17538_32519# 2.12e-19
C6640 a_526_44458# a_5437_45600# 2.03e-20
C6641 a_2324_44458# a_10210_45822# 3.44e-20
C6642 a_5257_43370# a_n2293_42834# 5.57e-19
C6643 a_n881_46662# a_14539_43914# 1.15e-20
C6644 a_12741_44636# a_20273_45572# 0.028616f
C6645 a_17339_46660# a_n913_45002# 4.56e-21
C6646 a_20528_46660# a_3357_43084# 0.002704f
C6647 a_5807_45002# a_4223_44672# 4.42e-21
C6648 a_768_44030# a_10157_44484# 0.00283f
C6649 a_11189_46129# a_11136_45572# 0.042798f
C6650 a_20202_43084# a_21188_45572# 0.013137f
C6651 a_11415_45002# a_21363_45546# 0.011178f
C6652 a_18597_46090# a_9313_44734# 0.029282f
C6653 a_10809_44734# a_12427_45724# 0.01284f
C6654 a_5732_46660# a_n2661_43370# 6.03e-21
C6655 a_n2956_39768# a_n2661_44458# 1.99e-20
C6656 a_n1630_35242# a_n2946_37690# 1.09e-19
C6657 a_6123_31319# a_2113_38308# 7.39e-20
C6658 a_13258_32519# a_22465_38105# 0.056749f
C6659 a_22400_42852# a_22545_38993# 0.038805f
C6660 a_14097_32519# a_22521_39511# 7.51e-21
C6661 a_8292_43218# VDD 0.08228f
C6662 a_1606_42308# a_7754_38470# 1.54e-19
C6663 a_n2109_47186# SMPL_ON_P 0.049302f
C6664 a_n1920_47178# a_n1741_47186# 0.173125f
C6665 a_n2497_47436# a_n815_47178# 0.003116f
C6666 a_6945_45028# DATA[4] 0.0111f
C6667 a_2382_45260# a_1755_42282# 4.8e-19
C6668 a_n1059_45260# a_4921_42308# 6.43e-19
C6669 a_n913_45002# a_4933_42558# 0.005299f
C6670 a_n2017_45002# a_5337_42558# 0.001525f
C6671 a_n967_46494# VDD 2.82e-20
C6672 a_n2810_45572# a_n4064_37440# 1.13e-20
C6673 a_9313_44734# a_743_42282# 0.024013f
C6674 a_n23_44458# a_n1853_43023# 4.42e-21
C6675 a_8103_44636# a_8037_42858# 2.12e-21
C6676 a_20159_44458# a_10341_43396# 3.98e-20
C6677 a_2998_44172# a_2896_43646# 0.001865f
C6678 a_n2661_42282# a_n2267_43396# 5.11e-21
C6679 en_comp a_5379_42460# 1.81e-20
C6680 a_12549_44172# a_13565_44260# 4.96e-19
C6681 a_12891_46348# a_13829_44260# 1.39e-19
C6682 a_768_44030# a_12710_44260# 6.85e-19
C6683 a_13759_46122# a_11691_44458# 7.99e-21
C6684 a_n755_45592# a_327_44734# 0.00429f
C6685 a_8697_45822# a_8696_44636# 1.69e-20
C6686 a_12741_44636# a_18989_43940# 0.002238f
C6687 a_4646_46812# a_6453_43914# 8.23e-20
C6688 a_2711_45572# a_3357_43084# 0.037825f
C6689 a_3483_46348# a_n699_43396# 2.82e-19
C6690 a_n443_42852# a_n2017_45002# 0.033337f
C6691 a_n906_45572# a_n913_45002# 1.9e-19
C6692 a_13259_45724# a_13556_45296# 0.019616f
C6693 a_18819_46122# a_18911_45144# 4e-21
C6694 a_1823_45246# a_5883_43914# 3.03e-19
C6695 a_19321_45002# a_20935_43940# 9.4e-19
C6696 a_5807_45002# a_15493_43940# 1.03e-20
C6697 a_13747_46662# a_11341_43940# 0.008288f
C6698 a_18597_46090# a_20974_43370# 0.025672f
C6699 a_n443_46116# a_2982_43646# 0.140614f
C6700 a_n2661_45546# a_5111_44636# 0.001037f
C6701 a_n971_45724# a_6755_46942# 0.185154f
C6702 a_2063_45854# a_8145_46902# 0.003229f
C6703 a_n237_47217# a_10554_47026# 3.85e-20
C6704 a_7227_47204# a_4646_46812# 0.01221f
C6705 a_12465_44636# a_n2293_46634# 0.012816f
C6706 a_n4209_38216# C8_P_btm 1.65e-20
C6707 a_7754_38470# a_8912_37509# 0.575911f
C6708 a_3754_38470# a_11206_38545# 0.078412f
C6709 a_4915_47217# a_5732_46660# 4.19e-20
C6710 a_6545_47178# a_4817_46660# 1.23e-20
C6711 a_n1151_42308# a_5429_46660# 4.3e-19
C6712 a_4791_45118# a_5072_46660# 7.69e-21
C6713 a_n2302_39072# VDD 0.355374f
C6714 a_8530_39574# VDAC_N 0.06498f
C6715 a_10227_46804# a_2107_46812# 0.002063f
C6716 a_n4064_39616# VREF_GND 0.241027f
C6717 a_n4064_37440# a_n4251_37440# 0.00105f
C6718 a_n2302_37690# a_n2216_37690# 0.011479f
C6719 a_n3565_38216# C10_P_btm 2.25e-20
C6720 a_3499_42826# a_n2293_42282# 0.058548f
C6721 a_3905_42865# a_4149_42891# 0.002034f
C6722 a_20193_45348# a_22465_38105# 7.48e-20
C6723 a_19721_31679# a_13258_32519# 0.054727f
C6724 a_9396_43370# a_9803_43646# 9.33e-19
C6725 a_18909_45814# VDD 0.205795f
C6726 a_21381_43940# a_21487_43396# 0.007531f
C6727 a_15682_43940# a_15567_42826# 1.02e-19
C6728 a_5891_43370# a_7227_42308# 8.82e-19
C6729 a_n2293_43922# a_2713_42308# 4.97e-20
C6730 a_11341_43940# a_10796_42968# 4.28e-19
C6731 a_20974_43370# a_743_42282# 1.42e-19
C6732 a_14401_32519# a_20556_43646# 2.02e-19
C6733 a_19479_31679# a_18194_35068# 8.48e-20
C6734 en_comp a_22821_38993# 1.42e-19
C6735 a_4185_45028# a_22223_43948# 9.96e-19
C6736 a_16375_45002# a_11967_42832# 9.56e-20
C6737 a_n913_45002# a_1307_43914# 0.298747f
C6738 a_768_44030# a_685_42968# 5.63e-19
C6739 a_10490_45724# a_10057_43914# 4.22e-20
C6740 a_8746_45002# a_8975_43940# 0.016889f
C6741 a_16333_45814# a_11827_44484# 3.46e-21
C6742 a_n2661_45010# a_1423_45028# 4.66e-19
C6743 a_9290_44172# a_12429_44172# 0.040422f
C6744 a_3316_45546# a_n2661_42834# 6.51e-21
C6745 a_3218_45724# a_n2661_43922# 3.16e-20
C6746 a_n1613_43370# a_7765_42852# 0.081834f
C6747 a_n2017_45002# a_375_42282# 0.03181f
C6748 a_10903_43370# a_10729_43914# 0.082892f
C6749 a_n2293_45010# a_626_44172# 0.024201f
C6750 a_5691_45260# a_6171_45002# 0.057463f
C6751 a_5111_44636# a_5205_44484# 0.200189f
C6752 a_526_44458# a_2479_44172# 0.08343f
C6753 a_948_46660# a_765_45546# 7.87e-19
C6754 a_19321_45002# a_20202_43084# 2.61e-20
C6755 a_11459_47204# a_6945_45028# 0.010682f
C6756 a_11599_46634# a_18819_46122# 0.314824f
C6757 a_n971_45724# a_8049_45260# 0.078318f
C6758 a_n237_47217# a_6633_46155# 0.002406f
C6759 a_6755_46942# a_8023_46660# 0.004684f
C6760 a_10554_47026# a_8270_45546# 9.49e-20
C6761 a_16327_47482# a_15682_46116# 0.050548f
C6762 a_2063_45854# a_5066_45546# 0.055269f
C6763 a_5807_45002# a_12741_44636# 0.041091f
C6764 a_n881_46662# a_1823_45246# 0.155149f
C6765 a_4007_47204# a_526_44458# 6.28e-22
C6766 a_10227_46804# a_14493_46090# 0.202633f
C6767 a_4883_46098# a_9823_46155# 0.046689f
C6768 a_13887_32519# a_5342_30871# 0.028465f
C6769 a_14209_32519# a_5534_30871# 0.057361f
C6770 a_4190_30871# a_19164_43230# 0.005605f
C6771 a_14021_43940# a_15890_42674# 3.09e-21
C6772 a_11341_43940# a_4958_30871# 2.27e-20
C6773 a_12607_44458# VDD 0.188171f
C6774 a_4361_42308# a_17701_42308# 0.004927f
C6775 a_1568_43370# a_1184_42692# 2.36e-19
C6776 a_1756_43548# a_1576_42282# 1e-20
C6777 a_1049_43396# a_961_42354# 1.08e-19
C6778 a_n1557_42282# a_196_42282# 0.031105f
C6779 a_9145_43396# a_13291_42460# 6.23e-20
C6780 a_743_42282# a_18599_43230# 1.85e-20
C6781 a_n4318_39768# a_n4334_39392# 3.4e-19
C6782 a_n755_45592# a_n1809_43762# 1.04e-19
C6783 a_1423_45028# a_8855_44734# 1.81e-20
C6784 a_n2661_45546# a_4235_43370# 0.088313f
C6785 a_413_45260# a_11967_42832# 4.85e-22
C6786 a_n2293_46634# a_8515_42308# 1.72e-21
C6787 a_19479_31679# a_22591_44484# 0.00246f
C6788 a_21513_45002# a_19237_31679# 4.7e-20
C6789 a_12549_44172# a_15051_42282# 1.32e-20
C6790 a_n863_45724# a_1209_43370# 8.74e-19
C6791 a_13348_45260# a_13213_44734# 1.03e-19
C6792 a_9482_43914# a_n2293_43922# 0.018115f
C6793 a_1138_42852# a_421_43172# 3.71e-20
C6794 a_13507_46334# a_21887_42336# 0.002462f
C6795 a_n913_45002# a_18579_44172# 7.45e-21
C6796 a_16388_46812# a_17715_44484# 0.032772f
C6797 a_n2293_46098# a_2202_46116# 0.002053f
C6798 a_n237_47217# a_2437_43646# 0.076344f
C6799 a_12861_44030# a_13297_45572# 8.01e-20
C6800 a_10227_46804# a_15903_45785# 0.00138f
C6801 a_765_45546# a_13925_46122# 4.47e-20
C6802 a_n2497_47436# a_n2661_45010# 0.281004f
C6803 a_16327_47482# a_16680_45572# 0.223571f
C6804 a_8023_46660# a_8049_45260# 1.59e-19
C6805 a_768_44030# a_7499_43078# 0.101779f
C6806 a_n901_46420# a_472_46348# 2.86e-20
C6807 a_n1076_46494# a_376_46348# 4.41e-20
C6808 a_20820_30879# a_4185_45028# 2.33e-19
C6809 a_1799_45572# a_3218_45724# 2.5e-21
C6810 a_n2293_46634# a_2711_45572# 0.003426f
C6811 a_12347_46660# a_10809_44734# 0.001417f
C6812 a_4883_46098# a_10306_45572# 1.7e-19
C6813 a_21855_43396# a_21887_42336# 1.39e-19
C6814 a_n2293_42282# a_3318_42354# 0.01699f
C6815 a_22591_43396# a_13258_32519# 1.79e-20
C6816 a_13467_32519# a_22775_42308# 0.016923f
C6817 a_4361_42308# a_21613_42308# 0.001002f
C6818 a_5649_42852# a_7174_31319# 0.025928f
C6819 a_10796_42968# a_10723_42308# 0.003077f
C6820 a_10835_43094# a_11323_42473# 3.74e-19
C6821 a_10341_42308# a_9885_42558# 0.003164f
C6822 a_10518_42984# a_5742_30871# 0.001042f
C6823 a_1793_42852# a_1606_42308# 2.01e-20
C6824 a_21101_45002# a_19862_44208# 0.00117f
C6825 a_3065_45002# a_3626_43646# 0.480498f
C6826 a_11827_44484# a_15493_43396# 0.00117f
C6827 a_7499_43078# a_5755_42852# 2.12e-20
C6828 a_n1925_42282# a_n4318_38216# 1.9e-19
C6829 a_n863_45724# a_3059_42968# 0.003162f
C6830 a_3232_43370# a_4905_42826# 4.37e-21
C6831 a_4185_45028# a_11323_42473# 6.87e-20
C6832 a_18911_45144# a_11341_43940# 2.97e-20
C6833 a_n2956_38680# a_n1630_35242# 6.62e-19
C6834 a_n357_42282# a_873_42968# 5.83e-19
C6835 a_n755_45592# a_133_42852# 0.020885f
C6836 a_n881_46662# DATA[2] 2.22e-20
C6837 a_n913_45002# a_9396_43370# 9.91e-20
C6838 a_n1613_43370# DATA[3] 3.98e-19
C6839 a_11691_44458# a_18079_43940# 4.05e-20
C6840 a_3537_45260# a_2982_43646# 7.1e-19
C6841 a_16388_46812# a_15861_45028# 1.87e-21
C6842 a_16721_46634# a_8696_44636# 2.23e-19
C6843 a_6419_46155# a_6511_45714# 3.42e-19
C6844 a_4915_47217# a_16112_44458# 7.03e-21
C6845 a_5257_43370# a_413_45260# 1.46e-20
C6846 a_8270_45546# a_2437_43646# 5.82e-21
C6847 a_n2438_43548# a_2304_45348# 2.8e-21
C6848 a_9625_46129# a_2711_45572# 0.019316f
C6849 a_12891_46348# a_13490_45394# 5.25e-19
C6850 a_19466_46812# a_19431_45546# 0.038922f
C6851 a_2107_46812# a_1307_43914# 0.015866f
C6852 a_n2956_38680# a_n2661_45546# 0.003946f
C6853 a_4646_46812# a_6171_45002# 0.032849f
C6854 a_5167_46660# a_5147_45002# 4.02e-21
C6855 a_4817_46660# a_4927_45028# 1.88e-20
C6856 a_18597_46090# a_18114_32519# 4.06e-20
C6857 a_10227_46804# a_n2661_44458# 0.034728f
C6858 a_3681_42891# VDD 0.223661f
C6859 a_n4318_38216# a_n4334_38528# 5.87e-19
C6860 a_1606_42308# a_1736_39587# 1.72e-20
C6861 a_15803_42450# a_15959_42545# 0.110532f
C6862 a_15764_42576# a_15890_42674# 0.181217f
C6863 a_7963_42308# a_7174_31319# 4.88e-21
C6864 a_15486_42560# a_15720_42674# 0.006453f
C6865 COMP_P comp_n 0.033828f
C6866 a_n3674_38680# a_n3690_38528# 0.071909f
C6867 a_5342_30871# EN_VIN_BSTR_N 0.010795f
C6868 a_2998_44172# a_1443_43940# 7.55e-21
C6869 a_2675_43914# a_2455_43940# 0.007392f
C6870 a_2479_44172# a_3353_43940# 4.3e-20
C6871 a_20193_45348# a_22591_43396# 0.001393f
C6872 a_n2661_42834# a_6197_43396# 1.61e-19
C6873 a_376_46348# VDD 0.116284f
C6874 a_20820_30879# VREF_GND 0.02097f
C6875 a_3537_45260# a_5837_42852# 0.042825f
C6876 a_11823_42460# a_13249_42558# 0.004086f
C6877 a_10193_42453# a_15959_42545# 1.6e-19
C6878 a_2711_45572# a_20107_42308# 0.164316f
C6879 a_n1059_45260# a_13291_42460# 0.03043f
C6880 a_n2017_45002# a_14635_42282# 0.025779f
C6881 a_n913_45002# a_13003_42852# 0.026478f
C6882 a_n356_44636# a_14205_43396# 6.46e-21
C6883 a_7499_43078# a_10149_42308# 3.73e-19
C6884 a_11415_45002# a_19778_44110# 0.030651f
C6885 a_20202_43084# a_18184_42460# 0.299795f
C6886 a_n443_46116# a_2253_43940# 0.011444f
C6887 a_15682_46116# a_14537_43396# 2.16e-21
C6888 a_2324_44458# a_14797_45144# 0.048583f
C6889 a_2711_45572# a_9159_45572# 0.003753f
C6890 a_6945_45028# a_8191_45002# 8.52e-21
C6891 a_10193_42453# a_8746_45002# 0.11003f
C6892 a_526_44458# a_2680_45002# 0.119733f
C6893 a_n1925_42282# a_2382_45260# 4.45e-19
C6894 a_10180_45724# a_10490_45724# 7.31e-21
C6895 a_15227_44166# a_15004_44636# 7.56e-19
C6896 a_3090_45724# a_18287_44626# 0.037072f
C6897 a_768_44030# a_3600_43914# 0.182408f
C6898 a_n1613_43370# a_n1644_44306# 0.001113f
C6899 a_n2312_39304# a_n2661_42282# 6.22e-20
C6900 a_7499_43078# a_11652_45724# 1.11e-20
C6901 a_6755_46942# a_9313_44734# 3.88e-20
C6902 a_1138_42852# a_n2661_43370# 0.023497f
C6903 a_12741_44636# a_18315_45260# 0.011294f
C6904 a_7227_45028# a_8697_45822# 3.36e-20
C6905 a_5164_46348# a_5093_45028# 0.003673f
C6906 a_16327_47482# a_20269_44172# 8.13e-19
C6907 a_15959_42545# VDD 0.19373f
C6908 a_15803_42450# RST_Z 1.82e-19
C6909 SMPL_ON_P a_n1925_46634# 1.71e-19
C6910 a_22465_38105# a_22609_37990# 3.5e-19
C6911 a_n237_47217# a_n2661_46634# 0.067716f
C6912 a_6151_47436# a_12891_46348# 0.169139f
C6913 a_18597_46090# a_12465_44636# 3.19e-19
C6914 a_19787_47423# a_4883_46098# 8.92e-21
C6915 a_7903_47542# a_8128_46384# 0.109077f
C6916 a_11031_47542# a_n881_46662# 0.183988f
C6917 a_10227_46804# a_11453_44696# 0.08211f
C6918 a_20990_47178# a_13507_46334# 0.017412f
C6919 a_n2109_47186# a_n2438_43548# 5.34e-19
C6920 a_4958_30871# C1_P_btm 9.46e-20
C6921 a_17737_43940# a_743_42282# 9.59e-21
C6922 a_9313_44734# a_16328_43172# 1.1e-19
C6923 a_n2810_45028# a_n4209_38216# 0.063751f
C6924 a_15493_43940# a_16867_43762# 6.77e-19
C6925 a_3905_42865# a_5111_42852# 0.079376f
C6926 a_742_44458# a_2713_42308# 7.64e-19
C6927 a_8746_45002# VDD 0.970181f
C6928 a_n97_42460# a_6031_43396# 0.002248f
C6929 a_1756_43548# a_1987_43646# 0.004999f
C6930 a_3422_30871# a_17333_42852# 1.02e-20
C6931 a_11750_44172# a_4361_42308# 1.32e-21
C6932 a_18079_43940# a_4190_30871# 4.22e-21
C6933 a_10193_42453# RST_Z 4.5e-19
C6934 a_14021_43940# a_16547_43609# 0.005885f
C6935 a_17339_46660# a_18451_43940# 0.012866f
C6936 a_2063_45854# a_10922_42852# 1.31e-20
C6937 a_13747_46662# a_10341_43396# 4.28e-20
C6938 a_18985_46122# a_11967_42832# 1.38e-21
C6939 a_8696_44636# a_14180_45002# 5.97e-21
C6940 a_2711_45572# a_16237_45028# 0.001569f
C6941 a_16680_45572# a_14537_43396# 3.12e-20
C6942 a_15765_45572# a_16019_45002# 0.001223f
C6943 a_15599_45572# a_16751_45260# 0.012353f
C6944 a_15903_45785# a_1307_43914# 8.62e-19
C6945 a_13507_46334# a_13467_32519# 0.043891f
C6946 a_2107_46812# a_9396_43370# 0.001284f
C6947 a_1823_45246# a_2889_44172# 3.93e-19
C6948 a_1848_45724# a_949_44458# 4.69e-19
C6949 a_n357_42282# a_n699_43396# 0.055761f
C6950 a_n755_45592# a_4223_44672# 3.55e-19
C6951 a_5066_45546# a_n2661_42834# 1.32e-20
C6952 a_18051_46116# a_18248_44752# 4.95e-21
C6953 a_11652_45724# a_11915_45394# 6.1e-19
C6954 a_8049_45260# a_9313_44734# 5.74e-21
C6955 a_n2293_46634# a_7466_43396# 2.46e-19
C6956 a_13507_46334# a_20273_46660# 0.026778f
C6957 a_21177_47436# a_20841_46902# 0.001161f
C6958 a_20990_47178# a_20623_46660# 0.004006f
C6959 C0_P_btm VREF_GND 0.350485f
C6960 C1_P_btm VCM 0.716121f
C6961 VDD RST_Z 4.72146f
C6962 a_2063_45854# a_5068_46348# 0.004281f
C6963 a_n237_47217# a_8199_44636# 0.089777f
C6964 a_n971_45724# a_8953_45546# 5.83e-21
C6965 a_11453_44696# a_17339_46660# 0.071641f
C6966 a_12465_44636# a_19123_46287# 1.94e-20
C6967 a_18597_46090# a_20528_46660# 8.24e-19
C6968 a_3877_44458# a_4817_46660# 0.017126f
C6969 a_4646_46812# a_4955_46873# 0.047208f
C6970 a_n1925_46634# a_8035_47026# 2.38e-20
C6971 a_n1151_42308# a_3483_46348# 8.25e-19
C6972 a_3160_47472# a_3699_46348# 0.109505f
C6973 a_2905_45572# a_4185_45028# 1.92e-21
C6974 a_768_44030# a_15227_44166# 3.48e-22
C6975 a_12549_44172# a_19333_46634# 3.59e-19
C6976 C0_dummy_N_btm VIN_N 0.544204f
C6977 a_n443_46116# a_1823_45246# 0.217935f
C6978 a_13747_46662# a_12991_46634# 1.32e-20
C6979 a_5807_45002# a_13607_46688# 0.002972f
C6980 a_n2661_46634# a_8270_45546# 0.037557f
C6981 a_n1741_47186# a_9290_44172# 9.99e-21
C6982 a_16327_47482# a_20719_46660# 5.41e-20
C6983 a_4883_46098# a_20107_46660# 1.93e-19
C6984 a_13467_32519# a_21855_43396# 0.003525f
C6985 a_21487_43396# a_5649_42852# 8.4e-20
C6986 a_4190_30871# a_14209_32519# 0.031783f
C6987 a_19721_31679# a_22609_37990# 7.56e-21
C6988 a_9145_43396# a_13460_43230# 0.002473f
C6989 a_20512_43084# a_20712_42282# 2.86e-20
C6990 a_10341_43396# a_10796_42968# 9.03e-20
C6991 a_1307_43914# a_n2661_44458# 0.007888f
C6992 a_8191_45002# a_8103_44636# 2.19e-19
C6993 a_3090_45724# a_9127_43156# 8.78e-19
C6994 a_8016_46348# a_9803_43646# 7.46e-19
C6995 a_3232_43370# a_8975_43940# 0.620589f
C6996 a_6171_45002# a_10057_43914# 1.53e-19
C6997 a_n967_45348# a_n356_44636# 2.16e-20
C6998 a_7499_43078# a_7845_44172# 0.112307f
C6999 a_4646_46812# a_8292_43218# 2.63e-20
C7000 a_2107_46812# a_8034_45724# 0.006608f
C7001 a_2864_46660# a_526_44458# 8.51e-20
C7002 a_8492_46660# a_2324_44458# 1.06e-20
C7003 a_n881_46662# a_n2293_45546# 0.004473f
C7004 a_20273_46660# a_20623_46660# 0.20669f
C7005 a_20107_46660# a_21188_46660# 0.102355f
C7006 a_19123_46287# a_20528_46660# 1.39e-20
C7007 a_n1613_43370# a_n1079_45724# 0.013012f
C7008 a_18597_46090# a_2711_45572# 2.61e-20
C7009 a_n743_46660# a_8379_46155# 1.92e-19
C7010 a_6755_46942# a_12594_46348# 1.41e-19
C7011 a_5807_45002# a_16375_45002# 0.042941f
C7012 a_8270_45546# a_8199_44636# 0.95539f
C7013 a_17339_46660# a_17639_46660# 0.081726f
C7014 a_n971_45724# a_8791_45572# 1.43e-20
C7015 a_5663_43940# VDD 0.133666f
C7016 a_3681_42891# a_n784_42308# 1.66e-21
C7017 a_15567_42826# a_16245_42852# 0.03084f
C7018 a_16547_43609# a_15764_42576# 2.95e-21
C7019 a_16243_43396# a_15803_42450# 2.1e-20
C7020 a_16137_43396# a_15959_42545# 0.001471f
C7021 a_5649_42852# a_5932_42308# 0.126438f
C7022 a_4361_42308# a_6761_42308# 0.042179f
C7023 a_743_42282# a_8515_42308# 0.005514f
C7024 a_10341_43396# a_4958_30871# 4.26e-20
C7025 a_18083_42858# a_18695_43230# 0.001881f
C7026 a_17333_42852# a_18504_43218# 0.157683f
C7027 a_n443_46116# DATA[2] 0.006001f
C7028 a_10193_42453# a_16243_43396# 2.07e-19
C7029 a_2711_45572# a_743_42282# 0.039036f
C7030 a_6171_45002# a_14021_43940# 5.61e-20
C7031 a_5891_43370# a_8238_44734# 9.85e-19
C7032 a_n1821_44484# a_n2661_42834# 0.001026f
C7033 a_22959_45036# a_19237_31679# 0.005799f
C7034 a_n863_45724# a_n722_43218# 6.21e-21
C7035 SMPL_ON_N a_22609_38406# 9.53e-21
C7036 a_2382_45260# a_3737_43940# 0.027805f
C7037 a_12883_44458# a_13296_44484# 5.31e-19
C7038 a_12607_44458# a_13940_44484# 5.31e-19
C7039 a_8375_44464# a_8333_44734# 7.47e-21
C7040 a_6851_47204# VDD 0.287724f
C7041 a_4791_45118# DATA[3] 5.9e-20
C7042 a_n2661_43370# a_n4318_39768# 0.068386f
C7043 a_13249_42308# a_12281_43396# 1.91e-19
C7044 a_13348_45260# a_11341_43940# 1.4e-21
C7045 w_11334_34010# a_18114_32519# 9.7e-19
C7046 a_8270_45546# a_8192_45572# 0.048422f
C7047 a_768_44030# a_4558_45348# 5.74e-21
C7048 a_11453_44696# a_1307_43914# 0.037741f
C7049 a_4883_46098# a_1423_45028# 0.022493f
C7050 a_9290_44172# a_10586_45546# 0.264957f
C7051 a_9625_46129# a_10037_46155# 0.006879f
C7052 a_n2293_46098# a_n1079_45724# 0.003233f
C7053 a_n2157_46122# a_n2293_45546# 6.79e-20
C7054 a_6755_46942# a_15037_45618# 1.85e-20
C7055 a_5807_45002# a_413_45260# 1.49e-19
C7056 a_9804_47204# a_6171_45002# 7.74e-21
C7057 a_n2293_46634# a_n2472_45002# 0.001349f
C7058 a_n881_46662# a_6709_45028# 0.011804f
C7059 a_12594_46348# a_8049_45260# 0.069217f
C7060 a_n2956_38680# a_n1533_46116# 9.67e-20
C7061 a_16243_43396# VDD 0.39865f
C7062 a_6171_42473# a_5934_30871# 1.01e-20
C7063 a_16137_43396# RST_Z 1.66e-20
C7064 a_1606_42308# a_13070_42354# 1.69e-20
C7065 a_3232_43370# a_2905_42968# 0.008509f
C7066 a_3537_45260# a_7871_42858# 8.33e-19
C7067 a_n913_45002# a_13635_43156# 0.036742f
C7068 a_n1059_45260# a_13460_43230# 0.004971f
C7069 a_18911_45144# a_10341_43396# 2.05e-21
C7070 a_13259_45724# a_17303_42282# 0.460497f
C7071 a_20640_44752# a_20623_43914# 0.003088f
C7072 a_20820_30879# a_22469_40625# 2.62e-20
C7073 a_3090_45724# CLK 0.001129f
C7074 a_n755_45592# a_5742_30871# 5.83e-20
C7075 a_n357_42282# a_11551_42558# 1.33e-19
C7076 a_19615_44636# a_11341_43940# 2.34e-21
C7077 a_14673_44172# a_14021_43940# 4.52e-19
C7078 a_n2661_42834# a_8415_44056# 1.54e-35
C7079 a_20766_44850# a_19862_44208# 1.08e-19
C7080 a_n699_43396# a_n144_43396# 1.99e-19
C7081 a_19692_46634# START 1.28e-19
C7082 a_18579_44172# a_18451_43940# 0.147572f
C7083 a_n2661_44458# a_9396_43370# 1.17e-21
C7084 a_5495_43940# a_5663_43940# 0.227135f
C7085 a_19279_43940# a_19478_44306# 0.03583f
C7086 a_5111_44636# a_4520_42826# 1.98e-19
C7087 a_5147_45002# a_5111_42852# 1.57e-20
C7088 a_13507_46334# a_22315_44484# 1.46e-19
C7089 a_13759_46122# a_2437_43646# 5.19e-20
C7090 a_3090_45724# a_17023_45118# 1.26e-20
C7091 a_8199_44636# a_n2017_45002# 0.020035f
C7092 a_8016_46348# a_n913_45002# 1.22e-20
C7093 a_1848_45724# a_1990_45572# 0.007833f
C7094 a_10586_45546# a_11064_45572# 6.98e-19
C7095 a_12741_44636# a_13017_45260# 9.29e-21
C7096 a_12005_46116# a_3357_43084# 8.11e-21
C7097 a_584_46384# a_3499_42826# 0.036739f
C7098 a_2698_46116# a_2382_45260# 4.99e-21
C7099 a_1823_45246# a_3537_45260# 0.482502f
C7100 a_12549_44172# a_12553_44484# 4.66e-19
C7101 a_11415_45002# a_9482_43914# 0.309633f
C7102 a_8049_45260# a_15037_45618# 0.001405f
C7103 a_2277_45546# a_2711_45572# 0.01233f
C7104 a_n784_42308# RST_Z 0.033698f
C7105 a_1606_42308# C2_N_btm 0.021793f
C7106 a_n327_42558# VDD 0.198414f
C7107 a_n4064_40160# a_n4334_38304# 0.013157f
C7108 a_n2946_39072# a_n2302_39072# 6.68e-19
C7109 a_n3690_39392# a_n3607_39392# 0.007692f
C7110 a_6545_47178# a_7227_47204# 0.001559f
C7111 a_5815_47464# a_6575_47204# 0.009009f
C7112 a_n1151_42308# a_13487_47204# 1.36e-19
C7113 a_4915_47217# a_9863_47436# 0.018512f
C7114 a_6151_47436# a_7903_47542# 7.86e-20
C7115 a_6491_46660# a_6851_47204# 0.132946f
C7116 a_3815_47204# a_n1435_47204# 2.24e-19
C7117 a_1443_43940# a_1568_43370# 4.63e-19
C7118 a_n2017_45002# a_19511_42282# 6.66e-20
C7119 a_n1059_45260# a_18548_42308# 0.001247f
C7120 a_21167_46155# VDD 8.63e-19
C7121 a_3422_30871# a_13678_32519# 0.452533f
C7122 a_n2293_43922# a_10796_42968# 2.47e-20
C7123 a_10729_43914# a_8685_43396# 5.97e-22
C7124 en_comp a_18907_42674# 1.94e-20
C7125 a_18184_42460# a_19326_42852# 1.25e-20
C7126 a_9313_44734# a_15279_43071# 0.007423f
C7127 a_20512_43084# a_20556_43646# 9.96e-19
C7128 a_5907_45546# a_1307_43914# 2.22e-20
C7129 a_18985_46122# a_18989_43940# 5.94e-20
C7130 a_8049_45260# a_18114_32519# 5.83e-20
C7131 a_11415_45002# a_20159_44458# 5.37e-19
C7132 a_12741_44636# a_19006_44850# 0.001054f
C7133 a_18175_45572# a_18691_45572# 0.105995f
C7134 a_18479_45785# a_18909_45814# 0.023226f
C7135 a_n1925_42282# a_5343_44458# 5.11e-21
C7136 a_8034_45724# a_n2661_44458# 7.74e-21
C7137 a_768_44030# a_1756_43548# 0.093469f
C7138 a_16375_45002# a_18315_45260# 4.03e-21
C7139 a_10193_42453# a_3232_43370# 0.016241f
C7140 a_10180_45724# a_6171_45002# 0.03378f
C7141 a_6755_46942# a_17737_43940# 5.46e-19
C7142 a_n1613_43370# a_2982_43646# 8.34e-20
C7143 w_11334_34010# a_13887_32519# 3.17e-19
C7144 a_10227_46804# a_9145_43396# 0.066362f
C7145 a_8953_45546# a_9313_44734# 3.9e-19
C7146 a_13259_45724# a_19778_44110# 1.81e-20
C7147 a_3483_46348# a_13857_44734# 0.005876f
C7148 a_n2956_38216# a_n2661_43370# 0.028301f
C7149 a_n755_45592# a_n2293_42834# 0.059468f
C7150 a_10227_46804# a_10384_47026# 1.7e-19
C7151 a_n237_47217# a_765_45546# 0.1364f
C7152 a_13717_47436# a_3090_45724# 2.02e-20
C7153 a_12861_44030# a_15009_46634# 0.058082f
C7154 a_13487_47204# a_14084_46812# 0.012167f
C7155 a_n1613_43370# a_6540_46812# 0.05541f
C7156 a_n1386_35608# a_n923_35174# 0.201937f
C7157 a_n1838_35608# EN_VIN_BSTR_P 2.62e-19
C7158 VDAC_N C3_N_btm 1.98783f
C7159 a_11599_46634# a_12991_46634# 4.06e-20
C7160 a_n2661_46634# a_1123_46634# 0.012266f
C7161 a_n2293_46634# a_33_46660# 6.74e-21
C7162 CAL_P a_21589_35634# 0.00593f
C7163 a_12465_44636# a_6755_46942# 0.021176f
C7164 a_n2860_37690# VDD 0.004184f
C7165 a_2063_45854# a_13059_46348# 5.17e-21
C7166 a_4915_47217# a_12978_47026# 1.2e-19
C7167 a_n1151_42308# a_14513_46634# 0.042579f
C7168 a_n1925_46634# a_n2438_43548# 0.166008f
C7169 a_n1021_46688# a_n743_46660# 0.11001f
C7170 a_4235_43370# a_4520_42826# 0.001794f
C7171 a_3080_42308# a_3681_42891# 5.97e-19
C7172 a_n97_42460# a_10796_42968# 3.04e-19
C7173 a_n3674_39768# a_n4318_37592# 0.023075f
C7174 a_10341_43396# a_15125_43396# 7.22e-20
C7175 a_3232_43370# VDD 2.96597f
C7176 a_16137_43396# a_16243_43396# 0.182209f
C7177 a_9313_44734# a_13258_32519# 0.003166f
C7178 a_3422_30871# a_6123_31319# 0.021957f
C7179 a_14401_32519# a_5342_30871# 0.062032f
C7180 a_584_46384# a_3318_42354# 1.04e-20
C7181 a_1138_42852# a_1568_43370# 9.74e-20
C7182 a_n1099_45572# a_453_43940# 2.55e-20
C7183 a_n357_42282# a_1467_44172# 0.002404f
C7184 a_n755_45592# a_1115_44172# 2.69e-21
C7185 a_15227_44166# a_16759_43396# 8.01e-19
C7186 a_10775_45002# a_10903_45394# 0.004764f
C7187 a_7229_43940# a_n2661_43370# 0.040132f
C7188 a_n863_45724# a_895_43940# 0.015488f
C7189 a_10586_45546# a_10807_43548# 1.23e-21
C7190 a_n2661_45546# a_3905_42865# 0.001705f
C7191 a_19479_31679# a_18114_32519# 0.182316f
C7192 a_16327_47482# a_20836_43172# 0.001598f
C7193 a_3090_45724# a_19268_43646# 0.003095f
C7194 a_22223_45572# a_19721_31679# 8.73e-19
C7195 a_6171_45002# a_13711_45394# 9.69e-20
C7196 a_n443_46116# a_1184_42692# 3.57e-21
C7197 a_2107_46812# a_8016_46348# 0.022583f
C7198 a_3160_47472# a_n755_45592# 0.001373f
C7199 a_n1151_42308# a_n357_42282# 0.009369f
C7200 a_15009_46634# a_14180_46812# 0.123843f
C7201 a_14976_45028# a_13885_46660# 6.33e-20
C7202 a_3090_45724# a_14035_46660# 6.08e-22
C7203 a_n743_46660# a_9290_44172# 0.048675f
C7204 a_n746_45260# a_n443_42852# 0.136813f
C7205 a_2063_45854# a_3218_45724# 0.004182f
C7206 a_584_46384# a_3316_45546# 1.77e-21
C7207 a_n971_45724# a_1609_45822# 1.47e-19
C7208 a_n443_46116# a_n2293_45546# 0.004986f
C7209 a_8270_45546# a_765_45546# 5.94e-19
C7210 a_4883_46098# a_9823_46482# 2.91e-19
C7211 a_10227_46804# a_14180_46482# 0.014179f
C7212 a_12465_44636# a_8049_45260# 0.027831f
C7213 a_n881_46662# a_n914_46116# 1.02e-19
C7214 a_2959_46660# a_3147_46376# 0.010696f
C7215 a_3177_46902# a_3483_46348# 2.05e-20
C7216 a_13569_47204# a_6945_45028# 6.5e-19
C7217 a_13661_43548# a_18819_46122# 0.02447f
C7218 a_13747_46662# a_17957_46116# 1.02e-19
C7219 a_5807_45002# a_18985_46122# 0.017912f
C7220 a_20974_43370# a_13258_32519# 7.54e-21
C7221 a_8791_43396# a_8685_42308# 1.69e-21
C7222 a_17595_43084# a_17701_42308# 0.141211f
C7223 a_16795_42852# a_18083_42858# 6.33e-21
C7224 a_16414_43172# a_17333_42852# 2.98e-20
C7225 a_5111_42852# a_5457_43172# 0.013377f
C7226 a_3626_43646# a_13575_42558# 0.008305f
C7227 a_n97_42460# a_4958_30871# 0.069553f
C7228 a_3422_30871# EN_VIN_BSTR_P 0.182769f
C7229 a_n2129_44697# a_7_44811# 1.23e-19
C7230 w_11334_34010# EN_VIN_BSTR_N 3.99277f
C7231 SMPL_ON_P a_n1838_35608# 0.399535f
C7232 a_n2956_39768# a_n4315_30879# 0.056491f
C7233 a_20528_45572# a_20365_43914# 4.03e-21
C7234 a_n1917_44484# a_n356_44636# 1.7e-20
C7235 a_20193_45348# a_9313_44734# 0.056112f
C7236 a_1823_45246# a_4649_43172# 3.11e-19
C7237 a_n2810_45028# a_n2661_42282# 2.09e-20
C7238 a_3232_43370# a_5495_43940# 0.060353f
C7239 a_5691_45260# a_5663_43940# 4.64e-21
C7240 a_n2433_44484# a_n1243_44484# 2.56e-19
C7241 a_15037_45618# a_15037_43940# 1.4e-21
C7242 a_n443_42852# a_8317_43396# 0.00203f
C7243 a_16327_47482# en_comp 3.13e-20
C7244 a_4791_45118# a_7705_45326# 9.46e-20
C7245 a_13059_46348# a_14383_46116# 3.09e-20
C7246 a_22731_47423# a_2437_43646# 3.67e-19
C7247 a_14311_47204# a_413_45260# 8.86e-20
C7248 a_10355_46116# a_11133_46155# 6.26e-20
C7249 a_n1423_46090# a_n1533_46116# 0.097745f
C7250 a_9290_44172# a_11189_46129# 0.199578f
C7251 a_6755_46942# a_2711_45572# 0.612305f
C7252 a_21811_47423# a_3357_43084# 9.16e-21
C7253 a_10227_46804# a_n1059_45260# 0.036978f
C7254 a_6545_47178# a_6171_45002# 3.78e-20
C7255 a_6151_47436# a_6431_45366# 8.2e-20
C7256 a_13661_43548# a_16223_45938# 3.77e-20
C7257 a_13747_46662# a_16020_45572# 0.016423f
C7258 a_n746_45260# a_375_42282# 0.41439f
C7259 a_3080_42308# RST_Z 0.00595f
C7260 a_17333_42852# a_7174_31319# 7.1e-21
C7261 a_n961_42308# a_n1630_35242# 0.028868f
C7262 a_10793_43218# a_5742_30871# 4.83e-21
C7263 a_19339_43156# a_19647_42308# 0.009735f
C7264 a_19164_43230# a_19511_42282# 0.001746f
C7265 a_196_42282# a_n3674_37592# 0.1528f
C7266 a_n4318_38680# a_n3690_38528# 1.96e-19
C7267 a_n784_42308# a_n327_42558# 5.3e-19
C7268 a_4905_42826# VDD 0.439034f
C7269 a_19479_31679# a_13887_32519# 0.051118f
C7270 a_9482_43914# a_9885_43646# 7.99e-20
C7271 a_1423_45028# a_8685_43396# 1.34e-21
C7272 a_14537_43396# a_14358_43442# 0.1418f
C7273 a_n2956_38216# COMP_P 1.9e-21
C7274 a_4223_44672# a_5326_44056# 4.3e-19
C7275 a_4651_46660# VDD 0.457722f
C7276 a_n2661_43922# a_2253_44260# 3.34e-19
C7277 a_n2661_42834# a_2537_44260# 1.37e-19
C7278 a_13556_45296# a_14955_43396# 8.22e-21
C7279 a_1307_43914# a_9145_43396# 0.003867f
C7280 a_18374_44850# a_15493_43940# 4.07e-21
C7281 a_n2293_42834# a_548_43396# 2.62e-19
C7282 a_19963_31679# a_13678_32519# 0.051335f
C7283 a_3422_30871# a_21073_44484# 3.97e-20
C7284 a_21398_44850# a_21145_44484# 4.61e-19
C7285 a_20193_45348# a_20974_43370# 0.026944f
C7286 a_12741_44636# a_20107_45572# 0.029025f
C7287 a_17339_46660# a_n1059_45260# 2.95e-19
C7288 a_768_44030# a_9838_44484# 0.00219f
C7289 a_9290_44172# a_11136_45572# 0.008811f
C7290 a_11189_46129# a_11064_45572# 7.76e-20
C7291 a_20202_43084# a_21363_45546# 0.029873f
C7292 a_11415_45002# a_20623_45572# 0.006621f
C7293 a_12991_46634# a_13348_45260# 7.26e-22
C7294 a_12816_46660# a_13159_45002# 3.88e-19
C7295 a_n2956_39768# a_n4318_40392# 0.023582f
C7296 a_10809_44734# a_11962_45724# 0.033571f
C7297 a_8049_45260# a_2711_45572# 2.31131f
C7298 a_6945_45028# a_11823_42460# 9.85e-22
C7299 a_n1630_35242# a_n3420_37440# 6.45e-19
C7300 a_n2288_47178# SMPL_ON_P 0.002143f
C7301 a_n2109_47186# a_n1741_47186# 0.18579f
C7302 a_n2497_47436# a_n1605_47204# 0.0417f
C7303 a_n3674_37592# a_n4064_37440# 0.651412f
C7304 a_19511_42282# a_21973_42336# 1.79e-19
C7305 a_22400_42852# a_22521_39511# 0.031206f
C7306 a_21887_42336# a_21613_42308# 0.071168f
C7307 a_5742_30871# a_n3420_38528# 0.004679f
C7308 a_2382_45260# a_1606_42308# 1.35e-20
C7309 a_n2017_45002# a_4921_42308# 0.006208f
C7310 a_n913_45002# a_3905_42558# 0.047606f
C7311 a_n1379_46482# VDD 1.08e-19
C7312 a_6945_45028# DATA[3] 0.014238f
C7313 a_5891_43370# a_4361_42308# 0.028094f
C7314 a_8103_44636# a_7765_42852# 4.51e-20
C7315 a_11827_44484# a_21356_42826# 5.05e-21
C7316 a_n2956_38216# a_n3565_37414# 0.001835f
C7317 a_2889_44172# a_2896_43646# 0.001151f
C7318 a_2479_44172# a_3626_43646# 3.71e-20
C7319 a_644_44056# a_648_43396# 2.15e-19
C7320 a_n2956_39304# CLK_DATA 0.003272f
C7321 a_5495_43940# a_4905_42826# 0.001789f
C7322 a_19615_44636# a_10341_43396# 2.09e-21
C7323 a_19321_45002# a_20623_43914# 0.294126f
C7324 a_13661_43548# a_11341_43940# 0.15891f
C7325 a_13747_46662# a_21115_43940# 0.02491f
C7326 a_12891_46348# a_13565_44260# 9.26e-19
C7327 a_12549_44172# a_12710_44260# 7.8e-19
C7328 a_768_44030# a_12603_44260# 0.00112f
C7329 a_19900_46494# a_16922_45042# 3.54e-21
C7330 a_n755_45592# a_413_45260# 0.032345f
C7331 a_n357_42282# a_327_44734# 0.078335f
C7332 a_n863_45724# a_3065_45002# 2.64e-21
C7333 a_12741_44636# a_18374_44850# 0.002579f
C7334 a_4646_46812# a_5663_43940# 2.23e-19
C7335 a_15227_44166# a_17517_44484# 0.104904f
C7336 a_13059_46348# a_n2661_42834# 2.13e-21
C7337 a_5066_45546# a_5093_45028# 5.33e-19
C7338 a_14275_46494# a_11827_44484# 2.75e-21
C7339 a_8016_46348# a_n2661_44458# 0.030129f
C7340 a_3483_46348# a_4223_44672# 4.16e-19
C7341 a_310_45028# a_1667_45002# 6.44e-21
C7342 a_11064_45572# a_11136_45572# 0.003395f
C7343 a_13163_45724# a_13485_45572# 0.001367f
C7344 a_n2293_45546# a_3537_45260# 8.32e-21
C7345 a_18597_46090# a_14401_32519# 3e-20
C7346 a_10193_42453# a_18341_45572# 6.23e-22
C7347 a_4791_45118# a_2982_43646# 0.002472f
C7348 a_n443_46116# a_2896_43646# 0.039985f
C7349 a_11823_42460# a_14127_45572# 3.38e-19
C7350 a_n2661_45546# a_5147_45002# 6.41e-20
C7351 a_18189_46348# a_19778_44110# 1.37e-20
C7352 a_13259_45724# a_9482_43914# 0.321549f
C7353 a_2063_45854# a_7577_46660# 0.032724f
C7354 a_n237_47217# a_10623_46897# 1.75e-20
C7355 a_6491_46660# a_4651_46660# 1.14e-20
C7356 a_n1435_47204# a_3524_46660# 7.47e-21
C7357 a_6851_47204# a_4646_46812# 8.39e-20
C7358 a_n4209_38216# C9_P_btm 1.91e-20
C7359 a_n4064_38528# C1_P_btm 4.13e-20
C7360 a_3754_38470# VDAC_P 0.323951f
C7361 a_4791_45118# a_6540_46812# 0.001459f
C7362 a_4915_47217# a_5907_46634# 1.88e-19
C7363 a_5129_47502# a_5167_46660# 6.56e-19
C7364 a_6151_47436# a_4817_46660# 1.46e-20
C7365 a_n1151_42308# a_5263_46660# 0.001012f
C7366 a_n881_46662# a_15928_47570# 2.48e-20
C7367 a_n4064_39072# VDD 1.74897f
C7368 a_7754_38470# VDAC_N 0.110573f
C7369 a_8530_39574# a_6886_37412# 0.616015f
C7370 a_n4064_39616# VREF 1.53e-20
C7371 a_n3420_39616# VCM 0.0424f
C7372 a_22959_47212# a_22612_30879# 0.156518f
C7373 a_n4064_37440# a_n2216_37690# 0.005567f
C7374 a_n3420_37440# a_n3607_37440# 0.001516f
C7375 a_3905_42865# a_3863_42891# 1.54e-19
C7376 a_18114_32519# a_13258_32519# 0.059438f
C7377 a_20193_45348# a_22397_42558# 0.00176f
C7378 a_9396_43370# a_9145_43396# 0.030617f
C7379 a_18341_45572# VDD 0.2432f
C7380 a_5891_43370# a_6761_42308# 0.010358f
C7381 a_11341_43940# a_10835_43094# 1.05e-19
C7382 a_19479_31679# EN_VIN_BSTR_N 0.007584f
C7383 a_20974_43370# a_20301_43646# 9.11e-21
C7384 a_17538_32519# a_4190_30871# 1.16e-20
C7385 en_comp a_22545_38993# 7.26e-21
C7386 a_n1613_43370# a_7871_42858# 0.659491f
C7387 a_3483_46348# a_15493_43940# 0.026486f
C7388 a_4185_45028# a_11341_43940# 1.23e-19
C7389 a_3537_45260# a_6709_45028# 5.94e-20
C7390 a_n1059_45260# a_1307_43914# 0.016622f
C7391 a_10193_42453# a_8975_43940# 0.023559f
C7392 a_8746_45002# a_10057_43914# 0.003098f
C7393 a_8049_45260# a_22485_44484# 2.49e-20
C7394 a_4927_45028# a_6171_45002# 8.82e-20
C7395 a_9290_44172# a_11750_44172# 0.001116f
C7396 a_3218_45724# a_n2661_42834# 1.7e-20
C7397 a_10903_43370# a_10405_44172# 0.026421f
C7398 a_15765_45572# a_11827_44484# 1.86e-20
C7399 a_5147_45002# a_5205_44484# 0.018671f
C7400 a_5691_45260# a_3232_43370# 0.123939f
C7401 a_526_44458# a_2127_44172# 0.001334f
C7402 a_3815_47204# a_526_44458# 4.06e-21
C7403 a_3785_47178# a_n1925_42282# 1.46e-20
C7404 a_1123_46634# a_765_45546# 0.025395f
C7405 a_13717_47436# a_20075_46420# 3.99e-21
C7406 a_9313_45822# a_6945_45028# 0.035455f
C7407 a_13747_46662# a_11415_45002# 0.099293f
C7408 a_n881_46662# a_1138_42852# 0.148785f
C7409 a_4883_46098# a_9569_46155# 0.008675f
C7410 a_11599_46634# a_17957_46116# 0.031252f
C7411 a_n237_47217# a_6347_46155# 0.001047f
C7412 a_n971_45724# a_8781_46436# 2.04e-19
C7413 a_10623_46897# a_8270_45546# 6.27e-20
C7414 a_11453_44696# a_8016_46348# 2.61e-20
C7415 a_16241_47178# a_15682_46116# 0.001179f
C7416 a_16327_47482# a_2324_44458# 1.53e-19
C7417 a_10227_46804# a_13925_46122# 0.635045f
C7418 a_n1613_43370# a_1823_45246# 1.96e-19
C7419 a_4190_30871# a_19339_43156# 0.002519f
C7420 a_14021_43940# a_15959_42545# 4.7e-21
C7421 a_n2661_42282# a_n2302_40160# 1.84e-20
C7422 a_19095_43396# a_18083_42858# 2.56e-19
C7423 a_5649_42852# a_15567_42826# 8.45e-21
C7424 a_4361_42308# a_17595_43084# 3.75e-20
C7425 a_1568_43370# a_1576_42282# 9.29e-19
C7426 a_1049_43396# a_1184_42692# 3.77e-21
C7427 a_4905_42826# a_n784_42308# 3.17e-21
C7428 a_n1557_42282# a_n473_42460# 0.077371f
C7429 a_743_42282# a_18817_42826# 1.5e-20
C7430 a_8975_43940# VDD 0.257588f
C7431 a_n2661_45546# a_4093_43548# 0.343267f
C7432 a_13507_46334# a_21335_42336# 2.39e-19
C7433 a_n2312_38680# a_6123_31319# 4.19e-21
C7434 a_n2293_46634# a_5934_30871# 2.22e-19
C7435 a_6755_46942# a_16877_42852# 1.98e-19
C7436 a_11136_45572# a_10807_43548# 5.02e-21
C7437 a_n863_45724# a_458_43396# 0.122956f
C7438 a_13159_45002# a_13213_44734# 2.87e-19
C7439 a_9482_43914# a_n2661_43922# 0.036658f
C7440 a_3090_45724# a_9306_43218# 2.03e-20
C7441 a_9290_44172# a_4361_42308# 0.1126f
C7442 a_3357_43084# a_20512_43084# 3.36e-21
C7443 a_19479_31679# a_22485_44484# 0.001111f
C7444 a_12978_47026# a_10809_44734# 1.72e-19
C7445 a_16388_46812# a_17583_46090# 0.033313f
C7446 a_16721_46634# a_15682_46116# 0.010175f
C7447 a_n2293_46098# a_1823_45246# 0.107882f
C7448 a_10227_46804# a_15599_45572# 0.001084f
C7449 a_11599_46634# a_16020_45572# 2.63e-20
C7450 a_383_46660# a_n443_42852# 1.35e-19
C7451 a_2609_46660# a_n755_45592# 4.05e-19
C7452 a_n743_46660# a_n89_45572# 0.003687f
C7453 a_765_45546# a_13759_46122# 9.6e-20
C7454 a_3090_45724# a_n1925_42282# 0.157861f
C7455 a_16327_47482# a_16855_45546# 0.305145f
C7456 a_n2661_46634# a_4099_45572# 2.95e-20
C7457 a_12549_44172# a_7499_43078# 1.93e-19
C7458 a_12741_44636# a_3483_46348# 0.023452f
C7459 a_n2661_46098# a_1848_45724# 5.47e-21
C7460 a_1799_45572# a_2957_45546# 7.87e-21
C7461 a_n2293_46634# a_1609_45572# 1.5e-19
C7462 a_4883_46098# a_10216_45572# 5.19e-19
C7463 a_n2293_42282# a_2903_42308# 0.005938f
C7464 a_14021_43940# RST_Z 0.007254f
C7465 a_5649_42852# a_20712_42282# 1.31e-19
C7466 a_13467_32519# a_21613_42308# 0.053076f
C7467 a_13887_32519# a_13258_32519# 0.054157f
C7468 a_13678_32519# a_7174_31319# 7.78e-20
C7469 a_10083_42826# a_5742_30871# 2.48e-19
C7470 a_10835_43094# a_10723_42308# 0.006083f
C7471 a_10796_42968# a_10533_42308# 8.22e-19
C7472 a_5342_30871# a_5934_30871# 0.018148f
C7473 a_1709_42852# a_1606_42308# 4.98e-19
C7474 a_18587_45118# a_11341_43940# 1.05e-21
C7475 a_18494_42460# a_20365_43914# 0.003336f
C7476 a_18184_42460# a_20623_43914# 4.99e-21
C7477 a_21005_45260# a_19862_44208# 6.37e-19
C7478 a_n881_46662# DATA[1] 8.44e-22
C7479 a_2382_45260# a_3539_42460# 0.110439f
C7480 a_3065_45002# a_3540_43646# 9.54e-20
C7481 a_11827_44484# a_19328_44172# 0.001549f
C7482 a_20202_43084# a_17303_42282# 0.00102f
C7483 a_16237_45028# a_15682_43940# 1.42e-19
C7484 a_11691_44458# a_17973_43940# 3.47e-19
C7485 a_16147_45260# a_16409_43396# 1.28e-21
C7486 a_n863_45724# a_2987_42968# 0.002594f
C7487 a_n1925_42282# a_n2472_42282# 2.81e-19
C7488 a_n2956_39304# a_n1630_35242# 0.001241f
C7489 a_8953_45546# a_8515_42308# 6.71e-19
C7490 a_4185_45028# a_10723_42308# 1.64e-19
C7491 a_n357_42282# a_133_42852# 0.011275f
C7492 a_n1613_43370# DATA[2] 3.98e-20
C7493 a_n1059_45260# a_9396_43370# 1.51e-19
C7494 a_3232_43370# a_3080_42308# 0.001461f
C7495 a_4646_46812# a_3232_43370# 0.305673f
C7496 a_768_44030# a_n2661_43370# 0.024666f
C7497 a_4817_46660# a_5111_44636# 2.19e-22
C7498 a_4651_46660# a_5691_45260# 1.21e-20
C7499 a_4955_46873# a_4927_45028# 7.8e-21
C7500 a_3877_44458# a_6171_45002# 1.79e-21
C7501 a_5385_46902# a_5147_45002# 9.06e-21
C7502 a_16388_46812# a_8696_44636# 2.13e-19
C7503 a_13059_46348# a_15861_45028# 2.15e-21
C7504 a_19333_46634# a_19431_45546# 4.38e-20
C7505 a_15227_44166# a_19256_45572# 2.59e-20
C7506 a_6419_46155# a_6472_45840# 6.52e-19
C7507 a_4915_47217# a_15004_44636# 0.008914f
C7508 a_12741_44636# a_14495_45572# 3.7e-20
C7509 a_33_46660# a_626_44172# 1.58e-20
C7510 a_8049_45260# a_10037_46155# 4.8e-19
C7511 a_8953_45546# a_2711_45572# 0.032277f
C7512 a_19466_46812# a_18691_45572# 2.36e-19
C7513 a_n2956_39304# a_n2661_45546# 5.38e-20
C7514 a_n2956_38680# a_n2810_45572# 5.73878f
C7515 a_2905_42968# VDD 0.142081f
C7516 a_n1630_35242# a_n3565_39304# 2.9e-19
C7517 a_1606_42308# a_1239_39587# 9.67e-20
C7518 a_n3674_37592# a_n3420_39072# 0.019892f
C7519 a_6123_31319# a_7174_31319# 13.9919f
C7520 a_15764_42576# a_15959_42545# 0.21686f
C7521 COMP_P a_1736_39043# 6.78e-21
C7522 a_13575_42558# a_13921_42308# 0.013377f
C7523 a_15486_42560# a_15890_42674# 0.051162f
C7524 a_n3674_38680# a_n3565_38502# 0.128677f
C7525 a_5342_30871# a_11530_34132# 0.012973f
C7526 a_n1853_46287# DATA[0] 2.73e-20
C7527 a_895_43940# a_2455_43940# 0.01899f
C7528 a_2998_44172# a_1241_43940# 1.39e-20
C7529 a_2479_44172# a_3052_44056# 9.94e-20
C7530 a_19615_44636# a_n97_42460# 5.97e-21
C7531 a_n2661_42834# a_6293_42852# 1.51e-19
C7532 a_n2661_43922# a_6031_43396# 1.84e-20
C7533 a_20193_45348# a_13887_32519# 0.277027f
C7534 a_20820_30879# VREF 0.195875f
C7535 a_5111_44636# a_8483_43230# 1.96e-19
C7536 a_n1076_46494# VDD 0.294742f
C7537 a_10949_43914# a_12429_44172# 0.156922f
C7538 a_11823_42460# a_14456_42282# 0.004505f
C7539 a_3537_45260# a_5193_42852# 0.012016f
C7540 a_10193_42453# a_15803_42450# 3.64e-19
C7541 a_2711_45572# a_13258_32519# 0.02914f
C7542 a_n2956_38216# a_n4209_39304# 0.020992f
C7543 a_n2017_45002# a_13291_42460# 0.042872f
C7544 a_n1059_45260# a_13003_42852# 0.004401f
C7545 a_n356_44636# a_14358_43442# 3.91e-21
C7546 a_7499_43078# a_9885_42308# 0.00284f
C7547 a_11415_45002# a_18911_45144# 0.006861f
C7548 a_20202_43084# a_19778_44110# 2.92e-20
C7549 a_16327_47482# a_19862_44208# 0.209324f
C7550 a_n443_46116# a_1443_43940# 2.66e-19
C7551 w_11334_34010# a_14401_32519# 0.023412f
C7552 a_12861_44030# a_22959_43948# 1.04e-19
C7553 a_2324_44458# a_14537_43396# 0.341957f
C7554 a_2711_45572# a_8791_45572# 6.36e-19
C7555 a_10053_45546# a_10490_45724# 0.084842f
C7556 a_526_44458# a_2382_45260# 0.072916f
C7557 a_10180_45724# a_8746_45002# 0.304016f
C7558 a_3483_46348# a_n2293_42834# 0.033766f
C7559 a_3090_45724# a_18248_44752# 0.027743f
C7560 a_768_44030# a_2998_44172# 0.571981f
C7561 a_n1613_43370# a_n3674_39768# 5.31e-19
C7562 a_n2312_40392# a_n2661_42282# 3.67e-19
C7563 a_1176_45822# a_n2661_43370# 4.9e-20
C7564 a_12741_44636# a_17719_45144# 0.011019f
C7565 a_5164_46348# a_5009_45028# 4.03e-19
C7566 a_7499_43078# a_11525_45546# 1.14e-21
C7567 a_15803_42450# VDD 0.448709f
C7568 a_15764_42576# RST_Z 1.86e-19
C7569 a_13258_32519# EN_VIN_BSTR_N 0.040234f
C7570 a_5742_30871# VIN_N 0.042613f
C7571 a_22465_38105# a_22705_38406# 0.003319f
C7572 a_7174_31319# EN_VIN_BSTR_P 0.053205f
C7573 a_4958_30871# C2_P_btm 9.53e-20
C7574 a_n1741_47186# a_n1925_46634# 0.012189f
C7575 SMPL_ON_P a_n2312_38680# 0.041837f
C7576 a_n746_45260# a_n2661_46634# 0.037885f
C7577 a_4915_47217# a_768_44030# 0.187438f
C7578 a_6151_47436# a_11309_47204# 0.065131f
C7579 a_7227_47204# a_8128_46384# 3.24e-20
C7580 a_9863_47436# a_n881_46662# 0.164043f
C7581 a_20894_47436# a_13507_46334# 0.00122f
C7582 a_18780_47178# a_12465_44636# 4.89e-19
C7583 a_20990_47178# a_21177_47436# 0.159555f
C7584 a_18479_47436# a_22223_47212# 7.85e-20
C7585 a_19386_47436# a_4883_46098# 7.49e-21
C7586 a_n2109_47186# a_n743_46660# 0.029623f
C7587 a_n2288_47178# a_n2438_43548# 9.47e-19
C7588 a_15682_43940# a_743_42282# 3.41e-20
C7589 a_5343_44458# a_1606_42308# 1.12e-20
C7590 a_9313_44734# a_15785_43172# 7.07e-19
C7591 a_15493_43940# a_16664_43396# 9.17e-19
C7592 a_3905_42865# a_4520_42826# 0.054799f
C7593 a_n2661_42282# a_n2840_42826# 0.001572f
C7594 a_10193_42453# VDD 2.18892f
C7595 a_3080_42308# a_4905_42826# 0.005659f
C7596 a_1756_43548# a_1891_43646# 0.008678f
C7597 a_3422_30871# a_18083_42858# 2.69e-20
C7598 a_15493_43396# a_16823_43084# 0.029968f
C7599 a_10807_43548# a_4361_42308# 0.006525f
C7600 a_14021_43940# a_16243_43396# 0.017079f
C7601 a_17339_46660# a_18326_43940# 0.006409f
C7602 a_2063_45854# a_10991_42826# 8.1e-19
C7603 a_4791_45118# a_7871_42858# 2.66e-21
C7604 a_13661_43548# a_10341_43396# 0.053085f
C7605 a_n2293_46634# a_7221_43396# 1.49e-19
C7606 a_310_45028# a_n699_43396# 9.49e-22
C7607 a_18819_46122# a_11967_42832# 5.34e-22
C7608 a_2711_45572# a_20193_45348# 5.96e-20
C7609 a_997_45618# a_949_44458# 5.82e-20
C7610 a_n755_45592# a_2779_44458# 1.49e-20
C7611 a_15903_45785# a_16019_45002# 0.139976f
C7612 a_15765_45572# a_15595_45028# 1.18e-19
C7613 a_15599_45572# a_1307_43914# 1.34e-19
C7614 a_8696_44636# a_13777_45326# 5.73e-20
C7615 a_13507_46334# a_19095_43396# 3.23e-19
C7616 a_1823_45246# a_2675_43914# 8.17e-19
C7617 a_1848_45724# a_742_44458# 1.5e-20
C7618 a_n357_42282# a_4223_44672# 7.15e-20
C7619 a_4646_46812# a_4905_42826# 5.08e-20
C7620 a_11652_45724# a_n2661_43370# 0.028174f
C7621 a_11322_45546# a_13105_45348# 6.34e-21
C7622 a_12549_44172# a_15781_43660# 0.062935f
C7623 C0_P_btm VREF 0.443926f
C7624 a_13507_46334# a_20411_46873# 0.035522f
C7625 a_21177_47436# a_20273_46660# 0.003694f
C7626 a_20990_47178# a_20841_46902# 1.82e-19
C7627 a_20894_47436# a_20623_46660# 4.85e-19
C7628 a_17591_47464# a_17639_46660# 1.72e-19
C7629 C1_P_btm VREF_GND 0.673422f
C7630 C2_P_btm VCM 0.716172f
C7631 a_4646_46812# a_4651_46660# 0.844575f
C7632 a_n237_47217# a_8349_46414# 0.047427f
C7633 a_n971_45724# a_5937_45572# 0.027865f
C7634 a_n443_46116# a_1138_42852# 0.017807f
C7635 a_13717_47436# a_21076_30879# 5.51e-19
C7636 a_12465_44636# a_18285_46348# 2.07e-20
C7637 a_11599_46634# a_11415_45002# 0.007504f
C7638 a_3877_44458# a_4955_46873# 0.029242f
C7639 a_3524_46660# a_3633_46660# 0.007416f
C7640 a_3699_46634# a_3878_46660# 0.007399f
C7641 a_n1925_46634# a_7832_46660# 0.00149f
C7642 a_2063_45854# a_4704_46090# 0.004146f
C7643 a_3160_47472# a_3483_46348# 0.154179f
C7644 a_n1151_42308# a_3147_46376# 0.001437f
C7645 a_2905_45572# a_3699_46348# 0.004136f
C7646 a_12549_44172# a_15227_44166# 0.354423f
C7647 a_4791_45118# a_1823_45246# 0.015359f
C7648 a_5807_45002# a_12816_46660# 0.004701f
C7649 a_18479_47436# a_20731_47026# 0.004016f
C7650 a_21487_43396# a_13678_32519# 7.05e-19
C7651 a_13467_32519# a_4361_42308# 0.121732f
C7652 a_9145_43396# a_13635_43156# 0.001181f
C7653 a_10341_43396# a_10835_43094# 1.26e-19
C7654 a_7499_43078# a_7542_44172# 0.069089f
C7655 a_4185_45028# a_10341_43396# 0.019539f
C7656 a_3090_45724# a_8387_43230# 2.71e-20
C7657 a_n357_42282# a_15493_43940# 2.07e-19
C7658 a_8016_46348# a_9145_43396# 2.69e-19
C7659 a_n2956_38680# a_n1557_42282# 1.47e-20
C7660 a_3232_43370# a_10057_43914# 0.025371f
C7661 en_comp a_n356_44636# 3.08e-20
C7662 a_7229_43940# a_5883_43914# 0.026061f
C7663 a_3524_46660# a_526_44458# 4.66e-19
C7664 a_2107_46812# a_8283_46482# 5.51e-19
C7665 a_8667_46634# a_2324_44458# 8.29e-21
C7666 a_n1151_42308# a_13249_42308# 2.6e-20
C7667 a_20107_46660# a_21363_46634# 0.043567f
C7668 a_20273_46660# a_20841_46902# 0.17072f
C7669 a_20411_46873# a_20623_46660# 0.007737f
C7670 a_n1613_43370# a_n2293_45546# 0.020156f
C7671 a_n743_46660# a_8062_46155# 1.71e-19
C7672 a_8270_45546# a_8349_46414# 0.002654f
C7673 a_13607_46688# a_3483_46348# 2.14e-20
C7674 a_n971_45724# a_8697_45572# 2.34e-19
C7675 a_13747_46662# a_13259_45724# 0.093177f
C7676 a_6755_46942# a_12005_46116# 1.39e-19
C7677 a_5495_43940# VDD 0.173477f
C7678 a_2905_42968# a_n784_42308# 4.32e-21
C7679 a_5342_30871# a_16245_42852# 8.35e-20
C7680 a_15567_42826# a_15953_42852# 0.006406f
C7681 a_16243_43396# a_15764_42576# 2.19e-20
C7682 a_16137_43396# a_15803_42450# 0.002599f
C7683 a_743_42282# a_5934_30871# 0.020602f
C7684 a_5649_42852# a_6171_42473# 0.00196f
C7685 a_13678_32519# a_5932_42308# 1.17e-19
C7686 a_4743_43172# a_4649_42852# 1.26e-19
C7687 a_17333_42852# a_17141_43172# 1.97e-19
C7688 a_18083_42858# a_18504_43218# 0.088127f
C7689 a_20193_45348# a_22485_44484# 0.027057f
C7690 a_4791_45118# DATA[2] 7.19e-19
C7691 a_10193_42453# a_16137_43396# 0.329316f
C7692 a_n2012_44484# a_n2293_43922# 9.53e-19
C7693 a_n755_45592# a_n13_43084# 0.113444f
C7694 a_n863_45724# a_n967_43230# 3.46e-21
C7695 SMPL_ON_N CAL_P 0.018369f
C7696 a_12607_44458# a_13296_44484# 0.002675f
C7697 a_19479_31679# a_14401_32519# 0.053843f
C7698 a_22959_45036# a_22959_44484# 0.025171f
C7699 a_22223_45036# a_19237_31679# 7.18e-19
C7700 a_6491_46660# VDD 0.436756f
C7701 a_4700_47436# DATA[3] 3.7e-20
C7702 a_15415_45028# a_15493_43396# 2.36e-21
C7703 a_526_44458# a_1709_42852# 3.71e-19
C7704 a_12005_46116# a_8049_45260# 0.006548f
C7705 a_765_45546# a_4099_45572# 1.94e-21
C7706 a_11453_44696# a_16019_45002# 0.006638f
C7707 a_10355_46116# a_10586_45546# 0.012906f
C7708 a_9625_46129# a_9751_46155# 0.005702f
C7709 a_n2293_46098# a_n2293_45546# 0.04779f
C7710 a_3483_46348# a_16375_45002# 5.28e-20
C7711 a_768_44030# a_4574_45260# 6.09e-21
C7712 a_n2293_46634# a_n2661_45010# 0.003275f
C7713 a_n2956_39768# a_n2017_45002# 1.08e-21
C7714 a_8128_46384# a_6171_45002# 4.91e-20
C7715 a_n881_46662# a_7229_43940# 0.002123f
C7716 a_n1613_43370# a_6709_45028# 0.037165f
C7717 a_n1991_46122# a_n2661_45546# 2.49e-20
C7718 a_16137_43396# VDD 0.483673f
C7719 a_4921_42308# a_4169_42308# 9.83e-20
C7720 a_2351_42308# a_5742_30871# 1.16e-20
C7721 a_5755_42308# a_5934_30871# 2.52e-20
C7722 a_5342_30871# a_7754_40130# 7.04e-19
C7723 a_6773_42558# a_6761_42308# 0.01129f
C7724 a_1606_42308# a_12563_42308# 3.31e-20
C7725 a_5932_42308# a_6123_31319# 1.49414f
C7726 a_n2661_44458# a_8791_43396# 2.51e-20
C7727 a_5013_44260# a_5663_43940# 0.083171f
C7728 a_3537_45260# a_7227_42852# 0.002978f
C7729 a_n1059_45260# a_13635_43156# 0.006041f
C7730 a_n913_45002# a_12895_43230# 0.029875f
C7731 a_n2017_45002# a_13460_43230# 2.95e-21
C7732 a_13259_45724# a_4958_30871# 0.054732f
C7733 a_20362_44736# a_20623_43914# 0.001795f
C7734 a_20820_30879# a_22521_40599# 3.31e-20
C7735 a_15009_46634# CLK 1.39e-20
C7736 a_n357_42282# a_5742_30871# 0.001298f
C7737 a_10193_42453# a_n784_42308# 1.64e-19
C7738 a_11967_42832# a_11341_43940# 0.046075f
C7739 a_n2661_42834# a_7499_43940# 5.15e-19
C7740 a_20835_44721# a_19862_44208# 0.00122f
C7741 a_19466_46812# START 9.72e-20
C7742 a_18579_44172# a_18326_43940# 0.096332f
C7743 a_19279_43940# a_15493_43396# 0.003821f
C7744 a_19692_46634# RST_Z 3.49e-20
C7745 a_11453_44696# a_18245_44484# 1.9e-19
C7746 a_13507_46334# a_3422_30871# 0.074924f
C7747 a_18597_46090# a_20512_43084# 0.023158f
C7748 a_1823_45246# a_3429_45260# 0.047931f
C7749 a_3090_45724# a_16922_45042# 0.206138f
C7750 a_14976_45028# a_16501_45348# 7.45e-21
C7751 a_8016_46348# a_n1059_45260# 2.52e-20
C7752 a_10586_45546# a_10544_45572# 3.58e-19
C7753 a_13351_46090# a_2437_43646# 1.08e-20
C7754 a_3483_46348# a_413_45260# 5.51e-19
C7755 a_10903_43370# a_3357_43084# 9.87e-21
C7756 a_n971_45724# a_8333_44056# 0.017284f
C7757 a_12549_44172# a_12189_44484# 6.62e-21
C7758 a_13661_43548# a_n2293_43922# 7.4e-20
C7759 a_11415_45002# a_13348_45260# 0.036052f
C7760 a_8049_45260# a_14033_45822# 0.004947f
C7761 a_5066_45546# a_8696_44636# 1.84e-20
C7762 a_n4315_30879# a_n3565_38216# 0.043307f
C7763 a_1343_38525# comp_n 0.004961f
C7764 a_1736_39587# a_2112_39137# 0.269796f
C7765 a_1606_42308# C1_N_btm 0.096405f
C7766 a_n237_47217# a_10227_46804# 0.00246f
C7767 a_n784_42308# VDD 0.597561f
C7768 a_n4064_40160# a_n4209_38216# 0.047163f
C7769 a_n3420_39616# a_n4064_38528# 0.048102f
C7770 a_n4064_39616# a_n3420_38528# 0.052176f
C7771 a_n3420_39072# a_n2302_39072# 2.77e-19
C7772 a_n3565_39304# a_n3607_39392# 0.001003f
C7773 a_n2946_39072# a_n4064_39072# 0.053263f
C7774 a_n1151_42308# a_12861_44030# 0.029342f
C7775 a_4915_47217# a_9067_47204# 0.061984f
C7776 a_6545_47178# a_6851_47204# 0.134581f
C7777 a_6151_47436# a_7227_47204# 3.14e-19
C7778 a_3785_47178# a_n1435_47204# 5.76e-19
C7779 a_5932_42308# EN_VIN_BSTR_P 0.067144f
C7780 a_20692_30879# RST_Z 0.051046f
C7781 a_1241_43940# a_1568_43370# 1.38e-20
C7782 a_5829_43940# a_n97_42460# 7.1e-20
C7783 a_19963_31679# a_22775_42308# 4.22e-21
C7784 a_n1059_45260# a_18310_42308# 0.006864f
C7785 a_3422_30871# a_21855_43396# 0.005365f
C7786 a_n2661_42834# a_10991_42826# 1.88e-20
C7787 a_n2293_43922# a_10835_43094# 1.05e-20
C7788 a_10405_44172# a_8685_43396# 4.99e-20
C7789 a_20850_46155# VDD 6.25e-20
C7790 en_comp a_18727_42674# 3.94e-20
C7791 a_18184_42460# a_14097_32519# 9.17e-19
C7792 a_6298_44484# a_7309_42852# 1.49e-22
C7793 a_9313_44734# a_5534_30871# 0.039673f
C7794 a_20512_43084# a_743_42282# 0.082751f
C7795 a_2324_44458# a_n356_44636# 0.00124f
C7796 a_20202_43084# a_20159_44458# 1.9e-19
C7797 a_12741_44636# a_18588_44850# 0.002114f
C7798 a_18175_45572# a_18909_45814# 0.053479f
C7799 a_18479_45785# a_18341_45572# 0.21997f
C7800 a_16147_45260# a_18691_45572# 9.71e-20
C7801 a_526_44458# a_5343_44458# 0.015378f
C7802 a_n1925_42282# a_4743_44484# 1.27e-19
C7803 a_13661_43548# a_n97_42460# 0.02781f
C7804 a_768_44030# a_1568_43370# 0.077231f
C7805 a_16375_45002# a_17719_45144# 0.201099f
C7806 a_n2472_45546# a_n2661_43370# 0.002286f
C7807 a_10053_45546# a_6171_45002# 5.53e-21
C7808 a_10180_45724# a_3232_43370# 1.58e-19
C7809 a_6755_46942# a_15682_43940# 0.028635f
C7810 a_4185_45028# a_n2293_43922# 0.093999f
C7811 a_4419_46090# a_n2661_43922# 4.13e-20
C7812 a_13259_45724# a_18911_45144# 9.82e-20
C7813 a_5937_45572# a_9313_44734# 0.006008f
C7814 a_9290_44172# a_5891_43370# 0.302383f
C7815 a_n357_42282# a_n2293_42834# 4.06139f
C7816 a_4883_46098# a_6969_46634# 1.82e-19
C7817 a_10227_46804# a_8270_45546# 1.67e-19
C7818 a_n746_45260# a_765_45546# 0.006723f
C7819 a_13717_47436# a_15009_46634# 9.67e-21
C7820 a_12861_44030# a_14084_46812# 0.003999f
C7821 a_13487_47204# a_13607_46688# 2.07e-19
C7822 a_n1613_43370# a_5732_46660# 0.268372f
C7823 a_n1386_35608# a_n1532_35090# 0.045378f
C7824 VDAC_N C2_N_btm 1.03255f
C7825 a_11599_46634# a_12251_46660# 7.45e-20
C7826 a_n2661_46634# a_383_46660# 0.007768f
C7827 CAL_P a_19864_35138# 0.003641f
C7828 a_n2302_37690# VDD 0.350133f
C7829 a_4915_47217# a_10933_46660# 1.75e-19
C7830 a_n1151_42308# a_14180_46812# 0.037471f
C7831 a_n1925_46634# a_n743_46660# 0.193773f
C7832 a_n2312_38680# a_n2438_43548# 0.046935f
C7833 a_14955_43396# a_15231_43396# 0.00119f
C7834 a_4235_43370# a_3935_42891# 0.082011f
C7835 a_4093_43548# a_4520_42826# 0.077799f
C7836 a_3080_42308# a_2905_42968# 3.9e-20
C7837 a_n97_42460# a_10835_43094# 7.73e-20
C7838 a_n4318_39768# a_n4318_37592# 0.023201f
C7839 a_n1557_42282# a_791_42968# 0.002272f
C7840 a_453_43940# a_1606_42308# 2.97e-21
C7841 a_895_43940# a_961_42354# 7.76e-22
C7842 a_10341_43396# a_15037_43396# 1.71e-21
C7843 a_5691_45260# VDD 0.205518f
C7844 a_9313_44734# a_19647_42308# 9.5e-20
C7845 a_1414_42308# a_1755_42282# 7.59e-19
C7846 w_11334_34010# a_5934_30871# 2.35e-19
C7847 a_584_46384# a_2903_42308# 1.37e-20
C7848 a_1138_42852# a_1049_43396# 0.022078f
C7849 a_n357_42282# a_1115_44172# 0.011627f
C7850 a_n755_45592# a_644_44056# 1.74e-20
C7851 a_n913_45002# a_11827_44484# 1.54e-19
C7852 a_3877_44458# a_3681_42891# 1.24e-20
C7853 a_15227_44166# a_16977_43638# 0.002041f
C7854 a_2324_44458# a_9165_43940# 1.24e-20
C7855 a_4185_45028# a_n97_42460# 0.022167f
C7856 a_7276_45260# a_n2661_43370# 0.007354f
C7857 a_n863_45724# a_2479_44172# 0.047943f
C7858 a_16327_47482# a_20573_43172# 0.001116f
C7859 a_3090_45724# a_15743_43084# 0.005519f
C7860 a_22223_45572# a_18114_32519# 4.88e-19
C7861 a_2437_43646# a_19721_31679# 3.14e-19
C7862 a_8049_45260# a_15682_43940# 6.17e-21
C7863 a_6171_45002# a_13490_45394# 1.03e-19
C7864 a_n443_46116# a_1576_42282# 2.01e-21
C7865 a_10227_46804# a_12638_46436# 3.98e-20
C7866 a_2107_46812# a_7920_46348# 0.006995f
C7867 a_2905_45572# a_n755_45592# 0.168143f
C7868 a_14084_46812# a_14180_46812# 0.318161f
C7869 a_3090_45724# a_13885_46660# 1.72e-19
C7870 a_4883_46098# a_9241_46436# 7.71e-20
C7871 a_11599_46634# a_13259_45724# 0.249721f
C7872 a_n743_46660# a_10355_46116# 0.011802f
C7873 a_n2293_46634# a_10903_43370# 0.046902f
C7874 a_n971_45724# a_n443_42852# 0.329303f
C7875 a_2063_45854# a_2957_45546# 0.002513f
C7876 a_n746_45260# a_509_45822# 4.34e-21
C7877 a_n1151_42308# a_310_45028# 2.08e-20
C7878 a_n1613_43370# a_n914_46116# 1.68e-19
C7879 a_n881_46662# a_739_46482# 3.69e-19
C7880 a_3177_46902# a_3147_46376# 0.003463f
C7881 a_2609_46660# a_3483_46348# 0.010427f
C7882 a_2959_46660# a_2804_46116# 2.23e-19
C7883 a_768_44030# a_10809_44734# 0.037504f
C7884 a_16119_47582# a_6945_45028# 2.34e-19
C7885 a_13747_46662# a_18189_46348# 0.022348f
C7886 a_5807_45002# a_18819_46122# 0.012467f
C7887 a_14401_32519# a_13258_32519# 0.053694f
C7888 a_16795_42852# a_17701_42308# 2.09e-19
C7889 a_5111_42852# a_5193_43172# 0.003935f
C7890 a_2982_43646# a_14456_42282# 2.19e-19
C7891 a_3626_43646# a_13070_42354# 0.001839f
C7892 a_3422_30871# a_n923_35174# 0.036845f
C7893 a_n2129_44697# a_n310_44811# 8.5e-19
C7894 w_11334_34010# a_11530_34132# 37.743603f
C7895 a_20623_45572# a_20935_43940# 1.84e-19
C7896 a_10057_43914# a_8975_43940# 0.069663f
C7897 a_n1699_44726# a_n356_44636# 1.11e-20
C7898 a_n1352_44484# a_n1190_44850# 0.006453f
C7899 a_n1917_44484# a_n1655_44484# 0.001705f
C7900 a_11691_44458# a_9313_44734# 5.15e-20
C7901 a_5111_44636# a_6453_43914# 2.3e-20
C7902 a_10903_43370# a_5342_30871# 2.1e-21
C7903 a_3232_43370# a_5013_44260# 0.081759f
C7904 a_5691_45260# a_5495_43940# 3.68e-21
C7905 a_n443_42852# a_8229_43396# 2.56e-19
C7906 a_9625_46129# a_10903_43370# 1.41e-19
C7907 a_n2293_46098# a_n914_46116# 1.25e-19
C7908 a_4791_45118# a_6709_45028# 0.017539f
C7909 a_13059_46348# a_15194_46482# 6.53e-22
C7910 a_13507_46334# a_19963_31679# 1.83e-19
C7911 a_10355_46116# a_11189_46129# 0.001778f
C7912 a_5204_45822# a_2324_44458# 2.51e-21
C7913 a_10249_46116# a_2711_45572# 9.85e-22
C7914 a_2063_45854# a_9482_43914# 0.018952f
C7915 a_n1151_42308# a_11787_45002# 2.96e-21
C7916 a_22223_47212# a_2437_43646# 0.001377f
C7917 a_4883_46098# a_3357_43084# 0.060164f
C7918 a_10227_46804# a_n2017_45002# 0.030377f
C7919 a_n881_46662# a_18596_45572# 1.26e-20
C7920 a_13487_47204# a_413_45260# 4.31e-19
C7921 a_6151_47436# a_6171_45002# 0.006279f
C7922 a_19692_46634# a_21167_46155# 0.005265f
C7923 a_13747_46662# a_17478_45572# 0.073886f
C7924 a_n1991_46122# a_n1533_46116# 0.034619f
C7925 a_n971_45724# a_375_42282# 1.02e-19
C7926 a_18083_42858# a_7174_31319# 1.26e-20
C7927 a_19339_43156# a_19511_42282# 4.61e-19
C7928 a_n473_42460# a_n3674_37592# 0.054584f
C7929 a_n4318_38680# a_n3565_38502# 5.19e-20
C7930 a_3080_42308# VDD 0.849483f
C7931 a_n1329_42308# a_n1630_35242# 0.043579f
C7932 a_14537_43396# a_14579_43548# 0.046172f
C7933 a_n2956_38216# a_n4318_37592# 0.023126f
C7934 a_17715_44484# a_17303_42282# 3.11e-21
C7935 a_4223_44672# a_5025_43940# 0.002864f
C7936 a_4646_46812# VDD 2.53408f
C7937 a_n2661_43922# a_1525_44260# 1.65e-19
C7938 a_n2661_42834# a_2253_44260# 3.6e-19
C7939 a_9482_43914# a_14955_43396# 5.1e-21
C7940 a_13556_45296# a_15095_43370# 6.47e-22
C7941 a_18443_44721# a_15493_43940# 1.61e-20
C7942 a_18989_43940# a_11341_43940# 0.004444f
C7943 a_5837_45028# a_6031_43396# 5.01e-21
C7944 a_n2293_42834# a_n144_43396# 3.51e-19
C7945 a_20447_31679# a_13467_32519# 0.051601f
C7946 a_5891_43370# a_10807_43548# 1.3e-19
C7947 a_20193_45348# a_14401_32519# 0.175398f
C7948 a_18479_47436# a_9313_44734# 4.54e-21
C7949 a_526_44458# a_4880_45572# 0.02064f
C7950 a_n881_46662# a_15004_44636# 9.62e-22
C7951 a_17339_46660# a_n2017_45002# 4.48e-20
C7952 a_768_44030# a_5883_43914# 0.087568f
C7953 a_8270_45546# a_1307_43914# 0.050297f
C7954 a_11415_45002# a_20841_45814# 0.004448f
C7955 a_20202_43084# a_20623_45572# 9.54e-19
C7956 a_14513_46634# a_413_45260# 1.94e-20
C7957 a_12991_46634# a_13159_45002# 2.16e-21
C7958 a_12816_46660# a_13017_45260# 2.41e-21
C7959 a_5167_46660# a_n2661_43370# 2.93e-21
C7960 a_5066_45546# a_7227_45028# 8.68e-20
C7961 a_10809_44734# a_11652_45724# 0.073342f
C7962 a_5934_30871# a_n4064_37984# 2.14e-19
C7963 a_21335_42336# a_21613_42308# 0.110671f
C7964 a_n1630_35242# a_n3690_37440# 1.11e-19
C7965 a_n2497_47436# SMPL_ON_P 0.131317f
C7966 a_n2109_47186# a_n1920_47178# 0.070142f
C7967 a_n2288_47178# a_n1741_47186# 0.001294f
C7968 a_n3674_37592# a_n2946_37690# 4.03e-21
C7969 a_13258_32519# a_21421_42336# 7.85e-19
C7970 COMP_P a_3726_37500# 0.00602f
C7971 a_22400_42852# a_22780_40081# 1.96e-20
C7972 a_5883_43914# a_5755_42852# 6.14e-21
C7973 a_n913_45002# a_3581_42558# 0.003935f
C7974 a_n2017_45002# a_4933_42558# 0.00112f
C7975 a_n1545_46494# VDD 1.74e-19
C7976 a_2479_44172# a_3540_43646# 5.31e-20
C7977 a_9313_44734# a_4190_30871# 0.02726f
C7978 a_18184_42460# a_22959_42860# 0.004934f
C7979 a_5013_44260# a_4905_42826# 3.52e-20
C7980 a_n2661_42282# a_n2433_43396# 1.4e-20
C7981 a_11967_42832# a_10341_43396# 0.076124f
C7982 a_19321_45002# a_20365_43914# 0.006039f
C7983 a_5807_45002# a_11341_43940# 0.002004f
C7984 a_13747_46662# a_20935_43940# 2.52e-19
C7985 a_12549_44172# a_12603_44260# 0.00397f
C7986 a_768_44030# a_12495_44260# 0.001355f
C7987 a_20075_46420# a_16922_45042# 9.42e-20
C7988 a_n357_42282# a_413_45260# 0.032207f
C7989 a_n755_45592# a_n37_45144# 0.050738f
C7990 a_n863_45724# a_2680_45002# 0.024737f
C7991 a_12741_44636# a_18443_44721# 0.002904f
C7992 a_15227_44166# a_17061_44734# 0.07208f
C7993 a_n2293_46634# a_14955_43940# 0.004724f
C7994 a_18479_47436# a_20974_43370# 0.008175f
C7995 a_5066_45546# a_5009_45028# 1.52e-19
C7996 a_12594_46348# a_11691_44458# 4.78e-21
C7997 a_7920_46348# a_n2661_44458# 4.63e-21
C7998 a_310_45028# a_327_44734# 0.006962f
C7999 a_13163_45724# a_13385_45572# 0.001684f
C8000 a_n443_42852# a_n2293_45010# 0.003134f
C8001 a_18597_46090# a_21381_43940# 0.080234f
C8002 a_10193_42453# a_18479_45785# 1.12e-19
C8003 a_n2293_45546# a_3429_45260# 3.77e-21
C8004 a_n2661_45546# a_4558_45348# 0.050441f
C8005 a_18189_46348# a_18911_45144# 1.91e-19
C8006 a_13259_45724# a_13348_45260# 0.016055f
C8007 a_n237_47217# a_10467_46802# 2.29e-19
C8008 a_2063_45854# a_7715_46873# 0.178294f
C8009 a_6851_47204# a_3877_44458# 8.01e-20
C8010 a_n1435_47204# a_3699_46634# 5.5e-20
C8011 a_6491_46660# a_4646_46812# 0.042695f
C8012 a_3754_38470# a_8912_37509# 1.88278f
C8013 a_4791_45118# a_5732_46660# 4.55e-19
C8014 a_5129_47502# a_5385_46902# 0.001505f
C8015 a_5815_47464# a_4817_46660# 0.00304f
C8016 a_9804_47204# a_10037_47542# 5.76e-19
C8017 a_n881_46662# a_768_44030# 0.057002f
C8018 a_n2946_39072# VDD 0.383374f
C8019 a_7754_38470# a_6886_37412# 0.180842f
C8020 a_4883_46098# a_n2293_46634# 0.046481f
C8021 a_n3420_39616# VREF_GND 0.117023f
C8022 a_11453_44696# a_22612_30879# 0.005655f
C8023 a_22959_47212# a_21588_30879# 0.018188f
C8024 a_n3420_37440# a_n4251_37440# 0.001432f
C8025 a_n4064_37440# a_n2860_37690# 0.003766f
C8026 a_n3690_37440# a_n3607_37440# 0.007692f
C8027 a_8530_39574# a_5700_37509# 0.947638f
C8028 a_n4209_38216# C10_P_btm 2.25e-20
C8029 en_comp a_22521_39511# 0.008551f
C8030 a_8791_43396# a_9145_43396# 0.092458f
C8031 a_18479_45785# VDD 0.536075f
C8032 a_14539_43914# a_14456_42282# 5.4e-20
C8033 a_14955_43940# a_5342_30871# 1.82e-19
C8034 a_n356_44636# a_9803_42558# 1.46e-19
C8035 a_21381_43940# a_743_42282# 4.2e-21
C8036 a_20974_43370# a_4190_30871# 0.214288f
C8037 a_n1613_43370# a_7227_42852# 0.007002f
C8038 a_n443_42852# a_9313_44734# 0.02484f
C8039 a_n1925_42282# a_1414_42308# 5.84e-21
C8040 a_3537_45260# a_7229_43940# 1.13e-19
C8041 a_n2017_45002# a_1307_43914# 0.001015f
C8042 a_8270_45546# a_9396_43370# 8.62e-19
C8043 a_22612_30879# a_17364_32525# 0.062457f
C8044 a_10193_42453# a_10057_43914# 4.92e-20
C8045 a_8746_45002# a_10440_44484# 0.027688f
C8046 a_10180_45724# a_8975_43940# 6.79e-20
C8047 a_15037_45618# a_11691_44458# 1.37e-19
C8048 a_8049_45260# a_20512_43084# 5.74e-21
C8049 a_5111_44636# a_6171_45002# 3.76e-19
C8050 a_4927_45028# a_3232_43370# 1.34e-20
C8051 a_9290_44172# a_10807_43548# 0.364112f
C8052 a_4791_45118# a_5193_42852# 0.004916f
C8053 a_n2293_45010# a_375_42282# 0.021456f
C8054 a_n2661_45010# a_626_44172# 0.0195f
C8055 a_15903_45785# a_11827_44484# 3.96e-21
C8056 a_12465_44636# a_5534_30871# 1.02e-21
C8057 a_526_44458# a_453_43940# 0.028123f
C8058 a_3785_47178# a_526_44458# 2.7e-22
C8059 a_383_46660# a_765_45546# 1.21e-19
C8060 a_13717_47436# a_19335_46494# 1.62e-21
C8061 a_11031_47542# a_6945_45028# 0.007285f
C8062 a_13661_43548# a_11415_45002# 0.107787f
C8063 a_13747_46662# a_20202_43084# 0.308003f
C8064 a_n881_46662# a_1176_45822# 0.048496f
C8065 a_n1613_43370# a_1138_42852# 1.35e-19
C8066 a_4883_46098# a_9625_46129# 0.164961f
C8067 a_11599_46634# a_18189_46348# 0.101491f
C8068 a_n237_47217# a_8034_45724# 0.0717f
C8069 a_10467_46802# a_8270_45546# 3.96e-20
C8070 a_6755_46942# a_6903_46660# 0.003896f
C8071 a_10428_46928# a_10384_47026# 1.46e-19
C8072 a_16327_47482# a_14840_46494# 6.83e-21
C8073 a_15673_47210# a_15682_46116# 6.62e-20
C8074 a_10227_46804# a_13759_46122# 0.920747f
C8075 a_n97_42460# a_n39_42308# 0.001449f
C8076 a_15493_43396# a_19332_42282# 3.15e-19
C8077 a_4190_30871# a_18599_43230# 0.008694f
C8078 a_14021_43940# a_15803_42450# 1.55e-20
C8079 a_15493_43940# a_15521_42308# 2.45e-20
C8080 a_n2661_42282# a_n4064_40160# 4.6e-21
C8081 a_5649_42852# a_5342_30871# 0.091782f
C8082 a_4361_42308# a_16795_42852# 2.38e-20
C8083 a_13887_32519# a_5534_30871# 0.047233f
C8084 a_458_43396# a_961_42354# 4.08e-20
C8085 a_1209_43370# a_1184_42692# 0.001053f
C8086 a_743_42282# a_18249_42858# 4.69e-20
C8087 a_1847_42826# a_3681_42891# 8.84e-21
C8088 a_2075_43172# a_2905_42968# 0.023236f
C8089 a_10057_43914# VDD 0.399284f
C8090 a_3080_42308# a_n784_42308# 0.170007f
C8091 a_n1557_42282# a_n961_42308# 0.041329f
C8092 a_4646_46812# a_n784_42308# 4.29e-21
C8093 a_3090_45724# a_9061_43230# 3.86e-21
C8094 a_10193_42453# a_14021_43940# 0.033291f
C8095 a_n755_45592# a_104_43370# 0.029812f
C8096 a_13507_46334# a_7174_31319# 0.041342f
C8097 a_18597_46090# a_21125_42558# 0.002227f
C8098 a_17339_46660# a_19164_43230# 9.04e-20
C8099 a_n2442_46660# a_5934_30871# 7.2e-21
C8100 a_11827_44484# a_n2661_44458# 0.003582f
C8101 a_10903_43370# a_743_42282# 0.029178f
C8102 a_n2293_46634# a_7963_42308# 2.47e-20
C8103 a_n2017_45002# a_18579_44172# 3.84e-19
C8104 a_20193_45348# a_20205_45028# 0.012189f
C8105 a_9482_43914# a_n2661_42834# 0.076592f
C8106 a_n863_45724# a_n229_43646# 4.39e-19
C8107 a_n2293_46634# a_1260_45572# 6.07e-19
C8108 a_16388_46812# a_15682_46116# 0.044769f
C8109 a_11415_45002# a_4185_45028# 5.21e-19
C8110 a_n971_45724# a_2437_43646# 0.204278f
C8111 a_11599_46634# a_17478_45572# 0.025658f
C8112 a_2443_46660# a_n755_45592# 5.37e-20
C8113 a_3090_45724# a_526_44458# 0.058033f
C8114 a_n2293_46098# a_1138_42852# 0.029886f
C8115 a_n881_46662# a_11652_45724# 4.56e-21
C8116 a_16327_47482# a_16115_45572# 0.163022f
C8117 a_n2661_46098# a_997_45618# 4.98e-22
C8118 a_8270_45546# a_8034_45724# 0.031124f
C8119 a_768_44030# a_8162_45546# 2.17e-21
C8120 a_765_45546# a_13351_46090# 9.37e-21
C8121 a_n1423_46090# a_472_46348# 3.09e-21
C8122 a_n901_46420# a_n1076_46494# 0.234322f
C8123 a_1799_45572# a_1848_45724# 0.080562f
C8124 a_4883_46098# a_9159_45572# 6.4e-19
C8125 a_n2293_42282# a_2713_42308# 0.002882f
C8126 a_14021_43940# VDD 1.60583f
C8127 a_13467_32519# a_21887_42336# 0.011781f
C8128 a_10518_42984# a_10723_42308# 6.75e-19
C8129 a_16328_43172# a_16245_42852# 1.48e-19
C8130 a_5649_42852# a_20107_42308# 1.31e-19
C8131 a_4361_42308# a_21335_42336# 0.013772f
C8132 a_743_42282# a_21125_42558# 3.76e-20
C8133 a_8953_45546# a_5934_30871# 0.113715f
C8134 a_4185_45028# a_10533_42308# 9.41e-20
C8135 a_17613_45144# a_15493_43940# 4.03e-21
C8136 a_18494_42460# a_20269_44172# 0.017863f
C8137 a_18184_42460# a_20365_43914# 2.05e-19
C8138 a_19778_44110# a_20623_43914# 3.52e-20
C8139 a_n881_46662# DATA[0] 0.003238f
C8140 a_3065_45002# a_2982_43646# 0.026494f
C8141 a_2382_45260# a_3626_43646# 0.041715f
C8142 a_n1613_43370# DATA[1] 7.06e-20
C8143 a_11827_44484# a_18451_43940# 0.006619f
C8144 a_n2956_38680# a_n3674_37592# 0.026013f
C8145 a_n2293_43922# a_11967_42832# 0.022597f
C8146 a_11691_44458# a_17737_43940# 1.76e-19
C8147 a_n863_45724# a_1793_42852# 5.96e-19
C8148 a_n2017_45002# a_9396_43370# 3.4e-20
C8149 a_n1059_45260# a_8791_43396# 0.196029f
C8150 a_n913_45002# a_8147_43396# 7.89e-20
C8151 a_5883_43914# a_7845_44172# 0.02286f
C8152 a_3232_43370# a_4699_43561# 9.73e-20
C8153 a_9804_47204# VDD 0.410522f
C8154 a_n2956_38680# a_n2840_45546# 2.65e-20
C8155 a_n2956_39304# a_n2810_45572# 0.043323f
C8156 a_4817_46660# a_5147_45002# 6.83e-20
C8157 a_3877_44458# a_3232_43370# 0.016642f
C8158 a_4646_46812# a_5691_45260# 1.06e-21
C8159 a_12549_44172# a_n2661_43370# 3e-20
C8160 a_13059_46348# a_8696_44636# 0.020156f
C8161 a_15227_44166# a_19431_45546# 2.07e-20
C8162 a_18479_47436# a_18114_32519# 3.09e-20
C8163 a_4915_47217# a_13720_44458# 0.006519f
C8164 a_12741_44636# a_13249_42308# 0.028381f
C8165 a_3090_45724# a_17668_45572# 0.071363f
C8166 a_11453_44696# a_11827_44484# 0.170003f
C8167 a_12465_44636# a_11691_44458# 0.15589f
C8168 a_2324_44458# a_3503_45724# 9.33e-22
C8169 a_8049_45260# a_9751_46155# 4.35e-19
C8170 a_5937_45572# a_2711_45572# 0.063757f
C8171 a_n746_45260# a_700_44734# 0.009437f
C8172 a_4651_46660# a_4927_45028# 5.26e-21
C8173 a_n2438_43548# a_1423_45028# 0.242599f
C8174 a_19466_46812# a_18909_45814# 0.001786f
C8175 a_n3674_38680# a_n4334_38528# 0.05024f
C8176 a_5534_30871# EN_VIN_BSTR_N 0.007335f
C8177 a_2075_43172# VDD 0.001106f
C8178 a_15764_42576# a_15803_42450# 0.901878f
C8179 a_7227_42308# a_7174_31319# 9.76e-21
C8180 COMP_P a_1239_39043# 0.001354f
C8181 a_5934_30871# a_13258_32519# 7.32e-19
C8182 a_13575_42558# a_13657_42308# 0.003935f
C8183 a_15486_42560# a_15959_42545# 7.99e-20
C8184 a_n356_44636# a_14579_43548# 5.95e-21
C8185 a_5891_43370# a_5837_43396# 1.86e-19
C8186 a_2479_44172# a_2455_43940# 0.025354f
C8187 a_895_43940# a_2253_43940# 0.053882f
C8188 a_11967_42832# a_n97_42460# 0.489711f
C8189 a_n2661_42834# a_6031_43396# 1.34e-19
C8190 a_20193_45348# a_22223_43396# 0.020364f
C8191 a_21076_30879# EN_OFFSET_CAL 0.2809f
C8192 a_1414_42308# a_3737_43940# 1.01e-19
C8193 a_n901_46420# VDD 0.518805f
C8194 a_10949_43914# a_11750_44172# 0.05299f
C8195 a_10729_43914# a_12429_44172# 1.01e-19
C8196 a_11823_42460# a_13575_42558# 0.075921f
C8197 a_3537_45260# a_4649_42852# 0.065656f
C8198 a_18989_43940# a_10341_43396# 2.68e-19
C8199 a_10193_42453# a_15764_42576# 2.52e-19
C8200 a_2711_45572# a_19647_42308# 0.046367f
C8201 a_n2810_45572# a_n3565_39304# 0.030572f
C8202 a_20820_30879# VIN_N 0.049556f
C8203 a_n2293_42834# a_8952_43230# 1.55e-19
C8204 a_7499_43078# a_11322_45546# 8.22e-21
C8205 a_22612_30879# a_19237_31679# 0.062542f
C8206 a_11415_45002# a_18587_45118# 0.005313f
C8207 a_12861_44030# a_15493_43940# 0.370814f
C8208 a_n443_46116# a_1241_43940# 1.44e-19
C8209 a_15015_46420# a_14797_45144# 2.32e-20
C8210 a_2324_44458# a_14180_45002# 0.026932f
C8211 a_6945_45028# a_6709_45028# 0.060282f
C8212 a_2711_45572# a_8697_45572# 3.48e-19
C8213 a_10053_45546# a_8746_45002# 0.075884f
C8214 a_10180_45724# a_10193_42453# 0.145672f
C8215 a_526_44458# a_2274_45254# 0.019853f
C8216 a_3090_45724# a_17970_44736# 1.26e-19
C8217 a_768_44030# a_2889_44172# 0.011283f
C8218 a_n1613_43370# a_n4318_39768# 1.98e-19
C8219 a_16327_47482# a_19478_44306# 3.2e-19
C8220 a_9049_44484# a_10490_45724# 1.71e-20
C8221 a_518_46155# a_413_45260# 3.64e-20
C8222 a_12741_44636# a_17613_45144# 0.006096f
C8223 a_4883_46098# a_9672_43914# 0.009886f
C8224 a_19787_47423# a_13507_46334# 5.57e-21
C8225 a_18597_46090# a_4883_46098# 0.084375f
C8226 a_15764_42576# VDD 0.258303f
C8227 a_15486_42560# RST_Z 5.88e-19
C8228 a_5742_30871# VIN_P 0.042613f
C8229 a_13258_32519# a_11530_34132# 0.002091f
C8230 a_n2109_47186# a_n1021_46688# 1.8e-21
C8231 a_n1920_47178# a_n1925_46634# 0.013665f
C8232 a_n4064_39072# a_n4064_37440# 0.046264f
C8233 a_22465_38105# a_22609_38406# 0.20695f
C8234 SMPL_ON_P a_n2104_46634# 3.11e-20
C8235 a_n971_45724# a_n2661_46634# 0.190714f
C8236 a_n443_46116# a_768_44030# 0.177051f
C8237 a_4915_47217# a_12549_44172# 0.316329f
C8238 a_9067_47204# a_n881_46662# 0.073421f
C8239 a_6575_47204# a_7989_47542# 6.62e-20
C8240 a_18479_47436# a_12465_44636# 7.24e-19
C8241 a_n2497_47436# a_n2438_43548# 0.206216f
C8242 a_7174_31319# a_n923_35174# 0.007133f
C8243 a_4958_30871# C3_P_btm 1.05e-19
C8244 en_comp a_1177_38525# 0.205977f
C8245 a_14955_43940# a_743_42282# 1.64e-22
C8246 a_9313_44734# a_14635_42282# 0.005265f
C8247 a_15493_43940# a_19700_43370# 5.37e-20
C8248 a_3905_42865# a_3935_42891# 0.240349f
C8249 a_10180_45724# VDD 0.336512f
C8250 a_19279_43940# a_21356_42826# 2.54e-19
C8251 a_18579_44172# a_19164_43230# 5.37e-20
C8252 a_3422_30871# a_17701_42308# 2.82e-20
C8253 a_14021_43940# a_16137_43396# 0.002723f
C8254 a_4699_43561# a_4905_42826# 1.43e-19
C8255 a_1568_43370# a_1891_43646# 7.4e-19
C8256 a_n97_42460# a_648_43396# 0.00481f
C8257 a_16147_45260# a_6171_45002# 0.072853f
C8258 a_2063_45854# a_10796_42968# 7.47e-21
C8259 a_5807_45002# a_10341_43396# 1.82e-19
C8260 a_n2293_46634# a_8685_43396# 0.335608f
C8261 a_15227_44166# a_15301_44260# 0.003263f
C8262 a_5257_43370# a_n97_42460# 0.167676f
C8263 a_16115_45572# a_14537_43396# 3.42e-21
C8264 a_2711_45572# a_11691_44458# 0.058464f
C8265 a_11322_45546# a_11915_45394# 3.21e-19
C8266 a_167_45260# a_2127_44172# 3.83e-20
C8267 a_22959_45572# a_20447_31679# 0.154273f
C8268 a_n755_45592# a_949_44458# 0.011024f
C8269 a_n357_42282# a_2779_44458# 8.49e-21
C8270 a_15599_45572# a_16019_45002# 0.001742f
C8271 a_15903_45785# a_15595_45028# 0.003784f
C8272 a_8696_44636# a_13556_45296# 0.022968f
C8273 a_13507_46334# a_21487_43396# 4.46e-21
C8274 a_4883_46098# a_743_42282# 1.38e-19
C8275 a_18597_46090# a_5649_42852# 9.18e-20
C8276 a_1823_45246# a_895_43940# 1.63e-20
C8277 a_4646_46812# a_3080_42308# 2.88e-19
C8278 a_18051_46116# a_17767_44458# 5.87e-22
C8279 a_12549_44172# a_15681_43442# 0.080982f
C8280 C1_P_btm VREF 0.98698f
C8281 a_13507_46334# a_20107_46660# 0.031344f
C8282 a_20990_47178# a_20273_46660# 1.7e-19
C8283 a_20894_47436# a_20841_46902# 2.44e-19
C8284 C2_P_btm VREF_GND 0.671742f
C8285 C3_P_btm VCM 0.716273f
C8286 a_3877_44458# a_4651_46660# 0.032518f
C8287 a_n971_45724# a_8199_44636# 0.247183f
C8288 a_n237_47217# a_8016_46348# 0.017823f
C8289 a_n443_46116# a_1176_45822# 0.092452f
C8290 a_9804_47204# a_10185_46660# 4.55e-19
C8291 a_n1925_46634# a_6086_46660# 2.66e-19
C8292 C0_dummy_P_btm VIN_P 0.544204f
C8293 a_2063_45854# a_4419_46090# 0.025095f
C8294 a_3160_47472# a_3147_46376# 0.208295f
C8295 a_2905_45572# a_3483_46348# 0.024106f
C8296 a_12549_44172# a_18834_46812# 0.01219f
C8297 a_5807_45002# a_12991_46634# 0.006904f
C8298 a_4700_47436# a_1823_45246# 1.11e-20
C8299 a_12861_44030# a_12741_44636# 0.366155f
C8300 a_n1741_47186# a_9823_46155# 1.05e-20
C8301 a_4883_46098# a_19123_46287# 0.022559f
C8302 a_3422_30871# a_21613_42308# 0.027998f
C8303 a_21487_43396# a_21855_43396# 7.52e-19
C8304 a_14579_43548# a_12379_42858# 2.62e-21
C8305 a_20512_43084# a_13258_32519# 2.41e-19
C8306 a_4190_30871# a_13887_32519# 0.032018f
C8307 a_743_42282# a_5649_42852# 0.030921f
C8308 a_8685_43396# a_5342_30871# 0.001246f
C8309 a_10341_43396# a_10518_42984# 5.04e-20
C8310 a_n467_45028# a_n2012_44484# 9.72e-23
C8311 a_8162_45546# a_7845_44172# 1.27e-21
C8312 a_7499_43078# a_7281_43914# 6.26e-21
C8313 a_7705_45326# a_6298_44484# 0.004597f
C8314 a_n2956_39304# a_n1557_42282# 1.75e-20
C8315 a_3232_43370# a_10440_44484# 0.042872f
C8316 a_12465_44636# a_n443_42852# 1.42e-19
C8317 a_3699_46634# a_526_44458# 1.66e-21
C8318 a_2107_46812# a_8062_46482# 2.73e-19
C8319 a_n1151_42308# a_13904_45546# 1.84e-19
C8320 a_20107_46660# a_20623_46660# 0.105914f
C8321 a_5732_46660# a_6945_45028# 1.4e-20
C8322 a_8270_45546# a_8016_46348# 0.036831f
C8323 a_6151_47436# a_8746_45002# 8.1e-20
C8324 a_12816_46660# a_3483_46348# 8.76e-22
C8325 a_n971_45724# a_8192_45572# 0.005205f
C8326 a_13747_46662# a_14383_46116# 2.43e-19
C8327 a_13661_43548# a_13259_45724# 0.250875f
C8328 a_6755_46942# a_10903_43370# 1.97e-19
C8329 a_n2661_46634# a_12005_46436# 8.72e-20
C8330 a_n1925_46634# a_8379_46155# 2.63e-19
C8331 a_18479_47436# a_2711_45572# 1.11e-19
C8332 a_5013_44260# VDD 0.198233f
C8333 a_685_42968# a_564_42282# 3.6e-19
C8334 a_15567_42826# a_15597_42852# 0.025037f
C8335 a_5342_30871# a_15953_42852# 5.76e-19
C8336 a_16137_43396# a_15764_42576# 0.008757f
C8337 a_5649_42852# a_5755_42308# 0.008092f
C8338 a_16409_43396# a_14113_42308# 1.57e-21
C8339 a_4649_43172# a_4649_42852# 6.96e-20
C8340 a_743_42282# a_7963_42308# 0.008222f
C8341 a_20193_45348# a_20512_43084# 0.160912f
C8342 a_4700_47436# DATA[2] 0.001637f
C8343 a_6151_47436# RST_Z 0.010195f
C8344 a_n1151_42308# CLK 0.022274f
C8345 a_n443_46116# DATA[0] 4.31e-19
C8346 a_8375_44464# a_5891_43370# 0.094782f
C8347 a_n2012_44484# a_n2661_43922# 0.00414f
C8348 a_2711_45572# a_4190_30871# 0.051595f
C8349 a_n357_42282# a_n13_43084# 0.194173f
C8350 a_n755_45592# a_n1076_43230# 2.49e-20
C8351 a_n863_45724# a_n1379_43218# 3.89e-21
C8352 a_12607_44458# a_12829_44484# 5.19e-19
C8353 a_n2293_42834# a_n1441_43940# 0.001195f
C8354 a_11827_44484# a_19237_31679# 3.81e-19
C8355 a_6545_47178# VDD 0.386368f
C8356 a_10903_43370# a_8049_45260# 0.114138f
C8357 a_19692_46634# a_10193_42453# 0.010323f
C8358 a_10185_46660# a_10180_45724# 7.92e-20
C8359 a_11453_44696# a_15595_45028# 0.007267f
C8360 a_n2472_46090# a_n2293_45546# 3.06e-19
C8361 a_n2293_46098# a_n2956_38216# 0.003979f
C8362 a_15368_46634# a_11823_42460# 0.014491f
C8363 a_768_44030# a_3537_45260# 0.341201f
C8364 a_n2442_46660# a_n2661_45010# 1.33e-20
C8365 a_n2293_46634# a_n2840_45002# 7.08e-19
C8366 a_8128_46384# a_3232_43370# 1.19e-20
C8367 a_n881_46662# a_7276_45260# 4.09e-20
C8368 a_n1613_43370# a_7229_43940# 0.059621f
C8369 a_n1853_46287# a_n2661_45546# 0.004849f
C8370 a_4185_45028# a_13259_45724# 0.194989f
C8371 a_4190_30871# EN_VIN_BSTR_N 0.043599f
C8372 a_2123_42473# a_5742_30871# 1.16e-20
C8373 a_4921_42308# a_3905_42308# 6.09e-20
C8374 a_6171_42473# a_6123_31319# 8.95e-21
C8375 a_5932_42308# a_7227_42308# 1.68e-20
C8376 a_19333_46634# START 3.38e-20
C8377 a_5013_44260# a_5495_43940# 0.251039f
C8378 a_3537_45260# a_5755_42852# 0.088502f
C8379 a_15227_44166# SINGLE_ENDED 3.5e-21
C8380 a_n443_42852# a_8515_42308# 2.59e-21
C8381 a_n2017_45002# a_13635_43156# 4.66e-19
C8382 a_n913_45002# a_13113_42826# 0.018663f
C8383 a_n1059_45260# a_12895_43230# 0.003645f
C8384 a_n2956_38680# a_n2302_39072# 2.87e-19
C8385 a_20362_44736# a_20365_43914# 0.012553f
C8386 a_20159_44458# a_20623_43914# 0.005333f
C8387 a_5343_44458# a_3626_43646# 0.001955f
C8388 a_742_44458# a_648_43396# 6.39e-22
C8389 a_5244_44056# a_5663_43940# 7.46e-20
C8390 a_n357_42282# a_11323_42473# 7.85e-20
C8391 a_11827_44484# a_9145_43396# 6.87e-20
C8392 a_n2661_42834# a_6671_43940# 6.64e-19
C8393 a_20679_44626# a_19862_44208# 0.001682f
C8394 a_19692_46634# VDD 2.53528f
C8395 a_19279_43940# a_19328_44172# 0.120319f
C8396 a_18579_44172# a_18079_43940# 3.67e-19
C8397 a_18989_43940# a_n97_42460# 1.52e-19
C8398 a_19466_46812# RST_Z 2.04e-20
C8399 a_11453_44696# a_18005_44484# 1e-19
C8400 a_13507_46334# a_21398_44850# 2.03e-20
C8401 a_18597_46090# a_21145_44484# 0.001307f
C8402 a_n1925_46634# a_5891_43370# 1.42e-20
C8403 a_1823_45246# a_3065_45002# 0.607468f
C8404 a_14976_45028# a_16405_45348# 1.42e-20
C8405 a_8016_46348# a_n2017_45002# 2.05e-20
C8406 a_10586_45546# a_10306_45572# 1.95e-19
C8407 a_3147_46376# a_413_45260# 0.015235f
C8408 a_12594_46348# a_2437_43646# 3.38e-20
C8409 a_167_45260# a_2382_45260# 0.002522f
C8410 a_n1151_42308# a_n630_44306# 0.001084f
C8411 a_n881_46662# a_17517_44484# 2.63e-20
C8412 a_768_44030# a_11541_44484# 0.003356f
C8413 a_11415_45002# a_13159_45002# 0.141106f
C8414 a_1609_45822# a_1609_45572# 0.009518f
C8415 a_n443_42852# a_2711_45572# 9.23e-22
C8416 a_2063_45854# a_11599_46634# 0.19861f
C8417 a_n3565_39590# a_n2302_38778# 8.95e-20
C8418 a_1343_38525# a_1736_39043# 0.310247f
C8419 a_1606_42308# C0_N_btm 0.029189f
C8420 a_196_42282# VDD 0.291844f
C8421 a_n4064_40160# a_n3607_38528# 5.58e-20
C8422 a_n3420_39072# a_n4064_39072# 4.93427f
C8423 a_n1151_42308# a_13717_47436# 2.89e-19
C8424 a_4915_47217# a_6575_47204# 0.849579f
C8425 a_6151_47436# a_6851_47204# 0.007871f
C8426 a_6545_47178# a_6491_46660# 0.181574f
C8427 a_3381_47502# a_n1435_47204# 4.12e-19
C8428 a_5932_42308# a_n923_35174# 0.006295f
C8429 a_20205_31679# RST_Z 0.049474f
C8430 a_20512_43084# a_20301_43646# 2.11e-20
C8431 a_1241_43940# a_1049_43396# 3.88e-19
C8432 a_19319_43548# a_18533_43940# 2.47e-20
C8433 a_5745_43940# a_n97_42460# 8.52e-20
C8434 a_n1059_45260# a_18220_42308# 0.00103f
C8435 a_n2293_43922# a_10518_42984# 5.88e-21
C8436 a_n2661_42834# a_10796_42968# 6.58e-21
C8437 a_n2661_43370# a_n1630_35242# 2.37e-20
C8438 a_9672_43914# a_8685_43396# 3.33e-20
C8439 en_comp a_18057_42282# 2.2e-20
C8440 a_20692_30879# VDD 0.499615f
C8441 a_18184_42460# a_22400_42852# 0.16156f
C8442 a_9313_44734# a_14543_43071# 0.00414f
C8443 a_3422_30871# a_4361_42308# 0.096125f
C8444 a_4099_45572# a_1307_43914# 1.48e-22
C8445 a_3316_45546# a_2809_45028# 9.97e-20
C8446 a_18175_45572# a_18341_45572# 0.577068f
C8447 a_16147_45260# a_18909_45814# 3.16e-20
C8448 a_526_44458# a_4743_44484# 5.55e-19
C8449 a_5807_45002# a_n97_42460# 1.62e-22
C8450 a_768_44030# a_1049_43396# 5.52e-20
C8451 a_16375_45002# a_17613_45144# 0.040514f
C8452 a_n2661_45546# a_n2661_43370# 0.145941f
C8453 a_11415_45002# a_11967_42832# 0.007699f
C8454 a_6755_46942# a_14955_43940# 0.00126f
C8455 a_4185_45028# a_n2661_43922# 0.022579f
C8456 a_9049_44484# a_6171_45002# 0.026882f
C8457 a_5937_45572# a_9241_44734# 9.79e-19
C8458 a_8199_44636# a_9313_44734# 0.016063f
C8459 a_13259_45724# a_18587_45118# 0.099974f
C8460 a_n1925_42282# a_n699_43396# 0.024581f
C8461 a_4883_46098# a_6755_46942# 0.060162f
C8462 a_n1925_46634# a_n1021_46688# 0.011448f
C8463 a_n2293_46634# a_n133_46660# 1.8e-21
C8464 a_n2104_46634# a_n2438_43548# 0.052991f
C8465 a_n971_45724# a_765_45546# 0.140618f
C8466 a_n881_46662# a_5167_46660# 7.84e-21
C8467 a_12861_44030# a_13607_46688# 0.019182f
C8468 a_n1613_43370# a_5907_46634# 0.338694f
C8469 CAL_P a_19120_35138# 0.00106f
C8470 a_n1838_35608# a_n1532_35090# 4.88e-19
C8471 VDAC_N C1_N_btm 0.55675f
C8472 a_11599_46634# a_12469_46902# 9.01e-21
C8473 a_n2661_46634# a_601_46902# 0.009214f
C8474 a_n4064_37440# VDD 1.65981f
C8475 a_n1151_42308# a_14035_46660# 0.026112f
C8476 a_n2312_38680# a_n743_46660# 0.001509f
C8477 a_14955_43396# a_15125_43396# 0.001675f
C8478 a_15095_43370# a_15231_43396# 0.001002f
C8479 a_4093_43548# a_3935_42891# 0.00342f
C8480 a_n97_42460# a_10518_42984# 1.55e-20
C8481 a_14401_32519# a_5534_30871# 0.339008f
C8482 a_4235_43370# a_3681_42891# 7.84e-21
C8483 a_8685_43396# a_743_42282# 1.88e-19
C8484 a_n1557_42282# a_685_42968# 0.003946f
C8485 a_895_43940# a_1184_42692# 2.55e-21
C8486 a_n3674_39768# a_n3674_38216# 0.02323f
C8487 a_4927_45028# VDD 0.159822f
C8488 a_15781_43660# a_16409_43396# 2.7e-19
C8489 a_10341_43396# a_16867_43762# 0.001683f
C8490 a_1414_42308# a_1606_42308# 0.056716f
C8491 a_9313_44734# a_19511_42282# 0.001387f
C8492 a_1138_42852# a_1209_43370# 0.01435f
C8493 a_n357_42282# a_644_44056# 0.007544f
C8494 a_n755_45592# a_175_44278# 0.01086f
C8495 en_comp a_18494_42460# 6.64e-20
C8496 a_n1059_45260# a_11827_44484# 9.98e-20
C8497 a_15227_44166# a_16409_43396# 0.003488f
C8498 a_13904_45546# a_13857_44734# 4.52e-21
C8499 a_13249_42308# a_13468_44734# 2.67e-20
C8500 a_5205_44484# a_n2661_43370# 0.033807f
C8501 a_8953_45002# a_8560_45348# 0.001921f
C8502 a_10586_45546# a_10729_43914# 2.76e-22
C8503 a_16327_47482# a_20256_43172# 0.054992f
C8504 a_21513_45002# a_19721_31679# 9.71e-20
C8505 a_n2661_45546# a_2998_44172# 0.060624f
C8506 a_6171_45002# a_13105_45348# 5.33e-20
C8507 a_11652_45724# a_11541_44484# 1.11e-20
C8508 a_13059_46348# a_14205_43396# 0.049915f
C8509 a_10227_46804# a_12379_46436# 0.001273f
C8510 a_n2661_46634# a_12594_46348# 7.33e-20
C8511 a_2107_46812# a_6419_46155# 0.007575f
C8512 a_13607_46688# a_14180_46812# 5.9e-19
C8513 a_14084_46812# a_14035_46660# 0.086342f
C8514 a_12816_46660# a_14513_46634# 1.47e-20
C8515 a_15009_46634# a_13885_46660# 2.97e-19
C8516 a_11813_46116# a_13059_46348# 0.001208f
C8517 a_4883_46098# a_8049_45260# 0.469963f
C8518 a_14955_47212# a_13259_45724# 7.31e-21
C8519 a_11599_46634# a_14383_46116# 0.026426f
C8520 a_n743_46660# a_9823_46155# 0.196587f
C8521 a_2063_45854# a_1848_45724# 0.057473f
C8522 a_n1151_42308# a_n1099_45572# 0.046104f
C8523 a_12861_44030# a_16375_45002# 0.033138f
C8524 a_n881_46662# a_518_46482# 5.79e-19
C8525 a_2443_46660# a_3483_46348# 1.28e-19
C8526 a_2609_46660# a_3147_46376# 4.21e-19
C8527 a_15928_47570# a_6945_45028# 0.004753f
C8528 a_12549_44172# a_10809_44734# 2.27272f
C8529 a_13747_46662# a_17715_44484# 0.025502f
C8530 a_13661_43548# a_18189_46348# 2.95e-19
C8531 a_5807_45002# a_17957_46116# 0.00544f
C8532 a_4520_42826# a_5193_43172# 1.24e-19
C8533 a_20974_43370# a_19511_42282# 1.07e-21
C8534 a_21381_43940# a_13258_32519# 1.65e-19
C8535 a_8147_43396# a_8325_42308# 8.68e-22
C8536 a_12281_43396# a_1606_42308# 1.94e-20
C8537 a_16795_42852# a_17595_43084# 0.010079f
C8538 a_n97_42460# a_16197_42308# 3.2e-21
C8539 a_2982_43646# a_13575_42558# 1.36e-19
C8540 a_3626_43646# a_12563_42308# 0.005049f
C8541 a_3232_43370# a_5244_44056# 0.017099f
C8542 a_20841_45814# a_20935_43940# 6.15e-21
C8543 a_18479_45785# a_14021_43940# 0.025329f
C8544 a_10440_44484# a_8975_43940# 0.045841f
C8545 a_n1917_44484# a_n1821_44484# 0.013793f
C8546 a_n1699_44726# a_n1655_44484# 3.69e-19
C8547 a_n2129_44697# a_n23_44458# 2.23e-19
C8548 a_n2267_44484# a_n356_44636# 1.82e-20
C8549 a_5111_44636# a_5663_43940# 0.001818f
C8550 a_3537_45260# a_7845_44172# 0.001398f
C8551 a_n913_45002# a_n2661_42282# 0.054259f
C8552 a_5691_45260# a_5013_44260# 9.29e-19
C8553 a_n2661_44458# a_7_44811# 3.19e-19
C8554 a_n443_42852# a_7466_43396# 2.62e-19
C8555 a_21496_47436# a_3357_43084# 2.47e-20
C8556 a_13507_46334# a_22591_45572# 9.32e-20
C8557 a_n746_45260# a_1307_43914# 1.91e-20
C8558 a_4791_45118# a_7229_43940# 0.026326f
C8559 a_13059_46348# a_14949_46494# 6.26e-19
C8560 a_5164_46348# a_2324_44458# 5.59e-20
C8561 a_10355_46116# a_9290_44172# 0.01806f
C8562 a_n1641_46494# a_n1379_46482# 0.001705f
C8563 a_n1423_46090# a_n967_46494# 4.2e-19
C8564 a_9823_46155# a_11189_46129# 6.08e-20
C8565 a_n1151_42308# a_10951_45334# 1.15e-20
C8566 a_19692_46634# a_20850_46155# 0.006879f
C8567 a_12465_44636# a_2437_43646# 0.18195f
C8568 a_12861_44030# a_413_45260# 2.92e-19
C8569 a_6151_47436# a_3232_43370# 7.33e-19
C8570 a_13747_46662# a_15861_45028# 0.021551f
C8571 a_n1853_46287# a_n1533_46116# 8.49e-19
C8572 a_17701_42308# a_7174_31319# 2.14e-20
C8573 a_n961_42308# a_n3674_37592# 0.005438f
C8574 a_n4318_38680# a_n4334_38528# 0.08371f
C8575 a_4699_43561# VDD 0.262218f
C8576 a_n473_42460# a_n327_42558# 0.171361f
C8577 a_196_42282# a_n784_42308# 0.00268f
C8578 COMP_P a_n1630_35242# 2.45645f
C8579 a_n913_45002# a_16823_43084# 1.15e-20
C8580 a_14180_45002# a_14579_43548# 9.2e-22
C8581 a_14537_43396# a_13667_43396# 2.79e-19
C8582 a_4223_44672# a_3992_43940# 1.9e-19
C8583 a_3877_44458# VDD 0.786903f
C8584 a_n2661_43922# a_1241_44260# 3.45e-19
C8585 a_n2661_42834# a_1525_44260# 1.72e-19
C8586 a_9482_43914# a_15095_43370# 1.57e-19
C8587 a_13556_45296# a_14205_43396# 0.012255f
C8588 a_n2956_38216# a_n1736_42282# 2.12e-20
C8589 a_18287_44626# a_15493_43940# 1.79e-20
C8590 a_n2293_42834# a_n998_43396# 1.67e-19
C8591 a_5891_43370# a_10949_43914# 0.005033f
C8592 a_20193_45348# a_21381_43940# 0.01388f
C8593 a_n357_42282# a_20753_42852# 0.013117f
C8594 a_7499_43078# a_8483_43230# 8.28e-19
C8595 a_10809_44734# a_11525_45546# 2.29e-19
C8596 a_526_44458# a_4808_45572# 0.005047f
C8597 a_20205_31679# a_21167_46155# 4.36e-20
C8598 a_21363_46634# a_3357_43084# 2.28e-20
C8599 a_768_44030# a_8701_44490# 0.00464f
C8600 a_3090_45724# a_8953_45002# 8.01e-20
C8601 a_11415_45002# a_20273_45572# 0.01364f
C8602 a_20202_43084# a_20841_45814# 0.001988f
C8603 a_14180_46812# a_413_45260# 1.15e-20
C8604 a_6633_46155# a_2711_45572# 1.05e-19
C8605 a_5066_45546# a_6598_45938# 1.62e-19
C8606 a_21335_42336# a_21887_42336# 0.001613f
C8607 a_n1630_35242# a_n3565_37414# 6.25e-19
C8608 a_n2833_47464# SMPL_ON_P 0.002772f
C8609 a_n2497_47436# a_n1741_47186# 0.098118f
C8610 a_n2288_47178# a_n1920_47178# 7.52e-19
C8611 a_n3674_37592# a_n3420_37440# 0.073321f
C8612 a_13258_32519# a_21125_42558# 0.002663f
C8613 a_22400_42852# a_22459_39145# 0.242947f
C8614 a_n784_42308# a_n4064_37440# 0.014901f
C8615 a_5742_30871# a_n3565_38502# 4.45e-21
C8616 a_n2017_45002# a_3905_42558# 0.006025f
C8617 a_n913_45002# a_3497_42558# 0.004643f
C8618 a_5244_44056# a_4905_42826# 0.002354f
C8619 a_11827_44484# a_19987_42826# 2.96e-20
C8620 a_n2956_38216# a_n4209_37414# 4.59e-21
C8621 a_2479_44172# a_2982_43646# 0.019219f
C8622 a_13259_45724# a_22469_40625# 1.39e-19
C8623 a_9313_44734# a_21259_43561# 1.06e-19
C8624 a_5343_44458# a_8037_42858# 0.019942f
C8625 a_1414_42308# a_3539_42460# 5.28e-20
C8626 a_14955_43940# a_15037_43940# 0.171361f
C8627 a_n1736_46482# VDD 0.083417f
C8628 a_18184_42460# a_22223_42860# 0.03037f
C8629 a_19321_45002# a_20269_44172# 6.92e-19
C8630 a_12549_44172# a_12495_44260# 0.002899f
C8631 a_768_44030# a_11816_44260# 5.23e-19
C8632 a_19335_46494# a_16922_45042# 1.17e-20
C8633 a_n755_45592# a_n143_45144# 0.07862f
C8634 a_n863_45724# a_2382_45260# 0.119625f
C8635 a_n357_42282# a_n37_45144# 1.32e-21
C8636 a_3147_46376# a_2779_44458# 2.99e-20
C8637 a_12741_44636# a_18287_44626# 0.004901f
C8638 a_14035_46660# a_13857_44734# 9.44e-21
C8639 a_n2661_45546# a_4574_45260# 0.014727f
C8640 a_15227_44166# a_16241_44734# 0.105126f
C8641 a_n2293_46634# a_13483_43940# 8.18e-21
C8642 a_18479_47436# a_14401_32519# 3.18e-21
C8643 a_13925_46122# a_11827_44484# 5.41e-21
C8644 a_6419_46155# a_n2661_44458# 1.98e-22
C8645 a_n1099_45572# a_327_44734# 3.5e-20
C8646 a_310_45028# a_413_45260# 0.025313f
C8647 a_13163_45724# a_13297_45572# 0.001089f
C8648 a_11415_45002# a_18989_43940# 2.61e-19
C8649 a_1609_45822# a_n2661_45010# 0.003846f
C8650 a_10193_42453# a_18175_45572# 5.07e-21
C8651 a_n2293_45546# a_3065_45002# 9.28e-21
C8652 a_12005_46116# a_11691_44458# 8.12e-21
C8653 a_18189_46348# a_18587_45118# 5.47e-19
C8654 a_17957_46116# a_18315_45260# 3.37e-20
C8655 a_13259_45724# a_13159_45002# 0.047761f
C8656 a_n237_47217# a_10428_46928# 1.3e-19
C8657 a_6545_47178# a_4646_46812# 0.02302f
C8658 a_6491_46660# a_3877_44458# 0.02519f
C8659 a_12465_44636# a_n2661_46634# 1.89e-19
C8660 a_n3565_39590# VCM 0.097317f
C8661 a_n3420_38528# C1_P_btm 5.88e-20
C8662 a_n4064_39616# VIN_P 0.048523f
C8663 VDAC_Ni VDAC_P 1.02e-19
C8664 a_2063_45854# a_7411_46660# 0.029159f
C8665 a_4791_45118# a_5907_46634# 0.016954f
C8666 a_4915_47217# a_5385_46902# 9.3e-21
C8667 a_5129_47502# a_4817_46660# 0.001806f
C8668 a_n881_46662# a_12549_44172# 0.225257f
C8669 a_n1613_43370# a_768_44030# 0.028683f
C8670 a_n3420_39072# VDD 1.01442f
C8671 a_3754_38470# VDAC_N 0.169096f
C8672 a_n2109_47186# a_5841_46660# 1.94e-19
C8673 a_22959_47212# a_20916_46384# 9.45e-20
C8674 SMPL_ON_N a_22612_30879# 5.16049f
C8675 a_11453_44696# a_21588_30879# 0.075738f
C8676 a_n3565_37414# a_n3607_37440# 0.001003f
C8677 a_n2946_37690# a_n2860_37690# 0.011479f
C8678 a_7754_38470# a_5700_37509# 0.971846f
C8679 a_n4064_37440# a_n2302_37690# 0.239588f
C8680 a_8530_39574# a_5088_37509# 0.166912f
C8681 a_20974_43370# a_21259_43561# 0.049502f
C8682 a_n97_42460# a_16867_43762# 1.22e-19
C8683 a_14401_32519# a_4190_30871# 0.10855f
C8684 en_comp a_22780_40081# 4.3e-20
C8685 a_8147_43396# a_9145_43396# 1.64e-19
C8686 a_18175_45572# VDD 0.38478f
C8687 a_n356_44636# a_9223_42460# 1.4e-19
C8688 a_3483_46348# a_11341_43940# 0.017129f
C8689 a_10907_45822# a_n2661_44458# 3.96e-19
C8690 a_526_44458# a_1414_42308# 0.097596f
C8691 a_2324_44458# a_3499_42826# 1.36e-21
C8692 a_3090_45724# a_3626_43646# 4.54e-20
C8693 a_8270_45546# a_8791_43396# 6.22e-19
C8694 a_21588_30879# a_17364_32525# 0.05857f
C8695 a_8746_45002# a_10334_44484# 0.019787f
C8696 a_10180_45724# a_10057_43914# 0.002709f
C8697 a_n755_45592# a_n2293_43922# 4.58e-19
C8698 a_13259_45724# a_11967_42832# 0.141918f
C8699 a_4927_45028# a_5691_45260# 0.018415f
C8700 a_5111_44636# a_3232_43370# 0.134191f
C8701 a_5147_45002# a_6171_45002# 3.36e-19
C8702 a_9290_44172# a_10949_43914# 0.113864f
C8703 a_16327_47482# a_21195_42852# 5.9e-20
C8704 a_4791_45118# a_4649_42852# 3.78e-19
C8705 a_15599_45572# a_11827_44484# 4.86e-21
C8706 a_12465_44636# a_14543_43071# 2.17e-22
C8707 a_n1151_42308# a_n1925_42282# 3.65e-19
C8708 a_n443_46116# a_518_46482# 6.82e-19
C8709 a_3381_47502# a_526_44458# 9.83e-20
C8710 a_601_46902# a_765_45546# 1.65e-19
C8711 a_12861_44030# a_18985_46122# 4.61e-20
C8712 a_13717_47436# a_19553_46090# 3.99e-21
C8713 a_9863_47436# a_6945_45028# 0.0046f
C8714 a_5807_45002# a_11415_45002# 0.05094f
C8715 a_13661_43548# a_20202_43084# 1.29e-19
C8716 a_n881_46662# a_1208_46090# 0.076994f
C8717 a_n1613_43370# a_1176_45822# 0.004031f
C8718 a_4883_46098# a_8953_45546# 0.078639f
C8719 a_10227_46804# a_13351_46090# 0.008909f
C8720 a_11599_46634# a_17715_44484# 0.031427f
C8721 a_n237_47217# a_8283_46482# 1.91e-19
C8722 a_10150_46912# a_10384_47026# 0.006453f
C8723 a_6755_46942# a_6682_46660# 9.82e-21
C8724 a_10428_46928# a_8270_45546# 1.48e-19
C8725 a_3160_47472# a_3873_46454# 5.76e-19
C8726 a_15811_47375# a_15682_46116# 0.002105f
C8727 a_15673_47210# a_2324_44458# 1.57e-19
C8728 a_768_44030# a_n2293_46098# 0.039783f
C8729 a_9145_43396# a_13569_43230# 1.23e-19
C8730 a_19328_44172# a_19332_42282# 1.13e-21
C8731 a_4190_30871# a_18817_42826# 0.011301f
C8732 a_15493_43940# a_17124_42282# 1.54e-21
C8733 a_n1557_42282# a_n1329_42308# 0.075734f
C8734 a_13678_32519# a_5342_30871# 0.028488f
C8735 a_9165_43940# a_9223_42460# 4.51e-21
C8736 a_743_42282# a_17333_42852# 8.08e-20
C8737 a_1847_42826# a_2905_42968# 0.097535f
C8738 a_10440_44484# VDD 0.159539f
C8739 a_458_43396# a_1184_42692# 1.51e-20
C8740 a_n755_45592# a_n97_42460# 1.02989f
C8741 a_n357_42282# a_104_43370# 0.026213f
C8742 a_13507_46334# a_20712_42282# 4.89e-19
C8743 a_n2293_46098# a_5755_42852# 4.28e-20
C8744 SMPL_ON_P a_n2302_37984# 5.6e-20
C8745 a_1423_45028# a_8238_44734# 2.37e-19
C8746 a_11136_45572# a_10729_43914# 1.39e-20
C8747 a_n2293_46634# a_6123_31319# 4.66e-20
C8748 a_n1059_45260# a_18005_44484# 5.53e-20
C8749 a_11691_44458# a_20205_45028# 2.19e-19
C8750 a_20193_45348# a_19929_45028# 4.23e-19
C8751 a_22959_45036# a_19721_31679# 0.156264f
C8752 a_n2661_46634# a_2711_45572# 0.032616f
C8753 a_n2293_46634# a_1176_45572# 4.47e-19
C8754 a_20202_43084# a_4185_45028# 2.38e-19
C8755 a_11453_44696# a_10907_45822# 3.71e-19
C8756 a_10227_46804# a_15225_45822# 7.94e-20
C8757 a_11599_46634# a_15861_45028# 4.02e-19
C8758 a_33_46660# a_n443_42852# 1.61e-19
C8759 a_n743_46660# a_2307_45899# 2.73e-19
C8760 a_n2293_46098# a_1176_45822# 0.027035f
C8761 a_16327_47482# a_16333_45814# 0.168559f
C8762 a_n2661_46098# a_n755_45592# 7.65e-20
C8763 a_765_45546# a_12594_46348# 7.51e-20
C8764 a_n1641_46494# a_n1076_46494# 7.99e-20
C8765 a_11309_47204# a_7499_43078# 3.32e-22
C8766 a_n2293_42282# a_2725_42558# 1.65e-19
C8767 a_21487_43396# a_21613_42308# 9.66e-20
C8768 a_10083_42826# a_10723_42308# 0.001074f
C8769 a_10518_42984# a_10533_42308# 0.001423f
C8770 a_10341_42308# a_9803_42558# 0.108853f
C8771 a_13467_32519# a_21335_42336# 0.005979f
C8772 a_4361_42308# a_7174_31319# 0.024432f
C8773 a_5649_42852# a_13258_32519# 0.040931f
C8774 a_5342_30871# a_6123_31319# 0.018227f
C8775 a_5534_30871# a_5934_30871# 0.018227f
C8776 a_3080_42308# a_n4064_37440# 1.61e-19
C8777 a_18184_42460# a_20269_44172# 0.002397f
C8778 a_19778_44110# a_20365_43914# 1.6e-19
C8779 a_3065_45002# a_2896_43646# 6.3e-21
C8780 a_2382_45260# a_3540_43646# 0.006906f
C8781 a_n1613_43370# DATA[0] 0.001615f
C8782 a_11827_44484# a_18326_43940# 0.001776f
C8783 a_n2956_39304# a_n3674_37592# 0.026377f
C8784 a_18494_42460# a_19862_44208# 0.019692f
C8785 a_5111_44636# a_4905_42826# 0.128918f
C8786 a_n2661_43922# a_11967_42832# 1.74e-20
C8787 a_11691_44458# a_15682_43940# 0.013321f
C8788 a_n863_45724# a_1709_42852# 7.55e-19
C8789 a_n2017_45002# a_8791_43396# 2.77e-21
C8790 a_n1059_45260# a_8147_43396# 4.32e-21
C8791 a_5063_47570# DATA[3] 3.18e-20
C8792 a_8128_46384# VDD 0.403575f
C8793 a_5883_43914# a_7542_44172# 0.187537f
C8794 a_3232_43370# a_4235_43370# 6.06e-20
C8795 a_n743_46660# a_1423_45028# 4.79e-20
C8796 a_n2956_39304# a_n2840_45546# 4.31e-19
C8797 a_3877_44458# a_5691_45260# 4.47e-21
C8798 a_13059_46348# a_16680_45572# 1.67e-21
C8799 a_16388_46812# a_16855_45546# 4.77e-21
C8800 a_15227_44166# a_18691_45572# 5.63e-21
C8801 a_n133_46660# a_626_44172# 1.1e-21
C8802 a_5204_45822# a_6511_45714# 2.92e-21
C8803 a_6419_46155# a_5907_45546# 2.91e-20
C8804 a_6165_46155# a_6194_45824# 5.54e-19
C8805 a_5807_45002# a_6945_45348# 2.54e-21
C8806 a_5167_46660# a_3537_45260# 9.28e-22
C8807 a_12741_44636# a_13904_45546# 2.6e-21
C8808 a_11415_45002# a_15143_45578# 0.003102f
C8809 a_3090_45724# a_17568_45572# 4.36e-20
C8810 a_2324_44458# a_3316_45546# 1.07e-19
C8811 a_33_46660# a_375_42282# 2.38e-20
C8812 a_8199_44636# a_2711_45572# 0.098064f
C8813 a_4419_46090# a_3775_45552# 2.91e-21
C8814 a_4651_46660# a_5111_44636# 7.15e-21
C8815 a_4883_46098# a_20193_45348# 3.03e-20
C8816 a_19692_46634# a_18479_45785# 5.23e-20
C8817 a_19466_46812# a_18341_45572# 0.02497f
C8818 a_765_45546# a_15037_45618# 3e-21
C8819 a_n3674_37592# a_n3565_39304# 6.52e-20
C8820 a_15486_42560# a_15803_42450# 0.102355f
C8821 a_14113_42308# a_15890_42674# 0.022182f
C8822 a_6761_42308# a_7174_31319# 4.88e-21
C8823 a_n3674_38680# a_n4209_38502# 0.04481f
C8824 a_5534_30871# a_11530_34132# 0.010307f
C8825 a_n1630_35242# a_n4209_39304# 4.66e-19
C8826 a_n784_42308# a_n3420_39072# 0.003982f
C8827 a_1847_42826# VDD 0.527555f
C8828 a_5342_30871# EN_VIN_BSTR_P 0.010795f
C8829 a_2479_44172# a_2253_43940# 0.010537f
C8830 a_2127_44172# a_2455_43940# 0.096132f
C8831 a_895_43940# a_1443_43940# 0.016028f
C8832 a_22959_46660# EN_OFFSET_CAL 0.050989f
C8833 a_n1641_46494# VDD 0.226065f
C8834 a_10729_43914# a_11750_44172# 0.144893f
C8835 a_10949_43914# a_10807_43548# 0.034945f
C8836 a_20193_45348# a_5649_42852# 0.052027f
C8837 a_11823_42460# a_13070_42354# 0.077142f
C8838 a_3537_45260# a_4149_42891# 2.78e-19
C8839 a_18374_44850# a_10341_43396# 3.04e-21
C8840 a_10193_42453# a_15486_42560# 8.28e-20
C8841 a_2711_45572# a_19511_42282# 0.234026f
C8842 a_n913_45002# a_11136_42852# 0.026537f
C8843 a_n2293_42834# a_9127_43156# 4.88e-19
C8844 a_6598_45938# a_6977_45572# 3.16e-19
C8845 a_526_44458# a_1667_45002# 2.21e-19
C8846 a_21588_30879# a_19237_31679# 0.055917f
C8847 a_11415_45002# a_18315_45260# 0.00724f
C8848 a_12741_44636# a_17023_45118# 0.005061f
C8849 a_19443_46116# a_19256_45572# 2.91e-19
C8850 a_16327_47482# a_15493_43396# 0.025969f
C8851 a_12861_44030# a_22223_43948# 0.001164f
C8852 a_14275_46494# a_14797_45144# 1.37e-19
C8853 a_15015_46420# a_14537_43396# 1.61e-20
C8854 a_6945_45028# a_7229_43940# 0.001224f
C8855 a_2711_45572# a_8192_45572# 0.005217f
C8856 a_10053_45546# a_10193_42453# 0.086012f
C8857 a_4185_45028# a_5837_45028# 1.38e-19
C8858 a_3090_45724# a_17767_44458# 1.66e-19
C8859 a_768_44030# a_2675_43914# 0.026212f
C8860 a_2324_44458# a_13777_45326# 0.002856f
C8861 a_7499_43078# a_10490_45724# 4.9e-20
C8862 a_5257_43370# a_n2661_43922# 0.030003f
C8863 a_9049_44484# a_8746_45002# 0.025877f
C8864 a_4883_46098# a_9028_43914# 0.002203f
C8865 a_n1613_43370# a_7845_44172# 5.96e-21
C8866 a_20894_47436# a_20990_47178# 0.313533f
C8867 a_15486_42560# VDD 0.275297f
C8868 a_15051_42282# RST_Z 0.001018f
C8869 a_n2109_47186# a_n1925_46634# 0.033276f
C8870 a_18143_47464# a_12465_44636# 0.001005f
C8871 a_19386_47436# a_13507_46334# 6.44e-21
C8872 a_18780_47178# a_4883_46098# 4.43e-20
C8873 a_18479_47436# a_21811_47423# 1.31e-19
C8874 a_2112_39137# a_3754_38470# 2.65e-20
C8875 a_22465_38105# CAL_P 0.026947f
C8876 SMPL_ON_P a_n2293_46634# 9.68e-20
C8877 a_n452_47436# a_n2661_46634# 0.001956f
C8878 a_n1605_47204# a_n2442_46660# 3.01e-19
C8879 a_4915_47217# a_12891_46348# 0.156543f
C8880 a_4791_45118# a_768_44030# 0.03019f
C8881 a_6491_46660# a_8128_46384# 6.19e-21
C8882 a_6575_47204# a_n881_46662# 0.708623f
C8883 a_7903_47542# a_7989_47542# 0.006584f
C8884 a_n2497_47436# a_n743_46660# 1.09e-19
C8885 a_7174_31319# a_n1532_35090# 1.2e-19
C8886 a_4958_30871# C4_P_btm 1.18e-19
C8887 a_13483_43940# a_743_42282# 4.27e-21
C8888 a_9313_44734# a_13291_42460# 0.003344f
C8889 a_3905_42865# a_3681_42891# 0.101054f
C8890 a_2998_44172# a_4520_42826# 5.74e-20
C8891 a_15037_43940# a_8685_43396# 6.84e-19
C8892 a_20679_44626# a_21671_42860# 3.31e-21
C8893 a_3422_30871# a_17595_43084# 6.38e-21
C8894 a_18579_44172# a_19339_43156# 3.57e-20
C8895 a_15493_43940# a_19268_43646# 9.38e-20
C8896 a_n97_42460# a_548_43396# 9.03e-19
C8897 a_4235_43370# a_4905_42826# 8.27e-21
C8898 a_1756_43548# a_n1557_42282# 1.14e-20
C8899 a_1568_43370# a_1427_43646# 0.046825f
C8900 a_4699_43561# a_3080_42308# 0.223965f
C8901 a_10053_45546# VDD 0.150582f
C8902 a_4646_46812# a_4699_43561# 2.54e-20
C8903 a_n2661_45546# a_5883_43914# 3.15e-21
C8904 a_1138_42852# a_895_43940# 0.017458f
C8905 a_2063_45854# a_10835_43094# 8.1e-21
C8906 a_n2293_46634# a_6809_43396# 3.99e-19
C8907 a_15227_44166# a_15037_44260# 6.14e-19
C8908 a_11453_44696# a_16823_43084# 7.31e-22
C8909 a_11322_45546# a_n2661_43370# 0.01285f
C8910 a_16333_45814# a_14537_43396# 4.99e-21
C8911 a_18189_46348# a_11967_42832# 2.07e-20
C8912 a_19963_31679# a_20447_31679# 0.069779f
C8913 a_13661_43548# a_14955_43396# 3.87e-20
C8914 a_n357_42282# a_949_44458# 0.016511f
C8915 a_n755_45592# a_742_44458# 3e-20
C8916 a_15599_45572# a_15595_45028# 2.01e-19
C8917 a_8696_44636# a_9482_43914# 0.042504f
C8918 a_1823_45246# a_2479_44172# 7.38e-19
C8919 a_19692_46634# a_14021_43940# 0.775991f
C8920 a_17339_46660# a_17973_43940# 8.68e-20
C8921 a_13717_47436# a_12741_44636# 5.57e-20
C8922 C2_P_btm VREF 0.987884f
C8923 a_21177_47436# a_20107_46660# 9.39e-19
C8924 a_20894_47436# a_20273_46660# 6.02e-20
C8925 a_13507_46334# a_19551_46910# 0.002438f
C8926 a_10227_46804# a_20731_47026# 0.016434f
C8927 C3_P_btm VREF_GND 0.67174f
C8928 C4_P_btm VCM 0.716447f
C8929 a_3877_44458# a_4646_46812# 0.056449f
C8930 a_n971_45724# a_8349_46414# 0.01782f
C8931 a_n1741_47186# a_9569_46155# 4.67e-20
C8932 a_n237_47217# a_7920_46348# 0.059304f
C8933 a_n443_46116# a_1208_46090# 1.26e-19
C8934 a_3524_46660# a_5072_46660# 5.75e-21
C8935 a_n1925_46634# a_5841_46660# 1.6e-19
C8936 a_2063_45854# a_4185_45028# 0.023928f
C8937 a_n1151_42308# a_2698_46116# 9.22e-21
C8938 a_2905_45572# a_3147_46376# 0.02017f
C8939 a_584_46384# a_4419_46090# 3.79e-21
C8940 a_3160_47472# a_2804_46116# 4.58e-19
C8941 a_12549_44172# a_17609_46634# 0.487224f
C8942 C0_P_btm VIN_P 0.529671f
C8943 a_n2661_46634# a_8654_47026# 1.14e-19
C8944 a_5807_45002# a_12251_46660# 0.003883f
C8945 a_4007_47204# a_1823_45246# 4.86e-22
C8946 a_4883_46098# a_18285_46348# 0.026239f
C8947 C10_N_btm VDD 2.40001f
C8948 a_12465_44636# a_765_45546# 0.019565f
C8949 a_3422_30871# a_21887_42336# 0.003456f
C8950 a_21487_43396# a_4361_42308# 0.077645f
C8951 a_8333_44056# a_5934_30871# 2.88e-21
C8952 a_8685_43396# a_15279_43071# 0.011343f
C8953 a_10341_43396# a_10083_42826# 0.002266f
C8954 a_5205_44484# a_5883_43914# 0.003713f
C8955 a_n443_42852# a_15682_43940# 0.002992f
C8956 a_2324_44458# a_6197_43396# 0.001135f
C8957 a_3483_46348# a_10341_43396# 2.31e-19
C8958 a_20692_30879# a_14021_43940# 1.18e-20
C8959 a_6709_45028# a_6298_44484# 0.006607f
C8960 a_5111_44636# a_8975_43940# 5.4e-19
C8961 a_12741_44636# a_19268_43646# 3.85e-21
C8962 a_3090_45724# a_8037_42858# 1.28e-20
C8963 a_n357_42282# a_11341_43940# 1.86e-19
C8964 a_4185_45028# a_14955_43396# 3.39e-21
C8965 a_8191_45002# a_5343_44458# 1.33e-19
C8966 a_6171_45002# a_10157_44484# 4.27e-20
C8967 a_3232_43370# a_10334_44484# 0.040395f
C8968 a_8953_45546# a_8685_43396# 0.062741f
C8969 a_n881_46662# a_n2661_45546# 0.02866f
C8970 a_n310_47243# a_n755_45592# 3.51e-20
C8971 a_2959_46660# a_526_44458# 6.06e-19
C8972 a_n1151_42308# a_13527_45546# 1.73e-20
C8973 a_20411_46873# a_20273_46660# 0.219954f
C8974 a_20107_46660# a_20841_46902# 0.053479f
C8975 a_n743_46660# a_9823_46482# 0.004996f
C8976 a_12549_44172# a_19443_46116# 3.9e-22
C8977 a_8270_45546# a_7920_46348# 5.66e-19
C8978 a_6151_47436# a_10193_42453# 5.26e-20
C8979 a_10249_46116# a_10903_43370# 7.46e-21
C8980 a_5807_45002# a_13259_45724# 0.096565f
C8981 a_3090_45724# a_167_45260# 5.35e-19
C8982 a_14035_46660# a_12741_44636# 8.27e-21
C8983 a_n1925_46634# a_8062_46155# 1.86e-19
C8984 a_5342_30871# a_15597_42852# 0.003587f
C8985 a_15781_43660# a_15890_42674# 2.11e-20
C8986 a_5244_44056# VDD 0.146618f
C8987 a_16547_43609# a_14113_42308# 6.85e-19
C8988 a_1847_42826# a_n784_42308# 0.001475f
C8989 a_4190_30871# a_5934_30871# 0.020923f
C8990 a_4361_42308# a_5932_42308# 0.072603f
C8991 a_743_42282# a_6123_31319# 0.018532f
C8992 a_6151_47436# VDD 4.39915f
C8993 a_14537_43396# a_15493_43396# 5.06e-19
C8994 a_4007_47204# DATA[2] 0.337596f
C8995 a_n2012_44484# a_n2661_42834# 0.001285f
C8996 a_n755_45592# a_n901_43156# 1.1e-19
C8997 a_n357_42282# a_n1076_43230# 0.001306f
C8998 a_12607_44458# a_12553_44484# 6.75e-20
C8999 a_7640_43914# a_5891_43370# 0.011186f
C9000 a_21359_45002# a_19237_31679# 8.84e-20
C9001 a_15227_44166# a_15890_42674# 0.001386f
C9002 a_11963_45334# a_11341_43940# 1.74e-20
C9003 a_11387_46155# a_8049_45260# 0.00421f
C9004 a_n2157_46122# a_n2661_45546# 5.14e-20
C9005 a_n2293_46098# a_n2472_45546# 0.015672f
C9006 a_11453_44696# a_15415_45028# 0.005374f
C9007 a_8199_44636# a_10037_46155# 4.91e-19
C9008 a_n2472_46090# a_n2956_38216# 5.66e-19
C9009 a_765_45546# a_2711_45572# 5.89e-20
C9010 a_14976_45028# a_11823_42460# 0.010375f
C9011 a_n881_46662# a_5205_44484# 0.013688f
C9012 a_2324_44458# a_5066_45546# 0.002463f
C9013 a_n1736_46482# a_n1545_46494# 4.61e-19
C9014 a_17364_32525# a_22469_39537# 1.61e-20
C9015 a_4190_30871# a_11530_34132# 0.031248f
C9016 a_1755_42282# a_5742_30871# 3.99e-20
C9017 a_1606_42308# a_11551_42558# 1.77e-20
C9018 a_14097_32519# a_4958_30871# 0.030871f
C9019 a_22400_42852# a_17303_42282# 0.004332f
C9020 a_5534_30871# a_7754_40130# 0.002632f
C9021 a_5755_42308# a_6123_31319# 2.22e-20
C9022 a_5932_42308# a_6761_42308# 0.001757f
C9023 a_15227_44166# START 0.001035f
C9024 a_175_44278# a_261_44278# 0.006584f
C9025 a_n984_44318# a_n822_43940# 0.006453f
C9026 a_19333_46634# RST_Z 1.4e-20
C9027 a_3537_45260# a_5111_42852# 0.123919f
C9028 a_n443_42852# a_5934_30871# 1.89e-19
C9029 a_n913_45002# a_12545_42858# 0.548984f
C9030 a_n1059_45260# a_13113_42826# 0.002702f
C9031 a_n2017_45002# a_12895_43230# 1.47e-19
C9032 a_n2956_39304# a_n2302_39072# 0.040755f
C9033 a_n2956_38680# a_n4064_39072# 0.001709f
C9034 a_20362_44736# a_20269_44172# 2.05e-20
C9035 a_20159_44458# a_20365_43914# 0.003347f
C9036 a_5244_44056# a_5495_43940# 0.107037f
C9037 a_18579_44172# a_17973_43940# 5.34e-19
C9038 a_13607_46688# CLK 2.1e-20
C9039 a_n357_42282# a_10723_42308# 7.12e-20
C9040 a_11967_42832# a_20935_43940# 9.08e-20
C9041 a_20640_44752# a_19862_44208# 0.001675f
C9042 a_19466_46812# VDD 0.664497f
C9043 a_18374_44850# a_n97_42460# 1.3e-21
C9044 a_21076_30879# VDAC_N 0.001403f
C9045 a_19279_43940# a_18451_43940# 3.9e-19
C9046 a_18597_46090# a_21073_44484# 6.09e-19
C9047 a_n755_45592# a_3733_45822# 4.98e-19
C9048 a_13259_45724# a_15143_45578# 0.060775f
C9049 a_n1925_46634# a_8375_44464# 1.53e-21
C9050 a_10809_44734# a_19431_45546# 5.65e-21
C9051 a_1823_45246# a_2680_45002# 0.073588f
C9052 a_14976_45028# a_16321_45348# 2.16e-20
C9053 a_11133_46155# a_3357_43084# 1.78e-21
C9054 a_18479_47436# a_20512_43084# 1.2e-19
C9055 a_10586_45546# a_10216_45572# 1.7e-19
C9056 a_5807_45002# a_n2661_43922# 1.32e-19
C9057 a_11415_45002# a_13017_45260# 0.100288f
C9058 a_768_44030# a_10809_44484# 1.65e-19
C9059 a_167_45260# a_2274_45254# 8.13e-20
C9060 a_n1151_42308# a_n875_44318# 5.38e-21
C9061 a_n3565_39590# a_n4064_38528# 0.031177f
C9062 a_n4315_30879# a_n4209_38216# 0.053149f
C9063 a_1343_38525# a_1239_39043# 0.01446f
C9064 a_n4334_39392# a_n4251_39392# 0.007692f
C9065 a_n4209_39304# a_n3607_39392# 0.002352f
C9066 a_1606_42308# C0_dummy_N_btm 0.007541f
C9067 a_n784_42308# C10_N_btm 1.34e-19
C9068 a_14097_32519# VCM 0.00888f
C9069 a_n4064_40160# a_n4251_38528# 0.001069f
C9070 a_n473_42460# VDD 0.27195f
C9071 a_n3420_39616# a_n3420_38528# 0.049464f
C9072 a_n4064_39616# a_n3565_38502# 0.02802f
C9073 a_n3565_39304# a_n2302_39072# 0.066757f
C9074 a_n3690_39392# a_n4064_39072# 0.085872f
C9075 a_n3420_39072# a_n2946_39072# 0.238708f
C9076 a_n443_46116# a_6575_47204# 2.21e-20
C9077 a_4915_47217# a_7903_47542# 0.042037f
C9078 a_6151_47436# a_6491_46660# 0.31912f
C9079 a_5815_47464# a_6851_47204# 1.23e-20
C9080 a_n1151_42308# a_n1435_47204# 0.002911f
C9081 a_5932_42308# a_n1532_35090# 1.05e-19
C9082 a_5742_30871# VDAC_P 0.030337f
C9083 a_20512_43084# a_4190_30871# 0.006642f
C9084 a_1241_43940# a_1209_43370# 3.49e-19
C9085 a_n1059_45260# a_18214_42558# 0.020063f
C9086 a_n913_45002# a_19332_42282# 2.77e-19
C9087 a_n2293_43922# a_10083_42826# 2.45e-20
C9088 a_375_42282# a_5934_30871# 1.48e-20
C9089 a_n2293_42834# a_1755_42282# 1.34e-19
C9090 a_9028_43914# a_8685_43396# 1.97e-20
C9091 en_comp a_17531_42308# 1.87e-20
C9092 a_20205_31679# VDD 0.737305f
C9093 a_9313_44734# a_13460_43230# 0.004332f
C9094 a_3422_30871# a_13467_32519# 0.421402f
C9095 w_11334_34010# a_13678_32519# 3.98e-19
C9096 a_2107_46812# a_9801_43940# 3.07e-19
C9097 a_17957_46116# a_18374_44850# 8.91e-21
C9098 a_7230_45938# a_7276_45260# 4.28e-19
C9099 a_12741_44636# a_17061_44484# 1.5e-19
C9100 a_18175_45572# a_18479_45785# 0.280208f
C9101 a_16147_45260# a_18341_45572# 0.001545f
C9102 a_10809_44734# a_13076_44458# 1.02e-19
C9103 a_768_44030# a_1209_43370# 1.23e-20
C9104 a_20202_43084# a_11967_42832# 0.02752f
C9105 a_7499_43078# a_6171_45002# 0.029896f
C9106 a_9049_44484# a_3232_43370# 0.17048f
C9107 a_4185_45028# a_n2661_42834# 0.023267f
C9108 a_13259_45724# a_18315_45260# 0.144632f
C9109 a_16375_45002# a_17023_45118# 0.014031f
C9110 a_n1925_42282# a_4223_44672# 0.053508f
C9111 a_526_44458# a_n699_43396# 0.285f
C9112 a_n2946_37690# VDD 0.38221f
C9113 a_4883_46098# a_10249_46116# 0.01923f
C9114 a_n2312_38680# a_n1021_46688# 7.19e-20
C9115 a_n2293_46634# a_n2438_43548# 0.807205f
C9116 a_n2104_46634# a_n743_46660# 6.41e-20
C9117 VDAC_P C0_dummy_P_btm 0.284358f
C9118 a_n881_46662# a_5385_46902# 5.4e-19
C9119 a_12861_44030# a_12816_46660# 7.2e-19
C9120 a_13717_47436# a_13607_46688# 6.92e-19
C9121 a_n1613_43370# a_5167_46660# 0.177362f
C9122 CAL_P a_18194_35068# 0.010626f
C9123 a_n1838_35608# a_n1386_35608# 0.150796f
C9124 VDAC_N C0_N_btm 0.324278f
C9125 a_11599_46634# a_11901_46660# 0.002693f
C9126 a_n2661_46634# a_33_46660# 0.050833f
C9127 a_4915_47217# a_12359_47026# 2.51e-19
C9128 a_n1151_42308# a_13885_46660# 0.333314f
C9129 a_8128_46384# a_4646_46812# 5.76e-21
C9130 a_14955_43396# a_15037_43396# 0.005781f
C9131 a_15095_43370# a_15125_43396# 0.007578f
C9132 a_n97_42460# a_10083_42826# 6.2e-20
C9133 a_413_45260# CLK 0.033653f
C9134 a_14673_44172# a_14113_42308# 2.36e-21
C9135 a_3080_42308# a_1847_42826# 2.31e-19
C9136 a_n1557_42282# a_421_43172# 3.1e-19
C9137 a_n4318_39768# a_n3674_38216# 0.023361f
C9138 a_5111_44636# VDD 1.28013f
C9139 a_15781_43660# a_16547_43609# 5.24e-19
C9140 a_10341_43396# a_16664_43396# 0.005311f
C9141 a_15681_43442# a_16409_43396# 3.1e-20
C9142 a_1467_44172# a_1606_42308# 2.54e-20
C9143 a_5891_43370# a_7174_31319# 9.47e-21
C9144 a_2232_45348# a_2304_45348# 0.003395f
C9145 a_11525_45546# a_11541_44484# 2.97e-20
C9146 a_6431_45366# a_n2661_43370# 0.009143f
C9147 a_n755_45592# a_n984_44318# 0.002789f
C9148 a_n357_42282# a_175_44278# 0.002018f
C9149 a_6171_45002# a_11915_45394# 7.98e-19
C9150 en_comp a_18184_42460# 2.88e-20
C9151 a_n2017_45002# a_11827_44484# 2.08e-20
C9152 a_15227_44166# a_16547_43609# 1.88e-20
C9153 w_11334_34010# a_6123_31319# 6.03e-19
C9154 a_3483_46348# a_n97_42460# 1.02e-19
C9155 a_7229_43940# a_7735_45067# 0.005614f
C9156 a_8191_45002# a_8560_45348# 0.03364f
C9157 a_6709_45028# a_7418_45067# 0.001659f
C9158 a_13249_42308# a_13213_44734# 1.19e-20
C9159 a_n863_45724# a_453_43940# 0.02533f
C9160 a_16327_47482# a_18707_42852# 0.012993f
C9161 a_21513_45002# a_18114_32519# 9.32e-20
C9162 a_10306_45572# a_5891_43370# 2.85e-21
C9163 a_13059_46348# a_14358_43442# 0.041731f
C9164 a_2107_46812# a_6165_46155# 0.003422f
C9165 a_2553_47502# a_n755_45592# 8.3e-22
C9166 a_n443_46116# a_n2661_45546# 0.136593f
C9167 a_14084_46812# a_13885_46660# 0.237373f
C9168 a_13607_46688# a_14035_46660# 0.003044f
C9169 a_12816_46660# a_14180_46812# 5.52e-19
C9170 a_4883_46098# a_8781_46436# 7.71e-20
C9171 a_n2661_46634# a_12005_46116# 0.038027f
C9172 a_584_46384# a_1848_45724# 3.13e-19
C9173 a_n971_45724# a_n906_45572# 0.001365f
C9174 a_1057_46660# a_1176_45822# 1.55e-19
C9175 a_2443_46660# a_3147_46376# 5.77e-19
C9176 a_n743_46660# a_9569_46155# 0.104962f
C9177 a_768_44030# a_6945_45028# 0.014703f
C9178 a_12891_46348# a_10809_44734# 0.102888f
C9179 a_13661_43548# a_17715_44484# 0.003425f
C9180 a_13747_46662# a_17583_46090# 1.47e-19
C9181 a_5807_45002# a_18189_46348# 0.033239f
C9182 a_14311_47204# a_13259_45724# 4.93e-21
C9183 a_4520_42826# a_4743_43172# 0.011458f
C9184 a_2982_43646# a_13070_42354# 7.37e-20
C9185 a_19237_31679# a_22469_39537# 2.75e-20
C9186 a_10903_43370# a_5534_30871# 0.134296f
C9187 a_n443_42852# a_7221_43396# 1.62e-19
C9188 a_n2433_44484# a_n23_44458# 2.38e-21
C9189 a_3232_43370# a_3905_42865# 0.027169f
C9190 a_10440_44484# a_10057_43914# 0.026774f
C9191 a_10334_44484# a_8975_43940# 0.044798f
C9192 a_n2129_44697# a_n356_44636# 0.009952f
C9193 a_n1699_44726# a_n1821_44484# 3.16e-19
C9194 a_5111_44636# a_5495_43940# 0.037006f
C9195 a_5147_45002# a_5663_43940# 0.019985f
C9196 a_3537_45260# a_7542_44172# 1.57e-19
C9197 a_n1059_45260# a_n2661_42282# 0.028862f
C9198 a_21188_45572# a_19862_44208# 1.49e-19
C9199 a_n2661_44458# a_n310_44811# 3.72e-19
C9200 a_n357_42282# a_10341_43396# 9.55e-19
C9201 a_13507_46334# a_3357_43084# 0.050295f
C9202 a_21811_47423# a_2437_43646# 0.025192f
C9203 a_18597_46090# a_21542_45572# 4.51e-19
C9204 a_n971_45724# a_1307_43914# 0.019541f
C9205 a_n2157_46122# a_n1533_46116# 9.73e-19
C9206 a_n1151_42308# a_10775_45002# 7.13e-22
C9207 a_4791_45118# a_7276_45260# 0.004255f
C9208 a_13059_46348# a_14537_46482# 0.002353f
C9209 a_n1641_46494# a_n1545_46494# 0.013793f
C9210 a_n1423_46090# a_n1379_46482# 3.69e-19
C9211 a_10623_46897# a_2711_45572# 8.62e-20
C9212 a_19692_46634# a_20692_30879# 4.77e-20
C9213 a_13717_47436# a_413_45260# 4.36729f
C9214 a_768_44030# a_14127_45572# 0.002434f
C9215 a_21363_46634# a_8049_45260# 3.11e-20
C9216 a_13661_43548# a_15861_45028# 0.047089f
C9217 a_5807_45002# a_17478_45572# 1.08e-20
C9218 a_13747_46662# a_8696_44636# 0.02273f
C9219 a_9625_46129# a_11133_46155# 4.63e-20
C9220 a_n1991_46122# a_n967_46494# 2.36e-20
C9221 a_17595_43084# a_7174_31319# 2.85e-21
C9222 a_22223_42860# a_17303_42282# 4.73e-19
C9223 a_n1329_42308# a_n3674_37592# 0.005224f
C9224 a_3080_42308# C10_N_btm 1.34e-19
C9225 a_4235_43370# VDD 0.229422f
C9226 a_n4318_37592# a_n1630_35242# 0.847279f
C9227 a_n473_42460# a_n784_42308# 0.020033f
C9228 a_4190_30871# a_7754_40130# 4.95e-20
C9229 a_n3674_39304# a_n4334_38528# 6.7e-20
C9230 a_n4318_38680# a_n4209_38502# 0.105064f
C9231 a_n1059_45260# a_16823_43084# 0.318918f
C9232 a_19963_31679# a_13467_32519# 0.051345f
C9233 a_4223_44672# a_3737_43940# 1.52e-19
C9234 a_11827_44484# a_21845_43940# 1.08e-19
C9235 a_n2661_42834# a_1241_44260# 3.84e-19
C9236 a_19279_43940# a_19237_31679# 5.63e-21
C9237 a_3422_30871# a_22315_44484# 0.19914f
C9238 a_19479_31679# a_13678_32519# 0.051236f
C9239 a_n1925_42282# a_5742_30871# 5.06e-20
C9240 a_9482_43914# a_14205_43396# 1.91e-22
C9241 a_n2956_38216# a_n3674_38216# 0.028821f
C9242 a_18248_44752# a_15493_43940# 8.91e-20
C9243 a_18443_44721# a_11341_43940# 2.01e-20
C9244 a_9290_44172# a_7174_31319# 2.43e-20
C9245 a_n2293_42834# a_n1243_43396# 1.39e-19
C9246 a_5891_43370# a_10729_43914# 0.001943f
C9247 a_n2810_45572# COMP_P 2.2e-21
C9248 a_n357_42282# a_20356_42852# 0.001192f
C9249 a_7499_43078# a_8292_43218# 7.98e-20
C9250 a_10809_44734# a_11322_45546# 0.22629f
C9251 a_526_44458# a_5024_45822# 1.2e-19
C9252 a_5257_43370# a_5837_45028# 0.008516f
C9253 a_12861_44030# a_13213_44734# 0.002516f
C9254 a_20623_46660# a_3357_43084# 0.013905f
C9255 a_10227_46804# a_9313_44734# 0.875947f
C9256 a_3090_45724# a_8191_45002# 7.02e-22
C9257 a_11415_45002# a_20107_45572# 0.019157f
C9258 a_20202_43084# a_20273_45572# 0.003019f
C9259 a_22000_46634# a_2437_43646# 0.010034f
C9260 a_14035_46660# a_413_45260# 2.37e-20
C9261 a_15227_44166# a_6171_45002# 0.021072f
C9262 a_20205_31679# a_20850_46155# 4.73e-21
C9263 a_768_44030# a_8103_44636# 0.004654f
C9264 a_4817_46660# a_n2661_43370# 6.7e-21
C9265 a_6347_46155# a_2711_45572# 1.62e-19
C9266 a_6945_45028# a_11652_45724# 2.08e-20
C9267 a_5066_45546# a_6667_45809# 1.76e-19
C9268 a_5934_30871# a_n3420_37984# 2.14e-19
C9269 a_n2288_47178# a_n2109_47186# 0.177673f
C9270 a_n2497_47436# a_n1920_47178# 0.049461f
C9271 a_n2833_47464# a_n1741_47186# 3.87e-20
C9272 a_6123_31319# a_n4064_37984# 1.56e-19
C9273 a_n3674_37592# a_n3690_37440# 0.071822f
C9274 a_19511_42282# a_21421_42336# 8.32e-19
C9275 a_22400_42852# a_22521_40055# 0.681186f
C9276 a_4223_44672# a_8387_43230# 4.84e-21
C9277 a_11691_44458# a_18249_42858# 5.39e-21
C9278 a_11967_42832# a_14955_43396# 2.03e-19
C9279 a_n913_45002# a_5379_42460# 0.179494f
C9280 a_n2017_45002# a_3581_42558# 0.001947f
C9281 a_n2810_45572# a_n3565_37414# 1.88e-20
C9282 a_3905_42865# a_4905_42826# 0.404829f
C9283 a_6298_44484# a_7227_42852# 2.52e-20
C9284 a_10809_44734# SINGLE_ENDED 0.008311f
C9285 a_11827_44484# a_19164_43230# 1.08e-21
C9286 a_5111_44636# a_n784_42308# 2.01e-20
C9287 a_2479_44172# a_2896_43646# 0.026857f
C9288 a_13259_45724# a_22521_40599# 3.75e-19
C9289 a_5343_44458# a_7765_42852# 0.010279f
C9290 a_1414_42308# a_3626_43646# 0.015112f
C9291 a_n2956_38680# VDD 0.871805f
C9292 a_18184_42460# a_22165_42308# 0.026631f
C9293 a_13829_44260# a_14021_43940# 1.97e-19
C9294 a_18597_46090# a_21205_44306# 6.68e-19
C9295 a_13747_46662# a_20365_43914# 1.31e-20
C9296 a_768_44030# a_11173_44260# 0.005635f
C9297 a_n755_45592# a_n467_45028# 0.26002f
C9298 a_n863_45724# a_2274_45254# 0.17549f
C9299 a_2804_46116# a_2779_44458# 9.85e-20
C9300 a_12741_44636# a_18248_44752# 0.00762f
C9301 a_n2661_45546# a_3537_45260# 0.780422f
C9302 a_15227_44166# a_14673_44172# 0.357896f
C9303 a_n2293_46634# a_12429_44172# 9.2e-20
C9304 a_18479_47436# a_21381_43940# 8.4e-20
C9305 a_19321_45002# a_19862_44208# 0.090113f
C9306 a_13759_46122# a_11827_44484# 4.47e-21
C9307 a_6165_46155# a_n2661_44458# 1.3e-22
C9308 a_1823_45246# a_5518_44484# 4.84e-19
C9309 a_n1099_45572# a_413_45260# 0.008675f
C9310 a_380_45546# a_327_44734# 6.27e-19
C9311 a_310_45028# a_n37_45144# 0.112458f
C9312 a_11415_45002# a_18374_44850# 6.96e-20
C9313 a_n443_42852# a_n2661_45010# 0.001666f
C9314 a_n971_45724# a_9396_43370# 2.62e-20
C9315 a_17339_46660# a_9313_44734# 2.43e-19
C9316 a_10193_42453# a_16147_45260# 0.193225f
C9317 a_584_46384# a_1512_43396# 7.9e-20
C9318 a_n443_46116# a_1427_43646# 0.05874f
C9319 a_n2293_45546# a_2680_45002# 3.47e-20
C9320 a_11823_42460# a_13385_45572# 1.28e-19
C9321 a_10903_43370# a_11691_44458# 0.020718f
C9322 a_n1925_42282# a_n2293_42834# 0.024873f
C9323 a_18189_46348# a_18315_45260# 0.101775f
C9324 a_17957_46116# a_17719_45144# 4.95e-21
C9325 a_13259_45724# a_13017_45260# 0.078313f
C9326 a_n237_47217# a_10150_46912# 2.7e-19
C9327 a_n1741_47186# a_6969_46634# 7.57e-20
C9328 a_5815_47464# a_4651_46660# 0.001772f
C9329 a_6151_47436# a_4646_46812# 0.153739f
C9330 a_6545_47178# a_3877_44458# 0.026367f
C9331 a_n3565_39590# VREF_GND 0.041931f
C9332 a_7754_38636# VDAC_P 3.34e-19
C9333 VDAC_Ni a_8912_37509# 4.77e-20
C9334 a_n4064_37984# EN_VIN_BSTR_P 0.031746f
C9335 a_2063_45854# a_5257_43370# 0.426517f
C9336 a_4915_47217# a_4817_46660# 2.69e-19
C9337 a_4791_45118# a_5167_46660# 0.008966f
C9338 a_n881_46662# a_12891_46348# 0.026595f
C9339 a_8128_46384# a_9804_47204# 0.001612f
C9340 a_n3690_39392# VDD 0.363068f
C9341 a_3754_38470# a_6886_37412# 7.59e-20
C9342 a_22731_47423# a_22612_30879# 9.38e-19
C9343 SMPL_ON_N a_21588_30879# 0.119129f
C9344 a_11453_44696# a_20916_46384# 0.021978f
C9345 a_8530_39574# a_4338_37500# 0.093669f
C9346 a_n3420_37440# a_n2860_37690# 0.002301f
C9347 a_n2946_37690# a_n2302_37690# 6.68e-19
C9348 a_7754_38470# a_5088_37509# 0.394117f
C9349 a_21381_43940# a_4190_30871# 0.023285f
C9350 a_14401_32519# a_21259_43561# 2.5e-19
C9351 a_n97_42460# a_16664_43396# 0.002303f
C9352 en_comp a_22459_39145# 0.415926f
C9353 a_8147_43396# a_8423_43396# 0.00119f
C9354 a_16147_45260# VDD 0.197706f
C9355 a_19319_43548# a_19095_43396# 0.006369f
C9356 a_n2293_43922# a_2351_42308# 3.54e-20
C9357 a_n356_44636# a_8791_42308# 2.77e-19
C9358 a_3626_43646# a_12281_43396# 0.001712f
C9359 a_5891_43370# a_5932_42308# 0.001048f
C9360 a_526_44458# a_1467_44172# 0.041836f
C9361 a_3537_45260# a_5205_44484# 7.92e-19
C9362 a_n2293_45010# a_1307_43914# 0.008547f
C9363 a_n755_45592# a_n2661_43922# 0.037767f
C9364 a_8746_45002# a_10157_44484# 0.003462f
C9365 a_10180_45724# a_10440_44484# 8.08e-21
C9366 a_n357_42282# a_n2293_43922# 0.02281f
C9367 a_5111_44636# a_5691_45260# 0.130044f
C9368 a_5147_45002# a_3232_43370# 0.253159f
C9369 a_9290_44172# a_10729_43914# 0.042243f
C9370 a_16327_47482# a_21356_42826# 0.003181f
C9371 a_22612_30879# a_14209_32519# 0.059911f
C9372 a_n2661_45010# a_375_42282# 0.017053f
C9373 a_9049_44484# a_8975_43940# 0.001423f
C9374 a_n1151_42308# a_526_44458# 0.003737f
C9375 a_3160_47472# a_n1925_42282# 2.98e-19
C9376 a_33_46660# a_765_45546# 4.44e-20
C9377 a_12861_44030# a_18819_46122# 0.001599f
C9378 a_13717_47436# a_18985_46122# 1.33e-21
C9379 a_9067_47204# a_6945_45028# 0.014009f
C9380 a_19594_46812# a_19636_46660# 0.009543f
C9381 a_n881_46662# a_805_46414# 0.011286f
C9382 a_n1613_43370# a_1208_46090# 0.002092f
C9383 a_4883_46098# a_5937_45572# 0.015486f
C9384 a_10227_46804# a_12594_46348# 0.001992f
C9385 a_11599_46634# a_17583_46090# 0.031836f
C9386 a_15507_47210# a_15682_46116# 3.39e-19
C9387 a_n971_45724# a_8034_45724# 0.027525f
C9388 a_n237_47217# a_8062_46482# 0.001342f
C9389 a_10150_46912# a_8270_45546# 4.81e-19
C9390 a_8492_46660# a_8601_46660# 0.007416f
C9391 a_8667_46634# a_8846_46660# 0.007399f
C9392 a_2063_45854# a_1337_46116# 4.29e-19
C9393 a_15811_47375# a_2324_44458# 0.001263f
C9394 a_1209_43370# a_1067_42314# 4.05e-20
C9395 a_15493_43396# a_18727_42674# 1.59e-21
C9396 a_1847_42826# a_2075_43172# 0.103349f
C9397 a_4190_30871# a_18249_42858# 0.029356f
C9398 a_14021_43940# a_15486_42560# 6.52e-22
C9399 a_n1557_42282# COMP_P 0.123881f
C9400 a_5649_42852# a_5534_30871# 0.234793f
C9401 a_743_42282# a_18083_42858# 1.7e-19
C9402 a_4361_42308# a_15567_42826# 3.24e-20
C9403 a_10334_44484# VDD 0.19332f
C9404 a_3090_45724# a_7309_42852# 1e-19
C9405 a_n755_45592# a_n447_43370# 0.017822f
C9406 a_n357_42282# a_n97_42460# 0.900712f
C9407 a_22223_45036# a_19721_31679# 2.55e-19
C9408 a_2437_43646# a_20512_43084# 3.76e-21
C9409 a_17339_46660# a_18599_43230# 0.001489f
C9410 SMPL_ON_P a_n4064_37984# 7.33e-21
C9411 a_1423_45028# a_5891_43370# 0.301629f
C9412 a_13507_46334# a_20107_42308# 5.01e-19
C9413 a_n2293_46634# a_7227_42308# 7.23e-22
C9414 a_n2442_46660# a_6123_31319# 6.51e-21
C9415 a_13249_42308# a_11341_43940# 0.032308f
C9416 a_11691_44458# a_19929_45028# 5.24e-19
C9417 a_22959_45036# a_18114_32519# 0.004401f
C9418 a_1307_43914# a_9313_44734# 0.021168f
C9419 a_n2438_43548# a_2277_45546# 9.99e-20
C9420 a_12359_47026# a_10809_44734# 0.010386f
C9421 a_13059_46348# a_2324_44458# 0.0606f
C9422 a_n1853_46287# a_472_46348# 1.54e-20
C9423 a_11415_45002# a_3483_46348# 0.057381f
C9424 a_10227_46804# a_15037_45618# 0.012118f
C9425 a_11599_46634# a_8696_44636# 0.003698f
C9426 a_171_46873# a_n443_42852# 5.11e-19
C9427 a_n743_46660# a_1990_45899# 5.84e-19
C9428 a_n2293_46098# a_1208_46090# 0.002845f
C9429 a_1799_45572# a_n755_45592# 0.024036f
C9430 a_n2661_46098# a_n357_42282# 6.61e-20
C9431 a_8035_47026# a_8049_45260# 6.19e-20
C9432 a_16327_47482# a_15765_45572# 0.048221f
C9433 a_n1741_47186# a_3357_43084# 0.03857f
C9434 a_n1423_46090# a_n1076_46494# 0.051162f
C9435 a_18504_43218# a_18695_43230# 4.61e-19
C9436 a_n97_42460# CAL_N 8.11e-21
C9437 a_10083_42826# a_10533_42308# 0.003061f
C9438 a_5649_42852# a_19647_42308# 1.31e-19
C9439 a_4361_42308# a_20712_42282# 0.013294f
C9440 a_13678_32519# a_13258_32519# 0.055554f
C9441 a_13467_32519# a_7174_31319# 6e-19
C9442 a_8199_44636# a_5934_30871# 0.159294f
C9443 a_17613_45144# a_11341_43940# 7.11e-21
C9444 a_19778_44110# a_20269_44172# 1.25e-19
C9445 a_2382_45260# a_2982_43646# 0.468592f
C9446 a_8103_44636# a_7845_44172# 2.71e-19
C9447 a_11827_44484# a_18079_43940# 0.002983f
C9448 a_16922_45042# a_15493_43940# 0.019907f
C9449 a_18184_42460# a_19862_44208# 0.028217f
C9450 a_5147_45002# a_4905_42826# 3.8e-19
C9451 a_9313_44734# a_18579_44172# 3.89e-19
C9452 a_n2661_42834# a_11967_42832# 2.11e-20
C9453 a_11691_44458# a_14955_43940# 0.00153f
C9454 a_n863_45724# a_945_42968# 0.003329f
C9455 a_5063_47570# DATA[2] 7.59e-20
C9456 a_n913_45002# a_7287_43370# 9.35e-21
C9457 a_5159_47243# VDD 2.18e-20
C9458 a_5883_43914# a_7281_43914# 0.029594f
C9459 a_3232_43370# a_4093_43548# 0.091441f
C9460 a_18494_42460# a_19478_44306# 6.46e-21
C9461 a_4955_46873# a_4558_45348# 2.33e-19
C9462 a_11309_47204# a_n2661_43370# 8.95e-20
C9463 a_15227_44166# a_18909_45814# 6.54e-21
C9464 a_18834_46812# a_18691_45572# 2.2e-20
C9465 a_10903_43370# a_n443_42852# 0.176275f
C9466 a_n2438_43548# a_626_44172# 0.025123f
C9467 a_n2293_46634# a_2903_45348# 5.43e-19
C9468 a_5164_46348# a_6511_45714# 4.12e-21
C9469 a_6165_46155# a_5907_45546# 6.1e-19
C9470 a_5807_45002# a_5837_45028# 0.006254f
C9471 a_5385_46902# a_3537_45260# 8.42e-22
C9472 a_12741_44636# a_13527_45546# 1.3e-21
C9473 a_2324_44458# a_3218_45724# 1.93e-20
C9474 a_8349_46414# a_2711_45572# 8.3e-21
C9475 a_n971_45724# a_n998_44484# 5.1e-19
C9476 a_4185_45028# a_3775_45552# 5.74e-20
C9477 a_4883_46098# a_11691_44458# 3.07e-20
C9478 a_19466_46812# a_18479_45785# 0.009818f
C9479 a_11415_45002# a_14495_45572# 1.03e-19
C9480 a_3877_44458# a_4927_45028# 1.65e-20
C9481 a_4646_46812# a_5111_44636# 0.078281f
C9482 a_4651_46660# a_5147_45002# 3e-19
C9483 a_15051_42282# a_15803_42450# 0.043619f
C9484 a_15486_42560# a_15764_42576# 0.118759f
C9485 a_14113_42308# a_15959_42545# 0.036113f
C9486 a_6123_31319# a_13258_32519# 0.00105f
C9487 a_791_42968# VDD 0.128737f
C9488 a_n3674_37592# a_n4334_39392# 6.37e-20
C9489 a_5342_30871# a_n923_35174# 0.00897f
C9490 a_2127_44172# a_2253_43940# 0.143754f
C9491 a_895_43940# a_1241_43940# 0.054548f
C9492 a_2479_44172# a_1443_43940# 8.09e-20
C9493 a_12741_44636# EN_OFFSET_CAL 0.230064f
C9494 a_n2810_45572# a_n4209_39304# 0.020327f
C9495 a_n1423_46090# VDD 0.227012f
C9496 a_9313_44734# a_9396_43370# 4.33e-20
C9497 a_10729_43914# a_10807_43548# 0.238591f
C9498 a_20193_45348# a_13678_32519# 0.055785f
C9499 a_11823_42460# a_12563_42308# 0.039858f
C9500 a_3537_45260# a_3863_42891# 5.22e-20
C9501 a_10193_42453# a_15051_42282# 5.96e-19
C9502 a_n2293_42834# a_8387_43230# 4.23e-19
C9503 a_18579_44172# a_20974_43370# 2.18e-20
C9504 a_n1059_45260# a_11136_42852# 0.004379f
C9505 a_9290_44172# a_1423_45028# 0.005536f
C9506 a_6667_45809# a_6977_45572# 0.013793f
C9507 a_6598_45938# a_6905_45572# 3.69e-19
C9508 a_6472_45840# a_8697_45822# 8.93e-21
C9509 a_526_44458# a_327_44734# 0.076983f
C9510 a_n1925_42282# a_413_45260# 4.11e-20
C9511 a_11415_45002# a_17719_45144# 0.006388f
C9512 a_12741_44636# a_16922_45042# 0.139755f
C9513 a_19443_46116# a_19431_45546# 1.05e-19
C9514 a_16327_47482# a_19328_44172# 0.0072f
C9515 a_12861_44030# a_11341_43940# 0.064865f
C9516 a_14275_46494# a_14537_43396# 9.72e-21
C9517 a_6945_45028# a_7276_45260# 0.00333f
C9518 a_2711_45572# a_8120_45572# 7.29e-19
C9519 a_10053_45546# a_10180_45724# 0.144403f
C9520 a_4185_45028# a_5093_45028# 9.16e-19
C9521 a_22612_30879# a_17730_32519# 0.060497f
C9522 a_8049_45260# a_21542_45572# 4.32e-19
C9523 a_768_44030# a_895_43940# 0.06559f
C9524 a_2324_44458# a_13556_45296# 0.026317f
C9525 a_7499_43078# a_8746_45002# 0.153858f
C9526 a_9049_44484# a_10193_42453# 6.5e-20
C9527 a_5257_43370# a_n2661_42834# 0.01982f
C9528 a_n1613_43370# a_7542_44172# 0.007527f
C9529 a_14976_45028# a_14539_43914# 2.57e-19
C9530 a_19787_47423# a_20990_47178# 4.61e-20
C9531 a_n2302_37984# a_n2216_37984# 0.011479f
C9532 a_15051_42282# VDD 0.461307f
C9533 a_14113_42308# RST_Z 2.01e-19
C9534 a_n2109_47186# a_n2312_38680# 4.37e-19
C9535 a_n2497_47436# a_n1021_46688# 9.22e-19
C9536 a_10227_46804# a_12465_44636# 0.057431f
C9537 a_18597_46090# a_13507_46334# 0.093881f
C9538 a_18479_47436# a_4883_46098# 0.038695f
C9539 a_n4064_39072# a_n3420_37440# 0.051893f
C9540 a_n3420_39072# a_n4064_37440# 0.047151f
C9541 a_n1920_47178# a_n2104_46634# 3.21e-19
C9542 a_n815_47178# a_n2661_46634# 0.003247f
C9543 SMPL_ON_P a_n2442_46660# 0.092029f
C9544 a_2063_45854# a_5807_45002# 0.074286f
C9545 a_4915_47217# a_11309_47204# 0.045252f
C9546 a_6151_47436# a_9804_47204# 0.095181f
C9547 a_6545_47178# a_8128_46384# 5.48e-21
C9548 a_7903_47542# a_n881_46662# 0.178742f
C9549 a_n4064_39616# VDAC_P 0.007212f
C9550 a_4958_30871# C5_P_btm 1.35e-19
C9551 a_6575_47204# a_n1613_43370# 0.005913f
C9552 a_20679_44626# a_21195_42852# 7.08e-20
C9553 a_18579_44172# a_18599_43230# 1.99e-20
C9554 a_19279_43940# a_19987_42826# 1.18e-19
C9555 a_3422_30871# a_16795_42852# 2.85e-21
C9556 a_n2956_37592# a_n2216_38778# 1.2e-19
C9557 a_9049_44484# VDD 0.680993f
C9558 a_12429_44172# a_743_42282# 3.38e-21
C9559 a_11341_43940# a_19700_43370# 4.45e-20
C9560 a_3905_42865# a_2905_42968# 2.41e-19
C9561 a_15493_43396# a_17486_43762# 3.67e-19
C9562 a_2998_44172# a_3935_42891# 3.35e-21
C9563 a_3600_43914# a_3681_42891# 2.17e-20
C9564 a_15493_43940# a_15743_43084# 0.206331f
C9565 a_n97_42460# a_n144_43396# 1.59e-19
C9566 a_4093_43548# a_4905_42826# 5.66e-20
C9567 a_1568_43370# a_n1557_42282# 3.82e-20
C9568 a_1049_43396# a_1427_43646# 0.010711f
C9569 a_4235_43370# a_3080_42308# 0.098951f
C9570 a_16375_45002# a_18248_44752# 1.65e-21
C9571 a_10490_45724# a_n2661_43370# 7.79e-21
C9572 a_13507_46334# a_743_42282# 0.026943f
C9573 a_1138_42852# a_2479_44172# 4.8e-21
C9574 a_n2293_46098# a_7542_44172# 5.6e-21
C9575 a_2437_43646# a_n2661_45010# 0.15182f
C9576 a_22591_45572# a_20447_31679# 7.75e-19
C9577 a_4791_45118# a_5111_42852# 0.012003f
C9578 a_16327_47482# a_20749_43396# 0.008166f
C9579 a_n2293_46634# a_6643_43396# 7e-19
C9580 a_15227_44166# a_14761_44260# 7.89e-21
C9581 a_13259_45724# a_18374_44850# 0.002311f
C9582 a_11322_45546# a_11361_45348# 9.02e-20
C9583 a_17715_44484# a_11967_42832# 0.081495f
C9584 a_13661_43548# a_15095_43370# 1.48e-20
C9585 a_n23_45546# a_n2661_44458# 5.06e-22
C9586 a_n755_45592# a_n452_44636# 0.015469f
C9587 a_n357_42282# a_742_44458# 0.085409f
C9588 a_15037_45618# a_1307_43914# 1.49e-21
C9589 a_15765_45572# a_14537_43396# 3.49e-19
C9590 a_15599_45572# a_15415_45028# 5.19e-19
C9591 a_8696_44636# a_13348_45260# 1.38e-20
C9592 a_19963_31679# a_22959_45572# 0.020087f
C9593 a_n2840_46090# a_n4318_39768# 9.97e-22
C9594 a_3815_47204# a_1823_45246# 6.25e-21
C9595 C3_P_btm VREF 0.984942f
C9596 a_13507_46334# a_19123_46287# 0.034113f
C9597 a_20990_47178# a_20107_46660# 2.98e-20
C9598 a_10227_46804# a_20528_46660# 1.1e-20
C9599 C4_P_btm VREF_GND 0.671882f
C9600 C5_P_btm VCM 0.719982f
C9601 a_n237_47217# a_6419_46155# 0.029086f
C9602 a_n1741_47186# a_9625_46129# 6.6e-20
C9603 a_n971_45724# a_8016_46348# 0.029312f
C9604 a_n443_46116# a_805_46414# 9.4e-20
C9605 a_11453_44696# a_16751_46987# 1.13e-21
C9606 a_3177_46902# a_3633_46660# 4.2e-19
C9607 a_n743_46660# a_6969_46634# 1.5e-19
C9608 a_2063_45854# a_3699_46348# 0.002997f
C9609 a_3160_47472# a_2698_46116# 4.19e-19
C9610 a_2905_45572# a_2804_46116# 3.04e-19
C9611 a_2952_47436# a_3147_46376# 1.09e-19
C9612 a_n1151_42308# a_2521_46116# 2.53e-20
C9613 a_584_46384# a_4185_45028# 5.71e-19
C9614 a_12549_44172# a_16292_46812# 0.013094f
C9615 C1_P_btm VIN_P 0.39234f
C9616 a_2107_46812# a_8492_46660# 2.24e-20
C9617 a_5807_45002# a_12469_46902# 0.003304f
C9618 C9_N_btm VDD 0.345685f
C9619 a_12465_44636# a_17339_46660# 6.05e-22
C9620 a_20512_43084# a_19511_42282# 7.2e-20
C9621 a_3422_30871# a_21335_42336# 0.002526f
C9622 a_21487_43396# a_13467_32519# 0.152042f
C9623 a_9145_43396# a_12545_42858# 6.25e-19
C9624 a_4905_42826# a_5457_43172# 2.02e-20
C9625 a_8685_43396# a_5534_30871# 4.59e-19
C9626 a_9885_43646# a_10083_42826# 1.33e-19
C9627 a_4190_30871# a_5649_42852# 0.434284f
C9628 a_n1613_43370# a_n1630_35242# 3.68e-19
C9629 a_2324_44458# a_6293_42852# 0.002463f
C9630 a_n443_42852# a_14955_43940# 5.77e-21
C9631 a_20205_31679# a_14021_43940# 1.01e-20
C9632 a_7229_43940# a_6298_44484# 0.028942f
C9633 a_5111_44636# a_10057_43914# 0.002052f
C9634 a_15861_45028# a_11967_42832# 6.28e-20
C9635 a_12741_44636# a_15743_43084# 2.11e-20
C9636 a_3090_45724# a_7765_42852# 2.34e-20
C9637 a_n357_42282# a_21115_43940# 1.83e-21
C9638 a_3232_43370# a_10157_44484# 0.049345f
C9639 a_6431_45366# a_5883_43914# 1.65e-19
C9640 a_7705_45326# a_5343_44458# 2.71e-19
C9641 a_5937_45572# a_8685_43396# 7.97e-21
C9642 a_2747_46873# a_n755_45592# 1.74e-20
C9643 a_n1613_43370# a_n2661_45546# 0.029057f
C9644 a_10227_46804# a_2711_45572# 0.130695f
C9645 a_3177_46902# a_526_44458# 0.001189f
C9646 a_7577_46660# a_2324_44458# 1.05e-20
C9647 a_14513_46634# a_11415_45002# 2.15e-20
C9648 a_20107_46660# a_20273_46660# 0.608339f
C9649 a_19123_46287# a_20623_46660# 1.73e-20
C9650 a_4883_46098# a_n443_42852# 0.074259f
C9651 a_6755_46942# a_11133_46155# 1.21e-19
C9652 a_6151_47436# a_10180_45724# 9.87e-21
C9653 a_5807_45002# a_14383_46116# 0.007691f
C9654 a_5342_30871# a_14853_42852# 5e-21
C9655 a_15781_43660# a_15959_42545# 2.85e-19
C9656 a_3905_42865# VDD 0.788273f
C9657 a_16243_43396# a_14113_42308# 3.98e-19
C9658 a_791_42968# a_n784_42308# 1.7e-19
C9659 a_13467_32519# a_5932_42308# 1.17e-19
C9660 a_743_42282# a_7227_42308# 0.008196f
C9661 a_4361_42308# a_6171_42473# 0.008302f
C9662 a_8975_43940# a_12553_44484# 1.95e-20
C9663 a_5815_47464# VDD 0.399354f
C9664 a_11827_44484# a_17730_32519# 0.009382f
C9665 a_3815_47204# DATA[2] 0.022461f
C9666 a_n443_42852# a_5649_42852# 8.75e-19
C9667 a_n357_42282# a_n901_43156# 0.008049f
C9668 a_10903_43370# a_14635_42282# 1.8e-20
C9669 SMPL_ON_N a_22469_39537# 0.017847f
C9670 a_14539_43914# a_15433_44458# 2.67e-20
C9671 a_15004_44636# a_15463_44811# 6.64e-19
C9672 a_12607_44458# a_12189_44484# 2.07e-20
C9673 a_6109_44484# a_5891_43370# 3.31e-20
C9674 a_7640_43914# a_8375_44464# 5.23e-19
C9675 a_11787_45002# a_11341_43940# 1.39e-22
C9676 a_13249_42308# a_10341_43396# 0.040208f
C9677 a_4185_45028# a_14097_32519# 0.020305f
C9678 a_n1151_42308# DATA[5] 0.006171f
C9679 a_16751_45260# a_15682_43940# 3.8e-19
C9680 a_n1613_43370# a_5205_44484# 0.551795f
C9681 a_n2472_46090# a_n2472_45546# 0.025171f
C9682 a_n2293_46098# a_n2661_45546# 3.03243f
C9683 a_n743_46660# a_3357_43084# 0.034228f
C9684 a_11453_44696# a_14797_45144# 0.002114f
C9685 a_8199_44636# a_9751_46155# 7.99e-20
C9686 a_n2840_46090# a_n2956_38216# 0.004667f
C9687 a_13607_46688# a_13527_45546# 8.43e-20
C9688 a_17339_46660# a_2711_45572# 0.02331f
C9689 a_765_45546# a_1609_45572# 1.84e-19
C9690 a_n881_46662# a_6431_45366# 0.177591f
C9691 a_11133_46155# a_8049_45260# 0.001208f
C9692 a_9625_46129# a_10586_45546# 9.22e-19
C9693 a_3483_46348# a_13259_45724# 0.230226f
C9694 a_3090_45724# a_11823_42460# 0.089008f
C9695 a_768_44030# a_3065_45002# 0.288972f
C9696 a_n2956_39304# a_n1379_46482# 9.59e-21
C9697 a_12465_44636# a_1307_43914# 0.022149f
C9698 a_1606_42308# a_5742_30871# 3.46204f
C9699 a_18707_42852# a_18727_42674# 2.69e-19
C9700 a_n784_42308# a_15051_42282# 1.37e-19
C9701 a_6171_42473# a_6761_42308# 3.88e-19
C9702 a_4921_42308# a_5934_30871# 3.08e-20
C9703 a_19333_46634# VDD 0.199048f
C9704 a_18834_46812# START 0.001199f
C9705 a_n2661_44458# a_7287_43370# 3.62e-21
C9706 a_15227_44166# RST_Z 2.45e-20
C9707 a_3537_45260# a_4520_42826# 0.066648f
C9708 a_n913_45002# a_12089_42308# 0.038293f
C9709 a_n1059_45260# a_12545_42858# 0.011705f
C9710 a_n2017_45002# a_13113_42826# 1.01e-19
C9711 a_n2956_39304# a_n4064_39072# 0.054199f
C9712 a_n2956_38680# a_n2946_39072# 0.004064f
C9713 a_20159_44458# a_20269_44172# 0.001015f
C9714 a_5343_44458# a_2982_43646# 1.31e-19
C9715 a_5244_44056# a_5013_44260# 0.094334f
C9716 a_3905_42865# a_5495_43940# 1.51e-20
C9717 a_18579_44172# a_17737_43940# 6.7e-20
C9718 a_12816_46660# CLK 6.39e-21
C9719 a_n443_42852# a_7963_42308# 4.91e-20
C9720 a_n357_42282# a_10533_42308# 7.55e-20
C9721 a_11691_44458# a_8685_43396# 5.46e-21
C9722 a_11967_42832# a_20623_43914# 7.1e-20
C9723 a_n699_43396# a_3626_43646# 2.23e-19
C9724 a_n755_45592# a_3638_45822# 9.05e-19
C9725 a_n2293_46098# a_5205_44484# 0.001237f
C9726 a_1823_45246# a_2382_45260# 0.801932f
C9727 a_11189_46129# a_3357_43084# 3.29e-22
C9728 a_13259_45724# a_14495_45572# 0.020864f
C9729 a_10586_45546# a_9159_45572# 1.71e-19
C9730 a_167_45260# a_1667_45002# 0.05322f
C9731 a_2698_46116# a_413_45260# 9.42e-21
C9732 a_5807_45002# a_n2661_42834# 5.92e-21
C9733 a_11415_45002# a_11963_45334# 0.031636f
C9734 a_584_46384# a_1241_44260# 1.06e-19
C9735 a_10903_43370# a_2437_43646# 5.87e-20
C9736 a_n4209_39304# a_n4251_39392# 0.00226f
C9737 a_1736_39587# comp_n 0.004824f
C9738 a_n4209_39590# a_n2302_38778# 7.57e-20
C9739 a_1606_42308# C0_dummy_P_btm 0.007541f
C9740 a_n784_42308# C9_N_btm 9.31e-20
C9741 a_14097_32519# VREF_GND 0.047244f
C9742 a_n3565_39304# a_n4064_39072# 0.344587f
C9743 a_n4064_39616# a_n4334_38528# 8.04e-19
C9744 a_7174_31319# a_2113_38308# 8.18e-20
C9745 a_n961_42308# VDD 0.24416f
C9746 a_5815_47464# a_6491_46660# 0.003594f
C9747 a_n1151_42308# a_13381_47204# 7.76e-20
C9748 a_4915_47217# a_7227_47204# 0.059062f
C9749 a_4791_45118# a_6575_47204# 8.32e-20
C9750 a_6151_47436# a_6545_47178# 0.39775f
C9751 a_3160_47472# a_n1435_47204# 5e-19
C9752 a_19479_31679# a_22775_42308# 3.61e-21
C9753 a_20062_46116# VDD 4.6e-19
C9754 a_20512_43084# a_21259_43561# 0.002989f
C9755 a_19808_44306# a_19319_43548# 1.05e-19
C9756 a_n2017_45002# a_18214_42558# 2.04e-19
C9757 a_n913_45002# a_18907_42674# 1.21e-19
C9758 a_n1059_45260# a_19332_42282# 8.78e-20
C9759 a_n2661_43922# a_10083_42826# 6.13e-21
C9760 a_n2293_43922# a_8952_43230# 2.5e-21
C9761 a_n2293_42834# a_1606_42308# 7.69e-19
C9762 a_8333_44056# a_8685_43396# 1.53e-20
C9763 en_comp a_17303_42282# 1.29e-19
C9764 a_20692_30879# C10_N_btm 2.44e-19
C9765 a_20835_44721# a_20749_43396# 2e-20
C9766 a_18494_42460# a_20256_43172# 0.052522f
C9767 a_n2661_43370# a_n3674_37592# 2.27e-20
C9768 a_1307_43914# a_8515_42308# 1.29e-21
C9769 a_9313_44734# a_13635_43156# 0.013436f
C9770 a_2107_46812# a_9420_43940# 1.23e-19
C9771 a_2957_45546# a_2809_45028# 6.81e-20
C9772 a_18985_46122# a_18248_44752# 4.72e-21
C9773 a_18819_46122# a_18287_44626# 3.39e-21
C9774 a_17715_44484# a_18989_43940# 1.14e-20
C9775 a_12741_44636# a_16789_44484# 0.009606f
C9776 a_16147_45260# a_18479_45785# 0.005418f
C9777 a_17786_45822# a_18341_45572# 3.4e-19
C9778 a_12861_44030# a_10341_43396# 0.018259f
C9779 a_22612_30879# a_17538_32519# 0.060018f
C9780 a_2711_45572# a_1307_43914# 0.187968f
C9781 a_10809_44734# a_12883_44458# 2.59e-19
C9782 a_768_44030# a_458_43396# 0.001002f
C9783 a_5164_46348# a_5608_44484# 4.14e-20
C9784 a_16375_45002# a_16922_45042# 0.170835f
C9785 a_13259_45724# a_17719_45144# 0.039832f
C9786 a_8199_44636# a_8855_44734# 0.002934f
C9787 a_8016_46348# a_9313_44734# 0.020204f
C9788 a_8568_45546# a_6171_45002# 0.005143f
C9789 a_7499_43078# a_3232_43370# 0.318423f
C9790 a_3483_46348# a_n2661_43922# 0.038814f
C9791 a_526_44458# a_4223_44672# 1.22e-19
C9792 a_n3420_37440# VDD 2.26579f
C9793 a_4883_46098# a_10554_47026# 1.36e-20
C9794 a_n2312_38680# a_n1925_46634# 0.004049f
C9795 a_n2293_46634# a_n743_46660# 0.001475f
C9796 a_n2442_46660# a_n2438_43548# 0.002667f
C9797 VDAC_P C0_P_btm 0.322595f
C9798 a_n881_46662# a_4817_46660# 1.02e-19
C9799 a_12861_44030# a_12991_46634# 0.001474f
C9800 a_n1435_47204# a_13607_46688# 7.18e-19
C9801 a_n1613_43370# a_5385_46902# 0.182522f
C9802 CAL_P EN_VIN_BSTR_N 0.049856f
C9803 VDAC_N C0_dummy_N_btm 0.287929f
C9804 a_13507_46334# a_6755_46942# 0.075659f
C9805 a_11599_46634# a_11813_46116# 0.106062f
C9806 a_n2661_46634# a_171_46873# 0.007801f
C9807 a_n1151_42308# a_13170_46660# 1.42e-19
C9808 a_4915_47217# a_12156_46660# 7.15e-20
C9809 a_8128_46384# a_3877_44458# 1.82e-21
C9810 a_15095_43370# a_15037_43396# 0.001617f
C9811 a_n97_42460# a_8952_43230# 6.13e-21
C9812 a_3905_42865# a_n784_42308# 7.08e-21
C9813 a_453_43940# a_961_42354# 2.06e-22
C9814 a_5147_45002# VDD 0.574918f
C9815 a_n3674_39768# a_n4318_38216# 0.032347f
C9816 a_413_45260# EN_OFFSET_CAL 0.114452f
C9817 a_10341_43396# a_19700_43370# 0.013451f
C9818 a_15781_43660# a_16243_43396# 7.62e-21
C9819 a_15681_43442# a_16547_43609# 2.74e-20
C9820 a_6171_45002# a_n2661_43370# 2.37006f
C9821 a_n755_45592# a_n809_44244# 0.404418f
C9822 a_n357_42282# a_n984_44318# 1.05e-19
C9823 a_2711_45572# a_18579_44172# 0.170319f
C9824 a_15227_44166# a_16243_43396# 0.002283f
C9825 a_7229_43940# a_7418_45067# 0.006955f
C9826 a_7276_45260# a_7735_45067# 6.64e-19
C9827 a_8191_45002# a_8488_45348# 0.004422f
C9828 a_13249_42308# a_n2293_43922# 6.65e-19
C9829 a_310_45028# a_175_44278# 1.47e-19
C9830 a_10216_45572# a_5891_43370# 3.99e-20
C9831 a_n863_45724# a_1414_42308# 0.711805f
C9832 a_n2661_45546# a_2675_43914# 1.1e-21
C9833 a_11823_42460# a_14815_43914# 2.04e-19
C9834 a_13059_46348# a_14579_43548# 0.171744f
C9835 a_16327_47482# a_19518_43218# 0.002315f
C9836 a_2107_46812# a_5497_46414# 0.003373f
C9837 a_584_46384# a_997_45618# 2.73e-20
C9838 a_2063_45854# a_n755_45592# 0.074611f
C9839 a_3524_46660# a_1823_45246# 2.12e-19
C9840 a_4791_45118# a_n2661_45546# 0.012117f
C9841 a_13487_47204# a_13259_45724# 1.12e-20
C9842 a_19466_46812# a_19692_46634# 0.001654f
C9843 a_12991_46634# a_14180_46812# 2e-20
C9844 a_13607_46688# a_13885_46660# 0.11044f
C9845 a_12816_46660# a_14035_46660# 5.75e-20
C9846 a_n2661_46634# a_10903_43370# 0.663878f
C9847 a_2124_47436# a_1848_45724# 6.36e-22
C9848 a_n971_45724# a_n1013_45572# 0.004752f
C9849 a_13507_46334# a_8049_45260# 0.086137f
C9850 a_n1613_43370# a_n1533_46116# 0.012221f
C9851 a_n881_46662# a_n722_46482# 6.07e-19
C9852 a_11309_47204# a_10809_44734# 5.65e-20
C9853 a_2443_46660# a_2804_46116# 0.006742f
C9854 a_2609_46660# a_2698_46116# 4.2e-21
C9855 a_n743_46660# a_9625_46129# 0.206271f
C9856 a_12549_44172# a_6945_45028# 0.028827f
C9857 a_13747_46662# a_15682_46116# 0.001312f
C9858 a_5807_45002# a_17715_44484# 0.045558f
C9859 a_14311_47204# a_14383_46116# 9.92e-21
C9860 a_4520_42826# a_4649_43172# 0.010132f
C9861 a_19741_43940# a_19647_42308# 5.24e-21
C9862 a_3539_42460# a_5742_30871# 2.25e-20
C9863 a_3626_43646# a_11551_42558# 0.005206f
C9864 a_5649_42852# a_14635_42282# 7.52e-20
C9865 a_16414_43172# a_16795_42852# 1.48e-19
C9866 a_2982_43646# a_12563_42308# 2.07e-19
C9867 a_n2017_45002# a_n2661_42282# 0.035164f
C9868 a_n443_42852# a_8685_43396# 0.281116f
C9869 a_13249_42308# a_n97_42460# 0.067568f
C9870 a_n2661_44458# a_n23_44458# 0.006363f
C9871 a_16375_45002# a_15743_43084# 1.19e-20
C9872 a_n1925_42282# a_n13_43084# 5.01e-21
C9873 a_20107_45572# a_20935_43940# 1.76e-21
C9874 a_16147_45260# a_14021_43940# 2.27e-20
C9875 a_10157_44484# a_8975_43940# 0.045547f
C9876 a_10334_44484# a_10057_43914# 0.002134f
C9877 a_n1917_44484# a_n1809_44850# 0.057222f
C9878 a_n1699_44726# a_n1190_44850# 2.6e-19
C9879 a_n2267_44484# a_n1821_44484# 2.28e-19
C9880 a_5111_44636# a_5013_44260# 0.029412f
C9881 a_5147_45002# a_5495_43940# 0.086203f
C9882 a_3232_43370# a_3600_43914# 0.087298f
C9883 a_21363_45546# a_19862_44208# 3.42e-20
C9884 a_4927_45028# a_5244_44056# 6.1e-21
C9885 a_3537_45260# a_7281_43914# 1.36e-20
C9886 a_22612_30879# a_22465_38105# 9.58e-19
C9887 a_4185_45028# a_22959_42860# 0.013205f
C9888 a_4883_46098# a_2437_43646# 0.458866f
C9889 a_13507_46334# a_19479_31679# 0.061466f
C9890 a_21177_47436# a_3357_43084# 5.54e-20
C9891 a_8199_44636# a_10903_43370# 8.9e-20
C9892 a_n1641_46494# a_n1736_46482# 0.049827f
C9893 a_n2293_46098# a_n1533_46116# 0.002776f
C9894 a_n2661_46634# a_12016_45572# 3.65e-19
C9895 a_4791_45118# a_5205_44484# 0.053467f
C9896 a_n1151_42308# a_8953_45002# 1.04e-19
C9897 a_13059_46348# a_12839_46116# 0.098052f
C9898 a_14513_46634# a_13259_45724# 2.83e-21
C9899 a_18597_46090# a_21297_45572# 4.45e-19
C9900 a_16327_47482# a_n913_45002# 0.137194f
C9901 a_9823_46155# a_10355_46116# 0.001471f
C9902 a_n1423_46090# a_n1545_46494# 3.16e-19
C9903 a_10467_46802# a_2711_45572# 2.47e-20
C9904 a_19692_46634# a_20205_31679# 0.001591f
C9905 a_n881_46662# a_18691_45572# 3.57e-20
C9906 a_n1435_47204# a_413_45260# 0.025027f
C9907 a_4915_47217# a_6171_45002# 0.022258f
C9908 a_12549_44172# a_14127_45572# 2.41e-19
C9909 a_768_44030# a_14033_45572# 7.13e-19
C9910 a_13661_43548# a_8696_44636# 0.049791f
C9911 a_13747_46662# a_16680_45572# 0.047612f
C9912 a_5807_45002# a_15861_45028# 3.23e-19
C9913 a_9625_46129# a_11189_46129# 0.003371f
C9914 a_2107_46812# a_9241_45822# 5.82e-21
C9915 a_22165_42308# a_17303_42282# 0.095988f
C9916 a_n1736_42282# a_n1630_35242# 0.071684f
C9917 COMP_P a_n3674_37592# 0.054748f
C9918 a_3080_42308# C9_N_btm 9.33e-20
C9919 a_4093_43548# VDD 0.216874f
C9920 a_n473_42460# a_196_42282# 2.5e-19
C9921 a_n961_42308# a_n784_42308# 0.154417f
C9922 a_n3674_39304# a_n4209_38502# 1.61e-20
C9923 a_n2017_45002# a_16823_43084# 5.82e-19
C9924 a_11787_45002# a_10341_43396# 1.52e-22
C9925 a_n699_43396# a_3052_44056# 1.83e-19
C9926 a_n2293_43922# a_n1441_43940# 1.93e-20
C9927 a_n2661_43922# a_261_44278# 3.53e-19
C9928 a_n2661_42834# a_n822_43940# 1.42e-19
C9929 a_526_44458# a_5742_30871# 2.52e-20
C9930 a_13777_45326# a_13667_43396# 1.06e-21
C9931 a_13556_45296# a_14579_43548# 1.57e-22
C9932 a_18287_44626# a_11341_43940# 8.01e-21
C9933 a_n2293_42834# a_3539_42460# 0.019435f
C9934 a_19279_43940# a_22959_44484# 6.44e-21
C9935 a_5891_43370# a_10405_44172# 0.15894f
C9936 a_20193_45348# a_21205_44306# 0.002474f
C9937 a_n2810_45572# a_n4318_37592# 0.023163f
C9938 a_n2956_38216# a_n2104_42282# 2.12e-20
C9939 a_n357_42282# a_20256_42852# 9.51e-19
C9940 a_7499_43078# a_7573_43172# 0.002331f
C9941 a_3357_43084# a_4361_42308# 3.35e-21
C9942 a_526_44458# a_3260_45572# 2.83e-20
C9943 a_5257_43370# a_5093_45028# 3.11e-21
C9944 a_4915_47217# a_14673_44172# 0.020025f
C9945 a_12861_44030# a_n2293_43922# 0.008309f
C9946 a_20841_46902# a_3357_43084# 0.001309f
C9947 a_13259_45724# a_n357_42282# 0.056511f
C9948 a_12594_46348# a_11682_45822# 4.71e-19
C9949 a_n743_46660# a_16237_45028# 0.038671f
C9950 a_22612_30879# a_19721_31679# 0.068873f
C9951 a_20202_43084# a_20107_45572# 0.002433f
C9952 a_11415_45002# a_18953_45572# 4.28e-19
C9953 a_21188_46660# a_2437_43646# 1.87e-22
C9954 a_13885_46660# a_413_45260# 1.99e-20
C9955 a_20205_31679# a_20692_30879# 0.055565f
C9956 a_768_44030# a_6298_44484# 0.015186f
C9957 a_10809_44734# a_10490_45724# 0.030973f
C9958 a_5066_45546# a_6511_45714# 2.64e-19
C9959 a_8034_45724# a_2711_45572# 0.035334f
C9960 a_n1630_35242# a_n4209_37414# 2.12e-19
C9961 a_n2497_47436# a_n2109_47186# 0.197671f
C9962 a_13258_32519# a_22775_42308# 6.32e-19
C9963 a_n3674_37592# a_n3565_37414# 0.129086f
C9964 a_19511_42282# a_21125_42558# 0.01129f
C9965 a_22400_42852# a_22780_40945# 2e-19
C9966 a_n784_42308# a_n3420_37440# 0.140549f
C9967 a_5932_42308# a_2113_38308# 9.09e-20
C9968 a_5742_30871# a_n4209_38502# 7.41e-22
C9969 a_11691_44458# a_17333_42852# 2.56e-21
C9970 a_11967_42832# a_15095_43370# 0.098499f
C9971 a_n913_45002# a_5267_42460# 0.081794f
C9972 a_n1059_45260# a_5379_42460# 2.17e-19
C9973 a_n2017_45002# a_3497_42558# 0.0024f
C9974 a_10809_44734# START 0.002613f
C9975 a_3905_42865# a_3080_42308# 0.029566f
C9976 a_22959_46124# RST_Z 0.001356f
C9977 a_6298_44484# a_5755_42852# 8.19e-21
C9978 a_13259_45724# CAL_N 0.005414f
C9979 a_1414_42308# a_3540_43646# 0.022584f
C9980 a_13483_43940# a_13565_43940# 0.171361f
C9981 a_n2956_39304# VDD 0.455981f
C9982 a_18184_42460# a_21671_42860# 0.021213f
C9983 a_5343_44458# a_7871_42858# 0.020081f
C9984 a_13661_43548# a_20365_43914# 0.020045f
C9985 a_768_44030# a_10555_44260# 0.00973f
C9986 a_18985_46122# a_16922_45042# 4.99e-21
C9987 a_2698_46116# a_2779_44458# 2.15e-19
C9988 a_12741_44636# a_17970_44736# 9.86e-19
C9989 a_5497_46414# a_n2661_44458# 6.51e-22
C9990 a_167_45260# a_n699_43396# 6.1e-22
C9991 a_1823_45246# a_5343_44458# 2.1e-19
C9992 a_380_45546# a_413_45260# 0.001298f
C9993 a_n1099_45572# a_n37_45144# 1.51e-19
C9994 a_310_45028# a_n143_45144# 1.85e-20
C9995 a_11415_45002# a_18443_44721# 7.02e-22
C9996 a_n2661_45546# a_3429_45260# 5.93e-20
C9997 a_4646_46812# a_3905_42865# 1.17e-19
C9998 a_3090_45724# a_15367_44484# 5.11e-19
C9999 a_n971_45724# a_8791_43396# 8.26e-19
C10000 a_12861_44030# a_n97_42460# 5.48e-20
C10001 a_n443_46116# a_n1557_42282# 0.006023f
C10002 a_584_46384# a_648_43396# 0.050476f
C10003 a_11823_42460# a_13297_45572# 3.1e-20
C10004 a_n2293_45546# a_2382_45260# 0.078874f
C10005 a_n863_45724# a_1667_45002# 0.20954f
C10006 a_11387_46155# a_11691_44458# 1.27e-22
C10007 a_526_44458# a_n2293_42834# 1.7774f
C10008 a_18189_46348# a_17719_45144# 0.002906f
C10009 a_19321_45002# a_19478_44306# 6.34e-21
C10010 a_n3565_39590# VREF 0.417978f
C10011 a_n1741_47186# a_6755_46942# 0.017537f
C10012 a_n237_47217# a_9863_46634# 0.008748f
C10013 a_n1435_47204# a_2609_46660# 5.42e-20
C10014 a_5129_47502# a_4651_46660# 0.002499f
C10015 a_5815_47464# a_4646_46812# 2.49e-19
C10016 a_6151_47436# a_3877_44458# 0.034088f
C10017 a_n4064_38528# C5_P_btm 0.042017f
C10018 a_n3420_39616# VIN_P 0.041227f
C10019 a_7754_38636# a_8912_37509# 5.52e-19
C10020 a_n4064_37984# a_n923_35174# 0.005035f
C10021 a_n1151_42308# a_5275_47026# 0.002003f
C10022 a_4791_45118# a_5385_46902# 0.007028f
C10023 a_n443_46116# a_4817_46660# 0.020386f
C10024 a_4915_47217# a_4955_46873# 0.00958f
C10025 a_2905_45572# a_3878_46660# 2.98e-19
C10026 a_n881_46662# a_11309_47204# 0.028783f
C10027 a_n3565_39304# VDD 0.888861f
C10028 a_n4209_39590# VCM 0.179761f
C10029 a_4883_46098# a_n2661_46634# 0.030655f
C10030 SMPL_ON_N a_20916_46384# 4.07e-20
C10031 a_22731_47423# a_21588_30879# 0.014331f
C10032 a_n3420_37440# a_n2302_37690# 1.28e-19
C10033 a_n4209_37414# a_n3607_37440# 0.002294f
C10034 a_8530_39574# a_3726_37500# 1.35509f
C10035 a_n4334_37440# a_n4251_37440# 0.007692f
C10036 a_7754_38470# a_4338_37500# 0.208284f
C10037 a_3754_38470# a_5700_37509# 0.124176f
C10038 a_n2946_37690# a_n4064_37440# 0.053228f
C10039 a_n97_42460# a_19700_43370# 0.154491f
C10040 a_21381_43940# a_21259_43561# 0.013931f
C10041 en_comp a_22521_40055# 0.260972f
C10042 a_n2293_43922# a_2123_42473# 3.54e-20
C10043 a_20193_45348# a_22775_42308# 1.84e-19
C10044 a_8147_43396# a_8317_43396# 0.001675f
C10045 a_17786_45822# VDD 0.007376f
C10046 a_n356_44636# a_8685_42308# 1.18e-19
C10047 a_5891_43370# a_6171_42473# 2.02e-20
C10048 a_526_44458# a_1115_44172# 0.009996f
C10049 a_3090_45724# a_2982_43646# 1.98e-20
C10050 a_n913_45002# a_14537_43396# 0.003001f
C10051 a_5111_44636# a_4927_45028# 0.134309f
C10052 a_10193_42453# a_10157_44484# 0.001446f
C10053 a_n755_45592# a_n2661_42834# 0.059506f
C10054 a_10180_45724# a_10334_44484# 7.3e-20
C10055 a_n357_42282# a_n2661_43922# 0.088336f
C10056 a_8746_45002# a_9838_44484# 6.4e-19
C10057 a_4558_45348# a_3232_43370# 6.67e-21
C10058 a_5147_45002# a_5691_45260# 0.035185f
C10059 a_9290_44172# a_10405_44172# 0.001407f
C10060 a_16327_47482# a_20922_43172# 0.001914f
C10061 a_21588_30879# a_14209_32519# 0.056208f
C10062 a_n2293_46634# a_4361_42308# 5.54e-21
C10063 a_3537_45260# a_6431_45366# 1.48e-19
C10064 a_15861_45028# a_18315_45260# 1.06e-20
C10065 a_17478_45572# a_17719_45144# 3.17e-19
C10066 a_12465_44636# a_13635_43156# 3.45e-20
C10067 a_7499_43078# a_8975_43940# 0.519621f
C10068 a_3503_45724# a_3363_44484# 8.59e-21
C10069 a_3160_47472# a_526_44458# 0.026069f
C10070 a_2905_45572# a_n1925_42282# 1.51e-21
C10071 a_13717_47436# a_18819_46122# 8.56e-21
C10072 a_12861_44030# a_17957_46116# 0.01013f
C10073 a_6575_47204# a_6945_45028# 0.06375f
C10074 a_19321_45002# a_19636_46660# 6.42e-19
C10075 a_n881_46662# a_472_46348# 0.022658f
C10076 a_n1613_43370# a_805_46414# 2.86e-19
C10077 a_4883_46098# a_8199_44636# 0.242f
C10078 a_11599_46634# a_15682_46116# 1.8289f
C10079 a_15507_47210# a_2324_44458# 4e-21
C10080 a_n237_47217# a_5527_46155# 0.001111f
C10081 a_n1741_47186# a_8049_45260# 0.003545f
C10082 a_6755_46942# a_7832_46660# 0.025487f
C10083 a_9863_46634# a_8270_45546# 7.01e-19
C10084 a_10227_46804# a_12005_46116# 8.43e-19
C10085 a_2063_45854# a_835_46155# 1.26e-20
C10086 a_584_46384# a_1337_46116# 0.044678f
C10087 a_18079_43940# a_18214_42558# 3.88e-21
C10088 a_4190_30871# a_17333_42852# 0.001829f
C10089 a_8685_43396# a_14635_42282# 2.12e-19
C10090 a_14021_43940# a_15051_42282# 1.01e-20
C10091 a_n1557_42282# a_n4318_37592# 0.004047f
C10092 a_13678_32519# a_5534_30871# 0.043974f
C10093 a_743_42282# a_17701_42308# 0.014357f
C10094 a_4361_42308# a_5342_30871# 0.047616f
C10095 a_5649_42852# a_14543_43071# 8.21e-22
C10096 a_10157_44484# VDD 0.174233f
C10097 a_19862_44208# a_17303_42282# 4.5e-20
C10098 a_9165_43940# a_8685_42308# 3.85e-21
C10099 a_n755_45592# a_n1352_43396# 3.17e-19
C10100 a_n357_42282# a_n447_43370# 0.00435f
C10101 a_6171_45002# a_11909_44484# 3.97e-20
C10102 a_22223_45036# a_18114_32519# 0.15655f
C10103 a_11827_44484# a_19721_31679# 6.72e-20
C10104 a_17339_46660# a_18817_42826# 3.49e-19
C10105 a_n2956_39768# a_5934_30871# 6.35e-21
C10106 a_1423_45028# a_8375_44464# 0.032906f
C10107 a_13507_46334# a_13258_32519# 0.049541f
C10108 a_8199_44636# a_5649_42852# 9.98e-20
C10109 a_9482_43914# a_10617_44484# 1.06e-19
C10110 a_11963_45334# a_n2661_43922# 4.65e-20
C10111 a_n743_46660# a_2277_45546# 8.23e-21
C10112 a_n2661_46098# a_310_45028# 5.46e-20
C10113 a_n133_46660# a_n443_42852# 0.001534f
C10114 a_n2438_43548# a_1609_45822# 0.002001f
C10115 a_n2293_46634# a_509_45572# 3.2e-19
C10116 a_12156_46660# a_10809_44734# 9.31e-19
C10117 a_765_45546# a_10903_43370# 1.58e-19
C10118 a_13059_46348# a_14840_46494# 0.031849f
C10119 a_n1991_46122# a_n1076_46494# 0.124988f
C10120 a_12861_44030# a_16020_45572# 9.09e-21
C10121 a_11599_46634# a_16680_45572# 0.002914f
C10122 a_n2293_46098# a_805_46414# 0.00328f
C10123 a_16327_47482# a_15903_45785# 0.005367f
C10124 a_6755_46942# a_10586_45546# 1.39e-19
C10125 a_4361_42308# a_20107_42308# 0.010379f
C10126 a_4190_30871# a_18997_42308# 6.68e-19
C10127 a_5534_30871# a_6123_31319# 0.01835f
C10128 a_13467_32519# a_20712_42282# 0.003044f
C10129 a_743_42282# a_21613_42308# 1.39e-19
C10130 a_21487_43396# a_21335_42336# 5.61e-19
C10131 a_21855_43396# a_13258_32519# 2.82e-20
C10132 a_5649_42852# a_19511_42282# 1.09e-19
C10133 a_3080_42308# a_n3420_37440# 7.3e-19
C10134 a_6298_44484# a_7845_44172# 0.007037f
C10135 a_n755_45592# a_n2293_42282# 0.208531f
C10136 a_3357_43084# a_7274_43762# 6.44e-21
C10137 a_19778_44110# a_19862_44208# 0.213467f
C10138 a_5147_45002# a_3080_42308# 1.53e-20
C10139 a_5111_44636# a_4699_43561# 9.88e-20
C10140 a_11691_44458# a_13483_43940# 7.11e-21
C10141 a_18494_42460# a_15493_43396# 7.22e-20
C10142 a_n863_45724# a_873_42968# 0.002982f
C10143 a_4842_47570# DATA[2] 1.24e-19
C10144 a_n1059_45260# a_7287_43370# 8.2e-20
C10145 a_n913_45002# a_6547_43396# 1.48e-20
C10146 a_11827_44484# a_17973_43940# 0.004848f
C10147 a_4842_47243# VDD 6.34e-20
C10148 a_5883_43914# a_6453_43914# 0.051468f
C10149 a_18184_42460# a_19478_44306# 7.63e-21
C10150 a_8049_45260# a_10586_45546# 0.038262f
C10151 a_1823_45246# a_4880_45572# 0.002594f
C10152 a_13059_46348# a_16115_45572# 1.11e-20
C10153 a_15227_44166# a_18341_45572# 0.017357f
C10154 a_18834_46812# a_18909_45814# 9e-22
C10155 a_6086_46660# a_3357_43084# 3.67e-19
C10156 a_13507_46334# a_20193_45348# 0.253904f
C10157 a_n2293_46634# a_2809_45348# 0.001204f
C10158 a_5204_45822# a_6194_45824# 4.22e-20
C10159 a_4817_46660# a_3537_45260# 4.15e-22
C10160 a_19466_46812# a_18175_45572# 7.28e-19
C10161 a_11415_45002# a_13249_42308# 0.071546f
C10162 a_3877_44458# a_5111_44636# 3.05e-20
C10163 a_4646_46812# a_5147_45002# 0.010619f
C10164 a_3699_46348# a_3775_45552# 1.45e-19
C10165 a_n746_45260# a_7_44811# 0.001383f
C10166 a_8016_46348# a_2711_45572# 0.028247f
C10167 a_15051_42282# a_15764_42576# 0.042737f
C10168 a_14113_42308# a_15803_42450# 0.289859f
C10169 a_5534_30871# EN_VIN_BSTR_P 0.007335f
C10170 a_685_42968# VDD 0.088446f
C10171 a_n3674_37592# a_n4209_39304# 5.44e-20
C10172 a_3065_45002# a_4149_42891# 4.76e-19
C10173 a_895_43940# a_726_44056# 8.79e-19
C10174 a_2479_44172# a_1241_43940# 7.25e-20
C10175 a_20820_30879# EN_OFFSET_CAL 0.107181f
C10176 a_5111_44636# a_6101_43172# 2.6e-20
C10177 a_1414_42308# a_2455_43940# 1.52e-20
C10178 a_10729_43914# a_10949_43914# 0.418928f
C10179 a_10405_44172# a_10807_43548# 0.004649f
C10180 a_20193_45348# a_21855_43396# 0.001332f
C10181 a_11823_42460# a_11633_42558# 0.039752f
C10182 a_18287_44626# a_10341_43396# 2.54e-20
C10183 a_10193_42453# a_14113_42308# 0.007003f
C10184 a_n2293_42834# a_8605_42826# 1.62e-19
C10185 a_n1991_46122# VDD 0.581018f
C10186 a_6598_45938# a_6469_45572# 4.2e-19
C10187 a_6667_45809# a_6905_45572# 0.001705f
C10188 a_6472_45840# a_8336_45822# 2.77e-20
C10189 a_6511_45714# a_6977_45572# 0.001881f
C10190 a_10809_44734# a_6171_45002# 0.244599f
C10191 a_526_44458# a_413_45260# 0.103799f
C10192 a_11415_45002# a_17613_45144# 0.004987f
C10193 a_16375_45002# a_17668_45572# 2.56e-19
C10194 a_16327_47482# a_18451_43940# 0.001635f
C10195 a_10227_46804# a_15682_43940# 0.003864f
C10196 a_12861_44030# a_21115_43940# 0.035299f
C10197 a_13925_46122# a_14797_45144# 1.91e-20
C10198 a_6945_45028# a_5205_44484# 0.058545f
C10199 a_2711_45572# a_11682_45822# 0.006243f
C10200 a_3483_46348# a_5837_45028# 0.00532f
C10201 a_4185_45028# a_5009_45028# 0.002751f
C10202 a_21588_30879# a_17730_32519# 0.05582f
C10203 a_768_44030# a_2479_44172# 0.056833f
C10204 a_14840_46494# a_13556_45296# 2.96e-19
C10205 a_2324_44458# a_9482_43914# 0.009807f
C10206 a_n1613_43370# a_7281_43914# 0.030229f
C10207 a_n881_46662# a_6453_43914# 2.61e-19
C10208 a_8049_45260# a_21297_45572# 2.09e-19
C10209 a_3090_45724# a_14539_43914# 0.040638f
C10210 a_376_46348# a_n2661_43370# 1.86e-21
C10211 a_9049_44484# a_10180_45724# 3.43e-20
C10212 a_8568_45546# a_8746_45002# 1.75e-19
C10213 a_7499_43078# a_10193_42453# 0.298293f
C10214 a_n4064_37984# a_n2216_37984# 0.005565f
C10215 a_14113_42308# VDD 0.365578f
C10216 a_n2497_47436# a_n1925_46634# 0.052533f
C10217 a_n2288_47178# a_n2312_38680# 4.65e-20
C10218 a_17591_47464# a_12465_44636# 0.001005f
C10219 a_19386_47436# a_20990_47178# 1.56e-20
C10220 a_n3565_39304# a_n2302_37690# 4.02e-19
C10221 a_2112_39137# VDAC_Ni 0.018166f
C10222 SMPL_ON_P a_n2472_46634# 2.91e-19
C10223 a_n2109_47186# a_n2104_46634# 0.009799f
C10224 a_n1741_47186# a_n2442_46660# 0.014004f
C10225 a_n1605_47204# a_n2661_46634# 0.006062f
C10226 a_4915_47217# a_11117_47542# 0.003021f
C10227 a_16327_47482# a_11453_44696# 0.038815f
C10228 a_6151_47436# a_8128_46384# 0.052868f
C10229 a_4958_30871# C6_P_btm 0.005441f
C10230 a_7227_47204# a_n881_46662# 0.001451f
C10231 a_18479_47436# a_21496_47436# 4.29e-19
C10232 a_18780_47178# a_13507_46334# 3.23e-20
C10233 a_18079_43940# a_16823_43084# 5.17e-20
C10234 a_2998_44172# a_3681_42891# 6.9e-21
C10235 a_20835_44721# a_20922_43172# 1.53e-20
C10236 a_20640_44752# a_21195_42852# 2.95e-22
C10237 a_19279_43940# a_19164_43230# 7.21e-21
C10238 a_20679_44626# a_21356_42826# 1.01e-20
C10239 en_comp a_n2302_38778# 1.86e-19
C10240 a_n2956_37592# a_n2860_38778# 3.22e-20
C10241 a_7499_43078# VDD 1.87959f
C10242 a_11750_44172# a_743_42282# 8.68e-22
C10243 a_742_44458# a_2123_42473# 9.65e-21
C10244 a_9313_44734# a_13814_43218# 1.02e-19
C10245 a_11341_43940# a_19268_43646# 5.82e-20
C10246 a_15493_43940# a_18783_43370# 1.32e-19
C10247 a_1209_43370# a_1427_43646# 0.08213f
C10248 a_1049_43396# a_n1557_42282# 0.211757f
C10249 a_n447_43370# a_n144_43396# 0.001377f
C10250 a_4093_43548# a_3080_42308# 0.08049f
C10251 a_4235_43370# a_4699_43561# 0.007134f
C10252 a_4646_46812# a_4093_43548# 3.43e-21
C10253 a_16375_45002# a_17970_44736# 0.00591f
C10254 a_8746_45002# a_n2661_43370# 0.052623f
C10255 a_10193_42453# a_11915_45394# 0.001156f
C10256 a_18597_46090# a_4361_42308# 0.024928f
C10257 a_3357_43084# a_20447_31679# 3.48e-19
C10258 a_4791_45118# a_4520_42826# 1.52e-19
C10259 a_n2293_46634# a_7274_43762# 1.42e-19
C10260 a_15227_44166# a_14485_44260# 4.39e-21
C10261 a_13259_45724# a_18443_44721# 0.004991f
C10262 a_17715_44484# a_19006_44850# 1.14e-20
C10263 a_22591_45572# a_22959_45572# 7.52e-19
C10264 a_13661_43548# a_14205_43396# 2.89e-19
C10265 a_8270_45546# a_9801_43940# 0.014887f
C10266 a_n356_45724# a_n2661_44458# 8.5e-21
C10267 a_n755_45592# a_n1352_44484# 1.52e-20
C10268 a_n863_45724# a_n699_43396# 0.23135f
C10269 a_15903_45785# a_14537_43396# 9.9e-21
C10270 a_8696_44636# a_13159_45002# 7.18e-20
C10271 a_13747_46662# a_11735_46660# 2.58e-21
C10272 a_5807_45002# a_11901_46660# 0.003131f
C10273 a_3785_47178# a_1823_45246# 4.37e-19
C10274 C4_P_btm VREF 0.98728f
C10275 a_13507_46334# a_18285_46348# 0.041986f
C10276 a_4883_46098# a_765_45546# 0.055532f
C10277 a_20894_47436# a_20107_46660# 3.26e-20
C10278 a_10227_46804# a_22000_46634# 5.39e-19
C10279 C5_P_btm VREF_GND 0.676559f
C10280 C6_P_btm VCM 0.877162f
C10281 a_3221_46660# a_3877_44458# 1.36e-19
C10282 a_n1741_47186# a_8953_45546# 2.11e-19
C10283 a_n237_47217# a_6165_46155# 0.021223f
C10284 a_n443_46116# a_472_46348# 0.025699f
C10285 a_13717_47436# a_22591_46660# 4.57e-19
C10286 a_12861_44030# a_11415_45002# 0.081894f
C10287 a_2609_46660# a_3633_46660# 2.36e-20
C10288 a_n743_46660# a_6755_46942# 0.044888f
C10289 a_2063_45854# a_3483_46348# 0.164542f
C10290 a_2905_45572# a_2698_46116# 2.3e-20
C10291 a_n1151_42308# a_167_45260# 8.02e-20
C10292 a_3160_47472# a_2521_46116# 1.93e-19
C10293 a_12549_44172# a_15559_46634# 0.012304f
C10294 a_768_44030# a_15368_46634# 6.08e-22
C10295 C2_P_btm VIN_P 0.502408f
C10296 a_2107_46812# a_8667_46634# 1.72e-19
C10297 C8_N_btm VDD 0.19922f
C10298 a_10695_43548# a_10341_42308# 1.31e-19
C10299 a_3422_30871# a_7174_31319# 2.22059f
C10300 a_4905_42826# a_5193_43172# 0.00336f
C10301 a_8685_43396# a_14543_43071# 4.35e-20
C10302 a_743_42282# a_4361_42308# 7.66647f
C10303 a_4190_30871# a_13678_32519# 0.032285f
C10304 a_21259_43561# a_5649_42852# 1.29e-20
C10305 a_n1925_42282# a_104_43370# 4.1e-21
C10306 a_2324_44458# a_6031_43396# 2.16e-20
C10307 a_n443_42852# a_13483_43940# 2.18e-20
C10308 a_n913_45002# a_n356_44636# 0.640597f
C10309 a_7276_45260# a_6298_44484# 0.007535f
C10310 a_8696_44636# a_11967_42832# 9.33e-19
C10311 a_12741_44636# a_18783_43370# 4.28e-21
C10312 a_3090_45724# a_7871_42858# 1.56e-20
C10313 a_n357_42282# a_20935_43940# 2.76e-19
C10314 a_3483_46348# a_14955_43396# 1.76e-19
C10315 a_4185_45028# a_14205_43396# 4.43e-21
C10316 a_6171_45002# a_5883_43914# 0.002503f
C10317 a_3232_43370# a_9838_44484# 0.053106f
C10318 a_8199_44636# a_8685_43396# 0.03394f
C10319 a_3357_43084# a_5891_43370# 0.013053f
C10320 a_n2293_45010# a_n1243_44484# 3.45e-19
C10321 a_2609_46660# a_526_44458# 2.13e-19
C10322 a_2107_46812# a_6640_46482# 8.98e-19
C10323 a_7715_46873# a_2324_44458# 2.47e-20
C10324 a_3090_45724# a_1823_45246# 0.038665f
C10325 a_14180_46812# a_11415_45002# 8.77e-22
C10326 a_20107_46660# a_20411_46873# 0.316529f
C10327 a_19551_46910# a_20273_46660# 2.93e-19
C10328 a_19123_46287# a_20841_46902# 3.69e-21
C10329 a_6755_46942# a_11189_46129# 6.12e-20
C10330 a_10249_46116# a_11133_46155# 0.007085f
C10331 a_n1151_42308# a_12791_45546# 1.07e-20
C10332 a_6151_47436# a_10053_45546# 2.75e-22
C10333 a_4915_47217# a_8746_45002# 9.87e-21
C10334 a_n743_46660# a_8049_45260# 2.07544f
C10335 a_10623_46897# a_10903_43370# 1.59e-19
C10336 a_4190_30871# a_6123_31319# 0.018095f
C10337 a_15781_43660# a_15803_42450# 1.76e-20
C10338 a_16137_43396# a_14113_42308# 2.26e-19
C10339 a_685_42968# a_n784_42308# 9.99e-21
C10340 a_10341_43396# a_17124_42282# 9.69e-21
C10341 a_16795_42852# a_17141_43172# 0.013377f
C10342 a_743_42282# a_6761_42308# 0.01018f
C10343 a_4361_42308# a_5755_42308# 0.010214f
C10344 a_5649_42852# a_4921_42308# 0.133152f
C10345 a_3600_43914# VDD 0.22716f
C10346 a_15227_44166# a_15803_42450# 0.006356f
C10347 a_8975_43940# a_12189_44484# 6.54e-20
C10348 a_5129_47502# VDD 0.20906f
C10349 a_20193_45348# a_20637_44484# 4.36e-19
C10350 a_11827_44484# a_22591_44484# 0.003361f
C10351 a_3785_47178# DATA[2] 0.119025f
C10352 a_4915_47217# RST_Z 5.15e-19
C10353 a_11823_42460# a_12281_43396# 0.049968f
C10354 a_n356_44636# a_556_44484# 0.001314f
C10355 a_n357_42282# a_n1641_43230# 2.03e-19
C10356 a_10903_43370# a_13291_42460# 0.135558f
C10357 SMPL_ON_N a_22821_38993# 2.28e-19
C10358 a_2274_45254# a_2253_43940# 2.55e-20
C10359 a_14539_43914# a_14815_43914# 0.099149f
C10360 a_15004_44636# a_15146_44811# 0.005572f
C10361 a_n1151_42308# DATA[4] 8.05e-22
C10362 a_10193_42453# a_15781_43660# 5.82e-21
C10363 a_4185_45028# a_22400_42852# 0.105692f
C10364 a_1307_43914# a_15682_43940# 0.028719f
C10365 a_15009_46634# a_11823_42460# 2.01e-21
C10366 a_4915_47217# a_14403_45348# 1.22e-19
C10367 a_768_44030# a_2680_45002# 0.028861f
C10368 a_n2293_46098# a_n2810_45572# 0.013787f
C10369 a_n2472_46090# a_n2661_45546# 0.00558f
C10370 a_11453_44696# a_14537_43396# 0.029591f
C10371 a_n2956_38680# a_n1736_46482# 1.43e-19
C10372 a_9823_46155# a_10044_46482# 0.007833f
C10373 a_8016_46348# a_10037_46155# 0.002633f
C10374 a_20202_43084# a_n357_42282# 0.062522f
C10375 a_15227_44166# a_10193_42453# 0.205591f
C10376 a_n2956_39768# a_n2661_45010# 1.22e-20
C10377 a_n133_46660# a_2437_43646# 3.38e-21
C10378 a_n881_46662# a_6171_45002# 0.090566f
C10379 a_n1613_43370# a_6431_45366# 0.006556f
C10380 a_n2956_39304# a_n1545_46494# 1.4e-20
C10381 a_11189_46129# a_8049_45260# 0.03932f
C10382 a_8953_45546# a_10586_45546# 2.02e-20
C10383 a_4190_30871# EN_VIN_BSTR_P 0.043599f
C10384 a_1606_42308# a_11323_42473# 1.34e-20
C10385 a_15781_43660# VDD 0.196099f
C10386 a_14209_32519# a_22469_39537# 1.36e-20
C10387 a_5755_42308# a_6761_42308# 2.13e-19
C10388 a_10341_43396# CLK 4.37e-20
C10389 a_9313_44734# a_10651_43940# 2.96e-19
C10390 a_18287_44626# a_n97_42460# 2.47e-20
C10391 a_15227_44166# VDD 2.69945f
C10392 a_17609_46634# START 4.81e-19
C10393 a_3537_45260# a_3935_42891# 0.001584f
C10394 a_n913_45002# a_12379_42858# 0.066604f
C10395 a_n2017_45002# a_12545_42858# 1.03e-19
C10396 a_n1059_45260# a_12089_42308# 0.022942f
C10397 a_n2956_39304# a_n2946_39072# 0.150476f
C10398 a_n2956_38680# a_n3420_39072# 0.001161f
C10399 a_3905_42865# a_5013_44260# 0.182997f
C10400 a_18579_44172# a_15682_43940# 1.06e-20
C10401 a_12991_46634# CLK 5.91e-20
C10402 a_n443_42852# a_6123_31319# 6.89e-19
C10403 a_11967_42832# a_20365_43914# 7.55e-20
C10404 a_n2661_42834# a_5326_44056# 2.01e-19
C10405 a_20159_44458# a_19862_44208# 8.53e-20
C10406 a_n699_43396# a_3540_43646# 7.76e-19
C10407 a_7499_43078# a_n784_42308# 6.51e-20
C10408 a_20202_43084# CAL_N 0.002046f
C10409 a_11309_47204# a_11541_44484# 3.58e-22
C10410 a_n881_46662# a_14673_44172# 1.47e-19
C10411 a_n755_45592# a_3775_45552# 0.100709f
C10412 a_22612_30879# a_9313_44734# 1.86e-20
C10413 a_10809_44734# a_18909_45814# 3.61e-23
C10414 a_1823_45246# a_2274_45254# 0.255985f
C10415 a_9290_44172# a_3357_43084# 5.59e-22
C10416 a_18479_47436# a_21073_44484# 5.66e-19
C10417 a_13259_45724# a_13249_42308# 0.358931f
C10418 a_14383_46116# a_14495_45572# 6.09e-19
C10419 a_n2293_46634# a_5891_43370# 0.105307f
C10420 a_167_45260# a_327_44734# 0.199136f
C10421 a_8049_45260# a_11136_45572# 8.45e-20
C10422 a_11415_45002# a_11787_45002# 0.072246f
C10423 a_5742_30871# VDAC_N 0.00823f
C10424 a_n3565_39590# a_n3420_38528# 0.031237f
C10425 a_14097_32519# VREF 2.43e-19
C10426 a_1736_39587# a_1736_39043# 1.92825f
C10427 a_1239_39587# comp_n 0.001233f
C10428 a_n4334_39392# a_n4064_39072# 0.410653f
C10429 a_n4209_39304# a_n2302_39072# 0.407162f
C10430 a_n4209_39590# a_n4064_38528# 0.032071f
C10431 a_n1329_42308# VDD 0.237697f
C10432 a_n784_42308# C8_N_btm 6.79e-20
C10433 a_1606_42308# C0_P_btm 0.029189f
C10434 a_2905_45572# a_n1435_47204# 5.63e-19
C10435 a_5815_47464# a_6545_47178# 0.001457f
C10436 a_4915_47217# a_6851_47204# 0.172567f
C10437 a_n1151_42308# a_11459_47204# 3.65e-19
C10438 a_5129_47502# a_6491_46660# 1.6e-20
C10439 a_n3690_39392# a_n3420_39072# 0.414961f
C10440 a_n3565_39304# a_n2946_39072# 0.410957f
C10441 a_n4064_39616# a_n4209_38502# 0.02801f
C10442 a_n3420_39616# a_n3565_38502# 0.028014f
C10443 COMP_P RST_Z 0.034203f
C10444 a_15493_43940# a_3626_43646# 3.83e-20
C10445 a_n2017_45002# a_19332_42282# 1.65e-19
C10446 a_n1059_45260# a_18907_42674# 0.001868f
C10447 a_n913_45002# a_18727_42674# 2.28e-19
C10448 a_n2661_43922# a_8952_43230# 6.16e-22
C10449 a_n2661_42834# a_10083_42826# 2.3e-20
C10450 a_n2293_43922# a_9127_43156# 6.49e-20
C10451 en_comp a_4958_30871# 0.086457f
C10452 a_20205_31679# C10_N_btm 2.25e-20
C10453 a_20692_30879# C9_N_btm 1.64e-19
C10454 a_375_42282# a_6123_31319# 1.31e-20
C10455 a_1307_43914# a_5934_30871# 3.28e-21
C10456 a_18184_42460# a_20256_43172# 0.043416f
C10457 a_9313_44734# a_12895_43230# 0.007885f
C10458 a_3422_30871# a_21487_43396# 0.003721f
C10459 a_20679_44626# a_20749_43396# 1.57e-21
C10460 a_2107_46812# a_9165_43940# 1.02e-19
C10461 a_17957_46116# a_18287_44626# 2.68e-21
C10462 a_18819_46122# a_18248_44752# 2.46e-21
C10463 a_17715_44484# a_18374_44850# 6.22e-20
C10464 a_6812_45938# a_5205_44484# 4.18e-20
C10465 a_16147_45260# a_18175_45572# 0.108647f
C10466 a_17339_46660# a_20512_43084# 1.02e-19
C10467 a_21588_30879# a_17538_32519# 0.055813f
C10468 a_2711_45572# a_16019_45002# 0.024255f
C10469 a_10809_44734# a_12607_44458# 0.0024f
C10470 a_526_44458# a_2779_44458# 0.090804f
C10471 a_n1613_43370# a_n1557_42282# 1.85e-19
C10472 a_13259_45724# a_17613_45144# 0.002217f
C10473 a_8199_44636# a_8783_44734# 0.00224f
C10474 a_16375_45002# a_16501_45348# 0.00327f
C10475 a_8568_45546# a_3232_43370# 4.2e-21
C10476 a_8162_45546# a_6171_45002# 0.008027f
C10477 a_3147_46376# a_n2661_43922# 3.32e-21
C10478 a_3483_46348# a_n2661_42834# 0.0234f
C10479 a_n3690_37440# VDD 0.363068f
C10480 a_4883_46098# a_10623_46897# 1.58e-19
C10481 a_n2661_46634# a_n133_46660# 0.022138f
C10482 a_n2472_46634# a_n2438_43548# 0.008762f
C10483 VDAC_P C1_P_btm 0.560533f
C10484 a_n881_46662# a_4955_46873# 0.066882f
C10485 a_n1435_47204# a_12816_46660# 7.47e-21
C10486 a_n1613_43370# a_4817_46660# 0.330391f
C10487 CAL_P a_11530_34132# 0.055606f
C10488 a_11599_46634# a_11735_46660# 0.268769f
C10489 a_n2293_46634# a_n1021_46688# 2.69e-22
C10490 a_n2104_46634# a_n1925_46634# 0.167849f
C10491 a_n1151_42308# a_12925_46660# 5.47e-20
C10492 a_768_44030# a_2864_46660# 1.39e-19
C10493 a_10341_43396# a_19268_43646# 0.010402f
C10494 a_n97_42460# a_9127_43156# 1.6e-19
C10495 a_3422_30871# a_5932_42308# 0.022048f
C10496 a_453_43940# a_1184_42692# 2.56e-21
C10497 a_4558_45348# VDD 0.25277f
C10498 a_n4318_39768# a_n4318_38216# 0.023318f
C10499 a_413_45260# DATA[5] 0.0381f
C10500 a_15681_43442# a_16243_43396# 6.39e-21
C10501 a_15781_43660# a_16137_43396# 0.089942f
C10502 a_3232_43370# a_n2661_43370# 0.077167f
C10503 a_n357_42282# a_n809_44244# 0.001553f
C10504 a_6171_45002# a_11361_45348# 8.73e-20
C10505 a_15227_44166# a_16137_43396# 0.002078f
C10506 a_n1613_43370# a_8483_43230# 5.99e-19
C10507 a_7276_45260# a_7418_45067# 0.005572f
C10508 a_8953_45002# a_n2293_42834# 1.18e-19
C10509 a_n863_45724# a_1467_44172# 0.021736f
C10510 a_13059_46348# a_13667_43396# 0.00451f
C10511 a_16327_47482# a_19273_43230# 9.01e-20
C10512 a_2107_46812# a_5204_45822# 0.002125f
C10513 a_n2293_46634# a_9290_44172# 0.102393f
C10514 a_584_46384# a_n755_45592# 0.020619f
C10515 a_2063_45854# a_n357_42282# 1.15e-20
C10516 a_3699_46634# a_1823_45246# 1.1e-20
C10517 a_n2661_46098# a_2804_46116# 1.71e-20
C10518 a_12861_44030# a_13259_45724# 0.435853f
C10519 a_12816_46660# a_13885_46660# 8.55e-20
C10520 a_n2661_46634# a_11387_46155# 0.0013f
C10521 a_1431_47204# a_1848_45724# 2.87e-19
C10522 a_n971_45724# a_7_45899# 3.69e-19
C10523 a_19333_46634# a_19692_46634# 0.005582f
C10524 a_n1613_43370# a_n722_46482# 0.002104f
C10525 a_n881_46662# a_n967_46494# 8.68e-20
C10526 a_n1151_42308# a_n863_45724# 0.081395f
C10527 a_2609_46660# a_2521_46116# 1.95e-19
C10528 a_2443_46660# a_2698_46116# 9.84e-20
C10529 a_n743_46660# a_8953_45546# 0.062066f
C10530 a_12891_46348# a_6945_45028# 0.013255f
C10531 a_13747_46662# a_2324_44458# 0.025909f
C10532 a_13661_43548# a_15682_46116# 1.42e-19
C10533 a_5807_45002# a_17583_46090# 0.008151f
C10534 a_15743_43084# a_20753_42852# 1.06e-19
C10535 a_17730_32519# a_22469_39537# 1.95e-20
C10536 a_3626_43646# a_5742_30871# 0.168508f
C10537 a_5649_42852# a_13291_42460# 5.5e-20
C10538 a_9396_43370# a_5934_30871# 4.98e-19
C10539 a_n97_42460# a_17124_42282# 5.78e-20
C10540 a_5111_44636# a_5244_44056# 0.01138f
C10541 a_4927_45028# a_3905_42865# 1.58e-19
C10542 a_3537_45260# a_6453_43914# 6.46e-19
C10543 a_10903_43370# a_13460_43230# 3.23e-19
C10544 a_n357_42282# a_14955_43396# 6.56e-20
C10545 a_n443_42852# a_6809_43396# 5.25e-19
C10546 a_n2661_44458# a_n356_44636# 0.055568f
C10547 a_526_44458# a_n13_43084# 2.42e-19
C10548 a_n1925_42282# a_n1076_43230# 1.95e-20
C10549 a_9290_44172# a_5342_30871# 6.73e-19
C10550 a_10334_44484# a_10440_44484# 0.313533f
C10551 a_9838_44484# a_8975_43940# 0.055678f
C10552 a_10157_44484# a_10057_43914# 6.36e-19
C10553 a_n1699_44726# a_n1809_44850# 0.097745f
C10554 a_n1917_44484# a_n2012_44484# 0.049827f
C10555 a_n2267_44484# a_n1190_44850# 1.46e-19
C10556 a_5147_45002# a_5013_44260# 0.189328f
C10557 a_3232_43370# a_2998_44172# 0.056614f
C10558 a_20623_45572# a_19862_44208# 7.47e-20
C10559 a_11827_44484# a_9313_44734# 1.07e-19
C10560 a_21588_30879# a_22465_38105# 7.99e-19
C10561 a_n2312_38680# a_7174_31319# 3.87e-21
C10562 a_4185_45028# a_22223_42860# 2.62e-20
C10563 a_20990_47178# a_3357_43084# 1.67e-19
C10564 a_4883_46098# a_21513_45002# 0.005388f
C10565 a_n2157_46122# a_n967_46494# 2.56e-19
C10566 a_n1641_46494# a_n2956_38680# 2.13e-19
C10567 a_4646_46812# a_7499_43078# 0.158236f
C10568 a_n1151_42308# a_8191_45002# 7.92e-19
C10569 a_14513_46634# a_14383_46116# 4.21e-20
C10570 a_14180_46812# a_13259_45724# 1.49e-21
C10571 a_21496_47436# a_2437_43646# 0.01965f
C10572 a_13507_46334# a_22223_45572# 0.015966f
C10573 a_16327_47482# a_n1059_45260# 0.235708f
C10574 a_10428_46928# a_2711_45572# 4.68e-20
C10575 a_5257_43370# a_7227_45028# 7.21e-21
C10576 a_13381_47204# a_413_45260# 1.38e-19
C10577 a_n881_46662# a_18909_45814# 1.16e-20
C10578 a_15227_44166# a_20850_46155# 8.44e-19
C10579 a_4791_45118# a_6431_45366# 1.75e-20
C10580 a_12549_44172# a_14033_45572# 2.6e-19
C10581 a_768_44030# a_13485_45572# 9.77e-20
C10582 a_20841_46902# a_8049_45260# 8.01e-21
C10583 a_13747_46662# a_16855_45546# 0.02676f
C10584 a_5807_45002# a_8696_44636# 0.024228f
C10585 a_3483_46348# a_17715_44484# 0.059106f
C10586 a_4419_46090# a_2324_44458# 2.42e-20
C10587 a_9625_46129# a_9290_44172# 4.14e-20
C10588 a_n1991_46122# a_n1545_46494# 2.28e-19
C10589 a_21671_42860# a_17303_42282# 3.64e-20
C10590 a_n4318_37592# a_n3674_37592# 3.06402f
C10591 a_n3674_38216# a_n1630_35242# 0.333493f
C10592 a_19164_43230# a_19332_42282# 0.002067f
C10593 a_n1329_42308# a_n784_42308# 9.6e-19
C10594 a_3080_42308# C8_N_btm 0.006767f
C10595 a_1756_43548# VDD 0.138878f
C10596 a_18579_44172# a_20512_43084# 3.29e-19
C10597 a_n2810_45572# a_n1736_42282# 2.3e-20
C10598 a_3686_47026# VDD 4.6e-19
C10599 a_22223_45036# a_14401_32519# 3.29e-20
C10600 a_11827_44484# a_20974_43370# 2.22e-20
C10601 a_3363_44484# a_3499_42826# 1.97e-20
C10602 a_n2661_42834# a_261_44278# 3.83e-19
C10603 a_21398_44850# a_3422_30871# 2.52e-19
C10604 a_13556_45296# a_13667_43396# 1.26e-20
C10605 a_14537_43396# a_9145_43396# 0.129182f
C10606 a_n357_42282# a_19326_42852# 1.44e-19
C10607 a_18248_44752# a_11341_43940# 6.59e-20
C10608 a_n2293_42834# a_3626_43646# 0.019674f
C10609 a_19279_43940# a_17730_32519# 1.25e-20
C10610 a_5891_43370# a_9672_43914# 0.009207f
C10611 a_n2956_38216# a_n4318_38216# 0.023519f
C10612 a_7499_43078# a_7309_43172# 0.001045f
C10613 a_768_44030# a_5518_44484# 0.00362f
C10614 a_20273_46660# a_3357_43084# 0.02704f
C10615 a_4651_46660# a_n2661_43370# 1.49e-21
C10616 a_21588_30879# a_19721_31679# 0.055771f
C10617 a_22612_30879# a_18114_32519# 0.061298f
C10618 a_3090_45724# a_6709_45028# 1.32e-20
C10619 a_11415_45002# a_18787_45572# 7.51e-19
C10620 a_21363_46634# a_2437_43646# 2.82e-19
C10621 a_3483_46348# a_15861_45028# 2.64e-19
C10622 a_10809_44734# a_8746_45002# 0.049227f
C10623 a_5066_45546# a_6472_45840# 2.68e-19
C10624 a_n1630_35242# a_8530_39574# 7.09e-20
C10625 a_n2497_47436# a_n2288_47178# 0.067981f
C10626 a_n2833_47464# a_n2109_47186# 0.002667f
C10627 a_6123_31319# a_n3420_37984# 0.00363f
C10628 a_13258_32519# a_21613_42308# 0.060546f
C10629 a_n3674_37592# a_n4334_37440# 0.050036f
C10630 a_22400_42852# a_22469_40625# 0.954861f
C10631 a_4223_44672# a_8037_42858# 9.39e-19
C10632 a_11967_42832# a_14205_43396# 1.68e-19
C10633 a_n1059_45260# a_5267_42460# 6.15e-20
C10634 a_n2017_45002# a_5379_42460# 0.003023f
C10635 a_n913_45002# a_3823_42558# 0.029622f
C10636 a_n2810_45572# a_n4209_37414# 3.74e-21
C10637 a_22959_46124# VDD 0.309939f
C10638 a_3905_42865# a_4699_43561# 0.001039f
C10639 a_10809_44734# RST_Z 0.00392f
C10640 a_6945_45028# SINGLE_ENDED 0.021393f
C10641 a_11827_44484# a_18599_43230# 5.4e-21
C10642 a_1307_43914# a_16245_42852# 1.03e-20
C10643 a_14673_44172# a_14621_43646# 6.57e-20
C10644 a_1414_42308# a_2982_43646# 0.071994f
C10645 a_18184_42460# a_21195_42852# 0.017258f
C10646 a_5891_43370# a_743_42282# 0.065685f
C10647 a_13661_43548# a_20269_44172# 0.001724f
C10648 a_768_44030# a_9895_44260# 9.29e-19
C10649 a_18819_46122# a_16922_45042# 9.18e-21
C10650 a_n755_45592# a_n659_45366# 4.7e-19
C10651 a_12741_44636# a_17767_44458# 2.58e-19
C10652 a_n2293_46634# a_10807_43548# 0.05087f
C10653 a_13747_46662# a_19862_44208# 0.15289f
C10654 a_1823_45246# a_4743_44484# 0.001634f
C10655 a_5204_45822# a_n2661_44458# 5e-21
C10656 a_n1099_45572# a_n143_45144# 8.04e-20
C10657 a_11415_45002# a_18287_44626# 9.88e-20
C10658 a_n2661_45546# a_3065_45002# 0.004264f
C10659 a_19321_45002# a_15493_43396# 1.18e-20
C10660 a_3090_45724# a_15146_44484# 7.43e-20
C10661 a_n971_45724# a_8147_43396# 0.116186f
C10662 a_584_46384# a_548_43396# 7.2e-19
C10663 a_n2293_45546# a_2274_45254# 0.07158f
C10664 a_n863_45724# a_327_44734# 0.353745f
C10665 a_12594_46348# a_11827_44484# 5.74e-21
C10666 a_17715_44484# a_17719_45144# 0.009296f
C10667 a_7754_40130# CAL_P 0.04831f
C10668 a_n237_47217# a_8492_46660# 0.002629f
C10669 a_n1741_47186# a_10249_46116# 5.18e-19
C10670 a_n1435_47204# a_2443_46660# 5.41e-20
C10671 a_4915_47217# a_4651_46660# 1.15e-19
C10672 a_5129_47502# a_4646_46812# 1.7e-20
C10673 a_5815_47464# a_3877_44458# 2.22e-20
C10674 a_n4334_39392# VDD 0.385989f
C10675 a_22223_47212# a_21588_30879# 0.164932f
C10676 a_12465_44636# a_22612_30879# 7.45e-19
C10677 a_n3420_38528# C4_P_btm 0.030945f
C10678 a_n4064_38528# C6_P_btm 0.001467f
C10679 a_n3420_37984# EN_VIN_BSTR_P 0.031779f
C10680 a_n443_46116# a_4955_46873# 0.126551f
C10681 a_4791_45118# a_4817_46660# 0.020367f
C10682 a_n1151_42308# a_5072_46660# 0.009494f
C10683 a_2905_45572# a_3633_46660# 3.11e-19
C10684 a_2063_45854# a_5263_46660# 1.33e-19
C10685 VDAC_Ni a_6886_37412# 0.178275f
C10686 a_7754_38636# VDAC_N 9.38e-20
C10687 a_n4209_39590# VREF_GND 0.083908f
C10688 a_n3420_37440# a_n4064_37440# 8.19012f
C10689 a_3754_38470# a_5088_37509# 0.632585f
C10690 a_7754_38470# a_3726_37500# 0.124796f
C10691 a_n4209_37414# a_n4251_37440# 0.00226f
C10692 a_n3565_37414# a_n2860_37690# 2.96e-19
C10693 a_22731_47423# a_20916_46384# 1.06e-19
C10694 a_n2293_43922# a_1755_42282# 1.6e-19
C10695 a_20193_45348# a_21613_42308# 0.137559f
C10696 a_8147_43396# a_8229_43396# 0.005781f
C10697 a_n97_42460# a_19268_43646# 0.002543f
C10698 a_n356_44636# a_8325_42308# 1.57e-19
C10699 a_2982_43646# a_12281_43396# 4.32e-19
C10700 a_5891_43370# a_5755_42308# 7.45e-19
C10701 a_12429_44172# a_5534_30871# 3.45e-20
C10702 a_22612_30879# a_13887_32519# 0.060052f
C10703 a_526_44458# a_644_44056# 3.05e-19
C10704 a_n2661_45010# a_1307_43914# 0.016415f
C10705 a_n1059_45260# a_14537_43396# 2.86e-21
C10706 a_5147_45002# a_4927_45028# 0.168157f
C10707 a_8746_45002# a_5883_43914# 2.04e-20
C10708 a_10180_45724# a_10157_44484# 0.001525f
C10709 a_n357_42282# a_n2661_42834# 0.239713f
C10710 a_4558_45348# a_5691_45260# 1.08e-19
C10711 a_9290_44172# a_9672_43914# 0.071844f
C10712 a_16327_47482# a_19987_42826# 0.053812f
C10713 a_3537_45260# a_6171_45002# 4.04e-19
C10714 a_4574_45260# a_3232_43370# 3.36e-21
C10715 a_8696_44636# a_18315_45260# 4.09e-21
C10716 a_15861_45028# a_17719_45144# 0.002134f
C10717 a_17478_45572# a_17613_45144# 3.37e-20
C10718 a_15037_45618# a_11827_44484# 3.23e-22
C10719 a_310_45028# a_n2661_43922# 2.83e-19
C10720 a_7499_43078# a_10057_43914# 0.262644f
C10721 a_3316_45546# a_3363_44484# 3.64e-20
C10722 a_2905_45572# a_526_44458# 0.142766f
C10723 a_3160_47472# a_2981_46116# 4.76e-19
C10724 a_12861_44030# a_18189_46348# 0.004513f
C10725 a_7903_47542# a_6945_45028# 0.005336f
C10726 a_n881_46662# a_376_46348# 0.016146f
C10727 a_n1613_43370# a_472_46348# 3.32e-19
C10728 a_4883_46098# a_8349_46414# 0.007204f
C10729 a_11599_46634# a_2324_44458# 0.428445f
C10730 a_n237_47217# a_5210_46155# 0.002744f
C10731 a_8492_46660# a_8270_45546# 0.007406f
C10732 a_10227_46804# a_10903_43370# 0.041882f
C10733 a_n133_46660# a_765_45546# 7.71e-20
C10734 a_584_46384# a_835_46155# 0.001103f
C10735 a_18451_43940# a_18727_42674# 1.72e-21
C10736 a_4190_30871# a_18083_42858# 0.023338f
C10737 a_8685_43396# a_13291_42460# 2.12e-19
C10738 a_14021_43940# a_14113_42308# 3.15e-20
C10739 a_n2293_43922# VDAC_P 6.46e-20
C10740 a_743_42282# a_17595_43084# 5.58e-20
C10741 a_13467_32519# a_5342_30871# 0.028573f
C10742 a_9838_44484# VDD 0.242131f
C10743 a_n1557_42282# a_n1736_42282# 0.170341f
C10744 a_n97_42460# a_1755_42282# 0.002698f
C10745 a_n357_42282# a_n1352_43396# 2.09e-19
C10746 a_n755_45592# a_n1177_43370# 3.74e-19
C10747 a_n2661_43370# a_8975_43940# 3.05e-19
C10748 a_3232_43370# a_11909_44484# 2.99e-20
C10749 a_11827_44484# a_18114_32519# 0.09907f
C10750 a_21359_45002# a_19721_31679# 2.35e-20
C10751 a_3357_43084# a_22315_44484# 1.44e-21
C10752 a_9290_44172# a_743_42282# 0.117511f
C10753 a_8953_45546# a_4361_42308# 0.012234f
C10754 a_17339_46660# a_18249_42858# 0.008924f
C10755 a_11322_45546# a_11173_44260# 2.01e-20
C10756 SMPL_ON_P a_n3420_37984# 6.62e-21
C10757 a_13507_46334# a_19647_42308# 5.23e-19
C10758 a_1423_45028# a_7640_43914# 0.105665f
C10759 a_11963_45334# a_n2661_42834# 9.32e-20
C10760 a_11787_45002# a_n2661_43922# 2.24e-20
C10761 a_16327_47482# a_15599_45572# 0.331892f
C10762 a_n2661_46098# a_n1099_45572# 7.03e-20
C10763 a_n2438_43548# a_n443_42852# 3.03e-19
C10764 a_n743_46660# a_1609_45822# 5.99e-19
C10765 a_n2293_46634# a_n89_45572# 4.13e-19
C10766 a_15227_46910# a_14840_46494# 2e-19
C10767 a_13059_46348# a_15015_46420# 0.002269f
C10768 a_n1853_46287# a_n1076_46494# 0.056078f
C10769 a_n1991_46122# a_n901_46420# 0.041816f
C10770 a_12861_44030# a_17478_45572# 3.55e-19
C10771 a_11599_46634# a_16855_45546# 0.002089f
C10772 a_2107_46812# a_3503_45724# 7.75e-22
C10773 a_n2293_46098# a_472_46348# 0.009446f
C10774 a_n2157_46122# a_376_46348# 2.25e-21
C10775 a_n2109_47186# a_3357_43084# 0.170493f
C10776 a_n1423_46090# a_n1641_46494# 0.209641f
C10777 a_10249_46116# a_10586_45546# 1.88e-19
C10778 a_5807_45002# a_7227_45028# 6.28e-20
C10779 a_13467_32519# a_20107_42308# 0.001069f
C10780 a_4361_42308# a_13258_32519# 0.076336f
C10781 a_n2293_42282# a_2351_42308# 6.05e-19
C10782 a_17538_32519# a_22469_39537# 1.77e-20
C10783 a_10083_42826# a_9885_42558# 0.001558f
C10784 a_n881_46662# RST_Z 0.351994f
C10785 a_6298_44484# a_7542_44172# 0.014735f
C10786 a_n1809_44850# a_n1761_44111# 7.57e-20
C10787 a_8696_44636# a_16867_43762# 1.57e-19
C10788 a_n357_42282# a_n2293_42282# 0.01064f
C10789 a_16922_45042# a_11341_43940# 0.028038f
C10790 a_14815_43914# a_15146_44484# 2.88e-19
C10791 a_11691_44458# a_12429_44172# 2.31e-20
C10792 a_18184_42460# a_15493_43396# 7.78e-20
C10793 a_n863_45724# a_133_42852# 1.03e-19
C10794 a_n2017_45002# a_7287_43370# 1.12e-20
C10795 a_11827_44484# a_17737_43940# 0.003402f
C10796 a_5883_43914# a_5663_43940# 0.153361f
C10797 a_3232_43370# a_1568_43370# 7.3e-19
C10798 a_19778_44110# a_19478_44306# 0.099524f
C10799 a_8049_45260# a_8379_46155# 1.85e-19
C10800 a_13059_46348# a_16333_45814# 3.56e-20
C10801 a_15227_44166# a_18479_45785# 0.035756f
C10802 a_5841_46660# a_3357_43084# 1.99e-19
C10803 a_13507_46334# a_11691_44458# 3.47e-20
C10804 a_17715_44484# a_n357_42282# 1.41e-20
C10805 a_n2438_43548# a_375_42282# 2.84e-20
C10806 a_n2293_46634# a_2304_45348# 0.00666f
C10807 a_5164_46348# a_6194_45824# 4.82e-20
C10808 a_5497_46414# a_5263_45724# 3.95e-21
C10809 a_12465_44636# a_11827_44484# 0.785011f
C10810 a_19466_46812# a_16147_45260# 3.68e-21
C10811 a_3877_44458# a_5147_45002# 1.31e-20
C10812 a_4646_46812# a_4558_45348# 7.53e-22
C10813 a_3483_46348# a_3775_45552# 3.9e-20
C10814 a_n746_45260# a_n310_44811# 0.002132f
C10815 a_7920_46348# a_2711_45572# 0.001215f
C10816 a_15051_42282# a_15486_42560# 0.234322f
C10817 a_14113_42308# a_15764_42576# 0.229529f
C10818 a_5534_30871# a_n923_35174# 0.007036f
C10819 a_5932_42308# a_7174_31319# 13.0265f
C10820 a_421_43172# VDD 1.56e-19
C10821 a_20193_45348# a_4361_42308# 7.54e-19
C10822 a_n2293_42834# a_8037_42858# 0.009778f
C10823 a_11823_42460# a_11551_42558# 0.138126f
C10824 a_453_43940# a_1443_43940# 0.009173f
C10825 a_n2661_42834# a_n144_43396# 2.02e-19
C10826 a_5111_44636# a_5837_43172# 1.31e-19
C10827 a_1414_42308# a_2253_43940# 1.35e-19
C10828 a_22591_46660# EN_OFFSET_CAL 0.047938f
C10829 a_10405_44172# a_10949_43914# 0.05348f
C10830 a_9672_43914# a_10807_43548# 2.13e-20
C10831 a_11415_45002# CLK 6.94e-20
C10832 a_18579_44172# a_21381_43940# 1.29e-21
C10833 a_n1853_46287# VDD 0.645231f
C10834 a_n913_45002# a_12800_43218# 0.016338f
C10835 a_10193_42453# a_13657_42558# 0.009218f
C10836 a_18248_44752# a_10341_43396# 3.47e-20
C10837 a_3537_45260# a_8292_43218# 1.01e-19
C10838 a_10903_43370# a_1307_43914# 0.065094f
C10839 a_6472_45840# a_6977_45572# 2.28e-19
C10840 a_10809_44734# a_3232_43370# 0.158726f
C10841 a_6945_45028# a_6431_45366# 0.00135f
C10842 a_2981_46116# a_413_45260# 0.002451f
C10843 a_16327_47482# a_18326_43940# 2.74e-20
C10844 a_10227_46804# a_14955_43940# 0.004814f
C10845 a_12861_44030# a_20935_43940# 0.02414f
C10846 a_13759_46122# a_14797_45144# 2.6e-20
C10847 a_14493_46090# a_14180_45002# 6.1e-20
C10848 a_13925_46122# a_14537_43396# 6.19e-21
C10849 a_2711_45572# a_11280_45822# 1.69e-19
C10850 a_3483_46348# a_5093_45028# 0.05597f
C10851 a_768_44030# a_2127_44172# 0.002861f
C10852 a_11415_45002# a_17023_45118# 0.004458f
C10853 a_14840_46494# a_9482_43914# 6.56e-21
C10854 a_2324_44458# a_13348_45260# 0.005924f
C10855 a_15015_46420# a_13556_45296# 2.21e-20
C10856 a_n1613_43370# a_6453_43914# 0.007952f
C10857 a_8049_45260# a_20447_31679# 0.009404f
C10858 a_14976_45028# a_15004_44636# 0.001535f
C10859 a_9049_44484# a_10053_45546# 0.005221f
C10860 a_13657_42558# VDD 0.195727f
C10861 a_n2497_47436# a_n2312_38680# 3.06e-19
C10862 a_16588_47582# a_12465_44636# 1.91e-19
C10863 a_n3565_39304# a_n4064_37440# 0.028266f
C10864 a_n4064_39072# a_n3565_37414# 0.031386f
C10865 a_n3420_39072# a_n3420_37440# 0.052876f
C10866 a_n4064_37984# a_n2860_37984# 0.003765f
C10867 a_22465_38105# a_22469_39537# 0.576946f
C10868 a_n2288_47178# a_n2104_46634# 3.21e-19
C10869 SMPL_ON_P a_n2661_46634# 0.0112f
C10870 a_n2109_47186# a_n2293_46634# 3.45e-19
C10871 a_n1920_47178# a_n2442_46660# 0.00281f
C10872 a_n1605_47204# a_n2956_39768# 2.5e-19
C10873 a_4915_47217# a_10037_47542# 1.22e-19
C10874 a_n3420_39616# VDAC_P 0.004488f
C10875 a_4958_30871# C7_P_btm 1.47e-19
C10876 a_7227_47204# a_n1613_43370# 2.15e-20
C10877 a_6851_47204# a_n881_46662# 0.002875f
C10878 a_18479_47436# a_13507_46334# 0.033523f
C10879 a_10227_46804# a_4883_46098# 0.200137f
C10880 a_2998_44172# a_2905_42968# 3.82e-19
C10881 a_3905_42865# a_1847_42826# 2.52e-20
C10882 a_18579_44172# a_18249_42858# 1.81e-20
C10883 a_20640_44752# a_21356_42826# 7.48e-22
C10884 a_19279_43940# a_19339_43156# 3.69e-21
C10885 a_n2956_37592# a_n2302_38778# 0.006499f
C10886 en_comp a_n4064_38528# 2.01e-21
C10887 a_8568_45546# VDD 0.182812f
C10888 a_n1441_43940# a_n1641_43230# 5.44e-21
C10889 a_10807_43548# a_743_42282# 0.011093f
C10890 a_3422_30871# a_15567_42826# 5.99e-21
C10891 a_742_44458# a_1755_42282# 0.013027f
C10892 a_9313_44734# a_13569_43230# 1.23e-19
C10893 a_14021_43940# a_15781_43660# 0.00563f
C10894 a_17973_43940# a_16823_43084# 1.54e-20
C10895 a_n699_43396# a_961_42354# 1.36e-21
C10896 a_11341_43940# a_15743_43084# 6.7e-19
C10897 a_15493_43940# a_18525_43370# 1.15e-19
C10898 a_1049_43396# a_766_43646# 6.4e-21
C10899 a_4093_43548# a_4699_43561# 7.24e-19
C10900 a_1209_43370# a_n1557_42282# 0.113851f
C10901 a_16375_45002# a_17767_44458# 0.00258f
C10902 a_10193_42453# a_n2661_43370# 3.69e-19
C10903 a_18597_46090# a_13467_32519# 0.002694f
C10904 a_1823_45246# a_1414_42308# 0.002939f
C10905 a_n2293_46098# a_6453_43914# 0.002061f
C10906 a_1138_42852# a_453_43940# 0.018298f
C10907 a_19479_31679# a_20447_31679# 0.05179f
C10908 a_n2293_46634# a_5837_43396# 1.35e-19
C10909 a_15227_44166# a_14021_43940# 0.052407f
C10910 a_13259_45724# a_18287_44626# 0.002131f
C10911 a_8049_45260# a_5891_43370# 0.00367f
C10912 a_n1925_42282# a_n2293_43922# 2.06056f
C10913 a_17715_44484# a_18588_44850# 4.47e-20
C10914 a_13507_46334# a_4190_30871# 0.186424f
C10915 a_10227_46804# a_5649_42852# 2.58e-19
C10916 a_3357_43084# a_22959_45572# 8.46e-19
C10917 a_22591_45572# a_19963_31679# 0.161955f
C10918 a_5807_45002# a_14205_43396# 9.38e-20
C10919 a_13661_43548# a_14358_43442# 1.8e-19
C10920 a_8270_45546# a_9420_43940# 0.007316f
C10921 a_2711_45572# a_11827_44484# 0.033351f
C10922 a_8696_44636# a_13017_45260# 1.73e-20
C10923 a_15599_45572# a_14537_43396# 3.89e-19
C10924 a_n755_45592# a_n1177_44458# 1.63e-19
C10925 a_3503_45724# a_n2661_44458# 4.06e-21
C10926 a_2107_46812# a_7927_46660# 5.88e-20
C10927 a_n1925_46634# a_6969_46634# 0.007338f
C10928 a_n2661_46634# a_8035_47026# 0.002111f
C10929 a_5807_45002# a_11813_46116# 0.037525f
C10930 a_n1151_42308# a_2202_46116# 1.13e-21
C10931 a_3381_47502# a_1823_45246# 1.03e-19
C10932 C5_P_btm VREF 0.987144f
C10933 a_11453_44696# a_16721_46634# 4.18e-21
C10934 a_4883_46098# a_17339_46660# 0.071433f
C10935 a_13507_46334# a_17829_46910# 8.95e-19
C10936 a_10227_46804# a_21188_46660# 0.22222f
C10937 C7_P_btm VCM 1.58335f
C10938 C6_P_btm VREF_GND 0.836236f
C10939 a_3055_46660# a_3877_44458# 2.12e-19
C10940 a_n237_47217# a_5497_46414# 0.021428f
C10941 a_n971_45724# a_6419_46155# 0.001374f
C10942 a_n1741_47186# a_5937_45572# 4.26e-20
C10943 a_n443_46116# a_376_46348# 0.025241f
C10944 a_13717_47436# a_11415_45002# 4.62e-20
C10945 a_12861_44030# a_20202_43084# 0.020377f
C10946 C9_N_btm C10_N_btm 37.815998f
C10947 a_18597_46090# a_20273_46660# 3.9e-19
C10948 a_2443_46660# a_3633_46660# 2.56e-19
C10949 a_n743_46660# a_10249_46116# 0.004613f
C10950 a_2063_45854# a_3147_46376# 0.005517f
C10951 a_584_46384# a_3483_46348# 0.00258f
C10952 a_3160_47472# a_167_45260# 2.66e-19
C10953 a_12549_44172# a_15368_46634# 0.012256f
C10954 C3_P_btm VIN_P 0.455045f
C10955 a_18479_47436# a_20623_46660# 0.005343f
C10956 C7_N_btm VDD 0.121904f
C10957 a_12465_44636# a_14447_46660# 1.13e-19
C10958 a_19721_31679# a_22469_39537# 3.67e-20
C10959 a_3422_30871# a_20712_42282# 0.016384f
C10960 a_n2661_43370# VDD 1.53673f
C10961 a_9145_43396# a_12379_42858# 0.001164f
C10962 a_4905_42826# a_4743_43172# 2.86e-19
C10963 a_8685_43396# a_13460_43230# 4.34e-20
C10964 a_743_42282# a_13467_32519# 0.003709f
C10965 a_n1925_42282# a_n97_42460# 0.021883f
C10966 a_8191_45002# a_4223_44672# 1.76e-20
C10967 a_n443_42852# a_12429_44172# 1.23e-19
C10968 a_n1059_45260# a_n356_44636# 0.07487f
C10969 a_n1613_43370# a_n3674_37592# 8.6e-20
C10970 a_5205_44484# a_6298_44484# 0.085118f
C10971 a_3090_45724# a_7227_42852# 3.82e-19
C10972 a_n357_42282# a_20623_43914# 1.2e-20
C10973 a_3483_46348# a_15095_43370# 1.36e-21
C10974 a_11415_45002# a_19268_43646# 2.56e-21
C10975 en_comp a_n2012_44484# 4.42e-20
C10976 a_7229_43940# a_5343_44458# 0.196399f
C10977 a_3232_43370# a_5883_43914# 0.337937f
C10978 a_10467_46802# a_10903_43370# 8.89e-21
C10979 a_6151_47436# a_9049_44484# 3.15e-20
C10980 a_11901_46660# a_3483_46348# 4.96e-21
C10981 a_2443_46660# a_526_44458# 3.42e-19
C10982 a_2609_46660# a_2981_46116# 0.001665f
C10983 a_14035_46660# a_11415_45002# 3.1e-21
C10984 a_19551_46910# a_20411_46873# 6.03e-20
C10985 a_19123_46287# a_20273_46660# 7.53e-20
C10986 a_16388_46812# a_18280_46660# 3.41e-20
C10987 a_4817_46660# a_6945_45028# 8.99e-21
C10988 a_2107_46812# a_6419_46482# 5.65e-19
C10989 a_7411_46660# a_2324_44458# 1.67e-21
C10990 a_6755_46942# a_9290_44172# 3.62e-19
C10991 a_10249_46116# a_11189_46129# 1.33e-19
C10992 a_n1151_42308# a_11823_42460# 9.67e-20
C10993 a_4915_47217# a_10193_42453# 1.89e-20
C10994 a_15681_43442# a_15803_42450# 3.32e-19
C10995 a_15781_43660# a_15764_42576# 3.57e-20
C10996 a_421_43172# a_n784_42308# 5.98e-21
C10997 a_16795_42852# a_16877_43172# 0.003935f
C10998 a_743_42282# a_6773_42558# 0.001159f
C10999 a_4361_42308# a_5421_42558# 7.13e-20
C11000 a_2998_44172# VDD 0.362233f
C11001 a_15227_44166# a_15764_42576# 0.003122f
C11002 a_8975_43940# a_11909_44484# 2.14e-19
C11003 a_4915_47217# VDD 3.43172f
C11004 a_n1151_42308# DATA[3] 5.14e-19
C11005 a_6109_44484# a_7640_43914# 0.002099f
C11006 a_3381_47502# DATA[2] 1.73e-19
C11007 a_413_45260# a_3052_44056# 4.96e-19
C11008 a_n913_45002# a_8487_44056# 1.53e-20
C11009 a_n2661_43370# a_5495_43940# 2.51e-21
C11010 a_11827_44484# a_22485_44484# 0.015798f
C11011 a_n357_42282# a_n1423_42826# 5.7e-19
C11012 a_10903_43370# a_13003_42852# 0.006128f
C11013 SMPL_ON_N a_22545_38993# 1.95e-21
C11014 a_526_44458# a_4156_43218# 2.93e-19
C11015 a_19929_45028# a_18579_44172# 6.24e-19
C11016 a_1307_43914# a_14955_43940# 0.00962f
C11017 a_16019_45002# a_15682_43940# 0.001434f
C11018 a_5937_45572# a_10586_45546# 1.5e-19
C11019 a_4915_47217# a_14309_45348# 0.002491f
C11020 a_768_44030# a_2382_45260# 0.094536f
C11021 a_4883_46098# a_1307_43914# 0.026965f
C11022 a_n2840_46090# a_n2661_45546# 0.003502f
C11023 a_n2293_46098# a_n2840_45546# 0.004047f
C11024 a_11453_44696# a_14180_45002# 0.005785f
C11025 a_n2956_39304# a_n1736_46482# 1.91e-20
C11026 a_8016_46348# a_9751_46155# 0.001112f
C11027 a_12816_46660# a_13163_45724# 1.14e-19
C11028 a_n2438_43548# a_2437_43646# 0.045715f
C11029 a_n1925_46634# a_3357_43084# 0.034378f
C11030 a_n881_46662# a_3232_43370# 0.001015f
C11031 a_9290_44172# a_8049_45260# 0.041148f
C11032 a_n1613_43370# a_6171_45002# 0.026867f
C11033 a_17364_32525# a_22521_39511# 9.72e-21
C11034 a_4190_30871# a_n923_35174# 0.025255f
C11035 a_4921_42308# a_6123_31319# 2.25e-19
C11036 a_1606_42308# a_10723_42308# 3.31e-20
C11037 a_6171_42473# a_6481_42558# 6.01e-20
C11038 a_15681_43442# VDD 0.159054f
C11039 a_9313_44734# a_10555_43940# 0.001497f
C11040 a_18248_44752# a_n97_42460# 1.22e-20
C11041 a_19615_44636# a_19862_44208# 8.86e-19
C11042 a_18834_46812# VDD 0.116625f
C11043 a_n1331_43914# a_n822_43940# 2.6e-19
C11044 a_3537_45260# a_3681_42891# 3.51e-19
C11045 a_n913_45002# a_10341_42308# 0.070067f
C11046 a_n1059_45260# a_12379_42858# 0.003827f
C11047 a_n2017_45002# a_12089_42308# 0.043278f
C11048 a_n863_45724# a_5742_30871# 2.35e-20
C11049 a_n2956_39304# a_n3420_39072# 0.208204f
C11050 a_13259_45724# a_17124_42282# 0.003167f
C11051 a_19279_43940# a_17973_43940# 5.98e-20
C11052 a_n443_42852# a_7227_42308# 8.04e-21
C11053 a_16922_45042# a_10341_43396# 0.048996f
C11054 a_11967_42832# a_20269_44172# 4.03e-20
C11055 a_n2661_42834# a_5025_43940# 1.83e-19
C11056 a_20820_30879# VDAC_N 4.55e-19
C11057 a_1307_43914# a_5649_42852# 2.47e-20
C11058 a_3905_42865# a_5244_44056# 0.002415f
C11059 a_n699_43396# a_2982_43646# 0.004394f
C11060 a_n2293_46098# a_6171_45002# 2.23e-21
C11061 a_n971_45724# a_n2661_42282# 3.65e-19
C11062 a_1823_45246# a_1667_45002# 0.24808f
C11063 a_21588_30879# a_9313_44734# 1.69e-20
C11064 a_10809_44734# a_18341_45572# 6.97e-21
C11065 a_4185_45028# en_comp 0.001836f
C11066 a_13259_45724# a_13904_45546# 0.007639f
C11067 a_14383_46116# a_13249_42308# 7.26e-20
C11068 a_n2293_46634# a_8375_44464# 1.16e-21
C11069 a_167_45260# a_413_45260# 0.120357f
C11070 a_11133_46155# a_2437_43646# 3.61e-22
C11071 a_5742_30871# a_6886_37412# 3.23e-19
C11072 a_14097_32519# VIN_N 0.053964f
C11073 a_1736_39587# a_1239_39043# 0.036194f
C11074 a_n4209_39304# a_n4064_39072# 0.19711f
C11075 COMP_P VDD 3.48893f
C11076 a_n784_42308# C7_N_btm 0.002308f
C11077 a_2952_47436# a_n1435_47204# 2.1e-19
C11078 a_5815_47464# a_6151_47436# 0.235454f
C11079 a_4915_47217# a_6491_46660# 0.19739f
C11080 a_n1151_42308# a_9313_45822# 0.024431f
C11081 a_5129_47502# a_6545_47178# 1.1e-19
C11082 a_4791_45118# a_7227_47204# 6.26e-19
C11083 a_n3565_39304# a_n3420_39072# 0.241179f
C11084 a_n3420_39616# a_n4334_38528# 4.91e-19
C11085 a_1606_42308# C1_P_btm 0.096405f
C11086 a_1307_43914# a_7963_42308# 3.36e-21
C11087 a_n1059_45260# a_18727_42674# 0.20226f
C11088 a_n2017_45002# a_18907_42674# 6.48e-20
C11089 a_n913_45002# a_18057_42282# 1.34e-19
C11090 a_18579_44172# a_5649_42852# 1.35e-22
C11091 a_n2661_43922# a_9127_43156# 2.21e-20
C11092 a_n2661_42834# a_8952_43230# 9.54e-21
C11093 a_n2293_43922# a_8387_43230# 9.06e-21
C11094 a_20447_31679# a_13258_32519# 0.054935f
C11095 a_20205_31679# C9_N_btm 1.91e-20
C11096 a_20692_30879# C8_N_btm 1.15e-19
C11097 a_18184_42460# a_18707_42852# 3.84e-20
C11098 a_9313_44734# a_13113_42826# 0.004011f
C11099 a_8162_45546# a_3232_43370# 8.68e-20
C11100 a_7230_45938# a_6171_45002# 0.001502f
C11101 a_2277_45546# a_2304_45348# 7.72e-19
C11102 a_17957_46116# a_18248_44752# 6.35e-20
C11103 a_18189_46348# a_18287_44626# 1.01e-19
C11104 a_17715_44484# a_18443_44721# 3.58e-20
C11105 a_13259_45724# a_17023_45118# 1.58e-19
C11106 a_8953_45546# a_5891_43370# 0.321625f
C11107 a_10227_46804# a_8685_43396# 0.227547f
C11108 w_11334_34010# a_13467_32519# 3.26e-19
C11109 a_22612_30879# a_14401_32519# 0.062739f
C11110 a_2711_45572# a_15595_45028# 7.51e-20
C11111 a_2981_46116# a_2779_44458# 2e-21
C11112 a_526_44458# a_949_44458# 0.03455f
C11113 a_n863_45724# a_n2293_42834# 0.107229f
C11114 a_n1925_42282# a_742_44458# 1.15e-20
C11115 a_10586_45546# a_11691_44458# 1e-20
C11116 a_12861_44030# a_14955_43396# 0.024664f
C11117 a_10809_44734# a_8975_43940# 0.169586f
C11118 a_16375_45002# a_16405_45348# 0.012425f
C11119 a_8199_44636# a_8333_44734# 0.002302f
C11120 a_4883_46098# a_9396_43370# 0.172323f
C11121 a_n3565_37414# VDD 0.783539f
C11122 a_4883_46098# a_10467_46802# 7.03e-19
C11123 a_n2661_46634# a_n2438_43548# 0.493975f
C11124 VDAC_P C2_P_btm 1.03235f
C11125 a_n1435_47204# a_12991_46634# 6.91e-20
C11126 a_n1613_43370# a_4955_46873# 0.051259f
C11127 a_11599_46634# a_11186_47026# 1.68e-20
C11128 a_n2104_46634# a_n2312_38680# 0.154937f
C11129 a_n2293_46634# a_n1925_46634# 0.051324f
C11130 a_n2442_46660# a_n1021_46688# 2.1e-20
C11131 a_n1151_42308# a_12513_46660# 1.2e-19
C11132 a_n881_46662# a_4651_46660# 1.63e-19
C11133 a_4574_45260# VDD 0.122256f
C11134 a_10341_43396# a_15743_43084# 0.464206f
C11135 a_n97_42460# a_8387_43230# 2.28e-20
C11136 a_1568_43370# a_2905_42968# 5.03e-21
C11137 a_n3674_39768# a_n3674_38680# 0.035445f
C11138 a_9396_43370# a_5649_42852# 6.62e-21
C11139 a_453_43940# a_1576_42282# 3.54e-21
C11140 a_413_45260# DATA[4] 0.037695f
C11141 a_1414_42308# a_1184_42692# 0.115223f
C11142 a_15681_43442# a_16137_43396# 2.85e-19
C11143 a_n863_45724# a_1115_44172# 0.008873f
C11144 a_n2661_45546# a_2479_44172# 6.41e-21
C11145 a_10903_43370# a_10867_43940# 0.004161f
C11146 a_5691_45260# a_n2661_43370# 0.015295f
C11147 a_8696_44636# a_18374_44850# 9.12e-20
C11148 a_n1613_43370# a_8292_43218# 0.011565f
C11149 a_7229_43940# a_8560_45348# 1.25e-19
C11150 a_380_45546# a_175_44278# 5.93e-21
C11151 a_n913_45002# a_18494_42460# 4.44e-19
C11152 a_11823_42460# a_13857_44734# 9.1e-21
C11153 a_8191_45002# a_n2293_42834# 0.084957f
C11154 a_10193_42453# a_11909_44484# 3.99e-20
C11155 a_n1151_42308# a_961_42354# 2.65e-22
C11156 a_16327_47482# a_18861_43218# 0.004178f
C11157 a_2107_46812# a_5164_46348# 0.002137f
C11158 a_584_46384# a_n357_42282# 0.107436f
C11159 a_n2661_46098# a_2698_46116# 3.89e-20
C11160 a_4007_47204# a_n2661_45546# 2.2e-21
C11161 a_13717_47436# a_13259_45724# 2.52e-20
C11162 a_12861_44030# a_14383_46116# 1.08e-19
C11163 a_12469_46902# a_14180_46812# 4.58e-22
C11164 a_4883_46098# a_8034_45724# 0.004608f
C11165 a_11599_46634# a_12839_46116# 0.042002f
C11166 a_n2109_47186# a_2277_45546# 3e-21
C11167 a_n746_45260# a_n23_45546# 0.004336f
C11168 a_n237_47217# a_n356_45724# 1.25e-20
C11169 a_n971_45724# a_n310_45899# 0.002723f
C11170 a_4955_46873# a_n2293_46098# 0.002285f
C11171 a_n1151_42308# a_n1079_45724# 0.012662f
C11172 a_15227_44166# a_19692_46634# 0.116169f
C11173 a_19333_46634# a_19466_46812# 0.167526f
C11174 a_n1613_43370# a_n967_46494# 2.95e-19
C11175 a_11309_47204# a_6945_45028# 0.010402f
C11176 a_2443_46660# a_2521_46116# 5.25e-19
C11177 a_n743_46660# a_5937_45572# 0.02494f
C11178 a_5807_45002# a_15682_46116# 0.062679f
C11179 a_13661_43548# a_2324_44458# 0.307974f
C11180 a_12549_44172# a_20708_46348# 1.12e-20
C11181 a_5342_30871# a_16795_42852# 2.89e-20
C11182 a_15567_42826# a_16414_43172# 0.001784f
C11183 a_19319_43548# a_20107_42308# 1.44e-20
C11184 a_3626_43646# a_11323_42473# 0.003176f
C11185 a_2982_43646# a_11551_42558# 1.36e-19
C11186 a_n2661_43922# CLK 1.98e-19
C11187 a_8147_43396# a_8515_42308# 6.85e-19
C11188 a_8791_43396# a_5934_30871# 5.94e-19
C11189 a_n97_42460# a_16522_42674# 2.08e-19
C11190 a_19237_31679# a_22521_39511# 1.89e-20
C11191 a_5111_44636# a_3905_42865# 0.006261f
C11192 a_5147_45002# a_5244_44056# 0.122327f
C11193 a_3537_45260# a_5663_43940# 1.06e-19
C11194 a_n2312_39304# a_n2302_38778# 5.35e-19
C11195 a_n913_45002# a_3499_42826# 6.51e-19
C11196 a_n357_42282# a_15095_43370# 0.034944f
C11197 a_n443_42852# a_6643_43396# 9.4e-19
C11198 a_n2433_44484# a_n1821_44484# 0.001881f
C11199 a_n1925_42282# a_n901_43156# 4.57e-20
C11200 a_5883_43914# a_8975_43940# 0.50976f
C11201 a_n2267_44484# a_n1809_44850# 0.027606f
C11202 a_n2129_44697# a_n1190_44850# 3.86e-19
C11203 a_4558_45348# a_5013_44260# 3.95e-20
C11204 a_4185_45028# a_22165_42308# 6.61e-20
C11205 a_20894_47436# a_3357_43084# 0.002793f
C11206 a_7715_46873# a_6511_45714# 9.45e-19
C11207 a_8016_46348# a_10903_43370# 6.55e-20
C11208 a_n1641_46494# a_n2956_39304# 2.7e-20
C11209 a_n1423_46090# a_n2956_38680# 7.5e-20
C11210 a_n2293_46098# a_n967_46494# 4.35e-20
C11211 a_4646_46812# a_8568_45546# 1.23e-19
C11212 a_n1151_42308# a_7705_45326# 0.042252f
C11213 a_14035_46660# a_13259_45724# 1.96e-19
C11214 a_14180_46812# a_14383_46116# 1.22e-20
C11215 a_13507_46334# a_2437_43646# 0.117533f
C11216 a_16327_47482# a_n2017_45002# 0.209709f
C11217 a_n2497_47436# a_1423_45028# 1.36987f
C11218 a_5257_43370# a_6598_45938# 2.41e-19
C11219 a_10150_46912# a_2711_45572# 1.65e-20
C11220 a_2063_45854# a_11787_45002# 2.33e-20
C11221 a_n1991_46122# a_n1736_46482# 0.06121f
C11222 a_15227_44166# a_20692_30879# 1.69e-19
C11223 a_11459_47204# a_413_45260# 4.35e-19
C11224 a_n881_46662# a_18341_45572# 1.2e-19
C11225 a_4791_45118# a_6171_45002# 0.031317f
C11226 a_n443_46116# a_3232_43370# 0.059286f
C11227 a_12549_44172# a_13485_45572# 0.004173f
C11228 a_20273_46660# a_8049_45260# 2.63e-21
C11229 a_13747_46662# a_16115_45572# 0.029803f
C11230 a_5807_45002# a_16680_45572# 0.006746f
C11231 a_8953_45546# a_9290_44172# 0.373944f
C11232 a_8199_44636# a_11133_46155# 2.47e-20
C11233 a_4185_45028# a_2324_44458# 0.015434f
C11234 a_9625_46129# a_10355_46116# 0.001354f
C11235 a_1568_43370# VDD 0.433732f
C11236 a_21195_42852# a_17303_42282# 3.32e-20
C11237 a_19339_43156# a_19332_42282# 0.004421f
C11238 a_n2104_42282# a_n1630_35242# 0.030917f
C11239 a_n1736_42282# a_n3674_37592# 0.006442f
C11240 COMP_P a_n784_42308# 0.10915f
C11241 a_3080_42308# C7_N_btm 0.002948f
C11242 a_n961_42308# a_n473_42460# 0.011409f
C11243 a_5891_43370# a_9028_43914# 0.001563f
C11244 a_n2956_38216# a_n2472_42282# 2.12e-20
C11245 a_n2810_45572# a_n3674_38216# 0.023322f
C11246 a_21359_45002# a_20974_43370# 5.16e-21
C11247 a_n2661_42834# a_n1441_43940# 0.004368f
C11248 a_n2661_43922# a_n630_44306# 3.27e-19
C11249 a_20679_44626# a_19237_31679# 1.41e-20
C11250 a_9482_43914# a_13667_43396# 1.67e-20
C11251 a_17970_44736# a_11341_43940# 3.63e-21
C11252 a_19279_43940# a_22591_44484# 1.13e-20
C11253 a_16979_44734# a_15493_43940# 6.95e-20
C11254 a_1307_43914# a_8685_43396# 4.34e-20
C11255 a_7499_43078# a_6101_43172# 3.94e-21
C11256 a_19479_31679# a_13467_32519# 0.051245f
C11257 a_2324_44458# a_6229_45572# 3.26e-19
C11258 a_768_44030# a_5343_44458# 0.066821f
C11259 a_12861_44030# a_n2661_42834# 1.42e-20
C11260 a_20411_46873# a_3357_43084# 0.157199f
C11261 a_4646_46812# a_n2661_43370# 0.028718f
C11262 a_n743_46660# a_11691_44458# 5.94e-20
C11263 a_21588_30879# a_18114_32519# 0.055884f
C11264 a_3090_45724# a_7229_43940# 0.054969f
C11265 a_20623_46660# a_2437_43646# 4.3e-20
C11266 a_3483_46348# a_8696_44636# 0.06521f
C11267 a_10903_43370# a_11682_45822# 0.071222f
C11268 a_10809_44734# a_10193_42453# 0.02204f
C11269 a_5066_45546# a_6194_45824# 5.14e-20
C11270 a_n1630_35242# a_7754_38470# 4.78e-20
C11271 a_n2833_47464# a_n2288_47178# 0.003549f
C11272 a_13258_32519# a_21887_42336# 8.1e-19
C11273 a_n3674_37592# a_n4209_37414# 0.044977f
C11274 a_20712_42282# a_7174_31319# 3.53e-19
C11275 a_n4318_37592# a_n2860_37690# 1.77e-20
C11276 a_22400_42852# a_22521_40599# 0.133947f
C11277 a_4223_44672# a_7765_42852# 2.94e-20
C11278 a_11967_42832# a_14358_43442# 8.52e-20
C11279 a_n2017_45002# a_5267_42460# 0.003851f
C11280 a_n913_45002# a_3318_42354# 0.03912f
C11281 a_n1059_45260# a_3823_42558# 2.04e-20
C11282 a_10809_44734# VDD 2.67671f
C11283 a_6945_45028# START 0.029602f
C11284 a_3905_42865# a_4235_43370# 0.041971f
C11285 a_22223_46124# RST_Z 1.13e-19
C11286 a_n2293_42834# a_7309_42852# 4.09e-20
C11287 a_2998_44172# a_3080_42308# 6.67e-19
C11288 a_1414_42308# a_2896_43646# 0.005191f
C11289 a_1467_44172# a_2982_43646# 8.78e-21
C11290 a_18184_42460# a_21356_42826# 0.016504f
C11291 a_5343_44458# a_5755_42852# 5.25e-22
C11292 a_5518_44484# a_5111_42852# 2.49e-21
C11293 a_9313_44734# a_16823_43084# 0.031008f
C11294 a_768_44030# a_9801_44260# 8.82e-19
C11295 a_17957_46116# a_16922_45042# 2.12e-21
C11296 a_n2293_46634# a_10949_43914# 0.001108f
C11297 a_n2661_46634# a_12429_44172# 1.5e-21
C11298 a_13661_43548# a_19862_44208# 2.53e-20
C11299 a_14180_46482# a_14180_45002# 2.55e-21
C11300 a_11189_46129# a_11691_44458# 1.61e-19
C11301 a_5164_46348# a_n2661_44458# 0.001579f
C11302 a_14495_45572# a_8696_44636# 3.04e-20
C11303 a_n1099_45572# a_n467_45028# 0.007609f
C11304 a_11682_45822# a_12016_45572# 2.43e-19
C11305 a_12741_44636# a_16979_44734# 0.008336f
C11306 a_11415_45002# a_18248_44752# 3.19e-20
C11307 a_n2661_45546# a_2680_45002# 0.004432f
C11308 a_n2293_45546# a_1667_45002# 0.07132f
C11309 a_19321_45002# a_19328_44172# 1.77e-19
C11310 a_3877_44458# a_3600_43914# 0.001072f
C11311 a_11823_42460# a_12649_45572# 5.54e-19
C11312 a_11962_45724# a_13297_45572# 0.001004f
C11313 a_12427_45724# a_12749_45572# 0.001367f
C11314 a_n863_45724# a_413_45260# 0.140312f
C11315 a_n755_45592# a_n967_45348# 2.3e-19
C11316 a_1823_45246# a_n699_43396# 0.08003f
C11317 a_17715_44484# a_17613_45144# 0.012898f
C11318 a_13507_46334# a_n2661_46634# 2.61e-20
C11319 a_n1741_47186# a_10554_47026# 1.58e-20
C11320 a_n237_47217# a_8667_46634# 0.171086f
C11321 a_n443_46116# a_4651_46660# 0.060179f
C11322 a_4915_47217# a_4646_46812# 1.43e-19
C11323 a_n4209_39304# VDD 0.984278f
C11324 a_12465_44636# a_21588_30879# 0.053175f
C11325 a_22223_47212# a_20916_46384# 4.95e-19
C11326 a_n3420_38528# C5_P_btm 0.001712f
C11327 a_n4064_38528# C7_P_btm 1.64e-19
C11328 a_n3420_37984# a_n923_35174# 0.002459f
C11329 a_n4209_39590# VREF 0.860047f
C11330 a_n1151_42308# a_6540_46812# 4.39e-20
C11331 a_4791_45118# a_4955_46873# 0.001577f
C11332 a_n1435_47204# a_n2661_46098# 6.55e-20
C11333 a_n3420_37440# a_n2946_37690# 0.236674f
C11334 a_n3690_37440# a_n4064_37440# 0.085414f
C11335 a_n3565_37414# a_n2302_37690# 0.046906f
C11336 a_3754_38470# a_4338_37500# 0.473597f
C11337 VDAC_Ni a_5700_37509# 0.079762f
C11338 a_n4209_37414# a_n2216_37690# 0.001361f
C11339 a_11453_44696# a_19594_46812# 0.041136f
C11340 a_n3565_39590# VIN_P 0.068367f
C11341 en_comp a_22469_40625# 0.021539f
C11342 a_n2293_43922# a_1606_42308# 0.080878f
C11343 a_20193_45348# a_21887_42336# 0.169001f
C11344 a_n97_42460# a_15743_43084# 0.205305f
C11345 a_9396_43370# a_8685_43396# 0.007917f
C11346 a_13483_43940# a_13460_43230# 2.1e-20
C11347 a_20447_31679# a_22609_37990# 9.79e-21
C11348 a_21588_30879# a_13887_32519# 0.056445f
C11349 a_n2017_45002# a_14537_43396# 3.09e-22
C11350 a_5147_45002# a_5111_44636# 0.562127f
C11351 a_4558_45348# a_4927_45028# 0.123258f
C11352 a_4185_45028# a_19862_44208# 1.38e-20
C11353 a_8746_45002# a_8701_44490# 1.65e-19
C11354 a_10053_45546# a_10157_44484# 1.49e-20
C11355 a_19321_45002# a_20749_43396# 2.22e-19
C11356 a_9290_44172# a_9028_43914# 0.169653f
C11357 a_16327_47482# a_19164_43230# 0.292734f
C11358 a_8953_45546# a_10807_43548# 5.44e-21
C11359 a_3537_45260# a_3232_43370# 0.530258f
C11360 a_8049_45260# a_22315_44484# 2.42e-21
C11361 a_8696_44636# a_17719_45144# 3.25e-19
C11362 a_15861_45028# a_17613_45144# 0.016666f
C11363 a_7499_43078# a_10440_44484# 3.35e-19
C11364 a_9049_44484# a_10334_44484# 2.09e-20
C11365 a_n1099_45572# a_n2661_43922# 2.98e-21
C11366 a_7227_47204# a_6945_45028# 0.01947f
C11367 a_12861_44030# a_17715_44484# 3.76e-19
C11368 a_20916_46384# a_20731_47026# 6.18e-20
C11369 a_n881_46662# a_n1076_46494# 0.018649f
C11370 a_n1613_43370# a_376_46348# 4.03e-19
C11371 a_4883_46098# a_8016_46348# 0.289691f
C11372 a_11599_46634# a_14840_46494# 0.051732f
C11373 a_8667_46634# a_8270_45546# 0.046604f
C11374 a_8145_46902# a_8601_46660# 4.2e-19
C11375 a_n743_46660# a_17829_46910# 1.56e-20
C11376 a_2747_46873# a_2804_46116# 0.001759f
C11377 a_16327_47482# a_13759_46122# 1.11e-21
C11378 a_n2438_43548# a_765_45546# 0.081258f
C11379 a_584_46384# a_518_46155# 0.002222f
C11380 a_4190_30871# a_17701_42308# 0.008836f
C11381 a_4361_42308# a_5534_30871# 0.049795f
C11382 a_458_43396# a_564_42282# 1.51e-20
C11383 a_3080_42308# COMP_P 4.43551f
C11384 a_5649_42852# a_13635_43156# 6.61e-20
C11385 a_743_42282# a_16795_42852# 1.32e-20
C11386 a_15493_43396# a_17303_42282# 1.81e-21
C11387 a_5883_43914# VDD 0.859221f
C11388 a_n1557_42282# a_n3674_38216# 1.82e-19
C11389 a_1568_43370# a_n784_42308# 8.96e-20
C11390 a_n97_42460# a_1606_42308# 1.2e-19
C11391 a_n755_45592# a_n1917_43396# 9.06e-20
C11392 a_n357_42282# a_n1177_43370# 7.33e-19
C11393 a_n2661_43370# a_10057_43914# 2.24e-19
C11394 a_3232_43370# a_11541_44484# 0.050289f
C11395 a_21359_45002# a_18114_32519# 2.21e-19
C11396 a_11827_44484# a_20205_45028# 5.4e-19
C11397 a_19479_31679# a_22315_44484# 7.36e-19
C11398 a_3357_43084# a_3422_30871# 1.8e-20
C11399 a_13507_46334# a_19511_42282# 0.004827f
C11400 a_18597_46090# a_21335_42336# 6.48e-21
C11401 en_comp a_11967_42832# 5.02e-20
C11402 a_1423_45028# a_6109_44484# 0.018788f
C11403 a_10951_45334# a_n2661_43922# 4.26e-20
C11404 a_526_44458# a_10341_43396# 0.005028f
C11405 a_n2956_39768# a_6123_31319# 5.77e-21
C11406 a_n743_46660# a_n443_42852# 0.378464f
C11407 a_n2293_46634# a_n310_45572# 1.08e-19
C11408 a_15227_46910# a_15015_46420# 3.17e-20
C11409 a_13059_46348# a_14275_46494# 0.036863f
C11410 a_n1853_46287# a_n901_46420# 0.049679f
C11411 a_n1991_46122# a_n1641_46494# 0.219633f
C11412 a_12861_44030# a_15861_45028# 0.015193f
C11413 a_n1741_47186# a_2437_43646# 4.86702f
C11414 a_11599_46634# a_16115_45572# 8.83e-19
C11415 a_15673_47210# a_15903_45785# 4.56e-21
C11416 a_n1925_46634# a_2277_45546# 1.47e-20
C11417 a_n2293_46098# a_376_46348# 0.004986f
C11418 a_n2157_46122# a_n1076_46494# 0.102355f
C11419 a_n881_46662# a_10193_42453# 6.12e-20
C11420 a_19692_46634# a_22959_46124# 1.54e-19
C11421 a_10554_47026# a_10586_45546# 8.4e-19
C11422 a_5807_45002# a_6598_45938# 0.002355f
C11423 a_n2293_42282# a_2123_42473# 1.62e-19
C11424 a_14635_42282# a_14853_42852# 0.01129f
C11425 a_743_42282# a_21335_42336# 2.86e-19
C11426 a_4361_42308# a_19647_42308# 0.007305f
C11427 a_13467_32519# a_13258_32519# 11.0084f
C11428 a_10341_42308# a_8325_42308# 1.07e-20
C11429 a_n913_45002# a_6197_43396# 2.11e-20
C11430 a_4185_45028# a_9803_42558# 8.71e-20
C11431 a_6298_44484# a_7281_43914# 0.010383f
C11432 a_n1809_44850# a_n2065_43946# 8.2e-20
C11433 a_n357_42282# a_22959_42860# 2.46e-20
C11434 a_3357_43084# a_5565_43396# 0.009914f
C11435 a_9313_44734# a_19279_43940# 3.78e-20
C11436 a_5343_44458# a_7845_44172# 0.103601f
C11437 a_11691_44458# a_11750_44172# 5.84e-19
C11438 a_18184_42460# a_19328_44172# 1.54e-19
C11439 a_19778_44110# a_15493_43396# 0.015561f
C11440 a_n2017_45002# a_6547_43396# 4.02e-20
C11441 a_11827_44484# a_15682_43940# 0.006752f
C11442 a_n881_46662# VDD 2.6692f
C11443 a_5883_43914# a_5495_43940# 0.09813f
C11444 a_4574_45260# a_3080_42308# 5.32e-21
C11445 a_3537_45260# a_4905_42826# 0.339989f
C11446 a_8049_45260# a_8062_46155# 1.21e-20
C11447 a_22959_46124# a_20692_30879# 0.155635f
C11448 a_n746_45260# a_n23_44458# 0.046452f
C11449 a_1823_45246# a_5024_45822# 6.21e-21
C11450 a_4651_46660# a_3537_45260# 4.86e-21
C11451 a_4646_46812# a_4574_45260# 1.08e-20
C11452 a_15227_44166# a_18175_45572# 0.018929f
C11453 a_n743_46660# a_375_42282# 8.64e-21
C11454 a_5164_46348# a_5907_45546# 5.55e-20
C11455 a_5204_45822# a_5263_45724# 0.109078f
C11456 a_13059_46348# a_15765_45572# 1.96e-19
C11457 a_3090_45724# a_18596_45572# 1.73e-19
C11458 a_11453_44696# a_18494_42460# 5.41e-22
C11459 a_19466_46812# a_17786_45822# 9.25e-23
C11460 a_12741_44636# a_11823_42460# 0.031865f
C11461 a_11415_45002# a_13527_45546# 3.65e-20
C11462 a_3877_44458# a_4558_45348# 0.028316f
C11463 a_3483_46348# a_7227_45028# 0.00331f
C11464 a_6419_46155# a_2711_45572# 0.002668f
C11465 a_n2293_46634# a_2232_45348# 8.56e-19
C11466 a_14113_42308# a_15486_42560# 0.039784f
C11467 a_n4318_37592# a_n4064_39072# 0.019896f
C11468 a_6171_42473# a_7174_31319# 4.88e-21
C11469 a_11551_42558# a_11897_42308# 0.013377f
C11470 a_133_43172# VDD 8.22e-19
C11471 a_20193_45348# a_13467_32519# 0.016015f
C11472 a_n2293_42834# a_7765_42852# 0.010796f
C11473 a_11823_42460# a_5742_30871# 9.73e-19
C11474 a_453_43940# a_1241_43940# 0.002487f
C11475 a_n2157_46122# VDD 0.42567f
C11476 a_n2293_43922# a_3539_42460# 6.26e-20
C11477 a_5111_44636# a_5457_43172# 0.002744f
C11478 a_1414_42308# a_1443_43940# 0.018064f
C11479 a_11415_45002# EN_OFFSET_CAL 0.14622f
C11480 a_10405_44172# a_10729_43914# 0.083277f
C11481 a_9672_43914# a_10949_43914# 2.19e-20
C11482 a_18579_44172# a_19741_43940# 0.005651f
C11483 a_19279_43940# a_20974_43370# 2.3e-20
C11484 a_n913_45002# a_10752_42852# 6.19e-19
C11485 a_n1059_45260# a_12800_43218# 0.002165f
C11486 a_3537_45260# a_7573_43172# 1e-19
C11487 a_6511_45714# a_6469_45572# 2.56e-19
C11488 a_6945_45028# a_6171_45002# 0.032875f
C11489 a_8049_45260# a_22959_45572# 0.176374f
C11490 a_17339_46660# a_18545_45144# 2.2e-19
C11491 a_16327_47482# a_18079_43940# 0.001128f
C11492 a_10227_46804# a_13483_43940# 8.62e-19
C11493 a_4915_47217# a_14021_43940# 4.68e-20
C11494 a_12861_44030# a_20623_43914# 0.033132f
C11495 a_13759_46122# a_14537_43396# 1.79e-20
C11496 a_13925_46122# a_14180_45002# 2.26e-20
C11497 a_2711_45572# a_10907_45822# 0.016608f
C11498 a_n357_42282# a_8696_44636# 4.53e-21
C11499 a_3483_46348# a_5009_45028# 0.029292f
C11500 a_11415_45002# a_16922_45042# 0.012903f
C11501 a_768_44030# a_453_43940# 0.110708f
C11502 a_10586_45546# a_2437_43646# 2.49e-20
C11503 a_3090_45724# a_15004_44636# 0.010872f
C11504 a_n901_46420# a_n2661_43370# 2.09e-20
C11505 a_2324_44458# a_13159_45002# 0.00216f
C11506 a_15015_46420# a_9482_43914# 1.28e-20
C11507 a_14275_46494# a_13556_45296# 3.84e-21
C11508 a_16763_47508# a_12465_44636# 8.56e-19
C11509 a_10227_46804# a_21496_47436# 0.007515f
C11510 a_n4209_39304# a_n2302_37690# 3.3e-19
C11511 a_n3420_37984# a_n2216_37984# 5.9e-20
C11512 a_13333_42558# VDD 0.008231f
C11513 a_n2833_47464# a_n2312_38680# 6.08e-20
C11514 a_18597_46090# a_20894_47436# 2.7e-21
C11515 a_19386_47436# a_19787_47423# 0.002814f
C11516 a_n3565_39304# a_n2946_37690# 2.71e-19
C11517 a_n4064_39072# a_n4334_37440# 3.19e-19
C11518 a_n2946_37984# a_n2860_37984# 0.011479f
C11519 a_22465_38105# a_22821_38993# 0.09356f
C11520 a_n2497_47436# a_n2104_46634# 0.002384f
C11521 a_n2109_47186# a_n2442_46660# 0.004864f
C11522 a_n2288_47178# a_n2293_46634# 0.011283f
C11523 a_n1741_47186# a_n2661_46634# 0.22396f
C11524 SMPL_ON_P a_n2956_39768# 0.039986f
C11525 a_4958_30871# C8_P_btm 0.001147f
C11526 a_6851_47204# a_n1613_43370# 2.26e-20
C11527 a_6491_46660# a_n881_46662# 1.53e-19
C11528 a_18479_47436# a_21177_47436# 0.001742f
C11529 a_17591_47464# a_4883_46098# 4.46e-20
C11530 a_4915_47217# a_9804_47204# 0.072476f
C11531 a_2889_44172# a_2905_42968# 5.52e-20
C11532 a_n3674_39768# a_n4318_38680# 0.024755f
C11533 a_n2956_37592# a_n4064_38528# 0.015398f
C11534 a_8162_45546# VDD 0.266272f
C11535 a_3422_30871# a_5342_30871# 0.026613f
C11536 a_742_44458# a_1606_42308# 0.001459f
C11537 a_n2810_45028# a_n2302_38778# 4.97e-19
C11538 a_14021_43940# a_15681_43442# 0.004196f
C11539 a_17737_43940# a_16823_43084# 1.26e-20
C11540 a_11341_43940# a_18783_43370# 3.91e-20
C11541 a_15493_43940# a_18429_43548# 4.75e-20
C11542 a_21115_43940# a_15743_43084# 3.08e-21
C11543 a_n97_42460# a_3539_42460# 0.021726f
C11544 a_458_43396# a_n1557_42282# 0.027865f
C11545 a_4093_43548# a_4235_43370# 0.515101f
C11546 a_n699_43396# a_1184_42692# 5.3e-21
C11547 a_10180_45724# a_n2661_43370# 0.038795f
C11548 a_n2293_46098# a_5663_43940# 0.142661f
C11549 a_21513_45002# a_21542_45572# 5.31e-19
C11550 a_n443_46116# a_2905_42968# 2.28e-19
C11551 a_n2293_46634# a_5565_43396# 2.79e-20
C11552 a_19900_46494# a_17517_44484# 2.41e-21
C11553 a_13259_45724# a_18248_44752# 0.003522f
C11554 a_16375_45002# a_16979_44734# 4.01e-20
C11555 a_8049_45260# a_8375_44464# 8.15e-22
C11556 a_n863_45724# a_2779_44458# 4.69e-21
C11557 a_n2293_45546# a_n699_43396# 4.61e-21
C11558 a_526_44458# a_n2293_43922# 1.43e-19
C11559 a_n1925_42282# a_n2661_43922# 0.028186f
C11560 a_2324_44458# a_11967_42832# 0.005512f
C11561 a_17715_44484# a_17325_44484# 1.25e-19
C11562 a_13507_46334# a_21259_43561# 1.05e-20
C11563 a_1138_42852# a_1414_42308# 4.35e-19
C11564 a_3357_43084# a_19963_31679# 0.009628f
C11565 a_19479_31679# a_22959_45572# 0.004153f
C11566 a_22223_45572# a_20447_31679# 2.46e-19
C11567 a_5807_45002# a_14358_43442# 4.13e-19
C11568 a_13661_43548# a_14579_43548# 8.17e-20
C11569 a_8696_44636# a_11963_45334# 5.44e-20
C11570 a_3316_45546# a_n2661_44458# 0.003189f
C11571 a_8270_45546# a_9165_43940# 0.063297f
C11572 a_2107_46812# a_8145_46902# 5.47e-21
C11573 a_n1925_46634# a_6755_46942# 0.12389f
C11574 a_n2661_46634# a_7832_46660# 0.001683f
C11575 a_5807_45002# a_11735_46660# 0.005164f
C11576 a_n1151_42308# a_1823_45246# 1.93e-19
C11577 a_3160_47472# a_2202_46116# 1.2e-19
C11578 a_12549_44172# a_14976_45028# 0.005173f
C11579 a_768_44030# a_3090_45724# 0.115303f
C11580 C6_P_btm VREF 1.41944f
C11581 a_11453_44696# a_16388_46812# 0.019353f
C11582 a_10227_46804# a_21363_46634# 0.273017f
C11583 C7_P_btm VREF_GND 1.61142f
C11584 C8_P_btm VCM 2.61094f
C11585 a_n237_47217# a_5204_45822# 0.019965f
C11586 a_n971_45724# a_6165_46155# 1.18e-20
C11587 a_n1741_47186# a_8199_44636# 4.26e-20
C11588 a_n443_46116# a_n1076_46494# 0.002776f
C11589 a_13717_47436# a_20202_43084# 1.46e-20
C11590 C8_N_btm C10_N_btm 0.878696f
C11591 a_13507_46334# a_765_45546# 0.045587f
C11592 a_18597_46090# a_20411_46873# 0.070431f
C11593 a_2905_45572# a_167_45260# 0.001572f
C11594 a_2063_45854# a_2804_46116# 0.007304f
C11595 a_584_46384# a_3147_46376# 6.53e-20
C11596 a_18479_47436# a_20841_46902# 0.006861f
C11597 a_16327_47482# a_16434_46660# 7.88e-19
C11598 C6_N_btm VDD 0.210613f
C11599 C4_P_btm VIN_P 0.50261f
C11600 a_4190_30871# a_4361_42308# 0.06171f
C11601 a_10695_43548# a_10991_42826# 8.2e-19
C11602 a_18114_32519# a_22469_39537# 2.15e-20
C11603 a_4905_42826# a_4649_43172# 9.93e-20
C11604 a_8685_43396# a_13635_43156# 3.19e-19
C11605 a_3422_30871# a_20107_42308# 3.36e-19
C11606 a_8016_46348# a_8685_43396# 7.84e-20
C11607 a_526_44458# a_n97_42460# 0.277959f
C11608 a_6431_45366# a_6298_44484# 0.006936f
C11609 a_6171_45002# a_8103_44636# 1.07e-20
C11610 a_n2017_45002# a_n356_44636# 0.036195f
C11611 a_6755_46942# a_16795_42852# 1.85e-20
C11612 a_5111_44636# a_10157_44484# 2.31e-20
C11613 a_16855_45546# a_11967_42832# 1.82e-21
C11614 a_3090_45724# a_5755_42852# 8.56e-21
C11615 a_4185_45028# a_14579_43548# 3.54e-21
C11616 a_3537_45260# a_8975_43940# 7.28e-19
C11617 a_5691_45260# a_5883_43914# 3.05e-21
C11618 a_5205_44484# a_5518_44484# 0.135771f
C11619 a_3232_43370# a_8701_44490# 0.062297f
C11620 a_n743_46660# a_6633_46155# 1.23e-19
C11621 a_10467_46802# a_11387_46155# 5.52e-19
C11622 a_10428_46928# a_10903_43370# 1.9e-19
C11623 a_5807_45002# a_14537_46482# 6.7e-19
C11624 a_6151_47436# a_7499_43078# 1.49e-19
C11625 a_6851_47204# a_7230_45938# 4.87e-21
C11626 a_11813_46116# a_3483_46348# 8.59e-21
C11627 a_2443_46660# a_2981_46116# 1.22e-19
C11628 a_n1925_46634# a_8049_45260# 0.088663f
C11629 a_n2661_46634# a_10586_45546# 0.001458f
C11630 a_19123_46287# a_20411_46873# 1.69e-20
C11631 a_18285_46348# a_20273_46660# 8.45e-20
C11632 a_16388_46812# a_17639_46660# 1.85e-19
C11633 a_2107_46812# a_5066_45546# 0.004218f
C11634 a_5257_43370# a_2324_44458# 0.067403f
C11635 a_6755_46942# a_10355_46116# 3.41e-20
C11636 a_10249_46116# a_9290_44172# 2.05e-19
C11637 a_12549_44172# a_18051_46116# 2.41e-20
C11638 a_4791_45118# a_8746_45002# 0.001033f
C11639 a_4915_47217# a_10180_45724# 1.08e-20
C11640 a_3090_45724# a_1176_45822# 5.71e-21
C11641 a_3080_42308# a_n4209_39304# 4.02e-21
C11642 a_743_42282# a_6481_42558# 0.001159f
C11643 a_15681_43442# a_15764_42576# 4.17e-19
C11644 a_14543_43071# a_14853_42852# 6.01e-20
C11645 a_5534_30871# a_13622_42852# 2.49e-19
C11646 a_2889_44172# VDD 0.1447f
C11647 a_15227_44166# a_15486_42560# 7.01e-19
C11648 a_8975_43940# a_11541_44484# 0.028558f
C11649 a_n443_46116# VDD 3.87014f
C11650 a_n1151_42308# DATA[2] 0.01294f
C11651 a_n863_45724# a_n13_43084# 0.041588f
C11652 a_2063_45854# CLK 0.271193f
C11653 a_n2312_38680# a_n2302_37984# 1.26e-19
C11654 a_3232_43370# a_11816_44260# 3.27e-19
C11655 a_3381_47502# DATA[1] 4.03e-22
C11656 a_9482_43914# a_15493_43396# 3.87e-21
C11657 a_n2661_43370# a_5013_44260# 3.07e-21
C11658 a_n2293_42834# a_n1644_44306# 5.64e-19
C11659 a_11827_44484# a_20512_43084# 0.030456f
C11660 a_20193_45348# a_22315_44484# 0.002679f
C11661 a_n443_42852# a_4361_42308# 0.016253f
C11662 a_2711_45572# a_16823_43084# 1.31e-19
C11663 a_n357_42282# a_n1991_42858# 8.06e-19
C11664 a_n755_45592# a_n1853_43023# 0.002072f
C11665 SMPL_ON_N a_22521_39511# 1.24e-19
C11666 a_526_44458# a_3935_43218# 6.08e-19
C11667 a_1307_43914# a_13483_43940# 0.00928f
C11668 a_18114_32519# a_19279_43940# 3.43e-19
C11669 a_15004_44636# a_14815_43914# 0.078606f
C11670 a_10355_46116# a_8049_45260# 0.003592f
C11671 a_8199_44636# a_10586_45546# 0.057648f
C11672 a_12816_46660# a_12791_45546# 3.25e-20
C11673 a_n1151_42308# a_14309_45028# 2.59e-21
C11674 a_768_44030# a_2274_45254# 0.001893f
C11675 a_8270_45546# a_8697_45822# 0.001837f
C11676 a_n2840_46090# a_n2810_45572# 4.48e-19
C11677 a_6545_47178# a_n2661_43370# 3.03e-20
C11678 a_n2956_39304# a_n2956_38680# 0.163045f
C11679 a_12991_46634# a_13163_45724# 3.39e-20
C11680 a_14226_46660# a_2711_45572# 3.51e-22
C11681 a_n743_46660# a_2437_43646# 0.031693f
C11682 a_11453_44696# a_13777_45326# 0.004241f
C11683 a_n1613_43370# a_3232_43370# 0.091534f
C11684 a_n881_46662# a_5691_45260# 1.46e-19
C11685 a_961_42354# a_5742_30871# 1.96e-20
C11686 a_4921_42308# a_7227_42308# 1.41e-19
C11687 a_6171_42473# a_5932_42308# 0.224949f
C11688 a_1606_42308# a_10533_42308# 1.94e-20
C11689 a_14621_43646# VDD 0.008139f
C11690 a_13887_32519# a_22469_39537# 1.15e-20
C11691 a_11967_42832# a_19862_44208# 3.19e-19
C11692 a_17609_46634# VDD 0.501057f
C11693 a_n984_44318# a_n875_44318# 0.007416f
C11694 a_n809_44244# a_n630_44306# 0.007399f
C11695 a_n1549_44318# a_n1441_43940# 0.057222f
C11696 a_n1899_43946# a_n822_43940# 1.46e-19
C11697 a_16292_46812# RST_Z 9.44e-21
C11698 a_n2661_44458# a_6197_43396# 1.22e-20
C11699 a_n913_45002# a_10922_42852# 0.01889f
C11700 a_n1059_45260# a_10341_42308# 0.032786f
C11701 a_n2017_45002# a_12379_42858# 2.94e-19
C11702 a_n2956_39304# a_n3690_39392# 0.016795f
C11703 a_n2956_38680# a_n3565_39304# 0.068534f
C11704 a_13259_45724# a_16522_42674# 9.98e-20
C11705 a_19615_44636# a_19478_44306# 0.004687f
C11706 a_3065_45002# a_3935_42891# 0.01149f
C11707 a_n443_42852# a_6761_42308# 0.00173f
C11708 a_n2661_42834# a_3992_43940# 3.11e-20
C11709 a_2998_44172# a_5013_44260# 0.004647f
C11710 a_n699_43396# a_2896_43646# 0.00787f
C11711 a_4646_46812# a_5883_43914# 0.019308f
C11712 a_12549_44172# a_15433_44458# 4.8e-20
C11713 a_n2293_46634# a_7640_43914# 7.73e-20
C11714 a_n2293_46098# a_3232_43370# 0.054403f
C11715 a_1823_45246# a_327_44734# 6.91e-21
C11716 a_n2438_43548# a_700_44734# 9.12e-20
C11717 a_6945_45028# a_18909_45814# 2.55e-22
C11718 a_10809_44734# a_18479_45785# 1.4e-21
C11719 a_9823_46155# a_3357_43084# 3.52e-21
C11720 a_18597_46090# a_3422_30871# 0.030159f
C11721 a_13259_45724# a_13527_45546# 0.00477f
C11722 a_167_45260# a_n37_45144# 0.277898f
C11723 a_509_45822# a_603_45572# 1.26e-19
C11724 a_n3565_39304# a_n3690_39392# 0.247167f
C11725 a_n3420_39616# a_n4209_38502# 0.028008f
C11726 a_n3565_39590# a_n3565_38502# 0.031189f
C11727 a_1239_39587# a_1239_39043# 0.054961f
C11728 a_n4334_39392# a_n3420_39072# 0.004849f
C11729 a_n4209_39304# a_n2946_39072# 0.022779f
C11730 a_n4209_39590# a_n3420_38528# 0.032196f
C11731 a_n4318_37592# VDD 0.919667f
C11732 a_n784_42308# C6_N_btm 5.52e-19
C11733 a_2553_47502# a_n1435_47204# 4.12e-19
C11734 a_4791_45118# a_6851_47204# 4.68e-20
C11735 a_4915_47217# a_6545_47178# 0.033555f
C11736 a_5129_47502# a_6151_47436# 1.77e-19
C11737 a_1606_42308# C2_P_btm 0.021793f
C11738 a_n913_45002# a_17531_42308# 2.07e-19
C11739 a_19443_46116# VDD 0.132317f
C11740 a_3422_30871# a_743_42282# 5.66e-19
C11741 a_4743_44484# a_4649_42852# 5.95e-21
C11742 a_15493_43940# a_2982_43646# 6.34e-20
C11743 a_11341_43940# a_3626_43646# 1.01e-21
C11744 a_n1059_45260# a_18057_42282# 0.141112f
C11745 a_n2017_45002# a_18727_42674# 8.71e-20
C11746 a_n2661_42834# a_9127_43156# 3.28e-20
C11747 a_n2661_43922# a_8387_43230# 4.36e-21
C11748 a_n2293_43922# a_8605_42826# 7.25e-21
C11749 a_n2293_42834# a_961_42354# 2.18e-20
C11750 a_9313_44734# a_12545_42858# 0.005689f
C11751 a_20692_30879# C7_N_btm 0.001136f
C11752 a_20205_31679# C8_N_btm 1.65e-20
C11753 a_5066_45546# a_n2661_44458# 8.22e-20
C11754 a_16375_45002# a_16321_45348# 0.009082f
C11755 a_18189_46348# a_18248_44752# 0.002127f
C11756 a_1609_45822# a_2304_45348# 0.002594f
C11757 a_17715_44484# a_18287_44626# 6.13e-20
C11758 a_5937_45572# a_5891_43370# 5.83e-19
C11759 a_13259_45724# a_16922_45042# 0.401687f
C11760 a_8199_44636# a_8238_44734# 0.003158f
C11761 a_12741_44636# a_15367_44484# 5.35e-20
C11762 a_3090_45724# a_7845_44172# 0.001391f
C11763 a_21588_30879# a_14401_32519# 0.058775f
C11764 a_2711_45572# a_15415_45028# 7.81e-20
C11765 a_526_44458# a_742_44458# 0.54618f
C11766 a_7499_43078# a_5111_44636# 0.753731f
C11767 a_12861_44030# a_15095_43370# 6.6e-19
C11768 a_10809_44734# a_10057_43914# 0.060542f
C11769 a_4883_46098# a_8791_43396# 0.001239f
C11770 a_n4334_37440# VDD 0.385859f
C11771 VDAC_P C3_P_btm 1.99006f
C11772 a_22717_37285# a_22717_36887# 0.003901f
C11773 a_n1613_43370# a_4651_46660# 0.686447f
C11774 a_4883_46098# a_10428_46928# 0.001889f
C11775 a_n2661_46634# a_n743_46660# 0.037388f
C11776 a_n2956_39768# a_n2438_43548# 8.21e-19
C11777 a_n1741_47186# a_765_45546# 0.536367f
C11778 a_13381_47204# a_12991_46634# 4.07e-19
C11779 a_n2293_46634# a_n2312_38680# 0.131017f
C11780 a_n2442_46660# a_n1925_46634# 6.55e-19
C11781 a_n1151_42308# a_12347_46660# 2.21e-19
C11782 a_n881_46662# a_4646_46812# 0.024758f
C11783 a_1115_44172# a_961_42354# 4.94e-20
C11784 a_1414_42308# a_1576_42282# 0.004774f
C11785 a_9313_44734# a_19332_42282# 2.91e-20
C11786 a_3537_45260# VDD 3.9063f
C11787 a_413_45260# DATA[3] 0.037695f
C11788 a_10341_43396# a_18783_43370# 0.010939f
C11789 a_n97_42460# a_8605_42826# 2.01e-20
C11790 a_n4318_39768# a_n3674_38680# 0.027425f
C11791 a_1568_43370# a_2075_43172# 0.006043f
C11792 a_1756_43548# a_1847_42826# 4.29e-19
C11793 a_8791_43396# a_5649_42852# 4.06e-22
C11794 a_10193_42453# a_11541_44484# 6.17e-19
C11795 a_7705_45326# a_n2293_42834# 0.071732f
C11796 a_n2293_46098# a_4905_42826# 0.004f
C11797 a_4927_45028# a_n2661_43370# 0.007616f
C11798 a_n863_45724# a_644_44056# 6.33e-20
C11799 a_10227_46804# a_15597_42852# 6.37e-19
C11800 a_2711_45572# a_19279_43940# 0.001969f
C11801 a_3232_43370# a_8704_45028# 3.4e-20
C11802 a_n755_45592# a_n1899_43946# 3.13e-19
C11803 a_8696_44636# a_18443_44721# 5.52e-20
C11804 a_10210_45822# a_9313_44734# 7.56e-21
C11805 a_n1099_45572# a_n809_44244# 2.33e-20
C11806 a_n1059_45260# a_18494_42460# 0.187733f
C11807 a_n913_45002# a_18184_42460# 3.93e-19
C11808 a_9290_44172# a_13565_43940# 1.77e-20
C11809 a_n443_46116# a_n784_42308# 2.29e-21
C11810 a_3090_45724# a_16759_43396# 7.41e-22
C11811 a_2107_46812# a_5068_46348# 0.007279f
C11812 a_n2661_46634# a_11189_46129# 1.44e-19
C11813 a_1431_47204# a_n755_45592# 1.62e-21
C11814 a_n2661_46098# a_2521_46116# 7.45e-20
C11815 a_3815_47204# a_n2661_45546# 1.03e-20
C11816 a_12816_46660# a_12925_46660# 0.007416f
C11817 a_12991_46634# a_13170_46660# 0.007399f
C11818 a_4883_46098# a_8283_46482# 7.98e-20
C11819 a_n746_45260# a_n356_45724# 0.030083f
C11820 a_n237_47217# a_3503_45724# 6.04e-21
C11821 a_n971_45724# a_n23_45546# 4.37e-19
C11822 a_584_46384# a_310_45028# 0.024195f
C11823 a_n1151_42308# a_n2293_45546# 0.01733f
C11824 a_15227_44166# a_19466_46812# 0.310201f
C11825 a_18834_46812# a_19692_46634# 1.69e-19
C11826 a_n1613_43370# a_n1379_46482# 0.001903f
C11827 a_2443_46660# a_167_45260# 0.012819f
C11828 a_n743_46660# a_8199_44636# 0.046048f
C11829 a_5807_45002# a_2324_44458# 0.232399f
C11830 a_16131_47204# a_15682_46116# 6.99e-20
C11831 a_13747_46662# a_15015_46420# 1.31e-19
C11832 a_13661_43548# a_14840_46494# 4.52e-20
C11833 a_5342_30871# a_16414_43172# 6.64e-20
C11834 a_3626_43646# a_10723_42308# 0.003809f
C11835 a_2982_43646# a_5742_30871# 0.196805f
C11836 a_11541_44484# VDD 0.004886f
C11837 a_16823_43084# a_16877_42852# 0.001502f
C11838 a_n2661_42834# CLK 3.56e-20
C11839 a_8147_43396# a_5934_30871# 1.84e-20
C11840 a_n97_42460# a_16104_42674# 0.007062f
C11841 a_4361_42308# a_14635_42282# 0.018479f
C11842 a_5147_45002# a_3905_42865# 0.048808f
C11843 a_3537_45260# a_5495_43940# 2.48e-20
C11844 a_n2312_39304# a_n4064_38528# 1.13e-20
C11845 a_n1059_45260# a_3499_42826# 0.002236f
C11846 a_10903_43370# a_12895_43230# 0.011631f
C11847 a_n357_42282# a_14205_43396# 6.12e-20
C11848 a_n1925_42282# a_n1641_43230# 1.11e-20
C11849 a_10157_44484# a_10334_44484# 0.159555f
C11850 a_8701_44490# a_8975_43940# 9.09e-19
C11851 a_5883_43914# a_10057_43914# 2.04e-20
C11852 a_n2267_44484# a_n2012_44484# 0.05936f
C11853 a_n2129_44697# a_n1809_44850# 0.026556f
C11854 a_3232_43370# a_2675_43914# 0.003881f
C11855 a_4185_45028# a_21671_42860# 2.44e-20
C11856 a_9290_44172# a_5534_30871# 0.472376f
C11857 a_13259_45724# a_15743_43084# 0.021493f
C11858 a_n881_46662# a_18479_45785# 9.48e-20
C11859 a_19787_47423# a_3357_43084# 0.001723f
C11860 a_n1423_46090# a_n2956_39304# 7.61e-21
C11861 a_n2157_46122# a_n1545_46494# 3.82e-19
C11862 a_n2293_46098# a_n1379_46482# 2.44e-19
C11863 a_4646_46812# a_8162_45546# 8.55e-19
C11864 a_n1151_42308# a_6709_45028# 0.286957f
C11865 a_13885_46660# a_13259_45724# 1.34e-21
C11866 a_13059_46348# a_14371_46494# 0.004662f
C11867 a_21177_47436# a_2437_43646# 0.014824f
C11868 a_13507_46334# a_21513_45002# 5.14e-19
C11869 a_5257_43370# a_6667_45809# 5.18e-20
C11870 a_9863_46634# a_2711_45572# 4.34e-20
C11871 a_2063_45854# a_10951_45334# 0.016425f
C11872 a_n1853_46287# a_n1736_46482# 0.170096f
C11873 a_n1991_46122# a_n2956_38680# 0.004896f
C11874 a_13747_46662# a_16333_45814# 0.018523f
C11875 a_5807_45002# a_16855_45546# 7.38e-19
C11876 a_13661_43548# a_16115_45572# 3.92e-20
C11877 a_20411_46873# a_8049_45260# 0.003303f
C11878 a_765_45546# a_10586_45546# 4.93e-20
C11879 a_12549_44172# a_13385_45572# 0.001759f
C11880 a_12891_46348# a_13485_45572# 4.18e-19
C11881 a_4791_45118# a_3232_43370# 0.268929f
C11882 a_15227_44166# a_20205_31679# 3.84e-19
C11883 a_9313_45822# a_413_45260# 2.11e-19
C11884 a_8953_45546# a_10355_46116# 3.1e-20
C11885 a_9625_46129# a_9823_46155# 0.321686f
C11886 a_8199_44636# a_11189_46129# 8.81e-19
C11887 a_1049_43396# VDD 0.196328f
C11888 a_21356_42826# a_17303_42282# 2.46e-20
C11889 a_5342_30871# a_7174_31319# 0.046616f
C11890 a_n3674_38216# a_n3674_37592# 0.048035f
C11891 a_n4318_38216# a_n1630_35242# 0.031712f
C11892 a_n4318_37592# a_n784_42308# 7e-20
C11893 COMP_P a_196_42282# 4.12e-21
C11894 a_3080_42308# C6_N_btm 2.67e-19
C11895 a_5891_43370# a_8333_44056# 0.070354f
C11896 a_19279_43940# a_22485_44484# 2.14e-20
C11897 a_13259_45724# a_1606_42308# 3.55e-20
C11898 a_n2956_38216# a_n3674_38680# 0.022975f
C11899 a_11827_44484# a_21381_43940# 0.002761f
C11900 a_n2661_43370# a_4699_43561# 4.75e-21
C11901 a_n2661_43922# a_n875_44318# 1.08e-19
C11902 a_n2661_42834# a_n630_44306# 3.44e-19
C11903 a_20640_44752# a_19237_31679# 7.45e-21
C11904 a_9482_43914# a_10695_43548# 1.47e-20
C11905 a_n357_42282# a_22400_42852# 1.12e-19
C11906 a_n2810_45572# a_n2104_42282# 2.3e-20
C11907 a_20692_30879# COMP_P 6.17e-20
C11908 a_n2293_42834# a_2982_43646# 0.019738f
C11909 a_20679_44626# a_22959_44484# 1.47e-21
C11910 a_18989_43940# a_19862_44208# 7.01e-21
C11911 a_20193_45348# a_19319_43548# 1.24e-19
C11912 a_8953_45002# a_10341_43396# 5.38e-21
C11913 a_14539_43914# a_15493_43940# 0.625897f
C11914 a_13777_45326# a_9145_43396# 1.2e-21
C11915 a_2324_44458# a_15143_45578# 0.002313f
C11916 a_526_44458# a_3733_45822# 3.36e-19
C11917 a_768_44030# a_4743_44484# 0.002819f
C11918 a_12741_44636# a_16789_45572# 1.15e-19
C11919 a_20107_46660# a_3357_43084# 0.025828f
C11920 a_3877_44458# a_n2661_43370# 0.038641f
C11921 a_3090_45724# a_7276_45260# 8.07e-21
C11922 a_n1613_43370# a_8975_43940# 4.75e-21
C11923 a_11415_45002# a_17668_45572# 0.002419f
C11924 a_20841_46902# a_2437_43646# 1.33e-20
C11925 w_11334_34010# a_3422_30871# 1.91172f
C11926 a_15559_46634# a_6171_45002# 3.5e-22
C11927 a_13059_46348# a_n913_45002# 2.23e-19
C11928 a_8199_44636# a_11136_45572# 0.001393f
C11929 a_11813_46116# a_11963_45334# 2.51e-19
C11930 a_10903_43370# a_11280_45822# 6.44e-19
C11931 a_10809_44734# a_10180_45724# 0.007361f
C11932 a_11387_46155# a_11682_45822# 2.23e-19
C11933 a_5527_46155# a_2711_45572# 1.62e-19
C11934 a_5066_45546# a_5907_45546# 9e-19
C11935 a_5934_30871# a_n4209_38216# 1.88e-21
C11936 a_n2833_47464# a_n2497_47436# 0.217831f
C11937 a_19511_42282# a_21613_42308# 0.001375f
C11938 a_13258_32519# a_21335_42336# 0.022004f
C11939 a_20107_42308# a_7174_31319# 0.175129f
C11940 a_22400_42852# CAL_N 0.001609f
C11941 a_4223_44672# a_7871_42858# 5.46e-20
C11942 a_11691_44458# a_17595_43084# 7.45e-21
C11943 a_11967_42832# a_14579_43548# 0.060711f
C11944 a_n913_45002# a_2903_42308# 0.041908f
C11945 a_n1059_45260# a_3318_42354# 3.58e-19
C11946 a_n2017_45002# a_3823_42558# 0.005755f
C11947 a_3357_43084# a_5932_42308# 2.19e-20
C11948 a_22223_46124# VDD 0.300745f
C11949 a_3905_42865# a_4093_43548# 0.032751f
C11950 a_6945_45028# RST_Z 0.022027f
C11951 a_20708_46348# SINGLE_ENDED 9.74e-21
C11952 a_11827_44484# a_18249_42858# 1.13e-20
C11953 a_n1441_43940# a_n1177_43370# 6.39e-20
C11954 a_3537_45260# a_n784_42308# 5.26e-20
C11955 a_18184_42460# a_20922_43172# 0.018236f
C11956 a_18494_42460# a_19987_42826# 0.098055f
C11957 a_5343_44458# a_5111_42852# 1.38e-21
C11958 a_768_44030# a_9248_44260# 2.63e-19
C11959 a_18189_46348# a_16922_45042# 0.015824f
C11960 a_10903_43370# a_11827_44484# 0.021644f
C11961 a_167_45260# a_949_44458# 0.021626f
C11962 a_1138_42852# a_n699_43396# 0.024181f
C11963 a_n2293_46634# a_10729_43914# 0.004608f
C11964 a_9290_44172# a_11691_44458# 3.23e-20
C11965 a_13249_42308# a_8696_44636# 0.021669f
C11966 a_12741_44636# a_14539_43914# 0.09527f
C11967 a_n2661_45546# a_2382_45260# 8.68e-19
C11968 a_n2293_45546# a_327_44734# 0.027309f
C11969 a_3090_45724# a_17517_44484# 0.020082f
C11970 a_13747_46662# a_15493_43396# 8.51e-22
C11971 a_3877_44458# a_2998_44172# 3.23e-20
C11972 a_4791_45118# a_4905_42826# 0.516502f
C11973 a_n443_46116# a_3080_42308# 3.12e-21
C11974 a_n755_45592# en_comp 1.09e-20
C11975 a_11823_42460# a_12561_45572# 0.004618f
C11976 a_12427_45724# a_12649_45572# 0.001658f
C11977 a_n357_42282# a_n967_45348# 0.003964f
C11978 a_n452_45724# a_n143_45144# 3.05e-21
C11979 a_n863_45724# a_n37_45144# 0.056531f
C11980 a_1823_45246# a_4223_44672# 0.008169f
C11981 a_17583_46090# a_17613_45144# 4.26e-20
C11982 a_12839_46116# a_13159_45002# 4.85e-20
C11983 a_13661_43548# a_19478_44306# 5.27e-20
C11984 a_n971_45724# a_8492_46660# 0.016456f
C11985 a_n237_47217# a_7927_46660# 0.008694f
C11986 a_n443_46116# a_4646_46812# 0.077958f
C11987 a_4915_47217# a_3877_44458# 8.8e-20
C11988 a_4791_45118# a_4651_46660# 0.020454f
C11989 a_1343_38525# VDD 3.25389f
C11990 a_12465_44636# a_20916_46384# 3.77e-19
C11991 a_n3420_38528# C6_P_btm 8.47e-20
C11992 a_n3565_38502# C4_P_btm 0.042623f
C11993 a_n3565_38216# EN_VIN_BSTR_P 0.005343f
C11994 a_n1151_42308# a_5732_46660# 9.82e-22
C11995 a_4700_47436# a_4955_46873# 0.001297f
C11996 a_n1435_47204# a_1799_45572# 3.59e-20
C11997 a_n881_46662# a_9804_47204# 0.061323f
C11998 a_7989_47542# a_8128_46384# 5.76e-19
C11999 a_4883_46098# a_22612_30879# 9.37e-21
C12000 a_21811_47423# a_21588_30879# 8.73e-19
C12001 a_n3565_37414# a_n4064_37440# 0.230258f
C12002 a_3754_38470# a_3726_37500# 0.554457f
C12003 VDAC_Ni a_5088_37509# 1.70462f
C12004 a_11453_44696# a_19321_45002# 0.023175f
C12005 en_comp a_22521_40599# 0.021604f
C12006 a_n2661_42834# a_1755_42282# 8.39e-21
C12007 a_16842_45938# VDD 4.6e-19
C12008 a_n97_42460# a_18783_43370# 0.00416f
C12009 a_3626_43646# a_10341_43396# 5.18e-20
C12010 a_20193_45348# a_21335_42336# 4.79e-20
C12011 a_8791_43396# a_8685_43396# 0.086218f
C12012 a_6452_43396# a_6643_43396# 4.61e-19
C12013 a_13483_43940# a_13635_43156# 4.94e-20
C12014 a_17478_45572# a_16922_45042# 3.77e-20
C12015 a_15861_45028# a_17023_45118# 0.076138f
C12016 a_3429_45260# a_3232_43370# 0.001753f
C12017 a_4558_45348# a_5111_44636# 0.009468f
C12018 a_n443_42852# a_5891_43370# 0.175668f
C12019 a_2382_45260# a_5205_44484# 1.09e-21
C12020 a_n913_45002# a_13556_45296# 7.49e-21
C12021 a_4574_45260# a_4927_45028# 0.047624f
C12022 a_16327_47482# a_19339_43156# 0.346029f
C12023 a_3357_43084# a_1423_45028# 0.02044f
C12024 a_3537_45260# a_5691_45260# 9.13e-19
C12025 a_8049_45260# a_3422_30871# 2.49e-20
C12026 a_8696_44636# a_17613_45144# 0.09062f
C12027 a_12465_44636# a_12545_42858# 1.55e-20
C12028 a_9049_44484# a_10157_44484# 1.97e-19
C12029 a_7499_43078# a_10334_44484# 1.72e-19
C12030 a_n1099_45572# a_n2661_42834# 2.37e-21
C12031 a_380_45546# a_n2661_43922# 1e-20
C12032 a_2063_45854# a_n1925_42282# 0.025501f
C12033 a_n1151_42308# a_n914_46116# 2.87e-19
C12034 a_6851_47204# a_6945_45028# 0.013916f
C12035 a_12861_44030# a_17583_46090# 2.84e-20
C12036 a_13661_43548# a_19636_46660# 3.05e-20
C12037 a_n881_46662# a_n901_46420# 0.053662f
C12038 a_n1613_43370# a_n1076_46494# 0.232314f
C12039 a_4883_46098# a_7920_46348# 0.006584f
C12040 a_11599_46634# a_15015_46420# 0.040858f
C12041 a_10227_46804# a_11133_46155# 0.019137f
C12042 a_14955_47212# a_14840_46494# 7.46e-21
C12043 a_7927_46660# a_8270_45546# 8.4e-21
C12044 a_7577_46660# a_8601_46660# 2.36e-20
C12045 a_2747_46873# a_2698_46116# 0.006795f
C12046 a_n743_46660# a_765_45546# 0.148721f
C12047 a_1239_47204# a_1337_46116# 6.31e-21
C12048 a_n1557_42282# a_n2104_42282# 3.45e-19
C12049 a_685_42968# a_791_42968# 0.13675f
C12050 a_4190_30871# a_17595_43084# 7.76e-19
C12051 a_13467_32519# a_5534_30871# 0.041703f
C12052 a_8701_44490# VDD 0.164475f
C12053 a_n2293_43922# VDAC_N 6.46e-20
C12054 a_3422_30871# a_n4064_37984# 0.031408f
C12055 a_15493_43396# a_4958_30871# 1.31e-20
C12056 a_5649_42852# a_12895_43230# 9.12e-21
C12057 a_743_42282# a_16414_43172# 5.93e-20
C12058 a_n4318_39768# a_n2860_39866# 4.42e-20
C12059 a_n2293_46634# a_5932_42308# 3.78e-20
C12060 a_10193_42453# a_11816_44260# 1.82e-19
C12061 a_n755_45592# a_n1699_43638# 1.23e-19
C12062 a_n357_42282# a_n1917_43396# 6.93e-20
C12063 a_n2661_43370# a_10440_44484# 9.47e-21
C12064 a_21101_45002# a_18114_32519# 1.7e-19
C12065 a_19479_31679# a_3422_30871# 2.13e-21
C12066 a_8199_44636# a_4361_42308# 0.024061f
C12067 a_17339_46660# a_18083_42858# 0.001069f
C12068 SMPL_ON_P a_n3565_38216# 6.6e-19
C12069 a_10775_45002# a_n2661_43922# 8.33e-21
C12070 a_1423_45028# a_5826_44734# 0.003941f
C12071 a_10951_45334# a_n2661_42834# 1.25e-20
C12072 a_n863_45724# a_104_43370# 0.046664f
C12073 a_12549_44172# a_12563_42308# 1.25e-20
C12074 a_526_44458# a_9885_43646# 0.008704f
C12075 a_n743_46660# a_509_45822# 0.039863f
C12076 a_2443_46660# a_n863_45724# 5.17e-22
C12077 a_13059_46348# a_14493_46090# 0.029059f
C12078 a_n1853_46287# a_n1641_46494# 0.033696f
C12079 a_n1991_46122# a_n1423_46090# 0.175891f
C12080 a_12861_44030# a_8696_44636# 0.046746f
C12081 a_11599_46634# a_16333_45814# 3.08e-19
C12082 a_15811_47375# a_15903_45785# 3.35e-20
C12083 a_n2293_46098# a_n1076_46494# 0.006462f
C12084 a_n2157_46122# a_n901_46420# 0.043559f
C12085 a_765_45546# a_11189_46129# 2.79e-21
C12086 a_19692_46634# a_10809_44734# 0.014397f
C12087 a_10623_46897# a_10586_45546# 5.93e-19
C12088 a_8035_47026# a_8034_45724# 1.67e-20
C12089 a_5807_45002# a_6667_45809# 2.91e-19
C12090 a_n2293_42282# a_1755_42282# 0.875855f
C12091 a_743_42282# a_7174_31319# 0.004769f
C12092 a_20556_43646# a_20712_42282# 1.47e-20
C12093 a_4361_42308# a_19511_42282# 0.071032f
C12094 a_5342_30871# a_5932_42308# 0.01856f
C12095 a_14401_32519# a_22469_39537# 1.48e-20
C12096 a_3315_47570# DATA[2] 9.25e-20
C12097 a_n1059_45260# a_6197_43396# 4.64e-20
C12098 a_4185_45028# a_9223_42460# 8.35e-20
C12099 a_6298_44484# a_6453_43914# 0.002276f
C12100 a_n2012_44484# a_n2065_43946# 7.1e-20
C12101 a_n357_42282# a_22223_42860# 4.11e-19
C12102 a_1823_45246# a_5742_30871# 4.25e-20
C12103 a_16922_45042# a_20935_43940# 1.08e-20
C12104 a_3357_43084# a_4181_43396# 1.16e-20
C12105 a_15463_44811# a_14673_44172# 0.001037f
C12106 a_n1177_44458# a_n1441_43940# 7.12e-20
C12107 a_5343_44458# a_7542_44172# 0.014194f
C12108 a_18911_45144# a_15493_43396# 2.88e-21
C12109 a_19778_44110# a_19328_44172# 0.064774f
C12110 a_18494_42460# a_18326_43940# 1.27e-19
C12111 a_n1613_43370# VDD 4.75085f
C12112 a_n913_45002# a_6293_42852# 0.001086f
C12113 a_11827_44484# a_14955_43940# 0.005645f
C12114 a_413_45260# a_2982_43646# 7.3e-22
C12115 a_5883_43914# a_5013_44260# 0.001282f
C12116 a_4574_45260# a_4699_43561# 3.74e-21
C12117 a_3537_45260# a_3080_42308# 0.02683f
C12118 a_9290_44172# a_n443_42852# 0.483812f
C12119 a_22959_46124# a_20205_31679# 0.012679f
C12120 a_10809_44734# a_20692_30879# 0.006707f
C12121 a_n746_45260# a_n356_44636# 0.418585f
C12122 a_n971_45724# a_n23_44458# 1.18e-20
C12123 a_4646_46812# a_3537_45260# 0.361823f
C12124 a_3877_44458# a_4574_45260# 0.010367f
C12125 a_8128_46384# a_n2661_43370# 3.48e-20
C12126 a_17609_46634# a_18479_45785# 4.93e-20
C12127 a_15227_44166# a_16147_45260# 0.282941f
C12128 a_16327_47482# a_19721_31679# 1.56e-20
C12129 a_2324_44458# a_n755_45592# 1.99e-20
C12130 a_5164_46348# a_5263_45724# 0.005959f
C12131 a_6945_45028# a_21167_46155# 7.16e-19
C12132 a_6540_46812# a_413_45260# 1.57e-21
C12133 a_13059_46348# a_15903_45785# 9.2e-19
C12134 a_3090_45724# a_19256_45572# 7.35e-19
C12135 a_4791_45118# a_8975_43940# 2.73e-20
C12136 a_3483_46348# a_6598_45938# 3.25e-21
C12137 a_6165_46155# a_2711_45572# 9.84e-19
C12138 a_n2293_46634# a_1423_45028# 0.025918f
C12139 a_n2438_43548# a_1307_43914# 0.006717f
C12140 a_n743_46660# a_16751_45260# 0.028358f
C12141 a_13657_42558# a_15486_42560# 1.21e-20
C12142 a_14113_42308# a_15051_42282# 0.077852f
C12143 a_n784_42308# a_1343_38525# 2.98e-20
C12144 a_5755_42308# a_7174_31319# 9.76e-21
C12145 a_11551_42558# a_11633_42308# 0.003935f
C12146 a_n1533_42852# VDD 0.142813f
C12147 a_n2293_42834# a_7871_42858# 0.027f
C12148 a_11823_42460# a_11323_42473# 0.0014f
C12149 a_2382_45260# a_3863_42891# 6.79e-20
C12150 a_453_43940# a_726_44056# 0.001159f
C12151 a_n2293_46098# VDD 1.7963f
C12152 a_n2293_43922# a_3626_43646# 0.03147f
C12153 a_n2661_42834# a_n1243_43396# 9.21e-20
C12154 a_1467_44172# a_1443_43940# 0.011516f
C12155 a_1414_42308# a_1241_43940# 0.005139f
C12156 a_20202_43084# EN_OFFSET_CAL 0.001606f
C12157 a_9672_43914# a_10729_43914# 1.18e-19
C12158 a_20766_44850# a_20974_43370# 4.78e-21
C12159 a_n1059_45260# a_10752_42852# 1.72e-19
C12160 a_n913_45002# a_11554_42852# 0.016237f
C12161 a_2711_45572# a_19332_42282# 0.004712f
C12162 a_3537_45260# a_7309_43172# 4.53e-19
C12163 a_16327_47482# a_17973_43940# 0.001972f
C12164 a_11599_46634# a_15493_43396# 2.13e-21
C12165 a_6472_45840# a_6469_45572# 2.36e-20
C12166 a_6945_45028# a_3232_43370# 2.77e-19
C12167 a_7499_43078# a_9049_44484# 8.37e-20
C12168 a_526_44458# a_n467_45028# 1.12e-20
C12169 a_8049_45260# a_19963_31679# 0.2062f
C12170 a_17339_46660# a_18450_45144# 3.54e-19
C12171 a_12861_44030# a_20365_43914# 0.044371f
C12172 a_13759_46122# a_14180_45002# 1.47e-20
C12173 a_2711_45572# a_10210_45822# 0.007317f
C12174 a_20202_43084# a_16922_45042# 1.58e-19
C12175 a_11415_45002# a_16501_45348# 9.97e-19
C12176 a_13259_45724# a_17668_45572# 0.050071f
C12177 a_20411_46873# a_20193_45348# 0.002202f
C12178 a_n1613_43370# a_5495_43940# 8.26e-21
C12179 a_768_44030# a_1414_42308# 0.072003f
C12180 a_3090_45724# a_13720_44458# 2.05e-21
C12181 a_1823_45246# a_n2293_42834# 0.031316f
C12182 a_n1641_46494# a_n2661_43370# 2.3e-20
C12183 a_5257_43370# a_5708_44484# 0.056224f
C12184 a_2324_44458# a_13017_45260# 0.021259f
C12185 a_14275_46494# a_9482_43914# 8.66e-21
C12186 a_16023_47582# a_12465_44636# 4.1e-19
C12187 a_10227_46804# a_13507_46334# 0.120657f
C12188 a_n4209_39304# a_n4064_37440# 0.029715f
C12189 a_13249_42558# VDD 0.009141f
C12190 a_n3565_39590# VDAC_P 0.001403f
C12191 a_18597_46090# a_19787_47423# 0.001396f
C12192 a_2684_37794# VDAC_Pi 0.133177f
C12193 a_n3565_39304# a_n3420_37440# 0.032339f
C12194 a_n4064_39072# a_n4209_37414# 0.030589f
C12195 a_n3420_39072# a_n3565_37414# 0.031846f
C12196 a_n4064_37984# a_n3607_38304# 4.68e-19
C12197 a_n3420_37984# a_n2860_37984# 0.003211f
C12198 a_22465_38105# a_22545_38993# 0.253407f
C12199 a_n2497_47436# a_n2293_46634# 0.174929f
C12200 SMPL_ON_P a_n2840_46634# 8.18e-19
C12201 a_n2288_47178# a_n2442_46660# 0.009097f
C12202 a_n1920_47178# a_n2661_46634# 1.7e-19
C12203 a_n1741_47186# a_n2956_39768# 1.86e-19
C12204 a_4958_30871# C9_P_btm 0.209166f
C12205 a_n1435_47204# a_2747_46873# 1.47e-19
C12206 a_6491_46660# a_n1613_43370# 0.071408f
C12207 a_6545_47178# a_n881_46662# 0.020203f
C12208 a_16588_47582# a_4883_46098# 6.92e-21
C12209 a_18479_47436# a_20990_47178# 0.003332f
C12210 a_4915_47217# a_8128_46384# 0.070866f
C12211 a_2675_43914# a_2905_42968# 9.88e-21
C12212 a_n4318_39768# a_n4318_38680# 0.02372f
C12213 a_n3674_39768# a_n3674_39304# 0.037712f
C12214 a_18579_44172# a_18083_42858# 2.69e-21
C12215 a_n2956_37592# a_n2946_38778# 2.49e-19
C12216 a_7230_45938# VDD 0.077608f
C12217 a_11967_42832# a_21671_42860# 1.16e-19
C12218 a_9313_44734# a_13157_43218# 1.2e-19
C12219 a_20935_43940# a_15743_43084# 6.65e-21
C12220 a_15493_43940# a_17324_43396# 1.55e-20
C12221 a_11341_43940# a_18525_43370# 1.4e-19
C12222 a_458_43396# a_766_43646# 0.017351f
C12223 a_n1177_43370# a_n998_43396# 0.007399f
C12224 a_n1352_43396# a_n1243_43396# 0.007416f
C12225 a_n97_42460# a_3626_43646# 0.394673f
C12226 a_n699_43396# a_1576_42282# 7.71e-23
C12227 a_15682_43940# a_16823_43084# 7.58e-19
C12228 a_14021_43940# a_14621_43646# 0.001689f
C12229 a_15903_45785# a_13556_45296# 1.89e-19
C12230 a_n2293_46098# a_5495_43940# 0.096987f
C12231 a_3357_43084# a_22591_45572# 0.181818f
C12232 a_n2293_46634# a_4181_43396# 3.92e-20
C12233 a_526_44458# a_n2661_43922# 0.154533f
C12234 a_20075_46420# a_17517_44484# 6e-21
C12235 a_n863_45724# a_949_44458# 0.034335f
C12236 a_16375_45002# a_14539_43914# 3.75e-20
C12237 a_13259_45724# a_17970_44736# 0.011308f
C12238 a_n1925_42282# a_n2661_42834# 0.029302f
C12239 a_1138_42852# a_1467_44172# 0.034446f
C12240 a_19479_31679# a_19963_31679# 0.104687f
C12241 a_2437_43646# a_20447_31679# 1.16e-19
C12242 a_21513_45002# a_21297_45572# 1.2e-19
C12243 a_n443_46116# a_2075_43172# 0.002146f
C12244 a_13661_43548# a_13667_43396# 0.168674f
C12245 a_167_45260# a_175_44278# 5.9e-20
C12246 a_n2661_45546# a_5343_44458# 1.16e-20
C12247 a_8696_44636# a_11787_45002# 5.52e-20
C12248 a_8049_45260# a_7640_43914# 0.003041f
C12249 a_15037_45618# a_14797_45144# 0.003975f
C12250 a_3218_45724# a_n2661_44458# 3.08e-20
C12251 a_8270_45546# a_8487_44056# 1.88e-19
C12252 C7_P_btm VREF 1.818f
C12253 C8_P_btm VREF_GND 2.58605f
C12254 C9_P_btm VCM 6.06251f
C12255 C7_N_btm C10_N_btm 0.680974f
C12256 C8_N_btm C9_N_btm 29.256199f
C12257 C5_N_btm VDD 0.267489f
C12258 C5_P_btm VIN_P 0.502041f
C12259 a_2107_46812# a_7577_46660# 1.05e-19
C12260 a_5807_45002# a_11186_47026# 0.003092f
C12261 a_3160_47472# a_1823_45246# 0.002764f
C12262 a_12549_44172# a_3090_45724# 0.082348f
C12263 a_11453_44696# a_13059_46348# 0.039573f
C12264 a_10227_46804# a_20623_46660# 0.156341f
C12265 a_n237_47217# a_5164_46348# 0.081549f
C12266 a_n2109_47186# a_5937_45572# 0.00225f
C12267 a_n443_46116# a_n901_46420# 0.367344f
C12268 a_n1151_42308# a_1138_42852# 1.84e-20
C12269 a_13507_46334# a_17339_46660# 0.05814f
C12270 a_18597_46090# a_20107_46660# 0.001674f
C12271 a_2443_46660# a_5072_46660# 1.72e-21
C12272 a_n743_46660# a_10623_46897# 7.67e-20
C12273 a_18479_47436# a_20273_46660# 0.018124f
C12274 a_584_46384# a_2804_46116# 1.93e-19
C12275 a_2553_47502# a_2521_46116# 7.08e-19
C12276 a_2063_45854# a_2698_46116# 0.006352f
C12277 a_21259_43561# a_4361_42308# 0.005186f
C12278 a_4190_30871# a_13467_32519# 0.032722f
C12279 a_10695_43548# a_10796_42968# 6.99e-20
C12280 a_8704_45028# VDD 0.004293f
C12281 a_3422_30871# a_13258_32519# 0.410904f
C12282 a_n2661_42282# a_5934_30871# 2.9e-20
C12283 a_3626_43646# a_3935_43218# 6.34e-19
C12284 a_13661_43548# a_20256_43172# 5.04e-19
C12285 w_11334_34010# a_7174_31319# 7.7e-19
C12286 a_6171_45002# a_6298_44484# 0.001994f
C12287 a_3232_43370# a_8103_44636# 0.013825f
C12288 a_n443_42852# a_10807_43548# 0.173997f
C12289 a_n2293_45010# a_n23_44458# 1.13e-19
C12290 a_n2017_45002# a_n1655_44484# 6.5e-19
C12291 a_3357_43084# a_6109_44484# 0.016236f
C12292 a_5111_44636# a_9838_44484# 1.88e-22
C12293 a_16115_45572# a_11967_42832# 1.12e-20
C12294 a_8696_44636# a_17325_44484# 5.02e-20
C12295 a_3090_45724# a_5111_42852# 5.57e-21
C12296 a_n357_42282# a_20269_44172# 1.22e-20
C12297 a_3483_46348# a_14358_43442# 1.32e-20
C12298 a_20202_43084# a_15743_43084# 0.021267f
C12299 a_3537_45260# a_10057_43914# 0.001231f
C12300 a_5205_44484# a_5343_44458# 0.129692f
C12301 a_n1613_43370# a_n784_42308# 0.002725f
C12302 a_n743_46660# a_6347_46155# 1.92e-19
C12303 a_6151_47436# a_8568_45546# 6.1e-21
C12304 a_11735_46660# a_3483_46348# 6.06e-21
C12305 a_4651_46660# a_6945_45028# 2.58e-21
C12306 a_19123_46287# a_20107_46660# 4.05e-20
C12307 a_18285_46348# a_20411_46873# 3.41e-21
C12308 a_2107_46812# a_5431_46482# 8.38e-19
C12309 a_10249_46116# a_10355_46116# 0.182836f
C12310 a_10467_46802# a_11133_46155# 0.001412f
C12311 a_10554_47026# a_9290_44172# 0.003141f
C12312 a_n1151_42308# a_11962_45724# 8.76e-37
C12313 a_16023_47582# a_2711_45572# 8.57e-20
C12314 a_4915_47217# a_10053_45546# 3.01e-22
C12315 a_3080_42308# a_1343_38525# 3.95e-19
C12316 a_743_42282# a_5932_42308# 0.024532f
C12317 a_4361_42308# a_4921_42308# 0.472085f
C12318 a_15681_43442# a_15486_42560# 2.96e-20
C12319 a_16414_43172# a_16328_43172# 0.001377f
C12320 a_2675_43914# VDD 0.200923f
C12321 a_15227_44166# a_15051_42282# 2.31e-20
C12322 a_8975_43940# a_10809_44484# 5.15e-19
C12323 a_4791_45118# VDD 3.05095f
C12324 a_1423_45028# a_9672_43914# 4.02e-19
C12325 a_3160_47472# DATA[2] 5.43e-20
C12326 a_n863_45724# a_n1076_43230# 1.91e-20
C12327 a_n1925_42282# a_n2293_42282# 0.234055f
C12328 a_526_44458# a_3445_43172# 2.76e-19
C12329 a_9290_44172# a_14635_42282# 3.64e-19
C12330 a_13249_42308# a_14205_43396# 5.12e-22
C12331 a_3232_43370# a_11173_44260# 0.002786f
C12332 a_n1151_42308# DATA[1] 0.009539f
C12333 a_21359_45002# a_20512_43084# 7.4e-21
C12334 a_20193_45348# a_3422_30871# 0.042753f
C12335 a_11827_44484# a_21145_44484# 0.001286f
C12336 a_n755_45592# a_n2157_42858# 1.64e-22
C12337 a_n357_42282# a_n1853_43023# 0.04297f
C12338 a_n2956_38216# a_n4318_38680# 0.023204f
C12339 a_18114_32519# a_20766_44850# 2.21e-19
C12340 a_20205_45028# a_19279_43940# 6.24e-19
C12341 a_1307_43914# a_12429_44172# 0.007436f
C12342 a_n2661_43370# a_5244_44056# 4.22e-21
C12343 a_9823_46155# a_8049_45260# 0.004922f
C12344 a_12991_46634# a_12791_45546# 5.89e-20
C12345 a_12816_46660# a_11823_42460# 1.3e-20
C12346 a_8270_45546# a_8336_45822# 0.009698f
C12347 a_n2840_46090# a_n2840_45546# 0.025171f
C12348 a_6151_47436# a_n2661_43370# 0.003024f
C12349 a_n881_46662# a_4927_45028# 0.001762f
C12350 a_13507_46334# a_1307_43914# 3.03e-20
C12351 a_12465_44636# a_14797_45144# 0.002814f
C12352 a_11453_44696# a_13556_45296# 0.027553f
C12353 a_n1613_43370# a_5691_45260# 5.61e-21
C12354 a_17364_32525# a_22459_39145# 1.15e-20
C12355 a_1184_42692# a_5742_30871# 1.12e-20
C12356 a_4921_42308# a_6761_42308# 9.41e-19
C12357 a_5755_42308# a_5932_42308# 0.196877f
C12358 a_14537_43646# VDD 0.008942f
C12359 a_14209_32519# a_22521_39511# 8.25e-21
C12360 a_3823_42558# a_4169_42308# 0.013377f
C12361 a_8696_44636# a_8495_42852# 8.39e-21
C12362 a_11827_44484# a_8685_43396# 3.35e-20
C12363 a_16292_46812# VDD 0.123916f
C12364 a_n1331_43914# a_n1441_43940# 0.097745f
C12365 a_n1761_44111# a_n822_43940# 2.49e-19
C12366 a_3600_43914# a_3905_42865# 1.98e-20
C12367 a_2998_44172# a_5244_44056# 3.3e-19
C12368 a_15559_46634# RST_Z 1.85e-21
C12369 a_n913_45002# a_10991_42826# 0.029878f
C12370 a_n1059_45260# a_10922_42852# 0.002568f
C12371 a_n2017_45002# a_10341_42308# 0.049998f
C12372 a_n2956_39304# a_n3565_39304# 0.307358f
C12373 a_11967_42832# a_19478_44306# 2.52e-19
C12374 a_2779_44458# a_2982_43646# 1.05e-20
C12375 a_742_44458# a_3626_43646# 3.38e-20
C12376 a_3065_45002# a_3681_42891# 1.71e-20
C12377 a_11901_46660# CLK 6.62e-20
C12378 a_n699_43396# a_1987_43646# 2.2e-19
C12379 a_n2661_42834# a_3737_43940# 3.81e-20
C12380 a_509_45822# a_509_45572# 6.96e-20
C12381 a_n443_42852# a_n89_45572# 5.42e-19
C12382 a_5807_45002# a_5708_44484# 3.53e-20
C12383 a_n2293_46634# a_6109_44484# 2.18e-19
C12384 a_12549_44172# a_14815_43914# 0.026324f
C12385 a_768_44030# a_14112_44734# 0.004013f
C12386 a_1823_45246# a_413_45260# 0.043122f
C12387 a_n443_46116# a_5013_44260# 7.51e-21
C12388 a_4791_45118# a_5495_43940# 8.22e-20
C12389 a_13507_46334# a_18579_44172# 2e-20
C12390 a_n2661_45546# a_4880_45572# 0.003682f
C12391 a_10809_44734# a_18175_45572# 1.39e-20
C12392 a_14976_45028# a_15060_45348# 0.005133f
C12393 a_3090_45724# a_15685_45394# 4.27e-20
C12394 a_1138_42852# a_327_44734# 1.41e-19
C12395 a_18597_46090# a_21398_44850# 0.002638f
C12396 a_3503_45724# a_4099_45572# 1.81e-19
C12397 a_13259_45724# a_13163_45724# 0.166368f
C12398 a_9569_46155# a_3357_43084# 1.93e-20
C12399 a_167_45260# a_n143_45144# 0.03701f
C12400 a_2063_45854# a_n1435_47204# 0.001106f
C12401 a_5129_47502# a_5815_47464# 4.88e-20
C12402 a_4791_45118# a_6491_46660# 0.002326f
C12403 a_4915_47217# a_6151_47436# 0.783303f
C12404 a_n443_46116# a_6545_47178# 0.001077f
C12405 a_7174_31319# a_n4064_37984# 0.003259f
C12406 a_n1736_42282# VDD 0.227152f
C12407 a_n4209_39304# a_n3420_39072# 0.071714f
C12408 a_n4334_39392# a_n3690_39392# 8.67e-19
C12409 a_n1741_47186# a_10227_46804# 0.020904f
C12410 a_1606_42308# C3_P_btm 5.68e-19
C12411 a_n784_42308# C5_N_btm 5.81e-19
C12412 a_n2661_44458# a_11554_42852# 3.79e-20
C12413 a_n1059_45260# a_17531_42308# 0.001278f
C12414 a_n913_45002# a_17303_42282# 1.81467f
C12415 a_19963_31679# a_13258_32519# 0.054679f
C12416 a_1307_43914# a_7227_42308# 7.17e-37
C12417 a_n2017_45002# a_18057_42282# 4.4e-19
C12418 a_9159_44484# a_8952_43230# 1.71e-20
C12419 a_n2293_43922# a_8037_42858# 1.82e-20
C12420 a_n2661_42834# a_8387_43230# 2.69e-20
C12421 a_n2293_42834# a_1184_42692# 6.11e-20
C12422 a_9313_44734# a_12089_42308# 0.011899f
C12423 a_20205_31679# C7_N_btm 1.43e-20
C12424 a_20692_30879# C6_N_btm 0.080378f
C12425 a_10809_44734# a_10440_44484# 0.002452f
C12426 a_18189_46348# a_17970_44736# 5.88e-19
C12427 a_17715_44484# a_18248_44752# 5.78e-20
C12428 a_8199_44636# a_5891_43370# 0.399007f
C12429 a_5937_45572# a_8375_44464# 1.42e-20
C12430 a_17478_45572# a_17668_45572# 0.045837f
C12431 a_3090_45724# a_7542_44172# 0.137368f
C12432 a_2277_45546# a_1423_45028# 9.3e-22
C12433 a_2711_45572# a_14797_45144# 4.99e-20
C12434 a_526_44458# a_n452_44636# 3.8e-20
C12435 a_8953_45546# a_7640_43914# 1.62e-20
C12436 a_12861_44030# a_14205_43396# 6.35e-20
C12437 a_4883_46098# a_8147_43396# 6.45e-20
C12438 a_n2497_47436# a_743_42282# 2.68e-22
C12439 a_n881_46662# a_3877_44458# 0.142507f
C12440 a_n1613_43370# a_4646_46812# 1.38979f
C12441 a_n4209_37414# VDD 0.817347f
C12442 a_4883_46098# a_10150_46912# 0.001971f
C12443 a_8530_39574# RST_Z 0.431385f
C12444 a_n2840_46634# a_n2438_43548# 0.002664f
C12445 VDAC_P C4_P_btm 3.9276f
C12446 a_n2661_46634# a_n1021_46688# 0.009022f
C12447 a_n2472_46634# a_n1925_46634# 0.001266f
C12448 a_n2442_46660# a_n2312_38680# 0.068683f
C12449 a_n2293_46634# a_n2104_46634# 0.042499f
C12450 a_n1151_42308# a_12978_47026# 1.07e-19
C12451 a_1115_44172# a_1184_42692# 1.35e-20
C12452 a_1467_44172# a_1576_42282# 1.16e-20
C12453 a_9313_44734# a_18907_42674# 4.46e-21
C12454 a_10341_43396# a_18525_43370# 0.015853f
C12455 a_413_45260# DATA[2] 0.048779f
C12456 a_n97_42460# a_8037_42858# 4.35e-19
C12457 a_n1761_44111# a_n327_42308# 1.97e-19
C12458 a_1414_42308# a_1067_42314# 0.100434f
C12459 a_3429_45260# VDD 0.142923f
C12460 a_1568_43370# a_1847_42826# 0.153113f
C12461 a_6709_45028# a_n2293_42834# 0.001466f
C12462 a_n2293_46098# a_3080_42308# 5.04e-19
C12463 a_5111_44636# a_n2661_43370# 0.075649f
C12464 a_n863_45724# a_175_44278# 0.113317f
C12465 a_13059_46348# a_9145_43396# 0.028786f
C12466 a_17478_45572# a_17970_44736# 3.84e-19
C12467 a_n755_45592# a_n1761_44111# 0.015303f
C12468 a_3232_43370# a_7735_45067# 0.001345f
C12469 a_8696_44636# a_18287_44626# 8.04e-20
C12470 a_n1613_43370# a_7309_43172# 7.87e-19
C12471 a_n1099_45572# a_n1549_44318# 2.98e-21
C12472 a_584_46384# a_1755_42282# 8.38e-21
C12473 a_4791_45118# a_n784_42308# 4.27e-20
C12474 a_9290_44172# a_11257_43940# 6.04e-19
C12475 a_626_44172# a_1423_45028# 0.014461f
C12476 w_11334_34010# a_5932_42308# 9.2e-19
C12477 a_13747_46662# a_21356_42826# 1.41e-19
C12478 a_19321_45002# a_19987_42826# 5.73e-20
C12479 a_n2017_45002# a_18494_42460# 0.002888f
C12480 a_n1059_45260# a_18184_42460# 0.52106f
C12481 a_n1613_43370# a_n1545_46494# 1.79e-19
C12482 a_15227_44166# a_19333_46634# 0.065741f
C12483 a_2747_46873# a_526_44458# 5.38e-20
C12484 a_n2661_46634# a_9290_44172# 2.69e-19
C12485 a_1239_47204# a_n755_45592# 4.63e-21
C12486 a_n2661_46098# a_167_45260# 1.31e-19
C12487 a_2609_46660# a_1823_45246# 3.24e-19
C12488 a_n1925_46634# a_5937_45572# 6.05e-20
C12489 a_4646_46812# a_n2293_46098# 1.72e-21
C12490 a_3785_47178# a_n2661_45546# 8.89e-21
C12491 a_13381_47204# a_13259_45724# 4.87e-21
C12492 a_4883_46098# a_8062_46482# 6.26e-20
C12493 a_10227_46804# a_10586_45546# 0.306536f
C12494 a_n2497_47436# a_2277_45546# 8.01e-22
C12495 a_n971_45724# a_n356_45724# 0.030873f
C12496 a_n237_47217# a_3316_45546# 1.38e-19
C12497 a_584_46384# a_n1099_45572# 0.021537f
C12498 a_2107_46812# a_4704_46090# 0.008508f
C12499 a_n1151_42308# a_n2956_38216# 4.1e-20
C12500 a_n881_46662# a_n1736_46482# 1.29e-19
C12501 a_17609_46634# a_19692_46634# 3.12e-20
C12502 a_13747_46662# a_14275_46494# 0.002369f
C12503 a_13661_43548# a_15015_46420# 0.001123f
C12504 a_5807_45002# a_14840_46494# 8.3e-21
C12505 a_n743_46660# a_8349_46414# 0.004029f
C12506 a_n97_42460# a_13921_42308# 0.003369f
C12507 a_2905_42968# a_3059_42968# 0.008678f
C12508 a_17730_32519# a_22521_39511# 1.16e-20
C12509 a_19319_43548# a_19647_42308# 1.57e-21
C12510 a_3626_43646# a_10533_42308# 0.002711f
C12511 a_2982_43646# a_11323_42473# 1.02e-19
C12512 a_5342_30871# a_15567_42826# 0.024331f
C12513 a_4190_30871# a_18695_43230# 1.55e-19
C12514 a_19237_31679# a_22459_39145# 1.6e-20
C12515 a_4361_42308# a_13291_42460# 0.029279f
C12516 a_8103_44636# a_8975_43940# 1.09e-20
C12517 a_20107_45572# a_19862_44208# 4.31e-20
C12518 a_4558_45348# a_3905_42865# 9.27e-19
C12519 a_3537_45260# a_5013_44260# 0.001173f
C12520 a_n2017_45002# a_3499_42826# 4.96e-19
C12521 a_10903_43370# a_13113_42826# 0.011891f
C12522 a_n357_42282# a_14358_43442# 3e-20
C12523 a_n443_42852# a_5837_43396# 2.02e-19
C12524 a_n2442_46660# a_7174_31319# 5.91e-21
C12525 a_n2433_44484# a_n1809_44850# 9.73e-19
C12526 a_n2661_44458# a_n1190_44850# 1.42e-19
C12527 a_5147_45002# a_3600_43914# 7.58e-20
C12528 a_16375_45002# a_17324_43396# 1.24e-20
C12529 a_n1925_42282# a_n1423_42826# 1.97e-20
C12530 a_n2129_44697# a_n2012_44484# 0.172424f
C12531 a_4185_45028# a_21195_42852# 2.22e-20
C12532 a_9290_44172# a_14543_43071# 0.005728f
C12533 a_11031_47542# a_413_45260# 1.03e-19
C12534 a_n881_46662# a_18175_45572# 1.17e-19
C12535 a_n2293_46098# a_n1545_46494# 4.26e-19
C12536 a_4646_46812# a_7230_45938# 0.005389f
C12537 a_2063_45854# a_10775_45002# 0.012226f
C12538 a_13747_46662# a_15765_45572# 0.5661f
C12539 a_9625_46129# a_9569_46155# 0.204034f
C12540 a_n1151_42308# a_7229_43940# 0.036511f
C12541 a_13885_46660# a_14383_46116# 2.54e-21
C12542 a_13059_46348# a_14180_46482# 0.025233f
C12543 a_20990_47178# a_2437_43646# 0.008979f
C12544 a_19386_47436# a_3357_43084# 4.09e-19
C12545 a_5257_43370# a_6511_45714# 9.68e-20
C12546 a_8492_46660# a_2711_45572# 8.18e-21
C12547 a_n1853_46287# a_n2956_38680# 6.64e-19
C12548 a_n1991_46122# a_n2956_39304# 2.14e-20
C12549 a_3090_45724# a_n2661_45546# 0.561435f
C12550 a_19692_46634# a_19443_46116# 1.33e-19
C12551 a_n443_46116# a_4927_45028# 5.42e-19
C12552 a_8953_45546# a_9823_46155# 6.18e-19
C12553 a_8199_44636# a_9290_44172# 0.516297f
C12554 a_3483_46348# a_2324_44458# 0.668551f
C12555 a_n2157_46122# a_n1736_46482# 0.086708f
C12556 a_13661_43548# a_16333_45814# 8.09e-19
C12557 a_20107_46660# a_8049_45260# 5.25e-21
C12558 a_12549_44172# a_13297_45572# 5.89e-19
C12559 a_12891_46348# a_13385_45572# 0.001139f
C12560 a_4791_45118# a_5691_45260# 0.001279f
C12561 a_15227_44166# a_20062_46116# 1.82e-19
C12562 a_n2497_47436# a_626_44172# 0.249352f
C12563 a_1209_43370# VDD 0.191694f
C12564 a_20922_43172# a_17303_42282# 1.39e-20
C12565 a_18249_42858# a_18214_42558# 2.84e-19
C12566 a_18599_43230# a_18907_42674# 0.001393f
C12567 a_n1329_42308# a_n961_42308# 0.001982f
C12568 COMP_P a_n473_42460# 1.25e-19
C12569 a_n1736_42282# a_n784_42308# 2.19e-19
C12570 a_n2104_42282# a_n3674_37592# 0.006157f
C12571 a_n2472_42282# a_n1630_35242# 0.040716f
C12572 a_3080_42308# C5_N_btm 3.03e-19
C12573 a_8375_44464# a_8333_44056# 2.14e-19
C12574 a_5891_43370# a_8018_44260# 8.02e-19
C12575 a_19279_43940# a_20512_43084# 1.32e-19
C12576 a_n2956_38216# a_n2840_42282# 2.12e-20
C12577 a_18989_43940# a_19478_44306# 1.12e-19
C12578 a_21005_45260# a_20974_43370# 3.69e-20
C12579 a_21359_45002# a_21381_43940# 5.38e-20
C12580 a_n2661_43922# a_n1287_44306# 5.84e-19
C12581 a_n2661_42834# a_n875_44318# 1.15e-19
C12582 a_8696_44636# a_9127_43156# 6.2e-21
C12583 a_n357_42282# a_20836_43172# 9.04e-20
C12584 a_n2810_45572# a_n4318_38216# 0.023144f
C12585 a_20205_31679# COMP_P 3.65e-20
C12586 a_20679_44626# a_17730_32519# 3.62e-21
C12587 a_16979_44734# a_11341_43940# 5.51e-20
C12588 a_16112_44458# a_15493_43940# 4.79e-19
C12589 a_8953_45002# a_9885_43646# 1.33e-20
C12590 a_11691_44458# a_19319_43548# 4.59e-19
C12591 a_13556_45296# a_9145_43396# 5.5e-21
C12592 a_9482_43914# a_9803_43646# 9.27e-20
C12593 a_13059_46348# a_n1059_45260# 2.69e-20
C12594 a_16327_47482# a_9313_44734# 0.169217f
C12595 a_n1925_42282# a_3775_45552# 2.95e-21
C12596 a_14840_46494# a_15143_45578# 1.28e-19
C12597 a_526_44458# a_3638_45822# 3.45e-19
C12598 a_19551_46910# a_3357_43084# 5.32e-20
C12599 a_2324_44458# a_14495_45572# 0.00152f
C12600 a_768_44030# a_n699_43396# 1.37533f
C12601 a_3090_45724# a_5205_44484# 0.005908f
C12602 a_11415_45002# a_17568_45572# 9.66e-19
C12603 a_20273_46660# a_2437_43646# 4.41e-20
C12604 a_11735_46660# a_11963_45334# 1.91e-21
C12605 a_11813_46116# a_11787_45002# 1.43e-19
C12606 a_8199_44636# a_11064_45572# 7.43e-21
C12607 a_15368_46634# a_6171_45002# 1.38e-19
C12608 a_6945_45028# a_10193_42453# 9.46e-20
C12609 a_10903_43370# a_10907_45822# 0.199567f
C12610 a_5066_45546# a_5263_45724# 0.022243f
C12611 a_n1630_35242# a_3754_38470# 9.47e-20
C12612 a_19511_42282# a_21887_42336# 2.03e-19
C12613 a_n4318_37592# a_n4064_37440# 0.04779f
C12614 a_5932_42308# a_n4064_37984# 0.003117f
C12615 a_3059_42968# VDD 8.13e-19
C12616 a_20107_42308# a_20712_42282# 0.008f
C12617 a_13258_32519# a_7174_31319# 0.02542f
C12618 a_5742_30871# comp_n 1.22e-19
C12619 a_10807_43548# a_11257_43940# 0.013221f
C12620 a_11691_44458# a_16795_42852# 1.42e-19
C12621 a_11967_42832# a_13667_43396# 6.68e-20
C12622 a_n913_45002# a_2713_42308# 0.291963f
C12623 a_n1059_45260# a_2903_42308# 0.003187f
C12624 a_n2017_45002# a_3318_42354# 0.01513f
C12625 a_6945_45028# VDD 1.30257f
C12626 a_11827_44484# a_17333_42852# 3.3e-21
C12627 a_n2293_42834# a_5193_42852# 2.39e-20
C12628 a_2998_44172# a_4235_43370# 2.06e-20
C12629 a_3600_43914# a_4093_43548# 4.01e-19
C12630 a_18494_42460# a_19164_43230# 5.14e-19
C12631 a_18184_42460# a_19987_42826# 0.208392f
C12632 a_n2956_38680# a_n2661_43370# 2.4e-20
C12633 a_17715_44484# a_16922_45042# 0.039816f
C12634 a_167_45260# a_742_44458# 9.2e-20
C12635 a_n2293_46634# a_10405_44172# 0.002468f
C12636 a_16327_47482# a_20974_43370# 0.004018f
C12637 a_8049_45260# a_1423_45028# 1.12e-19
C12638 a_13904_45546# a_8696_44636# 5.54e-21
C12639 a_10907_45822# a_12016_45572# 3.47e-20
C12640 a_1823_45246# a_2779_44458# 0.00892f
C12641 a_2202_46116# a_949_44458# 7.07e-21
C12642 a_11415_45002# a_17767_44458# 4.21e-20
C12643 a_12741_44636# a_16112_44458# 0.019518f
C12644 a_n2661_45546# a_2274_45254# 0.002096f
C12645 a_n2293_45546# a_413_45260# 0.066602f
C12646 a_13661_43548# a_15493_43396# 0.491785f
C12647 a_11823_42460# a_16223_45938# 3.12e-20
C12648 a_n452_45724# a_n467_45028# 0.001128f
C12649 a_n863_45724# a_n143_45144# 0.033306f
C12650 a_n357_42282# en_comp 2.96e-20
C12651 a_12427_45724# a_12561_45572# 0.001089f
C12652 a_4791_45118# a_3080_42308# 1.96e-19
C12653 a_n443_46116# a_4699_43561# 9.16e-21
C12654 a_10586_45546# a_1307_43914# 1.48e-20
C12655 a_12839_46116# a_13017_45260# 5.04e-21
C12656 a_5807_45002# a_19478_44306# 0.001092f
C12657 a_n4334_37440# a_n4064_37440# 0.448688f
C12658 a_n3690_37440# a_n3420_37440# 0.431074f
C12659 a_n3565_37414# a_n2946_37690# 0.407439f
C12660 a_n4209_37414# a_n2302_37690# 0.407594f
C12661 VDAC_Ni a_4338_37500# 0.640521f
C12662 a_7754_38636# a_5088_37509# 0.288061f
C12663 a_n4064_40160# VCM 0.121302f
C12664 a_n4209_39590# VIN_P 0.105382f
C12665 a_n1741_47186# a_10467_46802# 9.36e-19
C12666 a_n971_45724# a_8667_46634# 0.006462f
C12667 a_n237_47217# a_8145_46902# 3.42e-20
C12668 a_4700_47436# a_4651_46660# 4.72e-19
C12669 a_n443_46116# a_3877_44458# 0.06318f
C12670 a_4791_45118# a_4646_46812# 0.485113f
C12671 a_n3607_39616# VDD 2.79e-20
C12672 a_n3565_38502# C5_P_btm 0.00105f
C12673 a_n3420_38528# C7_P_btm 7.66e-20
C12674 a_10227_46804# a_n743_46660# 0.134234f
C12675 a_7754_38968# a_8912_37509# 6.06e-19
C12676 a_n881_46662# a_8128_46384# 0.206292f
C12677 a_4883_46098# a_21588_30879# 4.72e-19
C12678 a_21811_47423# a_20916_46384# 0.109084f
C12679 a_19319_43548# a_4190_30871# 0.188868f
C12680 en_comp CAL_N 0.024527f
C12681 a_19963_31679# a_22609_37990# 8.31e-21
C12682 a_3905_42865# a_5193_43172# 8.11e-19
C12683 a_7287_43370# a_7466_43396# 0.007399f
C12684 a_n97_42460# a_18525_43370# 0.005868f
C12685 a_8696_44636# CLK 0.006002f
C12686 a_8147_43396# a_8685_43396# 0.077232f
C12687 a_7112_43396# a_7221_43396# 0.007416f
C12688 a_10949_43914# a_5534_30871# 2.43e-20
C12689 a_20447_31679# a_22609_38406# 4.44e-21
C12690 a_n863_45724# a_n2293_43922# 7.65e-20
C12691 a_8696_44636# a_17023_45118# 0.064781f
C12692 a_15861_45028# a_16922_45042# 0.259169f
C12693 a_4558_45348# a_5147_45002# 0.09356f
C12694 a_3065_45002# a_3232_43370# 0.049451f
C12695 a_22612_30879# a_13678_32519# 0.060546f
C12696 a_n443_42852# a_8375_44464# 6.71e-19
C12697 a_n913_45002# a_9482_43914# 8.96e-20
C12698 a_3537_45260# a_4927_45028# 0.216859f
C12699 a_4574_45260# a_5111_44636# 1.69e-19
C12700 a_16327_47482# a_18599_43230# 0.182696f
C12701 a_2437_43646# a_2304_45348# 0.006164f
C12702 a_8199_44636# a_10807_43548# 6.84e-21
C12703 a_9049_44484# a_9838_44484# 8.16e-19
C12704 a_7499_43078# a_10157_44484# 4.34e-20
C12705 a_380_45546# a_n2661_42834# 3.2e-21
C12706 a_2063_45854# a_526_44458# 0.039908f
C12707 a_584_46384# a_n1925_42282# 0.194054f
C12708 a_6151_47436# a_10809_44734# 5.72e-19
C12709 a_6491_46660# a_6945_45028# 0.0023f
C12710 a_13717_47436# a_17583_46090# 1.18e-21
C12711 a_12861_44030# a_15682_46116# 0.030474f
C12712 a_13661_43548# a_18900_46660# 0.003751f
C12713 a_n881_46662# a_n1641_46494# 4.9e-19
C12714 a_n1613_43370# a_n901_46420# 0.406381f
C12715 a_4883_46098# a_6419_46155# 0.007342f
C12716 a_11599_46634# a_14275_46494# 0.029786f
C12717 a_10227_46804# a_11189_46129# 0.001224f
C12718 a_14955_47212# a_15015_46420# 4.84e-19
C12719 a_n1741_47186# a_8034_45724# 3.32e-21
C12720 a_8145_46902# a_8270_45546# 4.35e-20
C12721 a_8492_46660# a_8654_47026# 0.006453f
C12722 a_7927_46660# a_8189_46660# 0.001705f
C12723 a_2747_46873# a_2521_46116# 7.97e-20
C12724 a_n743_46660# a_17339_46660# 2.36e-19
C12725 a_n237_47217# a_5066_45546# 1.48406f
C12726 a_5649_42852# a_13113_42826# 3.48e-21
C12727 a_n1557_42282# a_n4318_38216# 2.95e-20
C12728 a_n3674_39768# a_n4064_39616# 0.464693f
C12729 a_18079_43940# a_18057_42282# 3.16e-21
C12730 a_8103_44636# VDD 0.124028f
C12731 a_743_42282# a_15567_42826# 7.68e-20
C12732 a_4190_30871# a_16795_42852# 3.12e-21
C12733 a_1209_43370# a_n784_42308# 3.67e-21
C12734 a_n2293_46634# a_6171_42473# 2.55e-21
C12735 a_n2442_46660# a_5932_42308# 5.39e-21
C12736 a_11823_42460# a_11341_43940# 0.087329f
C12737 a_n755_45592# a_n2267_43396# 2.31e-20
C12738 a_n357_42282# a_n1699_43638# 4.63e-20
C12739 a_n2661_43370# a_10334_44484# 7.92e-20
C12740 a_13259_45724# a_3626_43646# 0.037016f
C12741 a_21005_45260# a_18114_32519# 6.8e-20
C12742 a_10775_45002# a_n2661_42834# 1.02e-20
C12743 a_8953_45002# a_n2661_43922# 5.04e-19
C12744 a_22223_45572# a_3422_30871# 2.45e-20
C12745 a_17715_44484# a_15743_43084# 1.72e-19
C12746 a_18597_46090# a_20712_42282# 8.69e-19
C12747 a_1423_45028# a_5289_44734# 0.002441f
C12748 a_14537_43396# a_9313_44734# 1.05e-20
C12749 a_n863_45724# a_n97_42460# 0.581863f
C12750 a_4883_46098# a_10907_45822# 1.59e-21
C12751 a_8270_45546# a_5066_45546# 0.189476f
C12752 a_13059_46348# a_13925_46122# 0.056739f
C12753 a_14513_46634# a_2324_44458# 1.3e-19
C12754 a_n1853_46287# a_n1423_46090# 0.043126f
C12755 a_n2109_47186# a_2437_43646# 0.027184f
C12756 a_2107_46812# a_2957_45546# 1.23e-20
C12757 a_n1925_46634# a_n443_42852# 5.96e-20
C12758 a_n2661_46098# a_n863_45724# 4.3e-20
C12759 a_3699_46634# a_n2661_45546# 5.3e-21
C12760 a_n2293_46098# a_n901_46420# 0.007523f
C12761 a_n2157_46122# a_n1641_46494# 0.105995f
C12762 a_n881_46662# a_10053_45546# 4.53e-21
C12763 a_8128_46384# a_8162_45546# 2.64e-19
C12764 a_765_45546# a_9290_44172# 4.14e-20
C12765 a_19466_46812# a_10809_44734# 0.007455f
C12766 a_19692_46634# a_22223_46124# 0.001994f
C12767 a_10249_46116# a_10044_46482# 0.00124f
C12768 a_10467_46802# a_10586_45546# 5.92e-20
C12769 a_5807_45002# a_6511_45714# 0.012932f
C12770 a_11599_46634# a_15765_45572# 0.001673f
C12771 a_n2293_42282# a_1606_42308# 0.192228f
C12772 a_21487_43396# a_13258_32519# 9.88e-21
C12773 a_743_42282# a_20712_42282# 0.001163f
C12774 a_13467_32519# a_19511_42282# 0.003538f
C12775 a_4361_42308# a_18548_42308# 5.09e-19
C12776 a_17538_32519# a_22521_39511# 1.06e-20
C12777 a_11173_44260# VDD 0.005546f
C12778 a_10083_42826# a_9803_42558# 0.006054f
C12779 a_3094_47570# DATA[2] 6.24e-20
C12780 a_n2017_45002# a_6197_43396# 4.71e-20
C12781 a_4185_45028# a_8791_42308# 1.64e-19
C12782 a_3065_45002# a_4905_42826# 2.38e-20
C12783 a_5883_43914# a_5244_44056# 1.47e-19
C12784 a_3315_47570# DATA[1] 1.79e-21
C12785 a_3357_43084# a_3457_43396# 5.15e-19
C12786 a_n357_42282# a_22165_42308# 1.25e-19
C12787 a_n2956_38680# COMP_P 0.001147f
C12788 a_n2956_39304# a_n1329_42308# 6.85e-20
C12789 a_16922_45042# a_20623_43914# 0.001335f
C12790 a_4558_45348# a_4093_43548# 9.14e-21
C12791 a_15146_44811# a_14673_44172# 0.001224f
C12792 a_9313_44734# a_20835_44721# 4.17e-21
C12793 a_5343_44458# a_7281_43914# 8.75e-20
C12794 a_n967_45348# a_n998_43396# 4.97e-19
C12795 a_11691_44458# a_10949_43914# 4.22e-20
C12796 a_3411_47243# VDD 2.18e-20
C12797 a_n1059_45260# a_6293_42852# 0.002519f
C12798 a_n913_45002# a_6031_43396# 2.91e-20
C12799 a_11827_44484# a_13483_43940# 5.96e-19
C12800 a_3537_45260# a_4699_43561# 0.024682f
C12801 a_15861_45028# a_15743_43084# 1.08e-20
C12802 a_11453_44696# a_19778_44110# 8.76e-20
C12803 a_n2293_46634# a_1145_45348# 1.48e-19
C12804 a_10809_44734# a_20205_31679# 0.039075f
C12805 a_22223_46124# a_20692_30879# 2.55e-19
C12806 a_n971_45724# a_n356_44636# 1.4e-19
C12807 a_3877_44458# a_3537_45260# 0.12249f
C12808 a_14035_46660# a_8696_44636# 6.34e-21
C12809 a_4883_46098# a_21359_45002# 5.09e-22
C12810 a_16327_47482# a_18114_32519# 5.2e-20
C12811 a_2324_44458# a_n357_42282# 1.23e-19
C12812 a_2107_46812# a_9482_43914# 0.109711f
C12813 a_5068_46348# a_5263_45724# 2.95e-19
C12814 a_5732_46660# a_413_45260# 8.11e-21
C12815 a_13059_46348# a_15599_45572# 5.07e-19
C12816 a_6969_46634# a_3357_43084# 3.01e-20
C12817 a_3090_45724# a_19431_45546# 4.09e-21
C12818 a_13507_46334# a_22223_45036# 0.005873f
C12819 a_6151_47436# a_5883_43914# 8.07e-21
C12820 a_4419_46090# a_6194_45824# 7.7e-20
C12821 a_3483_46348# a_6667_45809# 3.14e-22
C12822 a_5497_46414# a_2711_45572# 0.001047f
C12823 a_n743_46660# a_1307_43914# 0.002676f
C12824 a_14456_42282# a_15803_42450# 5.2e-21
C12825 a_n4318_37592# a_n3420_39072# 0.02033f
C12826 a_5742_30871# a_11633_42308# 0.001223f
C12827 a_n3674_38216# a_n4064_39072# 0.019725f
C12828 a_22165_42308# CAL_N 8.8e-21
C12829 a_5932_42308# a_13258_32519# 5.13e-19
C12830 a_n722_43218# VDD 1.22e-19
C12831 a_20193_45348# a_21487_43396# 5.6e-20
C12832 a_n2293_42834# a_7227_42852# 0.008564f
C12833 a_11823_42460# a_10723_42308# 3.49e-19
C12834 a_16979_44734# a_10341_43396# 8.24e-21
C12835 a_n2956_38216# a_n2302_39866# 3.61e-19
C12836 a_n2472_46090# VDD 0.224658f
C12837 a_1467_44172# a_1241_43940# 0.011879f
C12838 a_1115_44172# a_1443_43940# 0.096132f
C12839 a_22365_46825# EN_OFFSET_CAL 0.195393f
C12840 a_9672_43914# a_10405_44172# 4.63e-19
C12841 a_5891_43370# a_6452_43396# 1.68e-20
C12842 a_18579_44172# a_19478_44056# 2.74e-19
C12843 a_20835_44721# a_20974_43370# 5.58e-21
C12844 a_n2956_38680# a_n3565_37414# 9.9e-21
C12845 a_n1059_45260# a_11554_42852# 0.002165f
C12846 a_2711_45572# a_18907_42674# 2.61e-19
C12847 a_10193_42453# a_14456_42282# 0.001037f
C12848 a_16327_47482# a_17737_43940# 3e-21
C12849 a_6194_45824# a_6469_45572# 0.007416f
C12850 a_5164_46348# a_5365_45348# 5.46e-19
C12851 a_8568_45546# a_9049_44484# 4.21e-19
C12852 a_1138_42852# a_n2293_42834# 0.015752f
C12853 a_n881_46662# a_5244_44056# 1.42e-21
C12854 a_12861_44030# a_20269_44172# 0.047709f
C12855 a_584_46384# a_3737_43940# 8.18e-19
C12856 a_2711_45572# a_9241_45822# 1.37e-19
C12857 a_8953_45546# a_1423_45028# 0.021907f
C12858 a_11415_45002# a_16405_45348# 9.91e-19
C12859 a_13259_45724# a_17568_45572# 0.005159f
C12860 a_21188_46660# a_21359_45002# 4.5e-21
C12861 a_20731_47026# a_20567_45036# 2.2e-21
C12862 a_8049_45260# a_22591_45572# 0.036446f
C12863 a_768_44030# a_1467_44172# 0.022755f
C12864 a_2324_44458# a_11963_45334# 0.001724f
C12865 a_13759_46122# a_13777_45326# 9.69e-19
C12866 a_13925_46122# a_13556_45296# 2.8e-21
C12867 a_16327_47482# a_12465_44636# 6.07e-19
C12868 a_10227_46804# a_21177_47436# 9.07e-19
C12869 a_17591_47464# a_13507_46334# 3.36e-20
C12870 a_n4209_39304# a_n2946_37690# 2.26e-19
C12871 a_n3565_38216# a_n2216_37984# 0.003076f
C12872 a_14456_42282# VDD 0.265543f
C12873 a_16763_47508# a_4883_46098# 8.86e-22
C12874 a_1736_39043# VDAC_Ni 5.86e-19
C12875 a_n3565_39304# a_n3690_37440# 2.75e-19
C12876 a_n3420_39072# a_n4334_37440# 2.36e-19
C12877 a_4958_30871# C10_P_btm 6.95e-19
C12878 a_n4064_37984# a_n4251_38304# 4.37e-19
C12879 a_22465_38105# a_22521_39511# 0.902378f
C12880 a_6545_47178# a_n1613_43370# 0.006198f
C12881 a_18597_46090# a_19386_47436# 0.007892f
C12882 a_18780_47178# a_19787_47423# 2.54e-20
C12883 a_6151_47436# a_n881_46662# 1.58776f
C12884 a_18479_47436# a_20894_47436# 0.032517f
C12885 a_4915_47217# a_5159_47243# 7.22e-19
C12886 a_n1151_42308# a_768_44030# 0.019901f
C12887 a_n1920_47178# a_n2956_39768# 6.13e-19
C12888 a_n2109_47186# a_n2661_46634# 0.038259f
C12889 a_n2288_47178# a_n2472_46634# 3.21e-19
C12890 a_n2497_47436# a_n2442_46660# 0.045496f
C12891 a_n4318_39768# a_n3674_39304# 0.024426f
C12892 a_2479_44172# a_3681_42891# 1.73e-19
C12893 a_19279_43940# a_18249_42858# 5.33e-20
C12894 a_n2956_37592# a_n3420_38528# 6.26e-20
C12895 a_6812_45938# VDD 0.132317f
C12896 a_10405_44172# a_743_42282# 1.09e-20
C12897 a_2675_43914# a_2075_43172# 3.57e-20
C12898 a_2889_44172# a_1847_42826# 6.94e-19
C12899 a_9313_44734# a_12991_43230# 2.5e-19
C12900 a_20623_43914# a_15743_43084# 1.72e-20
C12901 a_15493_43940# a_17499_43370# 2.64e-19
C12902 a_11341_43940# a_18429_43548# 2.54e-20
C12903 a_n97_42460# a_3540_43646# 0.027089f
C12904 a_3422_30871# a_5534_30871# 0.023427f
C12905 a_14021_43940# a_14537_43646# 0.001553f
C12906 a_n2661_42282# a_5649_42852# 0.052118f
C12907 a_n1099_45572# a_n1177_44458# 2.8e-19
C12908 a_15599_45572# a_13556_45296# 7.13e-22
C12909 a_n2293_46634# a_3457_43396# 8.01e-19
C12910 a_n2293_46098# a_5013_44260# 0.040459f
C12911 a_19479_31679# a_22591_45572# 0.011797f
C12912 a_12549_44172# a_12281_43396# 0.004094f
C12913 a_526_44458# a_n2661_42834# 0.06021f
C12914 a_n452_45724# a_n452_44636# 6.69e-19
C12915 a_19335_46494# a_17517_44484# 2.71e-21
C12916 a_16375_45002# a_16112_44458# 4.06e-20
C12917 a_13259_45724# a_17767_44458# 0.026768f
C12918 a_n863_45724# a_742_44458# 0.629795f
C12919 a_9049_44484# a_n2661_43370# 0.030026f
C12920 a_18597_46090# a_20556_43646# 1.94e-19
C12921 a_1138_42852# a_1115_44172# 0.012127f
C12922 a_21513_45002# a_20447_31679# 4.16e-20
C12923 a_n443_46116# a_1847_42826# 0.00118f
C12924 a_22223_45572# a_19963_31679# 0.00254f
C12925 a_10227_46804# a_4361_42308# 0.073929f
C12926 a_n2661_45546# a_4743_44484# 0.004404f
C12927 a_8696_44636# a_10951_45334# 0.001322f
C12928 a_15037_45618# a_14537_43396# 3.1e-20
C12929 a_2957_45546# a_n2661_44458# 5.79e-21
C12930 a_3090_45724# a_15301_44260# 9.33e-19
C12931 a_8270_45546# a_8415_44056# 1.57e-19
C12932 a_2107_46812# a_7715_46873# 0.032178f
C12933 a_2905_45572# a_1823_45246# 1.3e-19
C12934 a_12549_44172# a_15009_46634# 0.009008f
C12935 a_768_44030# a_14084_46812# 0.013767f
C12936 a_12891_46348# a_3090_45724# 1.19e-21
C12937 C8_P_btm VREF 3.6701f
C12938 a_10227_46804# a_20841_46902# 0.164019f
C12939 C9_P_btm VREF_GND 5.18245f
C12940 a_n237_47217# a_5068_46348# 0.033474f
C12941 a_n971_45724# a_5204_45822# 4.32e-20
C12942 a_n1741_47186# a_8016_46348# 3.91e-20
C12943 a_n1151_42308# a_1176_45822# 1.53e-19
C12944 C6_N_btm C10_N_btm 0.421276f
C12945 C7_N_btm C9_N_btm 0.227839f
C12946 a_13507_46334# a_15312_46660# 5.88e-21
C12947 a_3524_46660# a_4817_46660# 1.33e-19
C12948 C4_N_btm VDD 0.265463f
C12949 C10_P_btm VCM 10.3108f
C12950 a_18479_47436# a_20411_46873# 0.192791f
C12951 C6_P_btm VIN_P 0.391898f
C12952 a_584_46384# a_2698_46116# 1.53e-19
C12953 a_2063_45854# a_2521_46116# 0.011365f
C12954 a_n743_46660# a_10467_46802# 9.14e-20
C12955 a_3539_42460# a_n2293_42282# 0.010651f
C12956 a_4190_30871# a_19095_43396# 0.046015f
C12957 a_743_42282# a_20556_43646# 0.028541f
C12958 a_10695_43548# a_10835_43094# 5.89e-20
C12959 a_19721_31679# a_22521_39511# 2.63e-20
C12960 a_7735_45067# VDD 2.18e-20
C12961 a_16823_43084# a_5649_42852# 6.08e-21
C12962 a_3422_30871# a_19647_42308# 6.32e-20
C12963 a_n97_42460# a_7309_42852# 0.024142f
C12964 a_13661_43548# a_18707_42852# 1.38e-19
C12965 a_n357_42282# a_19862_44208# 0.138067f
C12966 a_n1925_42282# a_n1177_43370# 1.62e-22
C12967 a_3232_43370# a_6298_44484# 0.256727f
C12968 a_7229_43940# a_4223_44672# 0.014299f
C12969 a_n443_42852# a_10949_43914# 3.54e-20
C12970 a_n2293_45010# a_n356_44636# 0.031375f
C12971 a_n2017_45002# a_n1821_44484# 0.001578f
C12972 a_3357_43084# a_5826_44734# 2.81e-19
C12973 a_17339_46660# a_4361_42308# 3.78e-20
C12974 a_5111_44636# a_5883_43914# 0.281106f
C12975 a_16333_45814# a_11967_42832# 2.46e-21
C12976 a_8696_44636# a_17061_44484# 3.53e-19
C12977 a_6755_46942# a_15567_42826# 7.16e-21
C12978 a_3090_45724# a_4520_42826# 2.44e-19
C12979 a_5205_44484# a_4743_44484# 8.65e-19
C12980 a_9482_43914# a_n2661_44458# 0.017706f
C12981 a_n743_46660# a_8034_45724# 0.021079f
C12982 a_n971_45724# a_8697_45822# 0.002809f
C12983 a_6755_46942# a_9569_46155# 1.96e-19
C12984 a_6491_46660# a_6812_45938# 1.44e-21
C12985 a_6151_47436# a_8162_45546# 6.52e-20
C12986 a_4915_47217# a_9049_44484# 1.19e-20
C12987 a_4646_46812# a_6945_45028# 0.090679f
C12988 a_n2661_46098# a_1431_46436# 2.82e-19
C12989 a_2107_46812# a_5210_46482# 8.98e-19
C12990 a_16327_47482# a_2711_45572# 0.101699f
C12991 a_n1151_42308# a_11652_45724# 4.93e-20
C12992 a_10428_46928# a_11133_46155# 6.41e-19
C12993 a_10467_46802# a_11189_46129# 0.005012f
C12994 a_10249_46116# a_9823_46155# 0.082191f
C12995 a_10623_46897# a_9290_44172# 0.00174f
C12996 a_4361_42308# a_4933_42558# 4.55e-21
C12997 a_743_42282# a_6171_42473# 0.007484f
C12998 a_15567_42826# a_16328_43172# 1.3e-20
C12999 a_15781_43660# a_14113_42308# 2.97e-21
C13000 a_15681_43442# a_15051_42282# 1.21e-19
C13001 a_13460_43230# a_13622_42852# 0.006453f
C13002 a_895_43940# VDD 0.318652f
C13003 a_15227_44166# a_14113_42308# 4.65e-20
C13004 a_10057_43914# a_10809_44484# 2.31e-19
C13005 a_4700_47436# VDD 0.086132f
C13006 a_1423_45028# a_9028_43914# 7.39e-20
C13007 a_2905_45572# DATA[2] 5.19e-19
C13008 a_n863_45724# a_n901_43156# 1.75e-19
C13009 a_526_44458# a_n2293_42282# 0.010969f
C13010 a_9290_44172# a_13291_42460# 0.078684f
C13011 a_11823_42460# a_10341_43396# 0.088285f
C13012 a_13249_42308# a_14358_43442# 1.53e-20
C13013 a_n1151_42308# DATA[0] 0.088597f
C13014 a_3160_47472# DATA[1] 8.03e-22
C13015 a_11827_44484# a_21073_44484# 7.17e-19
C13016 a_n357_42282# a_n2157_42858# 1.01e-19
C13017 a_21076_30879# a_n1630_35242# 0.034943f
C13018 a_2063_45854# DATA[5] 0.001488f
C13019 a_n2956_38216# a_n3674_39304# 0.023342f
C13020 a_18114_32519# a_20835_44721# 9.39e-20
C13021 a_1307_43914# a_11750_44172# 0.007207f
C13022 a_n2661_43370# a_3905_42865# 6.49e-20
C13023 a_n356_44636# a_9313_44734# 2.11e-20
C13024 a_13720_44458# a_14112_44734# 0.016359f
C13025 SMPL_ON_N a_22459_39145# 0.00803f
C13026 a_8016_46348# a_10586_45546# 2.29e-19
C13027 a_n1925_46634# a_2437_43646# 0.02753f
C13028 a_n2293_46634# a_3357_43084# 0.963711f
C13029 a_4883_46098# a_15415_45028# 1.77e-20
C13030 a_9569_46155# a_8049_45260# 0.009377f
C13031 a_n881_46662# a_5111_44636# 0.00608f
C13032 a_n1613_43370# a_4927_45028# 6.4e-22
C13033 a_11453_44696# a_9482_43914# 0.042575f
C13034 a_12465_44636# a_14537_43396# 0.031033f
C13035 a_8128_46384# a_3537_45260# 0.001708f
C13036 a_768_44030# a_327_44734# 0.00311f
C13037 a_10467_46802# a_11136_45572# 1.63e-20
C13038 a_5379_42460# a_5934_30871# 5.78e-20
C13039 a_n784_42308# a_14456_42282# 3.86e-20
C13040 a_1576_42282# a_5742_30871# 2.87e-20
C13041 a_5755_42308# a_6171_42473# 0.017801f
C13042 a_5421_42558# a_5932_42308# 6.5e-19
C13043 a_3823_42558# a_3905_42308# 0.003935f
C13044 a_n443_42852# a_6481_42558# 0.001736f
C13045 a_n2956_38680# a_n4209_39304# 0.021073f
C13046 a_n2956_39304# a_n4334_39392# 6.77e-20
C13047 a_15559_46634# VDD 0.301657f
C13048 a_n2661_44458# a_6031_43396# 5.36e-21
C13049 a_n1899_43946# a_n1441_43940# 0.03441f
C13050 a_11967_42832# a_15493_43396# 0.02628f
C13051 a_19615_44636# a_19328_44172# 3.27e-21
C13052 a_2998_44172# a_3905_42865# 3.52e-19
C13053 a_15368_46634# RST_Z 3.47e-20
C13054 a_1307_43914# a_4361_42308# 7.03e-21
C13055 a_n913_45002# a_10796_42968# 0.545674f
C13056 a_n1059_45260# a_10991_42826# 0.004257f
C13057 a_n2017_45002# a_10922_42852# 1.02e-20
C13058 a_13259_45724# a_13921_42308# 9.76e-19
C13059 a_16979_44734# a_n97_42460# 1.23e-21
C13060 a_2779_44458# a_2896_43646# 6.83e-21
C13061 a_742_44458# a_3540_43646# 1.09e-20
C13062 a_2382_45260# a_3935_42891# 0.061675f
C13063 a_11813_46116# CLK 2.07e-20
C13064 a_n357_42282# a_9803_42558# 4.98e-21
C13065 a_n755_45592# a_9223_42460# 1.28e-19
C13066 a_n699_43396# a_1891_43646# 4.33e-19
C13067 a_13259_45724# a_12791_45546# 0.001427f
C13068 a_768_44030# a_13857_44734# 0.011246f
C13069 a_4791_45118# a_5013_44260# 0.02062f
C13070 a_4646_46812# a_8103_44636# 0.002138f
C13071 a_n2661_45546# a_4808_45572# 0.001338f
C13072 a_19335_46494# a_19256_45572# 5.26e-20
C13073 a_6945_45028# a_18479_45785# 4.52e-21
C13074 a_17715_44484# a_17668_45572# 0.006757f
C13075 a_14976_45028# a_14976_45348# 0.002418f
C13076 a_1138_42852# a_413_45260# 0.026098f
C13077 a_18597_46090# a_20980_44850# 0.005953f
C13078 a_10586_45546# a_11682_45822# 0.014019f
C13079 a_14537_46482# a_13249_42308# 1.3e-20
C13080 a_4883_46098# a_19279_43940# 3.51e-21
C13081 a_18479_47436# a_3422_30871# 1.58e-20
C13082 a_9625_46129# a_3357_43084# 1.12e-20
C13083 a_167_45260# a_n467_45028# 1.04e-19
C13084 a_n2293_46098# a_4927_45028# 0.015237f
C13085 a_584_46384# a_n1435_47204# 5e-19
C13086 a_4915_47217# a_5815_47464# 0.064955f
C13087 a_4791_45118# a_6545_47178# 0.112353f
C13088 a_n1151_42308# a_9067_47204# 6.01e-21
C13089 a_n443_46116# a_6151_47436# 1.3e-19
C13090 a_n4064_40160# a_n4064_38528# 0.055466f
C13091 a_n3674_38216# VDD 0.309006f
C13092 a_n3565_39590# a_n4209_38502# 0.0315f
C13093 a_n4209_39304# a_n3690_39392# 0.045342f
C13094 a_n4334_39392# a_n3565_39304# 0.001004f
C13095 a_n4209_39590# a_n3565_38502# 0.031792f
C13096 a_1606_42308# C4_P_btm 3.05e-19
C13097 a_n784_42308# C4_N_btm 0.001073f
C13098 a_n1059_45260# a_17303_42282# 0.001091f
C13099 a_n2017_45002# a_17531_42308# 0.00607f
C13100 a_n913_45002# a_4958_30871# 0.058702f
C13101 a_11341_43940# a_2982_43646# 0.002145f
C13102 a_9159_44484# a_9127_43156# 7.52e-21
C13103 a_n2661_43922# a_8037_42858# 4.47e-22
C13104 a_n2293_43922# a_7765_42852# 1.03e-20
C13105 a_3422_30871# a_4190_30871# 12.909901f
C13106 a_n2293_42834# a_1576_42282# 5e-20
C13107 a_18579_44172# a_4361_42308# 6.73e-20
C13108 a_9313_44734# a_12379_42858# 0.05039f
C13109 a_20692_30879# C5_N_btm 3.17e-19
C13110 a_20205_31679# C6_N_btm 1.26e-20
C13111 a_12861_44030# a_14358_43442# 1.87e-20
C13112 a_10809_44734# a_10334_44484# 0.002242f
C13113 a_167_45260# a_n2661_43922# 2.12e-19
C13114 a_3483_46348# a_5708_44484# 0.005523f
C13115 a_18189_46348# a_17767_44458# 3.29e-19
C13116 a_17715_44484# a_17970_44736# 0.001614f
C13117 a_8199_44636# a_8375_44464# 0.043989f
C13118 a_8349_46414# a_5891_43370# 7.96e-21
C13119 a_15861_45028# a_17668_45572# 0.065471f
C13120 a_3090_45724# a_7281_43914# 0.170855f
C13121 a_17478_45572# a_17568_45572# 0.008441f
C13122 a_2711_45572# a_14537_43396# 0.249285f
C13123 a_1609_45822# a_1423_45028# 2.44e-19
C13124 a_5937_45572# a_7640_43914# 2.38e-19
C13125 a_8162_45546# a_5111_44636# 1.13e-21
C13126 a_n1613_43370# a_3877_44458# 1.43013f
C13127 a_8530_39574# VDD 0.346613f
C13128 a_4883_46098# a_9863_46634# 0.007473f
C13129 a_7754_38470# RST_Z 0.034995f
C13130 a_n2109_47186# a_765_45546# 0.126431f
C13131 VDAC_P C5_P_btm 7.72471f
C13132 a_12861_44030# a_11735_46660# 4.6e-21
C13133 a_n1435_47204# a_11901_46660# 7.78e-20
C13134 a_5063_47570# a_4955_46873# 3.3e-22
C13135 a_22609_37990# a_22717_36887# 0.08947f
C13136 a_22705_37990# a_22717_37285# 9.87e-19
C13137 a_n2472_46634# a_n2312_38680# 0.039578f
C13138 a_n2661_46634# a_n1925_46634# 4.75867f
C13139 a_n2442_46660# a_n2104_46634# 0.001169f
C13140 a_1115_44172# a_1576_42282# 2.71e-21
C13141 a_9313_44734# a_18727_42674# 2.59e-20
C13142 a_10341_43396# a_18429_43548# 0.012565f
C13143 a_n97_42460# a_7765_42852# 0.002083f
C13144 a_453_43940# a_564_42282# 4.63e-21
C13145 a_1414_42308# a_n1630_35242# 2.24e-20
C13146 a_413_45260# DATA[1] 0.004906f
C13147 a_3065_45002# VDD 0.501045f
C13148 a_15095_43370# a_15743_43084# 0.022008f
C13149 a_9145_43396# a_15231_43396# 0.005861f
C13150 a_1568_43370# a_791_42968# 4.67e-20
C13151 a_9396_43370# a_4361_42308# 3.82e-20
C13152 a_8685_43396# a_16823_43084# 7.39e-20
C13153 a_9290_44172# a_11173_43940# 0.001076f
C13154 a_7229_43940# a_n2293_42834# 0.148023f
C13155 a_8192_45572# a_8375_44464# 1.55e-21
C13156 a_11823_42460# a_n2293_43922# 0.494696f
C13157 a_6709_45028# a_7639_45394# 0.004982f
C13158 a_n2293_46098# a_4699_43561# 0.001614f
C13159 a_n863_45724# a_n984_44318# 0.002194f
C13160 a_5147_45002# a_n2661_43370# 0.034793f
C13161 a_n452_45724# a_n809_44244# 4.69e-20
C13162 a_n2293_46634# a_5342_30871# 3.03e-20
C13163 a_15227_44166# a_15781_43660# 0.016739f
C13164 a_626_44172# a_1145_45348# 0.009374f
C13165 a_17478_45572# a_17767_44458# 6.59e-21
C13166 a_n755_45592# a_n2065_43946# 3.71e-20
C13167 a_n357_42282# a_n1761_44111# 0.004602f
C13168 a_3232_43370# a_7418_45067# 0.001221f
C13169 a_6171_45002# a_10903_45394# 5.41e-20
C13170 a_8696_44636# a_18248_44752# 7.61e-21
C13171 a_n2661_45546# a_1414_42308# 3.34e-20
C13172 a_20447_31679# a_22959_45036# 4.88e-19
C13173 a_584_46384# a_1606_42308# 2.19e-19
C13174 a_3090_45724# a_16409_43396# 4.65e-21
C13175 a_16327_47482# a_16877_42852# 7.73e-21
C13176 a_n2017_45002# a_18184_42460# 0.205351f
C13177 a_18834_46812# a_19333_46634# 3.48e-20
C13178 a_19386_47436# a_8049_45260# 2.52e-22
C13179 a_n2661_46634# a_10355_46116# 6.98e-21
C13180 a_n1925_46634# a_8199_44636# 0.007627f
C13181 a_2443_46660# a_1823_45246# 0.001195f
C13182 a_1799_45572# a_167_45260# 0.061186f
C13183 a_3877_44458# a_n2293_46098# 0.030683f
C13184 a_n971_45724# a_3503_45724# 0.011412f
C13185 a_n237_47217# a_3218_45724# 1.35e-20
C13186 a_n2497_47436# a_1609_45822# 1.24e-19
C13187 a_584_46384# a_380_45546# 0.0075f
C13188 a_2107_46812# a_4419_46090# 0.007223f
C13189 a_n2661_46098# a_2202_46116# 0.002327f
C13190 a_n881_46662# a_n2956_38680# 5.42e-20
C13191 a_n1613_43370# a_n1736_46482# 2.61e-19
C13192 a_12549_44172# a_19335_46494# 3.43e-19
C13193 a_13747_46662# a_14493_46090# 5.42e-19
C13194 a_5807_45002# a_15015_46420# 1.7e-19
C13195 a_n743_46660# a_8016_46348# 0.155955f
C13196 a_9804_47204# a_6945_45028# 0.028722f
C13197 a_n97_42460# a_13657_42308# 0.005924f
C13198 a_2905_42968# a_2987_42968# 0.004999f
C13199 a_19319_43548# a_19511_42282# 1.71e-21
C13200 a_2982_43646# a_10723_42308# 2.53e-19
C13201 a_15463_44811# VDD 6.37e-19
C13202 a_4190_30871# a_18504_43218# 9.82e-19
C13203 a_15743_43084# a_14097_32519# 0.001681f
C13204 a_15279_43071# a_15567_42826# 7.4e-20
C13205 a_10903_43370# a_12545_42858# 0.026404f
C13206 a_n357_42282# a_14579_43548# 0.049501f
C13207 a_n443_42852# a_5565_43396# 1.34e-19
C13208 a_n2433_44484# a_n2012_44484# 0.093133f
C13209 a_n2661_44458# a_n1809_44850# 0.003338f
C13210 a_3537_45260# a_5244_44056# 6.11e-20
C13211 a_5147_45002# a_2998_44172# 7.85e-20
C13212 a_16375_45002# a_17499_43370# 1.41e-19
C13213 a_n1925_42282# a_n1991_42858# 1.72e-19
C13214 a_11823_42460# a_n97_42460# 0.324041f
C13215 a_22612_30879# a_22775_42308# 8.11e-21
C13216 a_4185_45028# a_21356_42826# 1.61e-20
C13217 a_9290_44172# a_13460_43230# 0.005304f
C13218 a_13259_45724# a_18525_43370# 5.74e-20
C13219 a_3232_43370# a_2479_44172# 0.003118f
C13220 a_15227_44166# a_21071_46482# 0.004602f
C13221 a_9863_47436# a_413_45260# 1.03e-19
C13222 a_n881_46662# a_16147_45260# 3.57e-19
C13223 a_13747_46662# a_15903_45785# 0.022255f
C13224 a_8953_45546# a_9569_46155# 0.014447f
C13225 a_13661_43548# a_15765_45572# 1.83e-20
C13226 a_2063_45854# a_8953_45002# 2.32e-19
C13227 a_n1151_42308# a_7276_45260# 0.062423f
C13228 a_13059_46348# a_12638_46436# 0.053952f
C13229 a_20894_47436# a_2437_43646# 0.007723f
C13230 a_18597_46090# a_3357_43084# 0.160577f
C13231 a_5257_43370# a_6472_45840# 0.012073f
C13232 a_8667_46634# a_2711_45572# 3.36e-20
C13233 a_n1853_46287# a_n2956_39304# 8.18e-20
C13234 a_19466_46812# a_19443_46116# 0.004595f
C13235 a_4791_45118# a_4927_45028# 0.03353f
C13236 a_n1925_46634# a_8192_45572# 0.03394f
C13237 a_8199_44636# a_10355_46116# 0.176325f
C13238 a_3147_46376# a_2324_44458# 2.35e-21
C13239 a_n2293_46098# a_n1736_46482# 0.002983f
C13240 a_n2157_46122# a_n2956_38680# 0.001648f
C13241 a_8016_46348# a_11189_46129# 1.23e-20
C13242 a_5807_45002# a_16333_45814# 3.87e-19
C13243 a_12549_44172# a_12749_45572# 0.004689f
C13244 a_12891_46348# a_13297_45572# 3.27e-19
C13245 a_458_43396# VDD 0.431902f
C13246 a_19987_42826# a_17303_42282# 5.3e-20
C13247 a_14097_32519# a_1606_42308# 2.3e-20
C13248 a_17333_42852# a_18214_42558# 0.00105f
C13249 a_18249_42858# a_19332_42282# 4.14e-19
C13250 a_18599_43230# a_18727_42674# 1e-19
C13251 a_18817_42826# a_18907_42674# 7.77e-19
C13252 COMP_P a_n961_42308# 0.001912f
C13253 a_n4318_38216# a_n3674_37592# 0.077253f
C13254 a_n3674_38680# a_n1630_35242# 0.020981f
C13255 a_n3674_38216# a_n784_42308# 0.001581f
C13256 a_5534_30871# a_7174_31319# 0.038837f
C13257 a_3080_42308# C4_N_btm 5.72e-19
C13258 a_18989_43940# a_15493_43396# 2.4e-19
C13259 a_n2293_43922# a_n1644_44306# 1.12e-19
C13260 a_5891_43370# a_7911_44260# 2.91e-19
C13261 a_19279_43940# a_21145_44484# 0.004519f
C13262 a_3357_43084# a_743_42282# 1.72e-19
C13263 a_n699_43396# a_726_44056# 7.74e-20
C13264 a_3067_47026# VDD 0.132018f
C13265 a_11827_44484# a_21205_44306# 4.85e-19
C13266 a_n2661_43922# a_n1453_44318# 0.001188f
C13267 a_n2661_42834# a_n1287_44306# 6.06e-19
C13268 a_8696_44636# a_8387_43230# 7.22e-21
C13269 a_526_44458# a_9885_42558# 9.36e-19
C13270 a_13017_45260# a_13667_43396# 1.23e-20
C13271 a_9482_43914# a_9145_43396# 5.35e-19
C13272 a_14539_43914# a_11341_43940# 0.077754f
C13273 a_n2810_45572# a_n2472_42282# 2.3e-20
C13274 a_n356_44636# a_17737_43940# 3.52e-21
C13275 a_20679_44626# a_22591_44484# 4.6e-21
C13276 a_13059_46348# a_n2017_45002# 3.52e-20
C13277 a_526_44458# a_3775_45552# 0.015665f
C13278 a_15015_46420# a_15143_45578# 0.011172f
C13279 a_10809_44734# a_9049_44484# 9.15e-21
C13280 a_14976_45028# a_6171_45002# 0.024858f
C13281 a_19123_46287# a_3357_43084# 1.6e-20
C13282 a_2324_44458# a_13249_42308# 0.072143f
C13283 a_11189_46129# a_11682_45822# 0.00283f
C13284 a_4646_46812# a_7735_45067# 2.05e-19
C13285 a_768_44030# a_4223_44672# 0.136643f
C13286 a_11415_45002# a_17034_45572# 2.62e-19
C13287 a_20411_46873# a_2437_43646# 7.51e-20
C13288 a_10903_43370# a_10210_45822# 0.001155f
C13289 a_6945_45028# a_10180_45724# 2.08e-20
C13290 a_11735_46660# a_11787_45002# 1.9e-19
C13291 a_8199_44636# a_10544_45572# 1.89e-19
C13292 a_5066_45546# a_4099_45572# 4.69e-20
C13293 a_10227_46804# a_5891_43370# 0.2393f
C13294 a_n4318_37592# a_n2946_37690# 3.13e-20
C13295 a_5742_30871# a_1736_39043# 4.53e-20
C13296 a_19647_42308# a_7174_31319# 0.006018f
C13297 a_13258_32519# a_20712_42282# 0.016015f
C13298 a_19511_42282# a_21335_42336# 0.011904f
C13299 a_n784_42308# a_8530_39574# 1.98e-19
C13300 a_10807_43548# a_11173_43940# 0.013678f
C13301 a_10949_43914# a_11257_43940# 0.001366f
C13302 a_1414_42308# a_1427_43646# 0.006859f
C13303 a_4223_44672# a_5755_42852# 5.06e-21
C13304 a_3065_45002# a_n784_42308# 1.67e-20
C13305 a_n1059_45260# a_2713_42308# 0.002489f
C13306 a_n2017_45002# a_2903_42308# 0.013263f
C13307 a_n913_45002# a_2725_42558# 0.005368f
C13308 a_3357_43084# a_5755_42308# 2.11e-20
C13309 a_21137_46414# VDD 0.219745f
C13310 a_19900_46494# START 3.05e-20
C13311 a_20708_46348# RST_Z 5.4e-22
C13312 a_15682_46116# CLK 2.6e-19
C13313 a_11827_44484# a_18083_42858# 3.77e-21
C13314 a_n2293_42834# a_4649_42852# 4.54e-19
C13315 a_2998_44172# a_4093_43548# 2.37e-19
C13316 a_18184_42460# a_19164_43230# 0.001269f
C13317 a_18494_42460# a_19339_43156# 4.88e-20
C13318 a_4743_44484# a_4520_42826# 6.49e-21
C13319 a_12549_44172# a_22959_43948# 2.47e-20
C13320 a_n2956_39304# a_n2661_43370# 1.05e-20
C13321 a_15682_46116# a_17023_45118# 5.09e-19
C13322 a_n1099_45572# a_n967_45348# 3.54e-20
C13323 a_n2661_45546# a_1667_45002# 0.003128f
C13324 a_n2293_46634# a_9672_43914# 4.81e-20
C13325 a_4883_46098# a_9801_43940# 0.001598f
C13326 a_16327_47482# a_14401_32519# 2.02e-20
C13327 a_13527_45546# a_8696_44636# 2.77e-21
C13328 a_1823_45246# a_949_44458# 0.005758f
C13329 a_12741_44636# a_15004_44636# 0.008679f
C13330 a_n2293_45546# a_n37_45144# 0.042299f
C13331 a_14976_45028# a_14673_44172# 8.68e-20
C13332 a_5807_45002# a_15493_43396# 0.002975f
C13333 a_13661_43548# a_19328_44172# 2.29e-19
C13334 a_11823_42460# a_16020_45572# 5.14e-20
C13335 a_n863_45724# a_n467_45028# 0.037721f
C13336 a_11962_45724# a_12561_45572# 1.59e-19
C13337 a_4791_45118# a_4699_43561# 1.93e-20
C13338 a_584_46384# a_3539_42460# 9.82e-19
C13339 a_4419_46090# a_n2661_44458# 6.4e-20
C13340 a_11415_45002# a_16979_44734# 3.74e-20
C13341 a_n4209_37414# a_n4064_37440# 0.265895f
C13342 a_n3565_37414# a_n3420_37440# 0.307576f
C13343 VDAC_Ni a_3726_37500# 1.5261f
C13344 a_11453_44696# a_13747_46662# 0.046437f
C13345 a_n4064_40160# VREF_GND 0.493568f
C13346 a_21496_47436# a_21588_30879# 6.1e-19
C13347 a_n971_45724# a_7927_46660# 0.035261f
C13348 a_n1741_47186# a_10428_46928# 3.82e-19
C13349 a_n237_47217# a_7577_46660# 0.032223f
C13350 a_4700_47436# a_4646_46812# 0.010115f
C13351 a_4791_45118# a_3877_44458# 0.024145f
C13352 a_n4251_39616# VDD 3.95e-19
C13353 a_12465_44636# a_20843_47204# 8.77e-22
C13354 a_n3565_38502# C6_P_btm 1.26e-20
C13355 a_n3565_38216# a_n1532_35090# 1e-19
C13356 a_n4209_38216# EN_VIN_BSTR_P 0.004167f
C13357 a_n1151_42308# a_5167_46660# 0.011285f
C13358 a_584_46384# a_3633_46660# 1.85e-22
C13359 a_2063_45854# a_5275_47026# 1.75e-19
C13360 a_4883_46098# a_20916_46384# 0.471396f
C13361 en_comp a_11206_38545# 0.002407f
C13362 a_n2293_43922# a_961_42354# 5.68e-20
C13363 a_2813_43396# a_3457_43396# 0.026697f
C13364 a_n97_42460# a_18429_43548# 0.003367f
C13365 a_2982_43646# a_10341_43396# 0.029008f
C13366 a_20193_45348# a_20712_42282# 0.010791f
C13367 a_7112_43396# a_8685_43396# 2.65e-19
C13368 a_3626_43646# a_14955_43396# 4.11e-21
C13369 a_n356_44636# a_8515_42308# 1.17e-19
C13370 a_n2293_46634# a_743_42282# 4.23e-20
C13371 a_17339_46660# a_18533_43940# 0.006189f
C13372 a_n863_45724# a_n2661_43922# 0.115404f
C13373 a_16680_45572# a_17023_45118# 0.002499f
C13374 a_8696_44636# a_16922_45042# 0.10244f
C13375 a_2437_43646# a_2232_45348# 0.001172f
C13376 a_21588_30879# a_13678_32519# 0.056847f
C13377 a_3537_45260# a_5111_44636# 1.36722f
C13378 a_4574_45260# a_5147_45002# 0.001891f
C13379 a_16327_47482# a_18817_42826# 0.215236f
C13380 a_9049_44484# a_5883_43914# 0.025986f
C13381 a_7499_43078# a_9838_44484# 2.03e-20
C13382 a_n443_42852# a_7640_43914# 4e-21
C13383 a_12465_44636# a_12379_42858# 4.6e-19
C13384 a_8199_44636# a_10949_43914# 4.16e-20
C13385 a_584_46384# a_526_44458# 0.458472f
C13386 a_2063_45854# a_2981_46116# 0.001617f
C13387 a_6545_47178# a_6945_45028# 0.09952f
C13388 a_n1925_46634# a_765_45546# 0.029508f
C13389 a_13717_47436# a_15682_46116# 9.15e-21
C13390 a_12861_44030# a_2324_44458# 0.95556f
C13391 a_20916_46384# a_21188_46660# 0.003748f
C13392 a_13661_43548# a_18280_46660# 4.34e-19
C13393 a_n881_46662# a_n1423_46090# 4.07e-19
C13394 a_n1613_43370# a_n1641_46494# 0.152421f
C13395 a_4883_46098# a_6165_46155# 0.006098f
C13396 a_11599_46634# a_14493_46090# 0.018622f
C13397 a_10227_46804# a_9290_44172# 0.918064f
C13398 a_7577_46660# a_8270_45546# 1.63e-19
C13399 a_7927_46660# a_8023_46660# 0.013793f
C13400 a_8145_46902# a_8189_46660# 3.69e-19
C13401 a_768_44030# a_12741_44636# 0.03898f
C13402 a_n743_46660# a_15312_46660# 1.45e-21
C13403 a_7411_46660# a_8601_46660# 2.56e-19
C13404 a_6755_46942# a_6969_46634# 0.085936f
C13405 a_5649_42852# a_12545_42858# 3.24e-20
C13406 a_n4318_39768# a_n4064_39616# 0.047349f
C13407 a_n3674_39768# a_n2946_39866# 4.03e-21
C13408 a_6298_44484# VDD 1.21616f
C13409 a_4361_42308# a_13635_43156# 2.7e-19
C13410 a_743_42282# a_5342_30871# 0.035916f
C13411 a_16823_43084# a_17333_42852# 5.93e-19
C13412 a_17678_43396# a_17701_42308# 1.14e-19
C13413 a_14021_43940# a_14456_42282# 3.19e-21
C13414 a_n1557_42282# a_n2472_42282# 3.44e-20
C13415 a_15743_43084# a_22959_42860# 0.001327f
C13416 a_3422_30871# a_n3420_37984# 0.031681f
C13417 a_458_43396# a_n784_42308# 1.67e-20
C13418 a_n97_42460# a_961_42354# 5.71e-22
C13419 a_n2293_46634# a_5755_42308# 2.62e-20
C13420 a_n755_45592# a_n2129_43609# 0.001714f
C13421 a_n357_42282# a_n2267_43396# 8.73e-20
C13422 a_n2661_43370# a_10157_44484# 7.91e-20
C13423 a_1307_43914# a_5891_43370# 0.084799f
C13424 a_6171_45002# a_15433_44458# 2.27e-20
C13425 a_20567_45036# a_18114_32519# 1.7e-20
C13426 a_6755_46942# a_16877_43172# 2.09e-19
C13427 SMPL_ON_P a_n4209_38216# 8.15e-19
C13428 a_8191_45002# a_n2661_43922# 8.71e-21
C13429 a_8953_45002# a_n2661_42834# 2.09e-19
C13430 a_2437_43646# a_3422_30871# 4.22e-21
C13431 a_11691_44458# a_16981_45144# 1.91e-19
C13432 a_1423_45028# a_5205_44734# 0.001252f
C13433 a_n863_45724# a_n447_43370# 7e-19
C13434 a_1138_42852# a_n13_43084# 3.75e-20
C13435 a_4883_46098# a_10210_45822# 6.13e-19
C13436 a_n2661_46098# a_n1079_45724# 3.76e-21
C13437 a_13059_46348# a_13759_46122# 0.249771f
C13438 a_19333_46634# a_10809_44734# 0.011589f
C13439 a_15227_44166# a_22959_46124# 1.38e-19
C13440 a_14180_46812# a_2324_44458# 4.9e-20
C13441 a_12861_44030# a_16855_45546# 4.91e-19
C13442 a_10227_46804# a_11064_45572# 6.09e-20
C13443 a_171_46873# a_n23_45546# 1.53e-20
C13444 a_2107_46812# a_1848_45724# 2.4e-19
C13445 a_1799_45572# a_n863_45724# 7.63e-20
C13446 a_2959_46660# a_n2661_45546# 6.8e-21
C13447 a_n2293_46098# a_n1641_46494# 0.006575f
C13448 a_n2157_46122# a_n1423_46090# 0.053479f
C13449 a_n1853_46287# a_n1991_46122# 0.737461f
C13450 a_n881_46662# a_9049_44484# 4.56e-21
C13451 a_19692_46634# a_6945_45028# 0.669658f
C13452 a_10249_46116# a_9823_46482# 1.82e-19
C13453 a_10428_46928# a_10586_45546# 4.33e-19
C13454 a_5807_45002# a_6472_45840# 0.016039f
C13455 a_n2293_46634# a_2277_45546# 0.001814f
C13456 a_11599_46634# a_15903_45785# 0.00101f
C13457 a_5649_42852# a_19332_42282# 1.31e-19
C13458 a_4361_42308# a_18310_42308# 9.35e-19
C13459 a_10555_44260# VDD 0.004772f
C13460 a_5534_30871# a_5932_42308# 0.025879f
C13461 a_4190_30871# a_7174_31319# 0.153555f
C13462 a_743_42282# a_20107_42308# 0.00961f
C13463 a_4185_45028# a_8685_42308# 6.95e-20
C13464 a_3065_45002# a_3080_42308# 0.171466f
C13465 a_5883_43914# a_3905_42865# 5.97e-20
C13466 a_3094_47570# DATA[1] 2.62e-21
C13467 a_3357_43084# a_2813_43396# 3.3e-19
C13468 a_n357_42282# a_21671_42860# 0.001708f
C13469 a_n2956_39304# COMP_P 8.08e-19
C13470 a_n2956_38680# a_n4318_37592# 0.02321f
C13471 a_16922_45042# a_20365_43914# 0.021687f
C13472 a_15433_44458# a_14673_44172# 0.027789f
C13473 a_5518_44484# a_5663_43940# 3.51e-19
C13474 a_9313_44734# a_20679_44626# 1.18e-20
C13475 a_5343_44458# a_6453_43914# 1.64e-20
C13476 a_n967_45348# a_n1243_43396# 1.73e-19
C13477 a_11691_44458# a_10729_43914# 0.001834f
C13478 a_18184_42460# a_18079_43940# 2.26e-21
C13479 a_3537_45260# a_4235_43370# 0.010714f
C13480 a_4223_44672# a_7845_44172# 0.004668f
C13481 a_3094_47243# VDD 6.34e-20
C13482 a_n2017_45002# a_6293_42852# 2.51e-19
C13483 a_n1059_45260# a_6031_43396# 5.04e-20
C13484 a_11827_44484# a_12429_44172# 6.51e-20
C13485 a_8696_44636# a_15743_43084# 3.96e-21
C13486 a_11453_44696# a_18911_45144# 4.04e-19
C13487 a_8034_45724# a_8379_46155# 0.001152f
C13488 a_n2293_46634# a_626_44172# 0.005771f
C13489 a_22223_46124# a_20205_31679# 0.160234f
C13490 a_6945_45028# a_20692_30879# 6.72e-20
C13491 a_1823_45246# a_1990_45572# 0.001177f
C13492 a_11415_45002# a_11823_42460# 0.349238f
C13493 a_17609_46634# a_16147_45260# 2.56e-21
C13494 a_8049_45260# a_9241_46436# 0.009374f
C13495 a_20708_46348# a_21167_46155# 6.64e-19
C13496 a_768_44030# a_n2293_42834# 0.036156f
C13497 a_5907_46634# a_413_45260# 1.96e-20
C13498 a_3877_44458# a_3429_45260# 0.02987f
C13499 a_13059_46348# a_15297_45822# 0.002837f
C13500 a_6755_46942# a_3357_43084# 6.8e-20
C13501 a_3090_45724# a_18691_45572# 3.57e-19
C13502 a_13507_46334# a_11827_44484# 0.384415f
C13503 a_4791_45118# a_10440_44484# 1.07e-20
C13504 a_3483_46348# a_6511_45714# 8.76e-21
C13505 a_5204_45822# a_2711_45572# 0.021829f
C13506 a_n743_46660# a_16019_45002# 0.002622f
C13507 a_13657_42558# a_14113_42308# 0.001685f
C13508 a_14456_42282# a_15764_42576# 4.16e-21
C13509 a_17364_32525# VCM 0.035838f
C13510 a_11323_42473# a_11633_42308# 7.95e-20
C13511 a_5742_30871# a_10149_42308# 3.62e-19
C13512 a_n967_43230# VDD 2.82e-20
C13513 a_11827_44484# a_21855_43396# 1e-20
C13514 a_n2293_42834# a_5755_42852# 0.007961f
C13515 a_11823_42460# a_10533_42308# 0.002582f
C13516 a_14539_43914# a_10341_43396# 0.041922f
C13517 a_n443_42852# a_7174_31319# 4.88e-21
C13518 a_n2840_46090# VDD 0.295278f
C13519 a_n2661_42834# a_3626_43646# 2.47e-20
C13520 a_n2293_43922# a_2982_43646# 0.094429f
C13521 a_20193_45348# a_20556_43646# 0.009643f
C13522 a_1115_44172# a_1241_43940# 0.143754f
C13523 a_5891_43370# a_9396_43370# 0.004592f
C13524 a_19279_43940# a_19741_43940# 6.62e-20
C13525 a_18579_44172# a_18533_43940# 0.011624f
C13526 a_20679_44626# a_20974_43370# 1.79e-20
C13527 a_2711_45572# a_18727_42674# 1.2e-21
C13528 a_10193_42453# a_13575_42558# 0.175489f
C13529 a_3537_45260# a_5837_43172# 0.001f
C13530 a_21076_30879# SINGLE_ENDED 1.21e-19
C13531 a_18184_42460# a_14209_32519# 0.006261f
C13532 a_16327_47482# a_15682_43940# 0.002941f
C13533 a_5164_46348# a_5105_45348# 6.6e-20
C13534 a_8568_45546# a_7499_43078# 0.070368f
C13535 a_8162_45546# a_9049_44484# 6.68e-20
C13536 a_n1991_46122# a_n2661_43370# 8.66e-21
C13537 a_10227_46804# a_10807_43548# 0.025916f
C13538 a_n971_45724# a_8487_44056# 2.58e-21
C13539 a_2711_45572# a_8697_45822# 0.003205f
C13540 a_5937_45572# a_1423_45028# 0.083936f
C13541 a_2804_46116# a_2809_45028# 6.45e-21
C13542 a_11415_45002# a_16321_45348# 0.001041f
C13543 a_13259_45724# a_17034_45572# 0.002067f
C13544 a_8049_45260# a_3357_43084# 0.08902f
C13545 a_768_44030# a_1115_44172# 0.003218f
C13546 a_n1925_42282# a_n967_45348# 0.004046f
C13547 a_12861_44030# a_19862_44208# 0.721035f
C13548 a_9290_44172# a_1307_43914# 0.122831f
C13549 a_2324_44458# a_11787_45002# 0.002598f
C13550 a_13925_46122# a_9482_43914# 1.87e-19
C13551 a_13759_46122# a_13556_45296# 1.81e-20
C13552 a_n4209_39304# a_n3420_37440# 0.033347f
C13553 a_13575_42558# VDD 0.182133f
C13554 a_n3565_39304# a_n3565_37414# 0.029571f
C13555 a_n3420_39072# a_n4209_37414# 0.030579f
C13556 a_n4064_37984# a_n2302_37984# 0.250408f
C13557 a_n3420_37984# a_n3607_38304# 8.36e-19
C13558 a_n3565_38216# a_n2860_37984# 0.001043f
C13559 a_n4209_39590# VDAC_P 0.001941f
C13560 a_16241_47178# a_12465_44636# 2.08e-19
C13561 a_10227_46804# a_20990_47178# 0.004463f
C13562 a_16588_47582# a_13507_46334# 3.49e-21
C13563 a_18780_47178# a_19386_47436# 3.06e-19
C13564 a_11599_46634# a_11453_44696# 0.075707f
C13565 a_16023_47582# a_4883_46098# 5.48e-21
C13566 a_6151_47436# a_n1613_43370# 0.548675f
C13567 a_18479_47436# a_19787_47423# 0.029306f
C13568 a_4915_47217# a_4842_47243# 1.81e-19
C13569 a_n1151_42308# a_12549_44172# 0.466584f
C13570 a_n2109_47186# a_n2956_39768# 4.34e-19
C13571 a_n2288_47178# a_n2661_46634# 1.83e-19
C13572 a_n2497_47436# a_n2472_46634# 0.009668f
C13573 a_n2833_47464# a_n2442_46660# 0.055535f
C13574 a_19862_44208# a_19700_43370# 3.23e-19
C13575 a_15493_43396# a_16867_43762# 0.02646f
C13576 a_2479_44172# a_2905_42968# 0.163227f
C13577 a_20159_44458# a_19987_42826# 4.85e-21
C13578 a_n699_43396# a_n1630_35242# 1.22e-20
C13579 a_n2956_37592# a_n3690_38528# 1.91e-20
C13580 a_895_43940# a_2075_43172# 1.77e-19
C13581 a_2675_43914# a_1847_42826# 2.13e-20
C13582 a_11967_42832# a_21356_42826# 4.18e-21
C13583 a_9313_44734# a_12800_43218# 0.001591f
C13584 a_375_42282# a_7174_31319# 1.7e-20
C13585 a_n2810_45028# a_n3420_38528# 3.16e-21
C13586 a_20365_43914# a_15743_43084# 1.24e-20
C13587 a_15493_43940# a_16759_43396# 8.32e-19
C13588 a_11341_43940# a_17324_43396# 1.91e-20
C13589 a_n97_42460# a_2982_43646# 0.180648f
C13590 w_11334_34010# a_5342_30871# 0.00275f
C13591 a_6755_46942# a_18533_44260# 9.89e-21
C13592 a_n2293_45546# a_949_44458# 0.004678f
C13593 a_n2661_45546# a_n699_43396# 0.022358f
C13594 a_n2293_46634# a_2813_43396# 8.36e-19
C13595 a_19479_31679# a_3357_43084# 0.058337f
C13596 a_n863_45724# a_n452_44636# 0.01836f
C13597 a_8696_44636# a_10775_45002# 0.00249f
C13598 a_7499_43078# a_n2661_43370# 0.027764f
C13599 a_18597_46090# a_743_42282# 3.54e-19
C13600 a_n2293_46098# a_5244_44056# 6.1e-19
C13601 a_22223_45572# a_22591_45572# 7.52e-19
C13602 a_2437_43646# a_19963_31679# 5.48e-19
C13603 a_13259_45724# a_16979_44734# 3.78e-21
C13604 a_n755_45592# a_n2129_44697# 9.75e-19
C13605 a_1848_45724# a_n2661_44458# 3.76e-22
C13606 a_8270_45546# a_7499_43940# 5.55e-20
C13607 a_18479_47436# a_20107_46660# 0.019527f
C13608 a_n2661_46634# a_6999_46987# 2.56e-19
C13609 a_5807_45002# a_8846_46660# 6.99e-19
C13610 a_12549_44172# a_14084_46812# 0.007343f
C13611 a_768_44030# a_13607_46688# 2.12e-20
C13612 a_6151_47436# a_n2293_46098# 9.86e-20
C13613 C9_P_btm VREF 7.369471f
C13614 a_10227_46804# a_20273_46660# 0.037464f
C13615 a_15811_47375# a_16434_46660# 2.88e-19
C13616 a_2107_46812# a_7411_46660# 7.26e-20
C13617 a_n971_45724# a_5164_46348# 1.88e-20
C13618 a_n2293_46634# a_6755_46942# 1.78e-19
C13619 a_12465_44636# a_16721_46634# 9.65e-22
C13620 C5_N_btm C10_N_btm 0.285351f
C13621 C6_N_btm C9_N_btm 0.169882f
C13622 C7_N_btm C8_N_btm 23.7884f
C13623 a_18597_46090# a_19123_46287# 0.188676f
C13624 C3_N_btm VDD 0.26836f
C13625 C10_P_btm VREF_GND 10.3207f
C13626 C7_P_btm VIN_P 1.52449f
C13627 a_584_46384# a_2521_46116# 4.33e-19
C13628 a_2063_45854# a_167_45260# 0.359284f
C13629 a_n237_47217# a_4704_46090# 0.042359f
C13630 a_n743_46660# a_10428_46928# 4.37e-20
C13631 a_3699_46634# a_4817_46660# 1.58e-19
C13632 a_3524_46660# a_4955_46873# 7.68e-19
C13633 a_8685_43396# a_12545_42858# 5.31e-20
C13634 a_3626_43646# a_n2293_42282# 3.32e-19
C13635 a_n2661_42282# a_6123_31319# 0.017717f
C13636 a_4190_30871# a_21487_43396# 0.001675f
C13637 a_18114_32519# a_22521_39511# 1.28e-20
C13638 a_7418_45067# VDD 0.001744f
C13639 a_20301_43646# a_20556_43646# 0.114664f
C13640 a_3422_30871# a_19511_42282# 0.025144f
C13641 a_4093_43548# a_4743_43172# 8.1e-19
C13642 a_n97_42460# a_5837_42852# 0.011979f
C13643 a_10586_45546# a_10651_43940# 6.43e-22
C13644 a_n1925_42282# a_n1917_43396# 2.35e-19
C13645 a_17715_44484# a_3626_43646# 3.08e-21
C13646 a_n443_42852# a_10729_43914# 1.44e-20
C13647 a_n2661_45010# a_n23_44458# 0.049334f
C13648 a_n357_42282# a_19478_44306# 2.51e-20
C13649 a_3232_43370# a_5518_44484# 0.01014f
C13650 a_6171_45002# a_5343_44458# 2.23e-19
C13651 a_5147_45002# a_5883_43914# 0.008506f
C13652 a_9290_44172# a_9396_43370# 5.85e-20
C13653 a_12741_44636# a_16759_43396# 1.39e-19
C13654 a_3090_45724# a_3935_42891# 5.91e-20
C13655 a_15765_45572# a_11967_42832# 8.39e-21
C13656 a_3483_46348# a_13667_43396# 1.35e-19
C13657 a_13747_46662# a_14180_46482# 0.008333f
C13658 a_n1151_42308# a_11525_45546# 2.76e-20
C13659 a_6755_46942# a_9625_46129# 3.29e-19
C13660 a_6151_47436# a_7230_45938# 1.1e-20
C13661 a_6545_47178# a_6812_45938# 1.37e-19
C13662 a_10768_47026# a_3483_46348# 4.61e-20
C13663 a_3877_44458# a_6945_45028# 0.001558f
C13664 a_n2661_46098# a_1337_46436# 4.38e-19
C13665 a_2107_46812# a_4365_46436# 1.79e-19
C13666 a_10467_46802# a_9290_44172# 2.22e-19
C13667 a_10428_46928# a_11189_46129# 6.48e-21
C13668 a_n2293_46634# a_8049_45260# 1.91e-20
C13669 a_743_42282# a_5755_42308# 0.00936f
C13670 a_4361_42308# a_3905_42558# 0.001685f
C13671 a_15567_42826# a_15785_43172# 0.007234f
C13672 a_4190_30871# a_5932_42308# 0.018227f
C13673 a_n4318_38680# a_n1630_35242# 7.78e-20
C13674 a_19237_31679# VCM 0.03748f
C13675 a_5649_42852# a_5379_42460# 0.35554f
C13676 a_2479_44172# VDD 0.431428f
C13677 a_2063_45854# DATA[4] 3.07e-19
C13678 a_10334_44484# a_11541_44484# 4.15e-20
C13679 a_4007_47204# VDD 0.41212f
C13680 a_1423_45028# a_8333_44056# 1.17e-19
C13681 a_n1151_42308# CLK_DATA 1.24e-21
C13682 a_2952_47436# DATA[2] 2.12e-19
C13683 a_n863_45724# a_n1641_43230# 2.33e-21
C13684 a_9290_44172# a_13003_42852# 7.01e-20
C13685 a_2905_45572# DATA[1] 1.91e-21
C13686 a_11827_44484# a_20637_44484# 9.54e-20
C13687 a_10903_43370# a_13157_43218# 6.01e-19
C13688 a_18114_32519# a_20679_44626# 6.99e-19
C13689 a_1307_43914# a_10807_43548# 0.016974f
C13690 a_n2293_42834# a_7845_44172# 0.008819f
C13691 a_14537_43396# a_15682_43940# 0.01288f
C13692 a_14797_45144# a_14955_43940# 4.38e-20
C13693 a_13720_44458# a_13857_44734# 0.126609f
C13694 SMPL_ON_N a_22521_40055# 5.57e-20
C13695 a_8016_46348# a_8379_46155# 0.005265f
C13696 a_12251_46660# a_11823_42460# 2.92e-20
C13697 a_3090_45724# a_10490_45724# 1.78e-21
C13698 a_9625_46129# a_8049_45260# 0.04571f
C13699 a_8953_45546# a_9241_46436# 2.17e-19
C13700 a_n881_46662# a_5147_45002# 3.9e-19
C13701 a_n1613_43370# a_5111_44636# 0.601769f
C13702 a_13507_46334# a_15595_45028# 1.41e-20
C13703 a_12465_44636# a_14180_45002# 0.015526f
C13704 a_11453_44696# a_13348_45260# 0.005514f
C13705 a_13661_43548# a_n913_45002# 6.88e-20
C13706 a_768_44030# a_413_45260# 0.182253f
C13707 a_5267_42460# a_5934_30871# 1.28e-20
C13708 a_5342_30871# a_n4064_37984# 0.028465f
C13709 a_n784_42308# a_13575_42558# 2.06e-20
C13710 a_14635_42282# a_7174_31319# 4.88e-21
C13711 a_1067_42314# a_5742_30871# 1.17e-20
C13712 a_n443_42852# a_5932_42308# 4.07e-19
C13713 a_n2956_39304# a_n4209_39304# 0.328727f
C13714 a_15368_46634# VDD 0.324877f
C13715 a_n1549_44318# a_n1287_44306# 0.001705f
C13716 a_n1331_43914# a_n875_44318# 4.2e-19
C13717 a_n1761_44111# a_n1441_43940# 8.49e-19
C13718 a_11967_42832# a_19328_44172# 1.02e-19
C13719 a_626_44172# a_743_42282# 6.2e-19
C13720 a_n1059_45260# a_10796_42968# 0.01348f
C13721 a_n913_45002# a_10835_43094# 0.053818f
C13722 a_n2017_45002# a_10991_42826# 1.61e-19
C13723 a_13259_45724# a_13657_42308# 6.47e-20
C13724 a_14539_43914# a_n97_42460# 0.05616f
C13725 a_5518_44484# a_4905_42826# 7.14e-20
C13726 a_742_44458# a_2982_43646# 9.65e-20
C13727 a_2998_44172# a_3600_43914# 0.012242f
C13728 a_14976_45028# RST_Z 2.6e-20
C13729 a_2382_45260# a_3681_42891# 0.067836f
C13730 a_11735_46660# CLK 6.72e-20
C13731 a_n357_42282# a_9223_42460# 3.69e-20
C13732 a_n755_45592# a_8791_42308# 7.02e-19
C13733 a_n699_43396# a_1427_43646# 0.00477f
C13734 a_n2661_42834# a_3052_44056# 1.84e-19
C13735 a_17517_44484# a_15493_43940# 7.18e-20
C13736 a_3316_45546# a_3175_45822# 0.05019f
C13737 a_3503_45724# a_2711_45572# 0.058013f
C13738 a_13259_45724# a_11823_42460# 0.626941f
C13739 a_8049_45260# a_9159_45572# 1.83e-19
C13740 a_768_44030# a_13468_44734# 0.001477f
C13741 SMPL_ON_P a_n2661_42282# 0.003852f
C13742 a_n1151_42308# a_7542_44172# 2.32e-19
C13743 a_4646_46812# a_6298_44484# 1.65052f
C13744 a_526_44458# a_8696_44636# 5.2e-21
C13745 a_19553_46090# a_19256_45572# 1.97e-19
C13746 a_19335_46494# a_19431_45546# 0.002697f
C13747 a_18819_46122# a_18799_45938# 2.22e-19
C13748 a_6945_45028# a_18175_45572# 3.9e-21
C13749 a_17583_46090# a_17668_45572# 5.29e-21
C13750 a_17715_44484# a_17568_45572# 0.001302f
C13751 a_1176_45822# a_413_45260# 3.98e-20
C13752 a_4791_45118# a_5244_44056# 0.003487f
C13753 a_16327_47482# a_20512_43084# 0.118893f
C13754 a_8953_45546# a_3357_43084# 2.47e-20
C13755 a_4185_45028# a_n913_45002# 0.855072f
C13756 a_9823_46155# a_2437_43646# 1.23e-20
C13757 a_n2293_46098# a_5111_44636# 0.086926f
C13758 a_10586_45546# a_11280_45822# 1.28e-20
C13759 a_n1151_42308# a_6575_47204# 1.72e-19
C13760 a_2124_47436# a_n1435_47204# 2.1e-19
C13761 a_4915_47217# a_5129_47502# 0.070911f
C13762 a_4791_45118# a_6151_47436# 0.019937f
C13763 a_2063_45854# a_11459_47204# 8.65e-20
C13764 a_n443_46116# a_5815_47464# 5.77e-19
C13765 a_n4064_40160# a_n2946_38778# 1.87e-20
C13766 a_7174_31319# a_n3420_37984# 7.78e-20
C13767 a_n4315_30879# a_n2302_38778# 6.48e-20
C13768 a_5742_30871# a_3726_37500# 0.001929f
C13769 a_n2104_42282# VDD 0.280329f
C13770 a_1606_42308# C5_P_btm 1.89e-19
C13771 a_n784_42308# C3_N_btm 0.001962f
C13772 a_n3607_39616# a_n3420_39072# 3.77e-20
C13773 a_n4209_39304# a_n3565_39304# 6.82668f
C13774 a_9313_44734# a_10341_42308# 0.019286f
C13775 a_n1059_45260# a_4958_30871# 0.005345f
C13776 a_n2017_45002# a_17303_42282# 0.006515f
C13777 a_5343_44458# a_8292_43218# 0.01105f
C13778 a_21115_43940# a_2982_43646# 5.25e-20
C13779 a_10807_43548# a_9396_43370# 2.23e-20
C13780 a_n2661_43922# a_7765_42852# 2.66e-21
C13781 a_n2293_43922# a_7871_42858# 1.21e-20
C13782 a_n2661_42834# a_8037_42858# 7.33e-22
C13783 a_3422_30871# a_21259_43561# 1.69e-19
C13784 a_21398_44850# a_4190_30871# 8.73e-21
C13785 a_20692_30879# C4_N_btm 5.85e-20
C13786 a_20205_31679# C5_N_btm 0.00105f
C13787 en_comp a_17124_42282# 4.59e-20
C13788 a_12861_44030# a_14579_43548# 1.6e-20
C13789 a_10809_44734# a_10157_44484# 3.6e-19
C13790 a_3699_46348# a_3363_44484# 1.94e-21
C13791 a_3483_46348# a_5608_44484# 0.001851f
C13792 a_9049_44484# a_3537_45260# 1.31e-19
C13793 a_17715_44484# a_17767_44458# 0.07408f
C13794 a_8016_46348# a_5891_43370# 0.183035f
C13795 a_1823_45246# a_n2293_43922# 1.33e-19
C13796 a_12741_44636# a_17517_44484# 0.01998f
C13797 a_3090_45724# a_6453_43914# 0.00316f
C13798 a_15861_45028# a_17568_45572# 0.004094f
C13799 a_8696_44636# a_17668_45572# 2.03e-19
C13800 a_n2293_46634# a_15037_43940# 0.001262f
C13801 a_2711_45572# a_14180_45002# 0.147337f
C13802 a_n443_42852# a_1423_45028# 1.15e-19
C13803 a_5937_45572# a_6109_44484# 0.163331f
C13804 a_8199_44636# a_7640_43914# 0.003096f
C13805 a_n2442_46660# a_n2293_46634# 0.004958f
C13806 a_n2472_46634# a_n2104_46634# 7.52e-19
C13807 a_4915_47217# a_15227_44166# 1.46e-20
C13808 a_n1613_43370# a_3221_46660# 0.003155f
C13809 a_7754_38470# VDD 0.302129f
C13810 a_4883_46098# a_8492_46660# 4.2e-20
C13811 VDAC_P C6_P_btm 15.441001f
C13812 a_n1435_47204# a_11813_46116# 2.37e-20
C13813 a_n2661_46634# a_n2312_38680# 0.106815f
C13814 a_n2956_39768# a_n1925_46634# 1.65e-19
C13815 a_768_44030# a_2609_46660# 1.29e-19
C13816 a_8791_43396# a_4361_42308# 2.28e-21
C13817 a_9313_44734# a_18057_42282# 2.51e-20
C13818 a_10341_43396# a_17324_43396# 0.010417f
C13819 a_n97_42460# a_7871_42858# 0.001218f
C13820 a_1115_44172# a_1067_42314# 2.43e-21
C13821 a_2680_45002# VDD 0.145087f
C13822 a_9145_43396# a_15125_43396# 0.001605f
C13823 a_1049_43396# a_791_42968# 5.89e-19
C13824 a_1568_43370# a_685_42968# 1.82e-20
C13825 a_15681_43442# a_15781_43660# 0.167615f
C13826 a_7287_43370# a_5649_42852# 1.08e-21
C13827 a_15037_43940# a_5342_30871# 6.83e-20
C13828 a_1414_42308# a_564_42282# 1.31e-20
C13829 a_9290_44172# a_10867_43940# 2.47e-19
C13830 a_1823_45246# a_n97_42460# 0.006778f
C13831 a_11823_42460# a_n2661_43922# 0.005005f
C13832 a_7276_45260# a_n2293_42834# 1.85e-19
C13833 a_n863_45724# a_n809_44244# 0.016179f
C13834 a_4558_45348# a_n2661_43370# 0.018142f
C13835 a_21188_45572# a_19721_31679# 3.94e-20
C13836 a_n1151_42308# a_n1630_35242# 0.056434f
C13837 a_15227_44166# a_15681_43442# 0.015868f
C13838 a_6171_45002# a_8560_45348# 0.004926f
C13839 a_7499_43078# a_11909_44484# 7.77e-22
C13840 a_8696_44636# a_17970_44736# 4.11e-19
C13841 a_12465_44636# a_12800_43218# 4.53e-20
C13842 a_3357_43084# a_20193_45348# 1.08e-20
C13843 a_3090_45724# a_16547_43609# 3.84e-21
C13844 a_22959_45572# a_22959_45036# 0.026152f
C13845 a_17478_45572# a_16979_44734# 9.61e-20
C13846 w_1575_34946# a_4958_30871# 0.00296f
C13847 a_8128_46384# a_6945_45028# 0.010979f
C13848 a_18834_46812# a_15227_44166# 0.231715f
C13849 a_18597_46090# a_8049_45260# 0.047215f
C13850 a_n2661_46634# a_9823_46155# 1.75e-20
C13851 a_n1925_46634# a_8349_46414# 0.006458f
C13852 a_n1151_42308# a_n2661_45546# 0.044338f
C13853 a_12861_44030# a_12839_46116# 0.003823f
C13854 a_11735_46660# a_14035_46660# 4.06e-21
C13855 a_12816_46660# a_12978_47026# 0.006453f
C13856 a_12251_46660# a_12513_46660# 0.001705f
C13857 a_12469_46902# a_12925_46660# 4.2e-19
C13858 a_11599_46634# a_14180_46482# 0.016275f
C13859 a_n971_45724# a_3316_45546# 0.086835f
C13860 a_n237_47217# a_2957_45546# 5.41e-20
C13861 a_n2497_47436# a_n443_42852# 0.005218f
C13862 a_2107_46812# a_4185_45028# 0.008044f
C13863 a_n2661_46098# a_1823_45246# 9.15e-19
C13864 a_1799_45572# a_2202_46116# 6.85e-20
C13865 a_n2293_46634# a_8953_45546# 0.04453f
C13866 a_6999_46987# a_765_45546# 2.41e-19
C13867 a_13747_46662# a_13925_46122# 0.020304f
C13868 a_5807_45002# a_14275_46494# 0.013842f
C13869 a_12549_44172# a_19553_46090# 7.25e-21
C13870 a_n743_46660# a_7920_46348# 0.006742f
C13871 a_2063_45854# a_n863_45724# 4.66e-19
C13872 a_n97_42460# a_11897_42308# 7.16e-19
C13873 a_7112_43396# a_6123_31319# 1.32e-19
C13874 a_17730_32519# a_22459_39145# 1.35e-20
C13875 a_2982_43646# a_10533_42308# 1.49e-19
C13876 a_15146_44811# VDD 6.34e-20
C13877 a_10617_44484# CLK 6.69e-19
C13878 a_15743_43084# a_22400_42852# 0.010325f
C13879 a_15279_43071# a_5342_30871# 0.214197f
C13880 a_10903_43370# a_12089_42308# 3.79e-19
C13881 a_n443_42852# a_4181_43396# 1.39e-19
C13882 a_n2661_44458# a_n2012_44484# 0.003432f
C13883 a_n4318_40392# a_n1809_44850# 5.8e-21
C13884 a_18494_42460# a_9313_44734# 0.028817f
C13885 a_3537_45260# a_3905_42865# 0.258917f
C13886 a_4558_45348# a_2998_44172# 2.03e-19
C13887 a_n1925_42282# a_n1853_43023# 0.003483f
C13888 a_4185_45028# a_20922_43172# 9.67e-21
C13889 a_21588_30879# a_22775_42308# 7.29e-21
C13890 a_9290_44172# a_13635_43156# 0.394766f
C13891 a_n967_45348# a_n875_44318# 4.26e-20
C13892 w_1575_34946# VCM 0.001153f
C13893 a_19123_46287# a_8049_45260# 3.32e-19
C13894 a_12549_44172# a_12649_45572# 0.004247f
C13895 a_15227_44166# a_20850_46482# 9.67e-19
C13896 a_9067_47204# a_413_45260# 4.35e-19
C13897 a_n881_46662# a_17786_45822# 4.61e-20
C13898 a_3877_44458# a_6812_45938# 4.82e-21
C13899 a_13661_43548# a_15903_45785# 0.001692f
C13900 a_13747_46662# a_15599_45572# 0.041358f
C13901 a_5807_45002# a_15765_45572# 0.003059f
C13902 a_8953_45546# a_9625_46129# 0.009628f
C13903 a_n1151_42308# a_5205_44484# 1.12e-20
C13904 a_13059_46348# a_12379_46436# 9.42e-19
C13905 a_13507_46334# a_21350_45938# 2.55e-20
C13906 a_19787_47423# a_2437_43646# 0.006262f
C13907 a_18597_46090# a_19479_31679# 3e-20
C13908 a_5257_43370# a_6194_45824# 0.029055f
C13909 a_4955_46873# a_4880_45572# 1.35e-20
C13910 a_4791_45118# a_5111_44636# 1.11355f
C13911 a_n2497_47436# a_375_42282# 0.018989f
C13912 a_n1925_46634# a_8120_45572# 0.004093f
C13913 a_8199_44636# a_9823_46155# 0.001773f
C13914 a_2804_46116# a_2324_44458# 1.12e-21
C13915 a_n2157_46122# a_n2956_39304# 7.88e-20
C13916 a_n2293_46098# a_n2956_38680# 0.022177f
C13917 a_8016_46348# a_9290_44172# 0.020766f
C13918 a_18780_47178# a_3357_43084# 2.77e-19
C13919 a_n229_43646# VDD 0.278436f
C13920 a_19164_43230# a_17303_42282# 9.77e-21
C13921 COMP_P a_n1329_42308# 0.232443f
C13922 a_n2472_42282# a_n3674_37592# 0.007439f
C13923 a_n2104_42282# a_n784_42308# 8.09e-20
C13924 a_18083_42858# a_18214_42558# 0.001378f
C13925 a_18249_42858# a_18907_42674# 0.001692f
C13926 a_18817_42826# a_18727_42674# 0.001214f
C13927 a_n2840_42282# a_n1630_35242# 0.040623f
C13928 a_5342_30871# a_13258_32519# 0.030303f
C13929 a_3080_42308# C3_N_btm 0.027071f
C13930 a_949_44458# a_1443_43940# 2.54e-19
C13931 a_18374_44850# a_15493_43396# 3.95e-21
C13932 a_n2293_43922# a_n3674_39768# 0.018871f
C13933 a_18989_43940# a_19328_44172# 4.08e-19
C13934 a_5891_43370# a_7584_44260# 2.54e-20
C13935 a_n2661_43922# a_n1644_44306# 0.002488f
C13936 a_20835_44721# a_20512_43084# 1.67e-21
C13937 a_20679_44626# a_22485_44484# 8.1e-21
C13938 a_20766_44850# a_21145_44484# 3.16e-19
C13939 a_19279_43940# a_21073_44484# 0.002178f
C13940 a_10057_43914# a_10555_44260# 0.041594f
C13941 a_2864_46660# VDD 0.076834f
C13942 a_n2661_42834# a_n1453_44318# 0.001232f
C13943 a_7640_43914# a_8018_44260# 9.16e-20
C13944 a_8696_44636# a_8605_42826# 4.39e-21
C13945 a_n357_42282# a_20256_43172# 3.27e-19
C13946 a_13348_45260# a_9145_43396# 9.73e-20
C13947 a_n2810_45572# a_n3674_38680# 0.023027f
C13948 a_8199_44636# a_7174_31319# 4.88e-21
C13949 a_20640_44752# a_22591_44484# 8.79e-21
C13950 a_n356_44636# a_15682_43940# 3.38e-21
C13951 a_8128_46384# a_8103_44636# 8.65e-21
C13952 a_10809_44734# a_7499_43078# 0.053075f
C13953 a_768_44030# a_2779_44458# 0.014949f
C13954 a_3090_45724# a_6171_45002# 0.030689f
C13955 a_9313_45822# a_n2661_43922# 3.03e-20
C13956 a_18285_46348# a_3357_43084# 1.63e-20
C13957 a_2324_44458# a_13904_45546# 0.004897f
C13958 a_11133_46155# a_10907_45822# 8.41e-19
C13959 a_11189_46129# a_11280_45822# 0.001906f
C13960 a_4646_46812# a_7418_45067# 0.001853f
C13961 a_9290_44172# a_11682_45822# 0.00219f
C13962 a_11415_45002# a_16789_45572# 1.55e-19
C13963 a_20107_46660# a_2437_43646# 5.01e-21
C13964 a_6945_45028# a_10053_45546# 5.1e-22
C13965 a_n743_46660# a_11827_44484# 2.74e-20
C13966 a_8270_45546# a_9482_43914# 0.004867f
C13967 a_8953_45546# a_9159_45572# 0.004909f
C13968 a_8199_44636# a_10306_45572# 5.75e-19
C13969 a_14097_32519# VDAC_N 2.69e-19
C13970 a_n1630_35242# VDAC_Ni 2.54e-19
C13971 a_13258_32519# a_20107_42308# 0.021019f
C13972 a_17303_42282# a_21973_42336# 5.22e-19
C13973 a_n4318_37592# a_n3420_37440# 0.001831f
C13974 a_5742_30871# a_1239_39043# 5.42e-20
C13975 a_5932_42308# a_n3420_37984# 1.17e-19
C13976 a_1793_42852# VDD 6.57e-19
C13977 a_19511_42282# a_7174_31319# 0.240861f
C13978 a_n784_42308# a_7754_38470# 1.35e-19
C13979 a_n1441_43940# a_n2267_43396# 4.29e-19
C13980 a_10729_43914# a_11257_43940# 0.007166f
C13981 a_10949_43914# a_11173_43940# 4.93e-19
C13982 a_10807_43548# a_10867_43940# 9.12e-19
C13983 a_1467_44172# a_1427_43646# 0.104539f
C13984 a_1414_42308# a_n1557_42282# 2.99e-21
C13985 a_n699_43396# a_4520_42826# 8.42e-22
C13986 a_4223_44672# a_5111_42852# 3.04e-21
C13987 a_n1059_45260# a_2725_42558# 2.97e-19
C13988 a_n2017_45002# a_2713_42308# 0.011694f
C13989 a_20708_46348# VDD 0.093079f
C13990 a_2324_44458# CLK 0.035116f
C13991 a_n2661_44458# a_10835_43094# 8.47e-20
C13992 a_11691_44458# a_15567_42826# 4.44e-21
C13993 a_11827_44484# a_17701_42308# 5.54e-22
C13994 en_comp a_1755_42282# 9.98e-21
C13995 a_18184_42460# a_19339_43156# 0.004558f
C13996 a_9313_44734# a_15940_43402# 4.1e-19
C13997 a_2479_44172# a_3080_42308# 0.001674f
C13998 a_12549_44172# a_15493_43940# 0.932577f
C13999 a_15682_46116# a_16922_45042# 6.61e-19
C14000 a_n755_45592# a_n745_45366# 0.014023f
C14001 a_n2661_45546# a_327_44734# 7.19e-19
C14002 a_4883_46098# a_9420_43940# 0.001234f
C14003 a_16327_47482# a_21381_43940# 0.001197f
C14004 a_5066_45546# a_5105_45348# 1.87e-19
C14005 a_11280_45822# a_11136_45572# 6.84e-19
C14006 a_15143_45578# a_15765_45572# 1.5e-19
C14007 a_1823_45246# a_742_44458# 4.02e-19
C14008 a_12741_44636# a_13720_44458# 0.00841f
C14009 a_n356_45724# a_n2661_45010# 6.56e-21
C14010 a_n2293_45546# a_n143_45144# 0.012062f
C14011 a_n2438_43548# a_n2661_42282# 4.44e-20
C14012 a_3090_45724# a_14673_44172# 0.018197f
C14013 a_2307_45899# a_2437_43646# 4.14e-19
C14014 a_13661_43548# a_18451_43940# 0.129334f
C14015 a_5807_45002# a_19328_44172# 7.07e-21
C14016 a_584_46384# a_3626_43646# 0.195961f
C14017 a_4185_45028# a_n2661_44458# 0.030414f
C14018 a_1138_42852# a_949_44458# 0.013552f
C14019 a_11415_45002# a_14539_43914# 0.010769f
C14020 a_n3565_37414# a_n3690_37440# 0.247968f
C14021 a_n4334_37440# a_n3420_37440# 0.015567f
C14022 a_n4209_37414# a_n2946_37690# 0.023544f
C14023 a_1736_39587# VDD 3.14139f
C14024 a_n4209_38502# C5_P_btm 0.040445f
C14025 a_n3565_38502# C7_P_btm 1.43e-20
C14026 a_n4315_30879# VCM 0.473529f
C14027 a_n3565_38216# a_n1386_35608# 1.22e-21
C14028 a_n4064_40160# VREF 1.12e-19
C14029 a_11453_44696# a_13661_43548# 0.099457f
C14030 a_21496_47436# a_20916_46384# 0.113102f
C14031 a_13507_46334# a_21588_30879# 6.05e-19
C14032 a_n971_45724# a_8145_46902# 0.051701f
C14033 a_n1741_47186# a_10150_46912# 2.54e-20
C14034 a_n237_47217# a_7715_46873# 0.051915f
C14035 a_4700_47436# a_3877_44458# 4.34e-21
C14036 a_n443_46116# a_3055_46660# 0.002062f
C14037 a_12465_44636# a_19594_46812# 9.01e-20
C14038 a_16588_47582# a_n743_46660# 1.72e-19
C14039 a_n1151_42308# a_5385_46902# 0.0125f
C14040 en_comp VDAC_P 0.003461f
C14041 a_19963_31679# a_22609_38406# 3.67e-21
C14042 a_n2293_43922# a_1184_42692# 3.75e-20
C14043 a_n97_42460# a_17324_43396# 0.003115f
C14044 a_7287_43370# a_8685_43396# 7.31e-19
C14045 a_13483_43940# a_12545_42858# 6.25e-20
C14046 a_n356_44636# a_5934_30871# 0.095373f
C14047 a_3626_43646# a_15095_43370# 1.07e-19
C14048 a_3065_45002# a_4927_45028# 1.12e-20
C14049 a_3429_45260# a_5111_44636# 3.89e-22
C14050 a_8953_45546# a_9672_43914# 1.03e-19
C14051 a_8199_44636# a_10729_43914# 3.27e-20
C14052 a_8016_46348# a_10807_43548# 1.5e-19
C14053 a_12861_44030# a_21671_42860# 5.22e-22
C14054 a_17339_46660# a_19319_43548# 2.03e-19
C14055 a_n863_45724# a_n2661_42834# 0.094705f
C14056 a_16375_45002# a_17517_44484# 4.98e-19
C14057 a_n1925_42282# a_n1899_43946# 1.14e-19
C14058 a_16680_45572# a_16922_45042# 5.89e-20
C14059 a_16855_45546# a_17023_45118# 4.36e-19
C14060 a_2382_45260# a_3232_43370# 0.239776f
C14061 a_2437_43646# a_1423_45028# 0.023818f
C14062 a_n755_45592# a_3363_44484# 8.3e-21
C14063 a_n2017_45002# a_9482_43914# 2.97e-21
C14064 a_4574_45260# a_4558_45348# 0.19344f
C14065 a_3537_45260# a_5147_45002# 0.092965f
C14066 a_3483_46348# a_15493_43396# 1.59e-19
C14067 a_16327_47482# a_18249_42858# 0.315855f
C14068 a_9049_44484# a_8701_44490# 0.100038f
C14069 a_7499_43078# a_5883_43914# 0.100372f
C14070 a_n443_42852# a_6109_44484# 0.002868f
C14071 a_n1079_45724# a_n2661_43922# 9.64e-21
C14072 a_584_46384# a_2981_46116# 6.74e-20
C14073 a_n1151_42308# a_n1533_46116# 0.002268f
C14074 a_6151_47436# a_6945_45028# 0.335681f
C14075 a_13717_47436# a_2324_44458# 1.33e-21
C14076 a_12861_44030# a_14840_46494# 7.53e-20
C14077 a_20916_46384# a_21363_46634# 0.017401f
C14078 a_19321_45002# a_20731_47026# 3.86e-21
C14079 a_13661_43548# a_17639_46660# 2.94e-20
C14080 a_5807_45002# a_18280_46660# 3.71e-20
C14081 a_n1613_43370# a_n1423_46090# 0.15966f
C14082 a_4883_46098# a_5497_46414# 0.007657f
C14083 a_11599_46634# a_13925_46122# 0.549622f
C14084 a_10227_46804# a_10355_46116# 0.022564f
C14085 a_8145_46902# a_8023_46660# 3.16e-19
C14086 a_7715_46873# a_8270_45546# 2.04e-19
C14087 a_n881_46662# a_n1991_46122# 0.001102f
C14088 a_2487_47570# a_167_45260# 9.29e-23
C14089 a_12549_44172# a_12741_44636# 0.090958f
C14090 a_4955_46873# a_3090_45724# 9.92e-20
C14091 a_n971_45724# a_5066_45546# 0.045749f
C14092 a_14311_47204# a_14275_46494# 4.74e-21
C14093 a_5649_42852# a_12089_42308# 3.26e-20
C14094 a_n3674_39768# a_n3420_39616# 0.073948f
C14095 a_n4318_39768# a_n2946_39866# 7.88e-20
C14096 a_16823_43084# a_18083_42858# 4.78e-20
C14097 a_4361_42308# a_12895_43230# 5.63e-20
C14098 a_5518_44484# VDD 0.40715f
C14099 a_15743_43084# a_22223_42860# 0.021215f
C14100 a_743_42282# a_15279_43071# 4.98e-21
C14101 a_4190_30871# a_15567_42826# 6.55e-21
C14102 a_n97_42460# a_1184_42692# 8.23e-20
C14103 a_18479_47436# a_20712_42282# 1.22e-20
C14104 a_18597_46090# a_13258_32519# 0.023292f
C14105 a_n755_45592# a_n2433_43396# 5.17e-20
C14106 a_n357_42282# a_n2129_43609# 0.001046f
C14107 a_n2661_43370# a_9838_44484# 1.69e-20
C14108 a_1307_43914# a_8375_44464# 3.91e-20
C14109 a_13259_45724# a_2982_43646# 0.06616f
C14110 a_6171_45002# a_14815_43914# 2.54e-21
C14111 a_20567_45036# a_20205_45028# 2.35e-20
C14112 a_413_45260# a_17517_44484# 0.013023f
C14113 a_n913_45002# a_11967_42832# 0.156551f
C14114 a_4185_45028# a_17364_32525# 0.046035f
C14115 a_5907_45546# a_5829_43940# 5.47e-21
C14116 a_n2293_45546# a_n97_42460# 2.89e-21
C14117 a_21513_45002# a_3422_30871# 9.94e-20
C14118 a_n863_45724# a_n1352_43396# 9.43e-21
C14119 a_1423_45028# a_4181_44734# 0.002332f
C14120 a_8953_45546# a_743_42282# 0.032209f
C14121 a_16327_47482# a_21125_42558# 5.5e-19
C14122 a_13507_46334# a_18214_42558# 1.84e-19
C14123 a_491_47026# a_310_45028# 9.66e-21
C14124 a_n743_46660# a_7_45899# 0.001065f
C14125 a_n2661_46098# a_n2293_45546# 4.48e-20
C14126 a_6755_46942# a_8049_45260# 0.035035f
C14127 a_14035_46660# a_2324_44458# 2.63e-20
C14128 a_15227_44166# a_10809_44734# 0.034868f
C14129 a_n2497_47436# a_2437_43646# 0.027407f
C14130 a_10227_46804# a_10544_45572# 0.00205f
C14131 a_171_46873# a_n356_45724# 5.68e-21
C14132 a_13059_46348# a_13351_46090# 0.074689f
C14133 a_n2293_46098# a_n1423_46090# 0.00572f
C14134 a_n2157_46122# a_n1991_46122# 0.614266f
C14135 a_765_45546# a_9823_46155# 1.78e-20
C14136 a_19466_46812# a_6945_45028# 2.92e-19
C14137 a_19692_46634# a_21137_46414# 0.242332f
C14138 a_n2293_46634# a_1609_45822# 0.036096f
C14139 a_5807_45002# a_6194_45824# 0.02442f
C14140 a_11599_46634# a_15599_45572# 0.26676f
C14141 a_5649_42852# a_18907_42674# 5.66e-20
C14142 a_20301_43646# a_20107_42308# 5.1e-21
C14143 a_4361_42308# a_18220_42308# 6.69e-19
C14144 a_17538_32519# a_22459_39145# 1.25e-20
C14145 a_14401_32519# a_22521_39511# 8.94e-21
C14146 a_743_42282# a_13258_32519# 0.030886f
C14147 a_4190_30871# a_20712_42282# 1.12e-20
C14148 a_8952_43230# a_9223_42460# 2.08e-19
C14149 a_9127_43156# a_9803_42558# 0.001572f
C14150 a_n2017_45002# a_6031_43396# 5.49e-20
C14151 a_11827_44484# a_11750_44172# 8.34e-20
C14152 a_n443_42852# a_15567_42826# 3.58e-19
C14153 a_n863_45724# a_n2293_42282# 0.028166f
C14154 a_4185_45028# a_8325_42308# 9.41e-20
C14155 a_3065_45002# a_4699_43561# 1.24e-20
C14156 a_2382_45260# a_4905_42826# 7.37e-21
C14157 a_n357_42282# a_21195_42852# 0.09377f
C14158 a_n2956_39304# a_n4318_37592# 0.023347f
C14159 a_16922_45042# a_20269_44172# 0.010825f
C14160 a_14815_43914# a_14673_44172# 0.173231f
C14161 a_n2267_44484# a_n1441_43940# 1.52e-19
C14162 a_5518_44484# a_5495_43940# 3.48e-20
C14163 a_18587_45118# a_18451_43940# 1.13e-20
C14164 a_3537_45260# a_4093_43548# 0.001642f
C14165 a_4223_44672# a_7542_44172# 0.052366f
C14166 a_5937_45572# a_6171_42473# 8.33e-22
C14167 a_n2956_38680# a_n1736_42282# 2.5e-20
C14168 a_8034_45724# a_8062_46155# 0.002525f
C14169 a_n2293_46634# a_501_45348# 1.32e-19
C14170 a_6945_45028# a_20205_31679# 0.00545f
C14171 a_20708_46348# a_20850_46155# 0.005572f
C14172 a_1823_45246# a_3733_45822# 0.003114f
C14173 a_6545_47178# a_6298_44484# 2.86e-20
C14174 a_11415_45002# a_12427_45724# 1.12e-20
C14175 a_5807_45002# a_6517_45366# 5.73e-19
C14176 a_3877_44458# a_3065_45002# 0.287919f
C14177 a_5167_46660# a_413_45260# 1.29e-20
C14178 a_5257_43370# a_n913_45002# 9.26e-20
C14179 a_13059_46348# a_15225_45822# 0.002175f
C14180 a_10249_46116# a_3357_43084# 5.65e-20
C14181 a_3090_45724# a_18909_45814# 7.08e-19
C14182 a_4791_45118# a_10334_44484# 1.31e-20
C14183 a_167_45260# a_3775_45552# 1.19e-20
C14184 a_3483_46348# a_6472_45840# 1.46e-20
C14185 a_n2497_47436# a_4181_44734# 0.01129f
C14186 a_5164_46348# a_2711_45572# 0.031464f
C14187 a_n743_46660# a_15595_45028# 2.81e-20
C14188 a_18597_46090# a_20193_45348# 0.021804f
C14189 a_13507_46334# a_21359_45002# 6.77e-19
C14190 a_14456_42282# a_15486_42560# 6.85e-20
C14191 a_n784_42308# a_1736_39587# 3.17e-20
C14192 a_17364_32525# VREF_GND 0.048253f
C14193 a_5742_30871# a_9885_42308# 1.65e-19
C14194 a_n3674_38216# a_n3420_39072# 0.020386f
C14195 a_n4318_38216# a_n4064_39072# 0.023072f
C14196 a_4921_42308# a_7174_31319# 1.72e-20
C14197 a_n1630_35242# a_n2302_39866# 5.02e-20
C14198 a_n1379_43218# VDD 1.08e-19
C14199 a_18184_42460# a_22591_43396# 8.5e-19
C14200 a_n2293_42834# a_5111_42852# 0.009675f
C14201 a_11823_42460# a_10545_42558# 1.52e-20
C14202 a_n2956_38216# a_n2946_39866# 4.86e-20
C14203 a_11827_44484# a_4361_42308# 1.05e-20
C14204 a_20193_45348# a_743_42282# 0.007306f
C14205 a_9028_43914# a_9672_43914# 2.65e-19
C14206 a_20640_44752# a_20974_43370# 2.23e-21
C14207 a_18579_44172# a_19319_43548# 0.031277f
C14208 a_5891_43370# a_8791_43396# 0.194389f
C14209 a_n2956_38680# a_n4209_37414# 1.36e-21
C14210 a_n913_45002# a_9114_42852# 4.02e-19
C14211 a_10193_42453# a_13070_42354# 1.07e-19
C14212 a_3537_45260# a_5457_43172# 0.001869f
C14213 a_12594_46348# a_13777_45326# 0.00118f
C14214 a_12861_44030# a_19478_44306# 2.84e-20
C14215 a_5907_45546# a_6229_45572# 0.007399f
C14216 a_5164_46348# a_4640_45348# 1.3e-19
C14217 a_8162_45546# a_7499_43078# 0.021916f
C14218 a_518_46482# a_413_45260# 1.79e-21
C14219 a_18280_46660# a_18315_45260# 4.34e-22
C14220 a_10227_46804# a_10949_43914# 2.49e-20
C14221 a_2711_45572# a_8336_45822# 2.46e-19
C14222 a_8199_44636# a_1423_45028# 0.088277f
C14223 a_2698_46116# a_2809_45028# 2.22e-20
C14224 a_11415_45002# a_14309_45028# 0.040538f
C14225 a_13259_45724# a_16789_45572# 9.06e-19
C14226 a_8049_45260# a_19479_31679# 0.022565f
C14227 a_768_44030# a_644_44056# 0.177755f
C14228 a_n1925_42282# en_comp 4.02e-19
C14229 a_2324_44458# a_10951_45334# 0.002224f
C14230 a_13759_46122# a_9482_43914# 1e-20
C14231 a_10227_46804# a_20894_47436# 0.010908f
C14232 a_18780_47178# a_18597_46090# 0.175179f
C14233 a_18479_47436# a_19386_47436# 0.219411f
C14234 a_n4209_39304# a_n3690_37440# 2.3e-19
C14235 a_n4209_38216# a_n2216_37984# 0.001433f
C14236 a_13070_42354# VDD 0.18656f
C14237 a_15673_47210# a_12465_44636# 6.52e-19
C14238 a_16327_47482# a_4883_46098# 0.096832f
C14239 a_n3565_39304# a_n4334_37440# 5.28e-19
C14240 a_n3690_38304# a_n3607_38304# 0.007692f
C14241 a_n2946_37984# a_n2302_37984# 6.68e-19
C14242 a_n1435_47204# a_n89_47570# 2.3e-21
C14243 a_5815_47464# a_n1613_43370# 0.360237f
C14244 a_16763_47508# a_13507_46334# 8.88e-21
C14245 a_4915_47217# a_7989_47542# 9.72e-19
C14246 a_n443_46116# a_4842_47243# 0.001129f
C14247 a_4791_45118# a_5159_47243# 0.00545f
C14248 a_n1151_42308# a_12891_46348# 0.038292f
C14249 a_2905_45572# a_768_44030# 0.02789f
C14250 a_n2288_47178# a_n2956_39768# 0.001146f
C14251 a_n2497_47436# a_n2661_46634# 0.079801f
C14252 a_n2833_47464# a_n2472_46634# 0.001084f
C14253 a_22465_38105# a_22459_39145# 0.98555f
C14254 a_20269_44172# a_15743_43084# 8.8e-21
C14255 a_15493_43940# a_16977_43638# 5.19e-19
C14256 a_11341_43940# a_17499_43370# 2.28e-19
C14257 a_15493_43396# a_16664_43396# 0.016417f
C14258 a_19279_43940# a_18083_42858# 9.26e-20
C14259 a_n2956_37592# a_n3565_38502# 0.024508f
C14260 a_6428_45938# VDD 4.6e-19
C14261 a_19478_44306# a_19700_43370# 0.008781f
C14262 a_895_43940# a_1847_42826# 2.53e-19
C14263 a_2479_44172# a_2075_43172# 0.034186f
C14264 a_742_44458# a_1184_42692# 1.39e-19
C14265 a_n699_43396# a_564_42282# 1.29e-22
C14266 a_n2129_43609# a_n144_43396# 7.58e-20
C14267 a_n97_42460# a_2896_43646# 0.027089f
C14268 a_n1699_43638# a_n1243_43396# 4.2e-19
C14269 a_1568_43370# a_1756_43548# 0.094732f
C14270 a_13661_43548# a_9145_43396# 0.135139f
C14271 a_8746_45002# a_8560_45348# 0.044092f
C14272 a_n2293_45546# a_742_44458# 1.34e-19
C14273 a_n2661_45546# a_4223_44672# 0.041115f
C14274 a_2711_45572# a_18494_42460# 0.1183f
C14275 a_4185_45028# a_19237_31679# 0.004066f
C14276 a_16327_47482# a_5649_42852# 9.95e-20
C14277 a_18985_46122# a_17517_44484# 2.43e-21
C14278 a_n863_45724# a_n1352_44484# 1.83e-21
C14279 a_n755_45592# a_n2433_44484# 4.6e-21
C14280 a_10809_44734# a_12189_44484# 1.06e-19
C14281 a_8568_45546# a_n2661_43370# 6.03e-21
C14282 a_8696_44636# a_8953_45002# 0.018854f
C14283 a_n2293_46098# a_3905_42865# 0.237656f
C14284 a_2437_43646# a_22591_45572# 2.94e-19
C14285 a_22223_45572# a_3357_43084# 0.07533f
C14286 a_21513_45002# a_19963_31679# 3.07e-19
C14287 a_18479_47436# a_20556_43646# 9.29e-19
C14288 a_13259_45724# a_14539_43914# 0.002022f
C14289 a_14033_45822# a_14180_45002# 2.17e-20
C14290 a_18479_47436# a_19551_46910# 0.001789f
C14291 a_n2661_46634# a_6682_46987# 4.03e-19
C14292 a_5807_45002# a_8601_46660# 1.44e-19
C14293 a_2063_45854# a_2202_46116# 0.026352f
C14294 a_12549_44172# a_13607_46688# 0.013421f
C14295 a_10227_46804# a_20411_46873# 0.013631f
C14296 a_2107_46812# a_5257_43370# 0.039927f
C14297 a_3524_46660# a_4651_46660# 1.59e-19
C14298 a_n971_45724# a_5068_46348# 3.37e-21
C14299 a_12465_44636# a_16388_46812# 7.04e-20
C14300 C5_N_btm C9_N_btm 0.153949f
C14301 C4_N_btm C10_N_btm 0.348092f
C14302 C6_N_btm C8_N_btm 0.170091f
C14303 a_18597_46090# a_18285_46348# 0.012666f
C14304 C2_N_btm VDD 0.268945f
C14305 a_n881_46662# a_15227_44166# 1.74e-19
C14306 C8_P_btm VIN_P 0.907642f
C14307 C10_P_btm VREF 14.773f
C14308 a_584_46384# a_167_45260# 0.0321f
C14309 a_n237_47217# a_4419_46090# 0.049065f
C14310 a_n743_46660# a_10150_46912# 4e-20
C14311 a_3699_46634# a_4955_46873# 2.52e-20
C14312 a_8685_43396# a_12089_42308# 3.95e-19
C14313 a_n2661_42282# a_7227_42308# 3.35e-19
C14314 a_19177_43646# a_19095_43396# 8.13e-19
C14315 a_21259_43561# a_21487_43396# 0.08444f
C14316 a_10695_43548# a_10083_42826# 0.005272f
C14317 a_19721_31679# a_22459_39145# 1.93e-20
C14318 a_20301_43646# a_743_42282# 0.09203f
C14319 a_4190_30871# a_20556_43646# 0.021112f
C14320 a_9145_43396# a_10835_43094# 4.2e-20
C14321 a_n1557_42282# a_873_42968# 8.49e-21
C14322 a_4093_43548# a_4649_43172# 0.001356f
C14323 a_16751_45260# a_16981_45144# 0.004937f
C14324 a_5205_44484# a_4223_44672# 0.235572f
C14325 a_n443_42852# a_10405_44172# 7.35e-20
C14326 a_n357_42282# a_15493_43396# 9.67e-20
C14327 a_n2661_45010# a_n356_44636# 0.091266f
C14328 a_n2017_45002# a_n1809_44850# 0.001936f
C14329 a_17339_46660# a_19095_43396# 0.049229f
C14330 w_11334_34010# a_13258_32519# 2.64e-19
C14331 a_5691_45260# a_5518_44484# 8.35e-19
C14332 a_3232_43370# a_5343_44458# 0.654021f
C14333 a_5111_44636# a_8103_44636# 0.001535f
C14334 a_n1613_43370# a_n961_42308# 0.0058f
C14335 w_1575_34946# a_n4064_38528# 7.84e-19
C14336 a_5807_45002# a_14371_46494# 0.002046f
C14337 a_n971_45724# a_6977_45572# 4.78e-20
C14338 a_n1151_42308# a_11322_45546# 0.001795f
C14339 a_10249_46116# a_9625_46129# 0.009289f
C14340 a_6755_46942# a_8953_45546# 0.001323f
C14341 a_6969_46634# a_5937_45572# 0.001066f
C14342 a_6151_47436# a_6812_45938# 0.018338f
C14343 a_4791_45118# a_9049_44484# 0.009879f
C14344 a_15673_47210# a_2711_45572# 2.77e-20
C14345 a_n1925_46634# a_8034_45724# 0.206805f
C14346 a_18285_46348# a_19123_46287# 0.007333f
C14347 a_2063_45854# a_11823_42460# 8.26e-19
C14348 a_12549_44172# a_16375_45002# 0.001412f
C14349 a_10467_46802# a_10355_46116# 0.008762f
C14350 a_10428_46928# a_9290_44172# 1.43e-19
C14351 a_3080_42308# a_1736_39587# 1.8e-19
C14352 a_743_42282# a_5421_42558# 0.001222f
C14353 a_n3674_39304# a_n1630_35242# 2.14e-19
C14354 a_2127_44172# VDD 0.138239f
C14355 a_19237_31679# VREF_GND 0.0061f
C14356 a_5649_42852# a_5267_42460# 0.016079f
C14357 a_3815_47204# VDD 0.260661f
C14358 a_n2661_43370# a_2998_44172# 9.42e-20
C14359 a_2553_47502# DATA[2] 2.89e-20
C14360 a_n863_45724# a_n1423_42826# 4.06e-21
C14361 a_13249_42308# a_13667_43396# 0.004219f
C14362 a_2952_47436# DATA[1] 7.06e-21
C14363 a_11827_44484# a_20397_44484# 3.81e-19
C14364 a_n2810_45572# a_n4318_38680# 0.023234f
C14365 a_22223_45036# a_22315_44484# 0.011923f
C14366 a_18114_32519# a_20640_44752# 9.12e-19
C14367 a_1307_43914# a_10949_43914# 0.062121f
C14368 a_n2293_42834# a_7542_44172# 0.010138f
C14369 a_14537_43396# a_14955_43940# 0.104291f
C14370 a_12607_44458# a_14815_43914# 6.91e-21
C14371 a_11322_45546# a_12293_43646# 9.9e-20
C14372 a_11823_42460# a_14955_43396# 5.12e-19
C14373 a_10903_43370# a_12991_43230# 0.001102f
C14374 a_8016_46348# a_8062_46155# 0.006879f
C14375 a_7920_46348# a_8379_46155# 6.64e-19
C14376 a_8199_44636# a_9823_46482# 1.73e-22
C14377 a_12469_46902# a_11823_42460# 2.61e-20
C14378 a_11901_46660# a_12791_45546# 8.23e-19
C14379 a_12251_46660# a_12427_45724# 1.4e-20
C14380 a_3090_45724# a_8746_45002# 1.22e-19
C14381 a_14976_45028# a_10193_42453# 1.31e-20
C14382 a_22612_30879# a_20447_31679# 0.107874f
C14383 a_12465_44636# a_13777_45326# 4.66e-20
C14384 a_10809_44734# a_22959_46124# 0.172346f
C14385 a_2324_44458# a_n1925_42282# 0.018757f
C14386 a_8953_45546# a_8049_45260# 0.156816f
C14387 a_n881_46662# a_4558_45348# 3.03e-21
C14388 a_n1613_43370# a_5147_45002# 1.57e-20
C14389 a_13507_46334# a_15415_45028# 1.22e-20
C14390 a_11453_44696# a_13159_45002# 0.006266f
C14391 a_13661_43548# a_n1059_45260# 0.004019f
C14392 a_5807_45002# a_n913_45002# 2.94e-20
C14393 a_12549_44172# a_413_45260# 2.22e-19
C14394 a_3823_42558# a_5934_30871# 1.35e-20
C14395 a_n784_42308# a_13070_42354# 1.96e-20
C14396 a_5379_42460# a_6123_31319# 0.011994f
C14397 a_5421_42558# a_5755_42308# 1.68e-19
C14398 a_13291_42460# a_7174_31319# 4.88e-21
C14399 a_n1630_35242# a_5742_30871# 1.85829f
C14400 a_4921_42308# a_5932_42308# 0.194195f
C14401 a_3065_45002# a_1847_42826# 2.79e-20
C14402 a_n443_42852# a_6171_42473# 6.33e-20
C14403 a_n2065_43946# a_n1441_43940# 9.73e-19
C14404 a_n1549_44318# a_n1453_44318# 0.013793f
C14405 a_n1331_43914# a_n1287_44306# 3.69e-19
C14406 a_n1899_43946# a_n875_44318# 2.36e-20
C14407 a_11967_42832# a_18451_43940# 0.01235f
C14408 a_n913_45002# a_10518_42984# 0.058603f
C14409 a_n2017_45002# a_10796_42968# 1.01e-19
C14410 a_n1059_45260# a_10835_43094# 0.004669f
C14411 a_16112_44458# a_n97_42460# 1.17e-19
C14412 a_5343_44458# a_4905_42826# 7.39e-21
C14413 a_742_44458# a_2896_43646# 8.3e-20
C14414 a_14976_45028# VDD 0.484864f
C14415 a_3090_45724# RST_Z 1.8e-20
C14416 a_2382_45260# a_2905_42968# 7.68e-19
C14417 a_11186_47026# CLK 6.21e-21
C14418 a_n984_44318# a_n3674_39768# 4.73e-20
C14419 a_n699_43396# a_n1557_42282# 0.02911f
C14420 a_n2661_42834# a_2455_43940# 0.002019f
C14421 a_14815_43914# a_14761_44260# 1.48e-19
C14422 a_n755_45592# a_8685_42308# 0.001582f
C14423 a_n357_42282# a_8791_42308# 6.28e-20
C14424 a_18479_47436# a_20980_44850# 0.002954f
C14425 a_3316_45546# a_2711_45572# 0.065336f
C14426 a_3218_45724# a_3175_45822# 0.132424f
C14427 a_13259_45724# a_12427_45724# 6.07e-19
C14428 a_12891_46348# a_13857_44734# 7.81e-20
C14429 a_768_44030# a_13213_44734# 0.00651f
C14430 a_9569_46155# a_2437_43646# 2.04e-20
C14431 a_13507_46334# a_19279_43940# 1.3e-20
C14432 a_10227_46804# a_3422_30871# 2.07e-19
C14433 a_19321_45002# a_9313_44734# 7.03e-21
C14434 a_n2661_45546# a_3260_45572# 6.42e-20
C14435 a_19553_46090# a_19431_45546# 8.55e-19
C14436 a_18985_46122# a_19256_45572# 5.12e-19
C14437 a_765_45546# a_1423_45028# 3.01e-22
C14438 a_805_46414# a_327_44734# 2.28e-19
C14439 a_4791_45118# a_3905_42865# 0.208831f
C14440 a_11453_44696# a_11967_42832# 6.13e-20
C14441 a_16327_47482# a_21145_44484# 1.79e-19
C14442 a_4185_45028# a_n1059_45260# 0.027781f
C14443 a_5937_45572# a_3357_43084# 0.257963f
C14444 a_n2293_46098# a_5147_45002# 0.211057f
C14445 a_5257_43370# a_n2661_44458# 0.027109f
C14446 a_4646_46812# a_5518_44484# 2.19e-19
C14447 a_10586_45546# a_10907_45822# 0.05477f
C14448 a_1609_45822# a_2277_45546# 2.47e-20
C14449 a_1431_47204# a_n1435_47204# 0.001005f
C14450 a_n443_46116# a_5129_47502# 0.10632f
C14451 a_4791_45118# a_5815_47464# 0.003581f
C14452 a_n1151_42308# a_7903_47542# 8.5e-20
C14453 a_2063_45854# a_9313_45822# 0.042979f
C14454 a_n4064_40160# a_n3420_38528# 0.057096f
C14455 a_n4209_39304# a_n4334_39392# 0.253307f
C14456 a_n4315_30879# a_n4064_38528# 0.034153f
C14457 a_n4318_38216# VDD 0.538766f
C14458 a_1606_42308# C6_P_btm 2.33e-19
C14459 a_n784_42308# C2_N_btm 0.005178f
C14460 a_n4209_39590# a_n4209_38502# 0.031979f
C14461 a_18579_44172# a_19095_43396# 1.8e-19
C14462 a_9313_44734# a_10922_42852# 0.002978f
C14463 a_n2293_42834# a_n1630_35242# 0.007885f
C14464 a_n2017_45002# a_4958_30871# 0.053522f
C14465 a_n1059_45260# a_16269_42308# 1.17e-19
C14466 a_18051_46116# VDD 0.189782f
C14467 a_n2661_43922# a_7871_42858# 7.71e-21
C14468 a_n2661_42834# a_7765_42852# 2.1e-21
C14469 a_20692_30879# C3_N_btm 3.19e-20
C14470 a_20205_31679# C4_N_btm 0.042623f
C14471 a_19479_31679# a_13258_32519# 0.054577f
C14472 a_n2661_42282# a_6643_43396# 1.74e-19
C14473 a_12861_44030# a_13667_43396# 5.08e-21
C14474 a_2711_45572# a_13777_45326# 0.008866f
C14475 a_10809_44734# a_9838_44484# 1.37e-19
C14476 a_n443_42852# a_1145_45348# 2.98e-20
C14477 a_10903_43370# a_n356_44636# 2.05e-19
C14478 a_8049_45260# a_20193_45348# 6.42e-20
C14479 a_7499_43078# a_3537_45260# 0.586701f
C14480 a_17583_46090# a_17767_44458# 1.63e-20
C14481 a_310_45028# a_117_45144# 2.88e-35
C14482 a_8016_46348# a_8375_44464# 1.63e-20
C14483 a_13259_45724# a_14309_45028# 0.063402f
C14484 a_1823_45246# a_n2661_43922# 0.441151f
C14485 a_12741_44636# a_17061_44734# 0.003447f
C14486 a_16680_45572# a_17668_45572# 1.69e-19
C14487 a_3090_45724# a_5663_43940# 0.001711f
C14488 a_8696_44636# a_17568_45572# 2.55e-19
C14489 a_1138_42852# a_n2293_43922# 9.77e-21
C14490 a_8199_44636# a_6109_44484# 1.61e-22
C14491 a_17715_44484# a_16979_44734# 0.005407f
C14492 a_3754_38470# RST_Z 0.203816f
C14493 VDAC_P C7_P_btm 30.8442f
C14494 a_22609_37990# a_22705_37990# 0.087835f
C14495 a_768_44030# a_2443_46660# 2.94e-19
C14496 a_n2661_46634# a_n2104_46634# 0.030211f
C14497 a_n2472_46634# a_n2293_46634# 0.163804f
C14498 a_n1151_42308# a_12359_47026# 0.002059f
C14499 a_n1613_43370# a_3055_46660# 9.54e-19
C14500 a_4883_46098# a_8667_46634# 2.2e-19
C14501 a_n2497_47436# a_765_45546# 1.79e-20
C14502 a_n1435_47204# a_11735_46660# 7.87e-20
C14503 a_5807_45002# a_2107_46812# 1.5594f
C14504 a_n2956_39768# a_n2312_38680# 0.076511f
C14505 a_n2840_46634# a_n1925_46634# 5.18e-19
C14506 a_8147_43396# a_4361_42308# 2.94e-21
C14507 a_10341_43396# a_17499_43370# 0.022768f
C14508 a_n97_42460# a_7227_42852# 0.117893f
C14509 a_2382_45260# VDD 1.6285f
C14510 a_9145_43396# a_15037_43396# 5.99e-20
C14511 a_8685_43396# a_16855_43396# 8.49e-20
C14512 a_1414_42308# a_n3674_37592# 2.19e-21
C14513 a_9313_44734# a_17531_42308# 4.72e-20
C14514 a_9290_44172# a_10651_43940# 3.97e-19
C14515 a_12427_45724# a_n2661_43922# 1.65e-19
C14516 a_11823_42460# a_n2661_42834# 4.26e-20
C14517 a_5205_44484# a_n2293_42834# 4.84e-20
C14518 a_21363_45546# a_19721_31679# 2.83e-19
C14519 a_1138_42852# a_n97_42460# 0.015603f
C14520 a_7499_43078# a_11541_44484# 0.048175f
C14521 a_6171_45002# a_8488_45348# 8.23e-19
C14522 a_8696_44636# a_17767_44458# 3.64e-19
C14523 a_4574_45260# a_n2661_43370# 0.007993f
C14524 a_20202_43084# a_2982_43646# 0.034798f
C14525 a_n2293_46634# a_5534_30871# 9.88e-20
C14526 a_n1151_42308# a_564_42282# 3.17e-20
C14527 a_13661_43548# a_19987_42826# 1.73e-19
C14528 a_3090_45724# a_16243_43396# 1.04e-20
C14529 a_19963_31679# a_22959_45036# 0.002114f
C14530 a_n2293_45546# a_n984_44318# 1.81e-20
C14531 a_n1079_45724# a_n809_44244# 8.53e-21
C14532 a_15861_45028# a_16979_44734# 4.51e-19
C14533 a_5807_45002# a_14493_46090# 0.006666f
C14534 a_13747_46662# a_13759_46122# 0.02887f
C14535 a_13661_43548# a_13925_46122# 2.91e-21
C14536 a_12549_44172# a_18985_46122# 1.04e-20
C14537 a_n743_46660# a_6419_46155# 0.00636f
C14538 a_584_46384# a_n863_45724# 0.051089f
C14539 a_n2661_46098# a_1138_42852# 0.020229f
C14540 a_17609_46634# a_15227_44166# 0.04317f
C14541 a_n785_47204# a_n755_45592# 1.12e-20
C14542 a_327_47204# a_n357_42282# 1.62e-22
C14543 a_n1925_46634# a_8016_46348# 0.014574f
C14544 a_11735_46660# a_13885_46660# 5.87e-21
C14545 a_12251_46660# a_12347_46660# 0.013793f
C14546 a_12469_46902# a_12513_46660# 3.69e-19
C14547 a_11901_46660# a_12925_46660# 2.36e-20
C14548 a_4883_46098# a_6640_46482# 2.25e-19
C14549 a_18780_47178# a_8049_45260# 2.82e-21
C14550 a_11599_46634# a_12638_46436# 0.006285f
C14551 a_n971_45724# a_3218_45724# 2.69e-19
C14552 a_n237_47217# a_1848_45724# 0.232571f
C14553 a_2107_46812# a_3699_46348# 0.00528f
C14554 a_1799_45572# a_1823_45246# 0.003001f
C14555 a_n2661_46634# a_9569_46155# 8.52e-20
C14556 a_n2293_46634# a_5937_45572# 2.05e-19
C14557 a_6682_46987# a_765_45546# 3.8e-19
C14558 a_n1613_43370# a_n2956_39304# 4.39e-21
C14559 a_n97_42460# a_11633_42308# 0.00291f
C14560 a_7287_43370# a_6123_31319# 2.73e-19
C14561 a_7112_43396# a_7227_42308# 4.93e-21
C14562 a_15433_44458# VDD 0.201121f
C14563 a_19237_31679# a_22469_40625# 1.24e-20
C14564 a_3422_30871# CAL_P 0.083836f
C14565 a_15743_43084# a_20836_43172# 3.08e-19
C14566 a_5534_30871# a_5342_30871# 11.128201f
C14567 a_n443_42852# a_3457_43396# 0.009582f
C14568 a_n913_45002# a_n822_43940# 1.95e-19
C14569 a_10903_43370# a_12379_42858# 0.02509f
C14570 a_n2956_39768# a_7174_31319# 5.27e-21
C14571 a_5343_44458# a_8975_43940# 1.49e-20
C14572 a_n4318_40392# a_n2012_44484# 7.25e-20
C14573 a_18184_42460# a_9313_44734# 0.069472f
C14574 a_n1925_42282# a_n2157_42858# 1.51e-19
C14575 a_17339_46660# a_18504_43218# 6.4e-19
C14576 a_9290_44172# a_12895_43230# 3.44e-20
C14577 a_4185_45028# a_19987_42826# 3.48e-20
C14578 a_13259_45724# a_17324_43396# 2.64e-19
C14579 a_3537_45260# a_3600_43914# 0.157156f
C14580 a_4574_45260# a_2998_44172# 1.08e-19
C14581 a_2698_46116# a_2324_44458# 5.34e-22
C14582 a_n2472_46090# a_n2956_38680# 0.157373f
C14583 a_n2293_46098# a_n2956_39304# 0.001354f
C14584 a_18285_46348# a_8049_45260# 3.95e-19
C14585 a_12549_44172# a_12561_45572# 0.001714f
C14586 a_15227_44166# a_19443_46116# 7.48e-19
C14587 a_6575_47204# a_413_45260# 2.11e-19
C14588 a_4651_46660# a_4880_45572# 1.53e-20
C14589 a_13661_43548# a_15599_45572# 0.01321f
C14590 a_5807_45002# a_15903_45785# 5.55e-20
C14591 a_5937_45572# a_9625_46129# 1.78e-19
C14592 a_8199_44636# a_9569_46155# 1.7e-19
C14593 a_13747_46662# a_15297_45822# 0.001012f
C14594 a_2063_45854# a_7705_45326# 5.97e-19
C14595 a_14035_46660# a_12839_46116# 3.7e-20
C14596 a_13059_46348# a_12005_46436# 1.79e-21
C14597 a_5257_43370# a_5907_45546# 0.064039f
C14598 a_n443_46116# a_4558_45348# 1.56e-19
C14599 a_4791_45118# a_5147_45002# 0.10845f
C14600 a_18479_47436# a_3357_43084# 0.292061f
C14601 a_19386_47436# a_2437_43646# 0.00484f
C14602 a_n1655_43396# VDD 8.44e-20
C14603 a_19339_43156# a_17303_42282# 4.17e-21
C14604 a_n4318_37592# a_n1329_42308# 7.71e-21
C14605 a_n3674_38680# a_n3674_37592# 0.028019f
C14606 a_n4318_38216# a_n784_42308# 3.7e-22
C14607 a_18249_42858# a_18727_42674# 6.54e-20
C14608 a_3080_42308# C2_N_btm 0.108823f
C14609 a_n2810_45572# a_n2840_42282# 2.3e-20
C14610 a_5111_44636# a_10149_43396# 0.001625f
C14611 a_n2661_46098# DATA[1] 9e-20
C14612 a_949_44458# a_1241_43940# 3.56e-19
C14613 a_18443_44721# a_15493_43396# 1.69e-21
C14614 a_n2661_43922# a_n3674_39768# 0.152656f
C14615 a_18989_43940# a_18451_43940# 0.114286f
C14616 a_n2661_42834# a_n1644_44306# 0.006513f
C14617 a_n2293_43922# a_n4318_39768# 3.58e-19
C14618 a_5891_43370# a_6756_44260# 4.32e-21
C14619 a_20679_44626# a_20512_43084# 0.003019f
C14620 a_20835_44721# a_21145_44484# 0.013793f
C14621 a_20766_44850# a_21073_44484# 3.69e-19
C14622 a_19279_43940# a_20637_44484# 9.22e-19
C14623 a_20640_44752# a_22485_44484# 8.77e-20
C14624 en_comp a_15743_43084# 5.37e-21
C14625 a_21513_45002# a_21487_43396# 9.71e-22
C14626 a_10440_44484# a_10555_44260# 0.001321f
C14627 a_3524_46660# VDD 0.278519f
C14628 a_7640_43914# a_7911_44260# 1.97e-19
C14629 a_8696_44636# a_8037_42858# 2.6e-21
C14630 a_n357_42282# a_18707_42852# 0.003328f
C14631 a_18184_42460# a_20974_43370# 3.83e-20
C14632 a_14537_43396# a_8685_43396# 0.007467f
C14633 a_15004_44636# a_11341_43940# 2.28e-20
C14634 a_11967_42832# a_19237_31679# 2.2e-20
C14635 a_5807_45002# a_n2661_44458# 1.89e-19
C14636 a_5937_45572# a_9159_45572# 0.048183f
C14637 a_8199_44636# a_10216_45572# 4.45e-19
C14638 a_5066_45546# a_2711_45572# 0.090644f
C14639 a_6945_45028# a_9049_44484# 2.27e-20
C14640 a_768_44030# a_949_44458# 0.002011f
C14641 a_3090_45724# a_3232_43370# 0.024183f
C14642 a_12741_44636# a_19431_45546# 3.15e-20
C14643 a_2324_44458# a_13527_45546# 0.001831f
C14644 a_14275_46494# a_14495_45572# 0.003638f
C14645 a_11189_46129# a_10907_45822# 0.021145f
C14646 a_9290_44172# a_11280_45822# 2.36e-19
C14647 a_19321_45002# a_18114_32519# 1.08e-21
C14648 a_1709_42852# VDD 0.001589f
C14649 a_19511_42282# a_20712_42282# 0.05034f
C14650 a_5934_30871# a_1177_38525# 1.19e-19
C14651 a_19647_42308# a_20107_42308# 4.99e-19
C14652 a_17303_42282# a_22465_38105# 3.32e-19
C14653 a_18907_42674# a_18997_42308# 0.004764f
C14654 a_n4318_37592# a_n3690_37440# 1.65e-19
C14655 a_10729_43914# a_11173_43940# 0.00134f
C14656 a_10949_43914# a_10867_43940# 3.29e-19
C14657 a_10807_43548# a_10651_43940# 3.34e-19
C14658 a_1467_44172# a_n1557_42282# 7.5e-21
C14659 a_n699_43396# a_3935_42891# 9.41e-22
C14660 a_4223_44672# a_4520_42826# 6.71e-22
C14661 a_2382_45260# a_n784_42308# 1.58e-20
C14662 a_n2017_45002# a_2725_42558# 6.21e-19
C14663 a_19900_46494# VDD 0.279179f
C14664 a_19335_46494# START 6.85e-21
C14665 a_20075_46420# RST_Z 3.65e-21
C14666 a_14840_46494# CLK 5.5e-21
C14667 a_11827_44484# a_17595_43084# 1.44e-20
C14668 a_11691_44458# a_5342_30871# 1.35e-19
C14669 en_comp a_1606_42308# 0.022666f
C14670 a_11967_42832# a_9145_43396# 8.37e-19
C14671 a_15493_43940# a_15301_44260# 1.97e-19
C14672 a_18494_42460# a_18817_42826# 5.74e-19
C14673 a_18184_42460# a_18599_43230# 1.68e-19
C14674 a_9313_44734# a_15868_43402# 6.39e-20
C14675 a_n356_44636# a_5649_42852# 0.023625f
C14676 a_9290_44172# a_11827_44484# 1.72e-19
C14677 a_14495_45572# a_15765_45572# 1.19e-20
C14678 a_n443_46116# a_1756_43548# 0.046156f
C14679 a_584_46384# a_3540_43646# 0.045907f
C14680 a_n1151_42308# a_n1557_42282# 0.214486f
C14681 a_3699_46348# a_n2661_44458# 3.05e-21
C14682 a_1176_45822# a_949_44458# 4.19e-19
C14683 a_11415_45002# a_16112_44458# 2.93e-20
C14684 a_1138_42852# a_742_44458# 0.040731f
C14685 a_10490_45724# a_12749_45572# 4.85e-22
C14686 a_n443_42852# a_3357_43084# 0.042246f
C14687 a_768_44030# a_11341_43940# 0.005879f
C14688 a_12549_44172# a_22223_43948# 6.97e-19
C14689 a_2324_44458# a_16922_45042# 6.23e-21
C14690 a_n2661_45546# a_413_45260# 0.022797f
C14691 a_n755_45592# a_n913_45002# 0.347782f
C14692 a_n2293_46634# a_8333_44056# 2.16e-20
C14693 a_4883_46098# a_9165_43940# 0.00241f
C14694 a_10809_44734# a_n2661_43370# 0.077978f
C14695 a_15143_45578# a_15903_45785# 8.61e-19
C14696 a_10907_45822# a_11136_45572# 0.080042f
C14697 a_12741_44636# a_13076_44458# 0.010522f
C14698 a_n2293_45546# a_n467_45028# 0.067105f
C14699 a_13059_46348# a_9313_44734# 3.57e-19
C14700 a_13661_43548# a_18326_43940# 0.024789f
C14701 a_526_44458# a_2809_45028# 0.033247f
C14702 a_n4209_37414# a_n3420_37440# 0.245806f
C14703 a_n4334_37440# a_n3690_37440# 8.67e-19
C14704 a_11453_44696# a_5807_45002# 0.050036f
C14705 a_13507_46334# a_20916_46384# 0.123008f
C14706 a_21177_47436# a_21588_30879# 3.24e-19
C14707 a_n971_45724# a_7577_46660# 0.523694f
C14708 a_n1741_47186# a_9863_46634# 4.44e-20
C14709 a_4007_47204# a_3877_44458# 0.002042f
C14710 a_n443_46116# a_3686_47026# 4.1e-19
C14711 a_1239_39587# VDD 0.530104f
C14712 a_12465_44636# a_19321_45002# 4.94e-19
C14713 a_n4209_38502# C6_P_btm 0.001141f
C14714 a_n3565_38502# C8_P_btm 1.65e-20
C14715 a_n4315_30879# VREF_GND 0.168163f
C14716 a_n3565_38216# a_n1838_35608# 1.01e-19
C14717 a_n4209_38216# a_n1532_35090# 1.2e-19
C14718 a_n1151_42308# a_4817_46660# 0.029921f
C14719 a_n237_47217# a_7411_46660# 0.033907f
C14720 a_2063_45854# a_6540_46812# 1.36e-19
C14721 a_n881_46662# a_7989_47542# 2.79e-20
C14722 a_20193_45348# a_13258_32519# 0.001033f
C14723 a_n2661_42834# a_961_42354# 1.54e-21
C14724 a_n2293_43922# a_1576_42282# 8.6e-20
C14725 a_n356_44636# a_7963_42308# 1.17e-19
C14726 a_3905_42865# a_3059_42968# 4.87e-20
C14727 a_n97_42460# a_17499_43370# 0.005876f
C14728 a_6765_43638# a_7221_43396# 4.2e-19
C14729 a_3626_43646# a_14205_43396# 3.91e-21
C14730 a_2982_43646# a_14955_43396# 1.35e-20
C14731 a_3065_45002# a_5111_44636# 9.21e-21
C14732 a_8953_45546# a_9028_43914# 0.01093f
C14733 a_8016_46348# a_10949_43914# 3.79e-20
C14734 a_8199_44636# a_10405_44172# 1.31e-19
C14735 a_10227_46804# a_16414_43172# 4.57e-21
C14736 a_12861_44030# a_21195_42852# 1.78e-21
C14737 a_n1925_42282# a_n1761_44111# 5.08e-20
C14738 a_3090_45724# a_4905_42826# 4.85e-19
C14739 a_16855_45546# a_16922_45042# 0.002263f
C14740 a_n1613_43370# a_685_42968# 2.27e-20
C14741 a_3537_45260# a_4558_45348# 0.236111f
C14742 a_7499_43078# a_8701_44490# 0.011795f
C14743 a_n2293_45546# a_n2661_43922# 2.12e-19
C14744 a_n2956_38216# a_n2293_43922# 2.59e-20
C14745 a_4791_45118# a_5457_43172# 2.47e-19
C14746 a_22612_30879# a_13467_32519# 0.061222f
C14747 a_16327_47482# a_17333_42852# 0.006539f
C14748 SMPL_ON_N a_4185_45028# 3.43e-19
C14749 a_584_46384# a_1431_46436# 3.89e-19
C14750 a_4915_47217# a_10809_44734# 0.037616f
C14751 a_5815_47464# a_6945_45028# 9.9e-19
C14752 a_12861_44030# a_15015_46420# 7.95e-20
C14753 a_13717_47436# a_14840_46494# 2.21e-21
C14754 a_20916_46384# a_20623_46660# 9.66e-19
C14755 a_19321_45002# a_20528_46660# 3.62e-19
C14756 a_5807_45002# a_17639_46660# 4.64e-19
C14757 a_4883_46098# a_5204_45822# 0.041898f
C14758 a_14955_47212# a_13925_46122# 4.01e-20
C14759 a_11599_46634# a_13759_46122# 0.262969f
C14760 a_10227_46804# a_9823_46155# 0.004734f
C14761 a_8145_46902# a_8654_47026# 2.6e-19
C14762 a_7577_46660# a_8023_46660# 2.28e-19
C14763 a_4651_46660# a_3090_45724# 9.87e-21
C14764 a_n881_46662# a_n1853_46287# 0.229188f
C14765 a_n1613_43370# a_n1991_46122# 0.031697f
C14766 a_12891_46348# a_12741_44636# 0.038901f
C14767 a_7411_46660# a_8270_45546# 1.1e-19
C14768 a_10249_46116# a_6755_46942# 0.068878f
C14769 a_5649_42852# a_12379_42858# 5.88e-20
C14770 a_n4318_39768# a_n3420_39616# 0.002167f
C14771 a_16823_43084# a_17701_42308# 2.64e-19
C14772 a_4361_42308# a_13113_42826# 1.92e-20
C14773 a_n3674_39768# a_n3690_39616# 0.07198f
C14774 a_5343_44458# VDD 0.49245f
C14775 a_4190_30871# a_5342_30871# 0.0276f
C14776 a_743_42282# a_5534_30871# 0.030281f
C14777 a_15743_43084# a_22165_42308# 0.008223f
C14778 a_n2956_39768# a_5932_42308# 4.83e-21
C14779 a_11652_45724# a_11341_43940# 8.54e-21
C14780 a_n357_42282# a_n2433_43396# 2.74e-19
C14781 a_n2661_43370# a_5883_43914# 1.78e-19
C14782 a_n1059_45260# a_11967_42832# 0.627158f
C14783 a_10227_46804# a_7174_31319# 2.63e-20
C14784 a_7499_43078# a_11816_44260# 0.002269f
C14785 a_1307_43914# a_7640_43914# 0.006778f
C14786 a_8953_45002# a_9159_44484# 1.62e-19
C14787 a_18494_42460# a_20205_45028# 0.001453f
C14788 a_n863_45724# a_n1177_43370# 5.65e-20
C14789 a_4185_45028# a_22959_43396# 0.01521f
C14790 a_2324_44458# a_15743_43084# 9.18e-19
C14791 a_13507_46334# a_19332_42282# 0.001224f
C14792 a_2107_46812# a_n755_45592# 4.66e-20
C14793 a_948_46660# a_997_45618# 7.48e-19
C14794 a_n133_46660# a_n356_45724# 1.93e-19
C14795 a_n743_46660# a_n310_45899# 1.97e-19
C14796 a_288_46660# a_310_45028# 2.47e-19
C14797 a_19321_45002# a_2711_45572# 1.76e-19
C14798 a_1799_45572# a_n2293_45546# 4.04e-20
C14799 a_n2661_46098# a_n2956_38216# 0.001609f
C14800 a_10249_46116# a_8049_45260# 0.001129f
C14801 a_14513_46634# a_14275_46494# 0.001809f
C14802 a_19333_46634# a_6945_45028# 9.77e-20
C14803 a_18834_46812# a_10809_44734# 0.006086f
C14804 a_15227_44166# a_22223_46124# 0.002009f
C14805 a_14035_46660# a_14840_46494# 5.47e-21
C14806 a_765_45546# a_9569_46155# 2.88e-20
C14807 a_2609_46660# a_n2661_45546# 1.76e-20
C14808 a_13059_46348# a_12594_46348# 0.03479f
C14809 a_n2293_46098# a_n1991_46122# 0.01544f
C14810 a_n2157_46122# a_n1853_46287# 0.617317f
C14811 a_n1613_43370# a_7499_43078# 0.324998f
C14812 a_19692_46634# a_20708_46348# 0.318388f
C14813 a_5807_45002# a_5907_45546# 0.013402f
C14814 a_n2293_46634# a_n443_42852# 2.09483f
C14815 a_5649_42852# a_18727_42674# 1.1e-19
C14816 a_14209_32519# a_4958_30871# 0.030901f
C14817 a_10341_42308# a_5934_30871# 3.73e-20
C14818 a_4190_30871# a_20107_42308# 2.08e-20
C14819 a_n2293_42282# a_961_42354# 2.32e-19
C14820 a_4361_42308# a_18214_42558# 9.81e-20
C14821 a_743_42282# a_19647_42308# 0.005892f
C14822 a_8952_43230# a_8791_42308# 6.34e-19
C14823 a_9127_43156# a_9223_42460# 0.001251f
C14824 a_4223_44672# a_7281_43914# 0.01814f
C14825 a_n1059_45260# a_648_43396# 1.51e-19
C14826 a_n443_42852# a_5342_30871# 2.41e-19
C14827 a_2747_46873# DATA[2] 5.46e-20
C14828 a_7229_43940# a_n97_42460# 6.25e-19
C14829 a_2382_45260# a_3080_42308# 0.006891f
C14830 a_3065_45002# a_4235_43370# 2.44e-20
C14831 a_7_47243# DATA[0] 0.001094f
C14832 a_3357_43084# a_6655_43762# 3.75e-19
C14833 a_n357_42282# a_21356_42826# 0.156735f
C14834 a_14112_44734# a_14673_44172# 5.17e-20
C14835 a_5518_44484# a_5013_44260# 1.4e-19
C14836 a_5343_44458# a_5495_43940# 7.49e-21
C14837 a_5883_43914# a_2998_44172# 7.17e-21
C14838 a_17613_45144# a_15493_43396# 1.5e-21
C14839 a_16922_45042# a_19862_44208# 0.038132f
C14840 a_n2956_38680# a_n3674_38216# 0.02335f
C14841 a_n2956_39304# a_n1736_42282# 2.99e-20
C14842 a_11453_44696# a_18315_45260# 0.010513f
C14843 a_5066_45546# a_10037_46155# 9.67e-23
C14844 a_n2293_46634# a_375_42282# 0.004296f
C14845 a_21137_46414# a_20205_31679# 2.27e-19
C14846 a_1823_45246# a_3638_45822# 0.003923f
C14847 a_6151_47436# a_6298_44484# 1.58e-19
C14848 a_n881_46662# a_n2661_43370# 0.020731f
C14849 a_4883_46098# a_20567_45036# 1.52e-20
C14850 a_5807_45002# a_6125_45348# 0.00337f
C14851 a_5385_46902# a_413_45260# 1.97e-20
C14852 a_3877_44458# a_2680_45002# 2.18e-20
C14853 a_13059_46348# a_15037_45618# 0.064109f
C14854 a_5257_43370# a_n1059_45260# 2.6e-19
C14855 a_10554_47026# a_3357_43084# 2.24e-20
C14856 a_3090_45724# a_18341_45572# 0.016963f
C14857 a_6969_46634# a_2437_43646# 5.02e-20
C14858 a_4791_45118# a_10157_44484# 5.67e-20
C14859 a_4419_46090# a_4099_45572# 0.002575f
C14860 a_n2497_47436# a_700_44734# 3.92e-21
C14861 a_5068_46348# a_2711_45572# 9.3e-19
C14862 a_n743_46660# a_15415_45028# 3.05e-20
C14863 a_18597_46090# a_11691_44458# 2.38e-20
C14864 a_14456_42282# a_15051_42282# 2.66e-19
C14865 a_n784_42308# a_1239_39587# 6.81e-20
C14866 a_14209_32519# VCM 0.007464f
C14867 COMP_P a_n4209_39304# 1.25e-21
C14868 a_n4318_37592# a_n4334_39392# 7.52e-20
C14869 a_n1630_35242# a_n4064_39616# 7.67e-20
C14870 a_n1545_43230# VDD 1.95e-19
C14871 a_5891_43370# a_8147_43396# 0.029069f
C14872 a_18184_42460# a_13887_32519# 0.03303f
C14873 a_n2293_42834# a_4520_42826# 0.01065f
C14874 a_n2956_38216# a_n3420_39616# 1.85e-19
C14875 a_11827_44484# a_13467_32519# 1.16e-20
C14876 a_12741_44636# SINGLE_ENDED 1.02e-19
C14877 a_14539_43914# a_14955_43396# 0.00238f
C14878 a_2711_45572# a_17531_42308# 2.41e-21
C14879 a_644_44056# a_726_44056# 0.004767f
C14880 a_20679_44626# a_21381_43940# 0.001413f
C14881 a_18579_44172# a_19808_44306# 3.69e-19
C14882 a_n1059_45260# a_9114_42852# 1.72e-19
C14883 a_n2810_45572# a_n2302_39866# 2.61e-19
C14884 a_n356_44636# a_8685_43396# 2.93e-20
C14885 a_10193_42453# a_12563_42308# 2.67e-19
C14886 a_3537_45260# a_5193_43172# 0.003266f
C14887 a_20193_45348# a_20301_43646# 0.005382f
C14888 a_21076_30879# RST_Z 0.052228f
C14889 a_11599_46634# a_18079_43940# 3.46e-21
C14890 a_10903_43370# a_14180_45002# 0.008124f
C14891 a_13351_46090# a_9482_43914# 2.3e-19
C14892 a_12594_46348# a_13556_45296# 1.95e-21
C14893 a_5164_46348# a_4185_45348# 4.37e-22
C14894 a_8162_45546# a_8568_45546# 0.078784f
C14895 a_7230_45938# a_7499_43078# 2.81e-21
C14896 a_3090_45724# a_8975_43940# 0.003577f
C14897 a_19240_46482# a_18691_45572# 2.45e-19
C14898 a_8049_45260# a_22223_45572# 0.013885f
C14899 a_10227_46804# a_10729_43914# 3.09e-19
C14900 a_2324_44458# a_10775_45002# 0.003159f
C14901 a_2711_45572# a_6977_45572# 0.001232f
C14902 a_11415_45002# a_13807_45067# 0.001105f
C14903 a_12861_44030# a_15493_43396# 0.254093f
C14904 a_768_44030# a_175_44278# 6.16e-19
C14905 a_n1925_42282# a_n2956_37592# 2.26e-20
C14906 a_10227_46804# a_19787_47423# 0.03269f
C14907 a_18479_47436# a_18597_46090# 0.473843f
C14908 a_n4209_39304# a_n3565_37414# 0.030571f
C14909 a_12563_42308# VDD 0.254292f
C14910 a_15811_47375# a_12465_44636# 5.18e-19
C14911 a_16241_47178# a_4883_46098# 3.3e-21
C14912 a_n3565_39304# a_n4209_37414# 0.028483f
C14913 a_n2946_37984# a_n4064_37984# 0.053263f
C14914 a_n3565_38216# a_n3607_38304# 0.001003f
C14915 a_n3420_37984# a_n2302_37984# 2.4e-19
C14916 a_n1435_47204# a_n310_47570# 3.53e-21
C14917 a_5129_47502# a_n1613_43370# 0.002387f
C14918 a_16023_47582# a_13507_46334# 1.53e-21
C14919 a_16327_47482# a_21496_47436# 4.85e-21
C14920 a_4915_47217# a_n881_46662# 1.23372f
C14921 a_4700_47436# a_5159_47243# 6.64e-19
C14922 a_4791_45118# a_4842_47243# 0.006879f
C14923 a_n1151_42308# a_11309_47204# 0.546434f
C14924 a_n2497_47436# a_n2956_39768# 7.4e-19
C14925 a_n2833_47464# a_n2661_46634# 0.011033f
C14926 a_22465_38105# a_22521_40055# 0.214039f
C14927 a_15493_43940# a_16409_43396# 0.004011f
C14928 a_11341_43940# a_16759_43396# 1.49e-20
C14929 a_15493_43396# a_19700_43370# 0.001674f
C14930 a_n2661_42282# a_4361_42308# 0.034761f
C14931 en_comp a_n4209_38502# 0.006885f
C14932 a_4880_45572# VDD 0.004682f
C14933 a_19862_44208# a_15743_43084# 0.022478f
C14934 a_8333_44056# a_743_42282# 9.61e-22
C14935 a_2127_44172# a_2075_43172# 8.71e-21
C14936 a_2479_44172# a_1847_42826# 0.141223f
C14937 a_1414_42308# a_3681_42891# 0.001924f
C14938 a_895_43940# a_791_42968# 5.63e-21
C14939 a_11967_42832# a_19987_42826# 9.2e-21
C14940 a_742_44458# a_1576_42282# 8.56e-19
C14941 a_9313_44734# a_11554_42852# 0.001434f
C14942 a_n699_43396# a_n3674_37592# 3.66e-22
C14943 a_5343_44458# a_n784_42308# 1.26e-20
C14944 a_n2810_45028# a_n3565_38502# 0.031875f
C14945 a_19478_44306# a_19268_43646# 9.35e-20
C14946 a_n1809_43762# a_n1557_42282# 3.46e-21
C14947 a_n2267_43396# a_n1243_43396# 2.36e-20
C14948 a_n2129_43609# a_n998_43396# 0.002155f
C14949 a_n97_42460# a_1987_43646# 5.54e-19
C14950 a_5807_45002# a_9145_43396# 1.15e-19
C14951 a_15037_45618# a_13556_45296# 1.52e-19
C14952 a_n1079_45724# a_n1352_44484# 1.48e-20
C14953 a_n2293_45546# a_n452_44636# 1.06e-19
C14954 a_2711_45572# a_18184_42460# 0.367034f
C14955 a_10180_45724# a_10903_45394# 8.17e-20
C14956 a_n2293_46634# a_6655_43762# 0.003277f
C14957 w_11334_34010# a_5534_30871# 0.002185f
C14958 a_768_44030# a_10341_43396# 1.28e-19
C14959 a_n755_45592# a_n2661_44458# 0.023853f
C14960 a_n863_45724# a_n1177_44458# 1.65e-20
C14961 a_18819_46122# a_17517_44484# 5.47e-21
C14962 a_7499_43078# a_8704_45028# 0.001053f
C14963 a_4185_45028# a_22959_44484# 0.011365f
C14964 a_2437_43646# a_3357_43084# 0.424652f
C14965 a_22223_45572# a_19479_31679# 0.155323f
C14966 a_18597_46090# a_4190_30871# 0.022042f
C14967 a_n2661_45546# a_2779_44458# 4.85e-20
C14968 a_13259_45724# a_16112_44458# 1.59e-20
C14969 a_8034_45724# a_7640_43914# 1.7e-20
C14970 a_14976_45028# a_14021_43940# 2.27e-20
C14971 C1_N_btm VDD 0.264503f
C14972 a_4883_46098# a_16721_46634# 2.68e-20
C14973 a_18479_47436# a_19123_46287# 8.06e-20
C14974 a_18780_47178# a_18285_46348# 9.29e-19
C14975 a_16327_47482# a_21363_46634# 5.35e-21
C14976 a_2063_45854# a_1823_45246# 0.038948f
C14977 a_584_46384# a_2202_46116# 0.003336f
C14978 a_12549_44172# a_12816_46660# 0.0037f
C14979 a_12891_46348# a_13607_46688# 1.34e-20
C14980 a_10227_46804# a_20107_46660# 0.312495f
C14981 a_3699_46634# a_4651_46660# 3.85e-19
C14982 a_3524_46660# a_4646_46812# 0.001606f
C14983 a_2864_46660# a_3877_44458# 1.05e-19
C14984 a_2107_46812# a_5429_46660# 4.28e-19
C14985 a_n1741_47186# a_6165_46155# 4.48e-20
C14986 a_n2661_46634# a_6969_46634# 0.006553f
C14987 a_n1151_42308# a_472_46348# 1.23e-20
C14988 a_12465_44636# a_13059_46348# 0.163448f
C14989 C6_N_btm C7_N_btm 20.5296f
C14990 C5_N_btm C8_N_btm 0.148944f
C14991 C3_N_btm C10_N_btm 0.208539f
C14992 C4_N_btm C9_N_btm 0.1579f
C14993 C9_P_btm VIN_P 1.82823f
C14994 a_n443_46116# a_n1853_46287# 0.013261f
C14995 a_2124_47436# a_167_45260# 1.26e-19
C14996 a_n237_47217# a_4185_45028# 0.074951f
C14997 a_n743_46660# a_9863_46634# 0.00299f
C14998 a_8685_43396# a_12379_42858# 1.07e-19
C14999 a_2982_43646# a_n2293_42282# 0.010686f
C15000 a_n2661_42282# a_6761_42308# 0.001468f
C15001 a_16823_43084# a_4361_42308# 1.45e-19
C15002 a_18114_32519# a_22459_39145# 1.47e-20
C15003 a_19721_31679# a_22521_40055# 7.56e-21
C15004 a_18579_44172# a_7174_31319# 0.002404f
C15005 a_8560_45348# VDD 0.004463f
C15006 a_21259_43561# a_20556_43646# 9.91e-19
C15007 a_4190_30871# a_743_42282# 0.18536f
C15008 a_9803_43646# a_10083_42826# 0.008857f
C15009 a_9145_43396# a_10518_42984# 6.43e-20
C15010 a_n1557_42282# a_133_42852# 4.96e-19
C15011 a_n2293_46634# a_14635_42282# 2.07e-20
C15012 a_3483_46348# a_9803_43646# 5.4e-19
C15013 a_n1925_42282# a_n2267_43396# 6.35e-19
C15014 a_16751_45260# a_16886_45144# 0.008535f
C15015 a_1307_43914# a_16981_45144# 8.73e-21
C15016 a_4927_45028# a_5518_44484# 0.00158f
C15017 a_n443_42852# a_9672_43914# 8.44e-20
C15018 a_n2017_45002# a_n2012_44484# 0.013231f
C15019 a_n2293_45010# a_n1190_44850# 2.46e-19
C15020 a_12549_44172# a_20753_42852# 8.1e-20
C15021 a_n1613_43370# a_n1329_42308# 0.001867f
C15022 a_5691_45260# a_5343_44458# 4.08e-20
C15023 a_3232_43370# a_4743_44484# 1.9e-19
C15024 a_12741_44636# a_16409_43396# 2.16e-19
C15025 a_15599_45572# a_11967_42832# 1.11e-21
C15026 a_5111_44636# a_6298_44484# 8.64e-20
C15027 a_11361_45348# a_n2661_43370# 0.009376f
C15028 a_n743_46660# a_5527_46155# 1.92e-19
C15029 a_6755_46942# a_5937_45572# 3.17e-19
C15030 a_10249_46116# a_8953_45546# 3.6e-20
C15031 a_4791_45118# a_7499_43078# 0.024468f
C15032 a_15811_47375# a_2711_45572# 1.5e-20
C15033 a_n1925_46634# a_8283_46482# 5.81e-19
C15034 a_19692_46634# a_21542_46660# 4.63e-19
C15035 a_n1151_42308# a_10490_45724# 2.28e-20
C15036 a_10428_46928# a_10355_46116# 0.009109f
C15037 a_n2661_46098# a_739_46482# 4.97e-19
C15038 a_948_46660# a_1337_46116# 1.31e-19
C15039 a_n4318_38680# a_n3674_37592# 0.02489f
C15040 a_3080_42308# a_1239_39587# 3.4e-19
C15041 a_17730_32519# VCM 0.068103f
C15042 a_5342_30871# a_14635_42282# 0.012123f
C15043 a_743_42282# a_5337_42558# 0.001061f
C15044 a_n13_43084# a_n1630_35242# 3.65e-20
C15045 a_13113_42826# a_13622_42852# 2.6e-19
C15046 a_453_43940# VDD 0.225569f
C15047 a_19237_31679# VREF 0.046045f
C15048 a_n443_42852# a_743_42282# 0.03363f
C15049 a_n357_42282# a_20749_43396# 0.001735f
C15050 a_3785_47178# VDD 0.387755f
C15051 a_n863_45724# a_n1991_42858# 3.37e-21
C15052 a_20820_30879# a_n1630_35242# 2.91e-19
C15053 a_2553_47502# DATA[1] 5.06e-21
C15054 a_20193_45348# a_20596_44850# 1.95e-19
C15055 a_n2810_45572# a_n3674_39304# 0.023379f
C15056 a_11827_44484# a_22315_44484# 0.013f
C15057 a_18494_42460# a_20512_43084# 0.115057f
C15058 a_18184_42460# a_22485_44484# 1.09e-21
C15059 a_22223_45036# a_3422_30871# 0.011196f
C15060 a_1307_43914# a_10729_43914# 0.051086f
C15061 a_12607_44458# a_14112_44734# 2.6e-19
C15062 a_13076_44458# a_13468_44734# 0.016359f
C15063 SMPL_ON_N a_22469_40625# 0.03403f
C15064 a_11823_42460# a_15095_43370# 0.003619f
C15065 a_7920_46348# a_8062_46155# 0.005572f
C15066 a_8016_46348# a_10044_46482# 6.14e-19
C15067 a_11901_46660# a_11823_42460# 2.29e-20
C15068 a_12251_46660# a_11962_45724# 1.12e-21
C15069 a_21542_46660# a_20692_30879# 3.76e-20
C15070 a_3090_45724# a_10193_42453# 0.027088f
C15071 a_21588_30879# a_20447_31679# 0.055937f
C15072 a_n2661_46634# a_3357_43084# 0.032385f
C15073 a_12465_44636# a_13556_45296# 0.248126f
C15074 a_4883_46098# a_14180_45002# 7.48e-22
C15075 a_2324_44458# a_526_44458# 0.279023f
C15076 a_5937_45572# a_8049_45260# 0.103218f
C15077 a_13059_46348# a_2711_45572# 0.075233f
C15078 a_n443_46116# a_n2661_43370# 0.030763f
C15079 a_n2293_46634# a_2437_43646# 0.030387f
C15080 a_11453_44696# a_13017_45260# 0.004658f
C15081 a_n881_46662# a_4574_45260# 1.99e-20
C15082 a_13661_43548# a_n2017_45002# 9.71e-20
C15083 a_5807_45002# a_n1059_45260# 5.37e-20
C15084 a_12891_46348# a_413_45260# 5.52e-20
C15085 a_3318_42354# a_5934_30871# 1.28e-20
C15086 a_5342_30871# a_n3420_37984# 0.028488f
C15087 a_564_42282# a_5742_30871# 2.87e-20
C15088 a_n784_42308# a_12563_42308# 3.86e-20
C15089 a_5267_42460# a_6123_31319# 1.13e-20
C15090 a_1606_42308# a_9803_42558# 1.77e-20
C15091 a_5534_30871# a_n4064_37984# 0.047233f
C15092 a_5337_42558# a_5755_42308# 1.15e-19
C15093 a_4921_42308# a_6171_42473# 0.004176f
C15094 a_2382_45260# a_2075_43172# 3.99e-21
C15095 a_n443_42852# a_5755_42308# 4.68e-21
C15096 a_n1331_43914# a_n1453_44318# 3.16e-19
C15097 a_11967_42832# a_18326_43940# 0.058879f
C15098 a_11735_46660# DATA[5] 4.37e-19
C15099 a_375_42282# a_743_42282# 0.006396f
C15100 a_n913_45002# a_10083_42826# 0.052028f
C15101 a_n1059_45260# a_10518_42984# 0.004826f
C15102 a_n2017_45002# a_10835_43094# 1e-19
C15103 a_5891_43370# a_10555_43940# 2.09e-19
C15104 a_4743_44484# a_4905_42826# 2.27e-19
C15105 a_742_44458# a_1987_43646# 2.71e-19
C15106 a_3090_45724# VDD 2.05725f
C15107 a_2889_44172# a_2998_44172# 0.179664f
C15108 a_15009_46634# RST_Z 8.66e-21
C15109 a_n809_44244# a_n3674_39768# 1.06e-21
C15110 a_n1549_44318# a_n1644_44306# 0.049827f
C15111 a_n699_43396# a_766_43646# 0.001138f
C15112 a_n2661_42834# a_2253_43940# 0.004238f
C15113 a_17517_44484# a_11341_43940# 7.52e-20
C15114 a_15433_44458# a_14021_43940# 4.46e-21
C15115 a_n2810_45572# a_5742_30871# 4.02e-21
C15116 a_n357_42282# a_8685_42308# 1.11e-20
C15117 a_n755_45592# a_8325_42308# 0.040306f
C15118 a_10768_47026# CLK 0.005946f
C15119 a_4883_46098# a_20679_44626# 8.04e-21
C15120 a_3218_45724# a_2711_45572# 0.1731f
C15121 a_2957_45546# a_3175_45822# 0.08213f
C15122 a_13259_45724# a_11962_45724# 0.026896f
C15123 a_12891_46348# a_13468_44734# 0.001942f
C15124 a_768_44030# a_n2293_43922# 0.027199f
C15125 a_9625_46129# a_2437_43646# 5.97e-20
C15126 a_n2661_45546# a_2211_45572# 3.69e-19
C15127 a_18985_46122# a_19431_45546# 0.00184f
C15128 a_18819_46122# a_19256_45572# 9.17e-19
C15129 a_472_46348# a_327_44734# 1.53e-19
C15130 a_16327_47482# a_21073_44484# 0.001903f
C15131 a_8199_44636# a_3357_43084# 9.87e-21
C15132 a_4185_45028# a_n2017_45002# 0.029634f
C15133 a_3483_46348# a_n913_45002# 1.56e-20
C15134 a_n443_46116# a_2998_44172# 0.001009f
C15135 a_n2293_46098# a_4558_45348# 0.030863f
C15136 a_6755_46942# a_11691_44458# 0.192426f
C15137 a_4646_46812# a_5343_44458# 0.24395f
C15138 a_10586_45546# a_10210_45822# 0.042978f
C15139 a_n443_42852# a_2277_45546# 1.61e-20
C15140 a_1239_47204# a_n1435_47204# 2.24e-19
C15141 a_n443_46116# a_4915_47217# 0.395101f
C15142 a_4791_45118# a_5129_47502# 0.240381f
C15143 a_2063_45854# a_11031_47542# 9.91e-19
C15144 a_n1151_42308# a_7227_47204# 1.79e-19
C15145 a_n4064_40160# a_n3690_38528# 2.54e-19
C15146 a_1606_42308# C7_P_btm 0.00238f
C15147 a_n2472_42282# VDD 0.278905f
C15148 a_n784_42308# C1_N_btm 0.027772f
C15149 a_19279_43940# a_4361_42308# 4.21e-21
C15150 a_18579_44172# a_21487_43396# 2.15e-21
C15151 a_9313_44734# a_10991_42826# 0.007504f
C15152 a_n2661_43370# a_n4318_37592# 2.73e-20
C15153 a_15002_46116# VDD 4.6e-19
C15154 a_742_44458# a_4649_42852# 5.01e-21
C15155 a_n2293_42834# a_564_42282# 5.42e-20
C15156 a_n2661_42834# a_7871_42858# 1.63e-20
C15157 a_n2293_43922# a_5755_42852# 3.26e-21
C15158 a_20692_30879# C2_N_btm 1.93e-20
C15159 a_n2661_42282# a_7274_43762# 9.24e-21
C15160 a_1307_43914# a_5932_42308# 0.00164f
C15161 a_n443_42852# a_626_44172# 0.028669f
C15162 a_2711_45572# a_13556_45296# 0.00137f
C15163 a_8049_45260# a_11691_44458# 7.14e-20
C15164 a_3147_46376# a_3363_44484# 4e-21
C15165 w_11334_34010# a_4190_30871# 0.006418f
C15166 a_7227_45028# a_8191_45002# 8.51e-20
C15167 a_13259_45724# a_13807_45067# 1.17e-19
C15168 a_1823_45246# a_n2661_42834# 0.174801f
C15169 a_12741_44636# a_16241_44734# 0.006663f
C15170 a_3090_45724# a_5495_43940# 0.004468f
C15171 a_8696_44636# a_17034_45572# 4.18e-19
C15172 a_1138_42852# a_n2661_43922# 0.027736f
C15173 a_5437_45600# a_5111_44636# 3.47e-19
C15174 a_8016_46348# a_7640_43914# 2.21e-22
C15175 a_768_44030# a_n97_42460# 0.034422f
C15176 a_17715_44484# a_14539_43914# 6.56e-19
C15177 a_13747_46662# a_17538_32519# 1.11e-19
C15178 a_n2293_46634# a_11257_43940# 1.65e-19
C15179 a_n2472_46634# a_n2442_46660# 0.155358f
C15180 a_n2661_46634# a_n2293_46634# 0.060962f
C15181 a_n1151_42308# a_12156_46660# 0.003059f
C15182 a_n1613_43370# a_3686_47026# 2.49e-19
C15183 a_3754_38470# VDD 2.52245f
C15184 a_4883_46098# a_7927_46660# 5.28e-21
C15185 VDAC_P C8_P_btm 61.723297f
C15186 a_11459_47204# a_11813_46116# 1.67e-20
C15187 a_22609_38406# a_22717_37285# 0.08753f
C15188 a_22705_38406# a_22705_37990# 0.003483f
C15189 CAL_P a_22717_36887# 9.62e-21
C15190 a_n2840_46634# a_n2312_38680# 0.040373f
C15191 a_1414_42308# a_n327_42558# 2.72e-21
C15192 a_10341_43396# a_16759_43396# 0.010617f
C15193 a_n97_42460# a_5755_42852# 0.149651f
C15194 a_413_45260# SINGLE_ENDED 0.037852f
C15195 a_n356_44636# a_18997_42308# 1.66e-20
C15196 a_2274_45254# VDD 0.256655f
C15197 a_14579_43548# a_15743_43084# 1.21e-19
C15198 a_458_43396# a_791_42968# 3.18e-19
C15199 a_9313_44734# a_17303_42282# 9.64e-19
C15200 a_584_46384# a_961_42354# 9.03e-21
C15201 a_9290_44172# a_10555_43940# 4.56e-19
C15202 a_7276_45260# a_7418_45394# 0.007833f
C15203 a_11962_45724# a_n2661_43922# 2.11e-20
C15204 a_n863_45724# a_n1331_43914# 1.23e-20
C15205 a_1307_43914# a_1423_45028# 0.054616f
C15206 a_375_42282# a_626_44172# 0.017957f
C15207 a_7499_43078# a_10809_44484# 3.94e-19
C15208 a_3537_45260# a_n2661_43370# 0.087747f
C15209 a_n2293_46634# a_14543_43071# 9.13e-20
C15210 a_n1151_42308# a_n3674_37592# 0.007818f
C15211 a_3090_45724# a_16137_43396# 1.3e-20
C15212 a_13661_43548# a_19164_43230# 3.49e-19
C15213 a_22223_45572# a_20193_45348# 1.1e-19
C15214 a_n2293_45546# a_n809_44244# 5.56e-20
C15215 a_n1079_45724# a_n1549_44318# 1.64e-19
C15216 a_6171_45002# a_8137_45348# 1.04e-19
C15217 a_15861_45028# a_14539_43914# 2.35e-19
C15218 a_8696_44636# a_16979_44734# 0.005402f
C15219 a_5807_45002# a_13925_46122# 0.027158f
C15220 a_13661_43548# a_13759_46122# 8.09e-22
C15221 a_n743_46660# a_6165_46155# 0.004708f
C15222 a_n2661_46098# a_1176_45822# 0.144277f
C15223 a_6969_46634# a_765_45546# 0.001746f
C15224 a_n881_46662# a_10809_44734# 0.026121f
C15225 a_17609_46634# a_18834_46812# 0.001296f
C15226 a_n237_47217# a_997_45618# 1.85e-19
C15227 a_n1925_46634# a_7920_46348# 0.007001f
C15228 a_2905_45572# a_n2661_45546# 0.003174f
C15229 a_12469_46902# a_12347_46660# 3.16e-19
C15230 a_18479_47436# a_8049_45260# 0.047429f
C15231 a_11599_46634# a_12379_46436# 0.005949f
C15232 a_n971_45724# a_2957_45546# 8.45e-20
C15233 a_327_47204# a_310_45028# 1.58e-19
C15234 a_2107_46812# a_3483_46348# 0.100707f
C15235 a_n2661_46634# a_9625_46129# 3.03e-19
C15236 a_n2293_46634# a_8199_44636# 0.029753f
C15237 a_2063_45854# a_n2293_45546# 0.002045f
C15238 a_4883_46098# a_6419_46482# 7.98e-20
C15239 a_n2312_39304# a_n1925_42282# 6.33e-20
C15240 a_19237_31679# a_22521_40599# 1.41e-20
C15241 a_20974_43370# a_17303_42282# 5.91e-22
C15242 a_n97_42460# a_10149_42308# 8.69e-19
C15243 a_6547_43396# a_6123_31319# 1.98e-19
C15244 a_7287_43370# a_7227_42308# 1.42e-19
C15245 a_7112_43396# a_6761_42308# 1.62e-20
C15246 a_5534_30871# a_15279_43071# 0.00177f
C15247 a_743_42282# a_14635_42282# 0.02914f
C15248 a_14815_43914# VDD 0.307386f
C15249 a_1847_42826# a_1793_42852# 2.52e-20
C15250 a_15743_43084# a_20573_43172# 3.04e-20
C15251 a_14543_43071# a_5342_30871# 5.56e-19
C15252 a_n443_42852# a_2813_43396# 0.017355f
C15253 a_3232_43370# a_1414_42308# 0.248035f
C15254 a_1823_45246# a_n2293_42282# 0.03994f
C15255 a_9290_44172# a_13113_42826# 0.003778f
C15256 a_4185_45028# a_19164_43230# 6.39e-21
C15257 a_13259_45724# a_17499_43370# 0.018042f
C15258 a_3065_45002# a_3905_42865# 0.034773f
C15259 a_3537_45260# a_2998_44172# 0.059736f
C15260 a_8016_46348# a_9823_46155# 0.048283f
C15261 a_n2840_46090# a_n2956_38680# 0.050916f
C15262 a_2521_46116# a_2324_44458# 1.5e-20
C15263 a_n2472_46090# a_n2956_39304# 9.6e-19
C15264 a_n1151_42308# a_6171_45002# 0.02292f
C15265 a_n443_46116# a_4574_45260# 5.16e-20
C15266 a_7903_47542# a_413_45260# 1.03e-19
C15267 a_18143_47464# a_3357_43084# 5.7e-19
C15268 a_n2497_47436# a_1307_43914# 0.069365f
C15269 a_6755_46942# a_n443_42852# 1.03e-19
C15270 a_5807_45002# a_15599_45572# 0.002399f
C15271 a_8199_44636# a_9625_46129# 0.011574f
C15272 a_5937_45572# a_8953_45546# 0.3871f
C15273 a_13747_46662# a_15225_45822# 6.29e-19
C15274 a_2063_45854# a_6709_45028# 4.65e-20
C15275 a_16327_47482# a_21542_45572# 0.002879f
C15276 a_5257_43370# a_5263_45724# 0.088982f
C15277 a_7577_46660# a_2711_45572# 4.24e-20
C15278 a_n971_45724# a_9482_43914# 8.96e-21
C15279 a_4791_45118# a_4558_45348# 0.077256f
C15280 a_18597_46090# a_2437_43646# 0.006962f
C15281 a_18479_47436# a_19479_31679# 2.29e-20
C15282 a_n1821_43396# VDD 3.05e-20
C15283 a_4190_30871# a_n4064_37984# 0.032018f
C15284 a_18599_43230# a_17303_42282# 1.61e-20
C15285 a_5534_30871# a_13258_32519# 0.04166f
C15286 a_n2840_42282# a_n3674_37592# 0.007977f
C15287 a_n4318_37592# COMP_P 0.001501f
C15288 a_17538_32519# VCM 0.0424f
C15289 a_18249_42858# a_18057_42282# 1.52e-19
C15290 a_18083_42858# a_18907_42674# 1.44e-20
C15291 a_n1736_42282# a_n1329_42308# 0.050456f
C15292 a_n3674_39304# a_n4251_39392# 8.42e-19
C15293 a_n3674_38216# a_n961_42308# 7.46e-20
C15294 a_3080_42308# C1_N_btm 0.011373f
C15295 a_13720_44458# a_11341_43940# 2.52e-20
C15296 a_5111_44636# a_9885_43396# 0.004113f
C15297 a_n2661_46098# DATA[0] 4.59e-20
C15298 a_1799_45572# DATA[1] 0.004719f
C15299 a_11691_44458# a_15037_43940# 2.9e-20
C15300 a_1423_45028# a_9396_43370# 5.93e-21
C15301 a_18287_44626# a_15493_43396# 1.74e-20
C15302 a_18374_44850# a_18451_43940# 6.12e-19
C15303 a_n2661_43922# a_n4318_39768# 0.010131f
C15304 a_5891_43370# a_n2661_42282# 0.032052f
C15305 a_n2661_42834# a_n3674_39768# 0.150968f
C15306 a_18989_43940# a_18326_43940# 3.26e-20
C15307 a_11967_42832# a_22959_44484# 4.39e-22
C15308 a_20640_44752# a_20512_43084# 4.38e-19
C15309 a_20766_44850# a_20637_44484# 4.2e-19
C15310 a_20835_44721# a_21073_44484# 0.001705f
C15311 a_19279_43940# a_20397_44484# 0.002084f
C15312 a_20679_44626# a_21145_44484# 3.82e-19
C15313 a_n1059_45260# a_16867_43762# 1.11e-19
C15314 a_8975_43940# a_9248_44260# 0.001408f
C15315 a_3699_46634# VDD 0.347281f
C15316 a_11827_44484# a_19319_43548# 0.00137f
C15317 a_7640_43914# a_7584_44260# 5.72e-19
C15318 a_526_44458# a_9803_42558# 2.85e-19
C15319 a_n2293_42834# a_n1557_42282# 0.034384f
C15320 a_18184_42460# a_14401_32519# 4.69e-20
C15321 a_18494_42460# a_21381_43940# 2.36e-20
C15322 a_10768_47026# a_10951_45334# 8.49e-21
C15323 a_8199_44636# a_9159_45572# 0.049711f
C15324 a_5732_46660# a_5837_45028# 3.47e-21
C15325 a_6945_45028# a_7499_43078# 4.09e-22
C15326 a_5257_43370# a_5837_45348# 0.001158f
C15327 a_768_44030# a_742_44458# 0.216263f
C15328 a_3090_45724# a_5691_45260# 1.29e-22
C15329 a_2324_44458# a_13163_45724# 7.36e-21
C15330 a_14275_46494# a_13249_42308# 8.84e-19
C15331 a_14493_46090# a_14495_45572# 0.00228f
C15332 a_9290_44172# a_10907_45822# 0.262972f
C15333 a_11189_46129# a_10210_45822# 3.66e-19
C15334 a_19321_45002# a_20205_45028# 5.38e-19
C15335 a_13747_46662# a_19721_31679# 0.001393f
C15336 a_n881_46662# a_5883_43914# 2.63e-20
C15337 a_765_45546# a_3357_43084# 0.035297f
C15338 a_19123_46287# a_2437_43646# 7.12e-20
C15339 a_11415_45002# a_18596_45572# 9.68e-19
C15340 a_19647_42308# a_13258_32519# 0.153411f
C15341 a_19511_42282# a_20107_42308# 0.043647f
C15342 a_17303_42282# a_22397_42558# 0.012536f
C15343 a_n4318_37592# a_n3565_37414# 4.06e-19
C15344 a_17517_44484# a_10341_43396# 0.001868f
C15345 a_n1441_43940# a_n2433_43396# 2.36e-19
C15346 a_10405_44172# a_11173_43940# 7.97e-21
C15347 a_10729_43914# a_10867_43940# 0.00501f
C15348 a_10807_43548# a_10555_43940# 1.21e-19
C15349 a_1115_44172# a_n1557_42282# 3.9e-19
C15350 a_4223_44672# a_3935_42891# 8.13e-21
C15351 a_n2017_45002# a_n39_42308# 6.45e-19
C15352 a_n913_45002# a_2351_42308# 0.023646f
C15353 a_20075_46420# VDD 0.347847f
C15354 a_19553_46090# START 1.2e-21
C15355 a_19335_46494# RST_Z 1.49e-21
C15356 a_15015_46420# CLK 7.59e-21
C15357 a_n2661_44458# a_10083_42826# 9.84e-22
C15358 a_3357_43084# a_4921_42308# 2.67e-20
C15359 a_18494_42460# a_18249_42858# 8.63e-19
C15360 a_18184_42460# a_18817_42826# 6.72e-20
C15361 a_11691_44458# a_15279_43071# 1.05e-19
C15362 a_2479_44172# a_4235_43370# 1.29e-20
C15363 a_14495_45572# a_15903_45785# 3.7e-21
C15364 a_11823_42460# a_8696_44636# 0.026654f
C15365 a_n443_46116# a_1568_43370# 0.584982f
C15366 a_584_46384# a_2982_43646# 0.057754f
C15367 a_n971_45724# a_6031_43396# 4.44e-21
C15368 a_3483_46348# a_n2661_44458# 1.44355f
C15369 a_1208_46090# a_949_44458# 2.47e-20
C15370 a_11415_45002# a_15004_44636# 6.08e-19
C15371 a_10490_45724# a_12649_45572# 4.67e-19
C15372 a_12549_44172# a_11341_43940# 0.406618f
C15373 a_n755_45592# a_n1059_45260# 0.53237f
C15374 a_n2661_45546# a_n37_45144# 0.001732f
C15375 a_n357_42282# a_n913_45002# 0.309845f
C15376 a_2277_45546# a_2437_43646# 0.001212f
C15377 a_8034_45724# a_1423_45028# 2.81e-21
C15378 a_15143_45578# a_15599_45572# 2.96e-19
C15379 a_10907_45822# a_11064_45572# 0.007306f
C15380 a_12741_44636# a_12883_44458# 0.073263f
C15381 a_n863_45724# a_n967_45348# 4.28e-20
C15382 a_n2293_45546# a_n955_45028# 0.002208f
C15383 a_13661_43548# a_18079_43940# 0.028277f
C15384 a_526_44458# a_2448_45028# 7.21e-21
C15385 a_n4334_37440# a_n3565_37414# 0.001292f
C15386 a_n4209_37414# a_n3690_37440# 0.046103f
C15387 a_21177_47436# a_20916_46384# 4.75e-19
C15388 a_20990_47178# a_21588_30879# 2.92e-19
C15389 a_16023_47582# a_n743_46660# 0.004115f
C15390 a_n971_45724# a_7715_46873# 0.029319f
C15391 a_n4315_30879# VREF 1.73216f
C15392 a_3785_47178# a_4646_46812# 8.96e-19
C15393 a_3815_47204# a_3877_44458# 1.11e-19
C15394 a_n2216_39866# VDD 0.004696f
C15395 a_n4209_38502# C7_P_btm 7.54e-20
C15396 a_n3565_38502# C9_P_btm 1.91e-20
C15397 a_n4064_40160# VIN_P 0.06337f
C15398 a_n4209_38216# a_n1386_35608# 1.32e-19
C15399 a_n237_47217# a_5257_43370# 0.022234f
C15400 a_2063_45854# a_5732_46660# 2.69e-20
C15401 a_n1151_42308# a_4955_46873# 0.261025f
C15402 a_4883_46098# a_19594_46812# 3.17e-19
C15403 a_3626_43646# a_14358_43442# 1.37e-20
C15404 a_2982_43646# a_15095_43370# 4.05e-20
C15405 a_n2661_42834# a_1184_42692# 6.05e-21
C15406 a_n356_44636# a_6123_31319# 0.169259f
C15407 a_3905_42865# a_2987_42968# 4.66e-20
C15408 en_comp VDAC_N 7.58e-19
C15409 a_n97_42460# a_16759_43396# 0.003171f
C15410 a_n913_45002# CAL_N 0.002966f
C15411 a_n2293_43922# a_1067_42314# 3.58e-20
C15412 a_7112_43396# a_7274_43762# 0.006453f
C15413 a_6547_43396# a_6809_43396# 0.001705f
C15414 a_12429_44172# a_12089_42308# 1.7e-21
C15415 a_13483_43940# a_12379_42858# 5.33e-20
C15416 a_20447_31679# a_22469_39537# 5.38e-20
C15417 a_6197_43396# a_7221_43396# 2.36e-20
C15418 a_8162_45546# a_5883_43914# 1.03e-21
C15419 a_n2293_45546# a_n2661_42834# 4.84e-20
C15420 a_n2956_38216# a_n2661_43922# 2.48e-19
C15421 a_3537_45260# a_4574_45260# 0.234297f
C15422 a_3065_45002# a_5147_45002# 4.34e-21
C15423 a_5937_45572# a_9028_43914# 2.88e-19
C15424 a_8199_44636# a_9672_43914# 0.043804f
C15425 a_8016_46348# a_10729_43914# 0.006537f
C15426 a_12861_44030# a_21356_42826# 1.38e-20
C15427 a_7499_43078# a_8103_44636# 3.16e-19
C15428 a_9049_44484# a_6298_44484# 2.08e-21
C15429 a_16375_45002# a_16241_44734# 1.69e-19
C15430 a_3090_45724# a_3080_42308# 0.002565f
C15431 a_10227_46804# a_15567_42826# 0.008041f
C15432 a_13259_45724# a_18204_44850# 1.43e-19
C15433 a_2437_43646# a_626_44172# 2.83e-21
C15434 a_4791_45118# a_5193_43172# 8.86e-20
C15435 a_21588_30879# a_13467_32519# 0.057457f
C15436 a_16327_47482# a_18083_42858# 0.591108f
C15437 a_n881_46662# a_n2157_46122# 0.005335f
C15438 a_11453_44696# a_3483_46348# 0.027804f
C15439 a_n1151_42308# a_n967_46494# 4.11e-19
C15440 a_13717_47436# a_15015_46420# 4.43e-21
C15441 a_12861_44030# a_14275_46494# 1.23e-19
C15442 a_20916_46384# a_20841_46902# 2.67e-19
C15443 a_768_44030# a_11415_45002# 0.021062f
C15444 a_5807_45002# a_16655_46660# 0.006956f
C15445 a_4883_46098# a_5164_46348# 0.01685f
C15446 a_14955_47212# a_13759_46122# 2.05e-20
C15447 a_7577_46660# a_8654_47026# 1.46e-19
C15448 a_4646_46812# a_3090_45724# 0.199722f
C15449 a_n2293_46634# a_765_45546# 8.06e-22
C15450 a_n1613_43370# a_n1853_46287# 0.354256f
C15451 a_10554_47026# a_6755_46942# 0.005096f
C15452 a_n237_47217# a_1337_46116# 8.45e-19
C15453 a_10227_46804# a_9569_46155# 1.63e-20
C15454 a_14311_47204# a_13925_46122# 1.89e-21
C15455 a_11599_46634# a_13351_46090# 0.105205f
C15456 a_15493_43396# a_17124_42282# 2.88e-21
C15457 a_5649_42852# a_10341_42308# 1.31e-20
C15458 a_104_43370# a_n1630_35242# 5.25e-21
C15459 a_16823_43084# a_17595_43084# 8.04e-20
C15460 a_4361_42308# a_12545_42858# 1.78e-19
C15461 a_19721_31679# VCM 0.03544f
C15462 a_n3674_39768# a_n3565_39590# 0.128683f
C15463 a_n4318_39768# a_n3690_39616# 3.79e-19
C15464 a_4743_44484# VDD 0.266843f
C15465 a_17737_43940# a_17303_42282# 7.23e-21
C15466 a_743_42282# a_14543_43071# 2.19e-20
C15467 a_15743_43084# a_21671_42860# 0.004756f
C15468 a_18597_46090# a_19511_42282# 0.156698f
C15469 a_n2661_43370# a_8701_44490# 2.05e-19
C15470 a_9482_43914# a_9313_44734# 0.060868f
C15471 a_n2017_45002# a_11967_42832# 0.086561f
C15472 a_18479_47436# a_13258_32519# 1.35e-21
C15473 a_n2293_46634# a_4921_42308# 4.37e-20
C15474 a_11525_45546# a_11341_43940# 2.62e-20
C15475 a_7499_43078# a_11173_44260# 5.58e-19
C15476 a_1307_43914# a_6109_44484# 0.00821f
C15477 a_7229_43940# a_n2661_43922# 0.030151f
C15478 a_19778_44110# a_18114_32519# 5.95e-20
C15479 a_11691_44458# a_20193_45348# 0.003224f
C15480 a_18184_42460# a_20205_45028# 0.001438f
C15481 a_10907_45822# a_10807_43548# 0.002089f
C15482 a_4185_45028# a_14209_32519# 0.091175f
C15483 a_8199_44636# a_743_42282# 0.036554f
C15484 a_17715_44484# a_17324_43396# 0.002059f
C15485 a_18189_46348# a_17499_43370# 2.45e-20
C15486 a_13507_46334# a_18907_42674# 0.202065f
C15487 a_948_46660# a_n755_45592# 8.59e-22
C15488 a_n743_46660# a_n23_45546# 0.070296f
C15489 a_1123_46634# a_997_45618# 1.11e-20
C15490 a_n2438_43548# a_n356_45724# 5.71e-20
C15491 a_14513_46634# a_14493_46090# 0.00967f
C15492 a_14180_46812# a_14275_46494# 0.002474f
C15493 a_15227_44166# a_6945_45028# 0.548194f
C15494 a_17609_46634# a_10809_44734# 0.018125f
C15495 a_14035_46660# a_15015_46420# 1.29e-20
C15496 a_765_45546# a_9625_46129# 1.15e-19
C15497 a_9313_45822# a_8696_44636# 4.84e-20
C15498 a_2443_46660# a_n2661_45546# 1.59e-20
C15499 a_12861_44030# a_15765_45572# 0.026773f
C15500 a_19692_46634# a_19900_46494# 0.004501f
C15501 a_13059_46348# a_12005_46116# 3.28e-19
C15502 a_n2293_46098# a_n1853_46287# 0.02738f
C15503 a_n2472_46090# a_n1991_46122# 7.66e-19
C15504 a_n881_46662# a_8162_45546# 1.32e-20
C15505 a_n2661_46634# a_2277_45546# 8.59e-21
C15506 a_11453_44696# a_14495_45572# 7.3e-20
C15507 a_3080_42308# a_3754_38470# 3.23e-19
C15508 a_5649_42852# a_18057_42282# 6.29e-20
C15509 a_4190_30871# a_13258_32519# 0.039476f
C15510 a_n2293_42282# a_1184_42692# 1.61e-19
C15511 a_4361_42308# a_19332_42282# 0.009695f
C15512 a_13887_32519# a_17303_42282# 0.0067f
C15513 a_945_42968# a_n784_42308# 7.59e-20
C15514 a_743_42282# a_19511_42282# 0.00872f
C15515 a_8952_43230# a_8685_42308# 0.008199f
C15516 a_22959_43948# RST_Z 0.001362f
C15517 a_5518_44484# a_5244_44056# 2.08e-19
C15518 a_4223_44672# a_6453_43914# 0.019918f
C15519 a_11827_44484# a_10949_43914# 5.25e-20
C15520 a_2583_47243# VDD 2.18e-20
C15521 a_n2956_38680# a_n2104_42282# 2.5e-20
C15522 a_3065_45002# a_4093_43548# 0.003025f
C15523 a_2382_45260# a_4699_43561# 6.05e-21
C15524 a_n2433_44484# a_n1441_43940# 4.71e-20
C15525 a_n310_47243# DATA[0] 0.002781f
C15526 a_2747_46873# DATA[1] 3.15e-21
C15527 a_3357_43084# a_6452_43396# 5.12e-19
C15528 a_n443_42852# a_15279_43071# 8.83e-21
C15529 a_n357_42282# a_20922_43172# 0.059485f
C15530 a_13857_44734# a_14673_44172# 2.8e-20
C15531 a_5343_44458# a_5013_44260# 1.37e-19
C15532 a_9313_44734# a_20159_44458# 1.77e-20
C15533 en_comp a_3626_43646# 5.78e-20
C15534 a_n2956_39304# a_n3674_38216# 0.023505f
C15535 a_15861_45028# a_17324_43396# 1.36e-19
C15536 a_2437_43646# a_2813_43396# 0.012852f
C15537 a_11453_44696# a_17719_45144# 0.105851f
C15538 a_18479_47436# a_20193_45348# 0.021013f
C15539 a_5066_45546# a_9751_46155# 6.54e-21
C15540 a_20708_46348# a_20205_31679# 2.2e-19
C15541 a_6945_45028# a_21071_46482# 7.43e-19
C15542 a_1823_45246# a_3775_45552# 0.070347f
C15543 a_4704_46090# a_2711_45572# 1.41e-19
C15544 a_11415_45002# a_11652_45724# 0.128811f
C15545 a_n1613_43370# a_n2661_43370# 0.05744f
C15546 a_5807_45002# a_5837_45348# 0.003033f
C15547 a_8953_45546# a_n443_42852# 0.134632f
C15548 a_3877_44458# a_2382_45260# 0.395451f
C15549 a_4817_46660# a_413_45260# 1.37e-20
C15550 a_5257_43370# a_n2017_45002# 2.04e-19
C15551 a_3090_45724# a_18479_45785# 0.259218f
C15552 a_6755_46942# a_2437_43646# 2.3e-19
C15553 a_4791_45118# a_9838_44484# 1.34e-19
C15554 a_4185_45028# a_4099_45572# 0.025863f
C15555 a_3483_46348# a_5907_45546# 6.03e-20
C15556 a_n743_46660# a_14797_45144# 2.35e-21
C15557 a_4883_46098# a_18494_42460# 4.26e-20
C15558 a_14456_42282# a_14113_42308# 0.038993f
C15559 a_n3674_38680# a_n4064_39072# 0.020036f
C15560 a_n1736_43218# VDD 0.082445f
C15561 a_14209_32519# VREF_GND 0.034351f
C15562 a_n4318_38216# a_n3420_39072# 0.032825f
C15563 COMP_P a_1343_38525# 0.004705f
C15564 a_n1630_35242# a_n2946_39866# 6.3e-21
C15565 a_17364_32525# VIN_N 0.039314f
C15566 a_8375_44464# a_8147_43396# 3.2e-20
C15567 a_5891_43370# a_7112_43396# 5.95e-19
C15568 a_n2293_42834# a_3935_42891# 0.008823f
C15569 a_17517_44484# a_n97_42460# 7.31e-22
C15570 a_22959_46660# RST_Z 0.001115f
C15571 a_18494_42460# a_5649_42852# 1.97e-19
C15572 a_14539_43914# a_15095_43370# 4.59e-20
C15573 a_2711_45572# a_17303_42282# 3.67e-19
C15574 a_21076_30879# VDD 1.17389f
C15575 a_18579_44172# a_18797_44260# 4.08e-20
C15576 a_10193_42453# a_11633_42558# 0.017236f
C15577 a_3537_45260# a_4743_43172# 0.002397f
C15578 a_1307_43914# a_15567_42826# 2.68e-20
C15579 a_20193_45348# a_4190_30871# 0.02125f
C15580 a_8333_44056# a_9028_43914# 0.007993f
C15581 a_13351_46090# a_13348_45260# 1.28e-19
C15582 a_12594_46348# a_9482_43914# 5.94e-21
C15583 a_3090_45724# a_10057_43914# 0.230475f
C15584 a_18051_46116# a_18175_45572# 2.57e-19
C15585 a_n1925_42282# a_n2810_45028# 2.5e-20
C15586 a_8049_45260# a_2437_43646# 0.041161f
C15587 a_10227_46804# a_10405_44172# 0.011223f
C15588 a_10903_43370# a_13777_45326# 3.61e-19
C15589 a_2711_45572# a_6905_45572# 6.06e-19
C15590 a_8016_46348# a_1423_45028# 1.1e-20
C15591 a_2324_44458# a_8953_45002# 1.65784f
C15592 a_n2293_46098# a_n2661_43370# 0.027372f
C15593 a_11415_45002# a_13490_45067# 0.002913f
C15594 a_19123_46287# a_19113_45348# 1.62e-19
C15595 a_19321_45002# a_20512_43084# 1.07e-19
C15596 a_768_44030# a_n984_44318# 3.28e-20
C15597 a_20273_46660# a_21359_45002# 7.05e-22
C15598 a_12861_44030# a_19328_44172# 1.89e-19
C15599 a_n4209_39304# a_n4334_37440# 4.61e-19
C15600 a_11633_42558# VDD 0.193501f
C15601 a_1736_39043# a_3754_38802# 7.66e-20
C15602 a_10227_46804# a_19386_47436# 0.041193f
C15603 a_18479_47436# a_18780_47178# 0.056304f
C15604 a_18143_47464# a_18597_46090# 0.002913f
C15605 a_n3420_37984# a_n4064_37984# 8.18485f
C15606 a_n1435_47204# a_n2312_39304# 6.02e-19
C15607 a_4915_47217# a_n1613_43370# 0.195064f
C15608 a_16327_47482# a_13507_46334# 0.043159f
C15609 a_n443_46116# a_n881_46662# 0.114922f
C15610 a_15507_47210# a_12465_44636# 9.53e-19
C15611 a_4700_47436# a_4842_47243# 0.005572f
C15612 a_2553_47502# a_768_44030# 2.24e-19
C15613 a_n237_47217# a_5807_45002# 0.082779f
C15614 a_n2833_47464# a_n2956_39768# 0.008074f
C15615 a_15493_43940# a_16547_43609# 0.002713f
C15616 a_11341_43940# a_16977_43638# 6.41e-21
C15617 a_19328_44172# a_19700_43370# 1.6e-19
C15618 a_n2956_37592# a_n4209_38502# 0.090878f
C15619 en_comp a_2112_39137# 1.51e-20
C15620 a_15493_43396# a_19268_43646# 0.024436f
C15621 a_2127_44172# a_1847_42826# 8.79e-22
C15622 a_1414_42308# a_2905_42968# 0.00136f
C15623 a_19615_44636# a_19339_43156# 1.43e-21
C15624 a_11967_42832# a_19164_43230# 1.58e-20
C15625 a_9313_44734# a_11301_43218# 2.3e-19
C15626 a_n2129_43609# a_n1243_43396# 9.68e-19
C15627 a_n97_42460# a_1891_43646# 0.001075f
C15628 a_1049_43396# a_1568_43370# 2.09e-20
C15629 a_19478_44306# a_15743_43084# 7.05e-21
C15630 a_15037_45618# a_9482_43914# 2.11e-19
C15631 a_n1079_45724# a_n1177_44458# 6.5e-20
C15632 a_n2293_45546# a_n1352_44484# 1.39e-19
C15633 a_2711_45572# a_19778_44110# 0.003443f
C15634 a_n2293_46634# a_6452_43396# 0.00445f
C15635 a_12549_44172# a_10341_43396# 0.0385f
C15636 a_n357_42282# a_n2661_44458# 0.031616f
C15637 a_17957_46116# a_17517_44484# 2.11e-21
C15638 a_18189_46348# a_18204_44850# 2.34e-20
C15639 a_4185_45028# a_17730_32519# 0.097949f
C15640 a_13059_46348# a_15682_43940# 9.48e-20
C15641 a_2437_43646# a_19479_31679# 0.004873f
C15642 a_21513_45002# a_3357_43084# 0.04265f
C15643 a_18597_46090# a_21259_43561# 0.005266f
C15644 a_n2293_46098# a_2998_44172# 2.44e-19
C15645 a_n2661_45546# a_949_44458# 1.19e-19
C15646 a_13259_45724# a_15004_44636# 6.12e-19
C15647 a_3090_45724# a_14021_43940# 0.049176f
C15648 C0_N_btm VDD 1.02806f
C15649 a_4883_46098# a_16388_46812# 0.041939f
C15650 a_18597_46090# a_765_45546# 1.63e-19
C15651 a_18479_47436# a_18285_46348# 7.49e-21
C15652 a_5807_45002# a_8270_45546# 0.029164f
C15653 a_584_46384# a_1823_45246# 0.094654f
C15654 a_2124_47436# a_2202_46116# 4.23e-20
C15655 a_12891_46348# a_12816_46660# 0.024711f
C15656 a_12549_44172# a_12991_46634# 0.010497f
C15657 a_n443_46116# a_n2157_46122# 3.46e-20
C15658 a_21589_35634# VIN_N 0.029423f
C15659 C10_P_btm VIN_P 3.66034f
C15660 a_3699_46634# a_4646_46812# 2.69e-19
C15661 a_3524_46660# a_3877_44458# 0.008528f
C15662 a_2107_46812# a_5263_46660# 8.47e-19
C15663 a_n2661_46634# a_6755_46942# 1.40968f
C15664 a_2063_45854# a_1138_42852# 2.69e-19
C15665 a_12861_44030# a_18280_46660# 0.140921f
C15666 C5_N_btm C7_N_btm 0.15419f
C15667 C2_N_btm C10_N_btm 0.215144f
C15668 C3_N_btm C9_N_btm 0.138859f
C15669 C4_N_btm C8_N_btm 0.149948f
C15670 a_1431_47204# a_167_45260# 5.7e-22
C15671 a_n237_47217# a_3699_46348# 0.044064f
C15672 a_n971_45724# a_4419_46090# 2.52e-19
C15673 a_n743_46660# a_8492_46660# 1.3e-20
C15674 a_2609_46660# a_4817_46660# 0.00171f
C15675 a_8685_43396# a_10341_42308# 3.51e-19
C15676 a_21259_43561# a_743_42282# 2.87e-19
C15677 a_4190_30871# a_20301_43646# 0.00107f
C15678 a_9145_43396# a_10083_42826# 6.91e-20
C15679 a_3483_46348# a_9145_43396# 2.59e-19
C15680 a_n1925_42282# a_n2129_43609# 5.05e-20
C15681 a_1307_43914# a_16886_45144# 9.14e-21
C15682 a_5111_44636# a_5518_44484# 0.124556f
C15683 a_4927_45028# a_5343_44458# 1.54e-19
C15684 a_n357_42282# a_18451_43940# 4.34e-22
C15685 a_n2017_45002# a_18989_43940# 1.19e-20
C15686 a_12549_44172# a_20356_42852# 9.25e-21
C15687 a_n1613_43370# COMP_P 0.001404f
C15688 a_3232_43370# a_n699_43396# 0.074855f
C15689 a_3537_45260# a_5883_43914# 0.018824f
C15690 a_6171_45002# a_4223_44672# 1.27e-20
C15691 a_8704_45028# a_n2661_43370# 3.79e-19
C15692 a_12741_44636# a_16547_43609# 3.38e-20
C15693 w_1575_34946# a_n3420_38528# 5.84e-19
C15694 a_n743_46660# a_5210_46155# 1.05e-19
C15695 a_5807_45002# a_12638_46436# 0.006618f
C15696 a_768_44030# a_13259_45724# 0.315247f
C15697 a_6755_46942# a_8199_44636# 3.74e-19
C15698 a_4791_45118# a_8568_45546# 2.1e-20
C15699 a_19692_46634# a_21297_46660# 5.35e-19
C15700 a_15507_47210# a_2711_45572# 5.18e-21
C15701 a_n1151_42308# a_8746_45002# 6.07e-20
C15702 a_2063_45854# a_11962_45724# 0.011034f
C15703 a_10150_46912# a_10355_46116# 7.72e-19
C15704 a_n2661_46634# a_8049_45260# 0.027919f
C15705 a_n2661_46098# a_518_46482# 0.001429f
C15706 a_1123_46634# a_1337_46116# 1.76e-19
C15707 a_n3674_39304# a_n3674_37592# 0.024803f
C15708 a_1414_42308# VDD 0.657887f
C15709 a_17730_32519# VREF_GND 0.241027f
C15710 a_4361_42308# a_5379_42460# 0.045451f
C15711 a_n1533_42852# COMP_P 0.001038f
C15712 a_5342_30871# a_13291_42460# 0.031084f
C15713 a_19237_31679# VIN_N 0.029585f
C15714 a_743_42282# a_4921_42308# 0.015669f
C15715 a_n1076_43230# a_n1630_35242# 2.32e-20
C15716 a_12545_42858# a_13622_42852# 1.46e-19
C15717 a_15279_43071# a_14635_42282# 2.87e-19
C15718 a_3381_47502# VDD 0.197761f
C15719 a_n2661_43370# a_2675_43914# 6.77e-21
C15720 a_n1151_42308# RST_Z 0.004602f
C15721 a_n863_45724# a_n1853_43023# 0.007839f
C15722 a_9290_44172# a_11136_42852# 0.001309f
C15723 a_10193_42453# a_12281_43396# 0.006314f
C15724 a_6171_45002# a_15493_43940# 5.86e-20
C15725 a_2063_45854# DATA[1] 8.67e-20
C15726 a_11827_44484# a_3422_30871# 0.076229f
C15727 a_18184_42460# a_20512_43084# 0.00468f
C15728 a_1307_43914# a_10405_44172# 0.010378f
C15729 a_13076_44458# a_13213_44734# 0.126609f
C15730 a_12607_44458# a_13857_44734# 0.002706f
C15731 a_12883_44458# a_13468_44734# 2.6e-19
C15732 SMPL_ON_N a_22521_40599# 1.14e-19
C15733 a_11823_42460# a_14205_43396# 0.176571f
C15734 a_11813_46116# a_11823_42460# 6.35e-21
C15735 a_11901_46660# a_12427_45724# 1.11e-19
C15736 a_11735_46660# a_12791_45546# 4.28e-19
C15737 a_n1151_42308# a_14403_45348# 1.39e-20
C15738 a_3090_45724# a_10180_45724# 4.56e-20
C15739 a_12465_44636# a_9482_43914# 0.069673f
C15740 a_6945_45028# a_22959_46124# 4.91e-20
C15741 a_22223_46124# a_10809_44734# 0.005525f
C15742 a_8199_44636# a_8049_45260# 0.069189f
C15743 a_765_45546# a_2277_45546# 3.26e-20
C15744 a_4791_45118# a_n2661_43370# 0.408007f
C15745 a_22612_30879# a_19963_31679# 0.078731f
C15746 a_4883_46098# a_13777_45326# 4.67e-21
C15747 a_11453_44696# a_11963_45334# 0.002899f
C15748 a_n1613_43370# a_4574_45260# 1.03e-20
C15749 a_n881_46662# a_3537_45260# 0.004983f
C15750 a_11309_47204# a_413_45260# 8.07e-21
C15751 a_5807_45002# a_n2017_45002# 2.87e-20
C15752 a_2903_42308# a_5934_30871# 2.52e-20
C15753 a_3823_42558# a_6123_31319# 1.19e-20
C15754 a_5379_42460# a_6761_42308# 1.12e-19
C15755 a_1606_42308# a_9223_42460# 1.69e-20
C15756 a_12281_43396# VDD 0.341026f
C15757 a_4921_42308# a_5755_42308# 0.175841f
C15758 a_2382_45260# a_1847_42826# 8.82e-20
C15759 a_n1899_43946# a_n1453_44318# 2.28e-19
C15760 a_n2065_43946# a_n875_44318# 2.56e-19
C15761 a_11967_42832# a_18079_43940# 0.052453f
C15762 a_2479_44172# a_3905_42865# 1.7e-19
C15763 a_n1059_45260# a_10083_42826# 0.006796f
C15764 a_n913_45002# a_8952_43230# 0.04786f
C15765 a_n2017_45002# a_10518_42984# 4.7e-20
C15766 a_5891_43370# a_9801_43940# 8.91e-19
C15767 a_4743_44484# a_3080_42308# 5.3e-21
C15768 a_949_44458# a_1427_43646# 2.11e-19
C15769 a_742_44458# a_1891_43646# 8.56e-19
C15770 a_15009_46634# VDD 0.205396f
C15771 a_2675_43914# a_2998_44172# 0.173844f
C15772 a_14084_46812# RST_Z 2.99e-19
C15773 a_n1549_44318# a_n3674_39768# 1.64e-19
C15774 a_n2661_42834# a_1443_43940# 0.001546f
C15775 a_14673_44172# a_15493_43940# 4.52e-20
C15776 a_14815_43914# a_14021_43940# 6.02e-20
C15777 a_n1925_42282# a_n2302_40160# 4.76e-20
C15778 a_n755_45592# a_8337_42558# 0.003302f
C15779 a_n357_42282# a_8325_42308# 5.17e-20
C15780 a_2957_45546# a_2711_45572# 0.056166f
C15781 a_n356_45724# a_603_45572# 6.01e-19
C15782 a_8049_45260# a_8192_45572# 0.008707f
C15783 a_768_44030# a_n2661_43922# 1.9176f
C15784 a_12891_46348# a_13213_44734# 0.052195f
C15785 a_12549_44172# a_n2293_43922# 0.194293f
C15786 a_n2293_46098# a_4574_45260# 0.001761f
C15787 a_12741_44636# a_6171_45002# 0.08387f
C15788 a_8953_45546# a_2437_43646# 1.66e-19
C15789 a_n2661_45546# a_1990_45572# 1.2e-19
C15790 a_13747_46662# a_9313_44734# 4.75e-21
C15791 a_18819_46122# a_19431_45546# 5.53e-19
C15792 a_18985_46122# a_18691_45572# 1.16e-19
C15793 a_19335_46494# a_18341_45572# 7.48e-19
C15794 a_472_46348# a_413_45260# 1.26e-19
C15795 a_376_46348# a_327_44734# 8.78e-20
C15796 a_16327_47482# a_20637_44484# 2.95e-19
C15797 a_4791_45118# a_2998_44172# 1.23e-19
C15798 a_n443_46116# a_2889_44172# 8.63e-19
C15799 a_3877_44458# a_5343_44458# 3.14e-20
C15800 a_n2438_43548# a_n356_44636# 0.082195f
C15801 a_12839_46116# a_13163_45724# 5.88e-19
C15802 a_n443_42852# a_1609_45822# 1.4e-19
C15803 a_n2302_39866# a_n2302_39072# 0.052227f
C15804 a_n4064_40160# a_n3565_38502# 0.028121f
C15805 a_n4315_30879# a_n3420_38528# 0.034192f
C15806 a_1606_42308# C8_P_btm 6.73e-20
C15807 a_n3674_38680# VDD 0.503323f
C15808 a_n784_42308# C0_N_btm 0.281635f
C15809 a_1209_47178# a_n1435_47204# 5.76e-19
C15810 a_4791_45118# a_4915_47217# 0.226891f
C15811 a_2063_45854# a_9863_47436# 0.12173f
C15812 a_9313_44734# a_10796_42968# 0.009402f
C15813 a_16375_45002# START 1.03e-19
C15814 a_18579_44172# a_20556_43646# 2.61e-19
C15815 a_18989_43940# a_19164_43230# 1.22e-19
C15816 a_742_44458# a_4149_42891# 2.67e-20
C15817 a_n2293_42834# a_n3674_37592# 0.025586f
C15818 a_16922_45042# a_20256_43172# 0.001682f
C15819 a_20692_30879# C1_N_btm 1.3e-20
C15820 a_1307_43914# a_6171_42473# 5.75e-21
C15821 a_n2293_43922# a_5111_42852# 9.71e-21
C15822 a_2711_45572# a_9482_43914# 0.01017f
C15823 a_n443_42852# a_501_45348# 1.56e-19
C15824 a_8162_45546# a_3537_45260# 2.11e-19
C15825 a_3316_45546# a_3602_45348# 0.001923f
C15826 a_7227_45028# a_7705_45326# 1.68e-19
C15827 a_12741_44636# a_14673_44172# 0.178572f
C15828 a_13249_42308# a_n913_45002# 0.019571f
C15829 a_3090_45724# a_5013_44260# 0.009874f
C15830 a_8696_44636# a_16789_45572# 3.81e-20
C15831 a_11415_45002# a_17517_44484# 0.006394f
C15832 a_1138_42852# a_n2661_42834# 0.024191f
C15833 a_7920_46348# a_7640_43914# 5.65e-22
C15834 a_12549_44172# a_n97_42460# 1.69e-19
C15835 a_15682_46116# a_16979_44734# 1.74e-20
C15836 a_13747_46662# a_20974_43370# 6.03e-20
C15837 a_n2293_46634# a_11173_43940# 2.54e-19
C15838 a_19321_45002# a_21381_43940# 3e-20
C15839 a_n2661_46634# a_n2442_46660# 0.063483f
C15840 a_n2956_39768# a_n2293_46634# 3.22e-21
C15841 a_n881_46662# a_1302_46660# 1.67e-19
C15842 VDAC_Ni RST_Z 1.24e-19
C15843 a_768_44030# a_1799_45572# 9.95e-20
C15844 VDAC_P C9_P_btm 0.123386p
C15845 a_11459_47204# a_11735_46660# 0.010464f
C15846 a_22609_38406# a_22705_37990# 3.51e-20
C15847 CAL_P a_22717_37285# 1.35e-20
C15848 a_7287_43370# a_4361_42308# 2.93e-20
C15849 a_1414_42308# a_n784_42308# 0.017857f
C15850 a_1667_45002# VDD 0.315476f
C15851 a_413_45260# START 0.035622f
C15852 a_10341_43396# a_16977_43638# 0.008076f
C15853 a_n97_42460# a_5111_42852# 5.6e-19
C15854 a_n1557_42282# a_n13_43084# 0.006682f
C15855 a_10807_43548# a_11136_42852# 0.006177f
C15856 a_458_43396# a_685_42968# 5.82e-20
C15857 a_8685_43396# a_15940_43402# 3.06e-19
C15858 a_6197_43396# a_5649_42852# 4.06e-21
C15859 a_9313_44734# a_4958_30871# 5.59e-19
C15860 a_644_44056# a_564_42282# 9.77e-22
C15861 a_13661_43548# a_19339_43156# 2.81e-20
C15862 a_584_46384# a_1184_42692# 3.73e-20
C15863 a_n1151_42308# a_n327_42558# 1.68e-19
C15864 a_9290_44172# a_9801_43940# 0.091547f
C15865 a_11652_45724# a_n2661_43922# 3.34e-21
C15866 a_7229_43940# a_5837_45028# 5.34e-21
C15867 a_11962_45724# a_n2661_42834# 3.66e-22
C15868 a_n863_45724# a_n1899_43946# 9.54e-20
C15869 a_8049_45260# a_8018_44260# 5.72e-20
C15870 a_375_42282# a_501_45348# 0.009374f
C15871 a_n2293_46634# a_13460_43230# 4.99e-21
C15872 a_2437_43646# a_20193_45348# 2.74e-21
C15873 a_n2293_45546# a_n1549_44318# 4.49e-19
C15874 a_3429_45260# a_n2661_43370# 0.004377f
C15875 a_n1079_45724# a_n1331_43914# 1.3e-20
C15876 a_6171_45002# a_n2293_42834# 0.035829f
C15877 a_15861_45028# a_16112_44458# 2.52e-20
C15878 a_8696_44636# a_14539_43914# 0.005592f
C15879 a_4185_45028# a_17538_32519# 0.043989f
C15880 a_5807_45002# a_13759_46122# 0.022269f
C15881 a_12549_44172# a_17957_46116# 8.35e-19
C15882 a_n743_46660# a_5497_46414# 0.005602f
C15883 a_n2661_46098# a_1208_46090# 0.023477f
C15884 a_6755_46942# a_765_45546# 0.002909f
C15885 a_13747_46662# a_12594_46348# 1.1e-19
C15886 a_n237_47217# a_n755_45592# 0.286948f
C15887 a_n1925_46634# a_6419_46155# 4.08e-20
C15888 a_13487_47204# a_14180_46482# 1.57e-20
C15889 a_12469_46902# a_12978_47026# 2.6e-19
C15890 a_11901_46660# a_12347_46660# 2.28e-19
C15891 a_11735_46660# a_12925_46660# 2.56e-19
C15892 a_11599_46634# a_12005_46436# 2.27e-19
C15893 a_n971_45724# a_1848_45724# 6.57e-22
C15894 a_327_47204# a_n1099_45572# 1.03e-21
C15895 a_n785_47204# a_310_45028# 9.87e-21
C15896 a_2107_46812# a_3147_46376# 0.010901f
C15897 a_n2661_46634# a_8953_45546# 8.33e-19
C15898 a_584_46384# a_n2293_45546# 0.029113f
C15899 a_4883_46098# a_5066_45546# 0.00636f
C15900 a_n2312_40392# a_n1925_42282# 0.002171f
C15901 a_n97_42460# a_9885_42308# 0.003237f
C15902 a_6765_43638# a_6123_31319# 1.83e-19
C15903 a_14543_43071# a_15279_43071# 4.07e-20
C15904 a_743_42282# a_13291_42460# 0.068071f
C15905 a_3626_43646# a_9803_42558# 0.006512f
C15906 a_14112_44734# VDD 0.004001f
C15907 a_1847_42826# a_1709_42852# 7.79e-21
C15908 a_12281_43396# a_n784_42308# 2.26e-20
C15909 a_15743_43084# a_20256_43172# 0.006046f
C15910 a_4185_45028# a_19339_43156# 2.91e-21
C15911 a_n443_42852# a_2437_43396# 2.27e-19
C15912 a_3065_45002# a_3600_43914# 0.011102f
C15913 a_n2661_45010# a_2537_44260# 6.6e-20
C15914 a_1138_42852# a_n2293_42282# 1.83e-20
C15915 a_n357_42282# a_9145_43396# 5.37e-19
C15916 a_n755_45592# a_8423_43396# 2.83e-20
C15917 a_9290_44172# a_12545_42858# 4.43e-19
C15918 a_8701_44490# a_5883_43914# 1.13e-20
C15919 a_3483_46348# a_13925_46122# 2.92e-19
C15920 a_167_45260# a_2324_44458# 0.001084f
C15921 a_n2840_46090# a_n2956_39304# 0.158668f
C15922 a_n1151_42308# a_3232_43370# 0.003308f
C15923 a_n443_46116# a_3537_45260# 0.003861f
C15924 a_4791_45118# a_4574_45260# 0.091783f
C15925 a_7227_47204# a_413_45260# 4.35e-19
C15926 a_n881_46662# a_16842_45938# 2.49e-19
C15927 a_12861_44030# a_n913_45002# 2.55e-20
C15928 a_10227_46804# a_3357_43084# 0.305304f
C15929 a_18780_47178# a_2437_43646# 0.008266f
C15930 a_13747_46662# a_15037_45618# 0.009886f
C15931 a_8349_46414# a_9625_46129# 7.25e-20
C15932 a_8199_44636# a_8953_45546# 0.71291f
C15933 a_8016_46348# a_9569_46155# 0.044705f
C15934 a_2063_45854# a_7229_43940# 0.003495f
C15935 a_765_45546# a_8049_45260# 6.27e-19
C15936 a_7715_46873# a_2711_45572# 8.9e-19
C15937 a_5257_43370# a_4099_45572# 1.01e-19
C15938 a_16327_47482# a_21297_45572# 6.03e-19
C15939 a_18597_46090# a_21513_45002# 0.00344f
C15940 a_n1190_43762# VDD 7.62e-19
C15941 a_18817_42826# a_17303_42282# 2.65e-20
C15942 a_17538_32519# VREF_GND 0.117023f
C15943 a_17333_42852# a_18057_42282# 3.02e-19
C15944 a_18083_42858# a_18727_42674# 3.76e-20
C15945 a_n1736_42282# COMP_P 0.005447f
C15946 a_n3674_38216# a_n1329_42308# 2.22e-19
C15947 a_n4318_38680# a_n4064_39072# 0.050323f
C15948 a_3080_42308# C0_N_btm 0.018211f
C15949 a_4185_45028# a_22465_38105# 0.065539f
C15950 a_1423_45028# a_8791_43396# 1.85e-20
C15951 a_18248_44752# a_15493_43396# 1.52e-20
C15952 a_18443_44721# a_18451_43940# 5.21e-19
C15953 a_18287_44626# a_19328_44172# 0.011011f
C15954 a_18374_44850# a_18326_43940# 9.6e-19
C15955 a_n2661_42834# a_n4318_39768# 0.031793f
C15956 a_11967_42832# a_17730_32519# 9.29e-22
C15957 a_20640_44752# a_21145_44484# 2.28e-19
C15958 a_n913_45002# a_19700_43370# 4.09e-21
C15959 a_n1059_45260# a_16664_43396# 9.44e-22
C15960 a_2959_46660# VDD 0.19762f
C15961 a_11827_44484# a_19808_44306# 2.85e-19
C15962 a_19279_43940# a_22315_44484# 1.97e-20
C15963 a_8696_44636# a_7871_42858# 3.01e-21
C15964 a_526_44458# a_9223_42460# 1.63e-20
C15965 a_10951_45334# a_10695_43548# 1.93e-21
C15966 a_1307_43914# a_3457_43396# 0.005402f
C15967 a_18184_42460# a_21381_43940# 0.003589f
C15968 a_6755_46942# a_16751_45260# 1.98e-19
C15969 a_8199_44636# a_8791_45572# 0.003441f
C15970 a_3090_45724# a_4927_45028# 0.088804f
C15971 a_13507_46334# a_n356_44636# 2.44e-20
C15972 a_13925_46122# a_14495_45572# 2.46e-19
C15973 a_14493_46090# a_13249_42308# 6.35e-19
C15974 a_19321_45002# a_19929_45028# 5.38e-19
C15975 a_10768_47026# a_10775_45002# 3.67e-22
C15976 a_13747_46662# a_18114_32519# 1.55e-19
C15977 a_18285_46348# a_2437_43646# 6.42e-20
C15978 a_n1613_43370# a_5883_43914# 0.352323f
C15979 a_11415_45002# a_19256_45572# 0.003224f
C15980 a_19511_42282# a_13258_32519# 0.072135f
C15981 a_17303_42282# a_21421_42336# 1.17e-19
C15982 a_6123_31319# a_1177_38525# 1.36e-19
C15983 a_n4318_37592# a_n4334_37440# 0.083644f
C15984 a_n913_45002# a_2123_42473# 0.029944f
C15985 a_10729_43914# a_10651_43940# 0.004213f
C15986 a_10405_44172# a_10867_43940# 0.022925f
C15987 a_n1441_43940# a_n4318_39304# 1.27e-19
C15988 a_644_44056# a_n1557_42282# 5.83e-21
C15989 a_1414_42308# a_3080_42308# 1.53e-19
C15990 a_n699_43396# a_2905_42968# 2.16e-19
C15991 a_n2017_45002# a_n327_42308# 2.31e-19
C15992 a_n1059_45260# a_2351_42308# 0.001198f
C15993 a_19335_46494# VDD 0.198512f
C15994 a_18985_46122# START 0.001317f
C15995 a_19553_46090# RST_Z 3.65e-21
C15996 a_14275_46494# CLK 3.42e-21
C15997 a_n2293_42834# a_8292_43218# 1.73e-19
C15998 a_18184_42460# a_18249_42858# 0.003882f
C15999 a_18494_42460# a_17333_42852# 0.00528f
C16000 a_2479_44172# a_4093_43548# 1.25e-20
C16001 a_895_43940# a_1756_43548# 1.47e-19
C16002 a_n2293_46098# a_5883_43914# 0.069185f
C16003 a_14495_45572# a_15599_45572# 5.49e-21
C16004 a_11823_42460# a_16680_45572# 3.71e-20
C16005 a_12427_45724# a_8696_44636# 4.63e-21
C16006 a_16375_45002# a_6171_45002# 0.026914f
C16007 a_n443_46116# a_1049_43396# 0.085877f
C16008 a_584_46384# a_2896_43646# 0.00371f
C16009 a_3147_46376# a_n2661_44458# 7.41e-21
C16010 a_11415_45002# a_13720_44458# 0.001979f
C16011 a_10490_45724# a_12561_45572# 0.001961f
C16012 a_12891_46348# a_11341_43940# 8.37e-19
C16013 a_12549_44172# a_21115_43940# 0.211261f
C16014 a_n2661_45546# a_n143_45144# 8.29e-19
C16015 a_n755_45592# a_n2017_45002# 0.088948f
C16016 a_n357_42282# a_n1059_45260# 7.3759f
C16017 a_15227_44166# a_15463_44811# 4.61e-19
C16018 a_n1079_45724# a_n967_45348# 4.19e-20
C16019 a_1609_45822# a_2437_43646# 0.189329f
C16020 a_13661_43548# a_17973_43940# 0.031319f
C16021 a_6945_45028# a_n2661_43370# 0.006001f
C16022 a_15143_45578# a_15297_45822# 0.008535f
C16023 a_10907_45822# a_10544_45572# 4.32e-19
C16024 a_12741_44636# a_12607_44458# 0.134974f
C16025 a_4185_45028# a_19721_31679# 0.004653f
C16026 a_n3565_38502# C10_P_btm 2.25e-20
C16027 a_n4209_37414# a_n3565_37414# 6.90997f
C16028 a_20990_47178# a_20916_46384# 4.4e-19
C16029 a_20894_47436# a_21588_30879# 1.66e-19
C16030 a_13507_46334# a_20843_47204# 4.38e-21
C16031 a_16327_47482# a_n743_46660# 0.53683f
C16032 a_10227_46804# a_n2293_46634# 0.032913f
C16033 a_n1741_47186# a_8667_46634# 4.44e-20
C16034 a_n1151_42308# a_4651_46660# 0.028941f
C16035 a_3785_47178# a_3877_44458# 5.26e-20
C16036 a_n2860_39866# VDD 0.004232f
C16037 a_12465_44636# a_13747_46662# 0.039773f
C16038 a_n4209_38502# C8_P_btm 5.41e-20
C16039 a_n4209_38216# a_n1838_35608# 1.13e-19
C16040 a_n971_45724# a_7411_46660# 0.567031f
C16041 a_2063_45854# a_5907_46634# 1.01e-19
C16042 a_2747_46873# a_768_44030# 0.00308f
C16043 a_4883_46098# a_19321_45002# 0.026904f
C16044 a_n1613_43370# a_n881_46662# 1.06426f
C16045 a_12429_44172# a_12379_42858# 5.92e-19
C16046 a_3626_43646# a_14579_43548# 1.34e-19
C16047 a_2982_43646# a_14205_43396# 1.37e-20
C16048 a_18494_42460# a_18997_42308# 0.002891f
C16049 a_20193_45348# a_19511_42282# 1.04e-19
C16050 a_5891_43370# a_5379_42460# 1.75e-20
C16051 a_n356_44636# a_7227_42308# 2.77e-19
C16052 a_n97_42460# a_16977_43638# 0.002871f
C16053 a_n1059_45260# CAL_N 0.001614f
C16054 a_n2293_43922# a_n1630_35242# 0.019388f
C16055 a_2998_44172# a_3059_42968# 5.55e-20
C16056 a_6547_43396# a_6643_43396# 0.013793f
C16057 a_6765_43638# a_6809_43396# 3.69e-19
C16058 a_20447_31679# a_22821_38993# 7.74e-20
C16059 a_6197_43396# a_8685_43396# 6.89e-20
C16060 a_3065_45002# a_4558_45348# 0.001793f
C16061 a_2382_45260# a_5111_44636# 1.01e-20
C16062 a_5937_45572# a_8333_44056# 7.94e-19
C16063 a_8016_46348# a_10405_44172# 0.098226f
C16064 a_17339_46660# a_18533_44260# 0.002232f
C16065 a_7499_43078# a_6298_44484# 1.09e-19
C16066 a_3090_45724# a_4699_43561# 1.16e-20
C16067 a_10227_46804# a_5342_30871# 0.163388f
C16068 a_n755_45592# a_n89_44484# 3.83e-19
C16069 a_13259_45724# a_17517_44484# 0.028602f
C16070 a_n2472_45546# a_n2661_43922# 2.25e-19
C16071 a_21076_30879# a_14021_43940# 1.4e-20
C16072 a_16327_47482# a_17701_42308# 0.001161f
C16073 a_3357_43084# a_1307_43914# 0.197864f
C16074 a_n881_46662# a_n2293_46098# 0.291354f
C16075 a_n1613_43370# a_n2157_46122# 0.296124f
C16076 a_n1151_42308# a_n1379_46482# 3.56e-19
C16077 a_4915_47217# a_6945_45028# 0.207881f
C16078 a_13487_47204# a_13925_46122# 1.5e-19
C16079 a_12861_44030# a_14493_46090# 7.43e-20
C16080 a_20916_46384# a_20273_46660# 2.16e-19
C16081 a_12549_44172# a_11415_45002# 0.028008f
C16082 a_5807_45002# a_16434_46660# 9.16e-19
C16083 a_4883_46098# a_5068_46348# 0.031466f
C16084 a_7927_46660# a_8035_47026# 0.057222f
C16085 a_3877_44458# a_3090_45724# 0.23348f
C16086 a_n237_47217# a_835_46155# 3.57e-20
C16087 a_10554_47026# a_10249_46116# 0.023301f
C16088 a_10623_46897# a_6755_46942# 0.008749f
C16089 a_7411_46660# a_8023_46660# 3.82e-19
C16090 a_10227_46804# a_9625_46129# 4.82e-19
C16091 a_14311_47204# a_13759_46122# 2.53e-21
C16092 a_11599_46634# a_12594_46348# 0.085826f
C16093 a_n3674_39768# a_n4334_39616# 0.05081f
C16094 a_n699_43396# VDD 0.922998f
C16095 a_5649_42852# a_10922_42852# 1.52e-20
C16096 a_4190_30871# a_5534_30871# 0.020828f
C16097 a_n97_42460# a_n1630_35242# 0.035802f
C16098 a_2982_43646# a_22400_42852# 3.1e-21
C16099 a_16823_43084# a_16795_42852# 0.065873f
C16100 a_4361_42308# a_12089_42308# 0.006552f
C16101 a_18114_32519# VCM 0.121302f
C16102 a_19721_31679# VREF_GND 0.001975f
C16103 a_15493_43940# a_15959_42545# 1.59e-20
C16104 a_n4318_39768# a_n3565_39590# 9.85e-20
C16105 a_743_42282# a_13460_43230# 1.8e-20
C16106 a_15743_43084# a_21195_42852# 0.004294f
C16107 a_4185_45028# a_22591_43396# 0.008398f
C16108 a_n2661_45546# a_n97_42460# 0.038952f
C16109 a_626_44172# a_700_44734# 1.02e-19
C16110 a_11322_45546# a_11341_43940# 2.88e-20
C16111 a_7499_43078# a_10555_44260# 0.03816f
C16112 a_n2661_43370# a_8103_44636# 5.82e-21
C16113 a_7229_43940# a_n2661_42834# 0.023622f
C16114 a_18184_42460# a_19929_45028# 0.001333f
C16115 a_16327_47482# a_21613_42308# 1.68e-19
C16116 a_17715_44484# a_17499_43370# 0.001287f
C16117 a_13507_46334# a_18727_42674# 0.093566f
C16118 a_10907_45822# a_10949_43914# 2.73e-20
C16119 a_n881_46662# a_7230_45938# 8.9e-20
C16120 a_n1613_43370# a_8162_45546# 1.42e-20
C16121 a_n743_46660# a_n356_45724# 0.223429f
C16122 a_1123_46634# a_n755_45592# 1.46e-19
C16123 a_948_46660# a_n357_42282# 1.33e-19
C16124 a_13747_46662# a_2711_45572# 0.032065f
C16125 a_10623_46897# a_8049_45260# 9.22e-20
C16126 a_15227_44166# a_21137_46414# 0.081665f
C16127 a_14513_46634# a_13925_46122# 2.11e-19
C16128 a_14180_46812# a_14493_46090# 1.41e-20
C16129 a_18834_46812# a_6945_45028# 1.91e-20
C16130 a_16292_46812# a_10809_44734# 0.005743f
C16131 a_14035_46660# a_14275_46494# 3.12e-19
C16132 a_n2293_46098# a_n2157_46122# 0.015455f
C16133 a_765_45546# a_8953_45546# 3.61e-19
C16134 a_12861_44030# a_15903_45785# 0.156145f
C16135 a_n2293_46634# a_n906_45572# 5.29e-19
C16136 a_n2661_46098# a_n2661_45546# 0.011799f
C16137 a_19466_46812# a_19900_46494# 2.79e-19
C16138 a_19692_46634# a_20075_46420# 5.36e-19
C16139 a_13059_46348# a_10903_43370# 0.11738f
C16140 a_n2472_46090# a_n1853_46287# 8.45e-19
C16141 a_11599_46634# a_15037_45618# 1.12e-19
C16142 a_11453_44696# a_13249_42308# 0.026348f
C16143 a_21259_43561# a_13258_32519# 3.03e-20
C16144 a_4190_30871# a_19647_42308# 0.001077f
C16145 a_n2293_42282# a_1576_42282# 3.68e-19
C16146 a_4361_42308# a_18907_42674# 0.010379f
C16147 a_13887_32519# a_4958_30871# 0.030919f
C16148 a_22959_43948# VDD 0.297936f
C16149 a_5649_42852# a_17531_42308# 5.44e-20
C16150 a_8387_43230# a_8791_42308# 0.001415f
C16151 a_9127_43156# a_8685_42308# 2.44e-19
C16152 a_15493_43940# RST_Z 0.004544f
C16153 a_5343_44458# a_5244_44056# 8.23e-19
C16154 a_9313_44734# a_19615_44636# 1.67e-21
C16155 a_4223_44672# a_5663_43940# 0.01368f
C16156 a_n1059_45260# a_n144_43396# 8.85e-20
C16157 a_16922_45042# a_15493_43396# 5.34e-20
C16158 a_2266_47243# VDD 6.34e-20
C16159 a_n2956_39304# a_n2104_42282# 2.99e-20
C16160 a_n2956_38680# a_n4318_38216# 0.023189f
C16161 a_5205_44484# a_n97_42460# 1.83e-20
C16162 a_2382_45260# a_4235_43370# 0.006145f
C16163 a_n1352_44484# a_n4318_39768# 3e-19
C16164 a_2487_47570# DATA[1] 7.79e-21
C16165 SMPL_ON_N VIN_N 0.587565f
C16166 a_n443_42852# a_5534_30871# 8.98e-20
C16167 a_n357_42282# a_19987_42826# 0.016903f
C16168 a_n2661_43370# a_11173_44260# 2.7e-19
C16169 a_n2956_38216# a_n2293_42282# 2.83e-20
C16170 a_15861_45028# a_17499_43370# 6.09e-20
C16171 a_8696_44636# a_17324_43396# 5.68e-21
C16172 a_2437_43646# a_2437_43396# 0.009374f
C16173 a_10249_46116# a_2437_43646# 1.78e-19
C16174 a_11453_44696# a_17613_45144# 3.78e-19
C16175 a_2324_44458# a_n863_45724# 0.01106f
C16176 a_4419_46090# a_2711_45572# 0.026096f
C16177 a_10227_46804# a_16237_45028# 7.21e-19
C16178 a_n2293_46634# a_1307_43914# 0.184387f
C16179 a_5937_45572# a_n443_42852# 5.42e-20
C16180 a_3877_44458# a_2274_45254# 7.27e-21
C16181 a_4955_46873# a_413_45260# 2.73e-20
C16182 a_11415_45002# a_11525_45546# 1.34e-19
C16183 a_10467_46802# a_3357_43084# 1.38e-20
C16184 a_3090_45724# a_18175_45572# 0.130163f
C16185 a_14976_45028# a_16147_45260# 0.001993f
C16186 a_n2497_47436# a_n1243_44484# 2.69e-19
C16187 a_3483_46348# a_5263_45724# 9.89e-20
C16188 a_4791_45118# a_5883_43914# 7.11e-19
C16189 a_n743_46660# a_14537_43396# 6.18e-20
C16190 a_13507_46334# a_20567_45036# 2.05e-21
C16191 a_4883_46098# a_18184_42460# 6.32e-21
C16192 a_5342_30871# CAL_P 0.007017f
C16193 a_13575_42558# a_14113_42308# 0.11418f
C16194 a_n3674_37592# a_n4064_39616# 0.019733f
C16195 a_n3674_38216# a_n4334_39392# 9.02e-20
C16196 a_14209_32519# VREF 2.95e-20
C16197 a_n4318_38680# VDD 0.417422f
C16198 a_13887_32519# VCM 0.011087f
C16199 a_n1630_35242# a_n3420_39616# 0.001297f
C16200 a_19279_43940# a_19319_43548# 0.023499f
C16201 a_18579_44172# a_18533_44260# 0.001461f
C16202 a_5891_43370# a_7287_43370# 0.008619f
C16203 a_n2293_42834# a_3681_42891# 0.006112f
C16204 a_10193_42453# a_11551_42558# 0.228057f
C16205 a_22959_46660# VDD 0.299681f
C16206 a_12741_44636# RST_Z 0.004532f
C16207 a_11827_44484# a_21487_43396# 3.48e-20
C16208 a_18184_42460# a_5649_42852# 0.028842f
C16209 a_15004_44636# a_14955_43396# 6.17e-20
C16210 a_14539_43914# a_14205_43396# 0.001533f
C16211 a_10057_43914# a_12281_43396# 5.88e-20
C16212 a_n2956_38216# a_n3565_39590# 0.021271f
C16213 a_2711_45572# a_4958_30871# 1.35e-20
C16214 a_n2810_45572# a_n2946_39866# 4.32e-20
C16215 a_n913_45002# a_8495_42852# 0.030544f
C16216 a_3537_45260# a_4649_43172# 5.06e-19
C16217 a_1307_43914# a_5342_30871# 5.9e-20
C16218 a_11691_44458# a_4190_30871# 0.002426f
C16219 a_20193_45348# a_21259_43561# 6.39e-21
C16220 a_12861_44030# a_18451_43940# 0.001042f
C16221 a_12594_46348# a_13348_45260# 7.19e-21
C16222 a_7230_45938# a_8162_45546# 1.68e-19
C16223 a_3090_45724# a_10440_44484# 1.35e-20
C16224 a_19240_46482# a_18341_45572# 1.94e-19
C16225 a_18051_46116# a_16147_45260# 5.51e-19
C16226 a_8049_45260# a_21513_45002# 0.007177f
C16227 a_10227_46804# a_9672_43914# 6.27e-19
C16228 a_10903_43370# a_13556_45296# 2.71e-19
C16229 a_2711_45572# a_6469_45572# 2.38e-19
C16230 a_2324_44458# a_8191_45002# 0.120399f
C16231 a_167_45260# a_2448_45028# 1.54e-19
C16232 a_11415_45002# a_15685_45394# 1.56e-19
C16233 a_768_44030# a_n809_44244# 4.27e-19
C16234 a_20623_46660# a_20567_45036# 3.11e-20
C16235 a_13759_46122# a_13017_45260# 9.47e-21
C16236 a_n4064_40160# VDAC_P 0.001245f
C16237 a_4958_30871# EN_VIN_BSTR_N 0.021638f
C16238 a_n4209_39304# a_n4209_37414# 0.029637f
C16239 a_12861_44030# a_11453_44696# 0.173308f
C16240 a_13717_47436# a_22959_47212# 8.82e-19
C16241 a_10227_46804# a_18597_46090# 0.07604f
C16242 a_n3420_37984# a_n2946_37984# 0.238664f
C16243 a_n3690_38304# a_n4064_37984# 0.085872f
C16244 a_n3565_38216# a_n2302_37984# 0.067194f
C16245 a_n4334_38304# a_n4251_38304# 0.007692f
C16246 a_n4209_38216# a_n3607_38304# 0.002352f
C16247 a_11551_42558# VDD 0.192086f
C16248 a_n1435_47204# a_n2312_40392# 0.002491f
C16249 a_4791_45118# a_n881_46662# 0.429542f
C16250 a_15811_47375# a_4883_46098# 1.03e-21
C16251 a_16241_47178# a_13507_46334# 6.13e-21
C16252 a_n443_46116# a_n1613_43370# 0.410263f
C16253 a_4915_47217# a_3411_47243# 2.39e-21
C16254 a_18143_47464# a_18780_47178# 0.001596f
C16255 a_11599_46634# a_12465_44636# 0.018625f
C16256 a_2063_45854# a_768_44030# 0.027746f
C16257 a_n2833_47464# a_n2840_46634# 0.019713f
C16258 a_22465_38105# a_22469_40625# 0.072192f
C16259 a_5742_30871# RST_Z 0.003575f
C16260 a_15493_43940# a_16243_43396# 0.006124f
C16261 a_11341_43940# a_16409_43396# 4.02e-20
C16262 a_5024_45822# VDD 0.004293f
C16263 a_19328_44172# a_19268_43646# 9.49e-19
C16264 a_15493_43396# a_15743_43084# 0.517624f
C16265 a_11967_42832# a_19339_43156# 9.23e-20
C16266 a_9313_44734# a_11229_43218# 1.2e-19
C16267 a_18248_44752# a_18707_42852# 7.68e-22
C16268 a_n2810_45028# a_n4209_38502# 0.022376f
C16269 a_104_43370# a_n1557_42282# 6.03e-21
C16270 a_n2433_43396# a_n1243_43396# 2.56e-19
C16271 a_n97_42460# a_1427_43646# 0.047018f
C16272 a_1209_43370# a_1568_43370# 9.57e-19
C16273 a_2437_43646# a_22223_45572# 0.165664f
C16274 a_2711_45572# a_18911_45144# 3.83e-20
C16275 a_n2293_45546# a_n1177_44458# 3.48e-19
C16276 a_14033_45822# a_9482_43914# 8.97e-21
C16277 a_n443_42852# a_11691_44458# 4.69e-20
C16278 a_n2293_46634# a_9396_43370# 0.012588f
C16279 a_18479_47436# a_4190_30871# 1.1e-19
C16280 a_10227_46804# a_743_42282# 0.045325f
C16281 a_12891_46348# a_10341_43396# 7.46e-20
C16282 a_10809_44734# a_10809_44484# 0.009578f
C16283 a_18189_46348# a_17517_44484# 1.78e-19
C16284 a_4185_45028# a_22591_44484# 0.013394f
C16285 a_16327_47482# a_4361_42308# 0.029635f
C16286 a_13059_46348# a_14955_43940# 0.001717f
C16287 a_21513_45002# a_19479_31679# 0.005077f
C16288 a_310_45028# a_n2661_44458# 0.003131f
C16289 a_13259_45724# a_13720_44458# 0.016851f
C16290 a_4883_46098# a_13059_46348# 0.097406f
C16291 a_18597_46090# a_17339_46660# 0.018491f
C16292 a_16327_47482# a_20841_46902# 8.93e-20
C16293 a_5807_45002# a_8189_46660# 7.17e-19
C16294 a_2124_47436# a_1823_45246# 9.81e-21
C16295 a_12549_44172# a_12251_46660# 0.001402f
C16296 a_12891_46348# a_12991_46634# 0.018656f
C16297 a_n443_46116# a_n2293_46098# 0.251135f
C16298 a_19864_35138# VIN_N 0.367112f
C16299 a_13507_46334# a_16721_46634# 0.00543f
C16300 a_10227_46804# a_19123_46287# 9.33e-20
C16301 a_18143_47464# a_18285_46348# 2.02e-19
C16302 a_18780_47178# a_765_45546# 2.8e-19
C16303 a_3699_46634# a_3877_44458# 0.087244f
C16304 a_2864_46660# a_3055_46660# 4.61e-19
C16305 a_2959_46660# a_4646_46812# 8.56e-21
C16306 a_n1741_47186# a_5204_45822# 4.65e-20
C16307 a_n2661_46634# a_10249_46116# 0.055133f
C16308 a_584_46384# a_1138_42852# 0.491749f
C16309 a_n1151_42308# a_n1076_46494# 0.023834f
C16310 a_2063_45854# a_1176_45822# 2.25e-19
C16311 EN_VIN_BSTR_N VCM 0.927905f
C16312 a_12861_44030# a_17639_46660# 0.033515f
C16313 C4_N_btm C7_N_btm 0.148546f
C16314 C5_N_btm C6_N_btm 18.2841f
C16315 C1_N_btm C10_N_btm 0.204172f
C16316 C2_N_btm C9_N_btm 0.144261f
C16317 C3_N_btm C8_N_btm 0.13616f
C16318 a_1239_47204# a_167_45260# 2.52e-21
C16319 a_n237_47217# a_3483_46348# 0.090759f
C16320 a_n971_45724# a_4185_45028# 4.59e-19
C16321 a_n743_46660# a_8667_46634# 9.34e-20
C16322 a_2443_46660# a_4817_46660# 2.35e-21
C16323 a_11599_46634# a_20528_46660# 2.63e-20
C16324 a_20512_43084# a_17303_42282# 4.29e-20
C16325 a_19721_31679# a_22469_40625# 1.46e-20
C16326 a_n2661_42282# a_6481_42558# 0.001754f
C16327 a_9803_43646# a_9127_43156# 3.02e-19
C16328 a_9145_43396# a_8952_43230# 1.61e-20
C16329 a_n1925_42282# a_n2433_43396# 0.001028f
C16330 a_5111_44636# a_5343_44458# 0.477401f
C16331 a_4927_45028# a_4743_44484# 3.54e-19
C16332 a_5147_45002# a_5518_44484# 0.064422f
C16333 a_n443_42852# a_8333_44056# 3.11e-19
C16334 a_n357_42282# a_18326_43940# 6.84e-21
C16335 a_n2661_45010# a_n1190_44850# 2.49e-19
C16336 a_17478_45572# a_17517_44484# 7.16e-22
C16337 a_3232_43370# a_4223_44672# 0.033907f
C16338 a_3537_45260# a_8701_44490# 5.76e-20
C16339 a_5937_45572# a_6655_43762# 8.87e-19
C16340 a_7735_45067# a_n2661_43370# 2.56e-19
C16341 a_1307_43914# a_16237_45028# 0.056593f
C16342 a_17339_46660# a_743_42282# 4.84e-20
C16343 a_12741_44636# a_16243_43396# 5.87e-20
C16344 a_5807_45002# a_12379_46436# 0.006522f
C16345 a_12549_44172# a_13259_45724# 0.110646f
C16346 a_6755_46942# a_8349_46414# 0.001141f
C16347 a_10249_46116# a_8199_44636# 0.002313f
C16348 a_4791_45118# a_8162_45546# 3.59e-20
C16349 a_6151_47436# a_4880_45572# 9.96e-20
C16350 a_8270_45546# a_3483_46348# 0.058754f
C16351 a_11599_46634# a_2711_45572# 0.018466f
C16352 a_765_45546# a_18285_46348# 5.85e-19
C16353 a_n1151_42308# a_10193_42453# 0.238612f
C16354 a_2063_45854# a_11652_45724# 0.002983f
C16355 a_10150_46912# a_9823_46155# 5.05e-19
C16356 a_9863_46634# a_10355_46116# 0.00109f
C16357 a_2107_46812# a_3873_46454# 4.52e-19
C16358 a_n13_43084# a_n3674_37592# 1.17e-20
C16359 a_n2293_42282# a_4649_42852# 5.38e-20
C16360 a_17730_32519# VREF 1.53e-20
C16361 a_1467_44172# VDD 0.391994f
C16362 a_4361_42308# a_5267_42460# 0.005989f
C16363 a_743_42282# a_4933_42558# 0.001023f
C16364 a_5534_30871# a_14635_42282# 0.020227f
C16365 a_n901_43156# a_n1630_35242# 3e-19
C16366 a_n1151_42308# VDD 2.57238f
C16367 a_19610_45572# a_19319_43548# 1.39e-20
C16368 a_13777_45326# a_13483_43940# 5.57e-20
C16369 a_13556_45296# a_14955_43940# 0.059957f
C16370 a_n863_45724# a_n2157_42858# 7.79e-21
C16371 a_9290_44172# a_13157_43218# 8.98e-21
C16372 a_10193_42453# a_12293_43646# 9.47e-19
C16373 a_n2312_38680# a_n4209_38216# 2.66e-20
C16374 a_584_46384# DATA[1] 0.007084f
C16375 a_11691_44458# a_18753_44484# 0.005052f
C16376 a_n2293_42834# a_5663_43940# 4.43e-21
C16377 a_1307_43914# a_9672_43914# 0.007152f
C16378 a_11827_44484# a_21398_44850# 0.003647f
C16379 a_13076_44458# a_n2293_43922# 5.37e-19
C16380 a_12883_44458# a_13213_44734# 0.002706f
C16381 a_12607_44458# a_13468_44734# 1.09e-19
C16382 a_11823_42460# a_14358_43442# 0.122636f
C16383 a_13249_42308# a_9145_43396# 0.072489f
C16384 a_11735_46660# a_11823_42460# 6.67e-20
C16385 a_11901_46660# a_11962_45724# 3.74e-20
C16386 a_n881_46662# a_3429_45260# 1.13e-19
C16387 a_12465_44636# a_13348_45260# 1.39e-21
C16388 a_6945_45028# a_10809_44734# 0.953135f
C16389 a_9625_46129# a_8034_45724# 1.73e-19
C16390 a_8349_46414# a_8049_45260# 2.39e-20
C16391 a_8199_44636# a_8781_46436# 2.2e-19
C16392 a_765_45546# a_1609_45822# 0.021736f
C16393 a_6151_47436# a_8560_45348# 1.29e-20
C16394 a_21076_30879# a_20692_30879# 0.117886f
C16395 a_21588_30879# a_19963_31679# 0.055898f
C16396 a_13507_46334# a_14180_45002# 1.58e-22
C16397 a_n1613_43370# a_3537_45260# 0.095192f
C16398 a_11453_44696# a_11787_45002# 0.005756f
C16399 a_2713_42308# a_5934_30871# 1.48e-20
C16400 a_3318_42354# a_6123_31319# 1.13e-20
C16401 a_1606_42308# a_8791_42308# 3.31e-20
C16402 a_5534_30871# a_n3420_37984# 0.043974f
C16403 a_5267_42460# a_6761_42308# 6.68e-20
C16404 a_n784_42308# a_11551_42558# 2.06e-20
C16405 a_16877_42852# a_4958_30871# 6.91e-19
C16406 a_12293_43646# VDD 0.005635f
C16407 a_9803_43646# CLK 2.81e-19
C16408 a_n1059_45260# a_8952_43230# 0.010945f
C16409 a_n913_45002# a_9127_43156# 0.038139f
C16410 a_n2017_45002# a_10083_42826# 1.71e-19
C16411 a_5891_43370# a_9420_43940# 4.11e-19
C16412 a_4743_44484# a_4699_43561# 6.57e-20
C16413 a_949_44458# a_n1557_42282# 1.2e-19
C16414 a_742_44458# a_1427_43646# 5.41e-19
C16415 a_14084_46812# VDD 0.087769f
C16416 a_2675_43914# a_2889_44172# 0.083573f
C16417 a_895_43940# a_2998_44172# 2.2e-19
C16418 a_13607_46688# RST_Z 3.83e-19
C16419 a_1307_43914# a_743_42282# 5.15e-19
C16420 a_n1899_43946# a_n1644_44306# 0.06121f
C16421 a_n1331_43914# a_n3674_39768# 6.83e-20
C16422 a_11967_42832# a_17973_43940# 0.070514f
C16423 a_4223_44672# a_4905_42826# 3.85e-20
C16424 a_n699_43396# a_3080_42308# 0.001343f
C16425 a_n2661_42834# a_1241_43940# 0.003456f
C16426 a_17517_44484# a_20935_43940# 1.78e-20
C16427 a_n755_45592# a_4169_42308# 1.51e-19
C16428 a_n356_45724# a_509_45572# 9.76e-19
C16429 a_12839_46116# a_12791_45546# 2.39e-19
C16430 a_8049_45260# a_8120_45572# 0.0028f
C16431 a_768_44030# a_n2661_42834# 4.99505f
C16432 a_12549_44172# a_n2661_43922# 0.061277f
C16433 a_12891_46348# a_n2293_43922# 8.04e-19
C16434 a_n2293_46098# a_3537_45260# 0.019207f
C16435 a_12741_44636# a_3232_43370# 4.67e-19
C16436 a_5937_45572# a_2437_43646# 3.38e-20
C16437 a_n755_45592# a_4099_45572# 0.001267f
C16438 a_n2661_45546# a_3733_45822# 1.54e-35
C16439 a_13661_43548# a_9313_44734# 3.79e-19
C16440 a_18819_46122# a_18691_45572# 5.44e-20
C16441 a_376_46348# a_413_45260# 1.85e-19
C16442 a_11453_44696# a_17325_44484# 1.07e-19
C16443 a_8016_46348# a_3357_43084# 1.25e-21
C16444 a_n443_46116# a_2675_43914# 0.011921f
C16445 a_n743_46660# a_n356_44636# 4.32e-20
C16446 a_16327_47482# a_20397_44484# 0.001966f
C16447 a_18597_46090# a_18579_44172# 9.48e-21
C16448 a_22765_42852# RST_Z 1.67e-19
C16449 a_327_47204# a_n1435_47204# 0.001005f
C16450 a_4791_45118# a_n443_46116# 0.115639f
C16451 a_4700_47436# a_4915_47217# 0.07122f
C16452 a_2063_45854# a_9067_47204# 1.79e-19
C16453 a_n1151_42308# a_6491_46660# 1.03e-19
C16454 a_3785_47178# a_6151_47436# 4.24e-20
C16455 a_n3420_39616# a_n3607_39392# 6.01e-19
C16456 a_n4064_40160# a_n4334_38528# 0.007725f
C16457 a_1606_42308# C9_P_btm 9.33e-20
C16458 a_n2840_42282# VDD 0.294987f
C16459 a_n784_42308# C0_dummy_N_btm 2.62e-20
C16460 a_9313_44734# a_10835_43094# 0.050385f
C16461 a_19478_44306# a_3626_43646# 6.67e-20
C16462 a_n913_45002# a_17124_42282# 4.89e-19
C16463 a_19240_46482# VDD 0.077608f
C16464 a_18579_44172# a_743_42282# 9.34e-19
C16465 a_n356_44636# a_17701_42308# 0.065679f
C16466 a_742_44458# a_3863_42891# 4.92e-20
C16467 a_n2661_43370# a_n3674_38216# 1.63e-20
C16468 a_3232_43370# a_5742_30871# 6.51e-20
C16469 a_20692_30879# C0_N_btm 9.35e-21
C16470 a_n2293_42834# a_n327_42558# 0.001338f
C16471 a_1307_43914# a_5755_42308# 1.01e-20
C16472 a_3422_30871# a_16823_43084# 4.23e-21
C16473 a_n2661_42834# a_5755_42852# 1.12e-20
C16474 a_n2661_43922# a_5111_42852# 3.12e-21
C16475 a_n2293_43922# a_4520_42826# 1.13e-20
C16476 a_2711_45572# a_13348_45260# 7.14e-20
C16477 a_n443_42852# a_375_42282# 0.075658f
C16478 a_6945_45028# a_5883_43914# 1.46e-20
C16479 a_8049_45260# a_22959_45036# 0.002194f
C16480 a_12861_44030# a_9145_43396# 1.84e-19
C16481 a_3316_45546# a_3495_45348# 0.004904f
C16482 a_7227_45028# a_6709_45028# 0.115677f
C16483 a_4185_45028# a_9313_44734# 0.078424f
C16484 a_11823_42460# en_comp 8.68e-21
C16485 a_12741_44636# a_14581_44484# 2.79e-20
C16486 a_13249_42308# a_n1059_45260# 0.026496f
C16487 a_16680_45572# a_16789_45572# 0.007416f
C16488 a_16855_45546# a_17034_45572# 0.007399f
C16489 a_3090_45724# a_5244_44056# 0.002228f
C16490 a_20202_43084# a_17517_44484# 0.021286f
C16491 a_4880_45572# a_5111_44636# 3.99e-20
C16492 a_526_44458# a_n2129_44697# 4.74e-20
C16493 a_15682_46116# a_14539_43914# 2.11e-19
C16494 a_n2293_46634# a_10867_43940# 7.16e-19
C16495 VDAC_P C10_P_btm 0.24639p
C16496 a_n2840_46634# a_n2293_46634# 2.97e-19
C16497 a_n2661_46634# a_n2472_46634# 0.0842f
C16498 a_n2956_39768# a_n2442_46660# 6.5214f
C16499 a_n881_46662# a_1057_46660# 1.39e-19
C16500 a_n1613_43370# a_1302_46660# 0.001965f
C16501 VDAC_Ni VDD 0.288547f
C16502 a_4883_46098# a_7577_46660# 7.2e-20
C16503 a_22609_38406# a_22609_37990# 0.32625f
C16504 CAL_P a_22705_37990# 1.58e-20
C16505 a_10227_46804# a_6755_46942# 0.778648f
C16506 a_6547_43396# a_4361_42308# 2.77e-20
C16507 a_1414_42308# a_196_42282# 6.32e-21
C16508 a_327_44734# VDD 0.667364f
C16509 a_10341_43396# a_16409_43396# 0.028466f
C16510 a_12281_43396# a_13943_43396# 6.37e-21
C16511 a_413_45260# RST_Z 0.199496f
C16512 a_n97_42460# a_4520_42826# 4.68e-20
C16513 a_n1557_42282# a_n1076_43230# 3.53e-20
C16514 a_9396_43370# a_743_42282# 5.17e-20
C16515 a_n984_44318# a_n1630_35242# 1.73e-21
C16516 a_8685_43396# a_15868_43402# 4.99e-20
C16517 a_6293_42852# a_5649_42852# 2.33e-19
C16518 a_13661_43548# a_18599_43230# 0.001237f
C16519 a_768_44030# a_n2293_42282# 1.83e-20
C16520 a_584_46384# a_1576_42282# 6.73e-21
C16521 a_n1151_42308# a_n784_42308# 0.154055f
C16522 a_9290_44172# a_9420_43940# 0.002091f
C16523 a_n863_45724# a_n1761_44111# 6.9e-20
C16524 a_10227_46804# a_16328_43172# 1.46e-21
C16525 a_2107_46812# a_9127_43156# 6e-20
C16526 a_11525_45546# a_n2661_43922# 1.39e-20
C16527 a_n2661_45546# a_n984_44318# 1.23e-21
C16528 a_19479_31679# a_22959_45036# 0.018372f
C16529 a_n2293_46634# a_13635_43156# 1.15e-19
C16530 a_21513_45002# a_20193_45348# 3.14e-20
C16531 a_n1079_45724# a_n1899_43946# 1.2e-21
C16532 a_3065_45002# a_n2661_43370# 0.356646f
C16533 a_6171_45002# a_7639_45394# 3.69e-19
C16534 a_2711_45572# a_19615_44636# 2.24e-21
C16535 a_3232_43370# a_n2293_42834# 0.041207f
C16536 a_8696_44636# a_16112_44458# 0.004409f
C16537 a_16855_45546# a_16979_44734# 2.49e-21
C16538 a_16680_45572# a_14539_43914# 2.31e-19
C16539 a_4185_45028# a_20974_43370# 0.184625f
C16540 a_1307_43914# a_626_44172# 6.24e-19
C16541 a_13059_46348# a_8685_43396# 0.002513f
C16542 a_2324_44458# a_2455_43940# 1.69e-19
C16543 a_12549_44172# a_18189_46348# 2.08e-19
C16544 a_n743_46660# a_5204_45822# 0.034798f
C16545 a_n2661_46098# a_805_46414# 0.044109f
C16546 a_1799_45572# a_1208_46090# 0.008066f
C16547 a_10249_46116# a_765_45546# 0.005411f
C16548 a_n881_46662# a_6945_45028# 0.239384f
C16549 a_15368_46634# a_15227_44166# 0.002374f
C16550 a_3090_45724# a_19466_46812# 1.49e-19
C16551 a_5807_45002# a_13351_46090# 0.002035f
C16552 a_13661_43548# a_12594_46348# 1.57e-21
C16553 a_n971_45724# a_997_45618# 4.51e-22
C16554 a_n746_45260# a_n755_45592# 0.172774f
C16555 a_n237_47217# a_n357_42282# 4.85e-21
C16556 a_n1925_46634# a_6165_46155# 6.31e-20
C16557 a_11901_46660# a_12978_47026# 1.46e-19
C16558 a_10227_46804# a_8049_45260# 0.058336f
C16559 a_4883_46098# a_5431_46482# 2.13e-19
C16560 a_n2293_46634# a_8016_46348# 4.84e-19
C16561 a_n2661_46634# a_5937_45572# 2.16e-19
C16562 a_2107_46812# a_2804_46116# 0.008475f
C16563 a_n23_47502# a_310_45028# 6.86e-20
C16564 a_n785_47204# a_n1099_45572# 1.19e-20
C16565 a_327_47204# a_380_45546# 1.52e-21
C16566 a_21381_43940# a_17303_42282# 4.27e-20
C16567 a_14401_32519# a_4958_30871# 0.079459f
C16568 a_n97_42460# a_15720_42674# 5.52e-19
C16569 a_6547_43396# a_6761_42308# 1.18e-20
C16570 a_3935_42891# a_4156_43218# 0.007833f
C16571 a_14543_43071# a_5534_30871# 0.196814f
C16572 a_13460_43230# a_15279_43071# 2.03e-20
C16573 a_6197_43396# a_6123_31319# 1.52e-19
C16574 a_17730_32519# a_22521_40599# 1.2e-20
C16575 a_19319_43548# a_19332_42282# 8.34e-20
C16576 a_3626_43646# a_9223_42460# 0.002263f
C16577 a_13857_44734# VDD 0.18416f
C16578 a_13635_43156# a_5342_30871# 0.001254f
C16579 a_15743_43084# a_18707_42852# 8.78e-20
C16580 a_9290_44172# a_12089_42308# 0.047614f
C16581 a_4185_45028# a_18599_43230# 1.09e-20
C16582 a_3065_45002# a_2998_44172# 0.024536f
C16583 a_n2293_45010# a_1241_44260# 1.56e-19
C16584 a_n2661_45010# a_2253_44260# 5.46e-19
C16585 a_10903_43370# a_10991_42826# 9.88e-21
C16586 a_n967_45348# a_n3674_39768# 2.29e-20
C16587 w_11334_34010# CAL_P 0.063131f
C16588 a_n357_42282# a_8423_43396# 1.68e-19
C16589 a_n755_45592# a_8317_43396# 0.007502f
C16590 a_3537_45260# a_2675_43914# 2.19e-19
C16591 a_2382_45260# a_3905_42865# 0.291572f
C16592 a_4223_44672# a_8975_43940# 1.67e-19
C16593 w_1575_34946# VIN_P 2.57e-20
C16594 a_18597_46090# a_20885_45572# 0.002608f
C16595 a_16327_47482# a_20447_31679# 2.78e-20
C16596 a_7411_46660# a_2711_45572# 5.52e-20
C16597 a_3483_46348# a_13759_46122# 6.81e-19
C16598 a_12549_44172# a_17478_45572# 8.8e-20
C16599 a_n1151_42308# a_5691_45260# 1.4e-20
C16600 a_3160_47472# a_3232_43370# 2.79e-20
C16601 a_15227_44166# a_19597_46482# 6.67e-19
C16602 a_4791_45118# a_3537_45260# 0.33264f
C16603 a_6851_47204# a_413_45260# 9.63e-20
C16604 a_n881_46662# a_14127_45572# 7.26e-20
C16605 a_12861_44030# a_n1059_45260# 7.52e-20
C16606 a_4883_46098# a_21363_45546# 2.24e-20
C16607 a_17591_47464# a_3357_43084# 5.7e-19
C16608 a_18479_47436# a_2437_43646# 0.041425f
C16609 a_13661_43548# a_15037_45618# 0.001104f
C16610 a_8016_46348# a_9625_46129# 0.128435f
C16611 a_8199_44636# a_5937_45572# 0.573373f
C16612 a_13747_46662# a_14033_45822# 0.021007f
C16613 a_17339_46660# a_8049_45260# 0.023006f
C16614 a_14180_46812# a_14180_46482# 6.29e-19
C16615 a_21496_47436# a_21188_45572# 1.76e-21
C16616 a_6540_46812# a_6598_45938# 1.76e-21
C16617 a_8270_45546# a_n357_42282# 5.72e-20
C16618 a_n1809_43762# VDD 0.142403f
C16619 a_4190_30871# a_n3420_37984# 0.032285f
C16620 a_18249_42858# a_17303_42282# 4.65e-20
C16621 a_n4318_38216# a_n961_42308# 1.13e-20
C16622 a_14401_32519# VCM 0.007907f
C16623 a_18083_42858# a_18057_42282# 9.91e-19
C16624 a_n1736_42282# a_n4318_37592# 0.153911f
C16625 a_n3674_38216# COMP_P 2.04e-19
C16626 a_n3674_39304# a_n4064_39072# 0.539144f
C16627 a_3080_42308# C0_dummy_N_btm 1.48e-19
C16628 a_n443_42852# a_14635_42282# 4.48e-20
C16629 a_12883_44458# a_11341_43940# 9.36e-21
C16630 a_1423_45028# a_8147_43396# 2e-21
C16631 a_18443_44721# a_18326_43940# 0.007036f
C16632 a_18287_44626# a_18451_43940# 0.005619f
C16633 a_18248_44752# a_19328_44172# 1.49e-20
C16634 a_11967_42832# a_22591_44484# 2.53e-20
C16635 a_20159_44458# a_20512_43084# 9.66e-22
C16636 a_20679_44626# a_20637_44484# 2.56e-19
C16637 a_2107_46812# CLK 3e-20
C16638 a_10775_45002# a_10695_43548# 1.22e-21
C16639 a_13556_45296# a_8685_43396# 6.99e-19
C16640 a_3177_46902# VDD 0.200982f
C16641 a_11827_44484# a_18797_44260# 5.32e-19
C16642 a_n2661_43922# a_7542_44172# 5.03e-21
C16643 a_n2661_42834# a_7845_44172# 0.009718f
C16644 a_6109_44484# a_6756_44260# 2.02e-19
C16645 a_18579_44172# a_19789_44512# 0.003679f
C16646 a_19279_43940# a_3422_30871# 0.02352f
C16647 a_n913_45002# a_19268_43646# 1.96e-21
C16648 a_526_44458# a_8791_42308# 1.73e-21
C16649 a_18989_43940# a_17973_43940# 8.65e-20
C16650 a_1307_43914# a_2813_43396# 6.65e-19
C16651 a_n2293_42834# a_4905_42826# 0.046599f
C16652 a_18184_42460# a_19741_43940# 4.62e-19
C16653 a_2324_44458# a_11823_42460# 0.058835f
C16654 a_6755_46942# a_1307_43914# 0.076439f
C16655 a_8199_44636# a_8697_45572# 4.76e-19
C16656 a_3090_45724# a_5111_44636# 0.063636f
C16657 a_6945_45028# a_8162_45546# 2.68e-20
C16658 a_n2661_46634# a_11691_44458# 8.5e-20
C16659 a_12816_46660# a_6171_45002# 6.34e-21
C16660 a_12741_44636# a_18341_45572# 2.38e-20
C16661 a_11453_44696# a_18287_44626# 0.001467f
C16662 a_13759_46122# a_14495_45572# 2.94e-20
C16663 a_13925_46122# a_13249_42308# 0.001657f
C16664 a_10355_46116# a_10210_45822# 1.86e-19
C16665 a_19321_45002# a_18545_45144# 8.98e-21
C16666 a_20841_46902# a_20731_45938# 1.09e-20
C16667 a_21363_46634# a_21188_45572# 9.99e-20
C16668 a_n1613_43370# a_8701_44490# 2.9e-20
C16669 a_11415_45002# a_19431_45546# 0.005163f
C16670 a_133_42852# VDD 0.184203f
C16671 a_n3674_38216# a_n3565_37414# 3.9e-20
C16672 a_19511_42282# a_19647_42308# 0.038787f
C16673 COMP_P a_8530_39574# 2.33e-19
C16674 a_n4318_37592# a_n4209_37414# 0.105251f
C16675 a_22959_43948# a_14021_43940# 3.06e-19
C16676 a_11827_44484# a_15567_42826# 8.21e-22
C16677 a_18494_42460# a_18083_42858# 0.002227f
C16678 a_18184_42460# a_17333_42852# 1.09e-19
C16679 a_n913_45002# a_1755_42282# 0.169955f
C16680 a_n1059_45260# a_2123_42473# 0.002629f
C16681 a_10405_44172# a_10651_43940# 0.014272f
C16682 a_10729_43914# a_10555_43940# 6.54e-19
C16683 a_7281_43914# a_n97_42460# 4.63e-19
C16684 a_1414_42308# a_4699_43561# 4.09e-21
C16685 a_n356_44636# a_4361_42308# 0.030056f
C16686 a_n2017_45002# a_2351_42308# 0.0062f
C16687 a_19553_46090# VDD 0.204238f
C16688 a_18819_46122# START 8.36e-19
C16689 a_18985_46122# RST_Z 1.22e-21
C16690 a_n2661_44458# a_9127_43156# 6.51e-21
C16691 a_n2293_42834# a_7573_43172# 1.55e-19
C16692 a_742_44458# a_4520_42826# 9.98e-21
C16693 a_2479_44172# a_1756_43548# 1.44e-20
C16694 a_895_43940# a_1568_43370# 3.85e-20
C16695 a_n1644_44306# a_n1699_43638# 2.06e-19
C16696 a_3357_43084# a_3905_42558# 2.81e-19
C16697 a_13249_42308# a_15599_45572# 6.02e-22
C16698 a_13904_45546# a_15903_45785# 8.4e-22
C16699 a_n443_46116# a_1209_43370# 0.061682f
C16700 a_584_46384# a_1987_43646# 2.38e-19
C16701 a_2804_46116# a_n2661_44458# 4.17e-21
C16702 a_11415_45002# a_13076_44458# 3.9e-21
C16703 a_472_46348# a_949_44458# 7.78e-21
C16704 a_12741_44636# a_8975_43940# 3.01e-19
C16705 a_n2312_38680# a_n2661_42282# 4.25e-20
C16706 a_12549_44172# a_20935_43940# 0.110704f
C16707 a_8049_45260# a_1307_43914# 1.63e-19
C16708 a_n2661_45546# a_n467_45028# 0.002796f
C16709 a_n357_42282# a_n2017_45002# 0.580077f
C16710 a_n2293_45546# a_n967_45348# 0.119714f
C16711 a_15227_44166# a_15146_44811# 1.56e-20
C16712 a_n443_42852# a_2437_43646# 0.006604f
C16713 a_13747_46662# a_15682_43940# 3.79e-21
C16714 a_13661_43548# a_17737_43940# 0.031811f
C16715 a_16327_47482# a_18533_43940# 0.001702f
C16716 a_15143_45578# a_15225_45822# 0.004937f
C16717 a_10210_45822# a_10544_45572# 2.43e-19
C16718 a_10907_45822# a_10306_45572# 2.2e-19
C16719 a_10227_46804# a_15037_43940# 0.002378f
C16720 a_n1099_45572# a_n913_45002# 2.98e-19
C16721 a_4185_45028# a_18114_32519# 0.080343f
C16722 a_n1435_47204# a_1983_46706# 5.62e-21
C16723 a_n4209_37414# a_n4334_37440# 0.253282f
C16724 a_13507_46334# a_19594_46812# 0.007313f
C16725 a_20894_47436# a_20916_46384# 4.94e-19
C16726 a_16241_47178# a_n743_46660# 0.001102f
C16727 a_n1151_42308# a_4646_46812# 0.330834f
C16728 a_12465_44636# a_13661_43548# 0.106973f
C16729 a_n4209_38502# C9_P_btm 3.26e-20
C16730 a_n971_45724# a_5257_43370# 0.001362f
C16731 a_2063_45854# a_5167_46660# 6.73e-19
C16732 a_n4315_30879# VIN_P 0.187185f
C16733 a_n2302_39866# VDD 0.361509f
C16734 a_10807_43548# a_12089_42308# 0.002697f
C16735 a_n2293_43922# a_564_42282# 8.6e-20
C16736 a_2982_43646# a_14358_43442# 8.47e-21
C16737 a_18184_42460# a_18997_42308# 2.46e-19
C16738 a_19963_31679# a_22469_39537# 4.14e-20
C16739 a_n356_44636# a_6761_42308# 1.57e-19
C16740 a_n97_42460# a_16409_43396# 0.002137f
C16741 a_6031_43396# a_7221_43396# 2.56e-19
C16742 a_6765_43638# a_6643_43396# 3.16e-19
C16743 a_11967_42832# a_17665_42852# 4.85e-19
C16744 a_n755_45592# a_n310_44484# 0.001049f
C16745 a_413_45260# a_3232_43370# 0.004402f
C16746 a_8016_46348# a_9672_43914# 0.074243f
C16747 a_5937_45572# a_8018_44260# 1.38e-20
C16748 a_8199_44636# a_8333_44056# 2.67e-19
C16749 a_12861_44030# a_19987_42826# 1.24e-19
C16750 a_8162_45546# a_8103_44636# 5.17e-20
C16751 a_3090_45724# a_4235_43370# 1.99e-22
C16752 a_3429_45260# a_3537_45260# 0.138977f
C16753 a_3065_45002# a_4574_45260# 4.96e-19
C16754 a_n1613_43370# a_n1533_42852# 0.012196f
C16755 a_9049_44484# a_5343_44458# 1.3e-20
C16756 a_n2661_45546# a_n2661_43922# 0.028803f
C16757 a_10227_46804# a_15279_43071# 0.001583f
C16758 a_16327_47482# a_17595_43084# 0.007234f
C16759 a_15903_45785# a_17023_45118# 6.24e-21
C16760 a_n2810_45572# a_n2293_43922# 2.93e-20
C16761 a_n881_46662# a_n2472_46090# 1.56e-19
C16762 a_n1613_43370# a_n2293_46098# 0.037934f
C16763 a_11599_46634# a_12005_46116# 0.27095f
C16764 a_584_46384# a_739_46482# 0.004982f
C16765 a_n1151_42308# a_n1545_46494# 4.22e-19
C16766 a_12861_44030# a_13925_46122# 0.012485f
C16767 a_13487_47204# a_13759_46122# 1.3e-19
C16768 a_9313_45822# a_2324_44458# 0.004416f
C16769 a_20843_47204# a_20841_46902# 0.002074f
C16770 a_20916_46384# a_20411_46873# 0.004811f
C16771 a_12891_46348# a_11415_45002# 0.059955f
C16772 a_12549_44172# a_20202_43084# 0.028142f
C16773 a_13661_43548# a_20528_46660# 1.2e-20
C16774 a_8145_46902# a_8035_47026# 0.097745f
C16775 a_7927_46660# a_7832_46660# 0.049827f
C16776 a_n743_46660# a_16721_46634# 0.038286f
C16777 a_n237_47217# a_518_46155# 5.8e-20
C16778 a_10467_46802# a_6755_46942# 0.256039f
C16779 a_10623_46897# a_10249_46116# 0.032312f
C16780 a_4883_46098# a_4704_46090# 0.1774f
C16781 a_n4318_39768# a_n4334_39616# 0.084616f
C16782 a_n3674_39768# a_n4209_39590# 0.044895f
C16783 a_4223_44672# VDD 2.99073f
C16784 a_5649_42852# a_10991_42826# 3.31e-20
C16785 a_19721_31679# VREF 0.057702f
C16786 a_16823_43084# a_16414_43172# 0.024882f
C16787 a_4361_42308# a_12379_42858# 2.98e-19
C16788 a_18114_32519# VREF_GND 0.493553f
C16789 a_11341_43940# a_15890_42674# 3.39e-22
C16790 a_15493_43940# a_15803_42450# 1.43e-21
C16791 a_n2661_44458# CLK 2.88e-19
C16792 a_104_43370# a_n3674_37592# 2.95e-21
C16793 a_n97_42460# a_564_42282# 4.81e-20
C16794 a_743_42282# a_13635_43156# 4.32e-19
C16795 a_15743_43084# a_21356_42826# 0.004418f
C16796 a_15682_43940# a_4958_30871# 2.92e-20
C16797 a_n2661_42282# a_7174_31319# 2.04e-20
C16798 a_4185_45028# a_13887_32519# 0.044689f
C16799 a_10193_42453# a_15493_43940# 0.597095f
C16800 a_n2293_45546# a_n1917_43396# 9.31e-20
C16801 a_n2661_43370# a_6298_44484# 6.23e-19
C16802 a_5205_44484# a_n2661_43922# 0.032439f
C16803 a_8016_46348# a_743_42282# 1.7e-20
C16804 a_13507_46334# a_18057_42282# 6.56e-20
C16805 a_10907_45822# a_10729_43914# 0.00119f
C16806 a_19778_44110# a_19929_45028# 0.001438f
C16807 a_n2840_46090# a_n1853_46287# 2.2e-19
C16808 a_n881_46662# a_6812_45938# 1.43e-19
C16809 a_n743_46660# a_3503_45724# 1.13e-21
C16810 a_13661_43548# a_2711_45572# 0.552383f
C16811 a_6755_46942# a_8034_45724# 4.79e-20
C16812 a_10467_46802# a_8049_45260# 1.3e-20
C16813 a_15227_44166# a_20708_46348# 0.106656f
C16814 a_14513_46634# a_13759_46122# 3.91e-20
C16815 a_14180_46812# a_13925_46122# 4.05e-19
C16816 a_13885_46660# a_14275_46494# 5.27e-19
C16817 a_17609_46634# a_6945_45028# 4.21e-20
C16818 a_15559_46634# a_10809_44734# 0.004011f
C16819 a_14035_46660# a_14493_46090# 2.33e-20
C16820 a_n2472_46090# a_n2157_46122# 0.080495f
C16821 a_765_45546# a_5937_45572# 9.62e-20
C16822 a_12861_44030# a_15599_45572# 0.025507f
C16823 a_n2661_46634# a_n443_42852# 3.69e-19
C16824 a_n2293_46634# a_n1013_45572# 0.001008f
C16825 a_1799_45572# a_n2661_45546# 0.003948f
C16826 a_768_44030# a_3775_45552# 1.42e-21
C16827 a_19466_46812# a_20075_46420# 0.007984f
C16828 a_19692_46634# a_19335_46494# 0.002287f
C16829 a_14955_47212# a_15037_45618# 4.91e-20
C16830 a_3080_42308# VDAC_Ni 6.28e-19
C16831 a_4190_30871# a_19511_42282# 0.005903f
C16832 a_4361_42308# a_18727_42674# 0.006318f
C16833 a_17538_32519# a_22521_40599# 4.64e-21
C16834 a_n2293_42282# a_1067_42314# 1.58e-19
C16835 a_15493_43940# VDD 1.4617f
C16836 a_133_42852# a_n784_42308# 1.2e-19
C16837 a_5649_42852# a_17303_42282# 0.060649f
C16838 a_16823_43084# a_7174_31319# 7.12e-22
C16839 a_8605_42826# a_8791_42308# 0.001071f
C16840 a_8387_43230# a_8685_42308# 1.16e-19
C16841 a_22223_43948# RST_Z 7.78e-20
C16842 a_9313_44734# a_11967_42832# 0.216837f
C16843 a_4223_44672# a_5495_43940# 0.06577f
C16844 a_n2956_39304# a_n4318_38216# 0.023331f
C16845 a_1307_43914# a_15037_43940# 0.004228f
C16846 a_n1699_44726# a_n1644_44306# 3.98e-19
C16847 a_n1177_44458# a_n4318_39768# 1.8e-20
C16848 a_2266_47570# DATA[1] 1.59e-20
C16849 a_22959_47212# EN_OFFSET_CAL 0.007205f
C16850 a_n443_42852# a_14543_43071# 6.35e-20
C16851 a_n357_42282# a_19164_43230# 0.011328f
C16852 a_n2956_38680# a_n2472_42282# 2.5e-20
C16853 a_4185_45028# a_8515_42308# 6.87e-20
C16854 a_11453_44696# CLK 8.57e-19
C16855 a_8696_44636# a_17499_43370# 5.21e-19
C16856 a_17719_45144# a_18079_43940# 2.13e-20
C16857 en_comp a_2982_43646# 0.021697f
C16858 a_13507_46334# a_18494_42460# 0.234442f
C16859 a_19900_46494# a_20062_46116# 0.006453f
C16860 a_4185_45028# a_2711_45572# 0.102913f
C16861 a_4651_46660# a_413_45260# 3.36e-20
C16862 a_11453_44696# a_17023_45118# 1.62e-19
C16863 a_8034_45724# a_8049_45260# 0.141057f
C16864 a_18985_46122# a_21167_46155# 1.63e-20
C16865 a_8199_44636# a_n443_42852# 0.021145f
C16866 a_768_44030# a_5093_45028# 1.51e-19
C16867 a_11415_45002# a_11322_45546# 0.527707f
C16868 a_10428_46928# a_3357_43084# 1.41e-20
C16869 a_3090_45724# a_16147_45260# 0.076341f
C16870 a_n743_46660# a_14180_45002# 7.43e-22
C16871 a_3483_46348# a_4099_45572# 0.15767f
C16872 a_4791_45118# a_8701_44490# 0.138973f
C16873 a_12741_44636# a_10193_42453# 0.078619f
C16874 a_4883_46098# a_19778_44110# 3.83e-22
C16875 a_14209_32519# VIN_N 0.044892f
C16876 a_13575_42558# a_13657_42558# 0.171361f
C16877 a_13070_42354# a_14113_42308# 1.66e-20
C16878 a_n1630_35242# a_n3690_39616# 9.65e-20
C16879 a_n3674_38680# a_n3420_39072# 0.172947f
C16880 a_n3674_39304# VDD 0.587205f
C16881 a_5934_30871# a_4958_30871# 0.018095f
C16882 a_13887_32519# VREF_GND 0.047292f
C16883 a_19279_43940# a_19808_44306# 0.002998f
C16884 a_16922_45042# a_20749_43396# 0.106779f
C16885 a_5891_43370# a_6547_43396# 6.62e-20
C16886 a_n2293_42834# a_2905_42968# 0.010834f
C16887 a_10193_42453# a_5742_30871# 0.303452f
C16888 a_11967_42832# a_20974_43370# 2.01e-20
C16889 a_12741_44636# VDD 0.988199f
C16890 a_n2293_43922# a_n1557_42282# 2.21e-19
C16891 a_21076_30879# C10_N_btm 9.75e-19
C16892 a_20820_30879# RST_Z 0.048737f
C16893 a_18184_42460# a_13678_32519# 0.019189f
C16894 a_14539_43914# a_14358_43442# 2.26e-19
C16895 a_15004_44636# a_15095_43370# 9.09e-22
C16896 a_10057_43914# a_12293_43646# 3.63e-20
C16897 a_n2810_45572# a_n3420_39616# 1.68e-19
C16898 a_n1059_45260# a_8495_42852# 0.00552f
C16899 a_13351_46090# a_13017_45260# 1.33e-20
C16900 a_12594_46348# a_13159_45002# 2.01e-20
C16901 a_8953_45546# a_1307_43914# 0.022061f
C16902 a_6945_45028# a_3537_45260# 9.87e-21
C16903 a_16375_45002# a_18341_45572# 9.37e-19
C16904 a_n1925_42282# a_n913_45002# 0.017956f
C16905 a_8049_45260# a_20885_45572# 3.49e-19
C16906 a_584_46384# a_1241_43940# 0.007526f
C16907 a_10903_43370# a_9482_43914# 1.20611f
C16908 a_2711_45572# a_6229_45572# 4.93e-19
C16909 a_6419_46155# a_1423_45028# 3.69e-22
C16910 a_2324_44458# a_7705_45326# 0.029419f
C16911 a_167_45260# a_117_45144# 0.003885f
C16912 a_11415_45002# a_15060_45348# 0.001314f
C16913 a_9290_44172# a_14537_43396# 3.99e-19
C16914 a_1823_45246# a_2809_45028# 0.076288f
C16915 a_13747_46662# a_20512_43084# 5.53e-21
C16916 a_4958_30871# a_11530_34132# 0.020719f
C16917 a_15673_47210# a_13507_46334# 0.001528f
C16918 a_15507_47210# a_4883_46098# 4.76e-22
C16919 a_5934_30871# VCM 0.121361f
C16920 a_13717_47436# a_11453_44696# 0.041574f
C16921 a_17591_47464# a_18597_46090# 8.92e-19
C16922 a_n3565_38216# a_n4064_37984# 0.342209f
C16923 a_n4209_38216# a_n4251_38304# 0.00226f
C16924 a_5742_30871# VDD 0.556959f
C16925 a_14955_47212# a_12465_44636# 0.002323f
C16926 a_4791_45118# a_n1613_43370# 0.223884f
C16927 a_18143_47464# a_18479_47436# 0.238309f
C16928 a_10227_46804# a_18780_47178# 0.050298f
C16929 a_n1151_42308# a_9804_47204# 0.108722f
C16930 a_584_46384# a_768_44030# 0.105366f
C16931 a_n971_45724# a_5807_45002# 0.0339f
C16932 a_22465_38105# a_22521_40599# 0.132396f
C16933 a_1209_43370# a_1049_43396# 0.194938f
C16934 a_n97_42460# a_n1557_42282# 0.149645f
C16935 a_458_43396# a_1568_43370# 2.29e-20
C16936 a_11341_43940# a_16547_43609# 2.97e-19
C16937 a_15493_43940# a_16137_43396# 0.043956f
C16938 a_n1644_44306# a_n2157_42858# 2.8e-20
C16939 a_n2956_37592# a_n2216_39072# 1.2e-19
C16940 a_19328_44172# a_15743_43084# 2.2e-21
C16941 a_15493_43396# a_18783_43370# 0.029898f
C16942 a_453_43940# a_791_42968# 1.04e-20
C16943 a_11967_42832# a_18599_43230# 0.003648f
C16944 a_n699_43396# a_196_42282# 0.001148f
C16945 a_1414_42308# a_1847_42826# 7.16e-21
C16946 a_4185_45028# a_22485_44484# 0.080982f
C16947 a_21513_45002# a_22223_45572# 5.7e-19
C16948 a_19692_46634# a_22959_43948# 8.6e-20
C16949 a_2711_45572# a_18587_45118# 7.13e-22
C16950 a_n2293_45546# a_n1917_44484# 6.29e-19
C16951 a_n2293_46634# a_8791_43396# 0.010288f
C16952 a_526_44458# a_3363_44484# 0.119556f
C16953 a_17715_44484# a_17517_44484# 0.163303f
C16954 a_2324_44458# a_15367_44484# 3.72e-19
C16955 a_16327_47482# a_13467_32519# 0.004353f
C16956 a_13059_46348# a_13483_43940# 0.124566f
C16957 a_20719_45572# a_3357_43084# 2.25e-19
C16958 a_13259_45724# a_13076_44458# 0.188498f
C16959 a_n1099_45572# a_n2661_44458# 9.19e-21
C16960 a_12549_44172# a_14955_43396# 4.21e-19
C16961 a_19120_35138# VIN_N 0.001664f
C16962 a_n1925_46634# a_8492_46660# 9.51e-19
C16963 a_5807_45002# a_8023_46660# 0.001248f
C16964 a_12549_44172# a_12469_46902# 0.00102f
C16965 a_12891_46348# a_12251_46660# 0.003575f
C16966 a_4791_45118# a_n2293_46098# 0.411939f
C16967 a_11453_44696# a_14035_46660# 1.53e-20
C16968 a_13507_46334# a_16388_46812# 0.083261f
C16969 a_18143_47464# a_17829_46910# 2.74e-19
C16970 a_18479_47436# a_765_45546# 1.7e-19
C16971 a_10227_46804# a_18285_46348# 5.46e-20
C16972 a_3177_46902# a_4646_46812# 2.63e-20
C16973 a_2609_46660# a_4651_46660# 1.13e-19
C16974 a_2959_46660# a_3877_44458# 2.53e-19
C16975 a_2107_46812# a_3878_46660# 3.62e-19
C16976 a_n2109_47186# a_5497_46414# 0.017063f
C16977 a_n1741_47186# a_5164_46348# 3.78e-20
C16978 a_n2661_46634# a_10554_47026# 0.009556f
C16979 a_584_46384# a_1176_45822# 0.039976f
C16980 a_n1151_42308# a_n901_46420# 0.002158f
C16981 a_2063_45854# a_1208_46090# 4.06e-19
C16982 EN_VIN_BSTR_N VREF_GND 0.85739f
C16983 a_12861_44030# a_16655_46660# 6.9e-19
C16984 a_n881_46662# a_15559_46634# 3.94e-20
C16985 a_1209_47178# a_167_45260# 2.76e-21
C16986 a_n971_45724# a_3699_46348# 0.013334f
C16987 a_n237_47217# a_3147_46376# 0.052931f
C16988 a_2443_46660# a_4955_46873# 4.31e-21
C16989 C2_N_btm C8_N_btm 0.14124f
C16990 C1_N_btm C9_N_btm 0.133953f
C16991 C0_N_btm C10_N_btm 0.251079f
C16992 C4_N_btm C6_N_btm 0.145942f
C16993 C3_N_btm C7_N_btm 0.136068f
C16994 a_n2293_42834# VDD 0.853754f
C16995 a_21259_43561# a_4190_30871# 0.198353f
C16996 a_8685_43396# a_10991_42826# 1.51e-19
C16997 a_18114_32519# a_22469_40625# 9.95e-21
C16998 a_19721_31679# a_22521_40599# 1.69e-20
C16999 a_n2661_42282# a_5932_42308# 0.070536f
C17000 a_18579_44172# a_13258_32519# 3.63e-20
C17001 a_3422_30871# a_19332_42282# 6.32e-20
C17002 a_9145_43396# a_9127_43156# 0.001269f
C17003 a_5111_44636# a_4743_44484# 0.02485f
C17004 a_5147_45002# a_5343_44458# 0.063193f
C17005 a_3537_45260# a_8103_44636# 0.140404f
C17006 a_n357_42282# a_18079_43940# 1.54e-20
C17007 a_n2661_45010# a_n1809_44850# 0.006483f
C17008 a_3232_43370# a_2779_44458# 0.003663f
C17009 a_4880_45572# a_3905_42865# 1.35e-19
C17010 a_15861_45028# a_17517_44484# 0.003385f
C17011 a_8696_44636# a_18204_44850# 7.09e-21
C17012 a_10951_45334# a_n2661_44458# 2.65e-20
C17013 a_n1613_43370# a_n1736_42282# 1.08e-20
C17014 a_16751_45260# a_11691_44458# 1.98e-19
C17015 a_16019_45002# a_16237_45028# 0.053167f
C17016 a_7418_45067# a_n2661_43370# 4e-19
C17017 a_8953_45546# a_9396_43370# 0.007396f
C17018 a_8270_45546# a_8952_43230# 1.53e-20
C17019 a_12741_44636# a_16137_43396# 3.03e-20
C17020 a_2107_46812# a_n1925_42282# 0.006094f
C17021 a_5807_45002# a_12005_46436# 8.93e-20
C17022 a_12891_46348# a_13259_45724# 1.04614f
C17023 a_2063_45854# a_11525_45546# 0.001514f
C17024 a_6755_46942# a_8016_46348# 0.002347f
C17025 a_4791_45118# a_7230_45938# 0.010716f
C17026 a_6151_47436# a_4808_45572# 2.53e-20
C17027 a_2747_46873# a_n2661_45546# 1.72e-21
C17028 a_765_45546# a_17829_46910# 0.069261f
C17029 a_17339_46660# a_18285_46348# 0.184197f
C17030 a_n1151_42308# a_10180_45724# 6.68e-20
C17031 a_9863_46634# a_9823_46155# 9.52e-19
C17032 a_n2661_46098# a_n722_46482# 0.001878f
C17033 a_14955_47212# a_2711_45572# 1.19e-21
C17034 a_n1076_43230# a_n3674_37592# 4.57e-20
C17035 a_n2293_42282# a_4149_42891# 1.94e-19
C17036 a_1115_44172# VDD 0.165092f
C17037 a_4361_42308# a_3823_42558# 0.114877f
C17038 a_n13_43084# a_n327_42558# 2.86e-20
C17039 a_17730_32519# VIN_N 0.048461f
C17040 a_10341_43396# a_15890_42674# 7.05e-21
C17041 a_14543_43071# a_14635_42282# 0.075815f
C17042 a_5534_30871# a_13291_42460# 0.045073f
C17043 a_n1641_43230# a_n1630_35242# 6.83e-20
C17044 a_743_42282# a_3905_42558# 0.003412f
C17045 a_3160_47472# VDD 0.256092f
C17046 a_n356_44636# a_5891_43370# 4.5e-19
C17047 a_13556_45296# a_13483_43940# 0.001149f
C17048 a_9482_43914# a_14955_43940# 6.17e-19
C17049 a_18114_32519# a_11967_42832# 0.002218f
C17050 a_n2661_43370# a_2479_44172# 4.26e-20
C17051 a_9290_44172# a_12991_43230# 1.31e-20
C17052 a_7499_43078# a_8945_43396# 2.24e-19
C17053 a_6171_45002# a_11341_43940# 5.17e-20
C17054 a_3090_45724# a_15051_42282# 1.14e-20
C17055 a_584_46384# DATA[0] 3.21e-20
C17056 a_2124_47436# DATA[1] 0.00138f
C17057 a_20193_45348# a_18579_44172# 2.14e-20
C17058 a_11691_44458# a_18681_44484# 0.002372f
C17059 a_12883_44458# a_n2293_43922# 0.06281f
C17060 a_18989_43940# a_9313_44734# 1.23e-19
C17061 a_12607_44458# a_13213_44734# 1.94e-19
C17062 a_n2293_42834# a_5495_43940# 1.87e-21
C17063 a_1307_43914# a_9028_43914# 0.010468f
C17064 a_21359_45002# a_21398_44850# 0.001485f
C17065 a_11827_44484# a_20980_44850# 0.002088f
C17066 a_11823_42460# a_14579_43548# 0.106967f
C17067 a_11453_44696# a_10951_45334# 5.15e-19
C17068 a_11813_46116# a_11962_45724# 1.15e-19
C17069 a_22959_46660# a_20692_30879# 0.004672f
C17070 a_n881_46662# a_3065_45002# 1.23e-20
C17071 a_n1613_43370# a_3429_45260# 2.46e-21
C17072 a_12465_44636# a_13159_45002# 6.58e-20
C17073 a_21137_46414# a_10809_44734# 1.12e-20
C17074 a_6945_45028# a_22223_46124# 0.17119f
C17075 a_8016_46348# a_8049_45260# 0.09608f
C17076 a_8953_45546# a_8034_45724# 2.24e-19
C17077 a_765_45546# a_n443_42852# 0.232932f
C17078 a_21076_30879# a_20205_31679# 0.055235f
C17079 a_n2661_46634# a_2437_43646# 0.02989f
C17080 a_4883_46098# a_9482_43914# 0.025151f
C17081 a_2903_42308# a_6123_31319# 2.22e-20
C17082 a_1606_42308# a_8685_42308# 1.35e-20
C17083 a_n784_42308# a_5742_30871# 0.550812f
C17084 a_16245_42852# a_4958_30871# 6.84e-19
C17085 a_10849_43646# VDD 0.009276f
C17086 a_9145_43396# CLK 2.67e-21
C17087 a_11967_42832# a_17737_43940# 0.054562f
C17088 a_n2065_43946# a_n1453_44318# 0.001881f
C17089 a_413_45260# a_2905_42968# 1.46e-20
C17090 a_n1059_45260# a_9127_43156# 0.006366f
C17091 a_n913_45002# a_8387_43230# 0.024148f
C17092 a_n2017_45002# a_8952_43230# 4.34e-20
C17093 a_n443_42852# a_4921_42308# 4.12e-19
C17094 a_5891_43370# a_9165_43940# 8.35e-19
C17095 a_742_44458# a_n1557_42282# 6.13e-20
C17096 a_13607_46688# VDD 0.209568f
C17097 a_2479_44172# a_2998_44172# 0.004129f
C17098 a_n1761_44111# a_n1644_44306# 0.170098f
C17099 a_n1899_43946# a_n3674_39768# 4.83e-19
C17100 a_4223_44672# a_3080_42308# 2.46e-19
C17101 a_n699_43396# a_4699_43561# 6.51e-20
C17102 a_n2661_42834# a_726_44056# 6.09e-19
C17103 a_14673_44172# a_11341_43940# 0.001734f
C17104 a_n755_45592# a_3905_42308# 6.37e-19
C17105 a_10384_47026# CLK 9.6e-20
C17106 a_12465_44636# a_11967_42832# 1.63e-20
C17107 a_4883_46098# a_20159_44458# 4.39e-22
C17108 a_3877_44458# a_n699_43396# 0.061672f
C17109 a_4646_46812# a_4223_44672# 0.018453f
C17110 a_8049_45260# a_11682_45822# 0.011453f
C17111 a_12839_46116# a_11823_42460# 2.9e-19
C17112 a_12891_46348# a_n2661_43922# 1.94e-19
C17113 a_12549_44172# a_n2661_42834# 0.04571f
C17114 a_n746_45260# a_261_44278# 5.72e-19
C17115 a_n2497_47436# a_n2661_42282# 4.56e-21
C17116 a_n971_45724# a_n822_43940# 1.37e-19
C17117 a_8199_44636# a_2437_43646# 3.38e-20
C17118 a_13507_46334# a_20640_44752# 8.68e-20
C17119 a_13259_45724# a_11322_45546# 5.48e-21
C17120 a_n2661_45546# a_3638_45822# 2.27e-21
C17121 a_5807_45002# a_9313_44734# 7.63e-20
C17122 a_18985_46122# a_18341_45572# 7.1e-19
C17123 a_18819_46122# a_18909_45814# 0.003441f
C17124 a_19335_46494# a_18175_45572# 1.2e-19
C17125 a_n2293_46098# a_3429_45260# 2.13e-20
C17126 a_11453_44696# a_17061_44484# 3.88e-19
C17127 a_n443_46116# a_895_43940# 0.163929f
C17128 a_16375_45002# a_10193_42453# 0.125364f
C17129 a_509_45822# a_n443_42852# 0.035689f
C17130 a_n755_45592# a_3175_45822# 0.046968f
C17131 a_n785_47204# a_n1435_47204# 9.32e-19
C17132 a_4700_47436# a_n443_46116# 0.255594f
C17133 a_n1151_42308# a_6545_47178# 0.01616f
C17134 a_2063_45854# a_6575_47204# 0.002711f
C17135 a_3785_47178# a_5815_47464# 2.66e-19
C17136 a_4007_47204# a_4915_47217# 0.001046f
C17137 a_n4064_39616# a_n4064_39072# 0.062881f
C17138 a_n3420_39616# a_n4251_39392# 8.88e-19
C17139 a_n4064_40160# a_n4209_38502# 0.05515f
C17140 a_1606_42308# C10_P_btm 1.34e-19
C17141 a_n4315_30879# a_n3565_38502# 0.085594f
C17142 a_22765_42852# VDD 0.006527f
C17143 a_n784_42308# C0_dummy_P_btm 2.62e-20
C17144 a_4958_30871# a_7754_40130# 5.49e-20
C17145 a_20679_44626# a_4361_42308# 2.91e-20
C17146 a_9313_44734# a_10518_42984# 0.008938f
C17147 a_n1059_45260# a_17124_42282# 0.008817f
C17148 a_16375_45002# VDD 1.14948f
C17149 a_18989_43940# a_18599_43230# 5.3e-19
C17150 a_n356_44636# a_17595_43084# 2.73e-20
C17151 a_9028_43914# a_9396_43370# 3.1e-19
C17152 a_15493_43396# a_3626_43646# 2.49e-20
C17153 a_19862_44208# a_2982_43646# 0.005666f
C17154 a_n2293_42834# a_n784_42308# 8.13e-19
C17155 a_1307_43914# a_5421_42558# 4.2e-20
C17156 a_18579_44172# a_20301_43646# 3.55e-20
C17157 a_n2661_42834# a_5111_42852# 5.01e-22
C17158 a_n2293_43922# a_3935_42891# 1.63e-22
C17159 a_2711_45572# a_13159_45002# 9.08e-19
C17160 a_n2293_45546# a_2809_45028# 5.9e-20
C17161 a_n1925_42282# a_n2661_44458# 0.029506f
C17162 a_7227_45028# a_7229_43940# 0.019397f
C17163 a_6598_45938# a_6709_45028# 3.05e-21
C17164 a_13259_45724# a_15060_45348# 4.35e-19
C17165 a_13249_42308# a_n2017_45002# 0.030327f
C17166 a_3090_45724# a_3905_42865# 0.025179f
C17167 a_4880_45572# a_5147_45002# 3.65e-19
C17168 a_6419_46155# a_6109_44484# 1.19e-21
C17169 a_9290_44172# a_n356_44636# 8.05e-19
C17170 a_n863_45724# a_117_45144# 2.14e-19
C17171 a_2324_44458# a_14539_43914# 0.028976f
C17172 a_15682_46116# a_16112_44458# 2.03e-21
C17173 a_13747_46662# a_21381_43940# 0.030122f
C17174 a_n2293_46634# a_10651_43940# 6.07e-19
C17175 a_n2840_46634# a_n2442_46660# 0.007415f
C17176 a_n2956_39768# a_n2472_46634# 5e-19
C17177 a_4915_47217# a_15368_46634# 4.4e-21
C17178 a_n1613_43370# a_1057_46660# 2.95e-19
C17179 a_7754_38636# VDD 0.036155f
C17180 a_4883_46098# a_7715_46873# 0.01159f
C17181 a_6151_47436# a_15009_46634# 0.00896f
C17182 a_22609_38406# a_22705_38406# 0.090011f
C17183 CAL_P a_22609_37990# 0.205305f
C17184 a_22469_39537# a_22717_36887# 0.003149f
C17185 a_10227_46804# a_10249_46116# 0.137273f
C17186 a_n1761_44111# a_961_42354# 1.47e-22
C17187 a_1414_42308# a_n473_42460# 2.2e-21
C17188 a_413_45260# VDD 1.203f
C17189 a_10341_43396# a_16547_43609# 0.026476f
C17190 a_12281_43396# a_13837_43396# 7.31e-21
C17191 a_n97_42460# a_3935_42891# 5.1e-20
C17192 a_13565_43940# a_13460_43230# 6.29e-20
C17193 a_n1557_42282# a_n901_43156# 2.27e-19
C17194 a_8791_43396# a_743_42282# 2.77e-21
C17195 a_n809_44244# a_n1630_35242# 5.42e-21
C17196 a_8685_43396# a_15231_43396# 0.002861f
C17197 a_6031_43396# a_5649_42852# 4.06e-21
C17198 a_n1151_42308# a_196_42282# 1.47e-19
C17199 a_9290_44172# a_9165_43940# 0.01396f
C17200 a_11652_45724# a_11649_44734# 1.66e-19
C17201 a_n863_45724# a_n2065_43946# 4.6e-21
C17202 a_n913_45002# a_16922_45042# 6.18e-19
C17203 a_10227_46804# a_15785_43172# 4.06e-19
C17204 a_n971_45724# a_n327_42308# 0.001391f
C17205 a_584_46384# a_1067_42314# 4.65e-21
C17206 a_11525_45546# a_n2661_42834# 5.55e-21
C17207 a_11322_45546# a_n2661_43922# 0.001721f
C17208 a_n2661_45546# a_n809_44244# 2.15e-20
C17209 a_16327_47482# a_18695_43230# 0.003378f
C17210 a_3357_43084# a_11827_44484# 8.78e-20
C17211 a_19479_31679# a_22223_45036# 0.01502f
C17212 a_n2293_45546# a_n1899_43946# 2.4e-20
C17213 a_2680_45002# a_n2661_43370# 0.006576f
C17214 a_6171_45002# a_7418_45394# 1.2e-19
C17215 a_2711_45572# a_11967_42832# 0.068241f
C17216 a_8696_44636# a_15004_44636# 0.003323f
C17217 a_16855_45546# a_14539_43914# 8.46e-20
C17218 a_4185_45028# a_14401_32519# 0.040395f
C17219 a_2324_44458# a_2253_43940# 2.21e-19
C17220 a_10809_44734# a_10555_44260# 6.94e-19
C17221 a_n743_46660# a_5164_46348# 0.031878f
C17222 a_12549_44172# a_17715_44484# 0.03426f
C17223 a_n2661_46098# a_472_46348# 0.065456f
C17224 a_6755_46942# a_15312_46660# 2.66e-21
C17225 a_n1613_43370# a_6945_45028# 0.049203f
C17226 a_5807_45002# a_12594_46348# 0.001952f
C17227 a_n746_45260# a_n357_42282# 0.002027f
C17228 a_n971_45724# a_n755_45592# 0.347347f
C17229 a_n1925_46634# a_5497_46414# 6.78e-20
C17230 a_2063_45854# a_n2661_45546# 0.038547f
C17231 a_12861_44030# a_12638_46436# 6.45e-19
C17232 a_12251_46660# a_12359_47026# 0.057222f
C17233 a_11735_46660# a_12347_46660# 3.82e-19
C17234 a_14976_45028# a_15227_44166# 0.035507f
C17235 a_4883_46098# a_5210_46482# 2.25e-19
C17236 a_17591_47464# a_8049_45260# 1.43e-20
C17237 a_n2661_46634# a_8199_44636# 2.29e-19
C17238 a_2107_46812# a_2698_46116# 0.00811f
C17239 a_13747_46662# a_10903_43370# 0.027209f
C17240 a_n97_42460# a_15890_42674# 0.022679f
C17241 a_13460_43230# a_5534_30871# 0.052631f
C17242 a_6197_43396# a_7227_42308# 1.57e-20
C17243 a_3626_43646# a_8791_42308# 0.003196f
C17244 a_2982_43646# a_9803_42558# 1.36e-19
C17245 a_3080_42308# a_5742_30871# 0.097222f
C17246 a_13468_44734# VDD 0.004018f
C17247 a_791_42968# a_945_42968# 0.008535f
C17248 a_16823_43084# a_17141_43172# 1.56e-19
C17249 a_18783_43370# a_18707_42852# 1.34e-19
C17250 a_15743_43084# a_19518_43218# 0.00221f
C17251 a_9290_44172# a_12379_42858# 0.001587f
C17252 a_4185_45028# a_18817_42826# 1.72e-20
C17253 a_8103_44636# a_8701_44490# 5.82e-19
C17254 a_6298_44484# a_5883_43914# 0.003333f
C17255 a_n443_42852# a_6452_43396# 0.001812f
C17256 a_3065_45002# a_2889_44172# 1.06e-19
C17257 a_2382_45260# a_3600_43914# 0.158274f
C17258 a_2680_45002# a_2998_44172# 1.29e-20
C17259 a_n2661_45010# a_1525_44260# 5.65e-20
C17260 a_n2293_45010# a_n822_43940# 4.54e-19
C17261 a_n913_45002# a_n875_44318# 5.75e-19
C17262 a_10903_43370# a_10796_42968# 0.001425f
C17263 en_comp a_n3674_39768# 0.036087f
C17264 a_13259_45724# a_16409_43396# 7.07e-20
C17265 a_18479_45785# a_15493_43940# 0.016583f
C17266 a_n755_45592# a_8229_43396# 0.002439f
C17267 a_18597_46090# a_20719_45572# 0.005294f
C17268 a_5257_43370# a_2711_45572# 0.082068f
C17269 a_12549_44172# a_15861_45028# 7.24e-20
C17270 a_768_44030# a_8696_44636# 0.031444f
C17271 a_6491_46660# a_413_45260# 3.19e-19
C17272 a_n881_46662# a_14033_45572# 5.52e-20
C17273 a_12861_44030# a_n2017_45002# 6.5e-19
C17274 a_4883_46098# a_20623_45572# 2.03e-20
C17275 a_16588_47582# a_3357_43084# 1.09e-19
C17276 a_16327_47482# a_22959_45572# 5.96e-20
C17277 a_18479_47436# a_21513_45002# 4.09e-20
C17278 a_1823_45246# a_2324_44458# 0.069409f
C17279 a_3483_46348# a_13351_46090# 1.87e-20
C17280 a_5807_45002# a_15037_45618# 4.32e-21
C17281 a_8016_46348# a_8953_45546# 0.060003f
C17282 a_8349_46414# a_5937_45572# 6.5e-20
C17283 a_2063_45854# a_5205_44484# 1.89e-20
C17284 a_14035_46660# a_14180_46482# 0.157972f
C17285 a_n443_46116# a_3065_45002# 1.4e-20
C17286 a_4791_45118# a_3429_45260# 6.17e-21
C17287 a_21496_47436# a_21363_45546# 4.09e-21
C17288 a_13507_46334# a_21188_45572# 8.13e-19
C17289 a_18143_47464# a_2437_43646# 0.013364f
C17290 a_n1151_42308# a_4927_45028# 9.34e-21
C17291 a_19466_46812# a_19431_46494# 0.001367f
C17292 a_19692_46634# a_19240_46482# 4.58e-21
C17293 a_6540_46812# a_6667_45809# 2.06e-20
C17294 a_n4318_38680# a_n3420_39072# 0.310238f
C17295 a_n3674_39304# a_n2946_39072# 4.03e-21
C17296 a_n4318_38216# a_n1329_42308# 2.61e-20
C17297 a_n2104_42282# COMP_P 3.78e-19
C17298 a_17538_32519# VIN_N 0.041176f
C17299 a_n2012_43396# VDD 0.08228f
C17300 a_17333_42852# a_17303_42282# 5.44e-19
C17301 a_14401_32519# VREF_GND 0.066097f
C17302 a_17701_42308# a_18057_42282# 4e-19
C17303 a_3080_42308# C0_dummy_P_btm 1.48e-19
C17304 a_n3674_38216# a_n4318_37592# 2.7294f
C17305 a_n443_42852# a_13291_42460# 1.19e-21
C17306 a_12607_44458# a_11341_43940# 8.67e-21
C17307 a_17767_44458# a_15493_43396# 2.64e-21
C17308 a_18287_44626# a_18326_43940# 0.001026f
C17309 a_18248_44752# a_18451_43940# 5.78e-19
C17310 a_20640_44752# a_20637_44484# 2.36e-20
C17311 a_n2017_45002# a_19700_43370# 4.64e-20
C17312 a_9482_43914# a_8685_43396# 3.32e-20
C17313 a_5883_43914# a_10555_44260# 2.18e-20
C17314 a_2609_46660# VDD 0.312974f
C17315 a_11827_44484# a_18533_44260# 3.57e-19
C17316 a_n2661_43922# a_7281_43914# 1.21e-20
C17317 a_n2661_42834# a_7542_44172# 0.019328f
C17318 a_6109_44484# a_n2661_42282# 0.003425f
C17319 a_11967_42832# a_22485_44484# 3.29e-19
C17320 a_19279_43940# a_21398_44850# 0.183186f
C17321 a_20766_44850# a_3422_30871# 6.2e-20
C17322 a_n913_45002# a_15743_43084# 2.14e-19
C17323 a_526_44458# a_8685_42308# 6.82e-21
C17324 a_1307_43914# a_2437_43396# 2.02e-19
C17325 a_n2293_42834# a_3080_42308# 0.021566f
C17326 a_19778_44110# a_19741_43940# 0.054731f
C17327 a_6171_45002# a_10341_43396# 2.27e-20
C17328 a_n357_42282# a_17749_42852# 0.001128f
C17329 a_2324_44458# a_12427_45724# 0.001185f
C17330 a_14840_46494# a_11823_42460# 0.004799f
C17331 a_6755_46942# a_16019_45002# 0.005906f
C17332 a_4646_46812# a_n2293_42834# 0.152973f
C17333 a_8199_44636# a_8192_45572# 0.04905f
C17334 a_n881_46662# a_6298_44484# 0.002351f
C17335 a_3090_45724# a_5147_45002# 0.023629f
C17336 a_765_45546# a_2437_43646# 0.030322f
C17337 a_526_44458# a_6194_45824# 7.16e-21
C17338 a_6945_45028# a_7230_45938# 5.3e-19
C17339 a_12741_44636# a_18479_45785# 0.035678f
C17340 a_11453_44696# a_18248_44752# 0.004115f
C17341 a_13759_46122# a_13249_42308# 0.001706f
C17342 a_13925_46122# a_13904_45546# 5.43e-19
C17343 a_20528_46660# a_20273_45572# 9.08e-22
C17344 a_21363_46634# a_21363_45546# 0.001846f
C17345 a_11415_45002# a_18691_45572# 0.002376f
C17346 a_n2293_46634# a_11827_44484# 0.002225f
C17347 a_9823_46155# a_10210_45822# 0.001193f
C17348 a_n914_42852# VDD 7.75e-19
C17349 a_19332_42282# a_7174_31319# 7.74e-19
C17350 a_n3674_38216# a_n4334_37440# 6.7e-20
C17351 a_5934_30871# a_n4064_38528# 0.004208f
C17352 COMP_P a_7754_38470# 1.8e-19
C17353 a_2779_44458# a_2905_42968# 2.56e-20
C17354 a_742_44458# a_3935_42891# 1.81e-19
C17355 a_15493_43940# a_14021_43940# 0.08284f
C17356 a_11827_44484# a_5342_30871# 2.98e-20
C17357 a_18184_42460# a_18083_42858# 0.003624f
C17358 a_18494_42460# a_17701_42308# 4.02e-20
C17359 a_14673_44172# a_10341_43396# 1.61e-19
C17360 a_n1059_45260# a_1755_42282# 0.004197f
C17361 a_n913_45002# a_1606_42308# 0.025848f
C17362 a_n2017_45002# a_2123_42473# 0.0078f
C17363 a_10405_44172# a_10555_43940# 0.018661f
C17364 a_10729_43914# a_9801_43940# 7.39e-20
C17365 a_n984_44318# a_n1557_42282# 2.08e-21
C17366 a_1414_42308# a_4235_43370# 1.4e-19
C17367 a_16922_45042# a_20922_43172# 1.86e-19
C17368 a_18985_46122# VDD 0.253642f
C17369 a_18819_46122# RST_Z 7.83e-21
C17370 a_13925_46122# CLK 1.2e-20
C17371 a_n699_43396# a_1847_42826# 5.48e-20
C17372 a_n2293_42834# a_7309_43172# 5.7e-19
C17373 a_2479_44172# a_1568_43370# 0.001043f
C17374 a_11823_42460# a_16115_45572# 9.08e-20
C17375 a_11652_45724# a_8696_44636# 3.56e-19
C17376 a_584_46384# a_1891_43646# 4.57e-19
C17377 a_n443_46116# a_458_43396# 1.87e-21
C17378 a_2698_46116# a_n2661_44458# 1.03e-21
C17379 a_n452_45724# a_n745_45366# 0.00143f
C17380 a_12549_44172# a_20623_43914# 0.033887f
C17381 a_8049_45260# a_16019_45002# 2.24e-21
C17382 a_n755_45592# a_n2293_45010# 0.159033f
C17383 a_15227_44166# a_15433_44458# 0.026124f
C17384 a_n2293_45546# en_comp 2.1e-19
C17385 a_13661_43548# a_15682_43940# 0.055235f
C17386 a_16327_47482# a_19319_43548# 0.021453f
C17387 a_10227_46804# a_13565_43940# 5.26e-19
C17388 a_n1099_45572# a_n1059_45260# 2.72e-19
C17389 a_10907_45822# a_10216_45572# 1.14e-19
C17390 a_15143_45578# a_15037_45618# 0.13675f
C17391 a_n1435_47204# a_2107_46812# 5.14e-20
C17392 a_n4209_38502# C10_P_btm 2.25e-20
C17393 a_7754_39300# a_5700_37509# 2.64e-19
C17394 a_20990_47178# a_20843_47204# 0.003683f
C17395 a_13507_46334# a_19321_45002# 0.034054f
C17396 a_21177_47436# a_19594_46812# 4.79e-20
C17397 a_n1151_42308# a_3877_44458# 0.019733f
C17398 a_3160_47472# a_4646_46812# 2.88e-21
C17399 a_n443_46116# a_3067_47026# 0.030121f
C17400 a_12465_44636# a_5807_45002# 0.59474f
C17401 a_n4064_39072# C0_P_btm 8.17e-21
C17402 a_15673_47210# a_n743_46660# 0.002403f
C17403 a_4883_46098# a_13747_46662# 0.050962f
C17404 a_n4064_39616# VDD 1.6861f
C17405 a_n2293_43922# a_n3674_37592# 0.062473f
C17406 a_2982_43646# a_14579_43548# 5.95e-20
C17407 a_10057_43914# a_5742_30871# 3.08e-19
C17408 a_n97_42460# a_16547_43609# 0.066612f
C17409 a_n2661_42834# a_n1630_35242# 1.36e-19
C17410 a_20447_31679# a_22521_39511# 3.7e-20
C17411 a_6197_43396# a_6643_43396# 2.28e-19
C17412 a_6765_43638# a_7274_43762# 2.6e-19
C17413 a_11967_42832# a_16877_42852# 0.005423f
C17414 a_6031_43396# a_8685_43396# 9.68e-21
C17415 a_5937_45572# a_7911_44260# 2.23e-20
C17416 a_12861_44030# a_19164_43230# 5.09e-21
C17417 a_3090_45724# a_4093_43548# 0.00131f
C17418 a_15861_45028# a_15685_45394# 8.17e-20
C17419 a_3065_45002# a_3537_45260# 0.162384f
C17420 a_n1613_43370# a_n722_43218# 0.00237f
C17421 a_12741_44636# a_14021_43940# 2.11e-19
C17422 a_2711_45572# a_18989_43940# 0.006251f
C17423 a_10227_46804# a_5534_30871# 0.304847f
C17424 a_16327_47482# a_16795_42852# 6.73e-19
C17425 a_15903_45785# a_16922_45042# 5.01e-20
C17426 a_n2661_45546# a_n2661_42834# 0.029567f
C17427 a_7499_43078# a_5343_44458# 0.050528f
C17428 a_10623_46897# a_10554_47026# 0.209641f
C17429 a_10428_46928# a_6755_46942# 0.155315f
C17430 a_10467_46802# a_10249_46116# 0.12624f
C17431 a_n1613_43370# a_n2472_46090# 3.22e-20
C17432 a_11599_46634# a_10903_43370# 0.439916f
C17433 a_4791_45118# a_6945_45028# 0.493927f
C17434 a_13717_47436# a_13925_46122# 5.15e-19
C17435 a_12861_44030# a_13759_46122# 0.032694f
C17436 a_20916_46384# a_20107_46660# 8.05e-20
C17437 a_19321_45002# a_20623_46660# 3.43e-19
C17438 a_13747_46662# a_21188_46660# 2.57e-20
C17439 a_11309_47204# a_11415_45002# 0.001299f
C17440 a_7577_46660# a_8035_47026# 0.027606f
C17441 a_n743_46660# a_16388_46812# 0.035819f
C17442 a_3055_46660# a_3090_45724# 9.03e-20
C17443 a_n2661_46634# a_765_45546# 1.82448f
C17444 a_10227_46804# a_5937_45572# 2.11e-20
C17445 a_4883_46098# a_4419_46090# 0.006295f
C17446 a_19721_31679# VIN_N 0.029175f
C17447 a_n4318_39768# a_n4209_39590# 0.105246f
C17448 a_5649_42852# a_10796_42968# 3.16e-20
C17449 a_18114_32519# VREF 1.12e-19
C17450 a_4361_42308# a_10341_42308# 0.006315f
C17451 a_11341_43940# a_15959_42545# 1.71e-21
C17452 a_15493_43940# a_15764_42576# 1.53e-21
C17453 a_n97_42460# a_n3674_37592# 0.012074f
C17454 a_743_42282# a_12895_43230# 6.86e-20
C17455 a_15743_43084# a_20922_43172# 0.004395f
C17456 a_2779_44458# VDD 0.38604f
C17457 a_n863_45724# a_n2129_43609# 0.003134f
C17458 a_n2661_43370# a_5518_44484# 0.001247f
C17459 a_22223_45036# a_20193_45348# 2.8e-19
C17460 a_16327_47482# a_21335_42336# 0.081786f
C17461 a_4185_45028# a_22223_43396# 3.93e-19
C17462 a_3232_43370# a_13213_44734# 6.1e-21
C17463 a_13507_46334# a_17531_42308# 1.18e-20
C17464 a_526_44458# a_9803_43646# 0.170855f
C17465 a_n2293_45546# a_n1699_43638# 6.05e-20
C17466 a_5205_44484# a_n2661_42834# 0.030553f
C17467 w_1575_34946# VDAC_P 0.037571f
C17468 a_19692_46634# a_19553_46090# 1.1e-19
C17469 a_19466_46812# a_19335_46494# 0.017838f
C17470 a_n881_46662# a_5437_45600# 0.001471f
C17471 a_n1613_43370# a_6812_45938# 0.00201f
C17472 a_n743_46660# a_3316_45546# 2.86e-19
C17473 a_33_46660# a_997_45618# 7.11e-21
C17474 a_5807_45002# a_2711_45572# 0.065611f
C17475 a_10428_46928# a_8049_45260# 2.57e-20
C17476 a_15227_44166# a_19900_46494# 0.053335f
C17477 a_14035_46660# a_13925_46122# 0.207108f
C17478 a_14180_46812# a_13759_46122# 0.001754f
C17479 a_13885_46660# a_14493_46090# 0.001138f
C17480 a_16292_46812# a_6945_45028# 3.43e-20
C17481 a_15368_46634# a_10809_44734# 0.002169f
C17482 a_n2840_46090# a_n2157_46122# 7.58e-21
C17483 a_n2472_46090# a_n2293_46098# 0.176709f
C17484 a_765_45546# a_8199_44636# 8.72e-20
C17485 a_n2661_46098# a_n2840_45546# 3.06e-19
C17486 a_11453_44696# a_13527_45546# 4.99e-21
C17487 a_4190_30871# a_18548_42308# 0.001263f
C17488 a_13291_42460# a_14635_42282# 0.111986f
C17489 a_4361_42308# a_18057_42282# 0.008747f
C17490 a_n2293_42282# a_n1630_35242# 0.18361f
C17491 a_22223_43948# VDD 0.254313f
C17492 a_133_42852# a_196_42282# 4.15e-19
C17493 a_13678_32519# a_17303_42282# 0.008395f
C17494 a_5649_42852# a_4958_30871# 0.293366f
C17495 a_8387_43230# a_8325_42308# 0.003469f
C17496 a_8037_42858# a_8791_42308# 0.002879f
C17497 a_4743_44484# a_3905_42865# 3.75e-22
C17498 a_4223_44672# a_5013_44260# 0.07599f
C17499 a_n913_45002# a_3539_42460# 0.359316f
C17500 a_n2017_45002# a_n998_43396# 5.23e-20
C17501 a_1307_43914# a_13565_43940# 0.004697f
C17502 a_n1917_44484# a_n4318_39768# 6.9e-19
C17503 a_17719_45144# a_17973_43940# 6.82e-19
C17504 a_11453_44696# EN_OFFSET_CAL 7.26e-19
C17505 a_n357_42282# a_19339_43156# 0.008506f
C17506 a_n2956_39304# a_n2472_42282# 2.99e-20
C17507 a_n2956_38680# a_n3674_38680# 0.023107f
C17508 a_4185_45028# a_5934_30871# 0.060401f
C17509 a_1423_45028# a_9801_43940# 5.54e-20
C17510 a_8696_44636# a_16759_43396# 1.51e-21
C17511 a_13507_46334# a_18184_42460# 0.505552f
C17512 a_18597_46090# a_11827_44484# 0.039373f
C17513 a_n743_46660# a_13777_45326# 1.09e-20
C17514 a_20708_46348# a_20850_46482# 0.007833f
C17515 a_18985_46122# a_20850_46155# 4.3e-20
C17516 a_3699_46348# a_2711_45572# 2.78e-20
C17517 a_4791_45118# a_8103_44636# 0.048713f
C17518 a_4646_46812# a_413_45260# 3.52e-20
C17519 a_11415_45002# a_10490_45724# 1.25e-19
C17520 a_11453_44696# a_16922_45042# 0.07136f
C17521 a_10227_46804# a_11691_44458# 0.012084f
C17522 a_8034_45724# a_8781_46436# 0.009374f
C17523 a_5066_45546# a_10586_45546# 9.49e-20
C17524 a_10150_46912# a_3357_43084# 1.08e-20
C17525 a_3090_45724# a_17786_45822# 0.003629f
C17526 a_2324_44458# a_n2293_45546# 9.66e-19
C17527 a_4883_46098# a_18911_45144# 8.04e-21
C17528 a_n1630_35242# a_n3565_39590# 0.036902f
C17529 a_13575_42558# a_13333_42558# 3.68e-20
C17530 a_n3674_37592# a_n3420_39616# 0.019754f
C17531 a_5534_30871# CAL_P 0.006743f
C17532 a_n13_43084# VDD 0.260551f
C17533 a_n4318_38216# a_n4334_39392# 1.1e-19
C17534 a_5379_42460# a_7174_31319# 3.55e-20
C17535 COMP_P a_1736_39587# 0.007099f
C17536 a_13887_32519# VREF 3.68e-19
C17537 a_5891_43370# a_6765_43638# 7.33e-21
C17538 a_1307_43914# a_5534_30871# 3.06e-20
C17539 a_10193_42453# a_11323_42473# 0.034215f
C17540 a_14673_44172# a_n97_42460# 1.2e-19
C17541 a_20820_30879# VDD 0.719502f
C17542 a_21076_30879# C9_N_btm 0.001137f
C17543 a_7640_43914# a_7287_43370# 0.001047f
C17544 a_18184_42460# a_21855_43396# 1.51e-19
C17545 a_n2293_42834# a_2075_43172# 0.005552f
C17546 a_14539_43914# a_14579_43548# 0.002303f
C17547 a_10057_43914# a_10849_43646# 0.003423f
C17548 a_20202_43084# SINGLE_ENDED 1.07e-19
C17549 a_n2956_38216# a_n4209_39590# 0.021267f
C17550 a_18494_42460# a_4361_42308# 0.061307f
C17551 a_22591_46660# RST_Z 4.25e-19
C17552 a_19321_45002# a_20637_44484# 1.7e-20
C17553 a_13661_43548# a_20512_43084# 0.00101f
C17554 a_13747_46662# a_21145_44484# 8.01e-19
C17555 a_20273_46660# a_20567_45036# 4.15e-22
C17556 a_17339_46660# a_11691_44458# 0.018074f
C17557 a_12594_46348# a_13017_45260# 4.35e-20
C17558 a_5937_45572# a_1307_43914# 0.101589f
C17559 a_3090_45724# a_10157_44484# 5.31e-20
C17560 a_16375_45002# a_18479_45785# 1.81e-19
C17561 a_526_44458# a_n913_45002# 0.250864f
C17562 a_n1925_42282# a_n1059_45260# 0.023119f
C17563 a_8049_45260# a_20719_45572# 6.29e-19
C17564 a_10903_43370# a_13348_45260# 0.011259f
C17565 a_2711_45572# a_15143_45578# 0.009403f
C17566 a_6165_46155# a_1423_45028# 4.27e-22
C17567 a_2324_44458# a_6709_45028# 0.076559f
C17568 a_167_45260# a_45_45144# 0.002149f
C17569 a_4185_45028# a_4185_45348# 0.009825f
C17570 a_11415_45002# a_14976_45348# 7.17e-19
C17571 a_1823_45246# a_2448_45028# 7.38e-19
C17572 a_n1613_43370# a_895_43940# 8.02e-21
C17573 a_4700_47436# a_n1613_43370# 5.19e-21
C17574 a_4915_47217# a_5063_47570# 0.003687f
C17575 a_n443_46116# a_3094_47243# 4.19e-19
C17576 a_10227_46804# a_18479_47436# 1.40697f
C17577 a_14311_47204# a_12465_44636# 0.004308f
C17578 a_11599_46634# a_4883_46098# 0.261488f
C17579 a_15811_47375# a_13507_46334# 0.002419f
C17580 a_5934_30871# VREF_GND 0.002663f
C17581 a_13717_47436# SMPL_ON_N 0.132417f
C17582 a_n4315_30879# VDAC_P 0.003601f
C17583 a_n4334_38304# a_n4064_37984# 0.410244f
C17584 a_n3690_38304# a_n3420_37984# 0.414894f
C17585 a_n3565_38216# a_n2946_37984# 0.411006f
C17586 a_n4209_38216# a_n2302_37984# 0.407312f
C17587 a_2684_37794# a_2113_38308# 0.468006f
C17588 a_11323_42473# VDD 0.205172f
C17589 a_n1151_42308# a_8128_46384# 0.328697f
C17590 a_4007_47204# a_n881_46662# 4.68e-20
C17591 a_16327_47482# a_20894_47436# 4.5e-21
C17592 a_2063_45854# a_12891_46348# 4.37e-20
C17593 a_22465_38105# CAL_N 0.072253f
C17594 a_458_43396# a_1049_43396# 0.052073f
C17595 a_n97_42460# a_766_43646# 5.09e-19
C17596 a_11341_43940# a_16243_43396# 1.07e-19
C17597 en_comp comp_n 0.026896f
C17598 a_n2956_37592# a_n2860_39072# 3.22e-20
C17599 a_6511_45714# DATA[3] 1.62e-21
C17600 a_18451_43940# a_15743_43084# 0.005843f
C17601 a_15493_43396# a_18525_43370# 0.031354f
C17602 a_453_43940# a_685_42968# 1.15e-21
C17603 a_19006_44850# a_18599_43230# 2.2e-20
C17604 a_11967_42832# a_18817_42826# 6.37e-20
C17605 a_9313_44734# a_10793_43218# 1.08e-19
C17606 a_4185_45028# a_20512_43084# 2.96e-20
C17607 a_21513_45002# a_2437_43646# 0.009475f
C17608 a_19692_46634# a_15493_43940# 0.16692f
C17609 a_n2293_45546# a_n1699_44726# 0.001074f
C17610 a_n2293_46634# a_8147_43396# 0.011922f
C17611 a_21363_45546# a_21542_45572# 0.007399f
C17612 a_n863_45724# a_n2129_44697# 2.81e-19
C17613 a_526_44458# a_556_44484# 0.077901f
C17614 a_7499_43078# a_8560_45348# 0.006911f
C17615 a_17583_46090# a_17517_44484# 5.71e-21
C17616 a_10227_46804# a_4190_30871# 6.29e-20
C17617 a_16327_47482# a_19095_43396# 6.39e-19
C17618 a_13059_46348# a_12429_44172# 8.69e-20
C17619 a_11453_44696# a_15743_43084# 9.67e-22
C17620 a_380_45546# a_n2661_44458# 2.29e-20
C17621 a_13259_45724# a_12883_44458# 0.003043f
C17622 a_21350_45938# a_3357_43084# 3.05e-19
C17623 a_21188_45572# a_21297_45572# 0.007416f
C17624 C0_P_btm VDD 1.02806f
C17625 a_18194_35068# VIN_N 0.066301f
C17626 a_16327_47482# a_20411_46873# 5.72e-19
C17627 a_12549_44172# a_11901_46660# 0.001645f
C17628 a_12891_46348# a_12469_46902# 0.009064f
C17629 a_11309_47204# a_12251_46660# 1.48e-19
C17630 a_13507_46334# a_13059_46348# 0.192049f
C17631 a_10227_46804# a_17829_46910# 4.34e-19
C17632 a_18479_47436# a_17339_46660# 3.12e-20
C17633 a_2443_46660# a_4651_46660# 1.35e-19
C17634 a_3524_46660# a_3686_47026# 0.006453f
C17635 a_2959_46660# a_3221_46660# 0.001705f
C17636 a_2609_46660# a_4646_46812# 4.37e-20
C17637 a_3177_46902# a_3877_44458# 3.33e-19
C17638 a_2107_46812# a_3633_46660# 2.47e-19
C17639 a_n2109_47186# a_5204_45822# 7.25e-19
C17640 a_n1741_47186# a_5068_46348# 1.28e-20
C17641 a_n2661_46634# a_10623_46897# 0.006678f
C17642 a_584_46384# a_1208_46090# 0.034313f
C17643 a_1431_47204# a_1138_42852# 1.47e-19
C17644 a_n1151_42308# a_n1641_46494# 0.003575f
C17645 a_2063_45854# a_805_46414# 8.93e-20
C17646 a_12861_44030# a_16434_46660# 0.001465f
C17647 a_n881_46662# a_15368_46634# 0.023127f
C17648 a_n971_45724# a_3483_46348# 0.211534f
C17649 a_n237_47217# a_2804_46116# 0.039625f
C17650 a_11599_46634# a_21188_46660# 3.88e-21
C17651 a_18143_47464# a_765_45546# 0.001396f
C17652 C1_N_btm C8_N_btm 0.131002f
C17653 C0_N_btm C9_N_btm 0.14782f
C17654 C0_dummy_N_btm C10_N_btm 0.63636f
C17655 C4_N_btm C5_N_btm 15.915401f
C17656 C3_N_btm C6_N_btm 0.134599f
C17657 C2_N_btm C7_N_btm 0.139982f
C17658 a_18579_44172# a_19647_42308# 7.92e-19
C17659 a_3422_30871# a_18907_42674# 2.69e-20
C17660 a_8685_43396# a_10796_42968# 9.94e-21
C17661 a_18114_32519# a_22521_40599# 1.3e-20
C17662 a_n2661_42282# a_6171_42473# 0.013039f
C17663 a_1568_43370# a_1793_42852# 0.011559f
C17664 a_8953_45546# a_8791_43396# 0.012124f
C17665 a_17339_46660# a_4190_30871# 0.005828f
C17666 a_3537_45260# a_6298_44484# 0.001842f
C17667 a_n1059_45260# a_18248_44752# 2.77e-20
C17668 a_n2661_45010# a_n2012_44484# 1.82e-19
C17669 a_20692_30879# a_15493_43940# 1.18e-20
C17670 a_16375_45002# a_14021_43940# 3.38e-20
C17671 a_10775_45002# a_n2661_44458# 8.26e-21
C17672 a_4927_45028# a_4223_44672# 2.44e-19
C17673 a_3232_43370# a_949_44458# 1.95e-20
C17674 a_5111_44636# a_n699_43396# 0.016349f
C17675 a_8696_44636# a_17517_44484# 0.001184f
C17676 a_15861_45028# a_17061_44734# 2.19e-19
C17677 a_1307_43914# a_11691_44458# 0.024289f
C17678 a_13259_45724# a_15037_44260# 3.72e-21
C17679 a_8270_45546# a_9127_43156# 0.002724f
C17680 a_10227_46804# a_n443_42852# 0.043674f
C17681 a_14311_47204# a_2711_45572# 3.64e-21
C17682 a_2107_46812# a_526_44458# 0.008773f
C17683 a_2063_45854# a_11322_45546# 0.105268f
C17684 a_6755_46942# a_7920_46348# 1.43e-19
C17685 a_10623_46897# a_8199_44636# 3.42e-19
C17686 a_10150_46912# a_9625_46129# 2.39e-19
C17687 a_10249_46116# a_8016_46348# 0.001301f
C17688 a_n743_46660# a_5066_45546# 0.124676f
C17689 a_19692_46634# a_12741_44636# 0.022879f
C17690 a_17339_46660# a_17829_46910# 1.33e-19
C17691 a_n1151_42308# a_10053_45546# 2.02e-20
C17692 a_22612_30879# a_8049_45260# 7.79e-20
C17693 a_n2661_46098# a_n967_46494# 8.5e-19
C17694 a_n901_43156# a_n3674_37592# 2e-19
C17695 a_n2293_42282# a_3863_42891# 1.73e-19
C17696 a_644_44056# VDD 0.147321f
C17697 a_4361_42308# a_3318_42354# 8.57e-20
C17698 a_n13_43084# a_n784_42308# 1.77e-19
C17699 a_n1379_43218# COMP_P 1.55e-21
C17700 a_10341_43396# a_15959_42545# 3.32e-20
C17701 a_5534_30871# a_13003_42852# 0.001789f
C17702 a_14543_43071# a_13291_42460# 0.107887f
C17703 a_13460_43230# a_14635_42282# 6.39e-20
C17704 a_n1423_42826# a_n1630_35242# 2.25e-19
C17705 a_743_42282# a_3581_42558# 7.35e-19
C17706 a_18494_42460# a_20397_44484# 3.54e-19
C17707 a_11827_44484# a_19789_44512# 4.59e-19
C17708 a_2905_45572# VDD 1.22598f
C17709 a_9482_43914# a_13483_43940# 0.006325f
C17710 a_9290_44172# a_12800_43218# 1.74e-20
C17711 a_8746_45002# a_10341_43396# 0.002313f
C17712 a_3232_43370# a_11341_43940# 0.112367f
C17713 a_3090_45724# a_14113_42308# 2.41e-20
C17714 a_1431_47204# DATA[1] 0.334099f
C17715 a_2124_47436# DATA[0] 2.79e-21
C17716 a_11691_44458# a_18579_44172# 2.18e-19
C17717 a_18374_44850# a_9313_44734# 3.42e-21
C17718 a_12607_44458# a_n2293_43922# 0.078602f
C17719 a_n2293_42834# a_5013_44260# 3.56e-20
C17720 a_1307_43914# a_8333_44056# 0.006875f
C17721 a_7499_43078# a_8873_43396# 0.001075f
C17722 a_11823_42460# a_13667_43396# 0.107673f
C17723 a_11735_46660# a_11962_45724# 4.42e-20
C17724 a_12741_44636# a_20692_30879# 7.57e-19
C17725 a_22959_46660# a_20205_31679# 0.00182f
C17726 a_22612_30879# a_19479_31679# 0.064572f
C17727 a_n1613_43370# a_3065_45002# 1.12e-20
C17728 a_12465_44636# a_13017_45260# 1.71e-20
C17729 a_20708_46348# a_10809_44734# 1.69e-21
C17730 a_5937_45572# a_8034_45724# 0.052916f
C17731 a_7920_46348# a_8049_45260# 0.003857f
C17732 a_765_45546# a_509_45822# 0.008717f
C17733 a_14226_46987# a_2711_45572# 3.21e-22
C17734 a_3090_45724# a_7499_43078# 0.23734f
C17735 a_11453_44696# a_10775_45002# 6.82e-19
C17736 a_9804_47204# a_413_45260# 6.79e-20
C17737 a_10341_43396# RST_Z 2.8e-19
C17738 a_4190_30871# CAL_P 0.007081f
C17739 a_2713_42308# a_6123_31319# 1.31e-20
C17740 a_1606_42308# a_8325_42308# 1.94e-20
C17741 a_196_42282# a_5742_30871# 7.34e-20
C17742 a_n784_42308# a_11323_42473# 1.56e-20
C17743 a_10765_43646# VDD 0.00801f
C17744 a_5379_42460# a_5932_42308# 0.761308f
C17745 a_n2065_43946# a_n1644_44306# 0.090164f
C17746 a_n1761_44111# a_n3674_39768# 7.14e-19
C17747 a_11967_42832# a_15682_43940# 1.63211f
C17748 a_n755_45592# a_8515_42308# 0.003799f
C17749 a_n1925_42282# a_n4315_30879# 3.26e-20
C17750 a_n1059_45260# a_8387_43230# 0.005946f
C17751 a_n2017_45002# a_9127_43156# 3.46e-19
C17752 a_n913_45002# a_8605_42826# 0.019641f
C17753 a_10193_42453# a_20753_42852# 0.082713f
C17754 a_13259_45724# a_15890_42674# 8.67e-20
C17755 a_12816_46660# VDD 0.293798f
C17756 a_895_43940# a_2675_43914# 0.099822f
C17757 a_2127_44172# a_2998_44172# 0.001419f
C17758 a_2479_44172# a_2889_44172# 0.002826f
C17759 a_4223_44672# a_4699_43561# 2.12e-19
C17760 a_17517_44484# a_20365_43914# 4.82e-21
C17761 a_8270_45546# CLK 7.07e-21
C17762 a_18479_47436# a_18579_44172# 1.01e-20
C17763 a_16327_47482# a_3422_30871# 0.220296f
C17764 a_3877_44458# a_4223_44672# 0.007855f
C17765 a_8049_45260# a_11280_45822# 1.62e-19
C17766 a_13259_45724# a_10490_45724# 1.48e-19
C17767 a_768_44030# a_9159_44484# 0.003496f
C17768 a_12891_46348# a_n2661_42834# 9.68e-21
C17769 a_6755_46942# a_11827_44484# 0.529579f
C17770 a_11309_47204# a_n2661_43922# 1.06e-21
C17771 a_13507_46334# a_20362_44736# 5.2e-22
C17772 a_n2661_45546# a_3775_45552# 0.006201f
C17773 a_18985_46122# a_18479_45785# 1.04e-21
C17774 a_18819_46122# a_18341_45572# 0.00524f
C17775 a_n2293_46098# a_3065_45002# 2.43e-19
C17776 a_11415_45002# a_6171_45002# 1.05801f
C17777 a_167_45260# a_n745_45366# 7.9e-20
C17778 a_n443_46116# a_2479_44172# 0.732848f
C17779 a_n755_45592# a_2711_45572# 0.168218f
C17780 a_n23_47502# a_n1435_47204# 4.14e-19
C17781 a_4700_47436# a_4791_45118# 0.31818f
C17782 a_4007_47204# a_n443_46116# 0.006041f
C17783 a_n1151_42308# a_6151_47436# 0.026437f
C17784 a_2063_45854# a_7903_47542# 1.25e-20
C17785 a_3785_47178# a_5129_47502# 4.3e-19
C17786 a_3815_47204# a_4915_47217# 2.1e-19
C17787 a_5742_30871# a_n4064_37440# 0.004687f
C17788 a_n784_42308# C0_P_btm 0.281635f
C17789 a_20753_42852# VDD 0.193909f
C17790 a_19328_44172# a_3626_43646# 2.27e-20
C17791 a_20679_44626# a_13467_32519# 4.42e-21
C17792 a_9313_44734# a_10083_42826# 0.013808f
C17793 a_n2017_45002# a_17124_42282# 0.002905f
C17794 a_18374_44850# a_18599_43230# 1.49e-21
C17795 a_18989_43940# a_18817_42826# 2.61e-19
C17796 a_5891_43370# a_10341_42308# 2.08e-19
C17797 a_n356_44636# a_16795_42852# 8.61e-19
C17798 a_9028_43914# a_8791_43396# 0.001013f
C17799 a_n2661_43370# a_n4318_38216# 0.002734f
C17800 a_n2293_42834# a_196_42282# 5.62e-20
C17801 a_18579_44172# a_4190_30871# 0.052036f
C17802 a_n2293_43922# a_3681_42891# 7.77e-21
C17803 a_n2661_43922# a_3935_42891# 1.92e-21
C17804 a_2711_45572# a_13017_45260# 0.050114f
C17805 a_3090_45724# a_3600_43914# 3.95e-19
C17806 a_n443_42852# a_1307_43914# 0.05746f
C17807 a_526_44458# a_n2661_44458# 0.087308f
C17808 a_n2293_45546# a_2448_45028# 9.06e-19
C17809 a_7227_45028# a_7276_45260# 0.098279f
C17810 a_6667_45809# a_6709_45028# 0.001946f
C17811 a_6511_45714# a_7705_45326# 8.07e-19
C17812 a_8049_45260# a_11827_44484# 1.09e-19
C17813 a_3483_46348# a_9313_44734# 0.015646f
C17814 a_1823_45246# a_5708_44484# 5.34e-19
C17815 a_16680_45572# a_18596_45572# 3.21e-21
C17816 a_n1613_43370# a_458_43396# 4.14e-20
C17817 a_11415_45002# a_14673_44172# 0.229077f
C17818 a_4880_45572# a_4558_45348# 3.7e-19
C17819 a_n863_45724# a_45_45144# 2.41e-19
C17820 a_19321_45002# a_19478_44056# 1.84e-21
C17821 a_n2956_39768# a_n2661_46634# 0.006224f
C17822 a_n2840_46634# a_n2472_46634# 7.52e-19
C17823 a_n1741_47186# a_13059_46348# 0.001771f
C17824 a_2063_45854# a_12359_47026# 9.65e-22
C17825 a_n1613_43370# a_3067_47026# 0.013046f
C17826 a_6151_47436# a_14084_46812# 5.28e-21
C17827 a_11031_47542# a_11186_47026# 2.5e-19
C17828 a_4915_47217# a_14976_45028# 3.23e-21
C17829 a_22469_39537# a_22717_37285# 0.002793f
C17830 a_4883_46098# a_7411_46660# 4.36e-20
C17831 a_10227_46804# a_10554_47026# 0.166977f
C17832 a_8685_43396# a_15125_43396# 8.47e-19
C17833 a_12281_43396# a_13749_43396# 1.13e-20
C17834 a_n1761_44111# a_1184_42692# 5.67e-20
C17835 a_n37_45144# VDD 0.138f
C17836 a_6197_43396# a_4361_42308# 4.64e-20
C17837 a_10341_43396# a_16243_43396# 0.058241f
C17838 a_13565_43940# a_13635_43156# 7.88e-21
C17839 a_n1557_42282# a_n1641_43230# 7.08e-19
C17840 a_8147_43396# a_743_42282# 2.1e-21
C17841 a_n1549_44318# a_n1630_35242# 5.92e-22
C17842 a_16327_47482# a_18504_43218# 0.002118f
C17843 a_13661_43548# a_18249_42858# 2.04e-19
C17844 a_n1151_42308# a_n473_42460# 0.006908f
C17845 a_22223_45572# a_22223_45036# 0.026152f
C17846 a_10227_46804# a_14635_42282# 0.008414f
C17847 a_11322_45546# a_n2661_42834# 4.07e-19
C17848 a_n2661_45546# a_n1549_44318# 1.94e-21
C17849 a_3357_43084# a_21359_45002# 6.53e-21
C17850 a_19479_31679# a_11827_44484# 0.01397f
C17851 a_n2293_45546# a_n1761_44111# 2.91e-20
C17852 a_2382_45260# a_n2661_43370# 0.03415f
C17853 a_n1079_45724# a_n2065_43946# 5.59e-22
C17854 a_6171_45002# a_6945_45348# 1.2e-19
C17855 a_8696_44636# a_13720_44458# 0.004063f
C17856 a_16115_45572# a_14539_43914# 4.47e-19
C17857 a_4185_45028# a_21381_43940# 1.24e-20
C17858 a_1307_43914# a_375_42282# 1.11e-20
C17859 a_3090_45724# a_15781_43660# 5.85e-20
C17860 a_n743_46660# a_5068_46348# 0.005784f
C17861 a_12549_44172# a_17583_46090# 3.17e-20
C17862 a_1799_45572# a_472_46348# 5.48e-20
C17863 a_n2661_46098# a_376_46348# 0.060405f
C17864 a_1110_47026# a_1176_45822# 6.94e-20
C17865 a_6755_46942# a_14447_46660# 0.001822f
C17866 a_n971_45724# a_n357_42282# 0.271282f
C17867 a_n452_47436# a_n755_45592# 1.25e-21
C17868 a_n1925_46634# a_5204_45822# 2.89e-19
C17869 a_584_46384# a_n2661_45546# 0.100439f
C17870 a_12469_46902# a_12359_47026# 0.097745f
C17871 a_12251_46660# a_12156_46660# 0.049827f
C17872 a_3090_45724# a_15227_44166# 0.428743f
C17873 a_11599_46634# a_11608_46482# 7.81e-19
C17874 a_2107_46812# a_2521_46116# 0.008501f
C17875 a_1983_46706# a_167_45260# 2.62e-20
C17876 a_n746_45260# a_310_45028# 0.378188f
C17877 a_13661_43548# a_10903_43370# 9.73e-19
C17878 a_5807_45002# a_12005_46116# 0.004606f
C17879 a_15743_43084# a_19273_43230# 0.001058f
C17880 a_n97_42460# a_15959_42545# 0.005005f
C17881 a_6031_43396# a_6123_31319# 6.63e-20
C17882 a_13635_43156# a_5534_30871# 0.078849f
C17883 a_13460_43230# a_14543_43071# 0.001783f
C17884 a_6197_43396# a_6761_42308# 1.61e-19
C17885 a_2982_43646# a_9223_42460# 1.29e-19
C17886 a_3626_43646# a_8685_42308# 0.002659f
C17887 a_13213_44734# VDD 0.184239f
C17888 a_791_42968# a_873_42968# 0.004937f
C17889 a_4520_42826# a_n2293_42282# 3.87e-20
C17890 a_16823_43084# a_16877_43172# 0.001729f
C17891 a_n2293_43922# RST_Z 4.75e-21
C17892 a_13259_45724# a_16547_43609# 3.22e-20
C17893 a_9290_44172# a_10341_42308# 0.051084f
C17894 a_4185_45028# a_18249_42858# 3.07e-20
C17895 a_6298_44484# a_8701_44490# 2.01e-20
C17896 a_n443_42852# a_9396_43370# 0.039136f
C17897 a_3065_45002# a_2675_43914# 8.4e-22
C17898 a_2382_45260# a_2998_44172# 0.045272f
C17899 a_n2293_45010# a_261_44278# 1.74e-19
C17900 a_n2956_38680# a_n4318_38680# 0.023283f
C17901 a_10903_43370# a_10835_43094# 0.001283f
C17902 a_5518_44484# a_5883_43914# 5.07e-20
C17903 a_n2956_37592# a_n3674_39768# 0.024317f
C17904 en_comp a_n4318_39768# 2e-19
C17905 a_3357_43084# a_n2661_42282# 0.028477f
C17906 a_18175_45572# a_15493_43940# 6.32e-22
C17907 a_22612_30879# a_13258_32519# 0.065697f
C17908 a_16763_47508# a_3357_43084# 4.84e-19
C17909 a_12549_44172# a_8696_44636# 0.035105f
C17910 a_6545_47178# a_413_45260# 3.66e-19
C17911 a_4883_46098# a_20841_45814# 5.36e-20
C17912 a_16327_47482# a_19963_31679# 1.05e-19
C17913 a_18479_47436# a_20885_45572# 6.01e-19
C17914 a_3483_46348# a_12594_46348# 0.011082f
C17915 a_21542_46660# a_10809_44734# 4.32e-19
C17916 a_8016_46348# a_5937_45572# 0.021789f
C17917 a_8349_46414# a_8199_44636# 0.032352f
C17918 a_n443_46116# a_2680_45002# 0.009148f
C17919 a_4791_45118# a_3065_45002# 0.006346f
C17920 a_20894_47436# a_20731_45938# 3.6e-21
C17921 a_13507_46334# a_21363_45546# 3.97e-19
C17922 a_10227_46804# a_2437_43646# 0.150025f
C17923 a_n1151_42308# a_5111_44636# 8.63e-19
C17924 a_19466_46812# a_19240_46482# 0.003742f
C17925 a_1138_42852# a_2324_44458# 9.6e-21
C17926 a_4185_45028# a_10903_43370# 1.24e-19
C17927 a_n3674_39304# a_n3420_39072# 0.065079f
C17928 a_n2104_42282# a_n4318_37592# 0.033328f
C17929 a_n4318_38216# COMP_P 5.3e-20
C17930 a_n3674_38216# a_n1736_42282# 7.03e-19
C17931 a_104_43370# VDD 0.252393f
C17932 a_n97_42460# RST_Z 2.62e-20
C17933 a_18083_42858# a_17303_42282# 7.17e-20
C17934 a_17701_42308# a_17531_42308# 0.109201f
C17935 a_9114_42852# a_5934_30871# 5.71e-20
C17936 a_3080_42308# C0_P_btm 0.018211f
C17937 a_n443_42852# a_13003_42852# 1.06e-19
C17938 a_18287_44626# a_18079_43940# 0.007509f
C17939 a_18248_44752# a_18326_43940# 7.79e-19
C17940 a_20362_44736# a_20637_44484# 0.007416f
C17941 a_8975_43940# a_11341_43940# 1.83e-19
C17942 a_5883_43914# a_9895_44260# 2.92e-19
C17943 a_2443_46660# VDD 0.413663f
C17944 a_n2661_42834# a_7281_43914# 0.010117f
C17945 a_6109_44484# a_6101_44260# 1.75e-20
C17946 a_11967_42832# a_20512_43084# 0.106819f
C17947 a_20679_44626# a_22315_44484# 7.27e-21
C17948 a_20835_44721# a_3422_30871# 2.09e-19
C17949 a_n2017_45002# a_19268_43646# 4.82e-21
C17950 a_n913_45002# a_18783_43370# 2.32e-21
C17951 a_n1059_45260# a_15743_43084# 0.101833f
C17952 a_n2293_42834# a_4699_43561# 3.68e-20
C17953 a_3232_43370# a_10341_43396# 2.1e-19
C17954 a_8953_45002# a_9803_43646# 2.76e-20
C17955 a_n357_42282# a_17665_42852# 8.95e-19
C17956 a_2324_44458# a_11962_45724# 0.004603f
C17957 a_15015_46420# a_11823_42460# 0.001494f
C17958 a_12594_46348# a_14495_45572# 5.14e-20
C17959 a_6755_46942# a_15595_45028# 0.012879f
C17960 a_3877_44458# a_n2293_42834# 3.47e-22
C17961 a_8349_46414# a_8192_45572# 2.67e-20
C17962 a_9625_46129# a_10907_45822# 2.68e-19
C17963 a_3090_45724# a_4558_45348# 0.147318f
C17964 a_n1613_43370# a_6298_44484# 0.02075f
C17965 a_17339_46660# a_2437_43646# 3.78e-20
C17966 a_526_44458# a_5907_45546# 3.52e-20
C17967 a_6945_45028# a_6812_45938# 0.002475f
C17968 a_4915_47217# a_15433_44458# 3.72e-20
C17969 a_3483_46348# a_15037_45618# 1.96e-21
C17970 a_12741_44636# a_18175_45572# 7.5e-20
C17971 a_11453_44696# a_17970_44736# 0.008957f
C17972 a_20528_46660# a_20107_45572# 5.09e-21
C17973 a_11415_45002# a_18909_45814# 0.002265f
C17974 a_19692_46634# a_413_45260# 6.26e-20
C17975 a_13759_46122# a_13904_45546# 0.008324f
C17976 a_5742_30871# a_n3420_39072# 0.005978f
C17977 a_18907_42674# a_7174_31319# 2.21e-20
C17978 a_n3674_38216# a_n4209_37414# 1.61e-20
C17979 a_17303_42282# a_22775_42308# 0.005701f
C17980 a_18548_42308# a_19511_42282# 3.36e-20
C17981 a_n4318_38216# a_n3565_37414# 2.51e-20
C17982 a_742_44458# a_3681_42891# 4.15e-19
C17983 a_22223_43948# a_14021_43940# 2.65e-20
C17984 a_11691_44458# a_13635_43156# 2.7e-21
C17985 a_18184_42460# a_17701_42308# 0.001244f
C17986 a_n1059_45260# a_1606_42308# 0.008752f
C17987 a_n2017_45002# a_1755_42282# 0.012188f
C17988 a_n913_45002# a_1221_42558# 1.43e-20
C17989 a_5663_43940# a_n97_42460# 9.61e-20
C17990 a_n809_44244# a_n1557_42282# 1.48e-21
C17991 a_1414_42308# a_4093_43548# 6.35e-21
C17992 a_2779_44458# a_2075_43172# 1.85e-20
C17993 a_16922_45042# a_19987_42826# 0.00105f
C17994 a_18819_46122# VDD 0.453432f
C17995 a_13759_46122# CLK 2.17e-20
C17996 a_n699_43396# a_791_42968# 6.37e-19
C17997 a_n2293_42834# a_6101_43172# 2.77e-19
C17998 a_895_43940# a_1209_43370# 9.02e-21
C17999 a_2127_44172# a_1568_43370# 3.06e-19
C18000 a_1307_43914# a_14635_42282# 3.78e-20
C18001 a_14495_45572# a_15037_45618# 0.00244f
C18002 a_11823_42460# a_16333_45814# 1.07e-20
C18003 a_n971_45724# a_n144_43396# 0.010576f
C18004 a_584_46384# a_1427_43646# 0.003548f
C18005 a_12861_44030# a_17538_32519# 4.84e-19
C18006 a_11415_45002# a_12607_44458# 1.53e-19
C18007 a_10193_42453# a_16223_45938# 1.24e-19
C18008 a_n863_45724# a_n745_45366# 7.61e-20
C18009 a_20692_30879# a_413_45260# 0.111034f
C18010 a_12549_44172# a_20365_43914# 0.069119f
C18011 a_8049_45260# a_15595_45028# 2.98e-20
C18012 a_13259_45724# a_6171_45002# 0.068737f
C18013 a_11525_45546# a_8696_44636# 2.88e-21
C18014 a_n357_42282# a_n2293_45010# 0.020718f
C18015 a_15227_44166# a_14815_43914# 4.45e-19
C18016 a_n2956_38216# en_comp 1.61e-19
C18017 a_n2661_45546# a_n659_45366# 5.25e-19
C18018 a_n2293_46634# a_n2661_42282# 0.039408f
C18019 a_13661_43548# a_14955_43940# 0.010124f
C18020 a_16327_47482# a_19808_44306# 3.3e-21
C18021 a_8120_45572# a_8192_45572# 0.003395f
C18022 a_n1435_47204# a_948_46660# 7.47e-21
C18023 a_7754_39300# a_5088_37509# 1.3e-19
C18024 a_20990_47178# a_19594_46812# 9.2e-20
C18025 a_20894_47436# a_20843_47204# 0.134298f
C18026 a_10227_46804# a_n2661_46634# 0.030546f
C18027 a_n1741_47186# a_7577_46660# 1.46e-20
C18028 a_2905_45572# a_4646_46812# 2.42e-21
C18029 a_n443_46116# a_2864_46660# 0.006317f
C18030 a_3160_47472# a_3877_44458# 2.11e-19
C18031 a_n1151_42308# a_3221_46660# 8.15e-21
C18032 a_n4064_39072# C1_P_btm 9.59e-21
C18033 a_15811_47375# a_n743_46660# 8.06e-19
C18034 a_2063_45854# a_4817_46660# 8.38e-20
C18035 a_4883_46098# a_13661_43548# 0.032161f
C18036 a_n2946_39866# VDD 0.393552f
C18037 a_10807_43548# a_10341_42308# 0.099222f
C18038 a_10949_43914# a_12379_42858# 3.5e-20
C18039 a_n2661_42834# a_564_42282# 1.13e-20
C18040 a_16223_45938# VDD 0.132317f
C18041 a_n97_42460# a_16243_43396# 0.004882f
C18042 a_6197_43396# a_7274_43762# 1.46e-19
C18043 a_11967_42832# a_16245_42852# 0.002841f
C18044 a_11415_45002# a_14761_44260# 1.35e-19
C18045 a_n357_42282# a_9313_44734# 5.02008f
C18046 a_2437_43646# a_1307_43914# 0.160142f
C18047 a_5937_45572# a_7584_44260# 2.31e-20
C18048 a_12861_44030# a_19339_43156# 1.64e-21
C18049 a_7230_45938# a_6298_44484# 3.58e-20
C18050 a_2680_45002# a_3537_45260# 8.13e-20
C18051 a_3483_46348# a_17737_43940# 8.22e-21
C18052 a_13661_43548# a_5649_42852# 3.72e-21
C18053 a_n1613_43370# a_n967_43230# 2.95e-19
C18054 a_20820_30879# a_14021_43940# 1.28e-20
C18055 a_10227_46804# a_14543_43071# 0.00196f
C18056 a_3065_45002# a_3429_45260# 0.037292f
C18057 a_15903_45785# a_16501_45348# 2.45e-20
C18058 a_11682_45822# a_11691_44458# 2.81e-20
C18059 a_13259_45724# a_14673_44172# 0.006759f
C18060 a_2711_45572# a_18374_44850# 5.8e-21
C18061 w_1575_34946# a_1606_42308# 0.001337f
C18062 a_10150_46912# a_6755_46942# 0.006336f
C18063 a_10428_46928# a_10249_46116# 0.704177f
C18064 a_10467_46802# a_10554_47026# 0.07009f
C18065 a_5257_43370# a_6903_46660# 3.74e-20
C18066 a_11599_46634# a_11387_46155# 0.035936f
C18067 a_n237_47217# a_n1925_42282# 0.109762f
C18068 a_13717_47436# a_13759_46122# 3.79e-20
C18069 a_19594_46812# a_20273_46660# 1.32e-19
C18070 a_13747_46662# a_21363_46634# 8.65e-20
C18071 a_12465_44636# a_3483_46348# 0.210833f
C18072 a_7577_46660# a_7832_46660# 0.056391f
C18073 a_n743_46660# a_13059_46348# 0.060636f
C18074 a_12861_44030# a_13351_46090# 1.04e-19
C18075 a_10227_46804# a_8199_44636# 0.460391f
C18076 a_4883_46098# a_4185_45028# 7.37e-19
C18077 a_n97_42460# a_n327_42558# 0.020924f
C18078 a_18114_32519# VIN_N 0.063295f
C18079 a_5649_42852# a_10835_43094# 1.19e-20
C18080 a_n1177_43370# a_n1630_35242# 5.63e-22
C18081 a_19700_43370# a_19339_43156# 0.012115f
C18082 a_4361_42308# a_10922_42852# 4.19e-20
C18083 a_15493_43940# a_15486_42560# 4.05e-19
C18084 a_11341_43940# a_15803_42450# 1.77e-21
C18085 a_n447_43370# a_n3674_37592# 2.26e-21
C18086 a_16823_43084# a_5342_30871# 3.63e-37
C18087 a_743_42282# a_13113_42826# 3.77e-20
C18088 a_15743_43084# a_19987_42826# 0.008026f
C18089 a_19268_43646# a_19164_43230# 3.42e-20
C18090 a_949_44458# VDD 1.2275f
C18091 a_n863_45724# a_n2433_43396# 3.43e-22
C18092 a_n2661_43370# a_5343_44458# 7.17e-19
C18093 a_11827_44484# a_20193_45348# 0.051742f
C18094 a_16327_47482# a_7174_31319# 4.51e-19
C18095 a_10193_42453# a_11341_43940# 0.082222f
C18096 a_n357_42282# a_20974_43370# 7.13e-19
C18097 a_6171_45002# a_n2661_43922# 0.020767f
C18098 a_3232_43370# a_n2293_43922# 9.68e-21
C18099 a_3357_43084# a_19279_43940# 1.53e-20
C18100 a_13507_46334# a_17303_42282# 1.68549f
C18101 a_4185_45028# a_5649_42852# 8.049951f
C18102 a_526_44458# a_9145_43396# 0.004932f
C18103 SMPL_ON_P a_n2302_38778# 5.6e-20
C18104 a_11823_42460# a_15493_43396# 2.38e-20
C18105 a_n2293_45546# a_n2267_43396# 1.47e-20
C18106 a_19466_46812# a_19553_46090# 0.001855f
C18107 a_19692_46634# a_18985_46122# 4.31e-19
C18108 a_n881_46662# a_6428_45938# 4.11e-19
C18109 a_12465_44636# a_14495_45572# 0.019417f
C18110 a_n743_46660# a_3218_45724# 1.78e-20
C18111 a_601_46902# a_n357_42282# 7.55e-20
C18112 a_10150_46912# a_8049_45260# 2.18e-20
C18113 a_15227_44166# a_20075_46420# 0.060002f
C18114 a_14035_46660# a_13759_46122# 0.162408f
C18115 a_19333_46634# a_19335_46494# 4.28e-19
C18116 a_15559_46634# a_6945_45028# 1.52e-20
C18117 a_13885_46660# a_13925_46122# 0.004214f
C18118 a_n2840_46090# a_n2293_46098# 0.003755f
C18119 a_383_46660# a_310_45028# 4.66e-21
C18120 a_14976_45028# a_10809_44734# 0.001621f
C18121 a_13059_46348# a_11189_46129# 6.1e-21
C18122 a_4361_42308# a_17531_42308# 0.007428f
C18123 a_4190_30871# a_18310_42308# 0.001467f
C18124 a_n2293_42282# a_564_42282# 4.89e-19
C18125 a_743_42282# a_18214_42558# 0.005672f
C18126 a_13678_32519# a_4958_30871# 0.031033f
C18127 a_21855_43396# a_17303_42282# 1.3e-20
C18128 a_8605_42826# a_8325_42308# 2.47e-19
C18129 a_8037_42858# a_8685_42308# 3.44e-20
C18130 a_11341_43940# VDD 1.23655f
C18131 a_4185_45028# a_7963_42308# 6.87e-20
C18132 a_3232_43370# a_n97_42460# 0.113391f
C18133 a_n913_45002# a_3626_43646# 0.104422f
C18134 a_n1059_45260# a_3539_42460# 0.021504f
C18135 a_n2017_45002# a_n1243_43396# 6.69e-20
C18136 a_7_47243# VDD 7.01e-19
C18137 a_1307_43914# a_11257_43940# 7.05e-19
C18138 a_2382_45260# a_1568_43370# 2.74e-21
C18139 a_4223_44672# a_5244_44056# 0.019617f
C18140 a_n1699_44726# a_n4318_39768# 3.3e-19
C18141 a_17719_45144# a_17737_43940# 2.8e-20
C18142 a_n89_47570# DATA[0] 2.46e-19
C18143 a_3357_43084# a_7112_43396# 2.88e-19
C18144 SMPL_ON_N EN_OFFSET_CAL 0.066251f
C18145 a_n443_42852# a_13635_43156# 1.86e-19
C18146 a_n357_42282# a_18599_43230# 0.006999f
C18147 a_n2810_45572# a_n2293_42282# 3.09e-20
C18148 a_n2956_38680# a_n2840_42282# 2.5e-20
C18149 a_n2956_39304# a_n3674_38680# 0.023226f
C18150 a_8696_44636# a_16977_43638# 6.12e-20
C18151 a_15861_45028# a_16409_43396# 2.62e-21
C18152 a_22612_30879# a_22609_37990# 1.7e-20
C18153 a_10467_46802# a_2437_43646# 1.48e-20
C18154 a_13507_46334# a_19778_44110# 1.08e-20
C18155 a_18597_46090# a_21359_45002# 0.008859f
C18156 a_n743_46660# a_13556_45296# 3.23e-21
C18157 a_2107_46812# a_8953_45002# 0.016508f
C18158 a_n2497_47436# a_n23_44458# 4.12e-19
C18159 a_3483_46348# a_2711_45572# 0.167588f
C18160 a_3147_46376# a_3175_45822# 0.001132f
C18161 a_4791_45118# a_6298_44484# 0.033887f
C18162 a_n2293_46098# a_5437_45600# 4.86e-19
C18163 a_3877_44458# a_413_45260# 3.15e-19
C18164 a_5066_45546# a_8379_46155# 0.001042f
C18165 a_8062_46482# a_8049_45260# 2.78e-21
C18166 a_8016_46348# a_n443_42852# 1.96e-19
C18167 a_768_44030# a_2809_45028# 0.005501f
C18168 a_9863_46634# a_3357_43084# 1.66e-20
C18169 a_3090_45724# a_16377_45572# 3.99e-19
C18170 a_13070_42354# a_13333_42558# 0.011552f
C18171 a_13575_42558# a_13249_42558# 2.37e-20
C18172 a_6123_31319# a_4958_30871# 0.021709f
C18173 a_13678_32519# VCM 0.014539f
C18174 a_13887_32519# VIN_N 0.061374f
C18175 a_n1076_43230# VDD 0.292942f
C18176 a_5267_42460# a_7174_31319# 4.88e-21
C18177 COMP_P a_1239_39587# 0.388733f
C18178 a_n1059_45260# a_9061_43230# 1.7e-20
C18179 a_1307_43914# a_14543_43071# 7.06e-21
C18180 a_5891_43370# a_6197_43396# 0.003102f
C18181 a_7499_43078# a_11633_42558# 2.79e-19
C18182 a_10193_42453# a_10723_42308# 0.046812f
C18183 a_n2810_45572# a_n3565_39590# 0.020853f
C18184 a_n2293_43922# a_4905_42826# 2.78e-20
C18185 a_21076_30879# C8_N_btm 0.384801f
C18186 a_n2293_42834# a_1847_42826# 0.078127f
C18187 a_8975_43940# a_10341_43396# 5.7e-20
C18188 a_10057_43914# a_10765_43646# 0.005404f
C18189 a_18184_42460# a_4361_42308# 0.058569f
C18190 a_18494_42460# a_13467_32519# 1.67e-19
C18191 a_11415_45002# RST_Z 4.24e-19
C18192 a_22591_46660# VDD 0.251892f
C18193 a_20411_46873# a_20567_45036# 1.28e-19
C18194 a_9290_44172# a_13777_45326# 1.57e-20
C18195 a_18189_46348# a_6171_45002# 2.69e-20
C18196 a_8199_44636# a_1307_43914# 0.044343f
C18197 a_3090_45724# a_9838_44484# 2.74e-22
C18198 a_16375_45002# a_18175_45572# 0.001125f
C18199 a_526_44458# a_n1059_45260# 0.097646f
C18200 a_n1925_42282# a_n2017_45002# 0.041988f
C18201 a_20273_46660# a_18494_42460# 1.49e-19
C18202 a_8049_45260# a_21350_45938# 1.72e-19
C18203 a_n2312_39304# a_n3674_39768# 0.023328f
C18204 a_10903_43370# a_13159_45002# 2.53e-19
C18205 a_5497_46414# a_1423_45028# 2.85e-22
C18206 a_2324_44458# a_7229_43940# 0.008305f
C18207 a_3483_46348# a_4640_45348# 3.32e-19
C18208 a_11415_45002# a_14403_45348# 3.58e-19
C18209 a_2711_45572# a_14495_45572# 0.008699f
C18210 a_3815_47204# a_n881_46662# 0.001037f
C18211 a_4007_47204# a_n1613_43370# 7.26e-20
C18212 a_n443_46116# a_5063_47570# 0.006259f
C18213 a_16327_47482# a_19787_47423# 2.23e-19
C18214 a_17591_47464# a_18479_47436# 6.29e-19
C18215 a_4958_30871# EN_VIN_BSTR_P 0.021638f
C18216 a_14955_47212# a_4883_46098# 1.4e-20
C18217 a_10227_46804# a_18143_47464# 0.112443f
C18218 a_5742_30871# C10_N_btm 0.00237f
C18219 a_13717_47436# a_22731_47423# 0.109987f
C18220 a_15507_47210# a_13507_46334# 1.32e-19
C18221 a_1177_38525# a_2113_38308# 1.21e-19
C18222 a_n4209_38216# a_n4064_37984# 0.19304f
C18223 a_n3565_38216# a_n3420_37984# 0.238595f
C18224 a_n4064_39616# a_n4064_37440# 0.050913f
C18225 a_10723_42308# VDD 0.223902f
C18226 a_2063_45854# a_11309_47204# 0.141276f
C18227 a_n1151_42308# a_5159_47243# 2.93e-19
C18228 a_13487_47204# a_12465_44636# 0.001864f
C18229 a_6123_31319# VCM 0.144585f
C18230 a_458_43396# a_1209_43370# 0.0172f
C18231 a_n97_42460# a_4905_42826# 0.147727f
C18232 a_11341_43940# a_16137_43396# 3.22e-19
C18233 a_n3674_39768# a_n2472_42826# 1.25e-19
C18234 en_comp a_1736_39043# 2.01e-19
C18235 a_6472_45840# DATA[3] 2.3e-21
C18236 a_18451_43940# a_18783_43370# 0.001344f
C18237 a_15493_43396# a_18429_43548# 0.045352f
C18238 a_n2661_42282# a_743_42282# 0.043675f
C18239 a_11967_42832# a_18249_42858# 0.018824f
C18240 a_9313_44734# a_10553_43218# 7.54e-19
C18241 a_15682_43940# a_16867_43762# 0.001981f
C18242 a_n2661_45546# a_n1177_44458# 3.02e-20
C18243 a_19466_46812# a_15493_43940# 4.43e-22
C18244 a_19692_46634# a_22223_43948# 0.003538f
C18245 a_n452_45724# a_n2661_44458# 5.67e-21
C18246 a_n1079_45724# a_n2129_44697# 4.42e-21
C18247 a_n2293_45546# a_n2267_44484# 3.38e-19
C18248 a_n863_45724# a_n2433_44484# 1.5e-21
C18249 a_10903_43370# a_11967_42832# 0.02192f
C18250 a_n2293_46634# a_7112_43396# 0.012325f
C18251 a_584_46384# a_4520_42826# 0.001248f
C18252 a_13661_43548# a_8685_43396# 8.18e-19
C18253 a_526_44458# a_484_44484# 0.003617f
C18254 a_8568_45546# a_8560_45348# 0.001331f
C18255 SMPL_ON_N a_15743_43084# 4.69e-20
C18256 a_13259_45724# a_12607_44458# 0.132105f
C18257 a_12549_44172# a_14205_43396# 9.74e-21
C18258 a_21188_45572# a_20447_31679# 3.01e-20
C18259 C1_P_btm VDD 0.264503f
C18260 EN_VIN_BSTR_N VIN_N 1.41696f
C18261 a_16327_47482# a_20107_46660# 0.007614f
C18262 a_n1925_46634# a_7927_46660# 0.009262f
C18263 a_5807_45002# a_6903_46660# 5.51e-19
C18264 a_1209_47178# a_1823_45246# 4.52e-19
C18265 a_768_44030# a_11735_46660# 2.94e-21
C18266 a_12891_46348# a_11901_46660# 0.028795f
C18267 a_12549_44172# a_11813_46116# 2.08e-20
C18268 a_4007_47204# a_n2293_46098# 1.9e-21
C18269 a_n881_46662# a_14976_45028# 0.020069f
C18270 a_17591_47464# a_17829_46910# 8.36e-19
C18271 a_2959_46660# a_3055_46660# 0.013793f
C18272 a_3177_46902# a_3221_46660# 3.69e-19
C18273 a_2609_46660# a_3877_44458# 4.32e-19
C18274 a_2443_46660# a_4646_46812# 2.79e-21
C18275 a_n2109_47186# a_5164_46348# 0.603312f
C18276 a_n2661_46634# a_10467_46802# 0.033928f
C18277 a_2063_45854# a_472_46348# 3.39e-19
C18278 a_584_46384# a_805_46414# 0.135394f
C18279 a_1239_47204# a_1138_42852# 9.6e-21
C18280 a_n1151_42308# a_n1423_46090# 0.009064f
C18281 EN_VIN_BSTR_P VCM 0.929333f
C18282 a_n237_47217# a_2698_46116# 0.032015f
C18283 a_n971_45724# a_3147_46376# 0.001884f
C18284 a_n743_46660# a_7577_46660# 6.2e-20
C18285 a_11599_46634# a_21363_46634# 5.21e-21
C18286 a_18143_47464# a_17339_46660# 6.71e-19
C18287 a_10227_46804# a_765_45546# 0.038035f
C18288 C0_dummy_P_btm C10_N_btm 0.001369f
C18289 C3_N_btm C5_N_btm 0.136119f
C18290 C0_N_btm C8_N_btm 0.148433f
C18291 C0_dummy_N_btm C9_N_btm 0.11363f
C18292 C2_N_btm C6_N_btm 0.138423f
C18293 C1_N_btm C7_N_btm 0.129707f
C18294 a_12465_44636# a_14513_46634# 0.01549f
C18295 a_18579_44172# a_19511_42282# 2.1e-20
C18296 a_3422_30871# a_18727_42674# 5.4e-20
C18297 a_17678_43396# a_4190_30871# 5.27e-21
C18298 a_8685_43396# a_10835_43094# 1.12e-19
C18299 a_2982_43646# a_21195_42852# 0.034024f
C18300 a_n1557_42282# a_n2293_42282# 4.61e-19
C18301 a_n2661_42282# a_5755_42308# 0.002898f
C18302 a_16823_43084# a_743_42282# 2.26e-19
C18303 a_1568_43370# a_1709_42852# 0.015873f
C18304 a_3080_42308# a_4156_43218# 0.00153f
C18305 a_n357_42282# a_17737_43940# 1.35e-20
C18306 a_5937_45572# a_8791_43396# 2.23e-21
C18307 a_8199_44636# a_9396_43370# 0.004302f
C18308 a_4558_45348# a_4743_44484# 5.35e-20
C18309 a_n1059_45260# a_17970_44736# 3.79e-19
C18310 a_n2017_45002# a_18248_44752# 3.8e-22
C18311 a_20205_31679# a_15493_43940# 1.01e-20
C18312 a_4185_45028# a_8685_43396# 2.24e-20
C18313 a_5111_44636# a_4223_44672# 0.418299f
C18314 a_8953_45002# a_n2661_44458# 6.7e-19
C18315 a_8696_44636# a_17061_44734# 0.003665f
C18316 a_16019_45002# a_11691_44458# 6.26e-20
C18317 a_8560_45348# a_n2661_43370# 1.75e-19
C18318 a_12465_44636# a_n357_42282# 1.28e-20
C18319 a_2107_46812# a_2981_46116# 0.002293f
C18320 a_9863_46634# a_9625_46129# 0.001647f
C18321 a_10467_46802# a_8199_44636# 3.56e-19
C18322 a_6755_46942# a_6419_46155# 7.31e-19
C18323 a_n1151_42308# a_9049_44484# 1.64e-19
C18324 a_4791_45118# a_5437_45600# 0.001854f
C18325 a_6575_47204# a_7227_45028# 9.87e-21
C18326 a_17339_46660# a_765_45546# 0.244447f
C18327 a_n2312_39304# a_n2293_45546# 6.75e-19
C18328 a_19466_46812# a_12741_44636# 0.043645f
C18329 a_2063_45854# a_10490_45724# 0.082703f
C18330 a_21588_30879# a_8049_45260# 7.12e-20
C18331 a_n2661_46634# a_8034_45724# 1.89e-20
C18332 a_n2661_46098# a_n1379_46482# 0.002086f
C18333 a_n1641_43230# a_n3674_37592# 2.78e-20
C18334 a_175_44278# VDD 0.20887f
C18335 a_n901_43156# a_n327_42558# 0.001558f
C18336 a_n1076_43230# a_n784_42308# 9.15e-21
C18337 a_n13_43084# a_196_42282# 2.75e-19
C18338 a_10341_43396# a_15803_42450# 3.14e-20
C18339 a_12281_43396# a_14113_42308# 1.99e-20
C18340 a_13460_43230# a_13291_42460# 3.16e-19
C18341 a_n1991_42858# a_n1630_35242# 1.18e-19
C18342 a_743_42282# a_3497_42558# 0.001105f
C18343 a_21101_45002# a_20980_44850# 0.001202f
C18344 a_11827_44484# a_20596_44850# 1.17e-19
C18345 a_2952_47436# VDD 0.089131f
C18346 a_9482_43914# a_12429_44172# 0.0636f
C18347 a_n2293_42834# a_5244_44056# 6.01e-21
C18348 a_10193_42453# a_10341_43396# 0.064616f
C18349 a_1239_47204# DATA[1] 0.01925f
C18350 a_1431_47204# DATA[0] 3.79e-20
C18351 a_626_44172# a_n2661_42282# 6.14e-21
C18352 a_11691_44458# a_18245_44484# 8.73e-19
C18353 a_12607_44458# a_n2661_43922# 0.060913f
C18354 a_7499_43078# a_12281_43396# 9.62e-20
C18355 a_2711_45572# a_16664_43396# 0.001086f
C18356 a_n357_42282# a_13887_32519# 3.9e-20
C18357 a_13507_46334# a_9482_43914# 2.01e-19
C18358 a_20820_30879# a_20692_30879# 8.973741f
C18359 a_12741_44636# a_20205_31679# 0.003338f
C18360 a_20916_46384# a_3357_43084# 7.98e-19
C18361 a_21588_30879# a_19479_31679# 0.055797f
C18362 a_n881_46662# a_2382_45260# 6.99e-22
C18363 a_21137_46414# a_6945_45028# 0.042885f
C18364 a_19900_46494# a_10809_44734# 3.7e-20
C18365 a_8199_44636# a_8034_45724# 0.127067f
C18366 a_14513_46634# a_2711_45572# 3.9e-21
C18367 a_11901_46660# a_11322_45546# 8.73e-20
C18368 a_11813_46116# a_11525_45546# 6.46e-19
C18369 a_8128_46384# a_413_45260# 4.76e-20
C18370 a_11453_44696# a_8953_45002# 6.78e-19
C18371 a_4883_46098# a_13159_45002# 2.87e-21
C18372 a_4933_42558# a_4921_42308# 0.012385f
C18373 a_17364_32525# VDAC_N 0.002821f
C18374 a_n784_42308# a_10723_42308# 3.86e-20
C18375 a_10341_43396# VDD 0.401264f
C18376 a_5267_42460# a_5932_42308# 0.026805f
C18377 a_5379_42460# a_6171_42473# 0.110293f
C18378 a_n2065_43946# a_n3674_39768# 0.001814f
C18379 a_n1761_44111# a_n4318_39768# 2.23e-20
C18380 a_1414_42308# a_3600_43914# 0.012293f
C18381 a_11967_42832# a_14955_43940# 1.47e-21
C18382 a_n755_45592# a_5934_30871# 0.040823f
C18383 a_n357_42282# a_8515_42308# 2.87e-20
C18384 a_n913_45002# a_8037_42858# 0.316376f
C18385 a_n1059_45260# a_8605_42826# 0.007493f
C18386 a_n2017_45002# a_8387_43230# 4.99e-20
C18387 a_n2956_38680# a_n2302_39866# 2.07e-19
C18388 a_10193_42453# a_20356_42852# 4.95e-19
C18389 a_13259_45724# a_15959_42545# 1.16e-19
C18390 a_12991_46634# VDD 0.357655f
C18391 a_2127_44172# a_2889_44172# 7.46e-20
C18392 a_2479_44172# a_2675_43914# 0.061502f
C18393 a_453_43940# a_2998_44172# 1.49e-21
C18394 a_n699_43396# a_4093_43548# 2.73e-20
C18395 a_4223_44672# a_4235_43370# 5.04e-19
C18396 a_17517_44484# a_20269_44172# 5.36e-20
C18397 a_413_45260# a_1847_42826# 2.14e-20
C18398 a_16327_47482# a_21398_44850# 2.55e-19
C18399 a_8049_45260# a_10907_45822# 0.010337f
C18400 a_8034_45724# a_8192_45572# 0.002594f
C18401 a_768_44030# a_10617_44484# 0.001771f
C18402 a_n971_45724# a_n1441_43940# 7.56e-19
C18403 a_n881_46662# a_15433_44458# 3.48e-21
C18404 a_8016_46348# a_2437_43646# 3.18e-20
C18405 a_4883_46098# a_11967_42832# 5.15e-22
C18406 a_18985_46122# a_18175_45572# 0.009338f
C18407 a_18819_46122# a_18479_45785# 2.67e-20
C18408 a_17957_46116# a_18341_45572# 1.43e-19
C18409 a_11415_45002# a_3232_43370# 4.11e-19
C18410 a_n443_46116# a_2127_44172# 0.196411f
C18411 a_6165_46155# a_3357_43084# 0.009006f
C18412 a_3090_45724# a_n2661_43370# 0.101361f
C18413 a_n755_45592# a_1609_45572# 5.85e-19
C18414 a_997_45618# a_1260_45572# 0.010598f
C18415 a_n357_42282# a_2711_45572# 0.039058f
C18416 a_18597_46090# a_19279_43940# 0.021978f
C18417 a_n237_47217# a_n1435_47204# 0.001134f
C18418 a_4007_47204# a_4791_45118# 0.002181f
C18419 a_3815_47204# a_n443_46116# 9.13e-19
C18420 a_3785_47178# a_4915_47217# 0.006427f
C18421 a_n1151_42308# a_5815_47464# 0.001311f
C18422 a_n2946_39866# a_n2946_39072# 0.052227f
C18423 a_n4064_39616# a_n3420_39072# 0.05019f
C18424 a_n3420_39616# a_n4064_39072# 6.32746f
C18425 a_1736_39587# a_1343_38525# 0.289453f
C18426 a_n4315_30879# a_n4209_38502# 0.082287f
C18427 a_20356_42852# VDD 7.06e-19
C18428 a_n784_42308# C1_P_btm 0.027772f
C18429 a_2711_45572# CAL_N 6.22e-19
C18430 a_11967_42832# a_5649_42852# 1.63e-19
C18431 a_20640_44752# a_13467_32519# 1.11e-19
C18432 a_9313_44734# a_8952_43230# 1.48e-19
C18433 a_5111_44636# a_5742_30871# 1.17e-20
C18434 a_n2017_45002# a_16522_42674# 0.002301f
C18435 a_n913_45002# a_13921_42308# 2.11e-20
C18436 a_n1059_45260# a_16104_42674# 4.45e-19
C18437 a_18989_43940# a_18249_42858# 4.24e-19
C18438 a_18287_44626# a_19339_43156# 3.19e-19
C18439 a_n2293_42834# a_n473_42460# 0.001023f
C18440 a_18579_44172# a_21259_43561# 8.21e-19
C18441 a_n2661_43922# a_3681_42891# 5.11e-21
C18442 a_n2293_43922# a_2905_42968# 1.12e-20
C18443 a_n2661_42834# a_3935_42891# 3.28e-21
C18444 a_13259_45724# RST_Z 0.003467f
C18445 a_2711_45572# a_11963_45334# 1.25e-20
C18446 a_3733_45822# a_3232_43370# 5.07e-20
C18447 a_3090_45724# a_2998_44172# 0.001518f
C18448 a_6945_45028# a_6298_44484# 0.00332f
C18449 a_n2293_45546# a_117_45144# 6.33e-19
C18450 a_6511_45714# a_6709_45028# 0.001019f
C18451 a_8049_45260# a_21359_45002# 2.51e-22
C18452 a_13259_45724# a_14403_45348# 0.001862f
C18453 a_1823_45246# a_5608_44484# 3.64e-19
C18454 a_16333_45814# a_16789_45572# 4.2e-19
C18455 a_15599_45572# a_17668_45572# 1.29e-20
C18456 a_17339_46660# a_18681_44484# 5.66e-19
C18457 a_n1613_43370# a_n229_43646# 3.21e-19
C18458 a_11415_45002# a_14581_44484# 0.009374f
C18459 a_376_46348# a_n2661_43922# 2.93e-22
C18460 a_2324_44458# a_15004_44636# 2.94e-20
C18461 a_13747_46662# a_21205_44306# 5.28e-19
C18462 a_n2840_46634# a_n2661_46634# 0.180867f
C18463 a_2063_45854# a_12156_46660# 2.28e-19
C18464 a_n881_46662# a_3524_46660# 2.99e-19
C18465 a_n1613_43370# a_2864_46660# 0.014165f
C18466 a_6151_47436# a_13607_46688# 2.73e-20
C18467 a_4915_47217# a_3090_45724# 2.35e-20
C18468 a_22469_39537# a_22705_37990# 3.12e-20
C18469 CAL_P a_22609_38406# 2.83e-19
C18470 a_4883_46098# a_5257_43370# 0.026597f
C18471 a_10227_46804# a_10623_46897# 0.180903f
C18472 a_8685_43396# a_15037_43396# 1.41e-19
C18473 a_6293_42852# a_4361_42308# 1.16e-19
C18474 a_n143_45144# VDD 0.092f
C18475 a_10341_43396# a_16137_43396# 0.021507f
C18476 a_n1557_42282# a_n1423_42826# 9.17e-20
C18477 a_14955_43396# a_16547_43609# 5.64e-21
C18478 a_n356_44636# a_7174_31319# 2.55e-20
C18479 a_n809_44244# a_n3674_37592# 3.34e-21
C18480 a_6755_46942# a_16823_43084# 1.01e-19
C18481 a_13661_43548# a_17333_42852# 1.34e-20
C18482 a_n1151_42308# a_n961_42308# 0.109068f
C18483 a_1307_43914# a_16751_45260# 1.36e-19
C18484 a_13249_42308# a_9313_44734# 0.031106f
C18485 a_8746_45002# a_n2661_43922# 0.003872f
C18486 a_10193_42453# a_n2293_43922# 0.024214f
C18487 a_10490_45724# a_n2661_42834# 4.83e-22
C18488 a_2437_43646# a_22223_45036# 3.35e-19
C18489 a_22223_45572# a_11827_44484# 0.00211f
C18490 a_10227_46804# a_13291_42460# 0.002348f
C18491 a_5257_43370# a_5649_42852# 8.9e-19
C18492 a_5111_44636# a_n2293_42834# 0.110286f
C18493 a_3357_43084# a_21101_45002# 2.54e-21
C18494 a_21513_45002# a_22959_45036# 7.2e-21
C18495 a_19479_31679# a_21359_45002# 3.83e-19
C18496 a_n2293_45546# a_n2065_43946# 2.73e-20
C18497 a_2274_45254# a_n2661_43370# 0.019962f
C18498 a_6171_45002# a_5837_45028# 0.001502f
C18499 a_8696_44636# a_13076_44458# 0.003013f
C18500 a_16115_45572# a_16112_44458# 7.96e-20
C18501 a_3090_45724# a_15681_43442# 3.44e-19
C18502 a_584_46384# a_564_42282# 7.22e-21
C18503 a_n2293_46634# a_12545_42858# 3.58e-20
C18504 a_768_44030# a_2324_44458# 0.047942f
C18505 a_12549_44172# a_15682_46116# 6.67e-19
C18506 a_n2661_46098# a_n1076_46494# 0.037593f
C18507 a_1983_46706# a_2202_46116# 0.001054f
C18508 a_10467_46802# a_765_45546# 0.003784f
C18509 a_6755_46942# a_14226_46660# 0.001921f
C18510 a_n815_47178# a_n755_45592# 2.36e-20
C18511 a_n1925_46634# a_5164_46348# 2.7e-19
C18512 a_n743_46660# a_4704_46090# 0.011859f
C18513 a_11901_46660# a_12359_47026# 0.034619f
C18514 a_n2661_46634# a_8016_46348# 1.16e-19
C18515 a_2107_46812# a_167_45260# 0.012514f
C18516 a_n971_45724# a_310_45028# 4.56e-21
C18517 a_n237_47217# a_380_45546# 6.95e-20
C18518 a_n746_45260# a_n1099_45572# 0.015931f
C18519 a_5807_45002# a_10903_43370# 0.002924f
C18520 a_15743_43084# a_18861_43218# 3.78e-19
C18521 a_n97_42460# a_15803_42450# 0.004106f
C18522 a_6031_43396# a_7227_42308# 2.05e-20
C18523 a_13635_43156# a_14543_43071# 0.013803f
C18524 a_12895_43230# a_5534_30871# 0.004896f
C18525 a_3626_43646# a_8325_42308# 0.001817f
C18526 a_2982_43646# a_8791_42308# 2.53e-19
C18527 a_n2293_43922# VDD 0.735248f
C18528 a_685_42968# a_873_42968# 7.47e-21
C18529 a_3935_42891# a_n2293_42282# 8.93e-19
C18530 a_13259_45724# a_16243_43396# 1.45e-20
C18531 a_9290_44172# a_10922_42852# 0.028552f
C18532 a_4185_45028# a_17333_42852# 1.67e-20
C18533 a_n443_42852# a_8791_43396# 0.053902f
C18534 a_2680_45002# a_2675_43914# 0.001197f
C18535 a_n2293_45010# a_n1441_43940# 0.009441f
C18536 a_n2956_38680# a_n3674_39304# 0.023431f
C18537 a_n2956_39304# a_n4318_38680# 0.023405f
C18538 a_10903_43370# a_10518_42984# 8.08e-19
C18539 a_6298_44484# a_8103_44636# 0.016067f
C18540 a_5343_44458# a_5883_43914# 0.042199f
C18541 a_n2956_37592# a_n4318_39768# 0.029002f
C18542 a_3357_43084# a_6101_44260# 4.26e-19
C18543 a_2324_44458# a_5755_42852# 3.34e-19
C18544 a_n2810_45028# a_n3674_39768# 0.023163f
C18545 a_10193_42453# a_n97_42460# 0.304653f
C18546 a_18479_45785# a_11341_43940# 0.019493f
C18547 a_16147_45260# a_15493_43940# 2.22e-19
C18548 a_21588_30879# a_13258_32519# 0.062822f
C18549 a_18597_46090# a_19610_45572# 4.96e-19
C18550 a_16023_47582# a_3357_43084# 2.06e-19
C18551 a_16327_47482# a_22591_45572# 1.29e-19
C18552 a_n1925_46634# a_8336_45822# 0.003059f
C18553 a_12891_46348# a_8696_44636# 0.028033f
C18554 a_2063_45854# a_6171_45002# 0.029207f
C18555 a_15227_44166# a_19431_46494# 0.001203f
C18556 a_6151_47436# a_413_45260# 3.16e-19
C18557 a_4883_46098# a_20273_45572# 9.32e-20
C18558 a_n2661_46634# a_11682_45822# 0.010865f
C18559 a_7920_46348# a_5937_45572# 4.23e-21
C18560 a_8016_46348# a_8199_44636# 0.33718f
C18561 a_765_45546# a_8034_45724# 1.01e-21
C18562 a_n443_46116# a_2382_45260# 0.027844f
C18563 a_13507_46334# a_20623_45572# 1.7e-20
C18564 a_n1151_42308# a_5147_45002# 4.06e-20
C18565 a_19466_46812# a_16375_45002# 5.87e-21
C18566 a_21297_46660# a_10809_44734# 2.09e-19
C18567 a_3483_46348# a_12005_46116# 4.4e-21
C18568 a_21076_30879# a_22959_46124# 5.19e-19
C18569 a_6540_46812# a_6472_45840# 3.24e-21
C18570 a_17591_47464# a_2437_43646# 0.013209f
C18571 a_n3674_39304# a_n3690_39392# 0.071784f
C18572 a_n4318_38216# a_n4318_37592# 0.139499f
C18573 a_14401_32519# VIN_N 0.03172f
C18574 a_n97_42460# VDD 3.61113f
C18575 a_17595_43084# a_17531_42308# 0.001512f
C18576 a_17701_42308# a_17303_42282# 0.049097f
C18577 a_n2104_42282# a_n1736_42282# 7.52e-19
C18578 a_n2472_42282# COMP_P 1.38e-19
C18579 a_3080_42308# C1_P_btm 0.011373f
C18580 a_2107_46812# DATA[4] 2.5e-21
C18581 a_18248_44752# a_18079_43940# 6.24e-19
C18582 a_n2956_38680# a_5742_30871# 4.45e-21
C18583 a_5883_43914# a_9801_44260# 3.67e-19
C18584 a_10057_43914# a_11341_43940# 1e-19
C18585 a_n2661_42834# a_6453_43914# 0.007635f
C18586 a_14539_43914# a_15493_43396# 0.024653f
C18587 a_20766_44850# a_20980_44850# 0.097745f
C18588 a_20679_44626# a_3422_30871# 0.078371f
C18589 a_20835_44721# a_21398_44850# 0.049827f
C18590 a_20640_44752# a_22315_44484# 2.12e-19
C18591 a_n2293_42834# a_4235_43370# 0.009569f
C18592 a_18494_42460# a_19319_43548# 0.016978f
C18593 a_n2661_46098# VDD 0.979859f
C18594 a_8953_45002# a_9145_43396# 3.05e-20
C18595 a_n357_42282# a_16877_42852# 0.016936f
C18596 a_n1925_42282# a_4169_42308# 2.9e-19
C18597 a_n1059_45260# a_18783_43370# 7.13e-19
C18598 a_n2017_45002# a_15743_43084# 0.049212f
C18599 a_2324_44458# a_11652_45724# 0.034041f
C18600 a_14275_46494# a_11823_42460# 1.34e-19
C18601 a_12594_46348# a_13249_42308# 4.26e-20
C18602 a_6755_46942# a_15415_45028# 5.84e-21
C18603 a_4646_46812# a_7418_45394# 0.001071f
C18604 a_9625_46129# a_10210_45822# 0.002126f
C18605 a_n1925_42282# a_4099_45572# 0.009682f
C18606 a_526_44458# a_5263_45724# 5.01e-19
C18607 a_4817_46660# a_5093_45028# 5.47e-21
C18608 a_4915_47217# a_14815_43914# 0.006248f
C18609 a_3483_46348# a_14033_45822# 0.030627f
C18610 a_n881_46662# a_5343_44458# 6.79e-19
C18611 a_3090_45724# a_4574_45260# 0.002261f
C18612 a_12741_44636# a_16147_45260# 0.023061f
C18613 a_11453_44696# a_17767_44458# 0.010225f
C18614 a_21188_46660# a_20273_45572# 3.8e-20
C18615 a_20411_46873# a_20528_45572# 3.25e-21
C18616 a_20623_46660# a_20623_45572# 2.72e-19
C18617 a_20273_46660# a_21188_45572# 6.41e-21
C18618 a_11415_45002# a_18341_45572# 0.002269f
C18619 a_19466_46812# a_413_45260# 2.56e-20
C18620 a_12861_44030# a_9313_44734# 0.001011f
C18621 a_18727_42674# a_7174_31319# 4.47e-20
C18622 a_5934_30871# a_n3420_38528# 2.14e-19
C18623 a_17303_42282# a_21613_42308# 0.061584f
C18624 COMP_P a_3754_38470# 4.61e-19
C18625 a_9313_44734# a_19700_43370# 0.001757f
C18626 a_13351_46090# CLK 4.09e-21
C18627 a_742_44458# a_2905_42968# 0.15065f
C18628 a_11341_43940# a_14021_43940# 3.06514f
C18629 a_n967_45348# a_n1630_35242# 0.03295f
C18630 a_11967_42832# a_8685_43396# 0.005728f
C18631 a_n2017_45002# a_1606_42308# 0.04498f
C18632 a_n913_45002# a_1149_42558# 4.87e-21
C18633 a_n1059_45260# a_1221_42558# 1.28e-19
C18634 a_9672_43914# a_9801_43940# 0.062574f
C18635 a_5495_43940# a_n97_42460# 3.76e-20
C18636 a_n1549_44318# a_n1557_42282# 4.58e-21
C18637 a_1414_42308# a_1756_43548# 6.51e-20
C18638 a_949_44458# a_2075_43172# 1.09e-20
C18639 a_2779_44458# a_1847_42826# 1.85e-21
C18640 a_11827_44484# a_5534_30871# 2.07e-22
C18641 a_14673_44172# a_14955_43396# 2.24e-22
C18642 a_17957_46116# VDD 0.138777f
C18643 a_n699_43396# a_685_42968# 3.03e-20
C18644 a_895_43940# a_458_43396# 6.21e-19
C18645 a_453_43940# a_1568_43370# 1.29e-19
C18646 a_n2293_42834# a_5837_43172# 1.46e-19
C18647 a_13249_42308# a_15037_45618# 1.93e-21
C18648 a_14495_45572# a_14033_45822# 3.98e-20
C18649 a_12861_44030# a_20974_43370# 1.38e-19
C18650 a_584_46384# a_n1557_42282# 0.032459f
C18651 a_n971_45724# a_n998_43396# 1.52e-19
C18652 a_167_45260# a_n2661_44458# 4.36e-19
C18653 a_n452_45724# a_n1059_45260# 2.74e-19
C18654 a_n863_45724# a_n913_45002# 0.565852f
C18655 a_20205_31679# a_413_45260# 0.034773f
C18656 a_n2472_45546# en_comp 5.76e-19
C18657 a_n2661_45546# a_n967_45348# 0.001666f
C18658 a_12549_44172# a_20269_44172# 0.049822f
C18659 a_8049_45260# a_15415_45028# 2.92e-20
C18660 a_10586_45546# a_9482_43914# 1.67e-20
C18661 a_11823_42460# a_15765_45572# 1.14e-19
C18662 a_11322_45546# a_8696_44636# 6e-19
C18663 a_11415_45002# a_8975_43940# 6.59e-20
C18664 a_n755_45592# a_n2661_45010# 0.01648f
C18665 a_n2956_38216# a_n2956_37592# 0.103811f
C18666 a_n2442_46660# a_n2661_42282# 7.91e-20
C18667 a_13661_43548# a_13483_43940# 0.057042f
C18668 a_16327_47482# a_18797_44260# 1.19e-19
C18669 a_n2293_45546# a_n2810_45028# 8.06e-21
C18670 a_310_45028# a_n2293_45010# 2.43e-21
C18671 a_n1435_47204# a_1123_46634# 6.22e-20
C18672 a_20990_47178# a_19321_45002# 1.58e-19
C18673 a_20894_47436# a_19594_46812# 7.48e-20
C18674 a_13507_46334# a_13747_46662# 0.049663f
C18675 a_n1741_47186# a_7715_46873# 2.98e-19
C18676 a_n443_46116# a_3524_46660# 0.049574f
C18677 a_2905_45572# a_3877_44458# 6.4e-20
C18678 a_3160_47472# a_3221_46660# 8.54e-19
C18679 a_n4064_39072# C2_P_btm 1.14e-20
C18680 a_18597_46090# a_20916_46384# 6.92e-19
C18681 VDAC_Pi VDAC_P 2.7e-19
C18682 a_n4064_38528# EN_VIN_BSTR_P 0.032853f
C18683 a_2063_45854# a_4955_46873# 0.002567f
C18684 a_15507_47210# a_n743_46660# 0.003069f
C18685 a_4883_46098# a_5807_45002# 1.76125f
C18686 a_n3420_39616# VDD 0.568506f
C18687 a_20447_31679# a_22459_39145# 2.66e-20
C18688 a_19479_31679# a_22469_39537# 3.29e-20
C18689 a_10949_43914# a_10341_42308# 1.01e-22
C18690 a_10807_43548# a_10922_42852# 0.010566f
C18691 a_18184_42460# a_21887_42336# 1.63e-19
C18692 a_19963_31679# a_22521_39511# 2.93e-20
C18693 a_10057_43914# a_10723_42308# 2.38e-19
C18694 a_n2293_43922# a_n784_42308# 1.67292f
C18695 a_3626_43646# a_9145_43396# 9.28e-20
C18696 a_16020_45572# VDD 0.077625f
C18697 a_n97_42460# a_16137_43396# 0.134668f
C18698 a_11967_42832# a_15953_42852# 2.76e-20
C18699 a_6031_43396# a_6643_43396# 3.82e-19
C18700 a_2479_44172# a_3059_42968# 7.19e-19
C18701 a_n356_44636# a_5932_42308# 0.040714f
C18702 a_n971_45724# a_8495_42852# 1.66e-19
C18703 a_8049_45260# a_19279_43940# 2.89e-20
C18704 a_5937_45572# a_6756_44260# 0.010335f
C18705 a_12861_44030# a_18599_43230# 7.75e-20
C18706 a_6812_45938# a_6298_44484# 1.87e-20
C18707 a_n863_45724# a_556_44484# 0.002594f
C18708 a_2382_45260# a_3537_45260# 0.250657f
C18709 a_n1059_45260# a_8953_45002# 8.21e-22
C18710 a_3483_46348# a_15682_43940# 0.261013f
C18711 a_n1613_43370# a_n1379_43218# 0.001903f
C18712 a_10227_46804# a_13460_43230# 0.243111f
C18713 a_2680_45002# a_3429_45260# 4.16e-19
C18714 a_15903_45785# a_16405_45348# 4.53e-20
C18715 a_8162_45546# a_5343_44458# 7.23e-21
C18716 a_2711_45572# a_18443_44721# 2.09e-20
C18717 a_n2109_47186# a_5066_45546# 0.02651f
C18718 a_n971_45724# a_3873_46454# 6.84e-19
C18719 a_10428_46928# a_10554_47026# 0.181217f
C18720 a_9863_46634# a_6755_46942# 0.014818f
C18721 a_7411_46660# a_8035_47026# 9.73e-19
C18722 a_10467_46802# a_10623_46897# 0.107482f
C18723 a_10150_46912# a_10249_46116# 0.066949f
C18724 a_5257_43370# a_6682_46660# 1.27e-19
C18725 a_n237_47217# a_526_44458# 0.198088f
C18726 a_19594_46812# a_20411_46873# 1.02e-20
C18727 a_19321_45002# a_20273_46660# 0.001516f
C18728 a_7715_46873# a_7832_46660# 0.157972f
C18729 a_12861_44030# a_12594_46348# 0.43362f
C18730 a_4883_46098# a_3699_46348# 2.14e-19
C18731 a_104_43370# a_196_42282# 4.54e-20
C18732 a_n97_42460# a_n784_42308# 0.006645f
C18733 a_5649_42852# a_10518_42984# 7.51e-21
C18734 a_n1917_43396# a_n1630_35242# 3.12e-20
C18735 a_4361_42308# a_10991_42826# 2.13e-19
C18736 a_15493_43940# a_15051_42282# 1.93e-19
C18737 a_15743_43084# a_19164_43230# 0.0353f
C18738 a_743_42282# a_12545_42858# 8.12e-20
C18739 a_19268_43646# a_19339_43156# 0.001878f
C18740 a_742_44458# VDD 1.3845f
C18741 a_n2661_43370# a_4743_44484# 0.001974f
C18742 a_21359_45002# a_20193_45348# 3.23e-20
C18743 a_11827_44484# a_11691_44458# 0.881979f
C18744 a_16327_47482# a_20712_42282# 0.030215f
C18745 a_1423_45028# a_n356_44636# 2.19e-21
C18746 a_3232_43370# a_n2661_43922# 0.197944f
C18747 a_6171_45002# a_n2661_42834# 0.001465f
C18748 a_13507_46334# a_4958_30871# 6.72e-21
C18749 a_4185_45028# a_13678_32519# 0.037732f
C18750 SMPL_ON_P a_n4064_38528# 9.15e-21
C18751 a_18587_45118# a_18545_45144# 7.47e-21
C18752 a_n133_46660# a_997_45618# 3.7e-20
C18753 a_2107_46812# a_n863_45724# 3.26e-20
C18754 a_n2293_46634# a_n23_45546# 2.45e-19
C18755 a_19692_46634# a_18819_46122# 2.56e-19
C18756 a_19466_46812# a_18985_46122# 0.033782f
C18757 a_n881_46662# a_4880_45572# 2.99e-19
C18758 a_12465_44636# a_13249_42308# 0.541909f
C18759 a_4883_46098# a_15143_45578# 5.67e-21
C18760 a_n743_46660# a_2957_45546# 2.2e-20
C18761 a_n2438_43548# a_1848_45724# 1.12e-20
C18762 a_171_46873# a_n755_45592# 1.47e-22
C18763 a_33_46660# a_n357_42282# 9.6e-20
C18764 a_9863_46634# a_8049_45260# 1.3e-20
C18765 a_15227_44166# a_19335_46494# 0.024137f
C18766 a_19333_46634# a_19553_46090# 0.001209f
C18767 a_13885_46660# a_13759_46122# 0.002423f
C18768 a_15368_46634# a_6945_45028# 3.82e-19
C18769 a_n2840_46090# a_n2472_46090# 7.52e-19
C18770 a_765_45546# a_8016_46348# 6.75e-20
C18771 a_383_46660# a_n1099_45572# 9.12e-21
C18772 a_8270_45546# a_526_44458# 0.007312f
C18773 a_14035_46660# a_13351_46090# 1.44e-19
C18774 a_3090_45724# a_10809_44734# 0.002539f
C18775 a_13059_46348# a_9290_44172# 2.64e-19
C18776 a_13487_47204# a_14033_45822# 1.36e-20
C18777 a_12861_44030# a_15037_45618# 1.43e-20
C18778 a_4361_42308# a_17303_42282# 0.050893f
C18779 a_4190_30871# a_18220_42308# 0.00137f
C18780 a_13003_42852# a_13291_42460# 2.39e-20
C18781 a_8037_42858# a_8325_42308# 5.53e-19
C18782 a_7871_42858# a_8791_42308# 0.004922f
C18783 a_743_42282# a_19332_42282# 0.006778f
C18784 a_n2293_42282# a_n3674_37592# 0.08084f
C18785 a_21115_43940# VDD 0.145936f
C18786 a_4185_45028# a_6123_31319# 0.068372f
C18787 a_18479_45785# a_10341_43396# 0.038969f
C18788 a_n1059_45260# a_3626_43646# 0.025708f
C18789 a_n2017_45002# a_3539_42460# 0.042001f
C18790 a_n310_47243# VDD 2.4e-19
C18791 a_n310_47570# DATA[0] 6.14e-19
C18792 a_1307_43914# a_11173_43940# 3.43e-19
C18793 a_17339_46660# a_18548_42308# 1.37e-19
C18794 a_2274_45254# a_1568_43370# 1.33e-21
C18795 a_4223_44672# a_3905_42865# 0.019153f
C18796 a_n2267_44484# a_n4318_39768# 4.62e-19
C18797 a_17613_45144# a_17737_43940# 7.01e-20
C18798 a_3357_43084# a_7287_43370# 7.22e-20
C18799 a_22731_47423# EN_OFFSET_CAL 1.57e-20
C18800 a_n357_42282# a_18817_42826# 0.008235f
C18801 a_n443_42852# a_12895_43230# 1.14e-19
C18802 a_n2956_39304# a_n2840_42282# 2.99e-20
C18803 a_8696_44636# a_16409_43396# 4.05e-20
C18804 a_15861_45028# a_16547_43609# 4.56e-21
C18805 a_21588_30879# a_22609_37990# 1.43e-20
C18806 a_n699_43396# a_3600_43914# 1.42e-19
C18807 a_10428_46928# a_2437_43646# 3.53e-20
C18808 a_13507_46334# a_18911_45144# 1.16e-20
C18809 a_18597_46090# a_21101_45002# 0.033595f
C18810 a_n743_46660# a_9482_43914# 7.74e-21
C18811 a_19553_46090# a_20062_46116# 2.6e-19
C18812 a_n2497_47436# a_n356_44636# 0.019387f
C18813 a_3147_46376# a_2711_45572# 7.31e-20
C18814 a_3524_46660# a_3537_45260# 1.28e-20
C18815 a_n2293_46098# a_6428_45938# 5.88e-21
C18816 a_3221_46660# a_413_45260# 9.19e-19
C18817 a_11415_45002# a_10193_42453# 0.024787f
C18818 a_18479_47436# a_11827_44484# 0.035345f
C18819 a_5066_45546# a_8062_46155# 9.9e-19
C18820 a_4791_45118# a_5518_44484# 2.27e-19
C18821 a_4883_46098# a_18315_45260# 1.48e-20
C18822 a_3090_45724# a_16211_45572# 7.88e-19
C18823 a_3823_42558# a_7174_31319# 4.88e-21
C18824 a_n3674_38680# a_n4334_39392# 1.52e-19
C18825 a_13575_42558# a_14456_42282# 0.008255f
C18826 a_13070_42354# a_13249_42558# 0.010303f
C18827 a_13678_32519# VREF_GND 0.047887f
C18828 a_n901_43156# VDD 0.475947f
C18829 a_n3674_37592# a_n3565_39590# 4.6e-20
C18830 a_n1630_35242# a_n4209_39590# 0.12484f
C18831 a_9803_42558# a_10149_42308# 0.013377f
C18832 a_20885_46660# SINGLE_ENDED 2.32e-21
C18833 a_5891_43370# a_6293_42852# 0.107308f
C18834 a_20820_30879# C10_N_btm 4.87e-19
C18835 a_11827_44484# a_4190_30871# 3.39e-20
C18836 a_1307_43914# a_13460_43230# 1.02e-20
C18837 a_3232_43370# a_3445_43172# 1.88e-19
C18838 a_10193_42453# a_10533_42308# 0.101629f
C18839 a_n2661_43922# a_4905_42826# 9.3e-21
C18840 a_n2293_43922# a_3080_42308# 0.084673f
C18841 a_21076_30879# C7_N_btm 0.00198f
C18842 a_6109_44484# a_6547_43396# 0.001963f
C18843 a_n2293_42834# a_791_42968# 0.007944f
C18844 a_10057_43914# a_10341_43396# 0.055207f
C18845 a_7499_43078# a_11551_42558# 3.18e-19
C18846 a_21005_45260# a_20556_43646# 2.16e-21
C18847 a_18184_42460# a_13467_32519# 0.022572f
C18848 a_18494_42460# a_19095_43396# 3.48e-20
C18849 a_14537_43396# a_15567_42826# 4.38e-22
C18850 a_20202_43084# RST_Z 7.21e-20
C18851 a_11415_45002# VDD 1.84504f
C18852 a_n1899_43946# a_726_44056# 1.56e-20
C18853 a_2711_45572# a_13249_42308# 0.043493f
C18854 a_768_44030# a_n1761_44111# 2.61e-20
C18855 a_20107_46660# a_20567_45036# 5.96e-22
C18856 a_9290_44172# a_13556_45296# 2.5e-20
C18857 a_17715_44484# a_6171_45002# 5.11e-20
C18858 a_3090_45724# a_5883_43914# 0.132458f
C18859 a_16375_45002# a_16147_45260# 1.01554f
C18860 a_526_44458# a_n2017_45002# 0.028467f
C18861 a_n2312_40392# a_n3674_39768# 0.025146f
C18862 a_n2312_39304# a_n4318_39768# 0.02345f
C18863 a_10903_43370# a_13017_45260# 2.86e-19
C18864 a_12005_46116# a_11963_45334# 1.6e-19
C18865 a_5204_45822# a_1423_45028# 3.01e-21
C18866 a_2324_44458# a_7276_45260# 0.049304f
C18867 a_4646_46812# a_n2293_43922# 8.64e-21
C18868 a_13259_45724# a_18341_45572# 1.51e-19
C18869 a_n1151_42308# a_4842_47243# 8.14e-19
C18870 a_3785_47178# a_n881_46662# 6.74e-19
C18871 a_3815_47204# a_n1613_43370# 0.001154f
C18872 a_n443_46116# a_4842_47570# 0.001342f
C18873 a_4958_30871# a_n923_35174# 0.015856f
C18874 a_16327_47482# a_19386_47436# 3.57e-20
C18875 a_17591_47464# a_18143_47464# 0.003298f
C18876 a_5742_30871# C9_N_btm 0.003249f
C18877 a_14311_47204# a_4883_46098# 1.02e-20
C18878 a_11599_46634# a_13507_46334# 0.259318f
C18879 a_n3565_38216# a_n3690_38304# 0.247167f
C18880 a_n4334_38304# a_n3420_37984# 0.004718f
C18881 a_n4209_38216# a_n2946_37984# 0.022779f
C18882 a_10533_42308# VDD 0.216201f
C18883 a_5934_30871# VIN_N 0.009408f
C18884 a_13717_47436# a_22223_47212# 0.00262f
C18885 a_12861_44030# a_12465_44636# 0.242761f
C18886 a_6123_31319# VREF_GND 0.00207f
C18887 a_n1177_43370# a_n1557_42282# 4.78e-22
C18888 a_n97_42460# a_3080_42308# 0.353977f
C18889 a_14021_43940# a_10341_43396# 1.5617f
C18890 en_comp a_1239_39043# 0.007802f
C18891 a_3733_45822# VDD 5.25e-19
C18892 a_18079_43940# a_15743_43084# 6.36e-20
C18893 a_18451_43940# a_18525_43370# 3.66e-19
C18894 a_15493_43396# a_17324_43396# 0.047612f
C18895 a_n3674_39768# a_n2840_42826# 0.001686f
C18896 a_11967_42832# a_17333_42852# 0.14149f
C18897 a_742_44458# a_n784_42308# 4.46e-20
C18898 a_15682_43940# a_16664_43396# 0.001235f
C18899 a_1115_44172# a_791_42968# 7.5e-19
C18900 a_16327_47482# a_20556_43646# 0.014087f
C18901 a_21188_45572# a_22959_45572# 8.11e-21
C18902 a_19692_46634# a_11341_43940# 0.06f
C18903 a_4646_46812# a_n97_42460# 0.016161f
C18904 a_n863_45724# a_n2661_44458# 0.091002f
C18905 a_2711_45572# a_17613_45144# 1.8e-20
C18906 a_n2293_45546# a_n2129_44697# 3.68e-19
C18907 a_15861_45028# a_6171_45002# 0.09425f
C18908 a_n2293_46634# a_7287_43370# 0.016986f
C18909 a_584_46384# a_3935_42891# 4.23e-20
C18910 a_5807_45002# a_8685_43396# 9.36e-20
C18911 a_526_44458# a_n89_44484# 1.64e-20
C18912 a_15682_46116# a_17061_44734# 1.05e-20
C18913 a_n443_42852# a_11827_44484# 1.48e-19
C18914 a_4808_45572# a_n2661_43370# 2.36e-19
C18915 a_n1151_42308# a_685_42968# 9.34e-22
C18916 a_21363_45546# a_20447_31679# 5.34e-20
C18917 C2_P_btm VDD 0.268945f
C18918 a_11530_34132# VIN_N 1.547f
C18919 a_16327_47482# a_19551_46910# 1.05e-19
C18920 a_n1925_46634# a_8145_46902# 0.005351f
C18921 a_5807_45002# a_6682_46660# 6.46e-19
C18922 a_12549_44172# a_11735_46660# 1.77e-19
C18923 a_12891_46348# a_11813_46116# 1.48e-19
C18924 a_3815_47204# a_n2293_46098# 2.35e-20
C18925 a_11309_47204# a_11901_46660# 0.001315f
C18926 a_n881_46662# a_3090_45724# 0.107805f
C18927 a_2443_46660# a_3877_44458# 2.31e-19
C18928 a_3177_46902# a_3055_46660# 3.16e-19
C18929 a_2107_46812# a_5072_46660# 8.97e-19
C18930 a_n2109_47186# a_5068_46348# 1.71e-20
C18931 a_n2661_46634# a_10428_46928# 0.052586f
C18932 a_584_46384# a_472_46348# 0.31609f
C18933 a_1209_47178# a_1138_42852# 1.18e-20
C18934 a_1239_47204# a_1176_45822# 4.07e-21
C18935 a_2063_45854# a_376_46348# 3.28e-20
C18936 EN_VIN_BSTR_P VREF_GND 0.85739f
C18937 a_n1741_47186# a_4419_46090# 4.26e-20
C18938 a_n971_45724# a_2804_46116# 1.43e-19
C18939 a_n237_47217# a_2521_46116# 0.039248f
C18940 a_n1151_42308# a_n1991_46122# 0.027139f
C18941 a_n743_46660# a_7715_46873# 0.003347f
C18942 a_11599_46634# a_20623_46660# 4.44e-20
C18943 a_10227_46804# a_17339_46660# 2.73e-20
C18944 a_17591_47464# a_765_45546# 0.004682f
C18945 C0_P_btm C10_N_btm 0.00154f
C18946 C0_dummy_P_btm C9_N_btm 7.47e-19
C18947 C2_N_btm C5_N_btm 0.138678f
C18948 C3_N_btm C4_N_btm 7.90108f
C18949 C1_N_btm C6_N_btm 0.128559f
C18950 C0_dummy_N_btm C8_N_btm 0.236317f
C18951 C0_N_btm C7_N_btm 0.142187f
C18952 a_12465_44636# a_14180_46812# 0.026945f
C18953 a_3422_30871# a_18057_42282# 3.03e-20
C18954 a_19279_43940# a_13258_32519# 4.56e-21
C18955 a_17433_43396# a_4190_30871# 4.55e-21
C18956 a_8685_43396# a_10518_42984# 4.24e-19
C18957 a_2982_43646# a_21356_42826# 0.005304f
C18958 a_15743_43084# a_14209_32519# 4.59e-21
C18959 a_n97_42460# a_7309_43172# 0.002468f
C18960 a_1568_43370# a_945_42968# 1.47e-20
C18961 a_3080_42308# a_3935_43218# 4.27e-20
C18962 a_15595_45028# a_11691_44458# 2.85e-20
C18963 a_n357_42282# a_15682_43940# 1.36e-19
C18964 a_8199_44636# a_8791_43396# 1.65e-19
C18965 a_17339_46660# a_19177_43646# 2.77e-19
C18966 a_n1613_43370# a_n4318_38216# 1.48e-19
C18967 a_n1059_45260# a_17767_44458# 2.41e-19
C18968 a_3537_45260# a_5343_44458# 0.378482f
C18969 a_8191_45002# a_n2661_44458# 0.001306f
C18970 a_5147_45002# a_4223_44672# 0.047867f
C18971 a_4558_45348# a_n699_43396# 4.82e-22
C18972 a_8696_44636# a_16241_44734# 0.004986f
C18973 a_2107_46812# a_1431_46436# 1.17e-19
C18974 a_5807_45002# a_11608_46482# 5.69e-19
C18975 a_10428_46928# a_8199_44636# 5.81e-19
C18976 a_6575_47204# a_6598_45938# 1.53e-21
C18977 a_n1151_42308# a_7499_43078# 6.25e-20
C18978 a_n443_46116# a_4880_45572# 0.048165f
C18979 a_n2312_39304# a_n2956_38216# 0.060648f
C18980 a_12861_44030# a_2711_45572# 0.104124f
C18981 a_2063_45854# a_8746_45002# 0.058531f
C18982 a_20916_46384# a_8049_45260# 0.003776f
C18983 a_n1925_46634# a_5066_45546# 0.195997f
C18984 a_n2661_46098# a_n1545_46494# 0.004305f
C18985 a_14209_32519# a_1606_42308# 1.87e-20
C18986 a_n1423_42826# a_n3674_37592# 4.62e-20
C18987 a_n1533_42852# a_n4318_38216# 4.39e-19
C18988 a_n984_44318# VDD 0.281427f
C18989 a_4361_42308# a_2713_42308# 2.85e-20
C18990 a_n901_43156# a_n784_42308# 4.44e-19
C18991 a_n13_43084# a_n473_42460# 2.62e-19
C18992 a_10341_43396# a_15764_42576# 7.76e-21
C18993 a_12281_43396# a_13657_42558# 1.55e-21
C18994 a_13635_43156# a_13291_42460# 0.004222f
C18995 a_n1853_43023# a_n1630_35242# 1.28e-19
C18996 a_743_42282# a_5379_42460# 0.013947f
C18997 a_18287_44626# a_9313_44734# 6.97e-21
C18998 a_12607_44458# a_n2661_42834# 5.21e-19
C18999 a_21005_45260# a_20980_44850# 5.39e-19
C19000 a_11827_44484# a_18753_44484# 0.001286f
C19001 a_n755_45592# a_5649_42852# 0.02386f
C19002 a_21076_30879# COMP_P 1.25e-19
C19003 a_2553_47502# VDD 0.150286f
C19004 a_8975_43940# a_n2661_43922# 0.11532f
C19005 a_18479_45785# a_n97_42460# 0.072469f
C19006 a_n2293_42834# a_3905_42865# 0.039227f
C19007 a_9482_43914# a_11750_44172# 0.020902f
C19008 a_18184_42460# a_22315_44484# 1.48e-22
C19009 a_18494_42460# a_3422_30871# 7.81e-19
C19010 a_9290_44172# a_11554_42852# 0.031758f
C19011 a_1239_47204# DATA[0] 2.02e-19
C19012 a_1209_47178# DATA[1] 0.076054f
C19013 a_20193_45348# a_19279_43940# 0.021458f
C19014 a_n2661_43370# a_1414_42308# 9.45e-21
C19015 a_11691_44458# a_18005_44484# 0.001888f
C19016 a_2711_45572# a_19700_43370# 0.016505f
C19017 a_13507_46334# a_13348_45260# 7.06e-20
C19018 a_11901_46660# a_10490_45724# 1.82e-20
C19019 a_20820_30879# a_20205_31679# 0.087297f
C19020 a_n1613_43370# a_2382_45260# 2e-21
C19021 a_20708_46348# a_6945_45028# 0.002334f
C19022 a_20075_46420# a_10809_44734# 2.78e-20
C19023 a_8349_46414# a_8034_45724# 0.05863f
C19024 a_14180_46812# a_2711_45572# 2.03e-20
C19025 a_11735_46660# a_11525_45546# 1.78e-20
C19026 a_11813_46116# a_11322_45546# 3.46e-20
C19027 a_22591_46660# a_20692_30879# 0.001224f
C19028 a_22612_30879# a_2437_43646# 9.37e-20
C19029 a_20202_43084# a_21167_46155# 2.55e-19
C19030 a_10227_46804# a_1307_43914# 0.081555f
C19031 a_2351_42308# a_5934_30871# 1.01e-20
C19032 a_3905_42558# a_4921_42308# 4.04e-22
C19033 a_n784_42308# a_10533_42308# 2.26e-20
C19034 a_9885_43646# VDD 0.190473f
C19035 a_3823_42558# a_5932_42308# 4.34e-21
C19036 a_5379_42460# a_5755_42308# 0.004559f
C19037 a_n2472_43914# a_n3674_39768# 0.162742f
C19038 a_n2065_43946# a_n4318_39768# 3.52e-21
C19039 a_1414_42308# a_2998_44172# 0.447595f
C19040 a_11967_42832# a_13483_43940# 1.65e-20
C19041 a_n357_42282# a_5934_30871# 0.001326f
C19042 a_17517_44484# a_19862_44208# 2.23e-19
C19043 a_n1059_45260# a_8037_42858# 0.048776f
C19044 a_n913_45002# a_7765_42852# 4.6e-19
C19045 a_n755_45592# a_7963_42308# 0.003087f
C19046 a_n2956_39304# a_n2302_39866# 2.06e-19
C19047 a_10193_42453# a_20256_42852# 4.84e-19
C19048 a_13259_45724# a_15803_42450# 7.39e-19
C19049 a_5891_43370# a_7499_43940# 7.45e-20
C19050 a_742_44458# a_3080_42308# 5.11e-20
C19051 a_12251_46660# VDD 0.195617f
C19052 a_2479_44172# a_895_43940# 0.318312f
C19053 a_2127_44172# a_2675_43914# 0.090298f
C19054 a_10057_43914# a_n97_42460# 4.56e-21
C19055 a_n699_43396# a_1756_43548# 0.004876f
C19056 a_4223_44672# a_4093_43548# 1.33e-19
C19057 a_327_44734# a_685_42968# 4.03e-22
C19058 a_16327_47482# a_20980_44850# 0.012339f
C19059 a_8049_45260# a_10210_45822# 0.01041f
C19060 a_13259_45724# a_10193_42453# 0.284945f
C19061 a_768_44030# a_5708_44484# 0.003906f
C19062 a_n881_46662# a_14815_43914# 3.35e-21
C19063 a_12861_44030# a_22485_44484# 2.25e-19
C19064 a_n2293_46634# a_n23_44458# 2.19e-20
C19065 a_17957_46116# a_18479_45785# 7.94e-19
C19066 a_18819_46122# a_18175_45572# 3.23e-19
C19067 a_18189_46348# a_18341_45572# 0.001747f
C19068 a_n2293_46098# a_2382_45260# 1.97e-20
C19069 a_n443_46116# a_453_43940# 0.004377f
C19070 a_167_45260# a_n1059_45260# 1.04e-20
C19071 a_5497_46414# a_3357_43084# 0.005427f
C19072 a_n2438_43548# a_n2012_44484# 0.009651f
C19073 a_7_45899# a_n443_42852# 5.72e-19
C19074 a_n755_45592# a_1260_45572# 0.001566f
C19075 a_997_45618# a_1176_45572# 0.007688f
C19076 a_18597_46090# a_20766_44850# 0.00611f
C19077 a_n784_42308# C2_P_btm 0.005178f
C19078 a_n746_45260# a_n1435_47204# 5.74e-19
C19079 a_4007_47204# a_4700_47436# 0.010942f
C19080 a_3785_47178# a_n443_46116# 0.040847f
C19081 a_n1151_42308# a_5129_47502# 0.002765f
C19082 a_3815_47204# a_4791_45118# 6.07e-20
C19083 a_3381_47502# a_4915_47217# 9.99e-20
C19084 a_7174_31319# a_1177_38525# 1.57e-19
C19085 a_n1741_47186# a_11599_46634# 0.164599f
C19086 a_1239_39587# a_1343_38525# 0.011696f
C19087 a_n3565_39590# a_n2302_39072# 8.95e-20
C19088 a_5742_30871# a_n3420_37440# 0.004591f
C19089 a_20256_42852# VDD 0.001626f
C19090 a_11967_42832# a_13678_32519# 1.08e-19
C19091 a_20679_44626# a_21487_43396# 5.88e-19
C19092 a_9313_44734# a_9127_43156# 0.001322f
C19093 a_18494_42460# a_18504_43218# 8.04e-19
C19094 a_n2017_45002# a_16104_42674# 0.004413f
C19095 a_20835_44721# a_20556_43646# 9.48e-20
C19096 a_18287_44626# a_18599_43230# 2.95e-19
C19097 a_18374_44850# a_18249_42858# 3.5e-21
C19098 a_14021_43940# a_n97_42460# 0.002657f
C19099 a_13259_45724# VDD 2.41738f
C19100 a_n2293_42834# a_n961_42308# 0.001885f
C19101 a_n356_44636# a_15567_42826# 1.19e-20
C19102 a_n2661_42834# a_3681_42891# 1.08e-21
C19103 a_n2661_43922# a_2905_42968# 2.14e-21
C19104 a_8333_44056# a_8147_43396# 0.011009f
C19105 a_2711_45572# a_11787_45002# 2.49e-20
C19106 a_3638_45822# a_3232_43370# 1.51e-20
C19107 a_3090_45724# a_2889_44172# 6.33e-21
C19108 a_n2293_45546# a_45_45144# 5.47e-19
C19109 a_6472_45840# a_6709_45028# 8.56e-19
C19110 a_6598_45938# a_5205_44484# 5.22e-19
C19111 a_6511_45714# a_7229_43940# 6.9e-21
C19112 a_8049_45260# a_21101_45002# 9.79e-21
C19113 a_13259_45724# a_14309_45348# 3.49e-19
C19114 a_1823_45246# a_3363_44484# 0.046566f
C19115 a_17478_45572# a_18341_45572# 5.87e-19
C19116 a_n1076_46494# a_n2661_43922# 1.73e-21
C19117 a_11823_42460# a_n913_45002# 0.281323f
C19118 a_17339_46660# a_18579_44172# 0.016577f
C19119 a_15765_45572# a_16789_45572# 2.36e-20
C19120 a_n1613_43370# a_n1655_43396# 0.001903f
C19121 a_2324_44458# a_13720_44458# 1.95e-20
C19122 a_14840_46494# a_15004_44636# 2.04e-21
C19123 a_3503_45724# a_1423_45028# 5.37e-21
C19124 a_19321_45002# a_19319_43548# 3.41e-19
C19125 a_n4064_37440# C1_P_btm 0.031032f
C19126 a_n2840_46634# a_n2956_39768# 0.156182f
C19127 a_n881_46662# a_3699_46634# 0.001985f
C19128 a_n1613_43370# a_3524_46660# 0.28004f
C19129 a_3754_38802# VDD 0.002173f
C19130 a_7754_38968# RST_Z 9.75e-19
C19131 a_13747_46662# a_n743_46660# 0.042998f
C19132 a_n443_46116# a_3090_45724# 0.011392f
C19133 a_6151_47436# a_12816_46660# 6.67e-20
C19134 a_4915_47217# a_15009_46634# 1.25e-20
C19135 a_22469_39537# a_22609_37990# 0.490939f
C19136 a_10227_46804# a_10467_46802# 0.678578f
C19137 a_2982_43646# a_20749_43396# 0.00204f
C19138 a_6031_43396# a_4361_42308# 3.96e-20
C19139 a_n809_44244# a_n327_42558# 7.98e-21
C19140 a_175_44278# a_196_42282# 4.29e-21
C19141 a_n467_45028# VDD 0.385804f
C19142 a_10341_43396# a_13943_43396# 7.41e-20
C19143 a_n1557_42282# a_n1991_42858# 1.42e-19
C19144 a_7287_43370# a_743_42282# 2.89e-20
C19145 a_n1899_43946# a_n1630_35242# 1.8e-21
C19146 a_10807_43548# a_11554_42852# 0.002521f
C19147 a_15095_43370# a_16547_43609# 2.35e-21
C19148 a_9313_44734# a_17124_42282# 4.54e-20
C19149 a_13661_43548# a_18083_42858# 0.009269f
C19150 a_10193_42453# a_n2661_43922# 0.025533f
C19151 a_15765_45572# a_14539_43914# 1.95e-20
C19152 a_8746_45002# a_n2661_42834# 1.37e-19
C19153 a_2437_43646# a_11827_44484# 0.013953f
C19154 a_21513_45002# a_22223_45036# 7.29e-20
C19155 a_10227_46804# a_13003_42852# 0.012229f
C19156 a_19692_46634# a_10341_43396# 0.022785f
C19157 a_8953_45546# a_9801_43940# 9.11e-19
C19158 a_5147_45002# a_n2293_42834# 1.41e-21
C19159 a_n357_42282# a_20512_43084# 0.005311f
C19160 a_1667_45002# a_n2661_43370# 0.01f
C19161 a_n2661_45546# a_n1899_43946# 1.44e-21
C19162 a_3357_43084# a_21005_45260# 1.78e-20
C19163 a_19479_31679# a_21101_45002# 5.63e-19
C19164 a_8696_44636# a_12883_44458# 0.002403f
C19165 a_3232_43370# a_5837_45028# 0.01175f
C19166 a_16333_45814# a_16112_44458# 4.95e-21
C19167 a_3090_45724# a_14621_43646# 1.89e-20
C19168 a_n1151_42308# a_n1329_42308# 0.167748f
C19169 a_11599_46634# a_10586_45546# 1.89e-19
C19170 a_12549_44172# a_2324_44458# 0.506903f
C19171 a_n237_47217# a_n452_45724# 6.22e-21
C19172 a_n2661_46098# a_n901_46420# 0.054328f
C19173 a_1983_46706# a_1823_45246# 0.005043f
C19174 a_2107_46812# a_2202_46116# 0.008835f
C19175 a_10428_46928# a_765_45546# 0.003387f
C19176 a_15368_46634# a_15559_46634# 0.022471f
C19177 a_n1925_46634# a_5068_46348# 4.81e-20
C19178 a_n743_46660# a_4419_46090# 0.032595f
C19179 a_1431_47204# a_n2661_45546# 3.64e-21
C19180 a_11901_46660# a_12156_46660# 0.06121f
C19181 a_11186_47026# a_10933_46660# 4.61e-19
C19182 a_3090_45724# a_17609_46634# 9.39e-20
C19183 a_14976_45028# a_16292_46812# 1.49e-19
C19184 a_948_46660# a_167_45260# 8.29e-21
C19185 a_n746_45260# a_380_45546# 0.003276f
C19186 a_n971_45724# a_n1099_45572# 0.508925f
C19187 a_5807_45002# a_11387_46155# 0.005659f
C19188 a_n2497_47436# a_3503_45724# 4.5e-21
C19189 a_9313_44734# CLK 9.52e-20
C19190 a_n97_42460# a_15764_42576# 0.174403f
C19191 a_6031_43396# a_6761_42308# 3.22e-19
C19192 a_13635_43156# a_13460_43230# 0.234322f
C19193 a_13113_42826# a_5534_30871# 0.024339f
C19194 a_16137_43396# a_20256_42852# 1.75e-20
C19195 a_2982_43646# a_8685_42308# 1.03e-19
C19196 a_n2661_43922# VDD 0.611934f
C19197 a_3681_42891# a_n2293_42282# 0.012859f
C19198 a_13259_45724# a_16137_43396# 0.038525f
C19199 a_9290_44172# a_10991_42826# 0.045863f
C19200 a_4185_45028# a_18083_42858# 4.75e-20
C19201 a_n755_45592# a_8685_43396# 0.001034f
C19202 a_n443_42852# a_8147_43396# 0.060401f
C19203 a_2382_45260# a_2675_43914# 1.8e-20
C19204 a_3065_45002# a_2479_44172# 5.13e-21
C19205 a_n2956_39304# a_n3674_39304# 0.029162f
C19206 a_5343_44458# a_8701_44490# 8.47e-20
C19207 a_3357_43084# a_5841_44260# 2.14e-21
C19208 a_2324_44458# a_5111_42852# 2.92e-22
C19209 a_n2810_45028# a_n4318_39768# 0.027945f
C19210 a_18175_45572# a_11341_43940# 1.54e-21
C19211 a_16327_47482# a_3357_43084# 0.114502f
C19212 a_2063_45854# a_3232_43370# 0.056568f
C19213 a_15227_44166# a_19240_46482# 2.61e-19
C19214 a_11309_47204# a_8696_44636# 2.99e-21
C19215 a_5815_47464# a_413_45260# 4.35e-19
C19216 a_4883_46098# a_20107_45572# 5.13e-20
C19217 a_18479_47436# a_21350_45938# 1.16e-19
C19218 a_7920_46348# a_8199_44636# 5.3e-19
C19219 a_6419_46155# a_5937_45572# 1.25e-20
C19220 a_8016_46348# a_8349_46414# 0.232167f
C19221 a_22959_46660# a_22959_46124# 0.026152f
C19222 a_n237_47217# a_8953_45002# 9.06e-19
C19223 a_n443_46116# a_2274_45254# 0.041907f
C19224 a_4791_45118# a_2382_45260# 3.36e-20
C19225 a_13507_46334# a_20841_45814# 3.6e-20
C19226 a_3483_46348# a_10903_43370# 0.404121f
C19227 a_21076_30879# a_10809_44734# 0.002069f
C19228 a_16588_47582# a_2437_43646# 0.00737f
C19229 a_3080_42308# C2_P_btm 0.108823f
C19230 a_n3674_39304# a_n3565_39304# 0.128699f
C19231 a_n447_43370# VDD 0.204801f
C19232 a_17595_43084# a_17303_42282# 1.12e-19
C19233 a_17701_42308# a_4958_30871# 0.007602f
C19234 a_n2104_42282# a_n3674_38216# 0.155459f
C19235 a_n2472_42282# a_n4318_37592# 0.030006f
C19236 a_n4318_38216# a_n1736_42282# 1.83e-19
C19237 a_n3674_38680# COMP_P 2.55e-20
C19238 a_8495_42852# a_8515_42308# 2.45e-19
C19239 a_n4318_38680# a_n4334_39392# 1.76e-19
C19240 a_4185_45028# a_22775_42308# 0.023674f
C19241 a_2107_46812# DATA[3] 2.5e-21
C19242 a_17970_44736# a_18079_43940# 4.64e-19
C19243 a_20159_44458# a_20397_44484# 0.007399f
C19244 a_n2956_39304# a_5742_30871# 5.51e-21
C19245 a_13259_45724# a_n784_42308# 4.14e-20
C19246 a_5883_43914# a_9248_44260# 0.003192f
C19247 a_n2661_43922# a_5495_43940# 2.85e-20
C19248 a_n2661_42834# a_5663_43940# 0.01057f
C19249 a_20679_44626# a_21398_44850# 0.086708f
C19250 a_20835_44721# a_20980_44850# 0.057222f
C19251 a_20640_44752# a_3422_30871# 0.006762f
C19252 a_1307_43914# a_9396_43370# 4.91e-20
C19253 a_n2293_42834# a_4093_43548# 0.00711f
C19254 a_18184_42460# a_19319_43548# 0.032261f
C19255 a_1799_45572# VDD 0.381212f
C19256 a_n357_42282# a_16245_42852# 0.008838f
C19257 a_526_44458# a_4169_42308# 6.81e-19
C19258 a_n2017_45002# a_18783_43370# 1.92e-20
C19259 a_n1059_45260# a_18525_43370# 0.001977f
C19260 a_13351_46090# a_13527_45546# 4.9e-19
C19261 a_12594_46348# a_13904_45546# 0.077346f
C19262 a_14493_46090# a_11823_42460# 2.22e-20
C19263 a_18189_46348# a_10193_42453# 1.46e-20
C19264 a_5937_45572# a_10907_45822# 1.68e-21
C19265 a_19333_46634# a_413_45260# 1.81e-20
C19266 a_526_44458# a_4099_45572# 0.063912f
C19267 a_2324_44458# a_11525_45546# 0.005847f
C19268 a_4817_46660# a_5009_45028# 5.42e-22
C19269 a_10903_43370# a_14495_45572# 4.3e-19
C19270 a_4915_47217# a_14112_44734# 4.38e-19
C19271 a_11901_46660# a_6171_45002# 1.49e-20
C19272 a_3090_45724# a_3537_45260# 0.198803f
C19273 a_n1613_43370# a_5343_44458# 0.03714f
C19274 a_11453_44696# a_16979_44734# 0.009676f
C19275 a_20841_46902# a_20623_45572# 3.35e-20
C19276 a_21188_46660# a_20107_45572# 2.91e-21
C19277 a_20107_46660# a_20528_45572# 1.27e-20
C19278 a_20623_46660# a_20841_45814# 1.29e-20
C19279 a_21363_46634# a_20273_45572# 2.68e-21
C19280 a_11415_45002# a_18479_45785# 0.047896f
C19281 a_8270_45546# a_8953_45002# 0.004456f
C19282 a_n2661_46634# a_11827_44484# 3.03e-20
C19283 a_5742_30871# a_n3565_39304# 5.51e-21
C19284 a_5932_42308# a_1177_38525# 1.83e-19
C19285 a_18057_42282# a_7174_31319# 2.5e-20
C19286 a_17303_42282# a_21887_42336# 0.001033f
C19287 a_19332_42282# a_13258_32519# 7.57e-19
C19288 a_n3674_38680# a_n3565_37414# 1.14e-20
C19289 a_12594_46348# CLK 1.08e-20
C19290 a_21115_43940# a_14021_43940# 1.8e-20
C19291 en_comp a_n1630_35242# 2.31448f
C19292 a_n913_45002# a_961_42354# 4.8e-20
C19293 a_n1059_45260# a_1149_42558# 1.69e-19
C19294 a_n2017_45002# a_1221_42558# 4.86e-19
C19295 a_5013_44260# a_n97_42460# 1.01e-19
C19296 a_1414_42308# a_1568_43370# 0.01352f
C19297 a_1467_44172# a_1756_43548# 0.100052f
C19298 a_9313_44734# a_19268_43646# 1.06e-20
C19299 a_949_44458# a_1847_42826# 3.24e-19
C19300 a_742_44458# a_2075_43172# 0.002798f
C19301 a_18189_46348# VDD 0.211855f
C19302 a_n1644_44306# a_n4318_39304# 1.35e-19
C19303 a_n3674_39768# a_n2433_43396# 0.002677f
C19304 a_n2293_42834# a_5457_43172# 1.98e-19
C19305 a_n2661_44458# a_7765_42852# 5.2e-21
C19306 a_13249_42308# a_14033_45822# 0.006215f
C19307 a_584_46384# a_766_43646# 0.006798f
C19308 a_12861_44030# a_14401_32519# 2.77e-19
C19309 a_n863_45724# a_n1059_45260# 0.162875f
C19310 a_n2472_45546# a_n2956_37592# 4.88e-19
C19311 a_n2661_45546# en_comp 0.001261f
C19312 a_2324_44458# a_15685_45394# 0.002859f
C19313 a_11823_42460# a_15903_45785# 2.67e-19
C19314 a_n357_42282# a_n2661_45010# 0.017732f
C19315 a_5807_45002# a_13483_43940# 1.27e-19
C19316 a_n2956_38216# a_n2810_45028# 5.73989f
C19317 a_n2293_45546# a_n745_45366# 0.038459f
C19318 a_n1079_45724# a_n913_45002# 2.36e-19
C19319 a_n1099_45572# a_n2293_45010# 0.002597f
C19320 a_n2293_46098# a_5343_44458# 4.66e-20
C19321 a_9241_45822# a_9159_45572# 5.37e-19
C19322 a_12549_44172# a_19862_44208# 0.262561f
C19323 a_n1435_47204# a_383_46660# 4.95e-20
C19324 a_9313_45822# a_2107_46812# 0.298046f
C19325 a_n3690_39616# VDD 0.358567f
C19326 a_7754_38470# a_8530_39574# 0.143675f
C19327 a_20894_47436# a_19321_45002# 1.6e-20
C19328 a_13507_46334# a_13661_43548# 0.038602f
C19329 a_19787_47423# a_19594_46812# 0.108653f
C19330 a_7754_39964# VDAC_P 0.003276f
C19331 a_7754_40130# CAL_N 0.050321f
C19332 a_2063_45854# a_4651_46660# 1.12e-19
C19333 a_n443_46116# a_3699_46634# 0.036317f
C19334 a_n4064_39072# C3_P_btm 1.38e-20
C19335 a_n3420_39072# C1_P_btm 6.64e-20
C19336 VDAC_Pi a_8912_37509# 1.57e-19
C19337 a_n4064_38528# a_n923_35174# 0.004282f
C19338 a_18479_47436# a_21588_30879# 2.9e-20
C19339 a_11599_46634# a_n743_46660# 0.248412f
C19340 a_n971_45724# a_3878_46660# 0.00101f
C19341 a_n1741_47186# a_7411_46660# 8.61e-20
C19342 a_20447_31679# a_22521_40055# 9.79e-21
C19343 a_10807_43548# a_10991_42826# 0.01427f
C19344 a_11750_44172# a_10796_42968# 1.07e-21
C19345 a_10057_43914# a_10533_42308# 7.44e-20
C19346 a_n2293_43922# a_196_42282# 1.63e-19
C19347 a_18494_42460# a_7174_31319# 0.023968f
C19348 a_18184_42460# a_21335_42336# 8.18e-20
C19349 a_17478_45572# VDD 0.411207f
C19350 a_11967_42832# a_15597_42852# 0.004349f
C19351 a_6293_42852# a_5837_43396# 3.72e-20
C19352 a_n356_44636# a_6171_42473# 1.17e-19
C19353 a_11415_45002# a_14021_43940# 3.49e-20
C19354 a_7499_43078# a_4223_44672# 0.02232f
C19355 a_5937_45572# a_n2661_42282# 0.060993f
C19356 a_2274_45254# a_3537_45260# 3.29e-20
C19357 a_3483_46348# a_14955_43940# 0.242667f
C19358 a_n1613_43370# a_n1545_43230# 1.79e-19
C19359 a_13747_46662# a_4361_42308# 4.79e-20
C19360 a_10227_46804# a_13635_43156# 0.320228f
C19361 a_2382_45260# a_3429_45260# 0.011518f
C19362 a_2680_45002# a_3065_45002# 0.13328f
C19363 a_15903_45785# a_16321_45348# 1.49e-19
C19364 a_19692_46634# a_n97_42460# 1.45e-19
C19365 a_2711_45572# a_18287_44626# 1.79e-20
C19366 a_12741_44636# a_12710_44260# 1.22e-20
C19367 a_10428_46928# a_10623_46897# 0.21686f
C19368 a_9863_46634# a_10249_46116# 0.027588f
C19369 a_8492_46660# a_6755_46942# 0.024647f
C19370 a_7411_46660# a_7832_46660# 0.086708f
C19371 a_10150_46912# a_10554_47026# 0.051162f
C19372 a_13487_47204# a_10903_43370# 1.95e-20
C19373 a_13507_46334# a_4185_45028# 0.479559f
C19374 a_n971_45724# a_n1925_42282# 5.37e-19
C19375 a_n746_45260# a_526_44458# 0.096099f
C19376 a_n237_47217# a_2981_46116# 0.024703f
C19377 a_19594_46812# a_20107_46660# 0.001514f
C19378 a_19321_45002# a_20411_46873# 7.75e-19
C19379 a_13661_43548# a_20623_46660# 4.62e-21
C19380 a_4883_46098# a_3483_46348# 0.813604f
C19381 a_11599_46634# a_11189_46129# 0.0158f
C19382 a_10227_46804# a_8016_46348# 0.093061f
C19383 a_13717_47436# a_12594_46348# 4.38e-22
C19384 a_n1435_47204# a_13351_46090# 4.5e-21
C19385 a_n97_42460# a_196_42282# 0.002328f
C19386 a_19721_31679# EN_OFFSET_CAL 3.03e-20
C19387 a_5649_42852# a_10083_42826# 3.09e-20
C19388 a_n3674_39768# a_n4064_40160# 0.139482f
C19389 a_4361_42308# a_10796_42968# 1.44e-19
C19390 a_11341_43940# a_15486_42560# 2.91e-21
C19391 a_15493_43940# a_14113_42308# 1.63e-20
C19392 a_743_42282# a_12089_42308# 0.016016f
C19393 a_15743_43084# a_19339_43156# 0.128224f
C19394 a_n452_44636# VDD 0.112149f
C19395 a_n1177_43370# a_n3674_37592# 4.34e-22
C19396 a_10809_44734# a_12281_43396# 4.31e-19
C19397 a_21101_45002# a_20193_45348# 1.15e-19
C19398 a_n357_42282# a_21381_43940# 0.060125f
C19399 a_n2661_43370# a_n699_43396# 8.19e-19
C19400 a_5691_45260# a_n2661_43922# 5.88e-20
C19401 a_3232_43370# a_n2661_42834# 0.127534f
C19402 a_6171_45002# a_11649_44734# 8.52e-20
C19403 a_3357_43084# a_20835_44721# 5.14e-21
C19404 a_16327_47482# a_20107_42308# 4.96e-19
C19405 a_4185_45028# a_21855_43396# 7.09e-21
C19406 a_18315_45260# a_18545_45144# 0.004937f
C19407 a_9482_43914# a_5891_43370# 0.005232f
C19408 a_n2293_45546# a_n2433_43396# 9.87e-21
C19409 w_1575_34946# a_6886_37412# 0.001151f
C19410 a_n2438_43548# a_997_45618# 0.008987f
C19411 a_n133_46660# a_n755_45592# 2.19e-22
C19412 a_948_46660# a_n863_45724# 1.85e-20
C19413 a_n2293_46634# a_n356_45724# 6.18e-19
C19414 a_19466_46812# a_18819_46122# 0.02948f
C19415 a_11453_44696# a_11823_42460# 0.072491f
C19416 a_12465_44636# a_13904_45546# 1.36e-20
C19417 a_n743_46660# a_1848_45724# 0.003213f
C19418 a_8492_46660# a_8049_45260# 4.06e-21
C19419 a_15227_44166# a_19553_46090# 0.047784f
C19420 a_19333_46634# a_18985_46122# 0.002899f
C19421 a_4883_46098# a_14495_45572# 3.88e-20
C19422 a_383_46660# a_380_45546# 1.76e-21
C19423 a_33_46660# a_310_45028# 3.11e-20
C19424 a_12861_44030# a_14033_45822# 0.003617f
C19425 a_15009_46634# a_10809_44734# 0.00292f
C19426 a_14976_45028# a_6945_45028# 2.34e-19
C19427 a_14035_46660# a_12594_46348# 9.29e-22
C19428 a_3080_42308# a_3754_38802# 4.08e-21
C19429 a_8952_43230# a_5934_30871# 0.001535f
C19430 a_4361_42308# a_4958_30871# 0.087697f
C19431 a_4190_30871# a_18214_42558# 0.078091f
C19432 a_13467_32519# a_17303_42282# 0.040387f
C19433 a_7871_42858# a_8685_42308# 1.33e-20
C19434 a_743_42282# a_18907_42674# 0.00626f
C19435 a_20935_43940# VDD 0.184334f
C19436 a_4185_45028# a_7227_42308# 1.64e-19
C19437 a_12465_44636# CLK 0.795478f
C19438 a_n2433_44484# a_n3674_39768# 0.003677f
C19439 a_n913_45002# a_2982_43646# 0.498826f
C19440 a_n2017_45002# a_3626_43646# 0.023645f
C19441 a_2747_46873# VDD 0.626468f
C19442 a_n2312_39304# DATA[0] 0.001796f
C19443 a_14797_45144# a_15037_43940# 1.29e-20
C19444 a_1307_43914# a_10867_43940# 0.001506f
C19445 a_n2129_44697# a_n4318_39768# 1.04e-19
C19446 a_3357_43084# a_6547_43396# 8.19e-19
C19447 a_n357_42282# a_18249_42858# 0.047936f
C19448 a_n443_42852# a_13113_42826# 0.001005f
C19449 a_15861_45028# a_16243_43396# 5.52e-22
C19450 a_8696_44636# a_16547_43609# 2.74e-20
C19451 a_22612_30879# a_22609_38406# 8.17e-21
C19452 a_22223_47212# EN_OFFSET_CAL 0.011048f
C19453 a_4223_44672# a_3600_43914# 0.00242f
C19454 a_n699_43396# a_2998_44172# 0.127437f
C19455 a_n967_45348# a_n1557_42282# 0.092498f
C19456 a_n2293_43922# a_13296_44484# 3.07e-19
C19457 a_2063_45854# a_8975_43940# 0.149528f
C19458 a_10150_46912# a_2437_43646# 3.29e-20
C19459 a_18597_46090# a_21005_45260# 0.034207f
C19460 a_16327_47482# a_16237_45028# 1.67e-19
C19461 a_10903_43370# a_n357_42282# 0.028411f
C19462 a_18985_46122# a_20062_46116# 1.46e-19
C19463 a_2107_46812# a_7705_45326# 2.71e-20
C19464 a_n2497_47436# a_n1655_44484# 8.54e-19
C19465 a_2804_46116# a_2711_45572# 1.25e-20
C19466 a_n2293_46098# a_4880_45572# 0.013174f
C19467 a_3055_46660# a_413_45260# 0.002017f
C19468 a_20202_43084# a_10193_42453# 0.296862f
C19469 a_9313_45822# a_n2661_44458# 3.78e-20
C19470 a_n2293_46634# a_14537_43396# 0.036569f
C19471 a_2324_44458# a_n2661_45546# 0.019247f
C19472 a_n443_46116# a_4743_44484# 1.56e-21
C19473 a_4791_45118# a_5343_44458# 0.003901f
C19474 a_4883_46098# a_17719_45144# 1.23e-20
C19475 a_3090_45724# a_16842_45938# 1.14e-19
C19476 a_8667_46634# a_3357_43084# 2.31e-20
C19477 a_14180_46812# a_14033_45822# 3.48e-22
C19478 a_3318_42354# a_7174_31319# 4.88e-21
C19479 a_n3674_37592# a_n4334_39616# 6.44e-20
C19480 a_n3674_38680# a_n4209_39304# 8.12e-21
C19481 a_13678_32519# VREF 1.33e-19
C19482 a_n1641_43230# VDD 0.203991f
C19483 a_9803_42558# a_9885_42308# 0.003935f
C19484 a_n1059_45260# a_7309_42852# 0.006756f
C19485 a_5891_43370# a_6031_43396# 0.01824f
C19486 a_20820_30879# C9_N_btm 3.29e-19
C19487 a_21359_45002# a_4190_30871# 3.76e-20
C19488 a_11827_44484# a_21259_43561# 4.17e-22
C19489 a_1307_43914# a_13635_43156# 2.74e-20
C19490 a_3232_43370# a_n2293_42282# 0.00771f
C19491 a_2382_45260# a_3059_42968# 6.58e-20
C19492 a_n2956_38216# a_n2302_40160# 0.001018f
C19493 a_n2661_43922# a_3080_42308# 3.25e-20
C19494 a_n2661_42834# a_4905_42826# 3.66e-20
C19495 a_n2293_42834# a_685_42968# 0.006422f
C19496 a_10440_44484# a_10341_43396# 2.81e-20
C19497 a_10057_43914# a_9885_43646# 8.16e-19
C19498 a_7499_43078# a_5742_30871# 0.019993f
C19499 a_2711_45572# a_17124_42282# 1.5e-21
C19500 a_n2810_45572# a_n4209_39590# 0.020489f
C19501 a_22365_46825# RST_Z 1.22e-19
C19502 a_20567_45036# a_20556_43646# 6.02e-22
C19503 a_11691_44458# a_16823_43084# 5.66e-20
C19504 a_n2661_43370# a_n4318_38680# 0.001014f
C19505 a_14537_43396# a_5342_30871# 1.75e-19
C19506 a_20202_43084# VDD 0.987622f
C19507 a_2711_45572# a_13904_45546# 0.021385f
C19508 a_9290_44172# a_9482_43914# 0.135239f
C19509 a_8016_46348# a_1307_43914# 0.035949f
C19510 a_3090_45724# a_8701_44490# 1.21e-20
C19511 a_19321_45002# a_3422_30871# 6.52e-21
C19512 a_20107_46660# a_18494_42460# 1.14e-20
C19513 a_n2312_40392# a_n4318_39768# 0.025298f
C19514 a_10903_43370# a_11963_45334# 0.209081f
C19515 a_5164_46348# a_1423_45028# 8.94e-20
C19516 a_2324_44458# a_5205_44484# 0.523531f
C19517 a_4646_46812# a_n2661_43922# 0.06073f
C19518 a_n1613_43370# a_453_43940# 1.01e-19
C19519 a_12861_44030# a_15682_43940# 0.016729f
C19520 a_13259_45724# a_18479_45785# 0.004171f
C19521 a_3785_47178# a_n1613_43370# 0.006133f
C19522 a_13487_47204# a_4883_46098# 4.22e-20
C19523 a_1343_38525# a_3754_38470# 4.25e-20
C19524 a_16327_47482# a_18597_46090# 1.28053f
C19525 a_17591_47464# a_10227_46804# 0.292864f
C19526 a_16588_47582# a_18143_47464# 4.68e-20
C19527 a_5742_30871# C8_N_btm 0.003514f
C19528 a_14955_47212# a_13507_46334# 2.55e-20
C19529 a_22775_42308# a_22469_40625# 2.08e-20
C19530 a_5934_30871# VIN_P 0.009408f
C19531 a_13717_47436# a_12465_44636# 0.049141f
C19532 a_10545_42558# VDD 0.004307f
C19533 a_n4334_38304# a_n3690_38304# 8.67e-19
C19534 a_n3420_39616# a_n4064_37440# 0.047863f
C19535 a_n4064_39616# a_n3420_37440# 0.056826f
C19536 a_n4209_38216# a_n3420_37984# 0.067687f
C19537 a_n1917_43396# a_n1557_42282# 7.04e-19
C19538 a_n97_42460# a_4699_43561# 0.025323f
C19539 a_3638_45822# VDD 2.13e-19
C19540 a_18326_43940# a_18525_43370# 0.003065f
C19541 a_18451_43940# a_18429_43548# 0.001082f
C19542 a_15493_43396# a_17499_43370# 0.038093f
C19543 a_n4318_39768# a_n2840_42826# 5.83e-21
C19544 a_11967_42832# a_18083_42858# 0.472348f
C19545 a_18588_44850# a_18249_42858# 1.79e-21
C19546 a_2711_45572# CLK 0.032985f
C19547 a_15493_43940# a_15781_43660# 0.049304f
C19548 a_644_44056# a_791_42968# 3.17e-20
C19549 a_526_44458# a_n310_44484# 1.02e-20
C19550 a_n1079_45724# a_n2661_44458# 6.12e-21
C19551 a_n2293_45546# a_n2433_44484# 1.15e-19
C19552 a_7499_43078# a_n2293_42834# 0.352878f
C19553 a_16327_47482# a_743_42282# 0.026382f
C19554 a_21188_45572# a_19963_31679# 4.63e-19
C19555 a_19466_46812# a_11341_43940# 6.61e-22
C19556 a_19692_46634# a_21115_43940# 4.88e-20
C19557 a_3877_44458# a_n97_42460# 3.76e-22
C19558 a_8696_44636# a_6171_45002# 0.070776f
C19559 a_n2293_46634# a_6547_43396# 0.010751f
C19560 a_584_46384# a_3681_42891# 0.001938f
C19561 a_n971_45724# a_8387_43230# 0.001371f
C19562 a_15227_44166# a_15493_43940# 0.091653f
C19563 a_15682_46116# a_16241_44734# 2.24e-20
C19564 a_768_44030# a_13667_43396# 2.71e-19
C19565 a_12549_44172# a_14579_43548# 1.26e-21
C19566 a_20731_45938# a_3357_43084# 0.005715f
C19567 a_20841_45814# a_21297_45572# 4.2e-19
C19568 a_13059_46348# a_10949_43914# 1.57e-20
C19569 a_4883_46098# a_14513_46634# 3.52e-20
C19570 C3_P_btm VDD 0.26836f
C19571 a_16327_47482# a_19123_46287# 0.005309f
C19572 a_n743_46660# a_7411_46660# 5e-20
C19573 a_n1925_46634# a_7577_46660# 0.007837f
C19574 a_12891_46348# a_11735_46660# 0.034334f
C19575 a_3785_47178# a_n2293_46098# 1.6e-20
C19576 a_11309_47204# a_11813_46116# 0.007374f
C19577 a_n881_46662# a_15009_46634# 0.004074f
C19578 a_n1613_43370# a_3090_45724# 0.039515f
C19579 a_2107_46812# a_6540_46812# 5.62e-20
C19580 a_3177_46902# a_3686_47026# 2.6e-19
C19581 a_2609_46660# a_3055_46660# 2.28e-19
C19582 a_n2661_46634# a_10150_46912# 0.010702f
C19583 a_584_46384# a_376_46348# 0.232754f
C19584 a_1209_47178# a_1176_45822# 4.3e-19
C19585 a_1239_47204# a_1208_46090# 7.29e-20
C19586 a_n237_47217# a_167_45260# 0.280171f
C19587 a_n2109_47186# a_4704_46090# 4.15e-21
C19588 a_n971_45724# a_2698_46116# 0.001385f
C19589 a_n1741_47186# a_4185_45028# 4.26e-20
C19590 a_n1151_42308# a_n1853_46287# 0.024093f
C19591 a_11599_46634# a_20841_46902# 9.01e-21
C19592 a_10227_46804# a_15312_46660# 3.7e-20
C19593 a_17591_47464# a_17339_46660# 3.44e-20
C19594 a_16588_47582# a_765_45546# 0.004612f
C19595 C0_P_btm C9_N_btm 8.4e-19
C19596 C1_P_btm C10_N_btm 0.001745f
C19597 C0_dummy_P_btm C8_N_btm 6.22e-19
C19598 C2_N_btm C4_N_btm 7.19288f
C19599 C1_N_btm C5_N_btm 0.128021f
C19600 C0_N_btm C6_N_btm 0.140033f
C19601 C0_dummy_N_btm C7_N_btm 0.120543f
C19602 a_12465_44636# a_14035_46660# 6.36e-21
C19603 a_15743_43084# a_22591_43396# 0.016556f
C19604 a_5837_45028# VDD 0.191549f
C19605 a_16823_43084# a_4190_30871# 0.004047f
C19606 a_8685_43396# a_10083_42826# 0.007757f
C19607 a_2982_43646# a_20922_43172# 0.004571f
C19608 a_3626_43646# a_19164_43230# 2.65e-20
C19609 a_3080_42308# a_3445_43172# 2.6e-22
C19610 a_4235_43370# a_4156_43218# 9.61e-19
C19611 a_1568_43370# a_873_42968# 1.46e-20
C19612 a_3422_30871# a_17531_42308# 2.58e-20
C19613 a_15415_45028# a_11691_44458# 0.002488f
C19614 a_8560_45348# a_8704_45028# 6.84e-19
C19615 a_4574_45260# a_n699_43396# 1.24e-19
C19616 a_n357_42282# a_14955_43940# 2.08e-21
C19617 a_8199_44636# a_8147_43396# 6.26e-20
C19618 a_20202_43084# a_16137_43396# 5.95e-21
C19619 a_16751_45260# a_11827_44484# 7.2e-21
C19620 a_n443_42852# a_n2661_42282# 0.133617f
C19621 a_3483_46348# a_8685_43396# 6.46e-19
C19622 a_3537_45260# a_4743_44484# 0.01411f
C19623 a_4558_45348# a_4223_44672# 7.57e-20
C19624 a_7705_45326# a_n2661_44458# 1.38e-20
C19625 a_16855_45546# a_17061_44734# 2.71e-21
C19626 a_8696_44636# a_14673_44172# 0.017655f
C19627 a_13259_45724# a_14021_43940# 0.028871f
C19628 a_8270_45546# a_8037_42858# 9.4e-21
C19629 a_3357_43084# a_n356_44636# 3.56e-20
C19630 a_n913_45002# a_14539_43914# 0.003048f
C19631 a_n1059_45260# a_16979_44734# 4.85e-22
C19632 a_n2312_39304# a_n2472_45546# 0.001998f
C19633 a_2107_46812# a_1337_46436# 1.09e-19
C19634 a_n1151_42308# a_8568_45546# 4.03e-20
C19635 a_4791_45118# a_4880_45572# 0.006889f
C19636 a_15227_44166# a_12741_44636# 0.250453f
C19637 a_19692_46634# a_11415_45002# 0.033537f
C19638 a_n2312_40392# a_n2956_38216# 0.053778f
C19639 a_4883_46098# a_n357_42282# 4.03e-19
C19640 a_n2661_46098# a_n1736_46482# 0.024986f
C19641 a_n2438_43548# a_1337_46116# 0.008585f
C19642 a_n743_46660# a_4365_46436# 2.75e-20
C19643 a_5807_45002# a_11387_46482# 2.88e-19
C19644 a_3090_45724# a_n2293_46098# 0.642755f
C19645 a_2063_45854# a_10193_42453# 0.114552f
C19646 a_n1991_42858# a_n3674_37592# 6.3e-20
C19647 a_n809_44244# VDD 0.47719f
C19648 a_9145_43396# a_13657_42308# 1.47e-19
C19649 a_10341_43396# a_15486_42560# 4.67e-21
C19650 a_12895_43230# a_13291_42460# 0.002402f
C19651 a_n2157_42858# a_n1630_35242# 2.26e-19
C19652 a_743_42282# a_5267_42460# 0.010719f
C19653 a_13507_46334# a_22469_40625# 7e-21
C19654 a_18248_44752# a_9313_44734# 1.88e-21
C19655 a_5837_45028# a_5495_43940# 4.33e-21
C19656 a_11827_44484# a_18681_44484# 7.17e-19
C19657 a_2711_45572# a_19268_43646# 3.71e-19
C19658 a_n357_42282# a_5649_42852# 0.011202f
C19659 a_n237_47217# DATA[4] 0.001087f
C19660 a_11823_42460# a_9145_43396# 0.146085f
C19661 a_2063_45854# VDD 3.60498f
C19662 a_10057_43914# a_n2661_43922# 0.034016f
C19663 a_8975_43940# a_n2661_42834# 0.083892f
C19664 a_9482_43914# a_10807_43548# 0.002194f
C19665 a_13017_45260# a_13483_43940# 3.52e-21
C19666 a_18450_45144# a_11967_42832# 1.01e-19
C19667 a_18184_42460# a_3422_30871# 0.649102f
C19668 a_n443_42852# a_16823_43084# 2.55e-21
C19669 a_9290_44172# a_11301_43218# 0.005694f
C19670 a_n2312_38680# a_n2216_38778# 0.003477f
C19671 a_1209_47178# DATA[0] 3.05e-20
C19672 a_327_47204# DATA[1] 2.2e-19
C19673 a_375_42282# a_n2661_42282# 2.72e-19
C19674 a_20193_45348# a_20766_44850# 4.03e-19
C19675 a_10193_42453# a_14955_43396# 4.69e-21
C19676 a_7499_43078# a_10849_43646# 0.003558f
C19677 a_n881_46662# a_1667_45002# 1.43e-20
C19678 a_11813_46116# a_10490_45724# 1.58e-20
C19679 a_20843_47204# a_3357_43084# 0.006792f
C19680 a_19335_46494# a_10809_44734# 7.36e-20
C19681 a_9823_46155# a_5066_45546# 3.05e-20
C19682 a_8016_46348# a_8034_45724# 0.254614f
C19683 a_6419_46155# a_6633_46155# 0.005572f
C19684 a_14035_46660# a_2711_45572# 1.05e-19
C19685 a_11735_46660# a_11322_45546# 5.37e-20
C19686 a_n1151_42308# a_n2661_43370# 0.027798f
C19687 a_4791_45118# a_8560_45348# 6.07e-20
C19688 a_11415_45002# a_20692_30879# 7.79e-19
C19689 a_22591_46660# a_20205_31679# 0.004038f
C19690 a_21588_30879# a_2437_43646# 0.001621f
C19691 a_8667_46634# a_9159_45572# 1.89e-21
C19692 a_6545_47178# a_6945_45348# 2.91e-20
C19693 a_10227_46804# a_16019_45002# 0.001575f
C19694 a_4883_46098# a_11963_45334# 8.43e-21
C19695 a_14955_43396# VDD 0.401358f
C19696 a_5649_42852# CAL_N 0.005399f
C19697 a_13678_32519# a_22521_40599# 2.48e-21
C19698 a_16877_42852# a_17124_42282# 4.18e-19
C19699 a_5267_42460# a_5755_42308# 0.055455f
C19700 a_5379_42460# a_5421_42558# 0.002327f
C19701 a_3318_42354# a_5932_42308# 4.34e-21
C19702 a_2123_42473# a_5934_30871# 1.01e-20
C19703 a_14209_32519# VDAC_N 2.4e-19
C19704 a_n699_43396# a_1568_43370# 0.004191f
C19705 a_n2472_43914# a_n4318_39768# 3.22e-19
C19706 a_1414_42308# a_2889_44172# 0.128883f
C19707 a_1467_44172# a_2998_44172# 1.71e-20
C19708 a_11967_42832# a_12429_44172# 6.2e-19
C19709 a_10193_42453# a_19326_42852# 1.39e-19
C19710 a_n2840_43914# a_n3674_39768# 0.022122f
C19711 a_8270_45546# DATA[4] 0.003852f
C19712 a_n913_45002# a_7871_42858# 0.005608f
C19713 a_n2017_45002# a_8037_42858# 6.62e-20
C19714 a_n1059_45260# a_7765_42852# 0.004965f
C19715 a_n755_45592# a_6123_31319# 0.199766f
C19716 a_n357_42282# a_7963_42308# 4.75e-20
C19717 a_n2956_38680# a_n2946_39866# 3.86e-20
C19718 a_n2956_39304# a_n4064_39616# 3.3e-20
C19719 a_13259_45724# a_15764_42576# 2.69e-19
C19720 a_5891_43370# a_6671_43940# 1.15e-20
C19721 a_12469_46902# VDD 0.203316f
C19722 a_2127_44172# a_895_43940# 0.132679f
C19723 a_18479_47436# a_19279_43940# 0.017993f
C19724 a_16327_47482# a_19789_44512# 1.05e-19
C19725 a_14180_46482# a_11823_42460# 2.88e-20
C19726 a_12638_46436# a_12791_45546# 5.55e-20
C19727 a_8049_45260# a_9241_45822# 7.66e-19
C19728 a_11601_46155# a_11652_45724# 3.78e-19
C19729 a_768_44030# a_5608_44484# 0.001348f
C19730 a_n443_46116# a_1414_42308# 0.18376f
C19731 a_1823_45246# a_n913_45002# 0.041568f
C19732 a_12861_44030# a_20512_43084# 0.005139f
C19733 a_n2293_46634# a_n356_44636# 6.35e-20
C19734 a_17957_46116# a_18175_45572# 8.59e-20
C19735 a_18189_46348# a_18479_45785# 2.57e-19
C19736 a_17715_44484# a_18341_45572# 3.97e-20
C19737 a_n901_46420# a_n467_45028# 2.24e-19
C19738 a_n310_45899# a_n443_42852# 4.25e-19
C19739 a_n755_45592# a_1176_45572# 1.94e-19
C19740 a_18597_46090# a_20835_44721# 0.012854f
C19741 a_13507_46334# a_11967_42832# 0.004262f
C19742 a_n784_42308# C3_P_btm 0.001962f
C19743 a_n971_45724# a_n1435_47204# 2.23698f
C19744 a_3381_47502# a_n443_46116# 4.13e-20
C19745 a_3785_47178# a_4791_45118# 0.010875f
C19746 a_n1151_42308# a_4915_47217# 0.1374f
C19747 a_2063_45854# a_6491_46660# 9.61e-20
C19748 a_n3420_39616# a_n3420_39072# 0.115485f
C19749 a_n4064_39616# a_n3565_39304# 0.028003f
C19750 a_n3565_39590# a_n4064_39072# 0.033734f
C19751 a_19326_42852# VDD 4.6e-19
C19752 a_14097_32519# RST_Z 0.051182f
C19753 a_11967_42832# a_21855_43396# 0.002687f
C19754 a_20640_44752# a_21487_43396# 1.18e-19
C19755 a_n2293_43922# a_1847_42826# 1.69e-20
C19756 a_1307_43914# a_3905_42558# 4.45e-19
C19757 a_18184_42460# a_18504_43218# 3.21e-21
C19758 a_20679_44626# a_20556_43646# 1.59e-20
C19759 a_22591_44484# a_15743_43084# 1.16e-20
C19760 a_20512_43084# a_19700_43370# 7.17e-19
C19761 a_18248_44752# a_18599_43230# 2.16e-21
C19762 a_18989_43940# a_18083_42858# 9.56e-20
C19763 a_18443_44721# a_18249_42858# 3.84e-21
C19764 a_5891_43370# a_10796_42968# 8.14e-20
C19765 a_n2293_42834# a_n1329_42308# 0.002332f
C19766 a_14383_46116# VDD 0.132317f
C19767 a_n356_44636# a_5342_30871# 0.133551f
C19768 a_19279_43940# a_4190_30871# 4.5e-20
C19769 a_n2661_42834# a_2905_42968# 6.38e-21
C19770 a_n2661_42282# a_6655_43762# 4.97e-19
C19771 a_n1613_43370# a_n1821_43396# 1.79e-19
C19772 a_2711_45572# a_10951_45334# 5.77e-20
C19773 a_7227_45028# a_6171_45002# 0.029883f
C19774 a_3775_45552# a_3232_43370# 1.51e-20
C19775 a_6598_45938# a_6431_45366# 0.001277f
C19776 a_3090_45724# a_2675_43914# 3.49e-22
C19777 a_n443_42852# a_15415_45028# 1.77e-21
C19778 a_6511_45714# a_7276_45260# 1.03e-19
C19779 a_6667_45809# a_5205_44484# 1.28e-19
C19780 a_8049_45260# a_21005_45260# 1.99e-20
C19781 a_17478_45572# a_18479_45785# 3.4e-19
C19782 a_15861_45028# a_18341_45572# 9.93e-20
C19783 a_n901_46420# a_n2661_43922# 1.04e-20
C19784 a_11823_42460# a_n1059_45260# 0.100641f
C19785 a_6945_45028# a_5343_44458# 4.48e-20
C19786 a_2324_44458# a_13076_44458# 7.95e-21
C19787 a_3316_45546# a_1423_45028# 1.81e-19
C19788 a_n3420_37440# C0_P_btm 0.033333f
C19789 a_n4064_37440# C2_P_btm 0.001797f
C19790 a_n881_46662# a_2959_46660# 2.16e-20
C19791 a_n1613_43370# a_3699_46634# 0.344308f
C19792 a_7754_38968# VDD 0.041093f
C19793 a_16327_47482# a_6755_46942# 0.067305f
C19794 a_13661_43548# a_n743_46660# 1.74e-19
C19795 a_4915_47217# a_14084_46812# 0.038663f
C19796 a_6151_47436# a_12991_46634# 2.17e-19
C19797 a_4791_45118# a_3090_45724# 0.206257f
C19798 a_22521_39511# a_22717_37285# 2.12e-20
C19799 a_10227_46804# a_10428_46928# 0.060058f
C19800 a_20447_31679# VCM 0.035344f
C19801 a_8685_43396# a_16664_43396# 1.93e-19
C19802 a_n809_44244# a_n784_42308# 1.32e-20
C19803 a_n955_45028# VDD 0.004233f
C19804 a_10341_43396# a_13837_43396# 7.41e-20
C19805 a_13565_43940# a_12545_42858# 1.31e-20
C19806 a_n1557_42282# a_n1853_43023# 1.74e-20
C19807 a_6547_43396# a_743_42282# 3.34e-20
C19808 a_n1761_44111# a_n1630_35242# 0.060838f
C19809 a_10807_43548# a_11301_43218# 0.001467f
C19810 a_n97_42460# a_1847_42826# 2.77e-20
C19811 a_14955_43396# a_16137_43396# 7.94e-20
C19812 a_14205_43396# a_16547_43609# 8.78e-22
C19813 a_15095_43370# a_16243_43396# 2.69e-21
C19814 a_6755_46942# a_16855_43396# 6.28e-20
C19815 a_13661_43548# a_17701_42308# 3.31e-20
C19816 a_12549_44172# a_21671_42860# 0.001174f
C19817 a_16019_45002# a_1307_43914# 0.01609f
C19818 a_6709_45028# a_6517_45366# 5.76e-19
C19819 a_10193_42453# a_n2661_42834# 0.034215f
C19820 a_10180_45724# a_n2661_43922# 1.65e-19
C19821 a_21513_45002# a_11827_44484# 0.010541f
C19822 a_10227_46804# a_13814_43218# 0.001965f
C19823 a_8953_45546# a_9420_43940# 2.33e-19
C19824 a_327_44734# a_n2661_43370# 0.035472f
C19825 a_8696_44636# a_12607_44458# 0.005383f
C19826 a_5691_45260# a_5837_45028# 0.171361f
C19827 a_n2956_38216# a_n2472_43914# 7.64e-21
C19828 a_3357_43084# a_20567_45036# 4.77e-19
C19829 a_19479_31679# a_21005_45260# 3.22e-19
C19830 a_2324_44458# a_15301_44260# 1.99e-19
C19831 a_n1151_42308# COMP_P 0.034f
C19832 a_18189_46348# a_14021_43940# 2.08e-20
C19833 a_n2293_46634# a_12379_42858# 1.17e-19
C19834 a_12891_46348# a_2324_44458# 0.026746f
C19835 a_12549_44172# a_14840_46494# 9.46e-38
C19836 a_n237_47217# a_n863_45724# 3.43e-19
C19837 a_n746_45260# a_n452_45724# 3.79e-20
C19838 a_n2661_46098# a_n1641_46494# 0.035694f
C19839 a_2107_46812# a_1823_45246# 0.007836f
C19840 a_10150_46912# a_765_45546# 4.34e-20
C19841 a_5807_45002# a_11133_46155# 0.00164f
C19842 a_n743_46660# a_4185_45028# 0.036891f
C19843 a_3699_46634# a_n2293_46098# 1.64e-20
C19844 a_1239_47204# a_n2661_45546# 4.78e-21
C19845 a_11735_46660# a_12359_47026# 9.73e-19
C19846 a_11813_46116# a_12156_46660# 0.157972f
C19847 a_14976_45028# a_15559_46634# 0.001514f
C19848 a_n1925_46634# a_4704_46090# 2.8e-20
C19849 a_n2661_46634# a_6419_46155# 1.76e-21
C19850 a_1123_46634# a_167_45260# 0.003466f
C19851 a_n452_47436# a_n1099_45572# 3.76e-20
C19852 a_n2497_47436# a_3316_45546# 1.34e-19
C19853 a_16327_47482# a_8049_45260# 0.605463f
C19854 a_16137_43396# a_19326_42852# 1.63e-20
C19855 a_n97_42460# a_15486_42560# 0.055334f
C19856 a_12545_42858# a_5534_30871# 0.17182f
C19857 a_12895_43230# a_13460_43230# 7.99e-20
C19858 a_2982_43646# a_8325_42308# 1.03e-19
C19859 a_3626_43646# a_4169_42308# 6.63e-19
C19860 a_n2661_42834# VDD 1.00348f
C19861 a_17730_32519# VDAC_N 0.00723f
C19862 a_2905_42968# a_n2293_42282# 0.001495f
C19863 a_n913_45002# a_n3674_39768# 2.02e-20
C19864 a_13259_45724# a_13943_43396# 2.96e-20
C19865 a_9290_44172# a_10796_42968# 0.050429f
C19866 a_3483_46348# a_17333_42852# 1.51e-19
C19867 a_4185_45028# a_17701_42308# 5.35e-20
C19868 a_n357_42282# a_8685_43396# 0.319118f
C19869 a_10907_45822# a_11257_43940# 8.34e-20
C19870 a_n443_42852# a_7112_43396# 0.00494f
C19871 a_3537_45260# a_1414_42308# 1.29e-19
C19872 a_2274_45254# a_2675_43914# 1.86e-20
C19873 a_2680_45002# a_2479_44172# 1.33e-19
C19874 a_16922_45042# a_9313_44734# 5.83e-19
C19875 a_413_45260# a_3600_43914# 2.35e-19
C19876 a_5343_44458# a_8103_44636# 0.001348f
C19877 a_16147_45260# a_11341_43940# 2.74e-20
C19878 a_18597_46090# a_20731_45938# 1.8e-20
C19879 a_16241_47178# a_3357_43084# 1.11e-19
C19880 a_16327_47482# a_19479_31679# 1.04e-19
C19881 a_12549_44172# a_16115_45572# 1.27e-21
C19882 a_2063_45854# a_5691_45260# 6.94e-20
C19883 a_584_46384# a_3232_43370# 0.277433f
C19884 a_15227_44166# a_16375_45002# 0.117865f
C19885 a_5129_47502# a_413_45260# 1.79e-19
C19886 a_n443_46116# a_1667_45002# 4.2e-20
C19887 a_16763_47508# a_2437_43646# 0.014946f
C19888 a_n2661_46634# a_10907_45822# 6.03e-21
C19889 a_22959_46660# a_10809_44734# 0.015306f
C19890 a_6165_46155# a_5937_45572# 1.14e-20
C19891 a_12741_44636# a_22959_46124# 3.35e-19
C19892 a_13507_46334# a_20273_45572# 7.72e-20
C19893 a_3080_42308# C3_P_btm 0.027071f
C19894 a_n1352_43396# VDD 0.288329f
C19895 a_16795_42852# a_17303_42282# 0.010298f
C19896 a_17595_43084# a_4958_30871# 9.74e-19
C19897 a_n4318_38216# a_n3674_38216# 2.91597f
C19898 a_n3674_38680# a_n4318_37592# 0.084223f
C19899 a_n2840_42282# COMP_P 7.51e-20
C19900 a_8495_42852# a_5934_30871# 8.72e-19
C19901 a_n3674_39304# a_n4334_39392# 0.060327f
C19902 a_4185_45028# a_21613_42308# 0.028903f
C19903 a_16922_45042# a_20974_43370# 0.077191f
C19904 a_17767_44458# a_18079_43940# 3.68e-19
C19905 a_2107_46812# DATA[2] 5.18e-20
C19906 a_1423_45028# a_6197_43396# 4.8e-22
C19907 a_2324_44458# a_15720_42674# 2.94e-22
C19908 a_5111_44636# a_10341_43396# 0.009186f
C19909 a_n2661_43922# a_5013_44260# 7.36e-20
C19910 a_n2661_42834# a_5495_43940# 0.009774f
C19911 a_20679_44626# a_20980_44850# 9.73e-19
C19912 a_20640_44752# a_21398_44850# 0.056391f
C19913 a_20766_44850# a_20596_44850# 2.6e-19
C19914 a_20362_44736# a_3422_30871# 3.94e-20
C19915 a_1307_43914# a_8791_43396# 4.19e-20
C19916 a_17970_44736# a_17973_43940# 0.002178f
C19917 a_n2293_42834# a_1756_43548# 1.53e-20
C19918 a_19778_44110# a_19319_43548# 0.003354f
C19919 a_n357_42282# a_15953_42852# 0.00164f
C19920 a_n1059_45260# a_18429_43548# 0.002978f
C19921 a_n913_45002# a_17324_43396# 7.64e-21
C19922 a_11453_44696# a_14539_43914# 0.006758f
C19923 a_12594_46348# a_13527_45546# 0.100424f
C19924 a_13925_46122# a_11823_42460# 2.39e-19
C19925 a_13351_46090# a_13163_45724# 3.18e-19
C19926 a_4651_46660# a_5093_45028# 1.49e-21
C19927 a_6755_46942# a_14537_43396# 0.120241f
C19928 a_17715_44484# a_10193_42453# 0.074403f
C19929 a_4646_46812# a_5837_45028# 1.48e-21
C19930 a_8199_44636# a_10907_45822# 0.081841f
C19931 a_5937_45572# a_10210_45822# 2.86e-19
C19932 a_8953_45546# a_9241_45822# 2.68e-20
C19933 a_15227_44166# a_413_45260# 4.28e-20
C19934 a_2324_44458# a_11322_45546# 0.068998f
C19935 a_10903_43370# a_13249_42308# 0.211356f
C19936 a_4955_46873# a_5009_45028# 4.28e-21
C19937 a_11813_46116# a_6171_45002# 1.01e-20
C19938 a_16721_46634# a_3357_43084# 7.55e-22
C19939 a_20841_46902# a_20841_45814# 8.24e-19
C19940 a_20273_46660# a_20623_45572# 3.64e-20
C19941 a_20623_46660# a_20273_45572# 1.3e-20
C19942 a_20107_46660# a_21188_45572# 2.1e-20
C19943 a_11415_45002# a_18175_45572# 0.003704f
C19944 a_3090_45724# a_3429_45260# 0.004791f
C19945 a_n881_46662# a_n699_43396# 6.09e-22
C19946 a_8270_45546# a_8191_45002# 0.001376f
C19947 a_526_44458# a_3175_45822# 0.003323f
C19948 a_n1925_42282# a_2711_45572# 0.019937f
C19949 a_5934_30871# a_n3565_38502# 4.1e-21
C19950 a_n2293_42282# VDD 0.464485f
C19951 a_19332_42282# a_19647_42308# 0.084365f
C19952 a_18214_42558# a_19511_42282# 9.74e-21
C19953 a_22959_42860# RST_Z 0.001357f
C19954 COMP_P VDAC_Ni 9.79e-19
C19955 a_17303_42282# a_21335_42336# 2.99e-19
C19956 a_17531_42308# a_7174_31319# 2.13e-20
C19957 a_6123_31319# a_n3420_38528# 0.003315f
C19958 a_20935_43940# a_14021_43940# 7.94e-20
C19959 a_n2956_37592# a_n1630_35242# 5.5e-19
C19960 a_n1059_45260# a_961_42354# 0.07089f
C19961 a_n913_45002# a_1184_42692# 0.031137f
C19962 a_n2017_45002# a_1149_42558# 4.17e-19
C19963 a_9028_43914# a_9420_43940# 0.016359f
C19964 a_n1899_43946# a_n1557_42282# 1.37e-19
C19965 a_1467_44172# a_1568_43370# 0.055004f
C19966 a_1414_42308# a_1049_43396# 0.003017f
C19967 a_9313_44734# a_15743_43084# 1.48048f
C19968 a_12005_46116# CLK 8.86e-21
C19969 a_949_44458# a_791_42968# 3.01e-19
C19970 a_742_44458# a_1847_42826# 0.372436f
C19971 a_14673_44172# a_14205_43396# 7.49e-20
C19972 a_n967_45348# a_n3674_37592# 0.002659f
C19973 a_17715_44484# VDD 0.526119f
C19974 a_5244_44056# a_n97_42460# 2.33e-20
C19975 a_17583_46090# RST_Z 1.08e-21
C19976 a_n3674_39768# a_n4318_39304# 2.75695f
C19977 a_3357_43084# a_3823_42558# 3.77e-19
C19978 a_n2293_42834# a_5193_43172# 2.71e-19
C19979 a_n2661_44458# a_7871_42858# 6.62e-21
C19980 a_n356_44636# a_743_42282# 0.063042f
C19981 a_12549_44172# a_19478_44306# 0.010691f
C19982 a_5066_45546# a_1423_45028# 3.17e-20
C19983 a_13527_45546# a_15037_45618# 2.92e-22
C19984 a_13904_45546# a_14033_45822# 0.062574f
C19985 a_12861_44030# a_21381_43940# 0.019154f
C19986 a_n901_46420# a_n452_44636# 1.9e-20
C19987 a_8746_45002# a_8696_44636# 0.058163f
C19988 a_10193_42453# a_15861_45028# 0.432483f
C19989 a_n863_45724# a_n2017_45002# 0.111825f
C19990 a_n2661_45546# a_n2956_37592# 6.64e-20
C19991 a_n2810_45572# en_comp 2.18e-19
C19992 a_8049_45260# a_14537_43396# 3.16e-21
C19993 a_14493_46090# a_14309_45028# 1.04e-20
C19994 a_2324_44458# a_15060_45348# 0.004184f
C19995 a_11823_42460# a_15599_45572# 3.42e-19
C19996 a_1823_45246# a_n2661_44458# 0.036985f
C19997 a_n2293_45546# a_n913_45002# 0.043147f
C19998 a_n1079_45724# a_n1059_45260# 0.003242f
C19999 a_310_45028# a_n2661_45010# 1.15e-19
C20000 a_n2293_46098# a_4743_44484# 0.002464f
C20001 a_n3565_39590# VDD 1.26658f
C20002 a_13507_46334# a_5807_45002# 1.64614f
C20003 a_20990_47178# a_13747_46662# 1.78e-20
C20004 a_19787_47423# a_19321_45002# 0.029499f
C20005 a_7754_40130# a_11206_38545# 0.736866f
C20006 a_7754_39964# a_8912_37509# 0.003864f
C20007 a_2063_45854# a_4646_46812# 0.093604f
C20008 a_n443_46116# a_2959_46660# 0.036727f
C20009 a_12465_44636# a_16285_47570# 1.31e-20
C20010 a_n3565_39304# C0_P_btm 9.35e-21
C20011 a_n4064_39072# C4_P_btm 1.7e-20
C20012 a_19386_47436# a_19594_46812# 0.069651f
C20013 a_n3420_38528# EN_VIN_BSTR_P 0.031973f
C20014 a_18479_47436# a_20916_46384# 0.014237f
C20015 a_14955_47212# a_n743_46660# 6.75e-21
C20016 a_n971_45724# a_3633_46660# 2.76e-19
C20017 a_n1741_47186# a_5257_43370# 1.22e-19
C20018 a_10405_44172# a_10341_42308# 5.11e-21
C20019 a_10949_43914# a_10991_42826# 3.02e-20
C20020 a_10807_43548# a_10796_42968# 0.030352f
C20021 a_11750_44172# a_10835_43094# 2e-20
C20022 a_19963_31679# a_22459_39145# 2.14e-20
C20023 a_3905_42865# a_4156_43218# 7.76e-19
C20024 a_n2293_43922# a_n473_42460# 8.65e-20
C20025 a_2982_43646# a_9145_43396# 1.33e-20
C20026 a_18184_42460# a_7174_31319# 0.007789f
C20027 a_15861_45028# VDD 0.690795f
C20028 a_8791_43396# a_9396_43370# 0.011032f
C20029 a_20974_43370# a_15743_43084# 6.72e-19
C20030 a_n356_44636# a_5755_42308# 2.77e-19
C20031 a_20202_43084# a_14021_43940# 0.020234f
C20032 a_8049_45260# a_20835_44721# 3.74e-21
C20033 a_5937_45572# a_6101_44260# 9.35e-20
C20034 a_12861_44030# a_18249_42858# 6.95e-20
C20035 a_n1613_43370# a_n1736_43218# 2.47e-19
C20036 a_n863_45724# a_n89_44484# 8.7e-19
C20037 a_3483_46348# a_13483_43940# 0.194464f
C20038 a_13661_43548# a_4361_42308# 6.79e-20
C20039 a_10227_46804# a_12895_43230# 0.152365f
C20040 a_413_45260# a_4558_45348# 4.69e-20
C20041 a_2382_45260# a_3065_45002# 0.632538f
C20042 a_13259_45724# a_13296_44484# 0.002753f
C20043 a_2711_45572# a_18248_44752# 8.88e-20
C20044 a_8667_46634# a_6755_46942# 0.011524f
C20045 a_10428_46928# a_10467_46802# 0.820079f
C20046 a_10150_46912# a_10623_46897# 7.99e-20
C20047 a_5257_43370# a_7832_46660# 2.48e-21
C20048 a_12861_44030# a_10903_43370# 0.378457f
C20049 a_n971_45724# a_526_44458# 0.21769f
C20050 a_n1151_42308# a_10809_44734# 0.334692f
C20051 a_19321_45002# a_20107_46660# 0.003274f
C20052 a_19594_46812# a_19551_46910# 0.07027f
C20053 a_13747_46662# a_20273_46660# 1.3e-20
C20054 a_4883_46098# a_3147_46376# 1.86e-19
C20055 a_n1435_47204# a_12594_46348# 1.19e-20
C20056 a_13381_47204# a_13351_46090# 7.4e-20
C20057 a_7577_46660# a_6999_46987# 5.54e-20
C20058 a_n97_42460# a_n473_42460# 0.096579f
C20059 a_5649_42852# a_8952_43230# 3.14e-21
C20060 a_n1076_43230# a_791_42968# 4.35e-20
C20061 a_n13_43084# a_685_42968# 0.002159f
C20062 a_n2267_43396# a_n1630_35242# 2.12e-20
C20063 a_n4318_39768# a_n4064_40160# 0.293052f
C20064 a_4361_42308# a_10835_43094# 2.74e-20
C20065 a_8685_43396# a_10553_43218# 1.84e-19
C20066 a_743_42282# a_12379_42858# 2.73e-19
C20067 a_15743_43084# a_18599_43230# 0.001457f
C20068 a_n1352_44484# VDD 0.276725f
C20069 a_15682_43940# a_17124_42282# 8.07e-20
C20070 a_n3674_39768# a_n4334_40480# 0.004086f
C20071 a_n1917_43396# a_n3674_37592# 1.93e-20
C20072 a_11341_43940# a_15051_42282# 3.24e-20
C20073 a_4185_45028# a_4361_42308# 0.042181f
C20074 a_21101_45002# a_11691_44458# 1.41e-20
C20075 a_11827_44484# a_22959_45036# 4.91e-20
C20076 a_21005_45260# a_20193_45348# 3.32e-20
C20077 a_5111_44636# a_n2293_43922# 4.86e-20
C20078 a_13249_42308# a_14955_43940# 6.27e-21
C20079 a_10193_42453# a_20623_43914# 0.001477f
C20080 a_n2661_43370# a_4223_44672# 0.001914f
C20081 a_5691_45260# a_n2661_42834# 1.59e-21
C20082 a_3232_43370# a_11649_44734# 0.011508f
C20083 a_3357_43084# a_20679_44626# 5.72e-21
C20084 a_16327_47482# a_13258_32519# 0.019817f
C20085 a_n2293_46634# a_3823_42558# 8.78e-21
C20086 a_17715_44484# a_16137_43396# 1.22e-20
C20087 a_21363_45546# a_3422_30871# 9.12e-20
C20088 a_18315_45260# a_18450_45144# 0.008535f
C20089 a_626_44172# a_n356_44636# 0.249281f
C20090 SMPL_ON_P a_n3420_38528# 8.16e-21
C20091 a_n743_46660# a_997_45618# 2.04e-19
C20092 a_n2438_43548# a_n755_45592# 0.213107f
C20093 a_1123_46634# a_n863_45724# 2.27e-20
C20094 a_n133_46660# a_n357_42282# 1.78e-19
C20095 a_14180_46812# a_10903_43370# 7.73e-19
C20096 a_12465_44636# a_13527_45546# 6.66e-22
C20097 a_11453_44696# a_12427_45724# 5.75e-21
C20098 a_8667_46634# a_8049_45260# 0.00101f
C20099 a_19333_46634# a_18819_46122# 0.003156f
C20100 a_15227_44166# a_18985_46122# 0.287996f
C20101 a_13507_46334# a_15143_45578# 3.04e-21
C20102 a_4883_46098# a_13249_42308# 3.03e-20
C20103 a_n1925_46634# a_2957_45546# 1.1e-20
C20104 a_33_46660# a_n1099_45572# 5.76e-21
C20105 a_171_46873# a_310_45028# 1.19e-19
C20106 a_2107_46812# a_n2293_45546# 2.33e-20
C20107 a_14084_46812# a_10809_44734# 0.004861f
C20108 a_3090_45724# a_6945_45028# 2.98e-19
C20109 a_9127_43156# a_5934_30871# 0.003851f
C20110 a_8387_43230# a_8515_42308# 7.06e-20
C20111 a_4361_42308# a_16269_42308# 2.5e-19
C20112 a_4190_30871# a_19332_42282# 0.154377f
C20113 a_13467_32519# a_4958_30871# 0.031235f
C20114 a_n2293_42282# a_n784_42308# 0.055588f
C20115 a_7871_42858# a_8325_42308# 7.98e-19
C20116 a_743_42282# a_18727_42674# 0.006169f
C20117 a_17538_32519# VDAC_N 0.004499f
C20118 a_20623_43914# VDD 0.258478f
C20119 a_n2312_39304# CLK_DATA 0.003547f
C20120 a_4185_45028# a_6761_42308# 9.41e-20
C20121 a_n2661_44458# a_n3674_39768# 0.037999f
C20122 a_n2433_44484# a_n4318_39768# 0.00138f
C20123 a_n1059_45260# a_2982_43646# 0.020128f
C20124 a_13249_42308# a_5649_42852# 3.17e-20
C20125 a_14537_43396# a_15037_43940# 0.018234f
C20126 a_1307_43914# a_10651_43940# 0.001528f
C20127 a_3357_43084# a_6765_43638# 3.46e-19
C20128 a_n443_42852# a_12545_42858# 7.04e-20
C20129 a_n357_42282# a_17333_42852# 0.05273f
C20130 a_12465_44636# EN_OFFSET_CAL 2.39e-20
C20131 a_21588_30879# a_22609_38406# 6.34e-21
C20132 a_16922_45042# a_17737_43940# 6.1e-19
C20133 a_17023_45118# a_15682_43940# 8.14e-19
C20134 a_4223_44672# a_2998_44172# 0.035464f
C20135 a_n699_43396# a_2889_44172# 0.006735f
C20136 en_comp a_n1557_42282# 4.48e-20
C20137 a_n2293_43922# a_12829_44484# 0.009626f
C20138 a_5111_44636# a_n97_42460# 0.211832f
C20139 a_2063_45854# a_10057_43914# 0.06633f
C20140 a_n1151_42308# a_5883_43914# 1.46e-20
C20141 a_n443_46116# a_n699_43396# 0.042248f
C20142 a_12861_44030# a_19929_45028# 7.5e-19
C20143 a_9863_46634# a_2437_43646# 9.58e-21
C20144 a_13507_46334# a_18315_45260# 8.76e-37
C20145 a_18597_46090# a_20567_45036# 0.001626f
C20146 a_16327_47482# a_20193_45348# 0.359904f
C20147 a_n743_46660# a_13159_45002# 7.14e-21
C20148 a_19900_46494# a_20009_46494# 0.007416f
C20149 a_20075_46420# a_20254_46482# 0.007399f
C20150 a_19335_46494# a_19443_46116# 0.057222f
C20151 a_n2497_47436# a_n1821_44484# 0.001505f
C20152 a_2698_46116# a_2711_45572# 6.21e-20
C20153 a_n2293_46098# a_4808_45572# 0.001218f
C20154 a_11453_44696# a_14309_45028# 0.004516f
C20155 a_18479_47436# a_21101_45002# 0.001064f
C20156 a_10227_46804# a_11827_44484# 0.065169f
C20157 a_7927_46660# a_3357_43084# 1.64e-20
C20158 a_14035_46660# a_14033_45822# 0.001323f
C20159 a_4791_45118# a_4743_44484# 0.165321f
C20160 a_2903_42308# a_7174_31319# 9.76e-21
C20161 a_n3674_37592# a_n4209_39590# 3.94e-20
C20162 a_13070_42354# a_13575_42558# 1e-19
C20163 COMP_P a_n2302_39866# 1.42e-19
C20164 a_n1423_42826# VDD 0.211036f
C20165 a_9223_42460# a_9885_42308# 9.07e-20
C20166 a_13678_32519# VIN_N 0.069898f
C20167 a_13467_32519# VCM 0.020152f
C20168 a_14539_43914# a_9145_43396# 0.008138f
C20169 a_n1059_45260# a_5837_42852# 0.005989f
C20170 a_20159_44458# a_19319_43548# 6.17e-19
C20171 a_20820_30879# C8_N_btm 9.97e-19
C20172 a_2382_45260# a_2987_42968# 6.35e-20
C20173 a_10193_42453# a_9885_42558# 0.006254f
C20174 a_n2956_38216# a_n4064_40160# 9.27e-19
C20175 a_n2661_43922# a_4699_43561# 3.07e-20
C20176 a_n2661_42834# a_3080_42308# 2.61e-19
C20177 a_21076_30879# C5_N_btm 1.31e-19
C20178 a_18114_32519# a_15743_43084# 1.84e-21
C20179 a_n2293_42834# a_421_43172# 2.71e-19
C20180 a_6109_44484# a_6197_43396# 0.001019f
C20181 a_10334_44484# a_10341_43396# 4.4e-19
C20182 a_13720_44458# a_13667_43396# 2.79e-20
C20183 a_7499_43078# a_11323_42473# 5.37e-19
C20184 a_2711_45572# a_16522_42674# 8.16e-20
C20185 a_18184_42460# a_21487_43396# 5.5e-20
C20186 a_11691_44458# a_17021_43396# 1.04e-20
C20187 a_n2661_43370# a_n3674_39304# 0.002283f
C20188 a_22365_46825# VDD 0.193587f
C20189 a_2711_45572# a_13527_45546# 0.006151f
C20190 a_n743_46660# a_11967_42832# 7.36e-20
C20191 a_n967_46494# a_n967_45348# 1.79e-21
C20192 a_15682_46116# a_6171_45002# 2.79e-19
C20193 a_2324_44458# a_6431_45366# 0.046214f
C20194 a_22959_46124# a_413_45260# 0.020082f
C20195 a_526_44458# a_n2293_45010# 2.25e-19
C20196 a_20107_46660# a_18184_42460# 3.9e-21
C20197 a_17339_46660# a_11827_44484# 0.031147f
C20198 a_8049_45260# a_20731_45938# 0.005076f
C20199 a_20411_46873# a_19778_44110# 1.83e-20
C20200 a_10903_43370# a_11787_45002# 0.003455f
C20201 a_12861_44030# a_14955_43940# 0.001655f
C20202 a_20528_46660# a_16922_45042# 3.33e-20
C20203 a_13259_45724# a_18175_45572# 3.33e-19
C20204 a_4646_46812# a_n2661_42834# 0.030297f
C20205 a_3877_44458# a_n2661_43922# 0.021496f
C20206 a_2063_45854# a_9804_47204# 0.249806f
C20207 a_n1151_42308# a_n881_46662# 1.41446f
C20208 a_3381_47502# a_n1613_43370# 5.5e-21
C20209 a_4700_47436# a_4842_47570# 0.007833f
C20210 a_14311_47204# a_13507_46334# 1.05e-20
C20211 a_n3565_39590# a_n2302_37690# 2.81e-19
C20212 a_13717_47436# a_21811_47423# 6.87e-20
C20213 a_12861_44030# a_4883_46098# 0.076083f
C20214 a_6123_31319# VIN_N 0.01057f
C20215 a_16588_47582# a_10227_46804# 0.039575f
C20216 a_5742_30871# C7_N_btm 0.04157f
C20217 a_21613_42308# a_22469_40625# 1.4e-21
C20218 a_22775_42308# a_22521_40599# 1.89e-20
C20219 a_n1741_47186# a_5807_45002# 0.029376f
C20220 a_n1435_47204# a_12465_44636# 0.002293f
C20221 a_9885_42558# VDD 0.18767f
C20222 a_16327_47482# a_18780_47178# 5.16e-20
C20223 a_n3607_38528# a_n3420_37984# 3.77e-20
C20224 a_n4334_38304# a_n3565_38216# 0.001004f
C20225 a_n4209_38216# a_n3690_38304# 0.045342f
C20226 a_2112_39137# VDAC_Pi 0.01062f
C20227 a_644_44056# a_685_42968# 2.21e-19
C20228 a_n97_42460# a_4235_43370# 0.003683f
C20229 a_n1699_43638# a_n1557_42282# 3.96e-21
C20230 a_17737_43940# a_15743_43084# 1.41e-19
C20231 a_3775_45552# VDD 0.089667f
C20232 a_18326_43940# a_18429_43548# 9.67e-19
C20233 a_15493_43396# a_16759_43396# 0.029803f
C20234 a_14021_43940# a_14955_43396# 0.01294f
C20235 a_11967_42832# a_17701_42308# 0.030406f
C20236 a_15493_43940# a_15681_43442# 0.03571f
C20237 a_11453_44696# a_17324_43396# 1.49e-21
C20238 a_12839_46116# a_13076_44458# 4.31e-21
C20239 a_526_44458# a_9313_44734# 4.07e-20
C20240 a_n2661_45546# a_n2267_44484# 2.71e-20
C20241 a_n2956_38216# a_n2433_44484# 7.79e-19
C20242 a_n2293_45546# a_n2661_44458# 0.006992f
C20243 a_21363_45546# a_19963_31679# 2.99e-19
C20244 a_19692_46634# a_20935_43940# 6.93e-20
C20245 a_n2956_38680# a_n2293_43922# 3.35e-20
C20246 a_8696_44636# a_3232_43370# 0.169534f
C20247 a_16680_45572# a_6171_45002# 7.1e-19
C20248 a_n2293_46634# a_6765_43638# 0.011639f
C20249 a_16327_47482# a_20301_43646# 4.99e-19
C20250 a_584_46384# a_2905_42968# 3.05e-20
C20251 a_n971_45724# a_8605_42826# 0.001728f
C20252 a_2711_45572# a_16922_45042# 1.19e-19
C20253 a_768_44030# a_10695_43548# 3.8e-21
C20254 a_12861_44030# a_5649_42852# 1.34e-19
C20255 a_20528_45572# a_3357_43084# 5.18e-19
C20256 a_21188_45572# a_22591_45572# 1.52e-20
C20257 a_20273_45572# a_21297_45572# 2.36e-20
C20258 a_n2109_47186# a_4419_46090# 3.48e-20
C20259 a_n971_45724# a_2521_46116# 6.68e-20
C20260 a_n746_45260# a_167_45260# 0.234425f
C20261 a_n83_35174# VIN_P 0.001664f
C20262 a_4883_46098# a_14180_46812# 8.02e-20
C20263 C4_P_btm VDD 0.265463f
C20264 a_16327_47482# a_18285_46348# 3.07e-20
C20265 a_n743_46660# a_5257_43370# 0.036418f
C20266 a_n1925_46634# a_7715_46873# 0.01948f
C20267 a_5807_45002# a_7832_46660# 0.001677f
C20268 a_n237_47217# a_2202_46116# 0.049087f
C20269 a_n1151_42308# a_n2157_46122# 0.027101f
C20270 a_11309_47204# a_11735_46660# 0.003123f
C20271 a_4915_47217# a_12741_44636# 0.031734f
C20272 a_16763_47508# a_765_45546# 0.005699f
C20273 a_2107_46812# a_5732_46660# 0.00317f
C20274 a_2609_46660# a_3686_47026# 1.46e-19
C20275 a_2443_46660# a_3055_46660# 0.001881f
C20276 a_n2661_46634# a_9863_46634# 0.010932f
C20277 a_584_46384# a_n1076_46494# 5.23e-20
C20278 a_1209_47178# a_1208_46090# 7.67e-19
C20279 a_13717_47436# a_22000_46634# 3.86e-20
C20280 a_11599_46634# a_20273_46660# 0.003014f
C20281 a_10227_46804# a_14447_46660# 2.5e-20
C20282 C0_P_btm C8_N_btm 7e-19
C20283 C1_P_btm C9_N_btm 9.52e-19
C20284 C0_dummy_P_btm C7_N_btm 3.73e-19
C20285 C1_N_btm C4_N_btm 0.128692f
C20286 C0_N_btm C5_N_btm 0.138736f
C20287 C2_N_btm C3_N_btm 5.64696f
C20288 C0_dummy_N_btm C6_N_btm 0.120464f
C20289 a_12465_44636# a_13885_46660# 0.006386f
C20290 a_n97_42460# a_5837_43172# 0.006105f
C20291 a_4235_43370# a_3935_43218# 3.44e-20
C20292 a_1568_43370# a_133_42852# 1.19e-20
C20293 a_n2661_42282# a_4921_42308# 0.001195f
C20294 a_19700_43370# a_5649_42852# 1.35e-22
C20295 a_15743_43084# a_13887_32519# 0.075021f
C20296 a_5093_45028# VDD 0.168437f
C20297 a_8685_43396# a_8952_43230# 0.003917f
C20298 a_2982_43646# a_19987_42826# 7.49e-20
C20299 a_3626_43646# a_19339_43156# 0.001776f
C20300 a_3080_42308# a_n2293_42282# 0.122474f
C20301 a_3422_30871# a_17303_42282# 0.063198f
C20302 a_14797_45144# a_11691_44458# 1.53e-19
C20303 a_3537_45260# a_n699_43396# 0.025655f
C20304 a_4574_45260# a_4223_44672# 9.56e-20
C20305 a_3065_45002# a_5343_44458# 3.26e-21
C20306 a_n357_42282# a_13483_43940# 1.74e-20
C20307 a_n2312_39304# a_n1630_35242# 0.002065f
C20308 a_5937_45572# a_7287_43370# 8.77e-22
C20309 a_12549_44172# a_20256_43172# 5.03e-21
C20310 a_1307_43914# a_11827_44484# 0.025083f
C20311 a_n2293_42834# a_n2661_43370# 0.038946f
C20312 a_n1059_45260# a_14539_43914# 0.029964f
C20313 a_6709_45028# a_n2661_44458# 2.58e-21
C20314 a_16751_46987# a_17829_46910# 2.45e-20
C20315 a_n2312_39304# a_n2661_45546# 0.022905f
C20316 a_12891_46348# a_12839_46116# 0.038804f
C20317 a_9863_46634# a_8199_44636# 2.9e-20
C20318 a_8667_46634# a_8953_45546# 0.002384f
C20319 a_8492_46660# a_5937_45572# 0.002914f
C20320 a_6575_47204# a_6511_45714# 2.63e-21
C20321 a_n1151_42308# a_8162_45546# 0.004489f
C20322 a_n443_46116# a_5024_45822# 0.009847f
C20323 a_4791_45118# a_4808_45572# 0.00122f
C20324 a_19692_46634# a_20202_43084# 0.172738f
C20325 a_19466_46812# a_11415_45002# 0.037852f
C20326 a_15227_44166# a_20820_30879# 5.72e-19
C20327 a_n2661_46098# a_n2956_38680# 0.123968f
C20328 a_n743_46660# a_1337_46116# 0.004248f
C20329 a_5807_45002# a_10586_45546# 0.001693f
C20330 a_2063_45854# a_10180_45724# 0.002207f
C20331 a_3080_42308# a_n3565_39590# 4.45e-21
C20332 a_n1853_43023# a_n3674_37592# 8.55e-20
C20333 a_n4318_38680# a_n4318_37592# 0.027855f
C20334 a_n1549_44318# VDD 0.200608f
C20335 a_n901_43156# a_n473_42460# 0.006054f
C20336 a_n1076_43230# a_n961_42308# 2.85e-19
C20337 a_n1736_43218# a_n1736_42282# 8.52e-19
C20338 a_10341_43396# a_15051_42282# 4.87e-20
C20339 a_12895_43230# a_13003_42852# 0.057222f
C20340 a_13635_43156# a_13814_43218# 0.007399f
C20341 a_13460_43230# a_13569_43230# 0.007416f
C20342 a_13113_42826# a_13291_42460# 1.73e-19
C20343 a_n2472_42826# a_n1630_35242# 2.09e-20
C20344 a_743_42282# a_3823_42558# 0.015894f
C20345 a_13507_46334# a_22521_40599# 2.03e-20
C20346 a_11827_44484# a_18579_44172# 0.045146f
C20347 a_2711_45572# a_15743_43084# 0.075024f
C20348 a_n357_42282# a_13678_32519# 1.42e-19
C20349 a_13249_42308# a_8685_43396# 0.03355f
C20350 a_584_46384# VDD 2.50905f
C20351 a_n237_47217# DATA[3] 0.0265f
C20352 a_10440_44484# a_n2661_43922# 0.006052f
C20353 a_10057_43914# a_n2661_42834# 0.053564f
C20354 a_8975_43940# a_11649_44734# 3.69e-19
C20355 a_9482_43914# a_10949_43914# 0.025292f
C20356 a_9290_44172# a_11229_43218# 0.002961f
C20357 a_n2312_38680# a_n2860_38778# 6.16e-19
C20358 a_3090_45724# a_14456_42282# 4.19e-20
C20359 a_327_47204# DATA[0] 0.353891f
C20360 a_n785_47204# DATA[1] 2.65e-19
C20361 a_7499_43078# a_10765_43646# 0.002149f
C20362 a_n2293_42834# a_2998_44172# 6.49e-20
C20363 a_20193_45348# a_20835_44721# 1.49e-19
C20364 a_n881_46662# a_327_44734# 3.44e-20
C20365 a_13507_46334# a_13017_45260# 2.21e-20
C20366 a_11735_46660# a_10490_45724# 2.75e-20
C20367 a_11901_46660# a_10193_42453# 4.59e-19
C20368 a_19594_46812# a_3357_43084# 4.56e-19
C20369 a_19900_46494# a_21137_46414# 3.02e-20
C20370 a_20075_46420# a_6945_45028# 1.64e-20
C20371 a_19553_46090# a_10809_44734# 5.04e-21
C20372 a_7920_46348# a_8034_45724# 0.032141f
C20373 a_6419_46155# a_6347_46155# 6.64e-19
C20374 a_13885_46660# a_2711_45572# 1.07e-21
C20375 a_11415_45002# a_20205_31679# 0.070403f
C20376 a_20202_43084# a_20692_30879# 3.23e-19
C20377 a_20916_46384# a_2437_43646# 0.010579f
C20378 a_9569_46155# a_5066_45546# 2.22e-20
C20379 a_10227_46804# a_15595_45028# 0.002256f
C20380 a_4883_46098# a_11787_45002# 1.41e-20
C20381 a_5379_42460# a_5337_42558# 8.44e-19
C20382 COMP_P a_5742_30871# 0.1094f
C20383 a_15095_43370# VDD 0.169652f
C20384 a_13678_32519# CAL_N 1.36e-19
C20385 a_2351_42308# a_6123_31319# 8.95e-21
C20386 a_5267_42460# a_5421_42558# 0.010303f
C20387 a_2903_42308# a_5932_42308# 8.68e-21
C20388 a_1606_42308# a_8515_42308# 1.34e-20
C20389 a_1755_42282# a_5934_30871# 3.43e-20
C20390 a_7640_43914# a_7499_43940# 0.049504f
C20391 a_n699_43396# a_1049_43396# 0.006702f
C20392 a_1414_42308# a_2675_43914# 0.305556f
C20393 a_1115_44172# a_2998_44172# 6.12e-20
C20394 a_n2840_43914# a_n4318_39768# 0.170372f
C20395 a_17517_44484# a_15493_43396# 7.93e-20
C20396 a_n1059_45260# a_7871_42858# 0.032582f
C20397 a_n2017_45002# a_7765_42852# 7.13e-20
C20398 a_n443_42852# a_5379_42460# 9.94e-21
C20399 a_n357_42282# a_6123_31319# 0.004292f
C20400 a_n755_45592# a_7227_42308# 3.68e-19
C20401 a_n2956_39304# a_n2946_39866# 0.004782f
C20402 a_n2956_38680# a_n3420_39616# 1.52e-19
C20403 a_5891_43370# a_5829_43940# 1.98e-19
C20404 a_742_44458# a_4235_43370# 3.35e-20
C20405 a_11901_46660# VDD 0.57548f
C20406 a_453_43940# a_895_43940# 0.420851f
C20407 a_2127_44172# a_2479_44172# 0.168988f
C20408 a_5164_46348# a_3357_43084# 7.34e-20
C20409 a_18479_47436# a_20766_44850# 0.007835f
C20410 a_8049_45260# a_8697_45822# 0.003995f
C20411 a_n2293_46098# a_1667_45002# 3.65e-20
C20412 a_8128_46384# a_n2661_43922# 4.1e-21
C20413 a_n443_46116# a_1467_44172# 0.031058f
C20414 a_6165_46155# a_2437_43646# 3.75e-20
C20415 a_4185_45028# a_20447_31679# 1.09e-20
C20416 a_1823_45246# a_n1059_45260# 0.021319f
C20417 a_18189_46348# a_18175_45572# 0.018402f
C20418 a_17715_44484# a_18479_45785# 9.75e-21
C20419 a_1138_42852# a_n913_45002# 0.032304f
C20420 a_n356_45724# a_1609_45822# 5.07e-20
C20421 a_n23_45546# a_n443_42852# 0.039956f
C20422 a_n755_45592# a_603_45572# 4.44e-20
C20423 a_n357_42282# a_1176_45572# 4.74e-21
C20424 a_18597_46090# a_20679_44626# 0.025074f
C20425 a_n784_42308# C4_P_btm 0.001073f
C20426 a_1606_42308# EN_VIN_BSTR_N 0.035204f
C20427 a_n237_47217# a_9313_45822# 0.063143f
C20428 a_n452_47436# a_n1435_47204# 2.2e-19
C20429 a_3815_47204# a_4007_47204# 0.224415f
C20430 a_n1151_42308# a_n443_46116# 0.099874f
C20431 a_3785_47178# a_4700_47436# 0.090466f
C20432 a_3381_47502# a_4791_45118# 3.29e-20
C20433 a_2063_45854# a_6545_47178# 2.04e-19
C20434 a_n2946_39866# a_n3565_39304# 0.001251f
C20435 a_n3420_39616# a_n3690_39392# 0.018295f
C20436 a_5934_30871# VDAC_P 0.029175f
C20437 a_n3690_39616# a_n3420_39072# 8.87e-19
C20438 a_n3565_39590# a_n2946_39072# 0.001251f
C20439 a_14097_32519# VDD 0.284675f
C20440 a_n4334_39616# a_n4064_39072# 7.91e-19
C20441 a_n2302_39866# a_n4209_39304# 0.001254f
C20442 a_n4209_39590# a_n2302_39072# 0.00133f
C20443 a_n4064_39616# a_n4334_39392# 0.001768f
C20444 a_22400_42852# RST_Z 0.059674f
C20445 a_n2661_43922# a_1847_42826# 3.92e-22
C20446 a_1307_43914# a_3581_42558# 4.31e-20
C20447 a_20679_44626# a_743_42282# 7.32e-21
C20448 a_20640_44752# a_20556_43646# 1.74e-20
C20449 a_11967_42832# a_4361_42308# 0.012085f
C20450 a_18287_44626# a_18249_42858# 2.07e-21
C20451 a_18248_44752# a_18817_42826# 8.42e-22
C20452 a_5891_43370# a_10835_43094# 1.38e-20
C20453 a_n2293_42834# COMP_P 8.54e-19
C20454 en_comp a_15890_42674# 1.81e-20
C20455 a_20512_43084# a_19268_43646# 2.18e-19
C20456 a_19279_43940# a_21259_43561# 5.61e-22
C20457 a_22485_44484# a_15743_43084# 0.003457f
C20458 a_n2661_42282# a_6452_43396# 0.011968f
C20459 a_3499_42826# a_3457_43396# 0.005429f
C20460 a_11823_42460# a_n2017_45002# 0.098619f
C20461 a_15599_45572# a_16789_45572# 2.56e-19
C20462 a_n755_45592# a_2903_45348# 1.85e-20
C20463 a_6598_45938# a_6171_45002# 0.002784f
C20464 a_6667_45809# a_6431_45366# 0.002877f
C20465 a_7227_45028# a_3232_43370# 9.21e-19
C20466 a_n443_42852# a_14797_45144# 5.7e-22
C20467 a_6511_45714# a_5205_44484# 5.08e-20
C20468 a_6472_45840# a_7276_45260# 6.14e-21
C20469 a_8049_45260# a_20567_45036# 3.41e-20
C20470 a_17478_45572# a_18175_45572# 0.001484f
C20471 a_8696_44636# a_18341_45572# 1.27e-19
C20472 a_15861_45028# a_18479_45785# 3.3e-20
C20473 a_2711_45572# a_10775_45002# 1.05e-19
C20474 a_n1641_46494# a_n2661_43922# 2.64e-22
C20475 a_4185_45028# a_5891_43370# 2.79e-19
C20476 a_13747_46662# a_19319_43548# 2.08e-20
C20477 a_13661_43548# a_18533_43940# 0.046643f
C20478 a_3218_45724# a_1423_45028# 2.67e-20
C20479 a_12861_44030# a_8685_43396# 0.007455f
C20480 a_n4064_37440# C3_P_btm 1.74e-19
C20481 a_n3420_37440# C1_P_btm 0.001902f
C20482 a_22469_39537# a_22609_38406# 0.198764f
C20483 a_22459_39145# a_22717_36887# 0.011525f
C20484 a_22521_39511# a_22705_37990# 0.004065f
C20485 a_n1613_43370# a_2959_46660# 0.187029f
C20486 a_2747_46873# a_3877_44458# 8.98e-21
C20487 a_5807_45002# a_n743_46660# 0.669712f
C20488 a_4915_47217# a_13607_46688# 0.082884f
C20489 a_9313_45822# a_8270_45546# 0.0271f
C20490 a_10227_46804# a_10150_46912# 0.236747f
C20491 a_20447_31679# VREF_GND 0.00199f
C20492 a_10341_43396# a_13749_43396# 9.69e-20
C20493 a_n659_45366# VDD 2.89e-19
C20494 a_n1557_42282# a_n2157_42858# 0.007773f
C20495 a_n2065_43946# a_n1630_35242# 4.6e-22
C20496 a_10807_43548# a_11229_43218# 6.49e-19
C20497 a_n1761_44111# a_564_42282# 1.16e-19
C20498 a_n97_42460# a_791_42968# 0.039538f
C20499 a_15095_43370# a_16137_43396# 1.7e-19
C20500 a_19479_31679# a_20567_45036# 3.97e-20
C20501 a_13661_43548# a_17595_43084# 2.01e-20
C20502 a_12549_44172# a_21195_42852# 2.16e-19
C20503 a_584_46384# a_n784_42308# 7.55e-22
C20504 a_15595_45028# a_1307_43914# 4.87e-19
C20505 a_15599_45572# a_14539_43914# 2.3e-21
C20506 a_8696_44636# a_8975_43940# 0.003372f
C20507 a_10180_45724# a_n2661_42834# 5.55e-20
C20508 a_n2956_38216# a_n2840_43914# 3.88e-19
C20509 a_21513_45002# a_21359_45002# 0.289039f
C20510 a_10227_46804# a_13569_43230# 2.95e-19
C20511 a_8199_44636# a_9801_43940# 0.048015f
C20512 a_8953_45546# a_9165_43940# 9.62e-19
C20513 a_8016_46348# a_10651_43940# 1.82e-19
C20514 a_413_45260# a_n2661_43370# 1.31746f
C20515 a_2711_45572# a_16789_44484# 2.48e-19
C20516 a_17715_44484# a_14021_43940# 3.95e-19
C20517 a_n1151_42308# a_n4318_37592# 4.12e-21
C20518 a_5257_43370# a_4361_42308# 7.33e-20
C20519 a_12549_44172# a_15015_46420# 7.35e-20
C20520 a_n971_45724# a_n452_45724# 0.03667f
C20521 a_n746_45260# a_n863_45724# 0.664707f
C20522 a_n2661_46098# a_n1423_46090# 0.021984f
C20523 a_11309_47204# a_2324_44458# 2.57e-20
C20524 a_9863_46634# a_765_45546# 3.07e-20
C20525 a_n1741_47186# a_n755_45592# 1.26e-21
C20526 a_5807_45002# a_11189_46129# 0.001199f
C20527 a_13661_43548# a_9290_44172# 0.00745f
C20528 a_n743_46660# a_3699_46348# 0.010053f
C20529 a_2959_46660# a_n2293_46098# 5.68e-21
C20530 a_2107_46812# a_1138_42852# 1.62e-19
C20531 a_6151_47436# a_13259_45724# 1.86e-20
C20532 a_11735_46660# a_12156_46660# 0.086708f
C20533 a_3090_45724# a_15559_46634# 2.45e-20
C20534 a_14976_45028# a_15368_46634# 0.097092f
C20535 a_n1925_46634# a_4419_46090# 3.01e-19
C20536 a_n2661_46634# a_6165_46155# 2.58e-20
C20537 a_n815_47178# a_n1099_45572# 3.58e-22
C20538 a_n2109_47186# a_1848_45724# 5.91e-22
C20539 a_n2497_47436# a_3218_45724# 2.25e-20
C20540 a_1847_42826# a_3445_43172# 4.44e-21
C20541 a_15743_43084# a_16877_42852# 1.77e-20
C20542 a_n97_42460# a_15051_42282# 0.049661f
C20543 a_12089_42308# a_5534_30871# 0.012295f
C20544 a_13113_42826# a_13460_43230# 0.051162f
C20545 a_3626_43646# a_3905_42308# 0.002949f
C20546 a_6293_42852# a_5932_42308# 8.47e-19
C20547 a_11649_44734# VDD 0.003396f
C20548 a_3457_43396# a_3318_42354# 8.91e-20
C20549 a_6197_43396# a_6171_42473# 5.91e-20
C20550 a_413_45260# a_2998_44172# 0.161528f
C20551 a_n2017_45002# a_n1644_44306# 0.00478f
C20552 a_17668_45572# a_17737_43940# 2.42e-20
C20553 a_13259_45724# a_13837_43396# 0.007401f
C20554 a_9290_44172# a_10835_43094# 0.172486f
C20555 a_4185_45028# a_17595_43084# 1.06e-20
C20556 a_n443_42852# a_7287_43370# 0.010578f
C20557 a_2680_45002# a_2127_44172# 2.9e-20
C20558 a_2382_45260# a_2479_44172# 0.00555f
C20559 a_n2312_39304# a_n3607_39392# 5.97e-20
C20560 a_n2293_45010# a_n1287_44306# 8.54e-19
C20561 a_19256_45572# a_15493_43396# 2.21e-21
C20562 a_19321_45002# a_20712_42282# 2.03e-21
C20563 a_19431_45546# a_19478_44306# 9.3e-21
C20564 a_3429_45260# a_1414_42308# 1.27e-22
C20565 a_3357_43084# a_3499_42826# 0.134316f
C20566 a_5343_44458# a_6298_44484# 0.128602f
C20567 a_4223_44672# a_5883_43914# 0.967973f
C20568 a_15861_45028# a_14021_43940# 3.03e-20
C20569 a_2324_44458# a_3935_42891# 6.13e-22
C20570 a_18597_46090# a_20528_45572# 0.03478f
C20571 a_12549_44172# a_16333_45814# 3.97e-22
C20572 a_19466_46812# a_13259_45724# 5.7e-20
C20573 a_n1151_42308# a_3537_45260# 4.52e-19
C20574 a_4915_47217# a_413_45260# 7.6e-19
C20575 a_n443_46116# a_327_44734# 4.41e-19
C20576 a_15673_47210# a_3357_43084# 3.29e-19
C20577 a_16023_47582# a_2437_43646# 0.00865f
C20578 a_16327_47482# a_22223_45572# 2.78e-19
C20579 a_3483_46348# a_11133_46155# 0.001334f
C20580 a_7920_46348# a_8016_46348# 0.318386f
C20581 a_12741_44636# a_10809_44734# 0.088683f
C20582 a_4185_45028# a_9290_44172# 4.71e-19
C20583 a_20820_30879# a_22959_46124# 0.00389f
C20584 a_n237_47217# a_7705_45326# 5.12e-19
C20585 a_n971_45724# a_8953_45002# 1.78e-20
C20586 a_15928_47570# a_15903_45785# 6.16e-21
C20587 a_2063_45854# a_4927_45028# 5.82e-19
C20588 a_5732_46660# a_5907_45546# 1.37e-19
C20589 a_5907_46634# a_6194_45824# 8.2e-20
C20590 a_n743_46660# a_15143_45578# 7.03e-21
C20591 a_13507_46334# a_20107_45572# 1.59e-20
C20592 a_20894_47436# a_20623_45572# 2.94e-21
C20593 a_3080_42308# C4_P_btm 5.72e-19
C20594 a_n1177_43370# VDD 0.354704f
C20595 a_16795_42852# a_4958_30871# 0.001047f
C20596 a_n2840_42282# a_n4318_37592# 0.037154f
C20597 a_14097_32519# a_n784_42308# 0.005039f
C20598 a_n4318_38216# a_n2104_42282# 7.75e-19
C20599 a_n2472_42282# a_n3674_38216# 0.040147f
C20600 a_9306_43218# a_5934_30871# 4.18e-20
C20601 a_n3674_39304# a_n4209_39304# 0.059449f
C20602 a_526_44458# a_8515_42308# 3.38e-20
C20603 a_n1925_42282# a_5934_30871# 3.98e-20
C20604 a_n443_42852# a_13157_43218# 4.11e-20
C20605 a_4185_45028# a_21887_42336# 8e-20
C20606 a_16922_45042# a_14401_32519# 1.06e-19
C20607 a_5111_44636# a_9885_43646# 0.010527f
C20608 a_n2661_43370# a_n2012_43396# 1.88e-20
C20609 a_n2661_42834# a_5013_44260# 0.021017f
C20610 a_20640_44752# a_20980_44850# 0.027606f
C20611 a_20159_44458# a_3422_30871# 2.52e-20
C20612 a_n2293_42834# a_1568_43370# 0.037512f
C20613 a_1307_43914# a_8147_43396# 2.66e-20
C20614 a_17970_44736# a_17737_43940# 1.63e-19
C20615 a_17767_44458# a_17973_43940# 0.012863f
C20616 a_n2661_43922# a_5244_44056# 2.61e-20
C20617 a_n2293_43922# a_3905_42865# 2.09e-20
C20618 a_19778_44110# a_19808_44306# 0.004261f
C20619 a_18587_45118# a_18533_43940# 6.8e-22
C20620 a_479_46660# VDD 1.63e-19
C20621 a_n357_42282# a_15597_42852# 0.009386f
C20622 a_n913_45002# a_17499_43370# 2.4e-20
C20623 a_n1059_45260# a_17324_43396# 0.003177f
C20624 a_11453_44696# a_16112_44458# 8.57e-20
C20625 a_12594_46348# a_13163_45724# 0.053634f
C20626 a_13759_46122# a_11823_42460# 1.12e-19
C20627 a_2324_44458# a_10490_45724# 0.015189f
C20628 a_4651_46660# a_5009_45028# 6.47e-22
C20629 a_6755_46942# a_14180_45002# 2.19e-22
C20630 a_5937_45572# a_9241_45822# 0.010703f
C20631 a_8953_45546# a_8697_45822# 0.006215f
C20632 a_8199_44636# a_10210_45822# 0.012124f
C20633 a_4883_46098# a_18287_44626# 1.92e-21
C20634 a_10903_43370# a_13904_45546# 0.081466f
C20635 a_11735_46660# a_6171_45002# 1.67e-20
C20636 a_11813_46116# a_3232_43370# 6.78e-22
C20637 a_16388_46812# a_3357_43084# 5.22e-20
C20638 a_n1613_43370# a_n699_43396# 0.008801f
C20639 a_20841_46902# a_20273_45572# 5.17e-21
C20640 a_20623_46660# a_20107_45572# 1.34e-20
C20641 a_20411_46873# a_20623_45572# 6.29e-19
C20642 a_11415_45002# a_16147_45260# 0.058206f
C20643 a_n881_46662# a_4223_44672# 1.75e-20
C20644 a_3090_45724# a_3065_45002# 0.475346f
C20645 a_2609_46660# a_n2661_43370# 7.75e-21
C20646 a_526_44458# a_2711_45572# 0.392618f
C20647 a_22959_42860# VDD 0.30747f
C20648 a_19332_42282# a_19511_42282# 0.174683f
C20649 a_18214_42558# a_18548_42308# 2.43e-19
C20650 a_22223_42860# RST_Z 5.92e-20
C20651 a_17303_42282# a_7174_31319# 0.027048f
C20652 a_5742_30871# a_n4209_39304# 6.2e-21
C20653 a_20623_43914# a_14021_43940# 1.48e-19
C20654 a_n1059_45260# a_1184_42692# 0.019924f
C20655 a_n913_45002# a_1576_42282# 0.001393f
C20656 a_n2017_45002# a_961_42354# 0.00519f
C20657 a_9028_43914# a_9165_43940# 0.126609f
C20658 a_1467_44172# a_1049_43396# 0.002443f
C20659 a_1115_44172# a_1568_43370# 1.06e-19
C20660 a_n1761_44111# a_n1557_42282# 0.018977f
C20661 a_1414_42308# a_1209_43370# 0.003338f
C20662 a_9313_44734# a_18783_43370# 8.63e-20
C20663 a_10903_43370# CLK 0.018377f
C20664 a_742_44458# a_791_42968# 3.18e-19
C20665 a_11827_44484# a_13635_43156# 3.57e-21
C20666 a_14673_44172# a_14358_43442# 0.00447f
C20667 en_comp a_n3674_37592# 0.050998f
C20668 a_n2810_45028# a_n1630_35242# 4.11e-19
C20669 a_17583_46090# VDD 0.23578f
C20670 a_3905_42865# a_n97_42460# 0.071125f
C20671 a_15682_46116# RST_Z 8.37e-21
C20672 a_n4318_39768# a_n4318_39304# 0.042825f
C20673 a_n3674_39768# a_n2840_43370# 0.006059f
C20674 a_453_43940# a_458_43396# 9.25e-20
C20675 a_3357_43084# a_3318_42354# 2.7e-19
C20676 a_n967_45348# a_n327_42558# 5.76e-21
C20677 a_n2293_42834# a_4743_43172# 2.14e-19
C20678 a_n1925_42282# a_4185_45348# 1.16e-20
C20679 a_13163_45724# a_15037_45618# 7.32e-23
C20680 a_12861_44030# a_19741_43940# 2.77e-20
C20681 a_584_46384# a_3080_42308# 0.010326f
C20682 a_n971_45724# a_3626_43646# 4.16e-20
C20683 a_n1076_46494# a_n1177_44458# 3.46e-22
C20684 a_n2293_46098# a_n699_43396# 0.001069f
C20685 a_10193_42453# a_8696_44636# 0.225102f
C20686 a_n2810_45572# a_n2956_37592# 0.048284f
C20687 a_n881_46662# a_15493_43940# 4.43e-21
C20688 a_2324_44458# a_14976_45348# 0.002969f
C20689 a_15368_46634# a_15433_44458# 1.7e-19
C20690 a_n2293_46634# a_3499_42826# 0.022726f
C20691 a_n2956_39768# a_n2661_42282# 6.98e-20
C20692 a_12549_44172# a_15493_43396# 0.079226f
C20693 a_n2293_45546# a_n1059_45260# 0.076047f
C20694 a_n1099_45572# a_n2661_45010# 7.2e-21
C20695 a_1138_42852# a_n2661_44458# 0.026505f
C20696 a_8697_45822# a_8791_45572# 1.26e-19
C20697 a_n1435_47204# a_33_46660# 3.84e-20
C20698 a_3754_38470# a_8530_39574# 0.059662f
C20699 a_14311_47204# a_n743_46660# 6.88e-21
C20700 a_7754_40130# VDAC_P 0.334598f
C20701 a_2063_45854# a_3877_44458# 0.024649f
C20702 a_n443_46116# a_3177_46902# 0.019328f
C20703 a_2905_45572# a_3686_47026# 1.64e-19
C20704 a_n4334_39616# VDD 0.385881f
C20705 a_7754_39964# VDAC_N 2.46e-19
C20706 a_n3565_39304# C1_P_btm 1.3e-20
C20707 a_n4064_39072# C5_P_btm 2.13e-20
C20708 a_18597_46090# a_19594_46812# 6.44e-19
C20709 a_19386_47436# a_19321_45002# 0.086877f
C20710 VDAC_Pi a_6886_37412# 0.259481f
C20711 a_n971_45724# a_5275_47026# 6.84e-21
C20712 a_n3420_38528# a_n923_35174# 0.002965f
C20713 a_20447_31679# a_22469_40625# 1.91e-20
C20714 a_19479_31679# a_22521_39511# 2.38e-20
C20715 a_10949_43914# a_10796_42968# 9.1e-19
C20716 a_10807_43548# a_10835_43094# 0.02952f
C20717 a_10729_43914# a_10991_42826# 1.29e-20
C20718 a_19741_43940# a_19700_43370# 5.56e-19
C20719 a_19963_31679# a_22521_40055# 8.31e-21
C20720 a_10057_43914# a_9885_42558# 4.04e-21
C20721 a_3905_42865# a_3935_43218# 0.004982f
C20722 a_n2661_42834# a_196_42282# 1.99e-22
C20723 a_n2293_43922# a_n961_42308# 1.63e-19
C20724 a_18184_42460# a_20712_42282# 3.18e-19
C20725 a_8696_44636# VDD 1.12228f
C20726 a_14401_32519# a_15743_43084# 0.017308f
C20727 a_18494_42460# a_20107_42308# 0.035023f
C20728 a_5807_45002# a_4361_42308# 2.93e-22
C20729 a_n971_45724# a_8649_43218# 3.91e-20
C20730 a_8162_45546# a_4223_44672# 4.14e-21
C20731 a_5937_45572# a_5841_44260# 1.15e-20
C20732 a_413_45260# a_4574_45260# 7.73e-20
C20733 a_19321_45002# a_20556_43646# 4.6e-19
C20734 a_n1613_43370# a_n4318_38680# 1.09e-19
C20735 a_n443_42852# a_n23_44458# 0.002324f
C20736 a_2324_44458# a_6453_43914# 0.010794f
C20737 a_4883_46098# a_9127_43156# 0.011077f
C20738 a_3483_46348# a_12429_44172# 9.13e-22
C20739 a_10227_46804# a_13113_42826# 0.159547f
C20740 a_2382_45260# a_2680_45002# 0.023953f
C20741 a_n863_45724# a_n310_44484# 1.13e-19
C20742 a_2711_45572# a_17970_44736# 6.8e-21
C20743 a_10150_46912# a_10467_46802# 0.102355f
C20744 a_7927_46660# a_6755_46942# 0.036549f
C20745 a_5257_43370# a_6086_46660# 1.63e-19
C20746 a_n1435_47204# a_12005_46116# 9.73e-21
C20747 a_13717_47436# a_10903_43370# 0.001667f
C20748 a_n881_46662# a_12741_44636# 7.98e-20
C20749 a_13507_46334# a_3483_46348# 1.37e-19
C20750 a_19321_45002# a_19551_46910# 0.009214f
C20751 a_19594_46812# a_19123_46287# 0.002216f
C20752 a_13747_46662# a_20411_46873# 3.16e-20
C20753 a_13661_43548# a_20273_46660# 5.45e-20
C20754 a_13381_47204# a_12594_46348# 3.26e-21
C20755 a_3067_47026# a_3090_45724# 1.04e-20
C20756 a_7577_46660# a_6682_46987# 3.94e-20
C20757 a_14401_32519# a_1606_42308# 0.001872f
C20758 a_n1177_43370# a_n784_42308# 2.67e-21
C20759 a_5649_42852# a_9127_43156# 8.16e-20
C20760 a_n1076_43230# a_685_42968# 4.61e-19
C20761 a_n13_43084# a_421_43172# 0.003935f
C20762 a_3080_42308# a_14097_32519# 1.75e-20
C20763 a_15743_43084# a_18817_42826# 0.003018f
C20764 a_18783_43370# a_18599_43230# 6.07e-19
C20765 a_743_42282# a_10341_42308# 0.020229f
C20766 a_19268_43646# a_18249_42858# 7.34e-20
C20767 a_n1177_44458# VDD 0.347966f
C20768 a_n4318_39768# a_n4334_40480# 0.002408f
C20769 a_n3674_39768# a_n4315_30879# 7.29e-19
C20770 a_8685_43396# a_8495_42852# 2.66e-19
C20771 a_4185_45028# a_13467_32519# 0.033397f
C20772 a_n2661_43370# a_2779_44458# 1.59e-19
C20773 a_8953_45002# a_9313_44734# 0.001727f
C20774 a_20567_45036# a_20193_45348# 0.037561f
C20775 a_16922_45042# a_20205_45028# 0.0038f
C20776 a_5111_44636# a_n2661_43922# 0.061031f
C20777 a_13249_42308# a_13483_43940# 0.193724f
C20778 a_10193_42453# a_20365_43914# 1.25e-20
C20779 a_3232_43370# a_9159_44484# 0.005178f
C20780 a_11827_44484# a_22223_45036# 0.179208f
C20781 a_3357_43084# a_20640_44752# 4.03e-21
C20782 a_16327_47482# a_19647_42308# 1.59e-19
C20783 a_21513_45002# a_19279_43940# 0.003201f
C20784 a_21363_45546# a_21398_44850# 1.78e-21
C20785 a_n2293_42834# a_5883_43914# 0.015714f
C20786 a_n2956_38216# a_n4318_39304# 0.023138f
C20787 a_7499_43078# a_11341_43940# 0.00321f
C20788 a_n2293_46634# a_3318_42354# 2.67e-19
C20789 a_n743_46660# a_n755_45592# 0.020454f
C20790 a_n2438_43548# a_n357_42282# 0.026249f
C20791 a_n2293_46634# a_3316_45546# 0.067277f
C20792 a_19466_46812# a_18189_46348# 0.001238f
C20793 a_14035_46660# a_10903_43370# 2e-19
C20794 a_n133_46660# a_310_45028# 8.97e-20
C20795 a_7927_46660# a_8049_45260# 7.61e-20
C20796 a_15227_44166# a_18819_46122# 0.288885f
C20797 a_765_45546# a_6165_46155# 6.78e-20
C20798 a_4883_46098# a_13904_45546# 1.69e-20
C20799 a_10227_46804# a_10907_45822# 2.47e-19
C20800 a_13607_46688# a_10809_44734# 0.002497f
C20801 a_15009_46634# a_6945_45028# 5.03e-20
C20802 a_6969_46634# a_5066_45546# 1.41e-19
C20803 a_171_46873# a_n1099_45572# 5.56e-21
C20804 a_33_46660# a_380_45546# 1.08e-19
C20805 a_5649_42852# a_17124_42282# 1.31e-19
C20806 a_743_42282# a_18057_42282# 0.008889f
C20807 a_8605_42826# a_8515_42308# 0.001559f
C20808 a_8387_43230# a_5934_30871# 0.001004f
C20809 a_4361_42308# a_16197_42308# 1.2e-19
C20810 a_21487_43396# a_17303_42282# 4.02e-21
C20811 a_4190_30871# a_18907_42674# 0.040515f
C20812 a_n2293_42282# a_196_42282# 4.89e-19
C20813 a_20365_43914# VDD 0.261299f
C20814 a_8696_44636# a_16137_43396# 2.49e-20
C20815 a_n2312_40392# CLK_DATA 0.213071f
C20816 a_n4318_40392# a_n3674_39768# 0.026429f
C20817 a_742_44458# a_3905_42865# 0.002336f
C20818 a_n2661_44458# a_n4318_39768# 8.38e-19
C20819 a_n2017_45002# a_2982_43646# 0.023101f
C20820 a_1307_43914# a_10555_43940# 0.001112f
C20821 a_17339_46660# a_18214_42558# 8.1e-20
C20822 a_2779_44458# a_2998_44172# 0.007931f
C20823 a_4883_46098# CLK 0.032195f
C20824 a_n357_42282# a_18083_42858# 0.026806f
C20825 a_16922_45042# a_15682_43940# 0.001439f
C20826 a_n699_43396# a_2675_43914# 0.015641f
C20827 a_n2293_43922# a_12553_44484# 1.41e-19
C20828 a_5147_45002# a_n97_42460# 0.085495f
C20829 a_3357_43084# a_6197_43396# 0.001107f
C20830 a_n2293_46634# a_13777_45326# 1.56e-21
C20831 a_4791_45118# a_n699_43396# 0.024838f
C20832 a_19466_46812# a_17478_45572# 2.38e-21
C20833 a_12861_44030# a_18545_45144# 1.5e-19
C20834 a_13507_46334# a_17719_45144# 8.16e-21
C20835 a_16327_47482# a_11691_44458# 0.536141f
C20836 a_n743_46660# a_13017_45260# 6.48e-21
C20837 a_19553_46090# a_19443_46116# 0.097745f
C20838 a_10809_44734# a_16375_45002# 6.42e-20
C20839 a_2107_46812# a_7229_43940# 4.89e-21
C20840 a_n2497_47436# a_n1190_44850# 1.37e-19
C20841 a_167_45260# a_3175_45822# 2.8e-19
C20842 a_1823_45246# a_5263_45724# 2e-20
C20843 a_n2293_46098# a_5024_45822# 0.001497f
C20844 a_11453_44696# a_13807_45067# 2e-19
C20845 a_18597_46090# a_18494_42460# 3.29e-19
C20846 a_18479_47436# a_21005_45260# 0.015257f
C20847 a_n881_46662# a_n2293_42834# 4.05e-20
C20848 a_8145_46902# a_3357_43084# 2.87e-21
C20849 a_3699_46634# a_3065_45002# 8.84e-21
C20850 a_2959_46660# a_3429_45260# 5.07e-19
C20851 a_2713_42308# a_7174_31319# 4.88e-21
C20852 a_n1630_35242# a_n2302_40160# 1.59e-19
C20853 a_n1991_42858# VDD 0.575656f
C20854 a_13467_32519# VREF_GND 0.048151f
C20855 a_11691_44458# a_16855_43396# 4.36e-20
C20856 a_n1059_45260# a_5193_42852# 0.004497f
C20857 a_20820_30879# C7_N_btm 0.184297f
C20858 a_18494_42460# a_743_42282# 0.476713f
C20859 a_14537_43396# a_5534_30871# 2.84e-19
C20860 a_13556_45296# a_15567_42826# 4.05e-21
C20861 a_19615_44636# a_19319_43548# 0.001036f
C20862 a_11967_42832# a_18533_43940# 4.96e-19
C20863 a_n2661_42834# a_4699_43561# 6.89e-20
C20864 a_6109_44484# a_6293_42852# 3.01e-21
C20865 a_n2293_42834# a_133_43172# 4.3e-19
C20866 a_9313_44734# a_3626_43646# 2.37e-19
C20867 a_22000_46634# EN_OFFSET_CAL 3.46e-20
C20868 a_n2956_38216# a_n4334_40480# 6.67e-19
C20869 a_7499_43078# a_10723_42308# 0.029878f
C20870 a_2711_45572# a_13163_45724# 0.006905f
C20871 a_2324_44458# a_6171_45002# 2.73828f
C20872 a_10809_44734# a_413_45260# 0.333257f
C20873 a_19321_45002# a_20980_44850# 6.29e-21
C20874 a_13747_46662# a_3422_30871# 1.93e-19
C20875 a_5066_45546# a_3357_43084# 0.033559f
C20876 a_8049_45260# a_20528_45572# 0.004485f
C20877 a_10903_43370# a_10951_45334# 0.005295f
C20878 a_11387_46155# a_11787_45002# 3.57e-19
C20879 a_12861_44030# a_13483_43940# 1.39e-19
C20880 a_13259_45724# a_16147_45260# 0.033344f
C20881 a_3090_45724# a_6298_44484# 0.013998f
C20882 a_5257_43370# a_5891_43370# 0.001693f
C20883 a_3877_44458# a_n2661_42834# 2.79e-19
C20884 a_2063_45854# a_8128_46384# 0.032153f
C20885 a_3160_47472# a_n881_46662# 0.070909f
C20886 a_n1151_42308# a_n1613_43370# 1.19311f
C20887 a_n3565_39590# a_n4064_37440# 0.031724f
C20888 a_16763_47508# a_10227_46804# 0.070681f
C20889 a_13717_47436# a_4883_46098# 2.67e-19
C20890 a_6123_31319# VIN_P 0.01057f
C20891 a_1343_38525# VDAC_Ni 0.006713f
C20892 a_16588_47582# a_17591_47464# 0.001438f
C20893 a_5742_30871# C6_N_btm 0.170624f
C20894 a_13487_47204# a_13507_46334# 1.68e-19
C20895 a_21613_42308# a_22521_40599# 2.02e-20
C20896 a_9377_42558# VDD 0.007808f
C20897 a_16327_47482# a_18479_47436# 0.723416f
C20898 a_n3420_39616# a_n3420_37440# 0.053603f
C20899 a_n4064_39616# a_n3565_37414# 0.029074f
C20900 a_n4209_38216# a_n3565_38216# 6.80743f
C20901 a_11341_43940# a_15781_43660# 4.59e-21
C20902 a_5891_43370# a_9114_42852# 1.43e-19
C20903 a_14539_43914# a_18861_43218# 4.42e-20
C20904 a_n2267_43396# a_n1557_42282# 1.4e-20
C20905 a_n97_42460# a_4093_43548# 0.028602f
C20906 a_15682_43940# a_15743_43084# 6.12e-19
C20907 en_comp a_n2302_39072# 4.43e-20
C20908 a_7227_45028# VDD 0.501104f
C20909 a_15493_43396# a_16977_43638# 0.018523f
C20910 a_3499_42826# a_743_42282# 1.89e-19
C20911 a_14021_43940# a_15095_43370# 0.001284f
C20912 a_11967_42832# a_17595_43084# 0.0964f
C20913 a_3090_45724# a_10555_44260# 0.041801f
C20914 a_11453_44696# a_17499_43370# 8.56e-21
C20915 a_10907_45822# a_1307_43914# 5.29e-20
C20916 a_8162_45546# a_n2293_42834# 0.001469f
C20917 a_n2956_38216# a_n2661_44458# 0.009784f
C20918 a_9290_44172# a_11967_42832# 0.0995f
C20919 a_20623_45572# a_19963_31679# 8.99e-21
C20920 a_768_44030# a_9803_43646# 5.37e-20
C20921 a_19692_46634# a_20623_43914# 0.007357f
C20922 a_n2956_39304# a_n2293_43922# 4.52e-20
C20923 a_4185_45028# a_22315_44484# 0.002812f
C20924 a_16327_47482# a_4190_30871# 0.335014f
C20925 a_n971_45724# a_8037_42858# 7.81e-19
C20926 a_n2293_46634# a_6197_43396# 0.05355f
C20927 a_15227_44166# a_11341_43940# 0.04747f
C20928 a_12861_44030# a_13678_32519# 6.9e-20
C20929 a_21188_45572# a_3357_43084# 0.057919f
C20930 a_20107_45572# a_21297_45572# 2.56e-19
C20931 a_n2472_45546# a_n2433_44484# 3.17e-20
C20932 a_2711_45572# a_16501_45348# 4.66e-19
C20933 a_2324_44458# a_14673_44172# 0.015622f
C20934 EN_VIN_BSTR_P VIN_P 1.41696f
C20935 C5_P_btm VDD 0.267489f
C20936 C0_P_btm C7_N_btm 4.2e-19
C20937 C1_P_btm C8_N_btm 7.93e-19
C20938 C3_P_btm C10_N_btm 0.002331f
C20939 C0_dummy_P_btm C6_N_btm 2.49e-19
C20940 C0_N_btm C4_N_btm 0.138884f
C20941 C0_dummy_N_btm C5_N_btm 0.11443f
C20942 C1_N_btm C3_N_btm 7.40325f
C20943 a_n2109_47186# a_4185_45028# 1.33e-19
C20944 a_n971_45724# a_167_45260# 1.89e-19
C20945 a_n1741_47186# a_3483_46348# 4.84e-20
C20946 a_4883_46098# a_14035_46660# 0.019262f
C20947 a_16327_47482# a_17829_46910# 7.11e-21
C20948 a_5807_45002# a_6086_46660# 1.02e-19
C20949 a_n237_47217# a_1823_45246# 0.370766f
C20950 a_n1151_42308# a_n2293_46098# 0.040266f
C20951 a_11309_47204# a_11186_47026# 0.004771f
C20952 a_n881_46662# a_13607_46688# 2.29e-20
C20953 a_13507_46334# a_14513_46634# 9.96e-20
C20954 a_16023_47582# a_765_45546# 0.006051f
C20955 a_2107_46812# a_5907_46634# 0.003718f
C20956 a_n1925_46634# a_7411_46660# 0.047823f
C20957 a_n2661_46634# a_8492_46660# 0.009944f
C20958 a_584_46384# a_n901_46420# 3.34e-19
C20959 a_11599_46634# a_20411_46873# 0.00162f
C20960 a_10227_46804# a_14226_46660# 4.83e-20
C20961 a_18597_46090# a_16388_46812# 0.011997f
C20962 a_13717_47436# a_21188_46660# 2.12e-21
C20963 a_n97_42460# a_5457_43172# 4.93e-20
C20964 a_15743_43084# a_22223_43396# 0.004521f
C20965 a_5009_45028# VDD 0.151712f
C20966 a_8685_43396# a_9127_43156# 0.01312f
C20967 a_2982_43646# a_19164_43230# 1.37e-20
C20968 a_18114_32519# VDAC_N 0.001372f
C20969 a_3422_30871# a_4958_30871# 0.101017f
C20970 a_14537_43396# a_11691_44458# 0.092307f
C20971 a_3537_45260# a_4223_44672# 0.1907f
C20972 a_n357_42282# a_12429_44172# 5.79e-21
C20973 a_n2312_40392# a_n1630_35242# 0.033733f
C20974 a_5937_45572# a_6547_43396# 6.63e-19
C20975 a_17339_46660# a_16823_43084# 7.42e-19
C20976 a_13661_43548# a_18695_43230# 2.15e-19
C20977 a_16019_45002# a_11827_44484# 4.4e-20
C20978 a_8270_45546# a_7871_42858# 8.9e-21
C20979 a_n2017_45002# a_14539_43914# 0.01532f
C20980 a_7229_43940# a_n2661_44458# 0.028622f
C20981 a_2063_45854# a_10053_45546# 1.55e-19
C20982 a_n881_46662# a_16375_45002# 2.62e-19
C20983 a_16434_46987# a_17829_46910# 4.36e-20
C20984 a_n2312_40392# a_n2661_45546# 7.42e-20
C20985 a_n2312_39304# a_n2810_45572# 0.044713f
C20986 a_2107_46812# a_739_46482# 5.16e-20
C20987 a_8667_46634# a_5937_45572# 0.001106f
C20988 a_8492_46660# a_8199_44636# 2.51e-19
C20989 a_6851_47204# a_6598_45938# 1.17e-21
C20990 a_6575_47204# a_6472_45840# 6.84e-21
C20991 a_4791_45118# a_5024_45822# 1.87e-20
C20992 a_17609_46634# a_12741_44636# 5.71e-21
C20993 a_19466_46812# a_20202_43084# 2.86e-21
C20994 a_16751_46987# a_765_45546# 1.47e-19
C20995 a_n2661_46098# a_n2956_39304# 0.008823f
C20996 a_n743_46660# a_835_46155# 4.14e-19
C20997 a_15227_44166# a_22591_46660# 1.6e-20
C20998 a_16388_46812# a_19123_46287# 4.8e-20
C20999 a_16721_46634# a_18285_46348# 2.92e-20
C21000 a_19594_46812# a_8049_45260# 9.33e-20
C21001 a_16327_47482# a_n443_42852# 2.73e-21
C21002 a_13507_46334# a_n357_42282# 0.001222f
C21003 a_3422_30871# VCM 1.12142f
C21004 a_n2840_42826# a_n1630_35242# 2.09e-20
C21005 a_n2157_42858# a_n3674_37592# 0.001748f
C21006 a_n3674_39304# a_n4318_37592# 0.023516f
C21007 a_14955_43396# a_15486_42560# 1.53e-19
C21008 a_n1331_43914# VDD 0.203823f
C21009 a_n901_43156# a_n961_42308# 0.002229f
C21010 a_10341_43396# a_14113_42308# 1.45e-20
C21011 a_13113_42826# a_13003_42852# 0.097745f
C21012 a_12545_42858# a_13291_42460# 1.52e-19
C21013 a_5649_42852# a_1755_42282# 0.023826f
C21014 a_743_42282# a_3318_42354# 0.01411f
C21015 a_7499_43078# a_10341_43396# 0.061281f
C21016 a_10193_42453# a_14205_43396# 5.63e-21
C21017 a_20820_30879# COMP_P 8.52e-20
C21018 a_13507_46334# CAL_N 0.004017f
C21019 a_1307_43914# a_n2661_42282# 0.042336f
C21020 a_11827_44484# a_18245_44484# 1.94e-19
C21021 SMPL_ON_P VIN_P 0.587766f
C21022 a_2711_45572# a_18783_43370# 6.16e-20
C21023 a_2124_47436# VDD 0.086403f
C21024 a_10334_44484# a_n2661_43922# 0.008746f
C21025 a_10440_44484# a_n2661_42834# 7.54e-20
C21026 a_8975_43940# a_9159_44484# 0.00805f
C21027 a_9482_43914# a_10729_43914# 0.047853f
C21028 a_16922_45042# a_20512_43084# 0.055985f
C21029 a_n237_47217# DATA[2] 7.36e-22
C21030 a_n755_45592# a_4361_42308# 0.035265f
C21031 a_n2312_38680# a_n2302_38778# 0.161815f
C21032 a_n785_47204# DATA[0] 0.598846f
C21033 a_n23_47502# DATA[1] 1.93e-20
C21034 a_n2293_42834# a_2889_44172# 3.27e-21
C21035 a_20193_45348# a_20679_44626# 0.017743f
C21036 a_10467_46802# a_10907_45822# 4.68e-20
C21037 a_10623_46897# a_10210_45822# 3.91e-20
C21038 a_n443_46116# a_n2293_42834# 9.36e-19
C21039 a_768_44030# a_n913_45002# 2.6e-19
C21040 a_n881_46662# a_413_45260# 0.026808f
C21041 a_n1613_43370# a_327_44734# 3.68e-20
C21042 a_11813_46116# a_10193_42453# 0.02832f
C21043 a_19321_45002# a_3357_43084# 0.030763f
C21044 a_19900_46494# a_20708_46348# 2.56e-19
C21045 a_19335_46494# a_6945_45028# 1.78e-20
C21046 a_18985_46122# a_10809_44734# 9.49e-20
C21047 a_3483_46348# a_10586_45546# 0.099824f
C21048 a_765_45546# a_n23_45546# 8.66e-20
C21049 a_3090_45724# a_5437_45600# 5.24e-20
C21050 a_20202_43084# a_20205_31679# 1.27e-19
C21051 a_20916_46384# a_21513_45002# 1.63e-20
C21052 a_22365_46825# a_20692_30879# 7.03e-19
C21053 a_9625_46129# a_5066_45546# 1.5e-20
C21054 a_10227_46804# a_15415_45028# 0.001754f
C21055 a_4883_46098# a_10951_45334# 2.01e-20
C21056 a_13887_32519# VDAC_N 2.99e-19
C21057 a_2123_42473# a_6123_31319# 8.95e-21
C21058 a_5379_42460# a_4921_42308# 0.033756f
C21059 a_5267_42460# a_5337_42558# 0.011552f
C21060 a_14205_43396# VDD 0.311811f
C21061 a_5649_42852# VDAC_P 3.45e-20
C21062 a_1606_42308# a_5934_30871# 0.095492f
C21063 a_2713_42308# a_5932_42308# 4.34e-21
C21064 a_13467_32519# a_22469_40625# 1.21e-20
C21065 a_n2293_43922# a_12710_44260# 9.27e-19
C21066 a_n699_43396# a_1209_43370# 0.004475f
C21067 a_1414_42308# a_895_43940# 0.208524f
C21068 a_11967_42832# a_10807_43548# 1.1e-20
C21069 a_10193_42453# a_22400_42852# 3.3e-21
C21070 a_18989_43940# a_18533_43940# 0.001685f
C21071 a_17517_44484# a_19328_44172# 7.19e-21
C21072 a_n913_45002# a_5755_42852# 1.7e-20
C21073 a_n1059_45260# a_7227_42852# 0.005565f
C21074 a_n2017_45002# a_7871_42858# 1.28e-19
C21075 a_n443_42852# a_5267_42460# 7.84e-22
C21076 a_n755_45592# a_6761_42308# 2.19e-19
C21077 a_n357_42282# a_7227_42308# 7.15e-20
C21078 a_n2956_39304# a_n3420_39616# 9.34e-19
C21079 a_5891_43370# a_5745_43940# 2.82e-19
C21080 a_949_44458# a_1756_43548# 0.001231f
C21081 a_742_44458# a_4093_43548# 2.85e-20
C21082 a_11813_46116# VDD 0.434656f
C21083 a_453_43940# a_2479_44172# 0.003275f
C21084 a_18479_47436# a_20835_44721# 0.007754f
C21085 a_16327_47482# a_18753_44484# 7.32e-19
C21086 a_n1099_45572# a_1260_45572# 5.75e-20
C21087 a_12379_46436# a_11823_42460# 4.72e-19
C21088 a_8049_45260# a_8336_45822# 4e-19
C21089 a_768_44030# a_556_44484# 0.001175f
C21090 a_584_46384# a_5013_44260# 1.69e-19
C21091 a_n2293_46098# a_327_44734# 1.74e-19
C21092 a_n1076_46494# a_n967_45348# 4.41e-20
C21093 a_n443_46116# a_1115_44172# 6.13e-20
C21094 a_1823_45246# a_n2017_45002# 0.024027f
C21095 a_5066_45546# a_9159_45572# 0.040307f
C21096 a_18189_46348# a_16147_45260# 0.129202f
C21097 a_10809_44734# a_12561_45572# 1.38e-19
C21098 a_4185_45028# a_22959_45572# 3.35e-19
C21099 a_1138_42852# a_n1059_45260# 0.004009f
C21100 a_n356_45724# a_n443_42852# 0.056063f
C21101 a_n755_45592# a_509_45572# 1.66e-20
C21102 a_n357_42282# a_603_45572# 7.72e-19
C21103 a_18597_46090# a_20640_44752# 0.027095f
C21104 a_11453_44696# a_18204_44850# 1.39e-19
C21105 a_n784_42308# C5_P_btm 5.81e-19
C21106 a_1606_42308# a_11530_34132# 0.004863f
C21107 a_n815_47178# a_n1435_47204# 0.003452f
C21108 a_3160_47472# a_n443_46116# 0.018382f
C21109 a_3785_47178# a_4007_47204# 0.106797f
C21110 a_n1151_42308# a_4791_45118# 1.16458f
C21111 a_2063_45854# a_6151_47436# 0.448977f
C21112 a_2905_45572# a_4915_47217# 0.001556f
C21113 a_n1741_47186# a_13487_47204# 1.17e-19
C21114 a_n3420_39616# a_n3565_39304# 0.035199f
C21115 a_1239_39587# a_1736_39587# 0.105143f
C21116 a_n3690_39616# a_n3690_39392# 0.052468f
C21117 a_n3565_39590# a_n3420_39072# 0.033891f
C21118 a_22400_42852# VDD 0.829052f
C21119 a_n4064_39616# a_n4209_39304# 0.029393f
C21120 a_n4209_39590# a_n4064_39072# 0.03458f
C21121 en_comp a_15959_42545# 3.92e-20
C21122 a_n2661_42834# a_1847_42826# 6.72e-21
C21123 a_n2293_43922# a_685_42968# 8.95e-21
C21124 a_9313_44734# a_8037_42858# 5.36e-20
C21125 a_n356_44636# a_5534_30871# 0.054103f
C21126 a_11967_42832# a_13467_32519# 3.36e-21
C21127 a_18248_44752# a_18249_42858# 1.79e-20
C21128 a_18287_44626# a_17333_42852# 2.93e-20
C21129 a_5891_43370# a_10518_42984# 0.001688f
C21130 a_n2293_42834# a_n4318_37592# 0.003537f
C21131 a_3537_45260# a_5742_30871# 3.39e-20
C21132 a_14539_43914# a_19164_43230# 7.82e-21
C21133 a_20512_43084# a_15743_43084# 0.761578f
C21134 a_18579_44172# a_16823_43084# 1.17e-21
C21135 a_20835_44721# a_4190_30871# 1.12e-20
C21136 a_3499_42826# a_2813_43396# 2.45e-19
C21137 a_17737_43940# a_3626_43646# 5.73e-21
C21138 a_n1613_43370# a_n1809_43762# 0.012235f
C21139 a_n755_45592# a_2809_45348# 7.33e-20
C21140 a_6511_45714# a_6431_45366# 6.29e-19
C21141 a_6667_45809# a_6171_45002# 0.004899f
C21142 a_n443_42852# a_14537_43396# 0.03432f
C21143 a_6472_45840# a_5205_44484# 2.12e-20
C21144 a_13259_45724# a_13105_45348# 1.66e-19
C21145 a_16680_45572# a_18341_45572# 6.97e-20
C21146 a_17478_45572# a_16147_45260# 0.050291f
C21147 a_8696_44636# a_18479_45785# 1.47e-20
C21148 a_15861_45028# a_18175_45572# 8.48e-20
C21149 a_2957_45546# a_1423_45028# 1.39e-20
C21150 a_13661_43548# a_19319_43548# 0.189089f
C21151 a_2324_44458# a_12607_44458# 4.05e-20
C21152 a_2711_45572# a_8953_45002# 0.003719f
C21153 a_8049_45260# a_18494_42460# 1.4e-19
C21154 a_n2312_39304# a_n1557_42282# 1.92e-20
C21155 a_n4064_37440# C4_P_btm 1.74e-19
C21156 a_n3565_37414# C0_P_btm 0.040442f
C21157 a_n3420_37440# C2_P_btm 2.75e-19
C21158 a_n881_46662# a_2609_46660# 1.09e-19
C21159 a_n1613_43370# a_3177_46902# 0.209276f
C21160 a_4915_47217# a_12816_46660# 0.006808f
C21161 a_22821_38993# a_22609_38406# 8.2e-19
C21162 a_22469_39537# CAL_P 0.024901f
C21163 a_22521_39511# a_22609_37990# 0.333805f
C21164 a_22459_39145# a_22717_37285# 0.012249f
C21165 a_768_44030# a_2107_46812# 0.087742f
C21166 VDAC_N EN_VIN_BSTR_N 0.341021f
C21167 a_15673_47210# a_6755_46942# 1.86e-19
C21168 a_10227_46804# a_9863_46634# 0.278164f
C21169 a_n967_45348# VDD 0.556063f
C21170 en_comp RST_Z 4.34313f
C21171 a_10341_43396# a_15781_43660# 0.011941f
C21172 a_n809_44244# a_n473_42460# 1.26e-20
C21173 a_n984_44318# a_n961_42308# 1.84e-20
C21174 a_19963_31679# VCM 0.035453f
C21175 a_13565_43940# a_12379_42858# 1.27e-20
C21176 a_1568_43370# a_n13_43084# 1.85e-20
C21177 a_20447_31679# VREF 0.059621f
C21178 a_n1761_44111# a_n3674_37592# 0.002395f
C21179 a_n97_42460# a_685_42968# 0.034735f
C21180 a_14021_43940# a_22959_42860# 3.35e-19
C21181 a_14579_43548# a_16547_43609# 5.47e-21
C21182 a_6197_43396# a_743_42282# 3.82e-20
C21183 a_12549_44172# a_21356_42826# 2.29e-20
C21184 a_n1151_42308# a_n1736_42282# 1.63e-20
C21185 a_15595_45028# a_16019_45002# 0.017418f
C21186 a_15415_45028# a_1307_43914# 1.07e-19
C21187 a_15599_45572# a_16112_44458# 7.05e-19
C21188 a_8696_44636# a_10057_43914# 0.001707f
C21189 a_8746_45002# a_10617_44484# 0.01623f
C21190 a_21513_45002# a_21101_45002# 0.003301f
C21191 a_10227_46804# a_11136_42852# 0.012196f
C21192 a_12861_44030# a_15597_42852# 5.41e-19
C21193 a_8016_46348# a_10555_43940# 3.45e-19
C21194 a_5937_45572# a_9165_43940# 1.38e-20
C21195 a_5111_44636# a_5837_45028# 0.019542f
C21196 a_7499_43078# a_n2293_43922# 1.48e-19
C21197 a_4927_45028# a_5093_45028# 0.143754f
C21198 a_9049_44484# a_n2661_43922# 0.003185f
C21199 a_n37_45144# a_n2661_43370# 0.007073f
C21200 a_9482_43914# a_1423_45028# 0.014596f
C21201 a_2711_45572# a_16335_44484# 0.001233f
C21202 a_3537_45260# a_n2293_42834# 0.195818f
C21203 a_15227_44166# a_10341_43396# 0.068268f
C21204 a_12549_44172# a_14275_46494# 4.53e-20
C21205 a_n971_45724# a_n863_45724# 0.199707f
C21206 a_1123_46634# a_1823_45246# 1.41e-19
C21207 a_4883_46098# a_n1925_42282# 5.4e-19
C21208 a_n2109_47186# a_997_45618# 4.13e-22
C21209 a_5807_45002# a_9290_44172# 0.00233f
C21210 a_n743_46660# a_3483_46348# 0.050648f
C21211 a_n2661_46098# a_n1991_46122# 0.025798f
C21212 a_948_46660# a_1138_42852# 4.64e-20
C21213 a_2107_46812# a_1176_45822# 1.38e-19
C21214 a_327_47204# a_n2661_45546# 5.19e-21
C21215 a_15009_46634# a_15559_46634# 4.99e-19
C21216 a_3090_45724# a_15368_46634# 0.440843f
C21217 a_6755_46942# a_16388_46812# 0.002525f
C21218 a_n1925_46634# a_4185_45028# 2.83e-19
C21219 a_n746_45260# a_n1079_45724# 9.3e-19
C21220 a_n237_47217# a_n2293_45546# 0.002405f
C21221 a_n2661_46634# a_5497_46414# 2.47e-20
C21222 a_n2497_47436# a_2957_45546# 2.23e-21
C21223 a_1847_42826# a_n2293_42282# 4.45e-19
C21224 a_15743_43084# a_16245_42852# 4.92e-19
C21225 a_n97_42460# a_14113_42308# 0.356407f
C21226 a_12379_42858# a_5534_30871# 0.128429f
C21227 a_12545_42858# a_13460_43230# 0.118423f
C21228 a_6293_42852# a_6171_42473# 0.00101f
C21229 a_6031_43396# a_5932_42308# 3.68e-19
C21230 a_9159_44484# VDD 0.004886f
C21231 a_3539_42460# a_5934_30871# 1.41e-20
C21232 a_3626_43646# a_8515_42308# 0.003306f
C21233 a_413_45260# a_2889_44172# 0.127135f
C21234 a_n2017_45002# a_n3674_39768# 2.64e-19
C21235 a_n1925_42282# a_5649_42852# 0.001675f
C21236 a_9290_44172# a_10518_42984# 0.04331f
C21237 a_4185_45028# a_16795_42852# 4.48e-21
C21238 a_7499_43078# a_n97_42460# 0.212833f
C21239 a_5343_44458# a_5518_44484# 0.054464f
C21240 a_n443_42852# a_6547_43396# 0.006641f
C21241 a_n2293_45010# a_n1453_44318# 0.001505f
C21242 a_19431_45546# a_15493_43396# 1.48e-19
C21243 a_8953_45546# a_10341_42308# 0.006033f
C21244 a_2711_45572# a_3626_43646# 0.072582f
C21245 a_3065_45002# a_1414_42308# 4.93e-19
C21246 a_13259_45724# a_13749_43396# 0.002234f
C21247 a_8696_44636# a_14021_43940# 2.1e-19
C21248 a_2324_44458# a_3681_42891# 9.45e-22
C21249 a_18597_46090# a_21188_45572# 0.00956f
C21250 a_n743_46660# a_14495_45572# 6.59e-20
C21251 a_17609_46634# a_16375_45002# 2.49e-19
C21252 a_3160_47472# a_3537_45260# 1.25e-21
C21253 a_n443_46116# a_413_45260# 0.369976f
C21254 a_18479_47436# a_20731_45938# 0.007339f
C21255 a_15811_47375# a_3357_43084# 2.81e-19
C21256 a_16327_47482# a_2437_43646# 0.046662f
C21257 a_4646_46812# a_7227_45028# 0.305597f
C21258 a_3877_44458# a_3775_45552# 0.002726f
C21259 a_20820_30879# a_10809_44734# 0.234047f
C21260 a_3483_46348# a_11189_46129# 0.001012f
C21261 a_6419_46155# a_8016_46348# 1.19e-20
C21262 a_12741_44636# a_22223_46124# 1.14e-19
C21263 a_5204_45822# a_5937_45572# 2.47e-19
C21264 a_n971_45724# a_8191_45002# 0.015833f
C21265 a_12549_44172# a_15765_45572# 3.88e-21
C21266 a_2063_45854# a_5111_44636# 0.004291f
C21267 a_20894_47436# a_20841_45814# 3.24e-21
C21268 a_3080_42308# C5_P_btm 3.03e-19
C21269 a_n2472_42282# a_n2104_42282# 7.52e-19
C21270 a_n1917_43396# VDD 0.204644f
C21271 a_16414_43172# a_4958_30871# 8.46e-19
C21272 a_n3674_38680# a_n3674_38216# 0.059687f
C21273 a_9061_43230# a_5934_30871# 5.05e-21
C21274 a_17767_44458# a_17737_43940# 0.004352f
C21275 a_n2661_43922# a_3905_42865# 3.56e-19
C21276 a_n2661_42834# a_5244_44056# 0.00436f
C21277 a_11967_42832# a_22315_44484# 6.72e-19
C21278 a_526_44458# a_5934_30871# 3.53e-19
C21279 a_n443_42852# a_12991_43230# 1.9e-19
C21280 a_16922_45042# a_21381_43940# 0.003996f
C21281 a_20692_30879# a_14097_32519# 0.051423f
C21282 a_4185_45028# a_21335_42336# 8e-20
C21283 a_19279_43940# a_18579_44172# 0.372064f
C21284 a_n2293_42834# a_1049_43396# 0.001716f
C21285 a_1307_43914# a_7112_43396# 3.85e-21
C21286 a_1110_47026# VDD 4.6e-19
C21287 a_n357_42282# a_14853_42852# 5.87e-19
C21288 a_n1059_45260# a_17499_43370# 0.385066f
C21289 a_n2017_45002# a_17324_43396# 1.13e-19
C21290 a_n913_45002# a_16759_43396# 3.29e-21
C21291 a_11453_44696# a_15004_44636# 3.53e-21
C21292 a_2324_44458# a_8746_45002# 0.34917f
C21293 a_15682_46116# a_10193_42453# 7.91e-19
C21294 a_5937_45572# a_8697_45822# 0.019555f
C21295 a_16375_45002# a_19443_46116# 4.21e-20
C21296 a_8199_44636# a_9241_45822# 1.53e-20
C21297 a_8016_46348# a_10907_45822# 1.99e-20
C21298 a_768_44030# a_n2661_44458# 0.028401f
C21299 a_4883_46098# a_18248_44752# 1.47e-21
C21300 a_10903_43370# a_13527_45546# 0.035694f
C21301 a_12594_46348# a_12791_45546# 0.026771f
C21302 a_13351_46090# a_11823_42460# 1.2e-19
C21303 a_6755_46942# a_13777_45326# 1.05e-21
C21304 a_3483_46348# a_11136_45572# 0.020129f
C21305 a_n881_46662# a_2779_44458# 3.56e-21
C21306 a_13059_46348# a_3357_43084# 1.83e-20
C21307 a_3090_45724# a_2680_45002# 0.003269f
C21308 a_n1613_43370# a_4223_44672# 0.022154f
C21309 a_20273_46660# a_20273_45572# 4.74e-19
C21310 a_20107_46660# a_20623_45572# 2.63e-20
C21311 a_2443_46660# a_n2661_43370# 1.76e-21
C21312 a_5934_30871# a_n4209_38502# 6.81e-22
C21313 a_22223_42860# VDD 0.250812f
C21314 a_18907_42674# a_19511_42282# 0.001351f
C21315 a_22165_42308# RST_Z 4.44e-21
C21316 a_17303_42282# a_20712_42282# 3.71e-19
C21317 a_4958_30871# a_7174_31319# 0.107892f
C21318 a_1606_42308# a_7754_40130# 0.001975f
C21319 a_6123_31319# a_n3565_38502# 3.8e-21
C21320 a_5742_30871# a_1343_38525# 1.5e-19
C21321 a_n356_44636# a_4190_30871# 0.04771f
C21322 a_20365_43914# a_14021_43940# 0.003393f
C21323 a_n1059_45260# a_1576_42282# 0.003521f
C21324 a_n2017_45002# a_1184_42692# 0.040166f
C21325 a_1115_44172# a_1049_43396# 3.25e-19
C21326 a_1467_44172# a_1209_43370# 0.004302f
C21327 a_9313_44734# a_18525_43370# 8.26e-20
C21328 a_742_44458# a_685_42968# 9.87e-20
C21329 a_14673_44172# a_14579_43548# 2.2e-20
C21330 a_n2956_37592# a_n3674_37592# 0.025613f
C21331 a_n913_45002# a_1067_42314# 9.28e-20
C21332 a_15682_46116# VDD 1.25004f
C21333 a_2324_44458# RST_Z 1.22e-21
C21334 a_n4318_39768# a_n2840_43370# 7.62e-19
C21335 a_3600_43914# a_n97_42460# 3.85e-21
C21336 a_n967_45348# a_n784_42308# 0.007598f
C21337 a_14537_43396# a_14635_42282# 4.55e-19
C21338 a_n2293_42834# a_4649_43172# 2.27e-19
C21339 a_584_46384# a_4699_43561# 7.44e-19
C21340 a_12861_44030# a_21205_44306# 3.21e-19
C21341 a_n1641_46494# a_n1352_44484# 2.48e-20
C21342 a_n2293_46098# a_4223_44672# 0.422068f
C21343 a_10193_42453# a_16680_45572# 1.46e-20
C21344 a_10180_45724# a_8696_44636# 0.002551f
C21345 a_n863_45724# a_n2293_45010# 0.090522f
C21346 a_13759_46122# a_14309_45028# 1.57e-20
C21347 a_2324_44458# a_14403_45348# 0.0023f
C21348 a_n2661_45546# a_n745_45366# 0.00237f
C21349 a_n2810_45572# a_n2810_45028# 0.063288f
C21350 a_12549_44172# a_19328_44172# 0.012953f
C21351 a_n2293_45546# a_n2017_45002# 1.75e-19
C21352 a_3090_45724# a_15146_44811# 1.56e-19
C21353 a_380_45546# a_n2661_45010# 3.48e-21
C21354 a_1176_45822# a_n2661_44458# 8.11e-22
C21355 a_8697_45822# a_8697_45572# 6.96e-20
C21356 a_8049_45260# a_13777_45326# 4.46e-20
C21357 a_18479_47436# a_20843_47204# 0.021416f
C21358 a_18780_47178# a_19594_46812# 2.12e-19
C21359 a_n1435_47204# a_171_46873# 5.97e-20
C21360 a_9067_47204# a_2107_46812# 1.22e-20
C21361 VDAC_Pi a_5700_37509# 2.20213f
C21362 a_3754_38470# a_7754_38470# 3.02e-20
C21363 a_11453_44696# a_768_44030# 0.031665f
C21364 a_7174_31319# VCM 0.076834f
C21365 a_10227_46804# a_20916_46384# 0.013668f
C21366 a_19787_47423# a_13747_46662# 1.81e-19
C21367 a_7754_40130# a_8912_37509# 1.81084f
C21368 a_n443_46116# a_2609_46660# 0.349838f
C21369 a_3815_47204# a_3524_46660# 1.6e-20
C21370 a_4007_47204# a_3699_46634# 0.008067f
C21371 a_584_46384# a_3877_44458# 1.42e-20
C21372 a_n4209_39590# VDD 2.06918f
C21373 a_7754_39964# a_6886_37412# 0.035115f
C21374 a_n3565_39304# C2_P_btm 1.93e-20
C21375 a_n4064_39072# C6_P_btm 2.76e-20
C21376 a_18597_46090# a_19321_45002# 0.024487f
C21377 a_19386_47436# a_19452_47524# 0.006978f
C21378 a_13487_47204# a_n743_46660# 2.02e-20
C21379 a_n971_45724# a_5072_46660# 4.58e-21
C21380 a_n2109_47186# a_5257_43370# 0.153164f
C21381 a_n3565_38502# EN_VIN_BSTR_P 0.003421f
C21382 a_20447_31679# a_22521_40599# 2.27e-20
C21383 a_10729_43914# a_10796_42968# 7.16e-21
C21384 a_10949_43914# a_10835_43094# 4.11e-21
C21385 a_10807_43548# a_10518_42984# 7.97e-19
C21386 a_n2293_43922# a_n1329_42308# 4.07e-19
C21387 a_n97_42460# a_15781_43660# 0.001962f
C21388 a_16680_45572# VDD 0.275078f
C21389 a_8147_43396# a_8791_43396# 0.001846f
C21390 a_6547_43396# a_6655_43762# 0.057222f
C21391 a_n2956_37592# a_n2216_37690# 0.001674f
C21392 a_18494_42460# a_13258_32519# 0.298557f
C21393 a_18184_42460# a_20107_42308# 0.013525f
C21394 a_11967_42832# a_18695_43230# 0.001256f
C21395 a_21381_43940# a_15743_43084# 0.02274f
C21396 a_13747_46662# a_21487_43396# 0.009398f
C21397 a_13661_43548# a_19095_43396# 0.048302f
C21398 a_15227_44166# a_n97_42460# 0.044664f
C21399 a_8049_45260# a_20640_44752# 2.15e-21
C21400 a_413_45260# a_3537_45260# 3.32e-19
C21401 a_19321_45002# a_743_42282# 1.16e-19
C21402 a_12861_44030# a_18083_42858# 2.04e-22
C21403 a_n1613_43370# a_n3674_39304# 2.21e-20
C21404 a_5257_43370# a_5837_43396# 1.77e-21
C21405 a_n443_42852# a_n356_44636# 0.262144f
C21406 a_n755_45592# a_5891_43370# 0.062112f
C21407 a_2324_44458# a_5663_43940# 0.010841f
C21408 a_3483_46348# a_11750_44172# 2.37e-21
C21409 a_10227_46804# a_12545_42858# 0.03565f
C21410 a_2274_45254# a_2680_45002# 0.076507f
C21411 a_12549_44172# a_20749_43396# 0.018798f
C21412 a_10150_46912# a_10428_46928# 0.118759f
C21413 a_9863_46634# a_10467_46802# 0.043587f
C21414 a_8145_46902# a_6755_46942# 0.02566f
C21415 a_7577_46660# a_6969_46634# 6.14e-19
C21416 a_5257_43370# a_5841_46660# 5.15e-20
C21417 a_n1435_47204# a_10903_43370# 1.64e-20
C21418 a_n1151_42308# a_6945_45028# 0.024325f
C21419 a_19321_45002# a_19123_46287# 2.27e-20
C21420 a_13747_46662# a_20107_46660# 2.33e-21
C21421 a_13661_43548# a_20411_46873# 3e-19
C21422 a_n2293_46634# a_13059_46348# 0.207934f
C21423 a_12549_44172# a_18280_46660# 0.03199f
C21424 a_16750_47204# a_765_45546# 1.34e-19
C21425 a_n743_46660# a_14513_46634# 2.15e-20
C21426 a_n1809_43762# a_n1736_42282# 1.55e-20
C21427 a_3422_30871# a_n4064_38528# 0.031148f
C21428 a_5649_42852# a_8387_43230# 1.14e-20
C21429 a_n901_43156# a_685_42968# 1.06e-20
C21430 a_n13_43084# a_133_43172# 0.013377f
C21431 a_n3674_39304# a_n1533_42852# 8.15e-22
C21432 a_n2433_43396# a_n1630_35242# 2.03e-20
C21433 a_4361_42308# a_10083_42826# 1.21e-19
C21434 a_18525_43370# a_18599_43230# 4.07e-19
C21435 a_15743_43084# a_18249_42858# 0.002881f
C21436 a_18783_43370# a_18817_42826# 0.012757f
C21437 a_743_42282# a_10922_42852# 1.14e-20
C21438 a_n1917_44484# VDD 0.186988f
C21439 a_15682_43940# a_16104_42674# 1.03e-20
C21440 a_n4318_39768# a_n4315_30879# 0.002449f
C21441 a_n2267_43396# a_n3674_37592# 1.26e-20
C21442 a_8685_43396# a_9306_43218# 1.84e-19
C21443 a_n2661_43370# a_949_44458# 6.02e-19
C21444 a_16922_45042# a_19929_45028# 0.003656f
C21445 a_5111_44636# a_n2661_42834# 0.04935f
C21446 a_5147_45002# a_n2661_43922# 0.029995f
C21447 a_13904_45546# a_13483_43940# 2.98e-21
C21448 a_13249_42308# a_12429_44172# 5.54e-19
C21449 a_10193_42453# a_20269_44172# 3.41e-21
C21450 a_3232_43370# a_10617_44484# 0.020516f
C21451 a_18494_42460# a_20193_45348# 0.116597f
C21452 a_16327_47482# a_19511_42282# 0.089559f
C21453 a_17719_45144# a_17969_45144# 0.008267f
C21454 a_375_42282# a_n356_44636# 0.015238f
C21455 SMPL_ON_P a_n3565_38502# 8.06e-19
C21456 a_13059_46348# a_5342_30871# 1.53e-19
C21457 a_n743_46660# a_n357_42282# 0.03365f
C21458 a_n2293_46634# a_3218_45724# 0.001771f
C21459 a_768_44030# a_5907_45546# 1.57e-21
C21460 a_13885_46660# a_10903_43370# 5.54e-19
C21461 a_11453_44696# a_11652_45724# 0.01055f
C21462 a_n1925_46634# a_997_45618# 5.01e-21
C21463 a_n2438_43548# a_310_45028# 2.28e-20
C21464 a_n1021_46688# a_n755_45592# 1.15e-20
C21465 a_n133_46660# a_n1099_45572# 5.35e-21
C21466 a_8145_46902# a_8049_45260# 4.44e-19
C21467 a_15227_44166# a_17957_46116# 0.0045f
C21468 a_18834_46812# a_18819_46122# 3.09e-19
C21469 a_12465_44636# a_12791_45546# 5.57e-21
C21470 a_4883_46098# a_13527_45546# 9.93e-20
C21471 a_10227_46804# a_10210_45822# 0.006028f
C21472 a_13507_46334# a_13249_42308# 2.05e-20
C21473 a_12816_46660# a_10809_44734# 0.011603f
C21474 a_14084_46812# a_6945_45028# 5.12e-21
C21475 a_6755_46942# a_5066_45546# 1.35e-19
C21476 a_1123_46634# a_n2293_45546# 1.17e-21
C21477 a_19862_44208# RST_Z 4.49e-21
C21478 a_8605_42826# a_5934_30871# 6.8e-19
C21479 a_8037_42858# a_8515_42308# 6.68e-20
C21480 a_4361_42308# a_15761_42308# 1.23e-19
C21481 a_4190_30871# a_18727_42674# 0.035226f
C21482 a_n2293_42282# a_n473_42460# 2.57e-19
C21483 a_743_42282# a_17531_42308# 0.007539f
C21484 a_14401_32519# VDAC_N 2.6e-19
C21485 a_20269_44172# VDD 0.169009f
C21486 a_10903_43370# a_1606_42308# 1.35e-20
C21487 a_n2661_43370# a_11341_43940# 8.02e-20
C21488 a_n4318_40392# a_n4318_39768# 2.73673f
C21489 a_n2810_45028# a_n1557_42282# 9.47e-21
C21490 a_n89_47570# VDD 4.63e-19
C21491 a_4883_46098# EN_OFFSET_CAL 8.93e-21
C21492 a_1307_43914# a_9801_43940# 0.004166f
C21493 a_2779_44458# a_2889_44172# 0.005445f
C21494 a_3357_43084# a_6293_42852# 0.001183f
C21495 a_n443_42852# a_12379_42858# 2.06e-19
C21496 a_n357_42282# a_17701_42308# 0.026888f
C21497 a_n2840_44458# a_n3674_39768# 0.005491f
C21498 a_n699_43396# a_895_43940# 0.001028f
C21499 a_n2661_43922# a_12553_44484# 0.009634f
C21500 a_1823_45246# a_4169_42308# 0.002692f
C21501 a_5066_45546# a_8049_45260# 0.076918f
C21502 a_n2293_46634# a_13556_45296# 0.00155f
C21503 a_2063_45854# a_10334_44484# 4.46e-36
C21504 a_4791_45118# a_4223_44672# 0.399086f
C21505 a_8667_46634# a_2437_43646# 1.27e-20
C21506 a_4883_46098# a_16922_45042# 4.62e-20
C21507 a_16327_47482# a_19113_45348# 1.22e-19
C21508 a_18985_46122# a_19443_46116# 0.027606f
C21509 a_n2497_47436# a_n1809_44850# 0.00201f
C21510 a_1823_45246# a_4099_45572# 0.047087f
C21511 a_167_45260# a_2711_45572# 0.003442f
C21512 a_2609_46660# a_3537_45260# 4.52e-20
C21513 a_n1151_42308# a_8103_44636# 2.41e-19
C21514 a_11453_44696# a_13490_45067# 4.23e-19
C21515 a_18597_46090# a_18184_42460# 0.020766f
C21516 a_18479_47436# a_20567_45036# 2.48e-20
C21517 a_n1613_43370# a_n2293_42834# 0.123758f
C21518 a_7577_46660# a_3357_43084# 1.08e-20
C21519 a_11415_45002# a_7499_43078# 4.24e-20
C21520 a_n443_46116# a_2779_44458# 0.00406f
C21521 a_3177_46902# a_3429_45260# 3.58e-20
C21522 a_2959_46660# a_3065_45002# 2.84e-20
C21523 a_n2661_46634# a_14537_43396# 7.41e-21
C21524 a_n1630_35242# a_n4064_40160# 1.13e-19
C21525 a_n3674_37592# a_n4251_40480# 9.61e-20
C21526 a_12563_42308# a_13070_42354# 0.001596f
C21527 a_n4318_37592# a_n4064_39616# 0.021014f
C21528 a_13467_32519# VREF 1.56e-19
C21529 a_17701_42308# CAL_N 8.77e-20
C21530 a_5932_42308# a_4958_30871# 0.01835f
C21531 a_n1853_43023# VDD 0.370563f
C21532 a_16922_45042# a_5649_42852# 8.28e-21
C21533 a_15004_44636# a_9145_43396# 3.39e-20
C21534 a_n2810_45572# a_n2302_40160# 7.76e-19
C21535 a_n1059_45260# a_4649_42852# 0.003629f
C21536 a_20820_30879# C6_N_btm 0.001067f
C21537 a_18184_42460# a_743_42282# 0.126294f
C21538 a_9482_43914# a_15567_42826# 1.86e-19
C21539 a_14537_43396# a_14543_43071# 9.84e-19
C21540 a_1307_43914# a_12545_42858# 4.9e-21
C21541 a_13556_45296# a_5342_30871# 1.19e-20
C21542 a_11967_42832# a_19319_43548# 5.45e-20
C21543 a_n2661_43922# a_4093_43548# 4.66e-20
C21544 a_6109_44484# a_6031_43396# 0.007586f
C21545 a_n2293_42834# a_n1533_42852# 0.003489f
C21546 a_18494_42460# a_20301_43646# 0.006153f
C21547 a_n2956_38216# a_n4315_30879# 0.025091f
C21548 a_n357_42282# a_21613_42308# 3.71e-20
C21549 a_7499_43078# a_10533_42308# 0.225871f
C21550 a_4419_46090# a_1423_45028# 3.66e-20
C21551 a_3090_45724# a_5518_44484# 9.17e-21
C21552 a_10903_43370# a_10775_45002# 3.83e-19
C21553 a_2711_45572# a_12791_45546# 0.008464f
C21554 a_2324_44458# a_3232_43370# 0.410727f
C21555 a_526_44458# a_n2661_45010# 0.703081f
C21556 a_13747_46662# a_21398_44850# 0.011329f
C21557 a_8049_45260# a_21188_45572# 0.015577f
C21558 a_4915_47217# a_11341_43940# 3.68e-20
C21559 a_12861_44030# a_12429_44172# 0.108591f
C21560 a_13259_45724# a_17786_45822# 0.001706f
C21561 a_n2109_47186# a_5807_45002# 0.003143f
C21562 a_2905_45572# a_n881_46662# 0.050468f
C21563 a_3160_47472# a_n1613_43370# 0.043254f
C21564 a_3785_47178# a_5063_47570# 2.94e-19
C21565 a_n1151_42308# a_3411_47243# 2.47e-19
C21566 a_n3565_39590# a_n2946_37690# 1.92e-19
C21567 a_n443_46116# a_3094_47570# 3.58e-19
C21568 a_16763_47508# a_17591_47464# 0.010417f
C21569 a_16023_47582# a_10227_46804# 0.036076f
C21570 a_16327_47482# a_18143_47464# 1.35e-19
C21571 a_5932_42308# VCM 0.146001f
C21572 a_n1435_47204# a_4883_46098# 2.09e-20
C21573 a_1736_39587# a_3754_38470# 0.002438f
C21574 a_n4209_39590# a_n2302_37690# 2.4e-19
C21575 a_5742_30871# C5_N_btm 0.089375f
C21576 a_13717_47436# a_21496_47436# 6.95e-20
C21577 a_12861_44030# a_13507_46334# 0.315418f
C21578 a_21613_42308# CAL_N 1.44e-19
C21579 a_n4064_40160# a_n3607_37440# 5.58e-20
C21580 a_9293_42558# VDD 0.006879f
C21581 a_n4064_39616# a_n4334_37440# 8.04e-19
C21582 a_n4209_38216# a_n4334_38304# 0.253307f
C21583 a_11341_43940# a_15681_43442# 1.37e-20
C21584 a_14539_43914# a_17749_42852# 0.002266f
C21585 a_n97_42460# a_1756_43548# 0.052563f
C21586 a_n2129_43609# a_n1557_42282# 9.91e-21
C21587 a_n2956_37592# a_n2302_39072# 0.005021f
C21588 a_6598_45938# VDD 0.204705f
C21589 a_4099_45572# DATA[2] 9.72e-21
C21590 a_15493_43396# a_16409_43396# 0.566182f
C21591 a_14021_43940# a_14205_43396# 0.008914f
C21592 a_11967_42832# a_16795_42852# 0.061673f
C21593 a_n356_44636# a_14635_42282# 1.57e-19
C21594 a_n2956_38216# a_n4318_40392# 0.027558f
C21595 a_20841_45814# a_19963_31679# 5.16e-20
C21596 a_768_44030# a_9145_43396# 0.004455f
C21597 a_19692_46634# a_20365_43914# 0.001873f
C21598 a_n2956_39304# a_n2661_43922# 1.05e-20
C21599 a_n2293_46634# a_6293_42852# 0.014742f
C21600 a_16115_45572# a_6171_45002# 3.23e-20
C21601 a_4185_45028# a_3422_30871# 0.176529f
C21602 a_16327_47482# a_21259_43561# 4.28e-20
C21603 a_584_46384# a_1847_42826# 4.79e-19
C21604 a_n1151_42308# a_n722_43218# 3.54e-19
C21605 a_12861_44030# a_21855_43396# 9.83e-19
C21606 a_21188_45572# a_19479_31679# 3.41e-20
C21607 a_21363_45546# a_3357_43084# 0.061421f
C21608 a_n2661_45546# a_n2433_44484# 3.06e-20
C21609 a_13507_46334# a_19700_43370# 4.92e-21
C21610 a_2711_45572# a_16405_45348# 5.81e-19
C21611 a_2324_44458# a_14581_44484# 1.05e-20
C21612 a_10809_44734# a_13213_44734# 1.94e-20
C21613 a_14840_46494# a_14673_44172# 2.17e-21
C21614 a_n1741_47186# a_3147_46376# 1.56e-20
C21615 a_n923_35174# VIN_P 1.547f
C21616 a_4883_46098# a_13885_46660# 5.17e-20
C21617 C6_P_btm VDD 0.210613f
C21618 a_5807_45002# a_5841_46660# 2.18e-20
C21619 a_n971_45724# a_2202_46116# 3.09e-20
C21620 a_3160_47472# a_n2293_46098# 1.31e-19
C21621 a_n881_46662# a_12816_46660# 5.76e-20
C21622 a_13507_46334# a_14180_46812# 3.77e-20
C21623 a_16327_47482# a_765_45546# 0.043622f
C21624 a_2107_46812# a_5167_46660# 0.002706f
C21625 a_2959_46660# a_3067_47026# 0.057222f
C21626 a_n1925_46634# a_5257_43370# 0.01497f
C21627 a_n2661_46634# a_8667_46634# 0.007776f
C21628 a_n237_47217# a_1138_42852# 2.57e-19
C21629 C3_P_btm C9_N_btm 0.001271f
C21630 C1_P_btm C7_N_btm 4.76e-19
C21631 C0_P_btm C6_N_btm 2.8e-19
C21632 a_11599_46634# a_20107_46660# 0.266678f
C21633 C0_dummy_P_btm C5_N_btm 1.24e-19
C21634 C0_N_btm C3_N_btm 0.409996f
C21635 C1_N_btm C2_N_btm 5.0586f
C21636 C0_dummy_N_btm C4_N_btm 0.113746f
C21637 a_13717_47436# a_21363_46634# 3.19e-20
C21638 a_2809_45028# VDD 0.189682f
C21639 a_16823_43084# a_17678_43396# 0.001907f
C21640 a_8685_43396# a_8387_43230# 0.002391f
C21641 a_3626_43646# a_18817_42826# 1.64e-20
C21642 a_2982_43646# a_19339_43156# 6.56e-21
C21643 a_4235_43370# a_n2293_42282# 7.36e-20
C21644 a_15743_43084# a_5649_42852# 0.024346f
C21645 a_2382_45260# a_5343_44458# 1e-19
C21646 a_n357_42282# a_11750_44172# 2.28e-21
C21647 a_5937_45572# a_6765_43638# 9.53e-19
C21648 a_2437_43646# a_n356_44636# 1.45e-20
C21649 a_15595_45028# a_11827_44484# 9.92e-21
C21650 a_6511_45714# a_6453_43914# 4.5e-21
C21651 a_3065_45002# a_n699_43396# 0.020711f
C21652 a_n2312_39304# a_n3674_37592# 0.026622f
C21653 a_13059_46348# a_743_42282# 2.35e-20
C21654 a_4791_45118# a_5742_30871# 3.2e-20
C21655 a_n913_45002# a_13720_44458# 3.43e-23
C21656 a_16333_45814# a_16241_44734# 1.85e-20
C21657 a_7276_45260# a_n2661_44458# 1.14e-20
C21658 a_19321_45002# a_8049_45260# 0.030309f
C21659 a_n2312_40392# a_n2810_45572# 0.052551f
C21660 a_n2312_39304# a_n2840_45546# 0.003056f
C21661 a_768_44030# a_14180_46482# 0.00983f
C21662 a_9863_46634# a_8016_46348# 0.001599f
C21663 a_8667_46634# a_8199_44636# 0.005444f
C21664 a_7227_47204# a_6511_45714# 7.86e-21
C21665 a_6491_46660# a_6598_45938# 1.3e-21
C21666 a_n443_46116# a_2211_45572# 1.46e-19
C21667 a_2063_45854# a_9049_44484# 3.38e-20
C21668 a_19692_46634# a_20885_46660# 0.002303f
C21669 a_n743_46660# a_518_46155# 4.76e-19
C21670 a_11459_47204# a_2711_45572# 3.52e-21
C21671 a_16721_46634# a_17829_46910# 8.81e-20
C21672 a_16388_46812# a_18285_46348# 0.028532f
C21673 a_15227_44166# a_11415_45002# 0.047556f
C21674 a_12281_43396# a_13575_42558# 5.62e-20
C21675 a_3422_30871# VREF_GND 0.10463f
C21676 a_n2472_42826# a_n3674_37592# 0.00166f
C21677 a_n1076_43230# COMP_P 1.14e-20
C21678 a_14955_43396# a_15051_42282# 2.17e-19
C21679 a_15095_43370# a_15486_42560# 0.001728f
C21680 a_3080_42308# a_n4209_39590# 7.41e-22
C21681 a_n1899_43946# VDD 0.475205f
C21682 a_n1853_43023# a_n784_42308# 8.46e-21
C21683 a_n4318_38680# a_n3674_38216# 0.023866f
C21684 a_12379_42858# a_14635_42282# 3.89e-21
C21685 a_12545_42858# a_13003_42852# 0.027606f
C21686 a_5534_30871# a_12800_43218# 1.43e-19
C21687 a_12089_42308# a_13291_42460# 1.22e-19
C21688 a_743_42282# a_2903_42308# 0.010301f
C21689 a_7499_43078# a_9885_43646# 2.67e-20
C21690 a_10193_42453# a_14358_43442# 2.71e-21
C21691 a_1307_43914# a_6101_44260# 7.06e-19
C21692 a_11827_44484# a_18005_44484# 3.81e-19
C21693 a_2711_45572# a_18525_43370# 7.09e-20
C21694 a_n2956_38680# a_n2293_42282# 3.4e-20
C21695 a_1431_47204# VDD 0.423871f
C21696 a_n971_45724# DATA[3] 0.09508f
C21697 a_10157_44484# a_n2661_43922# 0.00841f
C21698 a_10334_44484# a_n2661_42834# 5.65e-20
C21699 a_16979_44734# a_9313_44734# 1.28e-21
C21700 a_8975_43940# a_10617_44484# 0.025058f
C21701 a_11963_45334# a_11750_44172# 5.86e-21
C21702 a_9482_43914# a_10405_44172# 0.01085f
C21703 a_n357_42282# a_4361_42308# 0.069224f
C21704 a_9290_44172# a_10793_43218# 0.001055f
C21705 a_n2312_38680# a_n4064_38528# 0.22404f
C21706 a_n23_47502# DATA[0] 0.022435f
C21707 a_n237_47217# DATA[1] 0.139838f
C21708 a_n2293_42834# a_2675_43914# 1.48e-20
C21709 a_20193_45348# a_20640_44752# 0.017592f
C21710 a_626_44172# a_2537_44260# 4.41e-22
C21711 a_8953_45546# a_5066_45546# 0.191859f
C21712 a_10428_46928# a_10907_45822# 4.91e-20
C21713 a_10467_46802# a_10210_45822# 4.57e-20
C21714 a_4791_45118# a_n2293_42834# 0.046352f
C21715 a_768_44030# a_n1059_45260# 2.61e-19
C21716 a_12549_44172# a_n913_45002# 7.26e-19
C21717 a_n881_46662# a_n37_45144# 3.17e-19
C21718 a_n1613_43370# a_413_45260# 0.046335f
C21719 a_11735_46660# a_10193_42453# 0.001441f
C21720 a_12741_44636# a_20254_46482# 3.54e-19
C21721 a_19452_47524# a_3357_43084# 1.74e-19
C21722 a_4883_46098# a_10775_45002# 1.52e-21
C21723 a_16327_47482# a_16751_45260# 1.87e-19
C21724 a_20075_46420# a_20708_46348# 0.017547f
C21725 a_19553_46090# a_6945_45028# 1.78e-21
C21726 a_18819_46122# a_10809_44734# 7.49e-20
C21727 a_7920_46348# a_8062_46482# 0.007833f
C21728 a_765_45546# a_n356_45724# 3.13e-19
C21729 a_20843_47204# a_2437_43646# 0.004179f
C21730 a_10227_46804# a_14797_45144# 0.003451f
C21731 a_22365_46825# a_20205_31679# 0.002648f
C21732 a_1755_42282# a_6123_31319# 0.033073f
C21733 a_5267_42460# a_4921_42308# 0.04229f
C21734 a_1606_42308# a_7963_42308# 1.34e-20
C21735 a_14358_43442# VDD 0.170277f
C21736 a_13467_32519# a_22521_40599# 1.43e-20
C21737 a_4361_42308# CAL_N 0.003501f
C21738 a_6109_44484# a_6671_43940# 0.008633f
C21739 a_n699_43396# a_458_43396# 0.064001f
C21740 a_1467_44172# a_895_43940# 0.017277f
C21741 a_1414_42308# a_2479_44172# 0.110442f
C21742 a_11967_42832# a_10949_43914# 2.29e-20
C21743 a_n2661_43370# a_10341_43396# 2.26e-20
C21744 a_10193_42453# a_20836_43172# 0.009033f
C21745 a_18374_44850# a_18533_43940# 8.18e-21
C21746 a_18989_43940# a_19319_43548# 3.72e-20
C21747 a_n913_45002# a_5111_42852# 2.26e-19
C21748 a_n1059_45260# a_5755_42852# 0.005901f
C21749 a_n443_42852# a_3823_42558# 9.86e-21
C21750 a_n357_42282# a_6761_42308# 5.14e-21
C21751 a_13259_45724# a_14113_42308# 0.00391f
C21752 a_13490_45067# a_9145_43396# 5.1e-21
C21753 a_n2956_38680# a_n3565_39590# 0.021577f
C21754 a_453_43940# a_2127_44172# 0.007699f
C21755 a_11735_46660# VDD 0.407307f
C21756 a_742_44458# a_1756_43548# 0.152145f
C21757 a_949_44458# a_1568_43370# 6.56e-19
C21758 a_n1151_42308# a_895_43940# 6.25e-21
C21759 a_18479_47436# a_20679_44626# 0.018117f
C21760 a_16327_47482# a_18681_44484# 0.001931f
C21761 a_1848_45724# a_2307_45899# 6.64e-19
C21762 a_310_45028# a_603_45572# 8.28e-19
C21763 a_n1099_45572# a_1176_45572# 5.07e-20
C21764 a_n2497_47436# a_1525_44260# 4.47e-19
C21765 a_n2293_46098# a_413_45260# 0.034414f
C21766 a_5204_45822# a_2437_43646# 3.52e-20
C21767 a_n2661_45546# a_6194_45824# 4.12e-20
C21768 a_17715_44484# a_16147_45260# 0.020415f
C21769 a_n356_45724# a_509_45822# 2.78e-19
C21770 a_3218_45724# a_2277_45546# 7.5e-20
C21771 a_3316_45546# a_1609_45822# 1.08e-19
C21772 a_n357_42282# a_509_45572# 3.18e-19
C21773 a_18597_46090# a_20362_44736# 3.05e-20
C21774 a_11453_44696# a_17517_44484# 0.014468f
C21775 a_4185_45028# a_19963_31679# 9.16e-19
C21776 a_1138_42852# a_n2017_45002# 1.31e-19
C21777 a_n2946_39866# a_n4209_39304# 5.32e-20
C21778 a_n3420_39616# a_n4334_39392# 0.014828f
C21779 a_n4209_39590# a_n2946_39072# 5.32e-20
C21780 a_n784_42308# C6_P_btm 5.52e-19
C21781 a_n4064_40160# a_n3607_39392# 5.58e-20
C21782 a_n3565_39590# a_n3690_39392# 7.97e-20
C21783 a_n3690_39616# a_n3565_39304# 7.97e-20
C21784 a_5934_30871# VDAC_N 0.007165f
C21785 a_6123_31319# VDAC_P 0.00959f
C21786 a_n1605_47204# a_n1435_47204# 0.110832f
C21787 a_3785_47178# a_3815_47204# 0.270823f
C21788 a_2905_45572# a_n443_46116# 0.14923f
C21789 a_n1151_42308# a_4700_47436# 0.01362f
C21790 a_n1741_47186# a_12861_44030# 5.74e-20
C21791 a_n2293_42834# a_n1736_42282# 0.002516f
C21792 en_comp a_15803_42450# 8.24e-20
C21793 a_n2661_43922# a_685_42968# 1.03e-21
C21794 a_n2661_42834# a_791_42968# 1.41e-20
C21795 a_n356_44636# a_14543_43071# 1.16e-21
C21796 a_1307_43914# a_5379_42460# 2.61e-20
C21797 a_5111_44636# a_9885_42558# 3.55e-21
C21798 a_20159_44458# a_20556_43646# 7.51e-20
C21799 a_18287_44626# a_18083_42858# 4.69e-21
C21800 a_18248_44752# a_17333_42852# 4.89e-19
C21801 a_5891_43370# a_10083_42826# 0.016347f
C21802 a_20679_44626# a_4190_30871# 8.87e-19
C21803 a_20835_44721# a_21259_43561# 7.23e-22
C21804 a_20512_43084# a_18783_43370# 8.84e-20
C21805 a_n699_43396# a_2987_42968# 8.45e-20
C21806 a_15682_43940# a_3626_43646# 5.73e-21
C21807 a_2711_45572# a_8191_45002# 0.003439f
C21808 a_8049_45260# a_18184_42460# 6.28e-23
C21809 a_3483_46348# a_5891_43370# 0.005051f
C21810 a_n1613_43370# a_n2012_43396# 2.53e-19
C21811 a_n755_45592# a_2304_45348# 2.24e-19
C21812 a_2324_44458# a_8975_43940# 0.005091f
C21813 a_6945_45028# a_4223_44672# 1.31e-20
C21814 a_6511_45714# a_6171_45002# 0.012882f
C21815 a_6472_45840# a_6431_45366# 4.9e-19
C21816 a_8199_44636# a_n356_44636# 2.05e-19
C21817 a_6194_45824# a_5205_44484# 1.42e-21
C21818 a_10193_42453# en_comp 1.87e-19
C21819 a_16680_45572# a_18479_45785# 5.64e-19
C21820 a_15861_45028# a_16147_45260# 0.146279f
C21821 a_8696_44636# a_18175_45572# 3.95e-21
C21822 a_17478_45572# a_17786_45822# 0.017351f
C21823 a_16855_45546# a_18341_45572# 7.24e-20
C21824 a_4915_47217# a_10341_43396# 2.29e-20
C21825 a_1848_45724# a_1423_45028# 8.69e-22
C21826 a_5807_45002# a_19319_43548# 1.9e-20
C21827 a_n2312_40392# a_n1557_42282# 2.63e-20
C21828 a_n3420_37440# C3_P_btm 2.18e-19
C21829 a_n4064_37440# C5_P_btm 1.49e-19
C21830 a_n3565_37414# C1_P_btm 0.001047f
C21831 a_21588_30879# a_22612_30879# 7.53611f
C21832 a_n881_46662# a_2443_46660# 1.1e-19
C21833 a_n1151_42308# a_15559_46634# 2.09e-19
C21834 a_n1613_43370# a_2609_46660# 0.631348f
C21835 a_3754_39134# VDD 0.004567f
C21836 a_6151_47436# a_11901_46660# 2.66e-19
C21837 a_4915_47217# a_12991_46634# 0.068619f
C21838 a_3815_47204# a_3090_45724# 6.61e-21
C21839 a_5807_45002# a_n1925_46634# 0.933976f
C21840 VDAC_N a_11530_34132# 0.022899f
C21841 a_15811_47375# a_6755_46942# 8.93e-20
C21842 a_10227_46804# a_8492_46660# 6.27e-21
C21843 a_22469_39537# a_22876_39857# 2.68e-19
C21844 a_22521_39511# a_22705_38406# 0.004065f
C21845 VDAC_P EN_VIN_BSTR_P 0.339793f
C21846 a_22459_39145# a_22705_37990# 7.75e-19
C21847 a_22545_38993# a_22609_38406# 2.17e-21
C21848 en_comp VDD 4.26539f
C21849 a_10341_43396# a_15681_43442# 0.008134f
C21850 a_n809_44244# a_n961_42308# 2.8e-19
C21851 a_n1761_44111# a_n327_42558# 0.004022f
C21852 a_n356_44636# a_19511_42282# 5.6e-21
C21853 a_19963_31679# VREF_GND 0.001997f
C21854 a_8685_43396# a_15743_43084# 1.67e-19
C21855 a_6293_42852# a_743_42282# 1.73e-19
C21856 a_20447_31679# VIN_N 0.028787f
C21857 a_n97_42460# a_421_43172# 0.003376f
C21858 a_2711_45572# a_16241_44484# 0.001104f
C21859 a_13661_43548# a_16414_43172# 2.69e-21
C21860 a_12549_44172# a_20922_43172# 6.03e-19
C21861 a_n1151_42308# a_n3674_38216# 6.62e-20
C21862 a_14797_45144# a_1307_43914# 6.81e-21
C21863 a_14537_43396# a_16751_45260# 0.011362f
C21864 a_8696_44636# a_10440_44484# 0.00348f
C21865 a_21513_45002# a_21005_45260# 3.98e-19
C21866 a_3357_43084# a_19778_44110# 1.15e-19
C21867 a_10227_46804# a_13157_43218# 0.001903f
C21868 a_8016_46348# a_9801_43940# 4.95e-19
C21869 a_11823_42460# a_9313_44734# 0.0934f
C21870 a_5111_44636# a_5093_45028# 0.021262f
C21871 a_7499_43078# a_n2661_43922# 0.087751f
C21872 a_4927_45028# a_5009_45028# 0.096132f
C21873 a_5147_45002# a_5837_45028# 0.001063f
C21874 a_n143_45144# a_n2661_43370# 0.002979f
C21875 a_n1613_43370# a_n914_42852# 1.3e-19
C21876 a_10809_44734# a_11341_43940# 1.55e-19
C21877 a_n2293_46634# a_10991_42826# 4.93e-20
C21878 a_768_44030# a_13925_46122# 0.02161f
C21879 a_12891_46348# a_14275_46494# 4.45e-21
C21880 a_8667_46634# a_765_45546# 1.37e-20
C21881 a_4883_46098# a_526_44458# 0.010154f
C21882 a_n2109_47186# a_n755_45592# 5.59e-21
C21883 a_5807_45002# a_10355_46116# 0.003081f
C21884 a_n743_46660# a_3147_46376# 0.016933f
C21885 a_n2661_46098# a_n1853_46287# 0.019613f
C21886 a_1123_46634# a_1138_42852# 0.00173f
C21887 a_2609_46660# a_n2293_46098# 1.8e-20
C21888 a_948_46660# a_1176_45822# 0.003207f
C21889 a_2107_46812# a_1208_46090# 5e-19
C21890 a_15009_46634# a_15368_46634# 7.72e-19
C21891 a_12861_44030# a_10586_45546# 9.62e-21
C21892 a_6755_46942# a_13059_46348# 0.239671f
C21893 a_3090_45724# a_14976_45028# 0.730613f
C21894 a_n746_45260# a_n2293_45546# 0.404324f
C21895 a_n971_45724# a_n1079_45724# 0.150623f
C21896 a_n2661_46634# a_5204_45822# 1.9e-19
C21897 a_33_46660# a_167_45260# 7.22e-22
C21898 a_n2497_47436# a_1848_45724# 7.52e-22
C21899 a_2813_43396# a_2903_42308# 6.21e-21
C21900 a_15743_43084# a_15953_42852# 0.006469f
C21901 a_n97_42460# a_13657_42558# 0.011259f
C21902 a_13113_42826# a_12895_43230# 0.209641f
C21903 a_12379_42858# a_14543_43071# 5.72e-21
C21904 a_12545_42858# a_13635_43156# 0.041762f
C21905 a_2982_43646# a_3905_42308# 4.18e-19
C21906 a_6031_43396# a_6171_42473# 2.49e-21
C21907 a_10617_44484# VDD 0.141193f
C21908 a_3626_43646# a_5934_30871# 0.192998f
C21909 a_n2661_43370# a_n2293_43922# 0.001105f
C21910 a_413_45260# a_2675_43914# 0.048283f
C21911 a_327_44734# a_895_43940# 3.3e-19
C21912 a_n2293_45010# a_n1644_44306# 3.56e-19
C21913 a_n2017_45002# a_n4318_39768# 9.4e-20
C21914 a_526_44458# a_5649_42852# 0.058712f
C21915 a_9290_44172# a_10083_42826# 0.136441f
C21916 a_4743_44484# a_5518_44484# 1.16e-19
C21917 a_4223_44672# a_8103_44636# 1.47e-19
C21918 a_n443_42852# a_6765_43638# 0.00334f
C21919 a_2274_45254# a_2127_44172# 5.57e-20
C21920 a_n2312_39304# a_n2302_39072# 0.130454f
C21921 a_n913_45002# a_7542_44172# 9.32e-22
C21922 a_13661_43548# a_7174_31319# 1.16e-20
C21923 a_2680_45002# a_1414_42308# 6.45e-20
C21924 a_2324_44458# a_2905_42968# 8.09e-22
C21925 a_18597_46090# a_21363_45546# 0.001567f
C21926 a_n743_46660# a_13249_42308# 4.93e-20
C21927 a_13059_46348# a_8049_45260# 0.068978f
C21928 a_n443_46116# a_n37_45144# 3.75e-19
C21929 a_4791_45118# a_413_45260# 2.6e-19
C21930 a_n881_46662# a_16223_45938# 8.49e-19
C21931 a_16241_47178# a_2437_43646# 0.004738f
C21932 a_16327_47482# a_21513_45002# 0.013118f
C21933 a_4646_46812# a_6598_45938# 6.19e-19
C21934 a_3483_46348# a_9290_44172# 0.207611f
C21935 a_12741_44636# a_6945_45028# 0.021699f
C21936 a_5164_46348# a_5937_45572# 3.66e-19
C21937 a_n237_47217# a_7229_43940# 4.29e-19
C21938 a_n971_45724# a_7705_45326# 5.33e-21
C21939 a_12549_44172# a_15903_45785# 3.38e-20
C21940 a_15227_44166# a_13259_45724# 0.916975f
C21941 a_3160_47472# a_3429_45260# 3.37e-21
C21942 a_2063_45854# a_5147_45002# 1.79e-19
C21943 a_11415_45002# a_22959_46124# 0.002009f
C21944 a_22591_46660# a_10809_44734# 0.013929f
C21945 a_15507_47210# a_3357_43084# 4.74e-19
C21946 a_20894_47436# a_20273_45572# 1.81e-21
C21947 a_3080_42308# C6_P_btm 2.67e-19
C21948 a_n2472_42282# a_n4318_38216# 0.157105f
C21949 a_n1699_43638# VDD 0.210236f
C21950 a_n2840_42282# a_n3674_38216# 0.03703f
C21951 a_15567_42826# a_4958_30871# 7.19e-21
C21952 a_1307_43914# a_7287_43370# 1.2e-19
C21953 a_n2661_42834# a_3905_42865# 0.018962f
C21954 a_17517_44484# a_19237_31679# 0.00388f
C21955 a_11967_42832# a_3422_30871# 0.139082f
C21956 a_10193_42453# a_22165_42308# 2.46e-21
C21957 a_n2661_43922# a_3600_43914# 8.69e-19
C21958 en_comp a_16137_43396# 1.88e-20
C21959 a_526_44458# a_7963_42308# 5.22e-20
C21960 a_n1925_42282# a_6123_31319# 3.21e-20
C21961 a_20692_30879# a_22400_42852# 8.51e-20
C21962 a_20205_31679# a_14097_32519# 0.051224f
C21963 a_1123_46634# DATA[1] 0.00365f
C21964 a_4185_45028# a_7174_31319# 0.027406f
C21965 a_n2661_43370# a_n97_42460# 6.42e-21
C21966 a_20640_44752# a_20596_44850# 1.46e-19
C21967 a_n935_46688# VDD 2.29e-19
C21968 a_n2293_42834# a_1209_43370# 0.001969f
C21969 a_n357_42282# a_13622_42852# 1.14e-19
C21970 a_n2017_45002# a_17499_43370# 4.8e-19
C21971 a_n1059_45260# a_16759_43396# 1.17e-19
C21972 a_n913_45002# a_16977_43638# 1.48e-21
C21973 a_16721_46634# a_2437_43646# 1.5e-22
C21974 a_11453_44696# a_13720_44458# 1.26e-20
C21975 a_2324_44458# a_10193_42453# 0.041338f
C21976 a_n2661_46098# a_n2661_43370# 1.87e-20
C21977 a_8199_44636# a_8697_45822# 0.067739f
C21978 a_8016_46348# a_10210_45822# 0.003734f
C21979 a_12549_44172# a_n2661_44458# 4.11e-20
C21980 a_16292_46812# a_413_45260# 1.24e-20
C21981 a_10903_43370# a_13163_45724# 0.06577f
C21982 a_12594_46348# a_11823_42460# 0.081079f
C21983 a_6755_46942# a_13556_45296# 0.103107f
C21984 a_19321_45002# a_20193_45348# 0.489018f
C21985 a_19594_46812# a_11691_44458# 1.96e-19
C21986 a_3483_46348# a_11064_45572# 0.002687f
C21987 a_n881_46662# a_949_44458# 1.39e-19
C21988 a_9313_45822# a_9313_44734# 1.19e-20
C21989 a_3090_45724# a_2382_45260# 0.002468f
C21990 a_11415_45002# a_16377_45572# 4.28e-19
C21991 a_20273_46660# a_20107_45572# 8.09e-19
C21992 a_20411_46873# a_20273_45572# 6.47e-19
C21993 a_20107_46660# a_20841_45814# 1.73e-21
C21994 a_8270_45546# a_7229_43940# 1.4e-36
C21995 a_13661_43548# a_16981_45144# 2.68e-21
C21996 a_17303_42282# a_20107_42308# 3.68e-19
C21997 a_22165_42308# VDD 0.336187f
C21998 a_18727_42674# a_19511_42282# 5.06e-19
C21999 a_21671_42860# RST_Z 4.49e-21
C22000 a_2998_44172# a_n97_42460# 4.27e-19
C22001 a_11133_46155# CLK 0.001561f
C22002 a_20269_44172# a_14021_43940# 5.52e-20
C22003 a_n2293_45010# a_961_42354# 2.42e-20
C22004 a_n2017_45002# a_1576_42282# 0.008099f
C22005 a_8333_44056# a_8487_44056# 0.008678f
C22006 a_1115_44172# a_1209_43370# 1.17e-19
C22007 a_18989_43940# a_19095_43396# 2.42e-19
C22008 a_9313_44734# a_18429_43548# 3.66e-20
C22009 a_n1059_45260# a_1067_42314# 0.006623f
C22010 a_n913_45002# a_n1630_35242# 3.81e-19
C22011 a_2324_44458# VDD 2.73366f
C22012 a_n2810_45028# a_n3674_37592# 0.025732f
C22013 en_comp a_n784_42308# 0.025103f
C22014 a_n967_45348# a_196_42282# 3.02e-20
C22015 a_14537_43396# a_13291_42460# 2.95e-20
C22016 a_n2293_42834# a_3059_42968# 1.04e-19
C22017 a_14840_46494# RST_Z 2.03e-21
C22018 a_526_44458# a_3602_45348# 7.3e-19
C22019 a_584_46384# a_4235_43370# 0.016368f
C22020 a_n971_45724# a_2982_43646# 3.56e-20
C22021 a_n2497_47436# a_1512_43396# 9.13e-21
C22022 a_n1641_46494# a_n1177_44458# 4.88e-19
C22023 a_10193_42453# a_16855_45546# 3.49e-20
C22024 a_n452_45724# a_n2661_45010# 4.16e-21
C22025 a_10586_45546# a_11787_45002# 3.84e-19
C22026 a_n881_46662# a_11341_43940# 6.61e-21
C22027 a_2324_44458# a_14309_45348# 0.001898f
C22028 a_11823_42460# a_15037_45618# 0.099829f
C22029 a_n2840_45546# a_n2810_45028# 5.19e-19
C22030 a_n2661_45546# a_n913_45002# 9.6e-19
C22031 a_3090_45724# a_15433_44458# 0.001223f
C22032 a_12549_44172# a_18451_43940# 0.013387f
C22033 a_n2293_46098# a_2779_44458# 2.44e-20
C22034 a_10907_45822# a_11280_45822# 0.001255f
C22035 a_8049_45260# a_13556_45296# 8.2e-22
C22036 a_18479_47436# a_19594_46812# 0.108004f
C22037 a_18780_47178# a_19321_45002# 4.23e-20
C22038 a_6575_47204# a_2107_46812# 1.07e-19
C22039 VDAC_Pi a_5088_37509# 0.391059f
C22040 VDAC_Ni a_8530_39574# 1.72e-20
C22041 a_11453_44696# a_12549_44172# 0.066205f
C22042 a_n443_46116# a_2443_46660# 0.041057f
C22043 a_n1151_42308# a_3067_47026# 7.63e-19
C22044 a_3785_47178# a_3524_46660# 0.002172f
C22045 a_3815_47204# a_3699_46634# 2.44e-19
C22046 a_584_46384# a_3221_46660# 6.04e-20
C22047 a_n2216_40160# VDD 0.00515f
C22048 a_7754_40130# VDAC_N 0.434929f
C22049 a_n3565_39304# C3_P_btm 3.19e-20
C22050 a_n4064_39072# C7_P_btm 0.072179f
C22051 a_n3420_39072# C5_P_btm 0.001006f
C22052 a_19386_47436# a_13747_46662# 0.145228f
C22053 a_7754_39964# a_5700_37509# 0.095724f
C22054 a_12861_44030# a_n743_46660# 0.100542f
C22055 a_n1435_47204# a_n133_46660# 2.75e-20
C22056 a_n971_45724# a_6540_46812# 0.31827f
C22057 a_19479_31679# a_22459_39145# 1.76e-20
C22058 a_10949_43914# a_10518_42984# 2.24e-21
C22059 a_10729_43914# a_10835_43094# 4.2e-21
C22060 a_10405_44172# a_10796_42968# 1.23e-20
C22061 a_n356_44636# a_4921_42308# 8e-19
C22062 a_n2293_43922# COMP_P 0.151768f
C22063 a_n2810_45028# a_n2216_37690# 0.003507f
C22064 a_19963_31679# a_22469_40625# 1.59e-20
C22065 a_n2661_42834# a_n961_42308# 1.03e-20
C22066 a_16855_45546# VDD 0.339227f
C22067 a_6765_43638# a_6655_43762# 0.097745f
C22068 a_6547_43396# a_6452_43396# 0.049827f
C22069 a_n2956_37592# a_n2860_37690# 0.001388f
C22070 a_18494_42460# a_19647_42308# 0.030348f
C22071 a_18184_42460# a_13258_32519# 0.038977f
C22072 a_11967_42832# a_18504_43218# 0.015494f
C22073 a_3905_42865# a_n2293_42282# 4.89e-19
C22074 a_19741_43940# a_15743_43084# 4.79e-20
C22075 a_2711_45572# a_16979_44734# 6.79e-20
C22076 a_13059_46348# a_15037_43940# 4.6e-20
C22077 a_8049_45260# a_20362_44736# 1.72e-21
C22078 a_n1613_43370# a_n13_43084# 4.63e-20
C22079 a_5257_43370# a_5565_43396# 2.14e-19
C22080 a_n357_42282# a_5891_43370# 0.304889f
C22081 a_11525_45546# a_n2661_44458# 1.89e-19
C22082 a_2324_44458# a_5495_43940# 8.3e-21
C22083 a_413_45260# a_3429_45260# 4.84e-19
C22084 a_n913_45002# a_5205_44484# 4.56e-21
C22085 a_3483_46348# a_10807_43548# 1.08e-20
C22086 a_2274_45254# a_2382_45260# 0.130215f
C22087 a_10227_46804# a_12089_42308# 5.68e-19
C22088 a_7577_46660# a_6755_46942# 0.035922f
C22089 a_7715_46873# a_6969_46634# 3.3e-19
C22090 a_9863_46634# a_10428_46928# 0.042509f
C22091 SMPL_ON_P a_n1925_42282# 1.26e-19
C22092 a_19321_45002# a_18285_46348# 4.63e-22
C22093 a_13661_43548# a_20107_46660# 2.78e-20
C22094 a_13747_46662# a_19551_46910# 0.001463f
C22095 a_5807_45002# a_20411_46873# 1.37e-19
C22096 a_12549_44172# a_17639_46660# 0.129285f
C22097 a_n743_46660# a_14180_46812# 4.96e-20
C22098 a_5829_43940# a_5932_42308# 1.65e-20
C22099 a_15493_43396# a_15890_42674# 1.56e-21
C22100 a_5649_42852# a_8605_42826# 9.36e-21
C22101 a_n4318_39304# a_n1630_35242# 2.74e-20
C22102 a_4361_42308# a_8952_43230# 1.43e-20
C22103 a_n1699_44726# VDD 0.198612f
C22104 a_18783_43370# a_18249_42858# 3.47e-20
C22105 a_15743_43084# a_17333_42852# 2.59e-20
C22106 a_743_42282# a_10991_42826# 1.68e-19
C22107 a_19268_43646# a_18083_42858# 1.18e-19
C22108 a_15231_43396# a_5342_30871# 2.63e-19
C22109 a_n97_42460# COMP_P 7.27e-21
C22110 a_8685_43396# a_9061_43230# 7.37e-20
C22111 a_18597_46090# a_17303_42282# 4.04e-19
C22112 a_4185_45028# a_21487_43396# 2.21e-21
C22113 a_10809_44734# a_10341_43396# 4.7e-21
C22114 a_526_44458# a_8685_43396# 0.04962f
C22115 a_n2293_42834# a_8103_44636# 0.006106f
C22116 a_n2661_43370# a_742_44458# 2.53e-19
C22117 a_16922_45042# a_18545_45144# 0.001431f
C22118 a_4558_45348# a_n2661_43922# 6.4e-20
C22119 a_5147_45002# a_n2661_42834# 0.060392f
C22120 a_13249_42308# a_11750_44172# 3.55e-20
C22121 a_18184_42460# a_20193_45348# 0.074414f
C22122 a_21359_45002# a_11827_44484# 0.005947f
C22123 a_18494_42460# a_11691_44458# 1.03e-19
C22124 a_n1059_45260# a_17517_44484# 1.46e-20
C22125 a_20623_45572# a_20980_44850# 1.83e-20
C22126 a_17719_45144# a_17896_45144# 0.004187f
C22127 a_10193_42453# a_19862_44208# 0.099944f
C22128 w_1575_34946# a_3726_37500# 0.007105f
C22129 a_13507_46334# a_13904_45546# 2.05e-20
C22130 a_33_46660# a_n863_45724# 5.8e-20
C22131 a_n2293_46634# a_2957_45546# 0.001699f
C22132 a_n1925_46634# a_n755_45592# 7.2e-20
C22133 a_n743_46660# a_310_45028# 0.143623f
C22134 a_n2438_43548# a_n1099_45572# 7.2e-20
C22135 a_7577_46660# a_8049_45260# 4.87e-20
C22136 a_2107_46812# a_n2661_45546# 9.54e-20
C22137 a_15227_44166# a_18189_46348# 0.066472f
C22138 a_765_45546# a_5204_45822# 1.06e-19
C22139 a_12465_44636# a_11823_42460# 0.127538f
C22140 a_11453_44696# a_11525_45546# 5.01e-19
C22141 a_12991_46634# a_10809_44734# 0.008021f
C22142 a_13607_46688# a_6945_45028# 3.26e-20
C22143 a_19862_44208# VDD 0.588967f
C22144 a_3080_42308# a_3754_39134# 1.67e-20
C22145 a_8037_42858# a_5934_30871# 7.18e-19
C22146 a_4361_42308# a_15521_42308# 1.42e-19
C22147 a_4190_30871# a_18057_42282# 0.02374f
C22148 a_n2293_42282# a_n961_42308# 4.89e-19
C22149 a_743_42282# a_17303_42282# 0.034786f
C22150 a_n310_47570# VDD 3.35e-19
C22151 a_22612_30879# a_22469_39537# 1.3e-19
C22152 a_4883_46098# DATA[5] 2.29e-20
C22153 a_4574_45260# a_n97_42460# 9.85e-22
C22154 a_327_44734# a_458_43396# 1.92e-21
C22155 a_4185_45028# a_5932_42308# 0.118319f
C22156 a_1307_43914# a_9420_43940# 9.31e-19
C22157 a_2779_44458# a_2675_43914# 1.27e-19
C22158 a_742_44458# a_2998_44172# 1.08e-19
C22159 a_3357_43084# a_6031_43396# 0.001792f
C22160 a_13249_42308# a_4361_42308# 0.009442f
C22161 a_n357_42282# a_17595_43084# 0.007854f
C22162 a_n443_42852# a_10341_42308# 2.65e-20
C22163 a_13507_46334# CLK 8.83e-20
C22164 a_n2840_44458# a_n4318_39768# 0.007737f
C22165 a_n699_43396# a_2479_44172# 0.063139f
C22166 en_comp a_3080_42308# 1.28517f
C22167 a_n2661_42834# a_12553_44484# 4.92e-20
C22168 a_n2661_43922# a_12189_44484# 1.22e-19
C22169 a_13556_45296# a_15037_43940# 0.001578f
C22170 a_13777_45326# a_13565_43940# 1.03e-20
C22171 a_1823_45246# a_3905_42308# 0.003168f
C22172 a_18479_47436# a_18494_42460# 2.53e-21
C22173 a_9290_44172# a_n357_42282# 0.138435f
C22174 a_n2293_46634# a_9482_43914# 6.32e-20
C22175 a_18819_46122# a_19443_46116# 9.73e-19
C22176 a_19335_46494# a_19597_46482# 0.001705f
C22177 a_19553_46090# a_20009_46494# 4.2e-19
C22178 a_6945_45028# a_16375_45002# 3.78e-20
C22179 a_2107_46812# a_5205_44484# 1.38e-20
C22180 a_167_45260# a_1609_45572# 2.26e-19
C22181 a_2443_46660# a_3537_45260# 3.5e-19
C22182 a_n1151_42308# a_6298_44484# 0.009717f
C22183 a_15227_44166# a_17478_45572# 0.009301f
C22184 a_18597_46090# a_19778_44110# 0.006796f
C22185 a_7715_46873# a_3357_43084# 6.39e-20
C22186 a_n443_46116# a_949_44458# 0.045448f
C22187 a_3177_46902# a_3065_45002# 8.4e-21
C22188 a_2609_46660# a_3429_45260# 6.06e-22
C22189 a_1823_45246# a_3175_45822# 2.41e-19
C22190 a_13467_32519# VIN_N 0.078487f
C22191 a_n3674_37592# a_n2302_40160# 6.29e-20
C22192 a_n2157_42858# VDD 0.424058f
C22193 a_13720_44458# a_9145_43396# 6.13e-21
C22194 a_n2810_45572# a_n4064_40160# 7.36e-19
C22195 a_n1059_45260# a_4149_42891# 4.67e-19
C22196 a_20820_30879# C5_N_btm 1.83e-19
C22197 a_11827_44484# a_16823_43084# 4.84e-20
C22198 a_9482_43914# a_5342_30871# 5.46e-21
C22199 a_10193_42453# a_9803_42558# 0.20198f
C22200 a_n2661_43922# a_1756_43548# 5.14e-21
C22201 a_n2661_42834# a_4093_43548# 1.69e-19
C22202 a_n2293_42834# a_n722_43218# 2.66e-19
C22203 a_18494_42460# a_4190_30871# 0.242908f
C22204 a_18184_42460# a_20301_43646# 6.85e-19
C22205 a_18900_46660# START 2.58e-19
C22206 a_21350_47026# VDD 4.6e-19
C22207 a_9313_44734# a_2982_43646# 0.027994f
C22208 a_21363_46634# EN_OFFSET_CAL 4.24e-21
C22209 a_7499_43078# a_10545_42558# 0.003046f
C22210 a_n357_42282# a_21887_42336# 3.8e-20
C22211 a_9838_44484# a_9885_43646# 4.23e-22
C22212 a_4185_45028# a_1423_45028# 0.016283f
C22213 a_3090_45724# a_5343_44458# 0.023693f
C22214 a_11415_45002# a_n2661_43370# 0.092334f
C22215 a_n1613_43370# a_644_44056# 1.52e-20
C22216 a_9290_44172# a_11963_45334# 1.31e-19
C22217 a_2711_45572# a_11823_42460# 0.065343f
C22218 a_15015_46420# a_6171_45002# 2.21e-20
C22219 a_2324_44458# a_5691_45260# 0.013607f
C22220 a_6945_45028# a_413_45260# 1.33e-19
C22221 a_13747_46662# a_20980_44850# 0.001171f
C22222 a_8049_45260# a_21363_45546# 0.013686f
C22223 a_13259_45724# a_16377_45572# 0.002102f
C22224 a_9625_46129# a_9482_43914# 2.09e-19
C22225 a_n746_45260# a_1443_43940# 3.72e-20
C22226 a_21887_42336# CAL_N 8.2e-19
C22227 a_n3565_39590# a_n3420_37440# 0.035128f
C22228 a_5932_42308# VREF_GND 0.001404f
C22229 a_n4209_39590# a_n4064_37440# 0.033425f
C22230 a_5742_30871# C4_N_btm 0.03103f
C22231 a_13258_32519# a_22459_39145# 2.2e-19
C22232 a_n4064_40160# a_n4251_37440# 0.001069f
C22233 a_9803_42558# VDD 0.253745f
C22234 a_n3420_39616# a_n3565_37414# 0.028804f
C22235 a_n4064_39616# a_n4209_37414# 0.028043f
C22236 a_n2302_38778# a_n2302_37984# 0.052227f
C22237 a_n237_47217# a_768_44030# 7.54e-19
C22238 a_2905_45572# a_n1613_43370# 0.044171f
C22239 a_3785_47178# a_4842_47570# 9.52e-19
C22240 a_3160_47472# a_3411_47243# 4.21e-19
C22241 a_n1151_42308# a_3094_47243# 3.77e-19
C22242 a_11599_46634# a_19386_47436# 1.17e-21
C22243 a_16763_47508# a_16588_47582# 0.233657f
C22244 a_16327_47482# a_10227_46804# 0.630403f
C22245 a_13381_47204# a_4883_46098# 7.29e-21
C22246 a_13717_47436# a_13507_46334# 3.3e-19
C22247 a_14539_43914# a_17665_42852# 0.003264f
C22248 a_n97_42460# a_1568_43370# 0.074153f
C22249 a_20974_43370# a_2982_43646# 0.051776f
C22250 a_n2433_43396# a_n1557_42282# 2.44e-21
C22251 a_n2956_37592# a_n4064_39072# 0.010695f
C22252 a_6667_45809# VDD 0.195842f
C22253 a_18079_43940# a_17499_43370# 0.001409f
C22254 a_15493_43396# a_16547_43609# 0.022221f
C22255 a_14021_43940# a_14358_43442# 0.007211f
C22256 a_n2810_45028# a_n2302_39072# 4.97e-19
C22257 a_n356_44636# a_13291_42460# 1.18e-19
C22258 a_17517_44484# a_19987_42826# 6.08e-21
C22259 a_11967_42832# a_16414_43172# 0.058563f
C22260 a_13507_46334# a_19268_43646# 2.35e-21
C22261 a_8696_44636# a_5111_44636# 3.25e-20
C22262 a_20273_45572# a_19963_31679# 0.001592f
C22263 a_21188_45572# a_22223_45572# 9.49e-20
C22264 a_20528_45572# a_2437_43646# 8.27e-22
C22265 a_12861_44030# a_4361_42308# 0.005354f
C22266 a_12549_44172# a_9145_43396# 6.67e-19
C22267 a_19466_46812# a_20365_43914# 5.98e-19
C22268 a_n2956_39304# a_n2661_42834# 5.57e-20
C22269 a_n2293_46634# a_6031_43396# 0.037881f
C22270 a_16333_45814# a_6171_45002# 3.41e-19
C22271 a_16327_47482# a_19177_43646# 7.13e-19
C22272 a_n971_45724# a_7871_42858# 2.7e-19
C22273 a_584_46384# a_791_42968# 4.57e-19
C22274 a_20623_45572# a_3357_43084# 0.041244f
C22275 a_n2956_38216# a_n2840_44458# 0.004419f
C22276 a_n2661_45546# a_n2661_44458# 0.032856f
C22277 a_2711_45572# a_16321_45348# 7.82e-19
C22278 a_10809_44734# a_n2293_43922# 2.24e-19
C22279 a_15015_46420# a_14673_44172# 2.63e-21
C22280 a_n2661_46098# a_2162_46660# 0.003322f
C22281 a_n2109_47186# a_3483_46348# 0.03221f
C22282 a_n1532_35090# VIN_P 0.066301f
C22283 C7_P_btm VDD 0.121904f
C22284 a_18479_47436# a_16388_46812# 5.74e-20
C22285 a_n971_45724# a_1823_45246# 0.514159f
C22286 a_768_44030# a_8270_45546# 0.03575f
C22287 a_2905_45572# a_n2293_46098# 0.028964f
C22288 a_n881_46662# a_12991_46634# 1.56e-19
C22289 a_13507_46334# a_14035_46660# 0.027121f
C22290 a_16327_47482# a_17339_46660# 0.058779f
C22291 a_16241_47178# a_765_45546# 0.004102f
C22292 a_2107_46812# a_5385_46902# 0.001613f
C22293 a_3177_46902# a_3067_47026# 0.097745f
C22294 a_3699_46634# a_3524_46660# 0.233657f
C22295 a_2959_46660# a_2864_46660# 0.049827f
C22296 a_n1925_46634# a_5429_46660# 4.33e-19
C22297 a_n2661_46634# a_7927_46660# 0.00501f
C22298 C3_P_btm C8_N_btm 0.001059f
C22299 C1_P_btm C6_N_btm 3.17e-19
C22300 C0_P_btm C5_N_btm 1.4e-19
C22301 a_11599_46634# a_19551_46910# 5.02e-19
C22302 C0_dummy_P_btm C4_N_btm 1.24e-19
C22303 C0_N_btm C2_N_btm 0.698973f
C22304 C0_dummy_N_btm C3_N_btm 0.087593f
C22305 a_13717_47436# a_20623_46660# 2.48e-20
C22306 a_4915_47217# a_11415_45002# 0.134061f
C22307 a_n237_47217# a_1176_45822# 3.23e-19
C22308 a_n746_45260# a_1138_42852# 6.98e-20
C22309 a_327_47204# a_472_46348# 7.59e-19
C22310 a_11967_42832# a_7174_31319# 5.83e-20
C22311 a_2448_45028# VDD 0.004293f
C22312 a_16823_43084# a_17433_43396# 8.76e-19
C22313 a_8685_43396# a_8605_42826# 0.001894f
C22314 a_3626_43646# a_18249_42858# 4.73e-20
C22315 a_2982_43646# a_18599_43230# 2.4e-20
C22316 a_4093_43548# a_n2293_42282# 5.81e-20
C22317 a_19700_43370# a_4361_42308# 7.65e-21
C22318 a_18783_43370# a_5649_42852# 1.76e-21
C22319 a_15743_43084# a_13678_32519# 0.020598f
C22320 a_10903_43370# a_3626_43646# 0.001928f
C22321 a_2382_45260# a_4743_44484# 5.73e-20
C22322 a_n357_42282# a_10807_43548# 0.031251f
C22323 a_5937_45572# a_6197_43396# 2.15e-19
C22324 a_2324_44458# a_3080_42308# 1.53e-21
C22325 a_13777_45326# a_11691_44458# 5.49e-20
C22326 a_15415_45028# a_11827_44484# 5.8e-21
C22327 a_n443_42852# a_3499_42826# 0.023367f
C22328 a_3065_45002# a_4223_44672# 0.001102f
C22329 a_2680_45002# a_n699_43396# 2.59e-19
C22330 a_n2312_40392# a_n3674_37592# 0.035844f
C22331 a_5205_44484# a_n2661_44458# 0.072981f
C22332 a_16721_46634# a_765_45546# 0.002907f
C22333 a_8492_46660# a_8016_46348# 7.47e-19
C22334 a_2063_45854# a_7499_43078# 0.478913f
C22335 a_7227_47204# a_6472_45840# 4.49e-20
C22336 a_6851_47204# a_6511_45714# 1.94e-21
C22337 a_6545_47178# a_6598_45938# 9.57e-19
C22338 a_6491_46660# a_6667_45809# 1.51e-21
C22339 a_n443_46116# a_1990_45572# 3.19e-20
C22340 a_6151_47436# a_7227_45028# 0.006424f
C22341 a_19692_46634# a_20719_46660# 0.004558f
C22342 a_n743_46660# a_3873_46454# 2.25e-19
C22343 a_4646_46812# a_2324_44458# 0.023652f
C22344 a_5807_45002# a_10044_46482# 5.69e-19
C22345 a_9313_45822# a_2711_45572# 0.016843f
C22346 a_16388_46812# a_17829_46910# 1.39e-19
C22347 a_15227_44166# a_20202_43084# 0.086371f
C22348 a_12281_43396# a_13070_42354# 5.19e-19
C22349 a_17364_32525# a_n1630_35242# 1.85e-20
C22350 a_n901_43156# COMP_P 8.12e-21
C22351 a_n1641_43230# a_n1329_42308# 0.004511f
C22352 a_15095_43370# a_15051_42282# 0.003143f
C22353 a_14955_43396# a_14113_42308# 1.29e-21
C22354 a_n1761_44111# VDD 0.620042f
C22355 a_n3674_39304# a_n3674_38216# 0.023464f
C22356 a_n1736_43218# a_n4318_38216# 3.63e-19
C22357 a_12379_42858# a_13291_42460# 6.47e-20
C22358 a_13113_42826# a_13569_43230# 4.2e-19
C22359 a_13678_32519# a_1606_42308# 6.06e-20
C22360 a_743_42282# a_2713_42308# 0.024879f
C22361 a_n4318_39304# a_n3607_39392# 8.54e-20
C22362 a_10193_42453# a_14579_43548# 5.04e-21
C22363 a_11827_44484# a_19279_43940# 0.078733f
C22364 a_6171_45002# a_15493_43396# 1.54e-20
C22365 a_2711_45572# a_18429_43548# 2.62e-20
C22366 a_n2956_39304# a_n2293_42282# 4.17e-20
C22367 a_1239_47204# VDD 0.278979f
C22368 a_10057_43914# a_10617_44484# 0.033364f
C22369 a_9838_44484# a_n2661_43922# 0.006262f
C22370 a_10157_44484# a_n2661_42834# 6.22e-20
C22371 a_14539_43914# a_9313_44734# 0.016028f
C22372 a_20107_45572# a_19319_43548# 3.02e-20
C22373 a_11787_45002# a_11750_44172# 8e-19
C22374 a_9482_43914# a_9672_43914# 0.122568f
C22375 a_5093_45028# a_3905_42865# 2.69e-19
C22376 a_19778_44110# a_19789_44512# 7.63e-19
C22377 a_n971_45724# DATA[2] 0.099284f
C22378 a_n357_42282# a_13467_32519# 0.002449f
C22379 a_n443_42852# a_15940_43402# 0.005303f
C22380 a_n1741_47186# CLK 0.028114f
C22381 a_9290_44172# a_10553_43218# 0.002152f
C22382 a_n2312_38680# a_n2946_38778# 0.024631f
C22383 a_3090_45724# a_12563_42308# 4.38e-21
C22384 a_n2293_42834# a_895_43940# 7.7e-20
C22385 a_n2661_43370# a_n984_44318# 7.79e-21
C22386 a_20193_45348# a_20362_44736# 0.013057f
C22387 a_626_44172# a_2253_44260# 6.94e-21
C22388 a_n356_44636# a_700_44734# 4.08e-19
C22389 a_n746_45260# DATA[1] 5.22e-20
C22390 a_n237_47217# DATA[0] 0.040942f
C22391 a_5937_45572# a_5066_45546# 0.419426f
C22392 a_10428_46928# a_10210_45822# 2.06e-20
C22393 a_768_44030# a_n2017_45002# 1.14e-19
C22394 a_12549_44172# a_n1059_45260# 2.03e-19
C22395 a_n881_46662# a_n143_45144# 7.46e-19
C22396 a_13747_46662# a_3357_43084# 7.23e-19
C22397 a_4883_46098# a_8953_45002# 0.013985f
C22398 a_16327_47482# a_1307_43914# 3.53e-20
C22399 a_20075_46420# a_19900_46494# 0.233657f
C22400 a_18985_46122# a_6945_45028# 1.4e-20
C22401 a_3090_45724# a_4880_45572# 0.002202f
C22402 a_10227_46804# a_14537_43396# 0.094463f
C22403 a_19594_46812# a_2437_43646# 0.003991f
C22404 a_1606_42308# a_6123_31319# 1.43958f
C22405 a_3823_42558# a_4921_42308# 0.001205f
C22406 a_14579_43548# VDD 0.278225f
C22407 a_5649_42852# VDAC_N 3.45e-20
C22408 a_n784_42308# a_9803_42558# 2.06e-20
C22409 a_16877_43172# a_4958_30871# 1.48e-19
C22410 a_13467_32519# CAL_N 2.02e-19
C22411 a_n863_45724# a_5934_30871# 2.07e-20
C22412 a_n2956_39304# a_n3565_39590# 0.072956f
C22413 a_13249_42308# a_13622_42852# 1.85e-19
C22414 a_5883_43914# a_n97_42460# 5.99e-19
C22415 a_n699_43396# a_n229_43646# 0.043893f
C22416 a_1115_44172# a_895_43940# 0.029554f
C22417 a_1414_42308# a_2127_44172# 0.091064f
C22418 a_1467_44172# a_2479_44172# 2.93e-20
C22419 a_18443_44721# a_18533_43940# 6.51e-20
C22420 a_18989_43940# a_19808_44306# 1.9e-20
C22421 a_n913_45002# a_4520_42826# 0.001583f
C22422 a_n1059_45260# a_5111_42852# 0.005242f
C22423 a_n2017_45002# a_5755_42852# 1.59e-20
C22424 a_n443_42852# a_3318_42354# 1.12e-21
C22425 a_13259_45724# a_13657_42558# 0.023664f
C22426 a_11186_47026# VDD 0.077608f
C22427 a_742_44458# a_1568_43370# 0.525694f
C22428 a_949_44458# a_1049_43396# 0.001408f
C22429 a_n755_45592# a_n310_45572# 0.001154f
C22430 a_n971_45724# a_n3674_39768# 2.61e-20
C22431 a_n1853_46287# a_n467_45028# 1.67e-19
C22432 a_167_45260# a_n2661_45010# 6.95e-20
C22433 a_18479_47436# a_20640_44752# 0.018112f
C22434 a_16327_47482# a_18579_44172# 0.043297f
C22435 a_1848_45724# a_1990_45899# 0.005572f
C22436 a_310_45028# a_509_45572# 1.27e-19
C22437 a_n1099_45572# a_603_45572# 3.32e-19
C22438 a_12839_46116# a_10193_42453# 2.22e-20
C22439 a_n2497_47436# a_1241_44260# 0.001773f
C22440 a_n2293_46098# a_n37_45144# 4.54e-20
C22441 a_5164_46348# a_2437_43646# 3.03e-20
C22442 a_n863_45724# a_1609_45572# 1.88e-19
C22443 a_n2661_45546# a_5907_45546# 3.27e-19
C22444 a_17583_46090# a_16147_45260# 1.41e-20
C22445 a_17715_44484# a_17786_45822# 0.001664f
C22446 a_18597_46090# a_20159_44458# 1.48e-20
C22447 a_11453_44696# a_17061_44734# 0.005756f
C22448 a_584_46384# a_3905_42865# 4.97e-20
C22449 a_n3420_39616# a_n4209_39304# 0.05141f
C22450 a_n4209_39590# a_n3420_39072# 0.034738f
C22451 a_n4064_39616# a_n3607_39616# 7.1e-19
C22452 a_n784_42308# C7_P_btm 0.002308f
C22453 a_1606_42308# EN_VIN_BSTR_P 0.035204f
C22454 a_2952_47436# a_n443_46116# 9.06e-19
C22455 a_2905_45572# a_4791_45118# 0.001355f
C22456 a_3381_47502# a_3815_47204# 0.021997f
C22457 a_n1151_42308# a_4007_47204# 0.015013f
C22458 a_n237_47217# a_9067_47204# 0.0235f
C22459 SMPL_ON_P a_n1435_47204# 0.082028f
C22460 a_2063_45854# a_5129_47502# 9.87e-20
C22461 a_n1741_47186# a_13717_47436# 6.56e-20
C22462 a_n4064_40160# a_n4251_39392# 0.001069f
C22463 a_n3565_39590# a_n3565_39304# 0.046203f
C22464 a_5934_30871# a_6886_37412# 3.68e-19
C22465 a_n1630_35242# a_21589_35634# 0.015148f
C22466 a_n2293_42834# a_n3674_38216# 0.001875f
C22467 a_3065_45002# a_5742_30871# 1.24e-20
C22468 en_comp a_15764_42576# 5.59e-20
C22469 a_10586_45546# CLK 0.125859f
C22470 a_n2661_42834# a_685_42968# 1.91e-21
C22471 a_9313_44734# a_7871_42858# 1.01e-19
C22472 a_1307_43914# a_5267_42460# 9.19e-21
C22473 a_11967_42832# a_21487_43396# 1.24e-20
C22474 a_18248_44752# a_18083_42858# 1.84e-20
C22475 a_5891_43370# a_8952_43230# 0.016573f
C22476 a_17970_44736# a_17333_42852# 5.58e-21
C22477 a_20640_44752# a_4190_30871# 5.05e-22
C22478 a_20679_44626# a_21259_43561# 9.33e-20
C22479 a_14539_43914# a_18599_43230# 1.28e-19
C22480 a_12839_46116# VDD 0.347766f
C22481 a_13925_46122# a_13720_44458# 1.08e-20
C22482 a_n443_42852# a_13777_45326# 1.94e-21
C22483 a_2711_45572# a_7705_45326# 0.001295f
C22484 a_8049_45260# a_19778_44110# 2.13e-20
C22485 a_3483_46348# a_8375_44464# 0.003197f
C22486 a_n1613_43370# a_104_43370# 1.95e-19
C22487 a_4883_46098# a_3626_43646# 4.8e-20
C22488 a_2324_44458# a_10057_43914# 1.41e-19
C22489 a_6511_45714# a_3232_43370# 5.46e-20
C22490 a_6472_45840# a_6171_45002# 0.005155f
C22491 a_11322_45546# a_n913_45002# 4.81e-21
C22492 a_n755_45592# a_2232_45348# 1.57e-19
C22493 a_5907_45546# a_5205_44484# 2.98e-20
C22494 a_12741_44636# a_15463_44811# 2.47e-19
C22495 a_13661_43548# a_18797_44260# 0.002056f
C22496 a_8270_45546# a_7845_44172# 1.29e-19
C22497 a_16020_45572# a_16211_45572# 4.61e-19
C22498 a_16855_45546# a_18479_45785# 1.38e-20
C22499 a_8696_44636# a_16147_45260# 0.284694f
C22500 a_16680_45572# a_18175_45572# 4.94e-20
C22501 a_n3420_37440# C4_P_btm 2.18e-19
C22502 a_n4064_37440# C6_P_btm 1.49e-19
C22503 a_15507_47210# a_6755_46942# 2.7e-19
C22504 a_20916_46384# a_22612_30879# 3.3e-20
C22505 a_n1741_47186# a_14035_46660# 2.61e-20
C22506 a_n1151_42308# a_15368_46634# 2.09e-19
C22507 a_n1613_43370# a_2443_46660# 0.917984f
C22508 a_7754_39300# VDD 0.048307f
C22509 a_n881_46662# a_n2661_46098# 0.096736f
C22510 a_6151_47436# a_11813_46116# 8.68e-20
C22511 a_9067_47204# a_8270_45546# 9.93e-19
C22512 a_3785_47178# a_3090_45724# 4.4e-22
C22513 a_4915_47217# a_12251_46660# 2.85e-19
C22514 a_9313_45822# a_8654_47026# 4.81e-20
C22515 a_10227_46804# a_8667_46634# 6.04e-20
C22516 a_22469_39537# a_22780_39857# 1.79e-19
C22517 VDAC_P a_n923_35174# 0.015621f
C22518 a_22459_39145# a_22609_37990# 0.172129f
C22519 a_22469_40625# a_22717_36887# 0.011861f
C22520 a_22521_40055# a_22705_37990# 0.016815f
C22521 a_22521_39511# a_22609_38406# 0.23688f
C22522 a_19237_31679# a_n1630_35242# 7.69e-20
C22523 a_n2956_37592# VDD 1.25966f
C22524 a_10341_43396# a_14621_43646# 4.92e-19
C22525 a_19963_31679# VREF 0.055795f
C22526 a_n1761_44111# a_n784_42308# 0.034368f
C22527 a_n356_44636# a_18548_42308# 4.18e-20
C22528 a_6031_43396# a_743_42282# 4.36e-20
C22529 a_14955_43396# a_15781_43660# 1.56e-19
C22530 a_3626_43646# a_5649_42852# 0.032897f
C22531 a_n97_42460# a_133_43172# 0.002798f
C22532 a_14021_43940# a_22165_42308# 6.79e-20
C22533 a_14579_43548# a_16137_43396# 6.3e-20
C22534 a_6431_45366# a_6517_45366# 0.006584f
C22535 a_21363_45546# a_20193_45348# 1.77e-22
C22536 a_12549_44172# a_19987_42826# 6.54e-20
C22537 a_n971_45724# a_1184_42692# 2.87e-20
C22538 a_15227_44166# a_14955_43396# 0.001876f
C22539 a_15415_45028# a_15595_45028# 0.185422f
C22540 a_14537_43396# a_1307_43914# 0.0516f
C22541 a_15037_45618# a_14539_43914# 4.54e-21
C22542 a_8696_44636# a_10334_44484# 0.001709f
C22543 a_3065_45002# a_n2293_42834# 0.021132f
C22544 a_19479_31679# a_19778_44110# 1.24e-19
C22545 a_21513_45002# a_20567_45036# 2e-19
C22546 a_10227_46804# a_12991_43230# 1.79e-19
C22547 a_13661_43548# a_15567_42826# 1.39e-23
C22548 a_5147_45002# a_5093_45028# 0.008723f
C22549 a_5111_44636# a_5009_45028# 8.57e-19
C22550 a_7499_43078# a_n2661_42834# 0.089963f
C22551 a_n467_45028# a_n2661_43370# 0.016799f
C22552 a_2324_44458# a_14021_43940# 8.72e-19
C22553 a_n2293_46634# a_10796_42968# 6.09e-20
C22554 a_15009_46634# a_14976_45028# 0.071873f
C22555 a_12549_44172# a_13925_46122# 5.78e-20
C22556 a_768_44030# a_13759_46122# 0.024686f
C22557 a_n815_47178# a_n863_45724# 2.42e-20
C22558 a_9804_47204# a_2324_44458# 1.14e-19
C22559 a_5807_45002# a_9823_46155# 0.005199f
C22560 a_n743_46660# a_2804_46116# 0.012952f
C22561 a_2443_46660# a_n2293_46098# 1.88e-20
C22562 a_1123_46634# a_1176_45822# 0.001261f
C22563 a_948_46660# a_1208_46090# 3.04e-19
C22564 a_2107_46812# a_805_46414# 1.28e-19
C22565 a_4915_47217# a_13259_45724# 0.04489f
C22566 a_n2661_46634# a_5164_46348# 1.31e-19
C22567 a_n971_45724# a_n2293_45546# 0.097168f
C22568 a_n1925_46634# a_3483_46348# 4.03e-19
C22569 a_n2661_46098# a_n2157_46122# 0.227082f
C22570 a_n1741_47186# a_n1099_45572# 2.08e-20
C22571 a_2982_43646# a_8515_42308# 1.02e-19
C22572 a_685_42968# a_n2293_42282# 2.16e-20
C22573 a_15743_43084# a_15597_42852# 0.055955f
C22574 a_n97_42460# a_13333_42558# 1.53e-20
C22575 a_3539_42460# a_6123_31319# 9e-21
C22576 a_3626_43646# a_7963_42308# 0.003306f
C22577 a_12545_42858# a_12895_43230# 0.215953f
C22578 a_12379_42858# a_13460_43230# 0.102325f
C22579 a_5708_44484# VDD 9.68e-19
C22580 a_n2661_43370# a_n2661_43922# 0.13591f
C22581 a_413_45260# a_895_43940# 0.001706f
C22582 a_n2293_45010# a_n3674_39768# 6.8e-20
C22583 a_2437_43646# a_3499_42826# 1.38e-20
C22584 a_2324_44458# a_2075_43172# 1.36e-20
C22585 a_9290_44172# a_8952_43230# 2.21e-19
C22586 a_5257_43370# a_5932_42308# 3.61e-20
C22587 a_4743_44484# a_5343_44458# 4.42e-19
C22588 a_4223_44672# a_6298_44484# 3.26e-19
C22589 a_18479_45785# a_19862_44208# 2.98e-20
C22590 a_n2312_39304# a_n4064_39072# 0.094407f
C22591 a_n1059_45260# a_7542_44172# 5.06e-21
C22592 a_n443_42852# a_6197_43396# 0.007993f
C22593 a_8199_44636# a_10341_42308# 1.19e-19
C22594 a_4185_45028# a_15567_42826# 9.4e-21
C22595 a_2711_45572# a_2982_43646# 9.28e-19
C22596 a_2382_45260# a_1414_42308# 0.005789f
C22597 a_18597_46090# a_20623_45572# 0.046479f
C22598 a_n743_46660# a_13904_45546# 1.24e-20
C22599 a_n443_46116# a_n143_45144# 0.001224f
C22600 a_4700_47436# a_413_45260# 8.97e-20
C22601 a_n881_46662# a_16020_45572# 0.013745f
C22602 a_18479_47436# a_21188_45572# 0.005114f
C22603 a_16327_47482# a_20885_45572# 0.002535f
C22604 a_4646_46812# a_6667_45809# 3.86e-19
C22605 a_3877_44458# a_6598_45938# 4.85e-19
C22606 a_12741_44636# a_21137_46414# 2.81e-21
C22607 a_3483_46348# a_10355_46116# 1.51e-21
C22608 a_12549_44172# a_15599_45572# 5.18e-22
C22609 a_2905_45572# a_3429_45260# 4.46e-19
C22610 a_3160_47472# a_3065_45002# 1.34e-21
C22611 a_11415_45002# a_10809_44734# 0.140489f
C22612 a_2063_45854# a_4558_45348# 8.06e-22
C22613 a_5167_46660# a_5263_45724# 4.57e-21
C22614 a_15673_47210# a_2437_43646# 0.007104f
C22615 a_11599_46634# a_3357_43084# 9.81e-19
C22616 a_10227_46804# a_20731_45938# 8.16e-20
C22617 a_20894_47436# a_20107_45572# 1.49e-21
C22618 a_11453_44696# a_19431_45546# 3.07e-21
C22619 a_3080_42308# C7_P_btm 0.002948f
C22620 a_n3674_38680# a_n4318_38216# 2.82961f
C22621 a_n2267_43396# VDD 0.570924f
C22622 a_17701_42308# a_17124_42282# 5.83e-19
C22623 a_5342_30871# a_4958_30871# 10.9366f
C22624 a_n3674_39304# a_n4251_39616# 5.77e-20
C22625 a_n2293_42834# a_458_43396# 0.003568f
C22626 a_1307_43914# a_6547_43396# 1.88e-19
C22627 a_11967_42832# a_21398_44850# 0.01381f
C22628 a_n743_46660# CLK 0.028835f
C22629 a_8953_45002# a_8685_43396# 6.4e-21
C22630 a_17517_44484# a_22959_44484# 0.00251f
C22631 a_n2661_43922# a_2998_44172# 0.003621f
C22632 a_n2661_42834# a_3600_43914# 0.012088f
C22633 a_16979_44734# a_15682_43940# 0.001729f
C22634 a_14539_43914# a_17737_43940# 5.43e-19
C22635 a_526_44458# a_6123_31319# 1.83e-19
C22636 a_20205_31679# a_22400_42852# 4.56e-20
C22637 a_4185_45028# a_20712_42282# 1.64e-19
C22638 a_5708_44484# a_5495_43940# 1.89e-19
C22639 a_20362_44736# a_20596_44850# 0.006453f
C22640 a_3537_45260# a_10341_43396# 4.95e-20
C22641 a_491_47026# VDD 0.132552f
C22642 a_n2017_45002# a_16759_43396# 1.39e-21
C22643 a_n913_45002# a_16409_43396# 9.35e-21
C22644 a_n1059_45260# a_16977_43638# 1.07e-19
C22645 a_20107_46660# a_20273_45572# 0.001469f
C22646 a_20411_46873# a_20107_45572# 0.001307f
C22647 a_16388_46812# a_2437_43646# 1.36e-19
C22648 a_11453_44696# a_13076_44458# 9.33e-21
C22649 a_2324_44458# a_10180_45724# 0.064932f
C22650 a_1799_45572# a_n2661_43370# 9.48e-20
C22651 a_9290_44172# a_13249_42308# 0.033421f
C22652 a_8199_44636# a_8336_45822# 2.62e-19
C22653 a_5937_45572# a_6977_45572# 4.29e-19
C22654 a_15559_46634# a_413_45260# 2.31e-21
C22655 a_12465_44636# a_14539_43914# 0.054102f
C22656 a_12594_46348# a_12427_45724# 0.040872f
C22657 a_6755_46942# a_9482_43914# 0.01168f
C22658 a_19321_45002# a_11691_44458# 0.064467f
C22659 a_n1613_43370# a_949_44458# 6.55e-22
C22660 a_13661_43548# a_16886_45144# 2.62e-21
C22661 a_11415_45002# a_16211_45572# 8.47e-19
C22662 a_n743_46660# a_17023_45118# 5.2e-19
C22663 a_12005_46116# a_11823_42460# 0.010777f
C22664 a_5257_43370# a_1423_45028# 0.020778f
C22665 a_10903_43370# a_12791_45546# 0.042213f
C22666 a_10227_46804# a_n356_44636# 4.54e-19
C22667 a_13507_46334# a_18248_44752# 1.76e-21
C22668 a_17303_42282# a_13258_32519# 0.064259f
C22669 a_5342_30871# VCM 0.325566f
C22670 a_21671_42860# VDD 0.229963f
C22671 a_18057_42282# a_19511_42282# 1.23e-20
C22672 a_21195_42852# RST_Z 4.44e-21
C22673 a_6123_31319# a_n4209_38502# 6.28e-22
C22674 a_2889_44172# a_n97_42460# 2.34e-20
C22675 a_11189_46129# CLK 3.69e-19
C22676 a_8333_44056# a_8415_44056# 0.004999f
C22677 a_9313_44734# a_17324_43396# 2.24e-20
C22678 a_11827_44484# a_12545_42858# 1.69e-22
C22679 a_19862_44208# a_14021_43940# 0.021104f
C22680 a_n1059_45260# a_n1630_35242# 0.007613f
C22681 a_n2017_45002# a_1067_42314# 0.01039f
C22682 a_14840_46494# VDD 0.275785f
C22683 a_n967_45348# a_n473_42460# 9.24e-19
C22684 a_n913_45002# a_564_42282# 1.62e-19
C22685 a_15015_46420# RST_Z 4.05e-21
C22686 a_526_44458# a_3495_45348# 0.002123f
C22687 a_n1151_42308# a_n229_43646# 4.13e-20
C22688 a_n443_46116# a_n97_42460# 0.131756f
C22689 a_584_46384# a_4093_43548# 0.00472f
C22690 a_12861_44030# a_18533_43940# 1.12e-19
C22691 a_n1423_46090# a_n1177_44458# 9.12e-21
C22692 a_10193_42453# a_16115_45572# 0.001215f
C22693 a_n863_45724# a_n2661_45010# 0.345234f
C22694 a_10586_45546# a_10951_45334# 2.24e-20
C22695 a_2324_44458# a_13711_45394# 6.14e-19
C22696 a_11823_42460# a_14033_45822# 0.093809f
C22697 a_9049_44484# a_8696_44636# 0.043734f
C22698 a_3316_45546# a_2437_43646# 7.08e-22
C22699 a_n2661_45546# a_n1059_45260# 0.003807f
C22700 a_n2293_46098# a_949_44458# 4.44e-20
C22701 a_3090_45724# a_14815_43914# 9.92e-21
C22702 a_n2293_45546# a_n2293_45010# 0.257189f
C22703 a_20692_30879# en_comp 2.56e-19
C22704 a_12549_44172# a_18326_43940# 0.013334f
C22705 a_8336_45822# a_8192_45572# 6.84e-19
C22706 a_8049_45260# a_9482_43914# 2.04e-21
C22707 VDAC_Ni a_7754_38470# 0.005657f
C22708 VDAC_Pi a_4338_37500# 1.92369f
C22709 a_n4251_40480# VDD 3.95e-19
C22710 a_7754_40130# a_6886_37412# 0.006212f
C22711 a_n3565_39304# C4_P_btm 5.85e-20
C22712 a_n3420_39072# C6_P_btm 0.054459f
C22713 a_n4064_39072# C8_P_btm 7.96e-19
C22714 a_7754_39964# a_5088_37509# 0.392826f
C22715 a_n4209_38502# EN_VIN_BSTR_P 0.002888f
C22716 a_n3565_38502# a_n1532_35090# 1.48e-19
C22717 a_18479_47436# a_19321_45002# 0.262984f
C22718 a_7903_47542# a_2107_46812# 1.01e-20
C22719 a_11453_44696# a_12891_46348# 0.029995f
C22720 a_10227_46804# a_20843_47204# 0.02328f
C22721 a_3160_47472# a_3067_47026# 0.002863f
C22722 a_3785_47178# a_3699_46634# 0.001286f
C22723 a_584_46384# a_3055_46660# 1.4e-19
C22724 a_12465_44636# a_16119_47582# 5.64e-20
C22725 a_18597_46090# a_13747_46662# 0.391702f
C22726 a_19386_47436# a_13661_43548# 1.13e-19
C22727 a_13717_47436# a_n743_46660# 7.97e-20
C22728 a_n1435_47204# a_n2438_43548# 1.05e-19
C22729 a_n443_46116# a_n2661_46098# 0.198865f
C22730 a_n971_45724# a_5732_46660# 0.004372f
C22731 a_n237_47217# a_5167_46660# 2.88e-21
C22732 a_10729_43914# a_10518_42984# 4.92e-21
C22733 a_10405_44172# a_10835_43094# 2.45e-20
C22734 a_n2293_43922# a_n4318_37592# 0.019728f
C22735 a_n2810_45028# a_n2860_37690# 6.28e-19
C22736 a_19963_31679# a_22521_40599# 1.85e-20
C22737 a_10057_43914# a_9803_42558# 5.35e-21
C22738 a_8975_43940# a_9223_42460# 8.9e-22
C22739 a_16115_45572# VDD 0.194492f
C22740 a_18494_42460# a_19511_42282# 0.047119f
C22741 a_18184_42460# a_19647_42308# 0.034507f
C22742 a_20193_45348# a_17303_42282# 0.013391f
C22743 a_n2956_37592# a_n2302_37690# 0.04217f
C22744 a_11967_42832# a_17141_43172# 0.001676f
C22745 a_3626_43646# a_8685_43396# 8.81e-20
C22746 a_6197_43396# a_6655_43762# 0.027317f
C22747 a_2711_45572# a_14539_43914# 0.199754f
C22748 a_13059_46348# a_13565_43940# 0.011241f
C22749 a_8049_45260# a_20159_44458# 6.75e-22
C22750 a_13661_43548# a_20556_43646# 8.75e-19
C22751 a_n1613_43370# a_n1076_43230# 0.224215f
C22752 a_11322_45546# a_n2661_44458# 0.005353f
C22753 a_2324_44458# a_5013_44260# 1.86e-20
C22754 a_413_45260# a_3065_45002# 0.027891f
C22755 a_1667_45002# a_2382_45260# 3.51e-19
C22756 a_n1059_45260# a_5205_44484# 3.03e-20
C22757 a_3483_46348# a_10949_43914# 1.95e-20
C22758 a_10227_46804# a_12379_42858# 0.298444f
C22759 a_4880_45572# a_4743_44484# 7.1e-20
C22760 a_19321_45002# a_4190_30871# 6.81e-20
C22761 w_1575_34946# a_n1630_35242# 3.10971f
C22762 a_n2497_47436# a_1337_46116# 8.17e-21
C22763 a_8667_46634# a_10467_46802# 2.84e-21
C22764 a_7715_46873# a_6755_46942# 0.089466f
C22765 a_9863_46634# a_10150_46912# 0.233657f
C22766 a_8492_46660# a_10428_46928# 8.55e-21
C22767 a_11459_47204# a_10903_43370# 1.51e-21
C22768 a_n746_45260# a_739_46482# 1.28e-19
C22769 a_n1741_47186# a_n1925_42282# 3.03e-20
C22770 a_7411_46660# a_6969_46634# 0.033891f
C22771 a_6545_47178# a_2324_44458# 2.07e-20
C22772 a_13747_46662# a_19123_46287# 0.191545f
C22773 a_13661_43548# a_19551_46910# 6.46e-20
C22774 a_12549_44172# a_16655_46660# 1.26e-19
C22775 a_n881_46662# a_11415_45002# 0.017774f
C22776 a_12861_44030# a_9290_44172# 0.09212f
C22777 a_n1435_47204# a_11133_46155# 2.19e-21
C22778 a_n743_46660# a_14035_46660# 0.007691f
C22779 a_18525_43370# a_18249_42858# 0.002332f
C22780 a_15743_43084# a_18083_42858# 0.00444f
C22781 a_743_42282# a_10796_42968# 1e-19
C22782 a_15125_43396# a_5342_30871# 3.56e-20
C22783 a_n1177_43370# a_n961_42308# 1.24e-19
C22784 a_15493_43396# a_15959_42545# 8.88e-21
C22785 a_3422_30871# a_n3420_38528# 0.031237f
C22786 a_5649_42852# a_8037_42858# 2.33e-20
C22787 a_n1736_43218# a_n1545_43230# 4.61e-19
C22788 a_n4318_38680# a_n1379_43218# 1.55e-20
C22789 a_4361_42308# a_9127_43156# 2.94e-19
C22790 a_n2267_44484# VDD 0.289888f
C22791 a_n2433_43396# a_n3674_37592# 5.99e-20
C22792 a_8685_43396# a_8649_43218# 7.48e-20
C22793 a_13059_46348# a_5534_30871# 1.92e-19
C22794 a_10193_42453# a_19478_44306# 4.96e-20
C22795 a_n2293_42834# a_6298_44484# 0.002718f
C22796 a_1307_43914# a_n356_44636# 0.013327f
C22797 a_n2661_43370# a_n452_44636# 0.002717f
C22798 a_16922_45042# a_18450_45144# 0.002084f
C22799 a_4558_45348# a_n2661_42834# 8.96e-21
C22800 a_n357_42282# a_19319_43548# 1.18e-21
C22801 a_12861_44030# a_21887_42336# 2.1e-21
C22802 a_n2810_45572# a_n4318_39304# 0.023142f
C22803 a_5691_45260# a_5708_44484# 5.85e-20
C22804 a_21101_45002# a_11827_44484# 0.006993f
C22805 a_19778_44110# a_20193_45348# 0.020562f
C22806 a_18184_42460# a_11691_44458# 2.38e-19
C22807 a_4574_45260# a_n2661_43922# 9.45e-20
C22808 a_3537_45260# a_n2293_43922# 1.59e-19
C22809 a_21513_45002# a_20679_44626# 0.001342f
C22810 a_17719_45144# a_17801_45144# 0.00659f
C22811 a_n443_42852# a_8415_44056# 1.8e-19
C22812 SMPL_ON_P a_n4209_38502# 0.001002f
C22813 a_4883_46098# a_12791_45546# 8.52e-20
C22814 a_13507_46334# a_13527_45546# 0.001293f
C22815 a_n2293_46634# a_1848_45724# 0.002657f
C22816 a_768_44030# a_4099_45572# 4.61e-22
C22817 a_n743_46660# a_n1099_45572# 0.108295f
C22818 a_n1925_46634# a_n357_42282# 5.15e-20
C22819 a_8667_46634# a_8034_45724# 0.001019f
C22820 a_15227_44166# a_17715_44484# 0.385336f
C22821 a_765_45546# a_5164_46348# 6.42e-20
C22822 a_11453_44696# a_11322_45546# 0.004775f
C22823 a_12465_44636# a_12427_45724# 1.45e-19
C22824 a_12251_46660# a_10809_44734# 0.023146f
C22825 a_12816_46660# a_6945_45028# 3.52e-20
C22826 a_4190_30871# a_17531_42308# 3.05e-20
C22827 a_n2293_42282# a_n1329_42308# 4.66e-19
C22828 a_7871_42858# a_8515_42308# 2.54e-20
C22829 a_4361_42308# a_17124_42282# 0.008373f
C22830 a_19478_44306# VDD 0.127794f
C22831 a_743_42282# a_4958_30871# 0.063224f
C22832 a_8037_42858# a_7963_42308# 8.28e-20
C22833 a_n2312_39304# VDD 0.587668f
C22834 a_22612_30879# a_22821_38993# 1.98e-19
C22835 a_21588_30879# a_22469_39537# 1.05e-19
C22836 a_3537_45260# a_n97_42460# 0.74108f
C22837 a_413_45260# a_458_43396# 1.25e-20
C22838 a_n913_45002# a_n1557_42282# 0.015193f
C22839 a_4883_46098# DATA[4] 2.04e-21
C22840 a_4185_45028# a_6171_42473# 6.87e-20
C22841 a_1307_43914# a_9165_43940# 0.003526f
C22842 a_17339_46660# a_18727_42674# 8.21e-21
C22843 a_742_44458# a_2889_44172# 2.44e-20
C22844 a_13507_46334# EN_OFFSET_CAL 0.00115f
C22845 a_n699_43396# a_2127_44172# 7.77e-20
C22846 a_11453_44696# SINGLE_ENDED 0.001844f
C22847 a_n2661_43922# a_11909_44484# 2.94e-20
C22848 a_n2661_42834# a_12189_44484# 0.010003f
C22849 a_9482_43914# a_15037_43940# 1.66e-20
C22850 a_13556_45296# a_13565_43940# 4.17e-20
C22851 a_n357_42282# a_16795_42852# 0.180926f
C22852 a_12465_44636# a_14309_45028# 0.001972f
C22853 a_5066_45546# a_6633_46155# 0.001122f
C22854 a_5807_45002# a_1423_45028# 2.15e-19
C22855 a_8145_46902# a_2437_43646# 8.67e-21
C22856 a_7411_46660# a_3357_43084# 2.31e-20
C22857 a_n743_46660# a_10951_45334# 3.01e-20
C22858 a_19553_46090# a_19597_46482# 3.69e-19
C22859 a_18985_46122# a_20009_46494# 2.36e-20
C22860 a_3067_47026# a_413_45260# 0.005586f
C22861 a_15227_44166# a_15861_45028# 0.208121f
C22862 a_13507_46334# a_16922_45042# 4.88e-20
C22863 a_18597_46090# a_18911_45144# 4.8e-20
C22864 a_n443_46116# a_742_44458# 0.018829f
C22865 a_2609_46660# a_3065_45002# 4.49e-20
C22866 a_2443_46660# a_3429_45260# 2.96e-21
C22867 a_1823_45246# a_2711_45572# 0.262616f
C22868 a_10809_44734# a_13259_45724# 1.7e-19
C22869 a_n3674_37592# a_n4064_40160# 0.022617f
C22870 a_n4318_37592# a_n3420_39616# 0.020563f
C22871 a_n1630_35242# a_n4315_30879# 0.129428f
C22872 a_n3674_38216# a_n4064_39616# 0.020042f
C22873 a_n2472_42826# VDD 0.229608f
C22874 a_13076_44458# a_9145_43396# 1.6e-19
C22875 a_n755_45592# a_7174_31319# 2.56e-20
C22876 a_n357_42282# a_21335_42336# 2.03e-19
C22877 a_n913_45002# a_8483_43230# 2.14e-19
C22878 a_n1059_45260# a_3863_42891# 4.31e-19
C22879 a_1307_43914# a_12379_42858# 2.23e-20
C22880 a_10193_42453# a_9223_42460# 6.94e-19
C22881 a_n2810_45572# a_n4334_40480# 5.22e-19
C22882 a_11967_42832# a_18797_44260# 3.24e-19
C22883 a_n2661_42834# a_1756_43548# 9.68e-20
C22884 a_n2661_43922# a_1568_43370# 4.28e-22
C22885 a_n356_44636# a_9396_43370# 1.18e-20
C22886 a_18280_46660# START 1.24e-19
C22887 a_7499_43078# a_9885_42558# 0.020607f
C22888 a_13556_45296# a_5534_30871# 1.32e-21
C22889 a_18184_42460# a_4190_30871# 0.630738f
C22890 a_n2293_42834# a_n967_43230# 7.58e-20
C22891 a_2324_44458# a_4927_45028# 3.2e-20
C22892 a_5257_43370# a_6109_44484# 0.001517f
C22893 a_3090_45724# a_4743_44484# 0.05313f
C22894 a_n881_46662# a_n984_44318# 8.92e-19
C22895 a_n1613_43370# a_175_44278# 2.35e-19
C22896 a_11189_46129# a_10951_45334# 4.23e-21
C22897 a_9290_44172# a_11787_45002# 4.62e-19
C22898 a_2711_45572# a_12427_45724# 0.014959f
C22899 a_14275_46494# a_6171_45002# 1.21e-20
C22900 a_4808_45572# a_4880_45572# 0.003395f
C22901 a_21137_46414# a_413_45260# 4e-22
C22902 a_8049_45260# a_20623_45572# 0.01128f
C22903 a_19123_46287# a_18911_45144# 7.75e-20
C22904 a_13059_46348# a_11691_44458# 0.015799f
C22905 a_13259_45724# a_16211_45572# 0.004313f
C22906 a_8953_45546# a_9482_43914# 1.61e-19
C22907 a_n746_45260# a_1241_43940# 4.29e-20
C22908 a_n746_45260# a_768_44030# 0.005354f
C22909 a_2952_47436# a_n1613_43370# 2.81e-19
C22910 a_2905_45572# a_3411_47243# 0.005614f
C22911 a_n1151_42308# a_5063_47570# 1.74e-19
C22912 a_n3565_39590# a_n3690_37440# 1.95e-19
C22913 a_11599_46634# a_18597_46090# 0.191253f
C22914 a_16241_47178# a_10227_46804# 0.022072f
C22915 a_16327_47482# a_17591_47464# 0.339529f
C22916 a_16023_47582# a_16588_47582# 7.99e-20
C22917 a_11459_47204# a_4883_46098# 2.08e-20
C22918 a_21335_42336# CAL_N 9.12e-19
C22919 a_1736_39587# VDAC_Ni 5.68e-19
C22920 a_n4209_39590# a_n2946_37690# 1.64e-19
C22921 a_15673_47210# a_18143_47464# 3.18e-20
C22922 a_5742_30871# C3_N_btm 0.030866f
C22923 a_n1435_47204# a_13507_46334# 1.53e-21
C22924 a_13717_47436# a_21177_47436# 6.95e-20
C22925 a_9223_42460# VDD 0.205797f
C22926 a_n3420_38528# a_n3607_38304# 6.01e-19
C22927 a_n3420_39616# a_n4334_37440# 4.91e-19
C22928 a_1736_39043# VDAC_Pi 0.001304f
C22929 a_11967_42832# a_15567_42826# 0.067391f
C22930 a_5891_43370# a_8495_42852# 3.14e-20
C22931 a_n97_42460# a_1049_43396# 0.195034f
C22932 a_14401_32519# a_2982_43646# 4.51e-20
C22933 a_17973_43940# a_17499_43370# 0.018568f
C22934 a_17737_43940# a_17324_43396# 0.001548f
C22935 a_n2956_37592# a_n2946_39072# 2.49e-19
C22936 a_6511_45714# VDD 0.405279f
C22937 a_n4318_40392# a_n1630_35242# 1.96e-19
C22938 a_14021_43940# a_14579_43548# 1.31e-19
C22939 a_15493_43396# a_16243_43396# 0.041358f
C22940 a_584_46384# a_685_42968# 0.00804f
C22941 a_11453_44696# a_16409_43396# 8.34e-21
C22942 a_13507_46334# a_15743_43084# 0.158635f
C22943 a_20107_45572# a_19963_31679# 3.1e-20
C22944 a_21188_45572# a_2437_43646# 0.00191f
C22945 a_12861_44030# a_13467_32519# 9.12e-21
C22946 a_12891_46348# a_9145_43396# 0.001541f
C22947 a_19466_46812# a_20269_44172# 2.46e-20
C22948 a_16327_47482# a_17678_43396# 0.001965f
C22949 a_20273_45572# a_22591_45572# 4.71e-20
C22950 a_20841_45814# a_3357_43084# 0.047766f
C22951 a_15765_45572# a_6171_45002# 0.001099f
C22952 a_10809_44734# a_n2661_43922# 0.073946f
C22953 a_2711_45572# a_14309_45028# 0.028068f
C22954 a_14275_46494# a_14673_44172# 3.31e-21
C22955 a_19692_46634# a_19862_44208# 0.027038f
C22956 a_11599_46634# a_19123_46287# 0.024241f
C22957 a_15673_47210# a_765_45546# 0.028544f
C22958 a_n2661_46098# a_1302_46660# 2.6e-19
C22959 a_n2497_47436# a_3699_46348# 6.3e-22
C22960 a_n2109_47186# a_3147_46376# 5.93e-20
C22961 a_n1741_47186# a_2698_46116# 9.05e-21
C22962 a_n1386_35608# VIN_P 0.367112f
C22963 C8_P_btm VDD 0.19922f
C22964 a_13507_46334# a_13885_46660# 5.84e-20
C22965 a_15811_47375# a_17829_46910# 2.1e-20
C22966 a_2107_46812# a_4817_46660# 0.002361f
C22967 a_2609_46660# a_3067_47026# 0.027317f
C22968 a_2959_46660# a_3524_46660# 7.99e-20
C22969 a_n1925_46634# a_5263_46660# 8.56e-19
C22970 C0_dummy_N_btm C2_N_btm 6.66125f
C22971 C0_N_btm C1_N_btm 10.8764f
C22972 C0_dummy_P_btm C3_N_btm 2.71e-19
C22973 C3_P_btm C7_N_btm 6.36e-19
C22974 C1_P_btm C5_N_btm 1.59e-19
C22975 C0_P_btm C4_N_btm 1.4e-19
C22976 a_13717_47436# a_20841_46902# 1.67e-20
C22977 a_n746_45260# a_1176_45822# 3.33e-20
C22978 a_n237_47217# a_1208_46090# 0.003284f
C22979 a_327_47204# a_376_46348# 1.5e-19
C22980 a_n971_45724# a_1138_42852# 1.34e-20
C22981 a_13747_46662# a_6755_46942# 0.316914f
C22982 a_n2661_46634# a_8145_46902# 0.008097f
C22983 a_18579_44172# a_18727_42674# 4.15e-22
C22984 a_117_45144# VDD 2.04e-19
C22985 a_8685_43396# a_8037_42858# 0.001875f
C22986 a_3626_43646# a_17333_42852# 2.21e-20
C22987 a_2982_43646# a_18817_42826# 3.67e-20
C22988 a_15743_43084# a_21855_43396# 0.001426f
C22989 a_19268_43646# a_4361_42308# 4.9e-21
C22990 a_8488_45348# a_8560_45348# 0.003395f
C22991 a_5937_45572# a_6293_42852# 1.17e-19
C22992 a_3775_45552# a_3600_43914# 9.84e-21
C22993 a_3065_45002# a_2779_44458# 0.001276f
C22994 w_11334_34010# a_4958_30871# 0.003841f
C22995 a_2324_44458# a_4699_43561# 1.33e-20
C22996 a_13556_45296# a_11691_44458# 0.399095f
C22997 a_14797_45144# a_11827_44484# 5.28e-21
C22998 a_5837_45028# a_n2661_43370# 0.005758f
C22999 a_6431_45366# a_n2661_44458# 7.71e-21
C23000 a_2382_45260# a_n699_43396# 0.075387f
C23001 SMPL_ON_N a_n1630_35242# 0.076872f
C23002 a_8696_44636# a_12553_44484# 8.86e-20
C23003 a_n2438_43548# a_526_44458# 0.107408f
C23004 a_n743_46660# a_n1925_42282# 0.010043f
C23005 a_13747_46662# a_8049_45260# 0.208778f
C23006 a_16388_46812# a_765_45546# 0.164902f
C23007 a_16721_46634# a_17339_46660# 0.005637f
C23008 a_12549_44172# a_12638_46436# 3.01e-19
C23009 a_12891_46348# a_14180_46482# 1.22e-21
C23010 a_8667_46634# a_8016_46348# 1.13e-19
C23011 a_7577_46660# a_5937_45572# 2.93e-19
C23012 a_7927_46660# a_8349_46414# 0.01072f
C23013 a_6151_47436# a_6598_45938# 0.173467f
C23014 a_6545_47178# a_6667_45809# 1.61e-19
C23015 a_6851_47204# a_6472_45840# 5.75e-21
C23016 a_6491_46660# a_6511_45714# 5.95e-22
C23017 a_n881_46662# a_13259_45724# 0.507296f
C23018 a_3877_44458# a_2324_44458# 0.153319f
C23019 a_5807_45002# a_9823_46482# 2.88e-19
C23020 a_15227_44166# a_22365_46825# 3.68e-20
C23021 a_17609_46634# a_11415_45002# 5.34e-21
C23022 a_12281_43396# a_12563_42308# 0.173003f
C23023 a_4361_42308# a_1755_42282# 0.015476f
C23024 a_n1641_43230# COMP_P 8.01e-19
C23025 a_n1423_42826# a_n1329_42308# 0.001077f
C23026 a_15095_43370# a_14113_42308# 6.79e-20
C23027 a_2982_43646# a_21421_42336# 9.11e-19
C23028 a_3626_43646# a_18997_42308# 8.14e-19
C23029 a_n2065_43946# VDD 0.4213f
C23030 a_n1991_42858# a_n961_42308# 0.001344f
C23031 a_12379_42858# a_13003_42852# 9.73e-19
C23032 a_n4318_38680# a_n4318_38216# 0.055776f
C23033 a_12895_43230# a_13157_43218# 0.001705f
C23034 a_12545_42858# a_13569_43230# 2.36e-20
C23035 a_3422_30871# VIN_N 0.057975f
C23036 a_n4318_39304# a_n4251_39392# 3.13e-19
C23037 a_8746_45002# a_10695_43548# 3.62e-21
C23038 a_10193_42453# a_13667_43396# 5.44e-20
C23039 a_3357_43084# a_5829_43940# 0.00562f
C23040 a_21359_45002# a_19279_43940# 8.47e-19
C23041 a_11827_44484# a_20766_44850# 0.004974f
C23042 a_2711_45572# a_17324_43396# 7.1e-20
C23043 a_1209_47178# VDD 0.38145f
C23044 a_5883_43914# a_n2661_43922# 0.028328f
C23045 a_10440_44484# a_10617_44484# 0.134298f
C23046 a_11963_45334# a_10949_43914# 1.06e-20
C23047 a_5009_45028# a_3905_42865# 1.03e-19
C23048 a_9482_43914# a_9028_43914# 0.092045f
C23049 a_n443_42852# a_15868_43402# 3.07e-19
C23050 a_11322_45546# a_9145_43396# 4.56e-21
C23051 a_n2312_38680# a_n3420_38528# 0.009774f
C23052 a_n2293_42834# a_2479_44172# 0.021799f
C23053 a_n2661_43370# a_n809_44244# 5.6e-20
C23054 a_20193_45348# a_20159_44458# 5.71e-19
C23055 w_11334_34010# VCM 0.001153f
C23056 a_626_44172# a_1525_44260# 2.9e-21
C23057 a_n2661_45010# a_2455_43940# 3.99e-19
C23058 a_n2293_45010# a_1443_43940# 3.99e-19
C23059 a_n971_45724# DATA[1] 0.050116f
C23060 a_n746_45260# DATA[0] 0.03466f
C23061 a_8199_44636# a_5066_45546# 0.178583f
C23062 a_12549_44172# a_n2017_45002# 5.58e-20
C23063 a_n881_46662# a_n467_45028# 0.008624f
C23064 a_n1613_43370# a_n143_45144# 4.99e-21
C23065 a_3094_47243# a_413_45260# 5.44e-19
C23066 a_13059_46348# a_n443_42852# 0.09278f
C23067 a_13661_43548# a_3357_43084# 2.72e-20
C23068 a_13747_46662# a_19479_31679# 8.06e-20
C23069 a_18819_46122# a_6945_45028# 4.66e-20
C23070 a_19335_46494# a_19900_46494# 7.99e-20
C23071 a_18985_46122# a_21137_46414# 5.31e-20
C23072 a_18189_46348# a_10809_44734# 8.9e-20
C23073 a_10227_46804# a_14180_45002# 0.002579f
C23074 a_19321_45002# a_2437_43646# 0.009654f
C23075 a_3090_45724# a_4808_45572# 2.21e-19
C23076 a_2063_45854# a_n2661_43370# 0.039988f
C23077 a_961_42354# a_5934_30871# 1.72e-20
C23078 a_5342_30871# a_n4064_38528# 0.028644f
C23079 a_3318_42354# a_4921_42308# 1.41e-19
C23080 a_1755_42282# a_6761_42308# 0.008867f
C23081 a_1606_42308# a_7227_42308# 3.31e-20
C23082 a_13667_43396# VDD 0.402378f
C23083 a_13678_32519# VDAC_N 3.33e-19
C23084 a_n784_42308# a_9223_42460# 1.96e-20
C23085 a_16328_43172# a_4958_30871# 1.29e-20
C23086 a_n755_45592# a_5932_42308# 0.040158f
C23087 a_n2661_43922# a_12495_44260# 2.04e-19
C23088 a_n2661_42834# a_12603_44260# 6.24e-19
C23089 a_1414_42308# a_453_43940# 0.248504f
C23090 a_644_44056# a_895_43940# 0.106452f
C23091 a_1115_44172# a_2479_44172# 9.15e-20
C23092 a_n2956_38680# a_n4209_39590# 0.020934f
C23093 a_18989_43940# a_18797_44260# 9.07e-19
C23094 a_n913_45002# a_3935_42891# 5.11e-21
C23095 a_n1059_45260# a_4520_42826# 0.004119f
C23096 a_n2017_45002# a_5111_42852# 1.11e-19
C23097 a_13259_45724# a_13333_42558# 8.98e-20
C23098 a_10768_47026# VDD 0.132317f
C23099 a_742_44458# a_1049_43396# 2.13e-19
C23100 a_949_44458# a_1209_43370# 6.32e-19
C23101 a_n755_45592# a_2307_45899# 9.75e-21
C23102 a_584_46384# a_3600_43914# 3.17e-19
C23103 a_18479_47436# a_20362_44736# 1.52e-20
C23104 a_16327_47482# a_18245_44484# 3.03e-19
C23105 a_380_45546# a_603_45572# 0.011458f
C23106 a_n1099_45572# a_509_45572# 0.001017f
C23107 a_11601_46155# a_10193_42453# 0.002905f
C23108 a_5807_45002# a_6109_44484# 3.89e-20
C23109 a_n2293_46098# a_n143_45144# 2.2e-21
C23110 a_5068_46348# a_2437_43646# 1.07e-20
C23111 a_n881_46662# a_n2661_43922# 4.12e-19
C23112 a_4185_45028# a_3357_43084# 0.027077f
C23113 a_n1613_43370# a_n2293_43922# 2.76e-19
C23114 a_5066_45546# a_8192_45572# 0.001238f
C23115 a_n2661_45546# a_5263_45724# 6.45e-19
C23116 a_n2293_46634# a_n2012_44484# 8.23e-19
C23117 a_10809_44734# a_17478_45572# 1.1e-21
C23118 a_1138_42852# a_n2293_45010# 9.98e-19
C23119 a_15682_46116# a_16147_45260# 2.64e-19
C23120 a_n4209_39590# a_n3690_39392# 2.69e-19
C23121 a_n4064_39616# a_n4251_39616# 0.001131f
C23122 a_6123_31319# VDAC_N 0.006984f
C23123 a_n784_42308# C8_P_btm 6.79e-20
C23124 a_1606_42308# a_n923_35174# 0.002555f
C23125 a_n1741_47186# a_n1435_47204# 0.047534f
C23126 a_2553_47502# a_n443_46116# 1.33e-19
C23127 a_3381_47502# a_3785_47178# 0.00589f
C23128 a_n1151_42308# a_3815_47204# 0.01223f
C23129 a_n237_47217# a_6575_47204# 0.0275f
C23130 a_2063_45854# a_4915_47217# 0.055521f
C23131 a_2905_45572# a_4700_47436# 4.48e-20
C23132 a_n3690_39616# a_n4209_39304# 2.69e-19
C23133 a_4958_30871# a_n4064_37984# 0.030919f
C23134 a_20256_43172# VDD 7.47e-19
C23135 a_n1630_35242# a_19864_35138# 0.020191f
C23136 en_comp a_15486_42560# 1.51e-21
C23137 a_n356_44636# a_13635_43156# 9.74e-20
C23138 a_1307_43914# a_3823_42558# 6.3e-20
C23139 a_n2293_42834# a_n2104_42282# 0.004809f
C23140 a_n913_45002# a_15890_42674# 1.94e-19
C23141 a_5891_43370# a_9127_43156# 0.457718f
C23142 a_17970_44736# a_18083_42858# 5.77e-21
C23143 a_20159_44458# a_20301_43646# 3.21e-20
C23144 a_20640_44752# a_21259_43561# 6.9e-19
C23145 a_14539_43914# a_18817_42826# 5.94e-20
C23146 a_11387_46482# DATA[5] 5.29e-20
C23147 a_n2661_42282# a_7112_43396# 1.53e-19
C23148 a_11601_46155# VDD 0.001563f
C23149 a_13661_43548# a_18533_44260# 7.69e-20
C23150 a_13759_46122# a_13720_44458# 1.69e-22
C23151 a_n443_42852# a_13556_45296# 2.5e-20
C23152 a_12549_44172# a_21845_43940# 0.003853f
C23153 a_2711_45572# a_6709_45028# 0.002223f
C23154 a_8049_45260# a_18911_45144# 1.78e-20
C23155 a_n1613_43370# a_n97_42460# 0.011527f
C23156 a_5907_45546# a_6431_45366# 9.96e-19
C23157 a_6194_45824# a_6171_45002# 0.006466f
C23158 a_6472_45840# a_3232_43370# 0.001072f
C23159 a_3483_46348# a_7640_43914# 0.003497f
C23160 a_3503_45724# a_1307_43914# 1.08e-21
C23161 a_n755_45592# a_1423_45028# 0.032517f
C23162 a_5263_45724# a_5205_44484# 4.99e-21
C23163 a_n2312_39304# a_3080_42308# 4.02e-21
C23164 a_3090_45724# a_1414_42308# 8.03e-21
C23165 a_6229_45572# a_3357_43084# 6.33e-19
C23166 a_8270_45546# a_7542_44172# 4.69e-19
C23167 a_16855_45546# a_18175_45572# 2.91e-21
C23168 a_16680_45572# a_16147_45260# 2.09e-19
C23169 a_12741_44636# a_15146_44811# 1.05e-19
C23170 a_n2293_46098# a_n2293_43922# 7.21e-22
C23171 a_n3420_37440# C5_P_btm 1.87e-19
C23172 a_n4209_37414# C1_P_btm 0.043983f
C23173 a_n4064_37440# C7_P_btm 1.83e-20
C23174 a_11599_46634# a_6755_46942# 0.321942f
C23175 a_20916_46384# a_21588_30879# 5.25e-19
C23176 a_13661_43548# a_n2293_46634# 0.055067f
C23177 a_n881_46662# a_1799_45572# 0.028083f
C23178 a_6151_47436# a_11735_46660# 1.81e-19
C23179 a_6575_47204# a_8270_45546# 9.19e-20
C23180 a_4915_47217# a_12469_46902# 5.76e-19
C23181 a_n1151_42308# a_14976_45028# 1.72e-19
C23182 a_n1613_43370# a_n2661_46098# 1.40554f
C23183 a_n4064_37984# VCM 0.011087f
C23184 a_4883_46098# a_5072_46660# 7.49e-20
C23185 a_22545_38993# a_22876_39857# 4.42e-19
C23186 a_22459_39145# a_22705_38406# 6.64e-21
C23187 a_22521_40599# a_22717_36887# 1.4e-19
C23188 a_22469_40625# a_22717_37285# 0.002464f
C23189 a_22521_40055# a_22609_37990# 0.234448f
C23190 a_22521_39511# CAL_P 0.027034f
C23191 a_19963_31679# VIN_N 0.029022f
C23192 a_19479_31679# VCM 0.03628f
C23193 a_n1761_44111# a_196_42282# 2.46e-19
C23194 a_n356_44636# a_18310_42308# 5.53e-19
C23195 a_n2810_45028# VDD 0.526631f
C23196 a_n1655_43396# a_n4318_38680# 7.29e-20
C23197 a_14955_43396# a_15681_43442# 9.54e-19
C23198 a_14021_43940# a_21671_42860# 6.16e-20
C23199 a_6431_45366# a_6125_45348# 7.37e-20
C23200 a_6171_45002# a_6517_45366# 6.95e-19
C23201 a_n357_42282# a_3422_30871# 0.122733f
C23202 a_20623_45572# a_20193_45348# 4.8e-19
C23203 a_12549_44172# a_19164_43230# 1.3e-20
C23204 a_15227_44166# a_15095_43370# 0.022423f
C23205 a_3090_45724# a_12281_43396# 0.027472f
C23206 a_14537_43396# a_16019_45002# 5.14e-20
C23207 a_n2293_46098# a_n97_42460# 0.333817f
C23208 a_8696_44636# a_10157_44484# 0.004815f
C23209 a_10227_46804# a_12800_43218# 2.53e-19
C23210 a_n1151_42308# a_n4318_38216# 9.61e-21
C23211 a_8162_45546# a_n2661_43922# 3.6e-21
C23212 a_4558_45348# a_5093_45028# 0.001257f
C23213 a_5147_45002# a_5009_45028# 0.007368f
C23214 a_9049_44484# a_9159_44484# 0.031707f
C23215 a_n2293_46634# a_10835_43094# 8.49e-20
C23216 a_21513_45002# a_18494_42460# 8.98e-20
C23217 a_n955_45028# a_n2661_43370# 6.51e-19
C23218 a_6755_46942# a_13693_46688# 0.001956f
C23219 a_15009_46634# a_3090_45724# 0.154981f
C23220 a_12549_44172# a_13759_46122# 5.27e-19
C23221 a_12891_46348# a_13925_46122# 2.71e-21
C23222 a_n2293_46634# a_4185_45028# 0.027799f
C23223 a_8128_46384# a_2324_44458# 2.07e-20
C23224 a_8145_46902# a_765_45546# 1.38e-20
C23225 a_n881_46662# a_18189_46348# 2.07e-20
C23226 a_11599_46634# a_8049_45260# 0.14064f
C23227 a_n2497_47436# a_n755_45592# 0.45034f
C23228 a_768_44030# a_13351_46090# 1.3e-19
C23229 a_n743_46660# a_2698_46116# 0.013101f
C23230 a_n2438_43548# a_2521_46116# 5.14e-19
C23231 a_1123_46634# a_1208_46090# 0.0037f
C23232 a_n133_46660# a_167_45260# 5.4e-22
C23233 a_2107_46812# a_472_46348# 2.45e-19
C23234 a_n237_47217# a_n2661_45546# 0.038356f
C23235 a_4915_47217# a_14383_46116# 9.48e-19
C23236 a_n2661_46634# a_5068_46348# 3.78e-20
C23237 a_n815_47178# a_n1079_45724# 7.01e-21
C23238 a_n971_45724# a_n2956_38216# 1.71e-19
C23239 a_n2661_46098# a_n2293_46098# 0.063852f
C23240 a_n1925_46634# a_3147_46376# 1.66e-19
C23241 a_5807_45002# a_9569_46155# 2.47e-19
C23242 a_n1435_47204# a_10586_45546# 4.56e-21
C23243 a_2982_43646# a_5934_30871# 0.178f
C23244 a_3422_30871# CAL_N 0.236929f
C23245 a_n97_42460# a_13249_42558# 5.74e-19
C23246 a_3626_43646# a_6123_31319# 0.109715f
C23247 a_12545_42858# a_13113_42826# 0.178024f
C23248 a_12379_42858# a_13635_43156# 0.043475f
C23249 a_12089_42308# a_12895_43230# 4.25e-19
C23250 a_5891_43370# CLK 8.38e-19
C23251 a_n2661_43370# a_n2661_42834# 0.306215f
C23252 a_413_45260# a_2479_44172# 0.008619f
C23253 a_n2472_45002# a_n3674_39768# 1.13e-19
C23254 a_n2293_45010# a_n4318_39768# 1.61e-21
C23255 a_n2661_45010# a_n1644_44306# 7.26e-19
C23256 a_2437_43646# a_2537_44260# 7.55e-20
C23257 a_2324_44458# a_1847_42826# 3.13e-21
C23258 a_9290_44172# a_9127_43156# 0.003077f
C23259 a_n443_42852# a_6293_42852# 0.033407f
C23260 a_n2312_39304# a_n2946_39072# 0.020842f
C23261 a_n2017_45002# a_7542_44172# 2.92e-21
C23262 a_n1925_42282# a_4361_42308# 0.08654f
C23263 a_8953_45546# a_10796_42968# 2.18e-20
C23264 a_4185_45028# a_5342_30871# 0.067871f
C23265 a_18479_45785# a_19478_44306# 0.005615f
C23266 a_4223_44672# a_5518_44484# 0.003606f
C23267 a_n699_43396# a_5343_44458# 9.51e-20
C23268 a_13661_43548# a_20107_42308# 3.89e-19
C23269 a_2274_45254# a_1414_42308# 1.01e-20
C23270 a_18597_46090# a_20841_45814# 0.024341f
C23271 a_n743_46660# a_13527_45546# 8.32e-20
C23272 a_5732_46660# a_2711_45572# 2.43e-20
C23273 a_2063_45854# a_4574_45260# 6.45e-20
C23274 a_n443_46116# a_n467_45028# 1.81e-19
C23275 a_4007_47204# a_413_45260# 4.35e-19
C23276 a_n881_46662# a_17478_45572# 0.11503f
C23277 a_18479_47436# a_21363_45546# 0.001869f
C23278 a_16327_47482# a_20719_45572# 0.001951f
C23279 a_4646_46812# a_6511_45714# 0.421269f
C23280 a_3877_44458# a_6667_45809# 7.89e-19
C23281 a_3483_46348# a_9823_46155# 2.75e-19
C23282 a_n237_47217# a_5205_44484# 1.8e-20
C23283 a_n971_45724# a_7229_43940# 7.24e-21
C23284 a_17609_46634# a_13259_45724# 9.09e-19
C23285 a_2905_45572# a_3065_45002# 0.004116f
C23286 a_11415_45002# a_22223_46124# 0.011454f
C23287 a_20202_43084# a_10809_44734# 0.014133f
C23288 a_584_46384# a_4558_45348# 2.74e-19
C23289 a_15811_47375# a_2437_43646# 0.006582f
C23290 a_14955_47212# a_3357_43084# 2.77e-19
C23291 a_3080_42308# C8_P_btm 0.006767f
C23292 a_n2840_42282# a_n4318_38216# 0.015074f
C23293 a_n2129_43609# VDD 0.400674f
C23294 a_17701_42308# a_16522_42674# 7.63e-21
C23295 a_n3674_38680# a_n2472_42282# 5e-19
C23296 a_n2293_42834# a_n229_43646# 0.001042f
C23297 a_1307_43914# a_6765_43638# 2.03e-20
C23298 a_19615_44636# a_19789_44512# 0.006584f
C23299 a_11967_42832# a_20980_44850# 8.49e-19
C23300 a_10193_42453# a_21195_42852# 0.005652f
C23301 a_3232_43370# a_10695_43548# 4.03e-21
C23302 a_14539_43914# a_15682_43940# 0.161926f
C23303 a_17517_44484# a_17730_32519# 0.00864f
C23304 a_n2661_43922# a_2889_44172# 0.001413f
C23305 a_n2661_42834# a_2998_44172# 0.790177f
C23306 a_526_44458# a_7227_42308# 5.53e-20
C23307 a_2324_44458# a_15486_42560# 5.07e-20
C23308 a_383_46660# DATA[0] 2.11e-19
C23309 a_n2661_43370# a_n1352_43396# 3.84e-21
C23310 a_5708_44484# a_5013_44260# 3.54e-19
C23311 a_3537_45260# a_9885_43646# 2e-19
C23312 a_4185_45028# a_20107_42308# 1.64e-19
C23313 a_288_46660# VDD 0.079457f
C23314 a_n357_42282# a_18504_43218# 0.003243f
C23315 a_n1059_45260# a_16409_43396# 4.57e-19
C23316 a_n913_45002# a_16547_43609# 4.63e-21
C23317 a_n2017_45002# a_16977_43638# 6.48e-21
C23318 a_20679_44626# a_18579_44172# 1.41e-20
C23319 a_20107_46660# a_20107_45572# 0.001171f
C23320 a_13059_46348# a_2437_43646# 7.82e-20
C23321 a_11453_44696# a_12883_44458# 1.4e-20
C23322 a_2324_44458# a_10053_45546# 0.008381f
C23323 a_5937_45572# a_6905_45572# 9.25e-20
C23324 a_11309_47204# a_n2661_44458# 1.64e-20
C23325 a_15368_46634# a_413_45260# 4.42e-20
C23326 a_12594_46348# a_11962_45724# 0.177228f
C23327 a_19321_45002# a_19113_45348# 0.147788f
C23328 a_13661_43548# a_16237_45028# 5.58e-19
C23329 a_13747_46662# a_20193_45348# 0.049365f
C23330 a_n443_46116# a_n2661_43922# 0.044169f
C23331 a_4791_45118# a_n2293_43922# 3.57e-19
C23332 a_12005_46116# a_12427_45724# 0.01091f
C23333 a_10903_43370# a_11823_42460# 1.16382f
C23334 a_n743_46660# a_16922_45042# 2.99e-19
C23335 a_5932_42308# a_n3420_38528# 0.001859f
C23336 a_17303_42282# a_19647_42308# 3.68e-19
C23337 a_4958_30871# a_13258_32519# 0.033151f
C23338 a_5342_30871# VREF_GND 0.055227f
C23339 a_21195_42852# VDD 0.285496f
C23340 a_18057_42282# a_18548_42308# 0.00278f
C23341 a_5742_30871# a_1736_39587# 7.65e-20
C23342 a_21356_42826# RST_Z 4.49e-21
C23343 a_2675_43914# a_n97_42460# 1.83e-19
C23344 a_9290_44172# CLK 0.151406f
C23345 a_11341_43940# a_11173_44260# 0.049235f
C23346 a_644_44056# a_458_43396# 2.18e-19
C23347 a_20512_43084# a_2982_43646# 0.029475f
C23348 a_9313_44734# a_17499_43370# 2.25e-19
C23349 a_n2017_45002# a_n1630_35242# 0.111641f
C23350 a_15015_46420# VDD 0.337162f
C23351 a_n967_45348# a_n961_42308# 0.174237f
C23352 a_n1059_45260# a_564_42282# 0.043244f
C23353 a_n913_45002# a_n3674_37592# 8.1e-20
C23354 a_19478_44306# a_14021_43940# 5.41e-20
C23355 a_n2293_42834# a_1793_42852# 1.98e-35
C23356 a_n2661_44458# a_3935_42891# 5.85e-22
C23357 a_11133_46155# DATA[5] 2.67e-20
C23358 a_10586_45546# a_10775_45002# 1.57e-19
C23359 a_4791_45118# a_n97_42460# 0.02536f
C23360 a_12861_44030# a_19319_43548# 0.024237f
C23361 a_584_46384# a_1756_43548# 0.00975f
C23362 a_n1076_46494# a_n2129_44697# 2.07e-21
C23363 a_10193_42453# a_16333_45814# 7.72e-20
C23364 a_2324_44458# a_13490_45394# 6.46e-19
C23365 a_11823_42460# a_12016_45572# 1.71e-19
C23366 a_n1991_46122# a_n1177_44458# 9.68e-22
C23367 a_7499_43078# a_8696_44636# 0.155392f
C23368 a_n2661_45546# a_n2017_45002# 0.001101f
C23369 a_10210_45822# a_10907_45822# 0.013775f
C23370 a_n1079_45724# a_n2661_45010# 5.36e-21
C23371 a_n2293_45546# a_n2472_45002# 3.35e-19
C23372 a_20205_31679# en_comp 1.91e-19
C23373 a_12549_44172# a_18079_43940# 0.008672f
C23374 a_8049_45260# a_13348_45260# 7.18e-21
C23375 a_n2302_40160# VDD 0.428934f
C23376 a_2747_46873# a_n881_46662# 5.46e-20
C23377 a_7754_40130# a_5700_37509# 0.037095f
C23378 a_7754_39964# a_4338_37500# 0.021449f
C23379 a_18780_47178# a_13747_46662# 0.028845f
C23380 a_18479_47436# a_19452_47524# 5.84e-19
C23381 a_7754_38636# a_7754_38470# 0.296258f
C23382 VDAC_Pi a_3726_37500# 1.17174f
C23383 a_11453_44696# a_11309_47204# 2.71e-19
C23384 a_10227_46804# a_19594_46812# 0.01518f
C23385 a_18143_47464# a_19321_45002# 2.46e-20
C23386 a_16588_47582# a_16750_47204# 0.006453f
C23387 a_n1151_42308# a_3524_46660# 4.19e-20
C23388 a_2905_45572# a_3067_47026# 1.43e-19
C23389 a_n3565_39304# C5_P_btm 3.17e-19
C23390 a_n3420_39072# C7_P_btm 9.48e-19
C23391 a_n4064_39072# C9_P_btm 7.29e-20
C23392 a_12465_44636# a_15928_47570# 5.23e-20
C23393 a_13258_32519# VCM 0.033198f
C23394 a_7174_31319# VIN_N 0.022822f
C23395 a_n1435_47204# a_n743_46660# 2.75e-20
C23396 a_n443_46116# a_1799_45572# 0.081828f
C23397 a_n2109_47186# a_5894_47026# 1.64e-19
C23398 a_n971_45724# a_5907_46634# 3.23e-19
C23399 a_n3565_38502# a_n1386_35608# 1.73e-19
C23400 a_18597_46090# a_13661_43548# 0.266647f
C23401 a_19386_47436# a_5807_45002# 2.36e-21
C23402 a_n2956_37592# a_n4064_37440# 0.070596f
C23403 a_11064_45572# CLK 6.18e-19
C23404 a_10729_43914# a_10083_42826# 5.47e-19
C23405 a_10405_44172# a_10518_42984# 2.78e-20
C23406 a_5891_43370# a_1755_42282# 3.89e-20
C23407 a_n2810_45028# a_n2302_37690# 0.162246f
C23408 a_19319_43548# a_19700_43370# 0.006809f
C23409 a_n2293_43922# a_n1736_42282# 4.89e-19
C23410 a_16333_45814# VDD 0.201203f
C23411 a_11967_42832# a_16877_43172# 0.003239f
C23412 a_19778_44110# a_19647_42308# 2.28e-21
C23413 a_18184_42460# a_19511_42282# 0.058931f
C23414 a_18494_42460# a_18548_42308# 0.005603f
C23415 a_6197_43396# a_6452_43396# 0.06121f
C23416 a_7287_43370# a_8147_43396# 2.55e-19
C23417 a_10227_46804# a_10341_42308# 0.004877f
C23418 a_2711_45572# a_16112_44458# 0.183744f
C23419 a_10490_45724# a_n2661_44458# 2.68e-21
C23420 a_n913_45002# a_6171_45002# 8.52e-21
C23421 a_13661_43548# a_743_42282# 0.132115f
C23422 a_n1613_43370# a_n901_43156# 0.281398f
C23423 a_413_45260# a_2680_45002# 0.01804f
C23424 a_n2017_45002# a_5205_44484# 2.49e-20
C23425 a_3483_46348# a_10729_43914# 1.6e-21
C23426 a_n357_42282# a_7640_43914# 8.82e-19
C23427 a_2324_44458# a_5244_44056# 1.7e-20
C23428 a_8492_46660# a_10150_46912# 0.00213f
C23429 a_8667_46634# a_10428_46928# 6.23e-20
C23430 a_11459_47204# a_11387_46155# 1.29e-20
C23431 a_n746_45260# a_518_46482# 7.09e-19
C23432 a_n1741_47186# a_526_44458# 3.03e-20
C23433 a_2063_45854# a_10809_44734# 0.169005f
C23434 a_7411_46660# a_6755_46942# 0.265786f
C23435 a_5257_43370# a_6969_46634# 6.29e-21
C23436 a_6151_47436# a_2324_44458# 0.002957f
C23437 a_13747_46662# a_18285_46348# 1.64e-19
C23438 a_n2661_46634# a_13059_46348# 1.84e-19
C23439 a_13661_43548# a_19123_46287# 0.073049f
C23440 a_5807_45002# a_19551_46910# 1.7e-20
C23441 a_12549_44172# a_16434_46660# 2.11e-19
C23442 a_n1435_47204# a_11189_46129# 9.06e-22
C23443 a_2959_46660# a_3090_45724# 4.18e-19
C23444 a_n743_46660# a_13885_46660# 1.96e-21
C23445 a_18597_46090# a_4185_45028# 1.12e-19
C23446 a_18783_43370# a_18083_42858# 9.54e-20
C23447 a_15743_43084# a_17701_42308# 1.11e-19
C23448 a_18429_43548# a_18249_42858# 0.001117f
C23449 a_743_42282# a_10835_43094# 8.66e-20
C23450 a_15037_43396# a_5342_30871# 9.74e-22
C23451 a_5829_43940# a_5755_42308# 9.03e-21
C23452 a_15493_43396# a_15803_42450# 8.19e-21
C23453 a_5649_42852# a_7765_42852# 1.28e-20
C23454 a_n4318_38680# a_n1545_43230# 2.34e-20
C23455 a_n2012_43396# a_n2104_42282# 2.27e-20
C23456 a_16664_43396# a_16414_43172# 4.88e-19
C23457 a_4361_42308# a_8387_43230# 5.06e-20
C23458 a_n2129_44697# VDD 1.4165f
C23459 a_n1352_43396# COMP_P 1.02e-19
C23460 a_n4318_39304# a_n3674_37592# 0.024848f
C23461 a_11341_43940# a_14456_42282# 4.56e-23
C23462 a_21513_45002# a_20640_44752# 1.55e-19
C23463 a_13059_46348# a_14543_43071# 4.18e-19
C23464 a_19692_46634# a_21671_42860# 1.06e-19
C23465 a_n2661_43370# a_n1352_44484# 0.001902f
C23466 a_16922_45042# a_17969_45144# 0.002405f
C23467 a_13249_42308# a_10949_43914# 3.22e-19
C23468 a_4185_45028# a_743_42282# 0.031243f
C23469 a_3232_43370# a_3363_44484# 0.103472f
C23470 a_21101_45002# a_21359_45002# 0.22264f
C23471 a_21005_45260# a_11827_44484# 0.005914f
C23472 a_19778_44110# a_11691_44458# 0.013164f
C23473 a_18911_45144# a_20193_45348# 5.06e-21
C23474 a_3537_45260# a_n2661_43922# 0.058875f
C23475 a_4574_45260# a_n2661_42834# 4.61e-21
C23476 a_11823_42460# a_14955_43940# 6.42e-21
C23477 a_n913_45002# a_14673_44172# 3.55e-20
C23478 a_17613_45144# a_17801_45144# 7.06e-21
C23479 a_10193_42453# a_15493_43396# 0.024143f
C23480 a_5837_45028# a_5883_43914# 4.44e-21
C23481 a_4883_46098# a_11823_42460# 1.64e-19
C23482 a_13507_46334# a_13163_45724# 4.48e-19
C23483 a_11453_44696# a_10490_45724# 6.39e-21
C23484 a_n743_46660# a_380_45546# 0.010247f
C23485 a_7927_46660# a_8034_45724# 9e-20
C23486 a_1123_46634# a_n2661_45546# 4.02e-20
C23487 a_17609_46634# a_18189_46348# 1.41e-19
C23488 a_15227_44166# a_17583_46090# 4.28e-21
C23489 a_765_45546# a_5068_46348# 3.71e-21
C23490 a_12465_44636# a_11962_45724# 1.34e-21
C23491 a_12469_46902# a_10809_44734# 0.014309f
C23492 a_12991_46634# a_6945_45028# 1.08e-19
C23493 a_7411_46660# a_8049_45260# 5.59e-20
C23494 a_n2293_46634# a_997_45618# 0.002767f
C23495 a_n2438_43548# a_n452_45724# 3.99e-20
C23496 a_n133_46660# a_n863_45724# 1.41e-19
C23497 a_n1021_46688# a_n1099_45572# 2.81e-21
C23498 a_n1925_46634# a_310_45028# 5.87e-20
C23499 a_15743_43084# a_21613_42308# 1.45e-19
C23500 a_4190_30871# a_17303_42282# 0.279034f
C23501 a_n2293_42282# COMP_P 0.026882f
C23502 a_10807_43548# CLK 8.86e-22
C23503 a_15493_43396# VDD 2.34659f
C23504 a_7871_42858# a_5934_30871# 0.001545f
C23505 a_4361_42308# a_16522_42674# 0.002806f
C23506 a_7765_42852# a_7963_42308# 9.95e-19
C23507 a_8037_42858# a_6123_31319# 5.06e-20
C23508 a_n2312_40392# VDD 0.947797f
C23509 a_21588_30879# a_22821_38993# 1.81e-19
C23510 a_1823_45246# a_5934_30871# 3.73e-20
C23511 a_n1059_45260# a_n1557_42282# 0.031252f
C23512 a_4883_46098# DATA[3] 2.04e-21
C23513 a_4185_45028# a_5755_42308# 1.64e-19
C23514 a_1307_43914# a_8487_44056# 4.35e-19
C23515 a_17339_46660# a_18057_42282# 1.93e-19
C23516 a_949_44458# a_895_43940# 0.002952f
C23517 a_2779_44458# a_2479_44172# 0.001425f
C23518 a_742_44458# a_2675_43914# 2.91e-21
C23519 a_n2661_43922# a_11541_44484# 0.004005f
C23520 a_n699_43396# a_453_43940# 0.006917f
C23521 a_22959_47212# RST_Z 0.001482f
C23522 a_9482_43914# a_13565_43940# 3.82e-19
C23523 a_11453_44696# START 8.37e-19
C23524 a_n357_42282# a_16414_43172# 0.005649f
C23525 a_n443_42852# a_10991_42826# 1.25e-19
C23526 a_11823_42460# a_5649_42852# 2.49e-19
C23527 a_18479_47436# a_19778_44110# 0.038618f
C23528 a_n743_46660# a_10775_45002# 1.84e-21
C23529 a_5066_45546# a_6347_46155# 7.61e-19
C23530 a_2107_46812# a_6171_45002# 0.023061f
C23531 a_5257_43370# a_3357_43084# 0.894879f
C23532 a_7577_46660# a_2437_43646# 1.39e-20
C23533 a_18819_46122# a_20009_46494# 2.56e-19
C23534 a_167_45260# a_1176_45572# 0.00195f
C23535 a_n2293_46098# a_3733_45822# 5.15e-19
C23536 a_2864_46660# a_413_45260# 9.11e-21
C23537 a_17609_46634# a_17478_45572# 8.56e-20
C23538 a_15227_44166# a_8696_44636# 0.203885f
C23539 a_n1613_43370# a_6945_45348# 1.51e-19
C23540 a_n443_46116# a_n452_44636# 1.47e-20
C23541 a_n1151_42308# a_5343_44458# 1.19e-19
C23542 a_2609_46660# a_2680_45002# 1.09e-20
C23543 a_2443_46660# a_3065_45002# 2.64e-21
C23544 a_16327_47482# a_11827_44484# 0.107078f
C23545 a_18597_46090# a_18587_45118# 6.25e-19
C23546 a_n2840_42826# VDD 0.302305f
C23547 a_2351_42308# a_7174_31319# 4.88e-21
C23548 COMP_P a_n3565_39590# 4.08e-21
C23549 a_n3674_37592# a_n4334_40480# 7.51e-19
C23550 a_11551_42558# a_12563_42308# 2.06e-19
C23551 a_8975_43940# a_10695_43548# 7.03e-21
C23552 a_n357_42282# a_7174_31319# 4.25e-19
C23553 a_n913_45002# a_8292_43218# 0.001438f
C23554 a_16922_45042# a_4361_42308# 0.00825f
C23555 a_10193_42453# a_8791_42308# 2.96e-20
C23556 a_n2810_45572# a_n4315_30879# 0.024132f
C23557 a_11967_42832# a_18533_44260# 0.001389f
C23558 a_n2661_43922# a_1049_43396# 2.6e-21
C23559 a_n2661_42834# a_1568_43370# 1.03e-19
C23560 a_n356_44636# a_8791_43396# 5.34e-22
C23561 a_7499_43078# a_9377_42558# 2.82e-19
C23562 a_9482_43914# a_5534_30871# 1.74e-21
C23563 a_18494_42460# a_19177_43646# 7.87e-20
C23564 a_19778_44110# a_4190_30871# 5.46e-20
C23565 a_18184_42460# a_21259_43561# 5.43e-20
C23566 a_n2293_42834# a_n1379_43218# 4.33e-19
C23567 a_3483_46348# a_1423_45028# 0.110369f
C23568 a_2324_44458# a_5111_44636# 0.090721f
C23569 a_5257_43370# a_5826_44734# 0.003375f
C23570 a_n881_46662# a_n809_44244# 3.25e-20
C23571 a_n1613_43370# a_n984_44318# 0.245331f
C23572 a_9290_44172# a_10951_45334# 0.136064f
C23573 a_2711_45572# a_11962_45724# 0.054424f
C23574 a_14493_46090# a_6171_45002# 6.27e-21
C23575 a_5024_45822# a_4880_45572# 6.84e-19
C23576 a_7227_45028# a_7499_43078# 5.28e-22
C23577 a_20708_46348# a_413_45260# 2.68e-21
C23578 a_20916_46384# a_19279_43940# 1.62e-21
C23579 a_3090_45724# a_n699_43396# 0.058797f
C23580 a_8049_45260# a_20841_45814# 0.008238f
C23581 a_12861_44030# a_10949_43914# 8.34e-19
C23582 a_17339_46660# a_18494_42460# 8.02e-20
C23583 a_n2293_46634# a_11967_42832# 6.03e-20
C23584 a_n2956_38680# en_comp 3.44e-19
C23585 a_n971_45724# a_768_44030# 0.069358f
C23586 a_2063_45854# a_n881_46662# 0.612456f
C23587 a_2553_47502# a_n1613_43370# 3.57e-20
C23588 a_2905_45572# a_3094_47243# 0.006879f
C23589 a_2952_47436# a_3411_47243# 6.64e-19
C23590 a_n3565_39590# a_n3565_37414# 0.032079f
C23591 a_n443_46116# a_2747_46873# 0.047485f
C23592 a_16327_47482# a_16588_47582# 0.276601f
C23593 a_9313_45822# a_4883_46098# 0.026043f
C23594 a_7174_31319# CAL_N 0.018266f
C23595 a_n4209_39590# a_n3420_37440# 0.038354f
C23596 a_15673_47210# a_10227_46804# 0.02634f
C23597 a_11599_46634# a_18780_47178# 3.49e-19
C23598 a_5742_30871# C2_N_btm 0.030783f
C23599 a_13717_47436# a_20990_47178# 9.85e-20
C23600 a_13381_47204# a_13507_46334# 0.001369f
C23601 a_8791_42308# VDD 0.226318f
C23602 a_n3420_38528# a_n4251_38304# 8.88e-19
C23603 a_n3420_39616# a_n4209_37414# 0.027966f
C23604 a_n4064_38528# a_n4064_37984# 0.057015f
C23605 a_5932_42308# VIN_N 0.023512f
C23606 a_11967_42832# a_5342_30871# 0.077151f
C23607 a_5891_43370# a_9306_43218# 5.41e-19
C23608 a_n97_42460# a_1209_43370# 0.027601f
C23609 a_21381_43940# a_2982_43646# 0.236232f
C23610 a_104_43370# a_458_43396# 0.07022f
C23611 a_17737_43940# a_17499_43370# 0.013048f
C23612 a_n2956_37592# a_n3420_39072# 6.43e-20
C23613 a_6472_45840# VDD 0.257073f
C23614 a_14021_43940# a_13667_43396# 4.76e-19
C23615 a_15493_43396# a_16137_43396# 0.023247f
C23616 a_11453_44696# a_16547_43609# 2.27e-20
C23617 a_13507_46334# a_18783_43370# 6.51e-20
C23618 a_21363_45546# a_2437_43646# 0.006526f
C23619 a_21188_45572# a_21513_45002# 0.002147f
C23620 a_n2661_45546# a_n2840_44458# 3.06e-19
C23621 a_16327_47482# a_17433_43396# 2.95e-19
C23622 a_20273_45572# a_3357_43084# 0.358383f
C23623 a_20107_45572# a_22591_45572# 3.89e-21
C23624 a_10227_46804# a_15940_43402# 1.75e-19
C23625 a_15903_45785# a_6171_45002# 0.011492f
C23626 a_n2840_45546# a_n2661_44458# 2.89e-19
C23627 a_n2810_45572# a_n4318_40392# 0.02461f
C23628 a_14493_46090# a_14673_44172# 4.72e-21
C23629 a_10809_44734# a_n2661_42834# 0.14417f
C23630 a_3775_45552# a_n2661_43370# 1.33e-21
C23631 a_19466_46812# a_19862_44208# 4.57e-20
C23632 C0_P_btm C3_N_btm 3.77e-19
C23633 C3_P_btm C6_N_btm 4.24e-19
C23634 C1_P_btm C4_N_btm 1.59e-19
C23635 a_11599_46634# a_18285_46348# 0.030958f
C23636 a_15811_47375# a_765_45546# 0.035109f
C23637 a_n2661_46098# a_1057_46660# 1.99e-19
C23638 a_n2293_46634# a_5257_43370# 0.061974f
C23639 a_n2497_47436# a_3483_46348# 4.12e-20
C23640 a_n1741_47186# a_2521_46116# 1.08e-20
C23641 a_584_46384# a_n1853_46287# 4.85e-21
C23642 a_n1838_35608# VIN_P 0.029423f
C23643 C9_P_btm VDD 0.345685f
C23644 a_2553_47502# a_n2293_46098# 4.34e-23
C23645 a_10227_46804# a_16388_46812# 8.39e-20
C23646 C0_dummy_N_btm C1_N_btm 1.2494f
C23647 a_13717_47436# a_20273_46660# 2.45e-21
C23648 a_n785_47204# a_376_46348# 1.57e-19
C23649 a_n746_45260# a_1208_46090# 3.58e-20
C23650 a_n237_47217# a_805_46414# 1.4e-19
C23651 a_n971_45724# a_1176_45822# 1.67e-19
C23652 a_13661_43548# a_6755_46942# 0.088986f
C23653 a_5807_45002# a_6969_46634# 0.003601f
C23654 a_n2661_46634# a_7577_46660# 0.047111f
C23655 a_3177_46902# a_3524_46660# 0.051162f
C23656 a_2609_46660# a_2864_46660# 0.055869f
C23657 a_2443_46660# a_3067_47026# 9.73e-19
C23658 a_2107_46812# a_4955_46873# 0.031068f
C23659 a_n2661_42282# a_5379_42460# 0.121051f
C23660 a_45_45144# VDD 3.5e-19
C23661 a_17021_43396# a_16823_43084# 0.002675f
C23662 a_1568_43370# a_n2293_42282# 3.41e-20
C23663 a_3626_43646# a_18083_42858# 9.29e-20
C23664 a_2982_43646# a_18249_42858# 6.61e-20
C23665 a_15743_43084# a_4361_42308# 0.020459f
C23666 a_10903_43370# a_2982_43646# 3.15e-19
C23667 a_5937_45572# a_6031_43396# 0.010894f
C23668 a_15903_45785# a_14673_44172# 1.01e-20
C23669 a_2680_45002# a_2779_44458# 1.99e-19
C23670 a_n357_42282# a_10729_43914# 4.51e-22
C23671 a_13661_43548# a_16328_43172# 1.62e-19
C23672 a_9482_43914# a_11691_44458# 0.616964f
C23673 a_14537_43396# a_11827_44484# 0.076354f
C23674 a_5093_45028# a_n2661_43370# 0.005328f
C23675 a_2274_45254# a_n699_43396# 1.36e-20
C23676 a_6171_45002# a_n2661_44458# 0.001196f
C23677 a_2382_45260# a_4223_44672# 5.91e-19
C23678 a_n2312_40392# a_n784_42308# 7.39e-19
C23679 a_n743_46660# a_526_44458# 0.020498f
C23680 a_13661_43548# a_8049_45260# 0.032643f
C23681 a_13059_46348# a_765_45546# 4.68e-19
C23682 a_16388_46812# a_17339_46660# 0.24887f
C23683 a_12549_44172# a_12379_46436# 3.71e-19
C23684 a_12891_46348# a_12638_46436# 0.13727f
C23685 a_8145_46902# a_8349_46414# 7.84e-19
C23686 a_7927_46660# a_8016_46348# 8.96e-19
C23687 a_7715_46873# a_5937_45572# 1.65e-20
C23688 a_7577_46660# a_8199_44636# 1.99e-19
C23689 a_6151_47436# a_6667_45809# 0.1609f
C23690 a_6491_46660# a_6472_45840# 7.23e-22
C23691 a_2063_45854# a_8162_45546# 2.61e-19
C23692 a_6545_47178# a_6511_45714# 4.48e-20
C23693 a_n881_46662# a_14383_46116# 1.43e-19
C23694 a_19692_46634# a_19636_46660# 3.77e-19
C23695 a_14976_45028# a_12741_44636# 3.06e-19
C23696 a_12895_43230# a_12991_43230# 0.013793f
C23697 a_n3674_39304# a_n4318_38216# 0.043431f
C23698 a_13113_42826# a_13157_43218# 3.69e-19
C23699 a_12281_43396# a_11633_42558# 4.33e-21
C23700 a_10341_43396# a_14456_42282# 2.53e-20
C23701 a_4361_42308# a_1606_42308# 1.99e-20
C23702 a_n1991_42858# a_n1329_42308# 0.001762f
C23703 a_n1423_42826# COMP_P 3.47e-19
C23704 a_n4318_38680# a_n2472_42282# 4.31e-19
C23705 a_n1736_43218# a_n3674_38680# 3.47e-20
C23706 a_2982_43646# a_21125_42558# 3.84e-19
C23707 a_n2472_43914# VDD 0.236691f
C23708 a_n1853_43023# a_n961_42308# 2.96e-20
C23709 a_3422_30871# VIN_P 0.057975f
C23710 a_3090_45724# a_11551_42558# 6.89e-20
C23711 a_3357_43084# a_5745_43940# 0.003915f
C23712 a_1307_43914# a_3499_42826# 0.532672f
C23713 a_21101_45002# a_19279_43940# 6.46e-20
C23714 a_11827_44484# a_20835_44721# 0.009929f
C23715 a_n1741_47186# DATA[5] 0.069294f
C23716 a_2711_45572# a_17499_43370# 2.44e-19
C23717 a_8746_45002# a_9803_43646# 1.37e-20
C23718 a_327_47204# VDD 0.367528f
C23719 a_8701_44490# a_n2661_43922# 0.00848f
C23720 a_5883_43914# a_n2661_42834# 0.106812f
C23721 a_10334_44484# a_10617_44484# 0.003683f
C23722 a_15004_44636# a_9313_44734# 6.27e-21
C23723 a_9482_43914# a_8333_44056# 6.18e-20
C23724 a_18494_42460# a_18579_44172# 2.2e-19
C23725 a_16922_45042# a_20397_44484# 3.67e-19
C23726 a_n443_42852# a_15231_43396# 4.71e-19
C23727 a_9290_44172# a_9306_43218# 1.97e-21
C23728 a_n2293_42834# a_2127_44172# 3.16e-21
C23729 a_n2661_43370# a_n1549_44318# 8.71e-21
C23730 a_626_44172# a_1241_44260# 1.9e-19
C23731 a_n2661_45010# a_2253_43940# 0.003669f
C23732 a_n2293_45010# a_1241_43940# 0.005122f
C23733 a_n971_45724# DATA[0] 0.213213f
C23734 a_n2312_38680# a_n3690_38528# 5.77e-19
C23735 a_11823_42460# a_8685_43396# 0.057344f
C23736 a_8349_46414# a_5066_45546# 0.005369f
C23737 a_9863_46634# a_10210_45822# 2.83e-20
C23738 a_4185_45028# a_8049_45260# 0.014062f
C23739 a_768_44030# a_n2293_45010# 0.03517f
C23740 a_n1613_43370# a_n467_45028# 0.004184f
C23741 a_10227_46804# a_13777_45326# 9.51e-19
C23742 a_5807_45002# a_3357_43084# 0.071743f
C23743 a_11453_44696# a_6171_45002# 1.39146f
C23744 a_4883_46098# a_7705_45326# 4.33e-20
C23745 a_18819_46122# a_21137_46414# 2.71e-21
C23746 a_19553_46090# a_19900_46494# 0.051162f
C23747 a_18985_46122# a_20708_46348# 2.48e-19
C23748 a_17715_44484# a_10809_44734# 1.44e-19
C23749 a_19452_47524# a_2437_43646# 0.001463f
C23750 a_19321_45002# a_21513_45002# 0.002479f
C23751 a_2063_45854# a_11361_45348# 6.44e-22
C23752 a_584_46384# a_n2661_43370# 0.034714f
C23753 a_1184_42692# a_5934_30871# 8.33e-21
C23754 a_2351_42308# a_5932_42308# 4.34e-21
C23755 a_1606_42308# a_6761_42308# 1.94e-20
C23756 a_3823_42558# a_3905_42558# 0.171361f
C23757 a_10695_43548# VDD 0.201247f
C23758 a_n784_42308# a_8791_42308# 3.86e-20
C23759 a_n357_42282# a_5932_42308# 6.58e-19
C23760 a_n755_45592# a_6171_42473# 1.56e-19
C23761 a_15433_44458# a_15493_43940# 0.001343f
C23762 a_n2661_42834# a_12495_44260# 8.52e-19
C23763 a_1467_44172# a_453_43940# 0.05905f
C23764 a_1115_44172# a_2127_44172# 2.04e-20
C23765 a_17517_44484# a_17973_43940# 4.57e-20
C23766 a_175_44278# a_895_43940# 2.38e-19
C23767 a_n863_45724# a_6123_31319# 8.96e-21
C23768 a_n2956_39304# a_n4209_39590# 0.022939f
C23769 a_10193_42453# a_18707_42852# 0.003123f
C23770 a_18287_44626# a_19319_43548# 1.07e-20
C23771 a_18989_43940# a_18533_44260# 3.53e-19
C23772 a_n913_45002# a_3681_42891# 1.8e-20
C23773 a_n1059_45260# a_3935_42891# 0.004841f
C23774 a_n2017_45002# a_4520_42826# 5.33e-20
C23775 a_742_44458# a_1209_43370# 1.04e-19
C23776 a_949_44458# a_458_43396# 0.001416f
C23777 a_13259_45724# a_13249_42558# 8.98e-20
C23778 a_1848_45724# a_1609_45822# 0.042695f
C23779 a_n356_45724# a_7_45899# 0.005265f
C23780 a_n755_45592# a_1990_45899# 9.01e-21
C23781 a_584_46384# a_2998_44172# 0.181241f
C23782 a_18479_47436# a_20159_44458# 3.97e-21
C23783 a_18597_46090# a_11967_42832# 0.021692f
C23784 a_16327_47482# a_18005_44484# 0.001967f
C23785 a_380_45546# a_509_45572# 0.010132f
C23786 a_n1099_45572# a_n89_45572# 9.15e-19
C23787 a_8034_45724# a_8336_45822# 8.44e-21
C23788 a_11315_46155# a_10193_42453# 7.86e-19
C23789 a_n2497_47436# a_261_44278# 0.002478f
C23790 a_n971_45724# a_7845_44172# 1.69e-20
C23791 a_n2293_46098# a_n467_45028# 2.4e-21
C23792 a_1823_45246# a_n2661_45010# 1.68e-19
C23793 a_n881_46662# a_n2661_42834# 6.26e-20
C23794 a_4185_45028# a_19479_31679# 0.03554f
C23795 a_n1613_43370# a_n2661_43922# 0.113996f
C23796 a_n2661_45546# a_4099_45572# 0.008087f
C23797 a_11453_44696# a_14673_44172# 0.001076f
C23798 a_12861_44030# a_3422_30871# 0.018986f
C23799 a_n1076_46494# a_n745_45366# 5.48e-20
C23800 a_n1991_46122# a_n967_45348# 1.72e-20
C23801 a_2324_44458# a_16147_45260# 1.7e-19
C23802 a_768_44030# a_9313_44734# 0.044729f
C23803 a_10809_44734# a_15861_45028# 8.82e-22
C23804 a_n4209_39590# a_n3565_39304# 0.032081f
C23805 a_n3420_39616# a_n3607_39616# 0.001546f
C23806 a_6123_31319# a_6886_37412# 4.22e-19
C23807 a_n784_42308# C9_P_btm 9.31e-20
C23808 a_2063_45854# a_n443_46116# 0.177177f
C23809 a_2905_45572# a_4007_47204# 0.001036f
C23810 a_n1151_42308# a_3785_47178# 0.029415f
C23811 a_n237_47217# a_7903_47542# 0.086772f
C23812 a_n1920_47178# a_n1435_47204# 0.001089f
C23813 a_3160_47472# a_3815_47204# 1.5e-19
C23814 a_n1741_47186# a_13381_47204# 4.11e-19
C23815 a_n3565_39590# a_n4209_39304# 5.4667f
C23816 a_n4064_40160# a_n4064_39072# 0.06545f
C23817 a_14097_32519# C7_N_btm 7.66e-20
C23818 a_n1630_35242# a_19120_35138# 7.97e-19
C23819 a_18707_42852# VDD 0.132317f
C23820 a_n4334_39616# a_n4334_39392# 0.052468f
C23821 a_20159_44458# a_4190_30871# 1.81e-20
C23822 a_11967_42832# a_743_42282# 0.043946f
C23823 a_16979_44734# a_17333_42852# 4.43e-22
C23824 a_14539_43914# a_18249_42858# 2.08e-19
C23825 a_2382_45260# a_5742_30871# 1.17e-20
C23826 en_comp a_15051_42282# 1.64e-19
C23827 a_n356_44636# a_12895_43230# 1.3e-20
C23828 a_1307_43914# a_3318_42354# 0.001768f
C23829 a_n2293_42834# a_n4318_38216# 7.97e-19
C23830 a_5111_44636# a_9803_42558# 2.44e-21
C23831 a_n1059_45260# a_15890_42674# 2.22e-20
C23832 a_n913_45002# a_15959_42545# 3.53e-19
C23833 a_n2017_45002# a_15720_42674# 1.72e-19
C23834 a_5891_43370# a_8387_43230# 0.010767f
C23835 a_17767_44458# a_18083_42858# 1.98e-19
C23836 a_742_44458# a_3059_42968# 1.47e-19
C23837 a_17517_44484# a_22591_43396# 7.11e-20
C23838 a_11315_46155# VDD 1.9e-20
C23839 a_13661_43548# a_15037_43940# 2.04e-19
C23840 a_n443_42852# a_9482_43914# 1.75e-19
C23841 a_n755_45592# a_1145_45348# 7.7e-19
C23842 a_997_45618# a_626_44172# 1.07e-19
C23843 a_12549_44172# a_17538_32519# 1.42e-19
C23844 a_2711_45572# a_7229_43940# 0.001392f
C23845 a_8049_45260# a_18587_45118# 2.06e-21
C23846 a_15765_45572# a_18341_45572# 0.001304f
C23847 a_n1613_43370# a_n447_43370# 7.94e-19
C23848 a_5907_45546# a_6171_45002# 0.001025f
C23849 a_6194_45824# a_3232_43370# 1.03e-19
C23850 a_3483_46348# a_6109_44484# 0.003232f
C23851 a_13507_46334# a_3626_43646# 0.04477f
C23852 a_3316_45546# a_1307_43914# 1.38e-19
C23853 a_n357_42282# a_1423_45028# 2.14e-20
C23854 a_10903_43370# a_14539_43914# 3.63e-21
C23855 a_n2312_40392# a_3080_42308# 5.51e-21
C23856 a_8270_45546# a_7281_43914# 1.81e-20
C23857 a_8696_44636# a_16377_45572# 2.13e-20
C23858 a_16855_45546# a_16147_45260# 1.95e-19
C23859 a_n2293_46098# a_n2661_43922# 0.026124f
C23860 a_12741_44636# a_15433_44458# 0.004093f
C23861 a_n3420_37440# C6_P_btm 1.87e-19
C23862 a_n4209_37414# C2_P_btm 0.001057f
C23863 a_n3565_37414# C4_P_btm 9.91e-21
C23864 a_14955_47212# a_6755_46942# 4.64e-19
C23865 a_11599_46634# a_10249_46116# 7.84e-19
C23866 a_5807_45002# a_n2293_46634# 9.62e-19
C23867 a_n1151_42308# a_3090_45724# 0.003613f
C23868 a_4915_47217# a_11901_46660# 0.004227f
C23869 a_6575_47204# a_8189_46660# 1.95e-20
C23870 a_n1613_43370# a_1799_45572# 0.008733f
C23871 a_n4064_37984# VREF_GND 0.047292f
C23872 a_4883_46098# a_6540_46812# 2.72e-20
C23873 a_22545_38993# a_22780_39857# 0.003614f
C23874 a_22521_39511# a_22876_39857# 0.011942f
C23875 a_22521_40599# a_22717_37285# 0.010048f
C23876 a_22459_39145# a_22609_38406# 0.12318f
C23877 a_22469_40625# a_22705_37990# 0.010408f
C23878 a_22521_40055# a_22705_38406# 0.010302f
C23879 a_22821_38993# a_22469_39537# 0.039707f
C23880 a_9145_43396# a_16547_43609# 2.43e-21
C23881 a_19479_31679# VREF_GND 0.00198f
C23882 a_3539_42460# a_4361_42308# 0.027414f
C23883 a_10341_43396# a_10149_43396# 7.68e-19
C23884 a_n1761_44111# a_n473_42460# 0.110251f
C23885 a_17730_32519# a_n1630_35242# 5.92e-20
C23886 a_n356_44636# a_18220_42308# 5.19e-19
C23887 a_n745_45366# VDD 0.20887f
C23888 a_n229_43646# a_n13_43084# 3.17e-20
C23889 a_n1821_43396# a_n4318_38680# 1.73e-19
C23890 a_n913_45002# RST_Z 2.65e-19
C23891 a_648_43396# a_743_42282# 4.53e-21
C23892 a_15095_43370# a_15681_43442# 3.23e-21
C23893 a_14205_43396# a_15781_43660# 9.18e-21
C23894 a_14021_43940# a_21195_42852# 8.07e-21
C23895 a_2982_43646# a_5649_42852# 0.205161f
C23896 a_13667_43396# a_13943_43396# 0.00119f
C23897 a_20447_31679# EN_OFFSET_CAL 2.14e-19
C23898 a_6171_45002# a_6125_45348# 4.58e-19
C23899 a_5257_43370# a_743_42282# 1.37e-19
C23900 a_12549_44172# a_19339_43156# 1.24e-20
C23901 a_15227_44166# a_14205_43396# 1.11e-19
C23902 a_14537_43396# a_15595_45028# 5.49e-20
C23903 a_15037_45618# a_15004_44636# 5.28e-20
C23904 a_8696_44636# a_9838_44484# 0.004732f
C23905 a_2382_45260# a_n2293_42834# 0.026697f
C23906 a_10227_46804# a_10752_42852# 1.7e-19
C23907 a_5807_45002# a_5342_30871# 1.35e-22
C23908 a_5937_45572# a_6671_43940# 0.06027f
C23909 a_13777_45326# a_1307_43914# 3.69e-21
C23910 a_n2293_46634# a_10518_42984# 4.29e-20
C23911 a_4558_45348# a_5009_45028# 0.013349f
C23912 a_5807_45002# a_9625_46129# 0.001468f
C23913 a_6755_46942# a_14543_46987# 4.62e-19
C23914 a_12891_46348# a_13759_46122# 2.87e-20
C23915 a_n2661_46634# a_4704_46090# 1.84e-20
C23916 a_7577_46660# a_765_45546# 0.002481f
C23917 a_n881_46662# a_17715_44484# 0.014166f
C23918 a_14955_47212# a_8049_45260# 1.17e-21
C23919 a_n2497_47436# a_n357_42282# 0.046314f
C23920 a_12549_44172# a_13351_46090# 0.014836f
C23921 a_768_44030# a_12594_46348# 0.001137f
C23922 a_n743_46660# a_2521_46116# 0.013075f
C23923 a_948_46660# a_472_46348# 7.34e-19
C23924 a_n2438_43548# a_167_45260# 0.050543f
C23925 a_2107_46812# a_376_46348# 7.16e-20
C23926 a_n746_45260# a_n2661_45546# 0.022378f
C23927 a_n971_45724# a_n2472_45546# 7.36e-20
C23928 a_n2109_47186# a_n1099_45572# 1.08e-20
C23929 a_n1925_46634# a_2804_46116# 3.92e-20
C23930 a_n2661_46098# a_n2472_46090# 0.094589f
C23931 a_1799_45572# a_n2293_46098# 0.014011f
C23932 a_16137_43396# a_18707_42852# 0.001058f
C23933 a_3422_30871# a_11206_38545# 1.36e-20
C23934 a_n97_42460# a_14456_42282# 0.067807f
C23935 a_3626_43646# a_7227_42308# 0.004361f
C23936 a_2982_43646# a_7963_42308# 8.09e-20
C23937 a_12379_42858# a_12895_43230# 0.109156f
C23938 a_12089_42308# a_13113_42826# 6.01e-19
C23939 a_5649_42852# a_5837_42852# 0.001623f
C23940 a_3363_44484# VDD 1.62e-19
C23941 a_n2661_44458# a_12607_44458# 1.59e-19
C23942 a_327_44734# a_453_43940# 8.52e-21
C23943 a_413_45260# a_2127_44172# 0.104737f
C23944 a_n2661_45010# a_n3674_39768# 0.001075f
C23945 a_2437_43646# a_2253_44260# 2.98e-19
C23946 a_9290_44172# a_8387_43230# 1.54e-20
C23947 a_5257_43370# a_5755_42308# 3.66e-19
C23948 a_19692_46634# a_20256_43172# 4.35e-19
C23949 a_n443_42852# a_6031_43396# 0.020526f
C23950 a_n2312_39304# a_n3420_39072# 6.52e-19
C23951 a_18479_45785# a_15493_43396# 0.235084f
C23952 a_526_44458# a_4361_42308# 0.072573f
C23953 a_8953_45546# a_10835_43094# 5.45e-21
C23954 a_3483_46348# a_15567_42826# 8.48e-21
C23955 a_13059_46348# a_13291_42460# 0.007788f
C23956 a_n699_43396# a_4743_44484# 0.235328f
C23957 a_4223_44672# a_5343_44458# 0.229803f
C23958 a_13661_43548# a_13258_32519# 6.71e-21
C23959 a_3483_46348# a_9569_46155# 1.05e-19
C23960 a_4419_46090# a_5937_45572# 8.29e-20
C23961 a_22365_46825# a_10809_44734# 0.010841f
C23962 a_18597_46090# a_20273_45572# 0.048762f
C23963 a_14311_47204# a_3357_43084# 1.17e-19
C23964 a_15507_47210# a_2437_43646# 0.027848f
C23965 a_n743_46660# a_13163_45724# 1.17e-20
C23966 a_2063_45854# a_3537_45260# 1.21e-20
C23967 a_584_46384# a_4574_45260# 0.001263f
C23968 a_3815_47204# a_413_45260# 5.94e-19
C23969 a_n881_46662# a_15861_45028# 0.153795f
C23970 a_18479_47436# a_20623_45572# 0.007543f
C23971 a_4646_46812# a_6472_45840# 0.129446f
C23972 a_12741_44636# a_19900_46494# 0.005543f
C23973 a_n971_45724# a_7276_45260# 2.9e-22
C23974 a_768_44030# a_15037_45618# 1.6e-21
C23975 a_14976_45028# a_16375_45002# 1.01e-20
C23976 a_3090_45724# a_19240_46482# 2.23e-19
C23977 a_4817_46660# a_5263_45724# 2.13e-19
C23978 a_2107_46812# a_8746_45002# 0.020783f
C23979 a_20202_43084# a_22223_46124# 1.62e-19
C23980 a_11415_45002# a_6945_45028# 0.002828f
C23981 a_10227_46804# a_21188_45572# 1.59e-21
C23982 a_3080_42308# C9_P_btm 9.33e-20
C23983 a_5534_30871# a_4958_30871# 0.024536f
C23984 a_7309_42852# a_6123_31319# 9.07e-19
C23985 a_14097_32519# COMP_P 7e-21
C23986 a_n2433_43396# VDD 0.416276f
C23987 a_16795_42852# a_17124_42282# 3.59e-19
C23988 a_17701_42308# a_16104_42674# 7.22e-21
C23989 a_n2840_42282# a_n2472_42282# 7.52e-19
C23990 a_4185_45028# a_13258_32519# 0.068774f
C23991 a_n2293_42834# a_n1655_43396# 3.89e-19
C23992 a_11967_42832# a_19789_44512# 5.08e-19
C23993 a_1307_43914# a_6197_43396# 7.34e-20
C23994 a_10193_42453# a_21356_42826# 1.27e-19
C23995 a_1983_46706# VDD 0.119964f
C23996 a_16112_44458# a_15682_43940# 0.006723f
C23997 a_17517_44484# a_22591_44484# 0.196232f
C23998 a_n2661_43922# a_2675_43914# 0.002037f
C23999 a_n2661_42834# a_2889_44172# 0.005688f
C24000 a_14539_43914# a_14955_43940# 0.064683f
C24001 a_2324_44458# a_15051_42282# 2.79e-19
C24002 a_6171_45002# a_9145_43396# 3.37e-21
C24003 a_3232_43370# a_9803_43646# 2.81e-21
C24004 a_601_46902# DATA[0] 2.35e-19
C24005 a_n2661_43370# a_n1177_43370# 3.12e-21
C24006 a_626_44172# a_648_43396# 0.04847f
C24007 a_n357_42282# a_17141_43172# 7.19e-19
C24008 a_n2017_45002# a_16409_43396# 1.12e-20
C24009 a_n913_45002# a_16243_43396# 3.59e-20
C24010 a_n1059_45260# a_16547_43609# 0.024317f
C24011 a_n743_46660# DATA[5] 5.08e-21
C24012 a_20766_44850# a_19279_43940# 0.021466f
C24013 a_11453_44696# a_12607_44458# 7.57e-20
C24014 a_16375_45002# a_18051_46116# 0.038793f
C24015 a_5937_45572# a_6469_45572# 1.2e-19
C24016 a_12594_46348# a_11652_45724# 5.18e-20
C24017 a_2324_44458# a_9049_44484# 0.102942f
C24018 a_6755_46942# a_13159_45002# 1.18e-21
C24019 a_13747_46662# a_11691_44458# 3.75e-19
C24020 a_13661_43548# a_20193_45348# 1.38e-20
C24021 a_n443_46116# a_n2661_42834# 0.075503f
C24022 a_4791_45118# a_n2661_43922# 0.034957f
C24023 a_14976_45028# a_413_45260# 3.29e-20
C24024 a_n1613_43370# a_n452_44636# 0.001807f
C24025 a_10903_43370# a_12427_45724# 0.083943f
C24026 a_12005_46116# a_11962_45724# 1.83e-19
C24027 a_n743_46660# a_16501_45348# 8.3e-19
C24028 a_17303_42282# a_19511_42282# 0.001918f
C24029 a_5934_30871# comp_n 1.4e-19
C24030 a_n1630_35242# VDAC_Pi 1.06e-19
C24031 a_21356_42826# VDD 0.225688f
C24032 a_18057_42282# a_18310_42308# 0.011913f
C24033 a_5534_30871# VCM 0.095752f
C24034 a_5742_30871# a_1239_39587# 1.45e-19
C24035 a_20922_43172# RST_Z 2.99e-22
C24036 a_n1059_45260# a_n3674_37592# 1.1e-19
C24037 a_n2017_45002# a_564_42282# 0.013024f
C24038 a_895_43940# a_n97_42460# 0.002734f
C24039 a_10355_46116# CLK 0.002305f
C24040 a_15367_44484# a_8685_43396# 2.8e-22
C24041 a_175_44278# a_458_43396# 4.64e-19
C24042 a_9313_44734# a_16759_43396# 8.78e-20
C24043 a_11827_44484# a_12379_42858# 2.49e-21
C24044 a_n967_45348# a_n1329_42308# 0.033651f
C24045 a_14275_46494# VDD 0.196859f
C24046 a_15493_43396# a_14021_43940# 0.139192f
C24047 a_14673_44172# a_9145_43396# 1.46e-19
C24048 en_comp a_n961_42308# 6.61e-20
C24049 a_n2293_42834# a_1709_42852# 2.82e-20
C24050 a_11189_46129# DATA[5] 1.65e-20
C24051 a_n2956_38216# a_n2472_45002# 0.00378f
C24052 a_n755_45592# a_3357_43084# 0.00172f
C24053 a_n2293_45546# a_n2661_45010# 0.014846f
C24054 a_526_44458# a_2809_45348# 0.001579f
C24055 a_6945_45028# a_6945_45348# 0.009798f
C24056 a_584_46384# a_1568_43370# 0.057089f
C24057 a_n1641_46494# a_n2267_44484# 4.94e-19
C24058 a_6755_46942# a_11967_42832# 0.030705f
C24059 a_2324_44458# a_13105_45348# 2.03e-19
C24060 a_11823_42460# a_11778_45572# 8.46e-20
C24061 a_n1853_46287# a_n1177_44458# 5.46e-23
C24062 a_10193_42453# a_15765_45572# 1.09e-19
C24063 a_8568_45546# a_8696_44636# 4.42e-20
C24064 a_4185_45028# a_20193_45348# 0.015456f
C24065 a_n2472_45546# a_n2293_45010# 3.35e-19
C24066 a_n2661_45546# a_n2109_45247# 0.003324f
C24067 a_12549_44172# a_17973_43940# 0.015874f
C24068 a_8049_45260# a_13159_45002# 4.59e-21
C24069 a_376_46348# a_n2661_44458# 9.54e-22
C24070 a_19123_46287# a_18989_43940# 2.88e-20
C24071 a_n4064_40160# VDD 2.37253f
C24072 a_7754_40130# a_5088_37509# 0.036831f
C24073 a_7754_39964# a_3726_37500# 0.030605f
C24074 a_2747_46873# a_n1613_43370# 0.03071f
C24075 a_18780_47178# a_13661_43548# 0.153988f
C24076 a_18479_47436# a_13747_46662# 0.083389f
C24077 a_n4064_39072# C10_P_btm 1.08e-19
C24078 VDAC_Ni a_3754_38470# 0.911632f
C24079 a_10227_46804# a_19321_45002# 0.111029f
C24080 a_n1151_42308# a_3699_46634# 1.12e-19
C24081 a_3381_47502# a_2959_46660# 0.005389f
C24082 a_3160_47472# a_3524_46660# 1.52e-20
C24083 a_584_46384# a_2162_46660# 0.001394f
C24084 a_n3565_39304# C6_P_btm 0.080378f
C24085 a_n3420_39072# C8_P_btm 8.3e-20
C24086 a_12465_44636# a_768_44030# 0.120859f
C24087 a_13381_47204# a_n743_46660# 1.37e-20
C24088 a_n971_45724# a_5167_46660# 3.91e-20
C24089 a_n237_47217# a_4817_46660# 6.61e-20
C24090 a_n4209_38502# a_n1532_35090# 9.11e-20
C24091 a_n3565_38502# a_n1838_35608# 1.42e-19
C24092 a_7174_31319# VIN_P 0.022822f
C24093 a_18597_46090# a_5807_45002# 0.005073f
C24094 a_13258_32519# VREF_GND 0.033872f
C24095 a_n2956_37592# a_n2946_37690# 0.148852f
C24096 a_15765_45572# VDD 0.249471f
C24097 a_19479_31679# a_22469_40625# 1.34e-20
C24098 a_10405_44172# a_10083_42826# 1.98e-19
C24099 a_5891_43370# a_1606_42308# 5.17e-20
C24100 a_5343_44458# a_5742_30871# 9.93e-21
C24101 a_n2661_42834# a_n4318_37592# 1.57e-19
C24102 a_n2810_45028# a_n4064_37440# 0.22413f
C24103 a_8975_43940# a_8685_42308# 1.95e-22
C24104 a_n2293_43922# a_n3674_38216# 0.032717f
C24105 a_2982_43646# a_8685_43396# 6.82e-20
C24106 a_11967_42832# a_16328_43172# 0.001925f
C24107 a_18494_42460# a_18310_42308# 0.001869f
C24108 a_19319_43548# a_19268_43646# 0.17076f
C24109 a_7287_43370# a_7112_43396# 0.234322f
C24110 a_6031_43396# a_6655_43762# 9.73e-19
C24111 a_6293_42852# a_6452_43396# 0.157972f
C24112 a_10227_46804# a_10922_42852# 0.159426f
C24113 a_2711_45572# a_15004_44636# 5.78e-22
C24114 a_8746_45002# a_n2661_44458# 0.017636f
C24115 a_n913_45002# a_3232_43370# 6.56e-20
C24116 a_5807_45002# a_743_42282# 2.41e-20
C24117 a_n443_46116# a_n2293_42282# 2.82e-20
C24118 a_n1613_43370# a_n1641_43230# 0.152896f
C24119 a_413_45260# a_2382_45260# 0.048205f
C24120 a_n357_42282# a_6109_44484# 1.45e-19
C24121 a_8696_44636# a_n2661_43370# 0.674122f
C24122 a_2324_44458# a_3905_42865# 1.55e-19
C24123 a_13661_43548# a_20301_43646# 0.072262f
C24124 a_13747_46662# a_4190_30871# 4.43e-21
C24125 a_8667_46634# a_10150_46912# 5.2e-20
C24126 a_8492_46660# a_9863_46634# 5.2e-20
C24127 a_6540_46812# a_6682_46660# 0.007833f
C24128 a_2747_46873# a_n2293_46098# 3.99e-20
C24129 a_4883_46098# a_1823_45246# 0.00603f
C24130 a_n2109_47186# a_n1925_42282# 2.07e-20
C24131 a_5257_43370# a_6755_46942# 8.35e-20
C24132 a_6151_47436# a_14840_46494# 4.06e-20
C24133 a_5807_45002# a_19123_46287# 0.006772f
C24134 a_13661_43548# a_18285_46348# 0.049064f
C24135 a_n1435_47204# a_9290_44172# 6.71e-22
C24136 a_19321_45002# a_17339_46660# 1.05e-20
C24137 a_18429_43548# a_17333_42852# 0.003673f
C24138 a_18525_43370# a_18083_42858# 0.016073f
C24139 a_15743_43084# a_17595_43084# 7.44e-20
C24140 a_743_42282# a_10518_42984# 2.81e-20
C24141 a_n4318_38680# a_n1736_43218# 4.04e-20
C24142 a_5745_43940# a_5755_42308# 5.58e-22
C24143 a_15493_43396# a_15764_42576# 1.23e-21
C24144 a_5649_42852# a_7871_42858# 1.53e-20
C24145 a_n1853_43023# a_685_42968# 1.6e-20
C24146 a_n1076_43230# a_n967_43230# 0.007416f
C24147 a_n901_43156# a_n722_43218# 0.007399f
C24148 a_n1641_43230# a_n1533_42852# 0.057222f
C24149 a_17538_32519# a_n1630_35242# 4.52e-20
C24150 a_n2433_44484# VDD 0.40658f
C24151 a_4361_42308# a_8605_42826# 3.01e-20
C24152 a_10193_42453# a_19328_44172# 4.1e-19
C24153 a_13059_46348# a_13460_43230# 5.21e-21
C24154 a_19692_46634# a_21195_42852# 6.29e-21
C24155 a_n2661_43370# a_n1177_44458# 0.002135f
C24156 a_16922_45042# a_17896_45144# 0.003722f
C24157 a_5111_44636# a_5708_44484# 0.002882f
C24158 a_13249_42308# a_10729_43914# 3.94e-20
C24159 a_n2293_42834# a_5343_44458# 0.165923f
C24160 a_18587_45118# a_20193_45348# 4.24e-21
C24161 a_18911_45144# a_11691_44458# 0.013593f
C24162 a_20567_45036# a_11827_44484# 0.004169f
C24163 a_21005_45260# a_21359_45002# 0.001885f
C24164 a_3537_45260# a_n2661_42834# 0.097192f
C24165 a_11823_42460# a_13483_43940# 0.029429f
C24166 a_n1059_45260# a_14673_44172# 7.92e-21
C24167 a_3065_45002# a_n2293_43922# 3.78e-20
C24168 a_n881_46662# a_3775_45552# 0.002767f
C24169 a_11453_44696# a_8746_45002# 0.002934f
C24170 a_768_44030# a_2711_45572# 0.529995f
C24171 a_15227_44166# a_15682_46116# 1.07e-20
C24172 a_17609_46634# a_17715_44484# 0.001359f
C24173 a_4915_47217# a_8696_44636# 0.02426f
C24174 a_765_45546# a_4704_46090# 7.8e-21
C24175 a_22959_46660# a_21076_30879# 0.165603f
C24176 a_11901_46660# a_10809_44734# 0.048084f
C24177 a_n2293_46634# a_n755_45592# 0.094759f
C24178 a_n2438_43548# a_n863_45724# 0.07341f
C24179 a_n743_46660# a_n452_45724# 0.070244f
C24180 a_n1925_46634# a_n1099_45572# 0.001556f
C24181 a_15743_43084# a_21887_42336# 3.74e-20
C24182 a_19700_43370# a_7174_31319# 2.53e-19
C24183 a_21259_43561# a_17303_42282# 9.51e-21
C24184 a_4190_30871# a_4958_30871# 11.510201f
C24185 a_n2293_42282# a_n4318_37592# 0.004341f
C24186 a_10949_43914# CLK 1.96e-21
C24187 a_19328_44172# VDD 0.263964f
C24188 a_n914_42852# a_n4318_38216# 5.63e-21
C24189 a_7765_42852# a_6123_31319# 6.64e-19
C24190 a_7871_42858# a_7963_42308# 3.99e-19
C24191 a_22612_30879# a_22521_39511# 9.02e-20
C24192 a_n357_42282# a_15567_42826# 0.008527f
C24193 a_n699_43396# a_1414_42308# 0.104607f
C24194 a_n913_45002# a_4905_42826# 0.101072f
C24195 a_n2017_45002# a_n1557_42282# 0.090464f
C24196 a_1307_43914# a_8415_44056# 5.17e-19
C24197 a_3065_45002# a_n97_42460# 0.019675f
C24198 a_949_44458# a_2479_44172# 3.43e-19
C24199 a_742_44458# a_895_43940# 0.025021f
C24200 a_10193_42453# a_20749_43396# 1.81e-19
C24201 a_n2661_43922# a_10809_44484# 1.69e-19
C24202 a_11453_44696# RST_Z 0.004685f
C24203 a_9290_44172# a_1606_42308# 9.18e-20
C24204 a_n443_42852# a_10796_42968# 1.54e-19
C24205 a_22959_47212# VDD 0.245964f
C24206 a_11599_46634# a_11691_44458# 7.06e-20
C24207 a_5066_45546# a_8034_45724# 0.242476f
C24208 a_n2661_46634# a_9482_43914# 9.45e-19
C24209 a_n743_46660# a_8953_45002# 0.001504f
C24210 a_2107_46812# a_3232_43370# 0.026265f
C24211 a_584_46384# a_5883_43914# 2.91e-20
C24212 a_7715_46873# a_2437_43646# 2.14e-19
C24213 a_19335_46494# a_19431_46494# 0.013793f
C24214 a_19900_46494# a_16375_45002# 9.97e-21
C24215 a_n2293_46098# a_3638_45822# 4.88e-19
C24216 a_3524_46660# a_413_45260# 4.83e-21
C24217 a_17609_46634# a_15861_45028# 2.54e-19
C24218 a_15368_46634# a_16223_45938# 6.08e-20
C24219 a_n881_46662# a_5093_45028# 8.78e-20
C24220 a_2443_46660# a_2680_45002# 3.28e-21
C24221 a_6945_45028# a_13259_45724# 7.64e-20
C24222 a_16327_47482# a_21359_45002# 2.1e-19
C24223 a_18597_46090# a_18315_45260# 1.77e-20
C24224 a_n4318_38216# a_n4064_39616# 0.024304f
C24225 a_17364_32525# RST_Z 0.050609f
C24226 a_20749_43396# VDD 7.57e-19
C24227 a_4190_30871# VCM 1.23535f
C24228 a_n3674_38216# a_n3420_39616# 0.02009f
C24229 a_n3674_37592# a_n4315_30879# 7.52e-19
C24230 a_2123_42473# a_7174_31319# 4.88e-21
C24231 a_11551_42558# a_11633_42558# 0.171361f
C24232 a_5742_30871# a_12563_42308# 1.19e-20
C24233 a_10057_43914# a_10695_43548# 0.148476f
C24234 a_12607_44458# a_9145_43396# 2.06e-20
C24235 a_n357_42282# a_20712_42282# 0.173926f
C24236 a_n1059_45260# a_8292_43218# 0.002071f
C24237 a_3537_45260# a_n2293_42282# 0.001815f
C24238 a_3065_45002# a_3935_43218# 5.01e-19
C24239 a_10193_42453# a_8685_42308# 3e-20
C24240 a_14539_43914# a_8685_43396# 5.25e-19
C24241 a_8975_43940# a_9803_43646# 8.14e-21
C24242 a_17517_44484# a_20974_43370# 1.2e-20
C24243 a_n2661_42834# a_1049_43396# 6.94e-20
C24244 a_n2661_43922# a_1209_43370# 1.01e-21
C24245 a_20273_46660# EN_OFFSET_CAL 3.18e-20
C24246 a_18280_46660# VDD 6.19e-19
C24247 a_n356_44636# a_8147_43396# 6.99e-22
C24248 a_7499_43078# a_9293_42558# 1.64e-19
C24249 a_13556_45296# a_13460_43230# 1.23e-19
C24250 a_18911_45144# a_4190_30871# 1.03e-21
C24251 a_n2293_42834# a_n1545_43230# 8.56e-19
C24252 a_1423_45028# a_8952_43230# 6.06e-21
C24253 a_9290_44172# a_10775_45002# 0.215292f
C24254 a_3147_46376# a_1423_45028# 8.68e-21
C24255 a_1823_45246# a_3602_45348# 0.001718f
C24256 a_2324_44458# a_5147_45002# 0.056065f
C24257 a_n1613_43370# a_n809_44244# 0.291484f
C24258 a_2711_45572# a_11652_45724# 0.013232f
C24259 a_13925_46122# a_6171_45002# 2.53e-20
C24260 a_19321_45002# a_18579_44172# 0.00855f
C24261 a_3090_45724# a_4223_44672# 0.269823f
C24262 a_8049_45260# a_20273_45572# 0.040989f
C24263 a_12861_44030# a_10729_43914# 3.15e-20
C24264 a_17339_46660# a_18184_42460# 3.97e-20
C24265 a_13259_45724# a_14127_45572# 2.92e-19
C24266 a_n2956_39304# en_comp 8.4e-19
C24267 a_n2956_38680# a_n2956_37592# 0.047258f
C24268 a_8199_44636# a_9482_43914# 0.276776f
C24269 a_584_46384# a_n881_46662# 0.286501f
C24270 a_2063_45854# a_n1613_43370# 0.04116f
C24271 a_2952_47436# a_3094_47243# 0.005572f
C24272 a_n3565_39590# a_n4334_37440# 3.56e-19
C24273 a_3785_47178# a_3315_47570# 2.31e-21
C24274 a_n1151_42308# a_2583_47243# 1.83e-19
C24275 a_16241_47178# a_16588_47582# 0.051162f
C24276 a_20712_42282# CAL_N 0.001755f
C24277 a_n4209_39590# a_n3690_37440# 1.67e-19
C24278 a_15811_47375# a_10227_46804# 0.019973f
C24279 a_11599_46634# a_18479_47436# 0.005025f
C24280 a_15673_47210# a_17591_47464# 1.51e-19
C24281 a_5742_30871# C1_N_btm 0.026156f
C24282 a_13717_47436# a_20894_47436# 6.95e-20
C24283 a_5932_42308# VIN_P 0.023512f
C24284 a_16327_47482# a_16763_47508# 0.338544f
C24285 a_8685_42308# VDD 0.286875f
C24286 a_13258_32519# a_22469_40625# 6.65e-19
C24287 a_5891_43370# a_9061_43230# 7.06e-20
C24288 a_n4318_40392# a_n3674_37592# 0.032206f
C24289 a_n97_42460# a_458_43396# 0.013064f
C24290 a_11967_42832# a_15279_43071# 0.027468f
C24291 a_19721_31679# a_n1630_35242# 1.04e-19
C24292 a_n2956_37592# a_n3690_39392# 1.91e-20
C24293 en_comp a_n3565_39304# 2.05e-19
C24294 a_6194_45824# VDD 0.274689f
C24295 a_n2810_45028# a_n3420_39072# 6.67e-21
C24296 a_3090_45724# a_15493_43940# 0.255251f
C24297 a_11453_44696# a_16243_43396# 1.19e-21
C24298 a_20623_45572# a_2437_43646# 2e-20
C24299 a_21363_45546# a_21513_45002# 0.06363f
C24300 a_20528_45572# a_20719_45572# 4.61e-19
C24301 a_12861_44030# a_21487_43396# 7.46e-20
C24302 a_526_44458# a_5891_43370# 1.12739f
C24303 a_8049_45260# a_18989_43940# 6.26e-20
C24304 a_n2293_46098# a_n809_44244# 1.32e-20
C24305 a_16327_47482# a_16823_43084# 0.535969f
C24306 a_19692_46634# a_15493_43396# 0.001909f
C24307 a_20107_45572# a_3357_43084# 0.308463f
C24308 a_20273_45572# a_19479_31679# 4.39e-20
C24309 a_10227_46804# a_15868_43402# 2.96e-20
C24310 a_15599_45572# a_6171_45002# 0.001026f
C24311 a_13925_46122# a_14673_44172# 2.92e-21
C24312 a_10809_44734# a_11649_44734# 2.53e-19
C24313 a_6945_45028# a_n2661_43922# 1.07e-19
C24314 a_7227_45028# a_n2661_43370# 0.026158f
C24315 C1_P_btm C3_N_btm 5.97e-19
C24316 C3_P_btm C5_N_btm 2.12e-19
C24317 a_15811_47375# a_17339_46660# 8.97e-20
C24318 a_n2497_47436# a_3147_46376# 7.92e-21
C24319 a_n1741_47186# a_167_45260# 4.69e-20
C24320 a_n2109_47186# a_2698_46116# 5.63e-21
C24321 a_15507_47210# a_765_45546# 0.00763f
C24322 a_2107_46812# a_4651_46660# 0.003567f
C24323 a_2063_45854# a_n2293_46098# 0.994164f
C24324 a_n881_46662# a_11901_46660# 1.99e-19
C24325 a_10227_46804# a_13059_46348# 0.656528f
C24326 a_16588_47582# a_16721_46634# 0.001918f
C24327 a_17591_47464# a_16388_46812# 2.32e-20
C24328 C10_P_btm VDD 2.40001f
C24329 C0_dummy_N_btm C0_N_btm 7.61701f
C24330 C0_dummy_P_btm C1_N_btm 2.22e-19
C24331 a_13717_47436# a_20411_46873# 1.46e-20
C24332 a_n746_45260# a_805_46414# 1.34e-19
C24333 a_n785_47204# a_n1076_46494# 9.42e-21
C24334 a_n237_47217# a_472_46348# 3.2e-19
C24335 a_5807_45002# a_6755_46942# 1.47519f
C24336 a_n2661_46634# a_7715_46873# 0.007284f
C24337 a_n1925_46634# a_3878_46660# 3.71e-19
C24338 a_2443_46660# a_2864_46660# 0.090164f
C24339 a_2609_46660# a_3524_46660# 0.118759f
C24340 a_n2661_42282# a_5267_42460# 2.34e-19
C24341 a_16855_43396# a_16823_43084# 0.005656f
C24342 a_8685_43396# a_7871_42858# 0.004749f
C24343 a_3626_43646# a_17701_42308# 0.003224f
C24344 a_2982_43646# a_17333_42852# 3.68e-20
C24345 a_17324_43396# a_5649_42852# 1.08e-21
C24346 a_19268_43646# a_19095_43396# 0.032587f
C24347 a_15743_43084# a_13467_32519# 0.02051f
C24348 a_18783_43370# a_4361_42308# 7.79e-21
C24349 a_3422_30871# a_17124_42282# 6.32e-20
C24350 a_15599_45572# a_14673_44172# 9.73e-20
C24351 a_2382_45260# a_2779_44458# 1.06e-19
C24352 a_n357_42282# a_10405_44172# 2.3e-20
C24353 a_3065_45002# a_742_44458# 2.17e-20
C24354 a_n913_45002# a_8975_43940# 4.06e-21
C24355 a_2324_44458# a_4093_43548# 1.63e-20
C24356 a_13348_45260# a_11691_44458# 2.44e-20
C24357 a_5009_45028# a_n2661_43370# 0.003943f
C24358 a_n2293_42834# a_8560_45348# 3.09e-20
C24359 a_5907_45546# a_5663_43940# 2.08e-20
C24360 a_3232_43370# a_n2661_44458# 0.468391f
C24361 a_n743_46660# a_2981_46116# 0.003499f
C24362 a_n2438_43548# a_1431_46436# 4.38e-20
C24363 a_5807_45002# a_8049_45260# 1.37423f
C24364 a_n1741_47186# a_12791_45546# 1.89e-19
C24365 a_n1925_46634# a_n1925_42282# 1.31e-19
C24366 a_12891_46348# a_12379_46436# 0.006296f
C24367 a_7927_46660# a_7920_46348# 3.44e-19
C24368 a_7577_46660# a_8349_46414# 0.001417f
C24369 a_7715_46873# a_8199_44636# 2.07e-21
C24370 a_n443_46116# a_3775_45552# 9.26e-22
C24371 a_6151_47436# a_6511_45714# 0.3215f
C24372 a_6545_47178# a_6472_45840# 6.79e-20
C24373 a_2063_45854# a_7230_45938# 0.016263f
C24374 a_4915_47217# a_7227_45028# 4.56e-21
C24375 a_19692_46634# a_18900_46660# 5.55e-20
C24376 a_3090_45724# a_12741_44636# 0.093609f
C24377 a_15559_46634# a_11415_45002# 1.37e-20
C24378 a_9067_47204# a_2711_45572# 1.64e-21
C24379 a_7411_46660# a_5937_45572# 2.28e-21
C24380 a_12895_43230# a_12800_43218# 0.049827f
C24381 a_13113_42826# a_12991_43230# 3.16e-19
C24382 a_12379_42858# a_13569_43230# 2.56e-19
C24383 a_19237_31679# RST_Z 0.050685f
C24384 a_13467_32519# a_1606_42308# 0.002946f
C24385 a_n1991_42858# COMP_P 1.96e-19
C24386 a_n4318_38680# a_n3674_38680# 3.04229f
C24387 a_14358_43442# a_14113_42308# 7.16e-21
C24388 a_12281_43396# a_11551_42558# 0.007065f
C24389 a_14579_43548# a_15051_42282# 0.002402f
C24390 a_n1641_43230# a_n1736_42282# 3.46e-19
C24391 a_n2840_43914# VDD 0.304745f
C24392 a_743_42282# a_n327_42308# 5.05e-21
C24393 a_n4318_39304# a_n4064_39072# 0.017224f
C24394 a_8953_45546# a_9114_42852# 1.98e-19
C24395 a_10180_45724# a_10695_43548# 1.07e-21
C24396 a_3090_45724# a_5742_30871# 7.9e-19
C24397 a_10775_45002# a_10807_43548# 1.41e-19
C24398 a_21005_45260# a_19279_43940# 4.39e-21
C24399 a_21101_45002# a_20766_44850# 0.01337f
C24400 a_21359_45002# a_20835_44721# 2.3e-19
C24401 a_20193_45348# a_11967_42832# 0.01602f
C24402 a_11691_44458# a_19615_44636# 0.001633f
C24403 a_11827_44484# a_20679_44626# 0.030022f
C24404 a_2711_45572# a_16759_43396# 6.88e-21
C24405 a_n1741_47186# DATA[4] 0.020035f
C24406 a_8746_45002# a_9145_43396# 1.83e-20
C24407 a_n785_47204# VDD 0.452945f
C24408 a_13720_44458# a_9313_44734# 1.1e-21
C24409 a_10951_45334# a_10949_43914# 8.94e-19
C24410 a_11787_45002# a_10729_43914# 3.79e-21
C24411 a_18114_32519# a_17517_44484# 0.055077f
C24412 a_18184_42460# a_18579_44172# 0.161593f
C24413 a_n755_45592# a_743_42282# 0.160592f
C24414 a_n357_42282# a_20556_43646# 4.02e-19
C24415 a_n2293_42834# a_453_43940# 1.92e-20
C24416 a_n356_44636# a_7_44811# 0.005265f
C24417 a_8103_44636# a_n2661_43922# 0.008682f
C24418 a_n2293_45010# a_726_44056# 8.78e-19
C24419 a_n452_47436# DATA[0] 0.039965f
C24420 a_n2312_38680# a_n3565_38502# 0.134976f
C24421 a_9290_44172# a_9061_43230# 2.91e-21
C24422 a_9290_44172# a_526_44458# 0.200352f
C24423 a_8016_46348# a_5066_45546# 0.054471f
C24424 a_6755_46942# a_15143_45578# 2.33e-21
C24425 a_4791_45118# a_5837_45028# 5.56e-20
C24426 a_n881_46662# a_n659_45366# 8.3e-19
C24427 a_10227_46804# a_13556_45296# 0.013693f
C24428 a_10384_47026# a_8746_45002# 5.86e-21
C24429 a_11453_44696# a_3232_43370# 0.132496f
C24430 a_18819_46122# a_20708_46348# 2.33e-20
C24431 a_18985_46122# a_19900_46494# 0.118759f
C24432 a_18189_46348# a_6945_45028# 4.84e-20
C24433 a_15811_47375# a_1307_43914# 1.46e-19
C24434 a_13747_46662# a_2437_43646# 0.008951f
C24435 a_3090_45724# a_3260_45572# 6.23e-19
C24436 a_6419_46155# a_6640_46482# 0.007833f
C24437 a_17583_46090# a_10809_44734# 2.89e-21
C24438 a_1576_42282# a_5934_30871# 2.52e-20
C24439 a_5342_30871# a_n3420_38528# 0.028503f
C24440 a_961_42354# a_6123_31319# 1.52e-20
C24441 a_3823_42558# a_3581_42558# 3.68e-20
C24442 a_5534_30871# a_n4064_38528# 0.057361f
C24443 a_n784_42308# a_8685_42308# 1.58e-20
C24444 a_2123_42473# a_5932_42308# 4.34e-21
C24445 a_1755_42282# a_6481_42558# 0.012532f
C24446 a_9803_43646# VDD 0.261557f
C24447 a_n357_42282# a_6171_42473# 0.010166f
C24448 a_n755_45592# a_5755_42308# 3.68e-19
C24449 a_14815_43914# a_15493_43940# 8.51e-20
C24450 a_n2661_42834# a_11816_44260# 1.53e-19
C24451 a_n984_44318# a_895_43940# 2.65e-20
C24452 a_1115_44172# a_453_43940# 0.150214f
C24453 a_17517_44484# a_17737_43940# 9.06e-20
C24454 a_14537_43396# a_16823_43084# 9.22e-21
C24455 a_18248_44752# a_19319_43548# 1.93e-20
C24456 a_6298_44484# a_n97_42460# 5.4e-19
C24457 a_1467_44172# a_1414_42308# 0.335735f
C24458 a_n913_45002# a_2905_42968# 0.009485f
C24459 a_n1059_45260# a_3681_42891# 0.003573f
C24460 a_n2017_45002# a_3935_42891# 4.3e-21
C24461 a_742_44458# a_458_43396# 4.92e-20
C24462 a_13259_45724# a_14456_42282# 5.4e-19
C24463 a_1848_45724# a_n443_42852# 5.35e-20
C24464 a_n356_45724# a_n310_45899# 0.006879f
C24465 a_2107_46812# a_8975_43940# 0.075583f
C24466 a_n2661_45546# a_3175_45822# 2.16e-19
C24467 a_13059_46348# a_1307_43914# 0.04241f
C24468 a_584_46384# a_2889_44172# 4.84e-20
C24469 a_18597_46090# a_19006_44850# 3.17e-20
C24470 a_16327_47482# a_19279_43940# 0.446333f
C24471 a_n1099_45572# a_n310_45572# 2.46e-19
C24472 a_8049_45260# a_15143_45578# 0.001756f
C24473 a_n2497_47436# a_n1441_43940# 0.004491f
C24474 a_3090_45724# a_n2293_42834# 0.023056f
C24475 a_n971_45724# a_7542_44172# 4.49e-21
C24476 a_3483_46348# a_3357_43084# 0.030022f
C24477 a_n1613_43370# a_n2661_42834# 0.112184f
C24478 a_4419_46090# a_2437_43646# 3.77e-20
C24479 a_12861_44030# a_21398_44850# 2.74e-20
C24480 a_1138_42852# a_n2661_45010# 0.017849f
C24481 a_n1076_46494# a_n913_45002# 8.43e-20
C24482 a_n901_46420# a_n745_45366# 7.11e-19
C24483 a_n1853_46287# a_n967_45348# 3.76e-21
C24484 a_17715_44484# a_16842_45938# 4.81e-20
C24485 a_12549_44172# a_9313_44734# 3.97e-19
C24486 a_10809_44734# a_8696_44636# 0.117876f
C24487 a_6945_45028# a_17478_45572# 2.17e-21
C24488 a_10586_45546# a_12791_45546# 9.22e-21
C24489 a_n863_45724# a_603_45572# 3.59e-21
C24490 a_n755_45592# a_2277_45546# 0.065177f
C24491 a_n2302_39866# a_n2216_39866# 0.011479f
C24492 a_n3420_39616# a_n4251_39616# 0.0016f
C24493 a_584_46384# a_n443_46116# 0.496286f
C24494 a_n971_45724# a_6575_47204# 0.01923f
C24495 a_n1151_42308# a_3381_47502# 0.051194f
C24496 a_2905_45572# a_3815_47204# 0.00535f
C24497 a_2063_45854# a_4791_45118# 0.039758f
C24498 a_n237_47217# a_7227_47204# 0.013654f
C24499 a_n1741_47186# a_11459_47204# 0.015445f
C24500 a_3160_47472# a_3785_47178# 2.34e-19
C24501 a_n2109_47186# a_n1435_47204# 0.041807f
C24502 a_n3690_39616# a_n3607_39616# 0.007692f
C24503 a_n4064_40160# a_n2946_39072# 2.04e-20
C24504 a_4958_30871# a_n3420_37984# 0.031033f
C24505 a_14097_32519# C6_N_btm 8.47e-20
C24506 a_n1630_35242# a_18194_35068# 0.465356f
C24507 a_5742_30871# a_3754_38470# 1.66e-19
C24508 a_n784_42308# C10_P_btm 1.34e-19
C24509 a_n4315_30879# a_n2302_39072# 6.48e-20
C24510 a_n4334_39616# a_n4209_39304# 3.3e-19
C24511 a_n4209_39590# a_n4334_39392# 3.3e-19
C24512 a_14539_43914# a_17333_42852# 0.072085f
C24513 en_comp a_14113_42308# 3.72e-20
C24514 a_19615_44636# a_4190_30871# 1.28e-21
C24515 a_22315_44484# a_15743_43084# 2.11e-21
C24516 a_n356_44636# a_13113_42826# 5.02e-21
C24517 a_1307_43914# a_2903_42308# 6.88e-22
C24518 a_5111_44636# a_9223_42460# 1.34e-20
C24519 a_n1059_45260# a_15959_42545# 0.002635f
C24520 a_n2017_45002# a_15890_42674# 0.00307f
C24521 a_n913_45002# a_15803_42450# 8.35e-19
C24522 a_8375_44464# a_8387_43230# 6.17e-22
C24523 a_5891_43370# a_8605_42826# 0.0011f
C24524 a_742_44458# a_2987_42968# 7.44e-19
C24525 a_n2661_42282# a_6547_43396# 0.00581f
C24526 a_n2293_42834# a_n2472_42282# 0.002489f
C24527 a_13661_43548# a_13565_43940# 0.017205f
C24528 a_n755_45592# a_626_44172# 0.100613f
C24529 a_n863_45724# a_2903_45348# 1.21e-20
C24530 a_n357_42282# a_1145_45348# 1.17e-20
C24531 a_12549_44172# a_20974_43370# 0.061866f
C24532 a_2711_45572# a_7276_45260# 0.00282f
C24533 a_8049_45260# a_18315_45260# 1.23e-20
C24534 a_7499_43078# en_comp 8.68e-21
C24535 a_10193_42453# a_n913_45002# 0.562004f
C24536 a_n1613_43370# a_n1352_43396# 0.244933f
C24537 a_4915_47217# a_14205_43396# 8.72e-21
C24538 a_13351_46090# a_13076_44458# 3.69e-21
C24539 a_2324_44458# a_10157_44484# 2.29e-21
C24540 a_5907_45546# a_3232_43370# 0.001196f
C24541 a_6194_45824# a_5691_45260# 1.08e-19
C24542 a_3775_45552# a_3537_45260# 1.46e-19
C24543 a_3483_46348# a_5826_44734# 8.07e-19
C24544 a_3218_45724# a_1307_43914# 6.18e-21
C24545 a_8696_44636# a_16211_45572# 2.41e-20
C24546 a_16115_45572# a_16147_45260# 6.95e-19
C24547 a_n2472_46090# a_n2661_43922# 5.03e-21
C24548 a_n2293_46098# a_n2661_42834# 0.029385f
C24549 a_12741_44636# a_14815_43914# 0.003697f
C24550 a_6886_37412# a_n923_35174# 0.003125f
C24551 a_n3565_37414# C5_P_btm 1.11e-20
C24552 a_n3420_37440# C7_P_btm 1.33e-20
C24553 a_11599_46634# a_10554_47026# 7.33e-21
C24554 a_20843_47204# a_21588_30879# 1e-19
C24555 a_3754_39466# VDD 0.009313f
C24556 a_14311_47204# a_6755_46942# 1.38e-20
C24557 a_7754_39632# RST_Z 0.030938f
C24558 a_n4064_37984# VREF 3.68e-19
C24559 a_n881_46662# a_479_46660# 3.54e-19
C24560 a_4915_47217# a_11813_46116# 1.35e-19
C24561 a_n1151_42308# a_15009_46634# 8.05e-19
C24562 a_6575_47204# a_8023_46660# 1.23e-19
C24563 a_9313_45822# a_8035_47026# 1.13e-19
C24564 a_6151_47436# a_10768_47026# 8.29e-20
C24565 a_n3420_37984# VCM 0.014539f
C24566 a_4883_46098# a_5732_46660# 3.05e-22
C24567 CAL_N a_22717_37285# 7.87e-21
C24568 a_22521_39511# a_22780_39857# 0.01318f
C24569 a_22469_40625# a_22609_37990# 0.130478f
C24570 a_22521_40055# a_22609_38406# 0.1922f
C24571 a_22521_40599# a_22705_37990# 1.29e-19
C24572 a_22459_39145# CAL_P 0.005678f
C24573 a_22545_38993# a_22469_39537# 0.049703f
C24574 a_n1613_43370# a_645_46660# 0.001903f
C24575 a_19479_31679# VREF 0.056254f
C24576 a_n1331_43914# COMP_P 5.76e-20
C24577 a_9145_43396# a_16243_43396# 2.75e-21
C24578 a_3626_43646# a_4361_42308# 5.20633f
C24579 a_10341_43396# a_9885_43396# 9.63e-20
C24580 a_n1761_44111# a_n961_42308# 0.002207f
C24581 a_n356_44636# a_18214_42558# 5.42e-19
C24582 a_n913_45002# VDD 9.190901f
C24583 a_n1059_45260# RST_Z 3.96e-20
C24584 a_14205_43396# a_15681_43442# 3.24e-20
C24585 a_12293_43646# a_12281_43396# 0.01129f
C24586 a_14021_43940# a_21356_42826# 6.95e-20
C24587 a_2982_43646# a_13678_32519# 2.63e-21
C24588 a_13667_43396# a_13837_43396# 0.001675f
C24589 a_3232_43370# a_6125_45348# 0.001449f
C24590 a_6171_45002# a_5837_45348# 9.51e-21
C24591 a_3537_45260# a_5093_45028# 0.009279f
C24592 a_20273_45572# a_20193_45348# 5.61e-19
C24593 a_6755_46942# a_16867_43762# 2.42e-19
C24594 a_12549_44172# a_18599_43230# 3.17e-20
C24595 a_n1613_43370# a_n2293_42282# 6.65e-20
C24596 a_14537_43396# a_15415_45028# 4.17e-20
C24597 a_8696_44636# a_5883_43914# 0.004598f
C24598 a_n967_45348# a_n2661_43370# 0.016831f
C24599 a_10227_46804# a_11554_42852# 2.46e-19
C24600 a_n971_45724# a_n1630_35242# 0.028303f
C24601 a_5937_45572# a_5829_43940# 0.006959f
C24602 a_13556_45296# a_1307_43914# 0.007672f
C24603 a_n2293_46634# a_10083_42826# 6.79e-20
C24604 a_13661_43548# a_5534_30871# 4.79e-20
C24605 a_21513_45002# a_19778_44110# 1.82e-19
C24606 a_7499_43078# a_10617_44484# 5.41e-19
C24607 a_n1925_46634# a_2698_46116# 8.92e-20
C24608 a_n2661_46098# a_n2840_46090# 0.170439f
C24609 a_5807_45002# a_8953_45546# 0.00249f
C24610 a_11459_47204# a_10586_45546# 1.75e-22
C24611 a_14084_46812# a_15009_46634# 4.66e-19
C24612 a_n2661_46634# a_4419_46090# 1.65e-19
C24613 a_n2293_46634# a_3483_46348# 0.157275f
C24614 a_7715_46873# a_765_45546# 0.001838f
C24615 a_n881_46662# a_17583_46090# 0.003148f
C24616 a_12891_46348# a_13351_46090# 0.019821f
C24617 a_12549_44172# a_12594_46348# 0.031894f
C24618 a_n743_46660# a_167_45260# 0.045398f
C24619 a_1123_46634# a_472_46348# 0.001483f
C24620 a_33_46660# a_1176_45822# 5.48e-19
C24621 a_383_46660# a_805_46414# 0.01072f
C24622 a_n971_45724# a_n2661_45546# 0.083094f
C24623 a_n2497_47436# a_310_45028# 4.48e-20
C24624 a_14311_47204# a_8049_45260# 4.71e-21
C24625 a_n2312_39304# a_n2956_38680# 0.048558f
C24626 a_16759_43396# a_16877_42852# 6.34e-20
C24627 a_15743_43084# a_18695_43230# 5.34e-19
C24628 a_3422_30871# VDAC_P 0.476038f
C24629 a_n97_42460# a_13575_42558# 0.179828f
C24630 a_3626_43646# a_6761_42308# 0.006571f
C24631 a_2982_43646# a_6123_31319# 0.163265f
C24632 a_12089_42308# a_12545_42858# 0.261463f
C24633 a_12379_42858# a_13113_42826# 0.06628f
C24634 a_5649_42852# a_5193_42852# 0.003625f
C24635 a_556_44484# VDD 0.004463f
C24636 a_13661_43548# a_19647_42308# 5.53e-21
C24637 a_20193_45348# a_18989_43940# 4.63e-22
C24638 a_n755_45592# a_2813_43396# 6.23e-21
C24639 a_413_45260# a_453_43940# 5.59e-20
C24640 a_n2840_45002# a_n3674_39768# 0.00158f
C24641 a_9290_44172# a_8605_42826# 9.78e-21
C24642 a_n443_42852# a_1512_43396# 3.67e-19
C24643 a_n2661_44458# a_8975_43940# 0.075732f
C24644 a_n2312_39304# a_n3690_39392# 4.25e-19
C24645 a_n913_45002# a_5495_43940# 4.51e-22
C24646 a_18479_45785# a_19328_44172# 0.003851f
C24647 a_8953_45546# a_10518_42984# 9.33e-20
C24648 a_8199_44636# a_10796_42968# 1.77e-20
C24649 a_3483_46348# a_5342_30871# 8.76e-19
C24650 a_4185_45028# a_5534_30871# 0.05188f
C24651 a_4223_44672# a_4743_44484# 0.043867f
C24652 w_1575_34946# RST_Z 0.001495f
C24653 a_n2293_46634# a_14495_45572# 5.19e-21
C24654 a_11415_45002# a_21137_46414# 6.03e-22
C24655 a_20202_43084# a_6945_45028# 0.02248f
C24656 a_3483_46348# a_9625_46129# 0.038063f
C24657 a_22365_46825# a_22223_46124# 0.011912f
C24658 a_20885_46660# a_10809_44734# 3.49e-19
C24659 a_18597_46090# a_20107_45572# 0.069963f
C24660 a_11599_46634# a_2437_43646# 0.006609f
C24661 a_5167_46660# a_2711_45572# 1.79e-20
C24662 a_n237_47217# a_6171_45002# 1.47e-19
C24663 a_584_46384# a_3537_45260# 0.108506f
C24664 a_3785_47178# a_413_45260# 7.03e-19
C24665 a_n881_46662# a_8696_44636# 0.178516f
C24666 a_18479_47436# a_20841_45814# 0.011134f
C24667 a_16327_47482# a_19610_45572# 0.00341f
C24668 a_n743_46660# a_12791_45546# 6.76e-20
C24669 a_4646_46812# a_6194_45824# 9.75e-21
C24670 a_3877_44458# a_6472_45840# 2.74e-20
C24671 a_12741_44636# a_20075_46420# 0.027561f
C24672 a_n971_45724# a_5205_44484# 9.71e-22
C24673 a_12549_44172# a_15037_45618# 7.69e-21
C24674 a_768_44030# a_14033_45822# 0.005149f
C24675 a_3090_45724# a_16375_45002# 0.026416f
C24676 a_15559_46634# a_13259_45724# 9.61e-21
C24677 a_2063_45854# a_3429_45260# 6.96e-22
C24678 a_10227_46804# a_21363_45546# 3.24e-21
C24679 a_11453_44696# a_18341_45572# 0.026938f
C24680 a_13487_47204# a_3357_43084# 5.65e-19
C24681 a_7309_42852# a_7227_42308# 4.85e-19
C24682 a_22400_42852# COMP_P 0.614467f
C24683 a_n4318_39304# VDD 0.643395f
C24684 a_4190_30871# a_n4064_38528# 0.031783f
C24685 a_n2840_42282# a_n3674_38680# 0.154001f
C24686 a_5342_30871# a_15761_42308# 1e-19
C24687 a_3080_42308# C10_P_btm 1.34e-19
C24688 a_4185_45028# a_19647_42308# 1.64e-19
C24689 a_n2293_42834# a_n1821_43396# 7.71e-19
C24690 a_1307_43914# a_6293_42852# 2.54e-19
C24691 a_n356_44636# a_n2661_42282# 2.54767f
C24692 a_11967_42832# a_20596_44850# 2.49e-19
C24693 a_10193_42453# a_20922_43172# 0.059157f
C24694 a_2107_46812# VDD 0.350275f
C24695 a_16922_45042# a_19319_43548# 1.84e-20
C24696 a_n2661_43922# a_895_43940# 0.002919f
C24697 a_n2661_42834# a_2675_43914# 0.024352f
C24698 a_14539_43914# a_13483_43940# 8.72e-20
C24699 a_3232_43370# a_9145_43396# 1.89e-19
C24700 a_33_46660# DATA[0] 1.05e-20
C24701 a_n2661_43370# a_n1917_43396# 3.88e-20
C24702 a_n1059_45260# a_16243_43396# 0.012252f
C24703 a_n2017_45002# a_16547_43609# 8.08e-20
C24704 a_n913_45002# a_16137_43396# 3.32e-19
C24705 a_n743_46660# DATA[4] 1.69e-21
C24706 a_17517_44484# a_22485_44484# 0.110643f
C24707 a_20835_44721# a_19279_43940# 0.036128f
C24708 a_20362_44736# a_18579_44172# 6.86e-20
C24709 a_19321_45002# a_22223_45036# 5.03e-20
C24710 a_12549_44172# a_18114_32519# 0.001232f
C24711 a_15227_44166# en_comp 4.89e-21
C24712 a_18280_46660# a_18479_45785# 5.88e-20
C24713 a_18243_46436# a_18051_46116# 6.96e-20
C24714 a_19240_46482# a_19431_46494# 4.61e-19
C24715 a_5937_45572# a_6229_45572# 5.31e-19
C24716 a_11453_44696# a_8975_43940# 0.027482f
C24717 a_12465_44636# a_13720_44458# 0.019702f
C24718 a_2324_44458# a_7499_43078# 0.018394f
C24719 a_13661_43548# a_11691_44458# 0.263889f
C24720 a_5807_45002# a_20193_45348# 1.07e-19
C24721 a_13747_46662# a_19113_45348# 2.83e-19
C24722 a_3483_46348# a_9159_45572# 0.006021f
C24723 a_8270_45546# a_6171_45002# 0.027058f
C24724 a_4791_45118# a_n2661_42834# 0.024946f
C24725 a_3090_45724# a_413_45260# 0.135828f
C24726 a_10903_43370# a_11962_45724# 0.357882f
C24727 a_12594_46348# a_11525_45546# 2.4e-19
C24728 a_n743_46660# a_16405_45348# 7.86e-19
C24729 a_14513_46634# a_3357_43084# 2.21e-20
C24730 a_n1613_43370# a_n1352_44484# 0.232498f
C24731 a_17124_42282# a_7174_31319# 5.22e-20
C24732 a_5934_30871# a_1736_39043# 5.23e-20
C24733 a_20922_43172# VDD 0.192467f
C24734 a_18907_42674# a_19332_42282# 0.017308f
C24735 a_18057_42282# a_18220_42308# 0.01135f
C24736 a_18727_42674# a_18214_42558# 0.035505f
C24737 a_5534_30871# VREF_GND 0.060532f
C24738 a_5342_30871# VIN_N 0.00693f
C24739 a_19987_42826# RST_Z 8.97e-21
C24740 a_n2017_45002# a_n3674_37592# 0.241068f
C24741 a_2479_44172# a_n97_42460# 0.196935f
C24742 a_n356_44636# a_16823_43084# 0.003531f
C24743 a_n913_45002# a_n784_42308# 0.005856f
C24744 a_n1059_45260# a_n327_42558# 6.01e-20
C24745 a_9313_44734# a_16977_43638# 1.9e-20
C24746 en_comp a_n1329_42308# 5.94e-20
C24747 a_n967_45348# COMP_P 0.00202f
C24748 a_n2293_45010# a_n1630_35242# 1.46e-20
C24749 a_14493_46090# VDD 0.203567f
C24750 a_19328_44172# a_14021_43940# 1.77e-20
C24751 a_n2661_44458# a_2905_42968# 1.46e-21
C24752 a_13925_46122# RST_Z 4.05e-21
C24753 a_n1076_46494# a_n2661_44458# 3.36e-21
C24754 a_n2956_38216# a_n2661_45010# 0.005195f
C24755 a_n357_42282# a_3357_43084# 0.010127f
C24756 a_584_46384# a_1049_43396# 0.148494f
C24757 a_n1641_46494# a_n2129_44697# 1.53e-21
C24758 a_n1423_46090# a_n2267_44484# 5.61e-21
C24759 a_11962_45724# a_12016_45572# 0.002378f
C24760 a_11823_42460# a_11688_45572# 8.92e-20
C24761 a_10193_42453# a_15903_45785# 2.18e-20
C24762 a_n2438_43548# a_n1644_44306# 1.68e-20
C24763 a_1848_45724# a_2437_43646# 0.007112f
C24764 a_n2472_45546# a_n2472_45002# 0.026152f
C24765 a_n2661_45546# a_n2293_45010# 0.003149f
C24766 a_12549_44172# a_17737_43940# 0.007227f
C24767 a_8049_45260# a_13017_45260# 4.13e-20
C24768 a_2324_44458# a_11915_45394# 8.14e-19
C24769 a_7754_40130# a_4338_37500# 0.030623f
C24770 a_2747_46873# a_3411_47243# 6.35e-21
C24771 a_16327_47482# a_20916_46384# 3.47e-19
C24772 a_18780_47178# a_5807_45002# 1.88e-20
C24773 a_18479_47436# a_13661_43548# 0.024025f
C24774 a_6491_46660# a_2107_46812# 7.39e-21
C24775 a_n1435_47204# a_n1925_46634# 1.17e-19
C24776 a_7754_38636# a_3754_38470# 0.037604f
C24777 a_n4334_40480# VDD 0.390668f
C24778 a_n4209_39304# C5_P_btm 1.83e-19
C24779 a_17591_47464# a_19321_45002# 6.33e-21
C24780 a_18143_47464# a_13747_46662# 3.2e-19
C24781 a_3160_47472# a_3699_46634# 7.39e-19
C24782 a_3381_47502# a_3177_46902# 2.56e-19
C24783 a_n1151_42308# a_2959_46660# 3.22e-19
C24784 a_2905_45572# a_3524_46660# 0.011982f
C24785 a_584_46384# a_1302_46660# 5.41e-21
C24786 a_13258_32519# VREF 9.37e-19
C24787 a_11459_47204# a_n743_46660# 3.96e-21
C24788 a_n443_46116# a_479_46660# 1.72e-19
C24789 a_n971_45724# a_5385_46902# 5.88e-20
C24790 a_n237_47217# a_4955_46873# 0.032268f
C24791 a_n4209_38502# a_n1386_35608# 1.52e-19
C24792 a_11599_46634# a_n2661_46634# 0.067552f
C24793 a_12465_44636# a_12549_44172# 0.093222f
C24794 a_n3420_39072# C9_P_btm 5.77e-20
C24795 a_n3565_39304# C7_P_btm 0.001136f
C24796 a_18494_42460# a_18220_42308# 7.47e-19
C24797 a_n2956_37592# a_n3420_37440# 0.233174f
C24798 a_15903_45785# VDD 0.291109f
C24799 a_19479_31679# a_22521_40599# 1.54e-20
C24800 a_9672_43914# a_10083_42826# 8.52e-20
C24801 a_n2810_45028# a_n2946_37690# 0.024678f
C24802 a_n2661_42834# a_n1736_42282# 6.4e-21
C24803 a_n2293_43922# a_n2104_42282# 0.009285f
C24804 a_11967_42832# a_15785_43172# 0.003242f
C24805 a_19319_43548# a_15743_43084# 0.035611f
C24806 a_18533_43940# a_18783_43370# 0.00197f
C24807 a_6547_43396# a_7112_43396# 7.99e-20
C24808 a_6031_43396# a_6452_43396# 0.086708f
C24809 a_10227_46804# a_10991_42826# 0.152133f
C24810 a_21076_30879# a_15493_43940# 1.4e-20
C24811 a_2711_45572# a_13720_44458# 0.001214f
C24812 a_10193_42453# a_n2661_44458# 3e-19
C24813 a_n1059_45260# a_3232_43370# 1.26e-19
C24814 a_n1613_43370# a_n1423_42826# 0.15981f
C24815 a_n23_45546# a_n23_44458# 6.98e-19
C24816 a_413_45260# a_2274_45254# 0.002353f
C24817 a_3483_46348# a_9672_43914# 0.125466f
C24818 a_12861_44030# a_15567_42826# 0.004897f
C24819 a_13661_43548# a_4190_30871# 0.147163f
C24820 a_n2109_47186# a_526_44458# 4.75e-20
C24821 a_2063_45854# a_6945_45028# 0.074119f
C24822 a_5807_45002# a_18285_46348# 0.006196f
C24823 a_11459_47204# a_11189_46129# 7.59e-19
C24824 a_13747_46662# a_765_45546# 7.33e-19
C24825 a_2609_46660# a_3090_45724# 2.67e-20
C24826 a_18429_43548# a_18083_42858# 1.96e-19
C24827 a_743_42282# a_10083_42826# 2.64e-19
C24828 a_15743_43084# a_16795_42852# 5.64e-20
C24829 a_n3674_39304# a_n1736_43218# 3.4e-21
C24830 a_10555_44260# a_10533_42308# 3.68e-22
C24831 a_15493_43396# a_15486_42560# 2.06e-19
C24832 a_n1423_42826# a_n1533_42852# 0.097745f
C24833 a_n2661_44458# VDD 1.06317f
C24834 a_4361_42308# a_8037_42858# 1.08e-19
C24835 a_18494_42460# a_11827_44484# 0.031498f
C24836 a_3065_45002# a_n2661_43922# 0.023551f
C24837 a_10193_42453# a_18451_43940# 0.20167f
C24838 a_13059_46348# a_13635_43156# 3.86e-20
C24839 a_19692_46634# a_21356_42826# 5.5e-20
C24840 a_n2661_43370# a_n1917_44484# 0.002293f
C24841 a_16922_45042# a_17801_45144# 0.005123f
C24842 a_17023_45118# a_16981_45144# 7.47e-21
C24843 a_5147_45002# a_5708_44484# 0.055267f
C24844 a_5111_44636# a_5608_44484# 0.002582f
C24845 a_3483_46348# a_743_42282# 2.47e-22
C24846 a_n2293_42834# a_4743_44484# 7.24e-21
C24847 a_8953_45002# a_5891_43370# 4.12e-19
C24848 a_18587_45118# a_11691_44458# 3.11e-20
C24849 a_21005_45260# a_21101_45002# 0.419086f
C24850 a_18911_45144# a_19113_45348# 0.054737f
C24851 a_11823_42460# a_12429_44172# 0.018664f
C24852 a_n2017_45002# a_14673_44172# 8.16e-21
C24853 a_12861_44030# a_20712_42282# 7.11e-22
C24854 a_2324_44458# a_15781_43660# 4.8e-19
C24855 a_768_44030# a_5934_30871# 3.24e-23
C24856 a_4185_45028# a_4190_30871# 0.16524f
C24857 a_10227_46804# a_17303_42282# 8.27e-21
C24858 a_16327_47482# a_19332_42282# 6.14e-19
C24859 a_4883_46098# a_11962_45724# 9.92e-21
C24860 a_n2661_46634# a_1848_45724# 2.19e-20
C24861 a_13661_43548# a_n443_42852# 0.045364f
C24862 a_n881_46662# a_7227_45028# 5.19e-19
C24863 a_n1613_43370# a_3775_45552# 1.56e-20
C24864 a_11453_44696# a_10193_42453# 0.071253f
C24865 a_13507_46334# a_11823_42460# 1.48e-19
C24866 a_n133_46660# a_n2293_45546# 1.48e-22
C24867 a_7577_46660# a_8034_45724# 1.64e-20
C24868 a_12549_44172# a_2711_45572# 2.05236f
C24869 a_15227_44166# a_2324_44458# 0.190521f
C24870 a_17609_46634# a_17583_46090# 0.008733f
C24871 a_12741_44636# a_21076_30879# 0.00607f
C24872 a_765_45546# a_4419_46090# 8e-20
C24873 a_11813_46116# a_10809_44734# 0.001353f
C24874 a_3090_45724# a_18985_46122# 1.47e-19
C24875 a_n2293_46634# a_n357_42282# 0.034749f
C24876 a_n743_46660# a_n863_45724# 0.007504f
C24877 a_3080_42308# a_3754_39466# 2.89e-20
C24878 a_18451_43940# VDD 0.172318f
C24879 a_15743_43084# a_21335_42336# 3.06e-20
C24880 a_4361_42308# a_13921_42308# 3.34e-19
C24881 a_n2293_42282# a_n1736_42282# 4.89e-19
C24882 a_7871_42858# a_6123_31319# 0.010286f
C24883 a_21588_30879# a_22521_39511# 7.63e-20
C24884 a_n357_42282# a_5342_30871# 0.039779f
C24885 a_17339_46660# a_17303_42282# 9.87e-21
C24886 a_n143_45144# a_n229_43646# 1.73e-21
C24887 a_22223_47212# SINGLE_ENDED 6.55e-19
C24888 a_n699_43396# a_1467_44172# 0.030347f
C24889 a_4223_44672# a_1414_42308# 2.93e-20
C24890 a_n913_45002# a_3080_42308# 0.044741f
C24891 a_n1059_45260# a_4905_42826# 0.027099f
C24892 a_1823_45246# a_6123_31319# 3.21e-20
C24893 a_1307_43914# a_7499_43940# 0.005916f
C24894 a_949_44458# a_2127_44172# 0.006932f
C24895 a_n2661_44458# a_5495_43940# 1.41e-20
C24896 a_742_44458# a_2479_44172# 0.019563f
C24897 a_13857_44734# a_14112_44734# 0.005172f
C24898 a_11649_44734# a_11541_44484# 5.37e-19
C24899 SMPL_ON_N RST_Z 2.43362f
C24900 a_4185_45028# a_5337_42558# 3.05e-19
C24901 a_n443_42852# a_10835_43094# 1.88e-19
C24902 a_11453_44696# VDD 3.75355f
C24903 a_2107_46812# a_5691_45260# 1.52e-20
C24904 a_n743_46660# a_8191_45002# 6.12e-22
C24905 a_4185_45028# a_n443_42852# 0.027973f
C24906 a_1138_42852# a_1260_45572# 0.001766f
C24907 a_n1151_42308# a_n699_43396# 0.022019f
C24908 a_19335_46494# a_19240_46482# 0.049827f
C24909 a_19553_46090# a_19431_46494# 3.16e-19
C24910 a_8953_45546# a_n755_45592# 3.44e-19
C24911 a_n2293_46098# a_3775_45552# 0.003338f
C24912 a_3699_46634# a_413_45260# 3.59e-20
C24913 a_15227_44166# a_16855_45546# 8.57e-19
C24914 a_4646_46812# a_n913_45002# 7.74e-20
C24915 a_15368_46634# a_16020_45572# 5.92e-20
C24916 a_7411_46660# a_2437_43646# 7.33e-20
C24917 a_2443_46660# a_2382_45260# 8.11e-22
C24918 a_16327_47482# a_21101_45002# 1.72e-19
C24919 a_17364_32525# VDD 0.511443f
C24920 a_5934_30871# a_10149_42308# 4.13e-20
C24921 a_n4318_37592# a_n4334_39616# 7.61e-20
C24922 COMP_P a_n4209_39590# 0.010869f
C24923 a_5342_30871# CAL_N 0.004302f
C24924 a_4190_30871# VREF_GND 0.105109f
C24925 a_22959_43396# RST_Z 0.001326f
C24926 a_1755_42282# a_7174_31319# 1.94e-20
C24927 a_20731_47026# SINGLE_ENDED 1.3e-20
C24928 a_5891_43370# a_3626_43646# 0.00315f
C24929 a_n2293_42834# a_n1736_43218# 0.005982f
C24930 a_1307_43914# a_10991_42826# 1.82e-20
C24931 a_2382_45260# a_4156_43218# 6.43e-19
C24932 a_10193_42453# a_8325_42308# 3.66e-20
C24933 a_8975_43940# a_9145_43396# 1.06e-19
C24934 a_10057_43914# a_9803_43646# 0.001251f
C24935 a_n357_42282# a_20107_42308# 5.18e-19
C24936 a_17517_44484# a_14401_32519# 8.5e-19
C24937 a_n2661_42834# a_1209_43370# 2.79e-20
C24938 a_17639_46660# VDD 0.001662f
C24939 a_7499_43078# a_9803_42558# 0.158876f
C24940 a_13556_45296# a_13635_43156# 8.03e-21
C24941 a_9482_43914# a_13460_43230# 1.07e-20
C24942 a_1423_45028# a_9127_43156# 2.04e-20
C24943 a_2804_46116# a_1423_45028# 1.3e-21
C24944 a_1823_45246# a_3495_45348# 2.54e-19
C24945 a_2324_44458# a_4558_45348# 9.57e-20
C24946 a_9290_44172# a_8953_45002# 0.002181f
C24947 a_n2293_46098# a_5093_45028# 0.00251f
C24948 a_3090_45724# a_2779_44458# 5.81e-20
C24949 a_n2956_38680# a_n2810_45028# 0.043221f
C24950 a_12549_44172# a_22485_44484# 2.07e-20
C24951 a_n1613_43370# a_n1549_44318# 0.16289f
C24952 a_7227_45028# a_8162_45546# 0.003048f
C24953 a_13759_46122# a_6171_45002# 4.55e-20
C24954 a_6667_45809# a_7499_43078# 2.77e-21
C24955 a_20075_46420# a_413_45260# 4.37e-21
C24956 a_13661_43548# a_18753_44484# 0.00166f
C24957 a_8049_45260# a_20107_45572# 0.024509f
C24958 a_18285_46348# a_18315_45260# 5.03e-22
C24959 a_20411_46873# a_16922_45042# 1.1e-20
C24960 a_13259_45724# a_14033_45572# 2.45e-19
C24961 a_n2956_39304# a_n2956_37592# 0.044994f
C24962 a_2711_45572# a_11525_45546# 0.0154f
C24963 a_2063_45854# a_11173_44260# 0.00917f
C24964 a_584_46384# a_n1613_43370# 0.085833f
C24965 a_n3565_39590# a_n4209_37414# 0.031279f
C24966 a_3785_47178# a_3094_47570# 1.78e-21
C24967 a_n1151_42308# a_2266_47243# 2.81e-19
C24968 a_9863_47436# a_4883_46098# 9.51e-21
C24969 a_7174_31319# VDAC_P 0.009122f
C24970 a_n4209_39590# a_n3565_37414# 0.032656f
C24971 a_15673_47210# a_16588_47582# 0.125324f
C24972 a_5742_30871# C0_N_btm 0.014563f
C24973 a_13717_47436# a_19787_47423# 6.87e-20
C24974 a_15507_47210# a_10227_46804# 0.23187f
C24975 a_16327_47482# a_16023_47582# 0.159305f
C24976 a_n4064_40160# a_n4064_37440# 0.056406f
C24977 a_8325_42308# VDD 0.313956f
C24978 a_n3420_38528# a_n4064_37984# 7.35343f
C24979 a_n4064_38528# a_n3420_37984# 0.044626f
C24980 a_n2946_38778# a_n2946_37984# 0.052227f
C24981 a_13258_32519# a_22521_40599# 4.4e-19
C24982 a_20107_42308# CAL_N 0.001744f
C24983 a_n1761_44111# a_685_42968# 5.14e-21
C24984 a_n97_42460# a_n229_43646# 0.046961f
C24985 a_n2012_43396# a_n1821_43396# 4.61e-19
C24986 a_15682_43940# a_16759_43396# 0.013707f
C24987 a_11967_42832# a_5534_30871# 0.017079f
C24988 a_18114_32519# a_n1630_35242# 6.72e-20
C24989 a_n2956_37592# a_n3565_39304# 0.0261f
C24990 a_5907_45546# VDD 0.390381f
C24991 a_18451_43940# a_16137_43396# 2.49e-19
C24992 a_14976_45028# a_11341_43940# 2.74e-20
C24993 a_11453_44696# a_16137_43396# 2.08e-20
C24994 a_20841_45814# a_2437_43646# 3.5e-21
C24995 a_20273_45572# a_22223_45572# 1.24e-19
C24996 a_526_44458# a_8375_44464# 5.01e-22
C24997 a_8696_44636# a_3537_45260# 1.04e-19
C24998 a_16327_47482# a_17021_43396# 0.001903f
C24999 a_18479_45785# a_n913_45002# 1.19e-20
C25000 a_19466_46812# a_15493_43396# 2.36e-21
C25001 a_20107_45572# a_19479_31679# 5.42e-21
C25002 a_10227_46804# a_15231_43396# 9.49e-20
C25003 a_6945_45028# a_n2661_42834# 4.26e-20
C25004 a_13759_46122# a_14673_44172# 1.65e-20
C25005 C0_dummy_P_btm C0_N_btm 1.93e-19
C25006 C2_P_btm C3_N_btm 1.05e-19
C25007 C0_P_btm C1_N_btm 2.85e-19
C25008 C3_P_btm C4_N_btm 2.12e-19
C25009 a_n2661_46098# a_2864_46660# 7.93e-22
C25010 a_n2661_46634# a_7411_46660# 0.023716f
C25011 a_n2497_47436# a_2804_46116# 8.29e-22
C25012 a_n2109_47186# a_2521_46116# 1.58e-20
C25013 a_11599_46634# a_765_45546# 0.332797f
C25014 a_16763_47508# a_16721_46634# 0.005734f
C25015 a_2107_46812# a_4646_46812# 0.03082f
C25016 a_n1741_47186# a_2202_46116# 6.06e-23
C25017 a_584_46384# a_n2293_46098# 0.039917f
C25018 a_n881_46662# a_11813_46116# 8.63e-20
C25019 a_21589_35634# VDD 0.525446f
C25020 a_16588_47582# a_16388_46812# 3.64e-19
C25021 a_10227_46804# a_15227_46910# 0.00877f
C25022 a_13717_47436# a_20107_46660# 1.28e-20
C25023 a_n237_47217# a_376_46348# 2.21e-19
C25024 a_n746_45260# a_472_46348# 0.002816f
C25025 a_5807_45002# a_10249_46116# 0.041839f
C25026 a_n1925_46634# a_3633_46660# 2.55e-19
C25027 a_2443_46660# a_3524_46660# 0.102325f
C25028 a_2609_46660# a_3699_46634# 0.042415f
C25029 a_3177_46902# a_2959_46660# 0.209641f
C25030 a_n2661_42282# a_3823_42558# 1.12e-19
C25031 a_3499_42826# a_3581_42558# 1.79e-19
C25032 a_1209_43370# a_n2293_42282# 3.21e-21
C25033 a_2982_43646# a_18083_42858# 1.03e-19
C25034 a_17499_43370# a_5649_42852# 8.65e-21
C25035 a_15743_43084# a_19095_43396# 0.012939f
C25036 a_18579_44172# a_17303_42282# 8.14e-21
C25037 a_n2293_43922# a_1736_39587# 3.88e-21
C25038 a_327_44734# a_n699_43396# 1.13e-20
C25039 a_2382_45260# a_949_44458# 2.24e-19
C25040 a_n913_45002# a_10057_43914# 1.12e-19
C25041 a_n1059_45260# a_8975_43940# 5.1e-19
C25042 a_13159_45002# a_11691_44458# 1.4e-19
C25043 a_2809_45028# a_n2661_43370# 0.003105f
C25044 a_n2293_42834# a_8488_45348# 1.54e-20
C25045 a_5691_45260# a_n2661_44458# 2.93e-20
C25046 a_19692_46634# a_20749_43396# 3.6e-20
C25047 a_8696_44636# a_11541_44484# 1.04e-19
C25048 a_9290_44172# a_3626_43646# 0.014922f
C25049 w_1575_34946# a_n4064_39072# 0.016546f
C25050 a_n743_46660# a_1431_46436# 0.004109f
C25051 a_n2438_43548# a_1337_46436# 0.001827f
C25052 a_n1741_47186# a_11823_42460# 9.63e-19
C25053 a_13059_46348# a_15312_46660# 3.94e-19
C25054 a_18597_46090# a_n357_42282# 0.250702f
C25055 a_n1925_46634# a_526_44458# 1.65e-19
C25056 a_n2312_38680# a_n1925_42282# 4.88e-20
C25057 a_7577_46660# a_8016_46348# 0.003484f
C25058 a_8145_46902# a_7920_46348# 8.72e-19
C25059 a_4915_47217# a_6598_45938# 1.39e-21
C25060 a_6151_47436# a_6472_45840# 0.045851f
C25061 a_2063_45854# a_6812_45938# 0.026385f
C25062 a_19692_46634# a_18280_46660# 2.23e-20
C25063 a_22959_47212# a_20692_30879# 1.9e-19
C25064 a_19333_46634# a_19636_46660# 0.001377f
C25065 a_15368_46634# a_11415_45002# 0.001587f
C25066 a_6755_46942# a_3483_46348# 0.014154f
C25067 a_7411_46660# a_8199_44636# 1.09e-20
C25068 a_5257_43370# a_5937_45572# 0.262028f
C25069 a_743_42282# a_2351_42308# 0.00729f
C25070 a_n1076_43230# a_n4318_38216# 2.24e-19
C25071 a_12545_42858# a_12991_43230# 2.28e-19
C25072 a_n1991_42858# a_n4318_37592# 3.9e-19
C25073 a_n1853_43023# COMP_P 5.05e-20
C25074 a_n2157_42858# a_n1329_42308# 1.45e-20
C25075 a_n3674_39304# a_n3674_38680# 0.17962f
C25076 a_22959_44484# RST_Z 0.001339f
C25077 a_14579_43548# a_14113_42308# 9.55e-20
C25078 a_12281_43396# a_5742_30871# 9.39e-19
C25079 a_19237_31679# VDD 0.746512f
C25080 a_n4318_39304# a_n2946_39072# 4.19e-20
C25081 a_n357_42282# a_743_42282# 0.067793f
C25082 a_3090_45724# a_11323_42473# 4.17e-20
C25083 a_1307_43914# a_2253_44260# 7.63e-19
C25084 a_20567_45036# a_19279_43940# 1.73e-21
C25085 a_21005_45260# a_20766_44850# 1.08e-19
C25086 a_21101_45002# a_20835_44721# 4.69e-19
C25087 a_21359_45002# a_20679_44626# 9.5e-19
C25088 a_11691_44458# a_11967_42832# 0.041904f
C25089 a_11827_44484# a_20640_44752# 0.016882f
C25090 a_n2293_42834# a_1414_42308# 0.02233f
C25091 a_10775_45002# a_10949_43914# 1.24e-19
C25092 a_2711_45572# a_16977_43638# 2.53e-20
C25093 w_11334_34010# VIN_N 2.57e-20
C25094 a_4185_45028# a_14635_42282# 9.41e-20
C25095 a_10180_45724# a_9803_43646# 8.22e-23
C25096 a_10193_42453# a_9145_43396# 0.02642f
C25097 a_n23_47502# VDD 0.152616f
C25098 a_n1741_47186# DATA[3] 0.033504f
C25099 a_5883_43914# a_9159_44484# 0.049132f
C25100 a_18597_46090# CAL_N 0.001283f
C25101 a_10951_45334# a_10729_43914# 2.14e-21
C25102 a_19778_44110# a_18579_44172# 0.268475f
C25103 a_16922_45042# a_3422_30871# 5.99e-20
C25104 a_n2661_43370# a_n1899_43946# 6.55e-21
C25105 a_n356_44636# a_n310_44811# 0.006879f
C25106 a_8103_44636# a_n2661_42834# 6.31e-20
C25107 a_6298_44484# a_n2661_43922# 0.048814f
C25108 a_n913_45002# a_14021_43940# 2.81e-19
C25109 a_n815_47178# DATA[0] 0.068508f
C25110 a_n2312_38680# a_n4334_38528# 6.16e-20
C25111 a_7920_46348# a_5066_45546# 0.04093f
C25112 a_3483_46348# a_8049_45260# 0.012066f
C25113 a_n443_46116# a_5009_45028# 4.3e-20
C25114 a_4791_45118# a_5093_45028# 0.007375f
C25115 a_n1151_42308# a_8137_45348# 5.47e-21
C25116 a_n743_46660# a_17034_45572# 2.11e-19
C25117 a_768_44030# a_n2661_45010# 0.015059f
C25118 a_n1613_43370# a_n659_45366# 0.001198f
C25119 a_10227_46804# a_9482_43914# 0.032461f
C25120 a_6755_46942# a_14495_45572# 2.1e-21
C25121 a_8270_45546# a_8746_45002# 0.017581f
C25122 a_4883_46098# a_7229_43940# 6.78e-21
C25123 a_n881_46662# a_n967_45348# 6.86e-19
C25124 a_13747_46662# a_21513_45002# 0.02166f
C25125 a_13661_43548# a_2437_43646# 0.003998f
C25126 a_19321_45002# a_20719_45572# 1.72e-19
C25127 a_20916_46384# a_20731_45938# 8.76e-21
C25128 a_3090_45724# a_2211_45572# 1.16e-19
C25129 a_765_45546# a_1848_45724# 2.79e-19
C25130 a_15682_46116# a_10809_44734# 4.63e-19
C25131 a_17715_44484# a_6945_45028# 8.4e-20
C25132 a_19553_46090# a_19335_46494# 0.209641f
C25133 a_18819_46122# a_19900_46494# 0.102355f
C25134 a_18985_46122# a_20075_46420# 0.042415f
C25135 a_13467_32519# VDAC_N 3.73e-19
C25136 a_743_42282# CAL_N 4.51e-19
C25137 a_1067_42314# a_5934_30871# 1.02e-20
C25138 a_5267_42460# a_5379_42460# 0.156424f
C25139 a_1184_42692# a_6123_31319# 7.32e-21
C25140 a_3318_42354# a_3581_42558# 0.011552f
C25141 a_3823_42558# a_3497_42558# 2.37e-20
C25142 a_9145_43396# VDD 2.43736f
C25143 a_n784_42308# a_8325_42308# 2.26e-20
C25144 a_1755_42282# a_5932_42308# 0.046344f
C25145 a_n913_45002# a_2075_43172# 0.175893f
C25146 a_n357_42282# a_5755_42308# 4.82e-20
C25147 a_n1925_42282# a_7174_31319# 2.64e-20
C25148 a_15433_44458# a_11341_43940# 4.01e-21
C25149 a_n2661_42834# a_11173_44260# 0.002687f
C25150 a_644_44056# a_453_43940# 0.077973f
C25151 a_n809_44244# a_895_43940# 1.44e-19
C25152 a_11823_42460# a_14853_42852# 9.4e-19
C25153 a_n2661_44458# a_3080_42308# 1.4e-21
C25154 a_1115_44172# a_1414_42308# 0.134389f
C25155 a_10384_47026# VDD 4.6e-19
C25156 a_n2956_38680# a_n2302_40160# 6.16e-19
C25157 a_13259_45724# a_13575_42558# 0.097619f
C25158 a_n2017_45002# a_3681_42891# 1.04e-20
C25159 a_n1059_45260# a_2905_42968# 0.002465f
C25160 a_n356_45724# a_n23_45546# 0.360492f
C25161 a_2107_46812# a_10057_43914# 7.24e-20
C25162 a_n2661_45546# a_2711_45572# 0.359276f
C25163 a_13059_46348# a_16019_45002# 4.51e-21
C25164 SMPL_ON_P a_n3674_39768# 0.03705f
C25165 a_584_46384# a_2675_43914# 7.8e-20
C25166 a_n2157_46122# a_n967_45348# 1.95e-20
C25167 a_16327_47482# a_20766_44850# 0.17113f
C25168 a_n2497_47436# a_n630_44306# 3.9e-19
C25169 a_18479_47436# a_11967_42832# 0.017885f
C25170 a_12861_44030# a_20980_44850# 7.8e-21
C25171 a_n901_46420# a_n913_45002# 6.07e-19
C25172 a_n1076_46494# a_n1059_45260# 3.89e-20
C25173 a_21076_30879# a_413_45260# 0.141502f
C25174 a_12891_46348# a_9313_44734# 2.52e-21
C25175 a_6945_45028# a_15861_45028# 5.7e-21
C25176 a_4646_46812# a_n2661_44458# 0.05901f
C25177 a_8049_45260# a_14495_45572# 0.004043f
C25178 a_10586_45546# a_11823_42460# 0.005505f
C25179 a_n863_45724# a_509_45572# 3.95e-21
C25180 a_n755_45592# a_1609_45822# 0.12055f
C25181 a_997_45618# a_n443_42852# 0.093108f
C25182 a_n4064_39616# a_n2216_39866# 0.005567f
C25183 a_5934_30871# a_3726_37500# 0.002188f
C25184 a_5932_42308# VDAC_P 0.009978f
C25185 a_2905_45572# a_3785_47178# 0.013619f
C25186 a_2124_47436# a_n443_46116# 6.88e-22
C25187 a_3160_47472# a_3381_47502# 0.099936f
C25188 a_n237_47217# a_6851_47204# 8.46e-19
C25189 a_n971_45724# a_7903_47542# 7.01e-19
C25190 a_n1741_47186# a_9313_45822# 0.102019f
C25191 a_n2288_47178# a_n1435_47204# 2.38e-19
C25192 a_n4064_40160# a_n3420_39072# 0.052668f
C25193 a_n3565_39590# a_n3607_39616# 0.001003f
C25194 a_14097_32519# C5_N_btm 0.001712f
C25195 a_n1630_35242# EN_VIN_BSTR_N 0.009773f
C25196 a_n4315_30879# a_n4064_39072# 0.036792f
C25197 a_n4209_39590# a_n4209_39304# 0.045123f
C25198 a_14539_43914# a_18083_42858# 0.00221f
C25199 a_n699_43396# a_133_42852# 1.03e-19
C25200 a_3422_30871# a_15743_43084# 0.022574f
C25201 a_11967_42832# a_4190_30871# 0.002622f
C25202 a_n356_44636# a_12545_42858# 4.75e-20
C25203 a_1307_43914# a_2713_42308# 4.75e-19
C25204 a_n1059_45260# a_15803_42450# 0.008866f
C25205 a_n2017_45002# a_15959_42545# 0.004519f
C25206 a_n913_45002# a_15764_42576# 5.85e-19
C25207 a_5891_43370# a_8037_42858# 0.12253f
C25208 a_n2661_42282# a_6765_43638# 2.44e-19
C25209 a_10807_43548# a_3626_43646# 0.001709f
C25210 a_14180_46482# VDD 0.077608f
C25211 a_n2293_42834# a_n3674_38680# 0.010983f
C25212 a_742_44458# a_1793_42852# 0.010622f
C25213 a_n357_42282# a_626_44172# 0.551369f
C25214 a_n755_45592# a_501_45348# 5.21e-19
C25215 a_n863_45724# a_2809_45348# 1.93e-19
C25216 a_n443_42852# a_13159_45002# 1.23e-20
C25217 a_12549_44172# a_14401_32519# 0.004427f
C25218 a_2711_45572# a_5205_44484# 8.29e-19
C25219 a_8049_45260# a_17719_45144# 3.83e-20
C25220 a_15599_45572# a_18341_45572# 1.38e-21
C25221 a_10193_42453# a_n1059_45260# 0.440111f
C25222 a_15765_45572# a_18175_45572# 6.29e-20
C25223 a_n1613_43370# a_n1177_43370# 0.325171f
C25224 a_4915_47217# a_14358_43442# 3.86e-20
C25225 a_2324_44458# a_9838_44484# 4.19e-20
C25226 a_12594_46348# a_13076_44458# 4.02e-22
C25227 a_n2661_45546# a_4640_45348# 0.003021f
C25228 a_5907_45546# a_5691_45260# 0.001013f
C25229 a_4185_45028# a_4181_44734# 5.69e-19
C25230 a_3483_46348# a_5289_44734# 5.06e-20
C25231 a_13507_46334# a_2982_43646# 0.063751f
C25232 a_8696_44636# a_16842_45938# 1.95e-20
C25233 a_16333_45814# a_16147_45260# 1.26e-19
C25234 a_12741_44636# a_14112_44734# 7.78e-19
C25235 a_3775_45552# a_3429_45260# 0.001061f
C25236 a_2957_45546# a_1307_43914# 1.73e-20
C25237 a_9804_47204# a_2107_46812# 0.033493f
C25238 a_13487_47204# a_6755_46942# 1.18e-19
C25239 a_n4209_37414# C4_P_btm 9.91e-21
C25240 a_n3565_37414# C6_P_btm 1.26e-20
C25241 a_11599_46634# a_10623_46897# 3.51e-20
C25242 a_3726_37500# a_11530_34132# 3.03e-19
C25243 a_20843_47204# a_20916_46384# 8.16e-20
C25244 a_5700_37509# a_n923_35174# 3.61e-19
C25245 a_n237_47217# a_10425_46660# 2.5e-20
C25246 a_2747_46873# a_3067_47026# 4.09e-19
C25247 a_7754_39632# VDD 0.205733f
C25248 a_n3420_37984# VREF_GND 0.047887f
C25249 a_4883_46098# a_5907_46634# 5.32e-21
C25250 a_22469_40625# a_22705_38406# 1.29e-19
C25251 a_22521_40599# a_22609_37990# 0.021352f
C25252 a_22521_40055# CAL_P 0.001469f
C25253 a_22521_39511# a_22469_39537# 1.02751f
C25254 a_22545_38993# a_22821_38993# 0.235701f
C25255 a_n1613_43370# a_479_46660# 1.79e-19
C25256 a_6151_47436# a_8846_46660# 0.002879f
C25257 a_2905_45572# a_3090_45724# 0.006554f
C25258 a_4915_47217# a_11735_46660# 3.49e-19
C25259 a_n1151_42308# a_14084_46812# 0.063788f
C25260 a_2982_43646# a_21855_43396# 2.81e-19
C25261 a_n4318_40392# a_n4064_39072# 2.29e-21
C25262 a_n1761_44111# a_n1329_42308# 7.38e-20
C25263 a_n1899_43946# COMP_P 4.56e-21
C25264 a_19963_31679# EN_OFFSET_CAL 4.91e-20
C25265 a_n1059_45260# VDD 4.75361f
C25266 a_n229_43646# a_n901_43156# 3.1e-19
C25267 a_n2017_45002# RST_Z 1.48e-20
C25268 a_14205_43396# a_14621_43646# 2.64e-19
C25269 a_14021_43940# a_20922_43172# 6.69e-20
C25270 a_19479_31679# VIN_N 0.029355f
C25271 a_3422_30871# a_1606_42308# 0.022481f
C25272 a_n2293_43922# a_13070_42354# 0.002481f
C25273 a_13667_43396# a_13749_43396# 0.005781f
C25274 a_3483_46348# a_15037_43940# 0.007725f
C25275 a_5691_45260# a_6125_45348# 0.003935f
C25276 a_3537_45260# a_5009_45028# 0.001769f
C25277 a_20107_45572# a_20193_45348# 8.83e-19
C25278 a_15227_44166# a_14579_43548# 7.96e-19
C25279 a_3090_45724# a_10765_43646# 6.96e-19
C25280 a_14537_43396# a_14797_45144# 0.082443f
C25281 a_8696_44636# a_8701_44490# 0.095858f
C25282 en_comp a_n2661_43370# 0.164814f
C25283 a_21188_45572# a_11827_44484# 1.57e-20
C25284 a_10227_46804# a_11301_43218# 1.79e-19
C25285 a_n2293_46634# a_8952_43230# 1.4e-20
C25286 a_5807_45002# a_5534_30871# 3.81e-20
C25287 a_n443_42852# a_11967_42832# 0.00555f
C25288 a_9482_43914# a_1307_43914# 0.010221f
C25289 a_5937_45572# a_5745_43940# 4.36e-20
C25290 a_n2497_47436# a_n1099_45572# 0.004833f
C25291 a_768_44030# a_10903_43370# 0.082359f
C25292 SMPL_ON_P a_n2293_45546# 8.05e-20
C25293 a_n743_46660# a_2202_46116# 0.012092f
C25294 a_n1925_46634# a_2521_46116# 8.92e-20
C25295 a_n2438_43548# a_1823_45246# 0.002972f
C25296 a_5807_45002# a_5937_45572# 0.038681f
C25297 a_9313_45822# a_10586_45546# 6.08e-20
C25298 a_6755_46942# a_14513_46634# 0.036712f
C25299 a_n2661_46634# a_4185_45028# 1.65e-19
C25300 a_n2293_46634# a_3147_46376# 1.96e-19
C25301 a_13487_47204# a_8049_45260# 1.12e-20
C25302 a_n881_46662# a_15682_46116# 7.66e-19
C25303 a_12891_46348# a_12594_46348# 0.088156f
C25304 a_601_46902# a_805_46414# 7.84e-19
C25305 a_383_46660# a_472_46348# 8.96e-19
C25306 a_171_46873# a_1176_45822# 5.65e-20
C25307 a_7411_46660# a_765_45546# 0.003093f
C25308 a_n2312_39304# a_n2956_39304# 6.38528f
C25309 a_n2312_40392# a_n2956_38680# 0.052782f
C25310 a_16977_43638# a_16877_42852# 6.98e-20
C25311 a_15743_43084# a_18504_43218# 2.23e-19
C25312 a_n97_42460# a_13070_42354# 0.02477f
C25313 a_2982_43646# a_7227_42308# 6.66e-20
C25314 a_12379_42858# a_12545_42858# 0.810394f
C25315 a_13661_43548# a_19511_42282# 4.91e-21
C25316 a_4223_44672# a_n699_43396# 0.217586f
C25317 a_11691_44458# a_18989_43940# 0.066207f
C25318 a_n2840_45002# a_n4318_39768# 0.002422f
C25319 a_9290_44172# a_8037_42858# 2.48e-20
C25320 a_n443_42852# a_648_43396# 0.002995f
C25321 a_n2661_44458# a_10057_43914# 0.007497f
C25322 a_n2312_39304# a_n3565_39304# 0.104981f
C25323 a_413_45260# a_1414_42308# 0.12534f
C25324 a_n913_45002# a_5013_44260# 7.77e-21
C25325 a_n1059_45260# a_5495_43940# 1.76e-21
C25326 a_16147_45260# a_15493_43396# 9.87e-21
C25327 a_8953_45546# a_10083_42826# 8.07e-20
C25328 a_8199_44636# a_10835_43094# 4.6e-21
C25329 a_3483_46348# a_15279_43071# 5.23e-21
C25330 a_4185_45028# a_14543_43071# 9.15e-22
C25331 w_11334_34010# CAL_N 1.49e-19
C25332 w_1575_34946# VDD 1.58877f
C25333 a_5257_43370# a_n443_42852# 0.016836f
C25334 a_n2293_46634# a_13249_42308# 0.027384f
C25335 a_11415_45002# a_20708_46348# 5.4e-21
C25336 a_20202_43084# a_21137_46414# 0.006423f
C25337 a_3483_46348# a_8953_45546# 0.133493f
C25338 a_4185_45028# a_8199_44636# 1.24e-19
C25339 a_20719_46660# a_10809_44734# 6.1e-19
C25340 a_14955_47212# a_2437_43646# 0.009063f
C25341 a_6755_46942# a_n357_42282# 3.13e-20
C25342 a_n237_47217# a_3232_43370# 7.83e-20
C25343 a_3381_47502# a_413_45260# 0.001239f
C25344 a_n1151_42308# a_327_44734# 8.48e-19
C25345 a_n881_46662# a_16680_45572# 0.051767f
C25346 a_n1613_43370# a_8696_44636# 5.83e-19
C25347 a_18479_47436# a_20273_45572# 0.028755f
C25348 a_16327_47482# a_19365_45572# 4.87e-19
C25349 a_4646_46812# a_5907_45546# 3.34e-21
C25350 a_n743_46660# a_11823_42460# 5.08e-19
C25351 a_12741_44636# a_19335_46494# 1.88e-20
C25352 a_15368_46634# a_13259_45724# 0.0178f
C25353 a_2063_45854# a_3065_45002# 4.37e-20
C25354 a_584_46384# a_3429_45260# 4.23e-21
C25355 a_10227_46804# a_20623_45572# 4e-20
C25356 a_11453_44696# a_18479_45785# 0.003588f
C25357 a_12861_44030# a_3357_43084# 3.68e-19
C25358 a_n2840_43370# VDD 0.246858f
C25359 a_16414_43172# a_16522_42674# 6.05e-20
C25360 a_5342_30871# a_15521_42308# 2.73e-19
C25361 a_5111_44636# a_10695_43548# 6.49e-20
C25362 a_4185_45028# a_19511_42282# 9.41e-20
C25363 a_n743_46660# DATA[3] 1.69e-21
C25364 a_n2293_42834# a_n1190_43762# 8.33e-20
C25365 a_1307_43914# a_6031_43396# 0.002834f
C25366 a_13249_42308# a_5342_30871# 7.46e-20
C25367 a_10193_42453# a_19987_42826# 0.164153f
C25368 a_948_46660# VDD 0.278482f
C25369 a_9482_43914# a_9396_43370# 0.011522f
C25370 a_15004_44636# a_14955_43940# 2.26e-20
C25371 a_n2661_43922# a_2479_44172# 0.002669f
C25372 a_n2661_42834# a_895_43940# 0.095907f
C25373 a_171_46873# DATA[0] 9.78e-20
C25374 a_n2017_45002# a_16243_43396# 9.54e-20
C25375 a_n1059_45260# a_16137_43396# 0.438785f
C25376 a_n1925_42282# a_5932_42308# 0.004062f
C25377 a_526_44458# a_6481_42558# 0.001415f
C25378 a_20159_44458# a_18579_44172# 4.88e-19
C25379 a_17517_44484# a_20512_43084# 0.027951f
C25380 a_20835_44721# a_20766_44850# 0.209641f
C25381 a_20679_44626# a_19279_43940# 0.279785f
C25382 a_375_42282# a_648_43396# 9.82e-19
C25383 a_n2661_43370# a_n1699_43638# 7.67e-21
C25384 a_10903_43370# a_11652_45724# 0.010404f
C25385 a_12594_46348# a_11322_45546# 1.17e-19
C25386 a_n743_46660# a_16321_45348# 7.66e-19
C25387 a_19321_45002# a_11827_44484# 0.037739f
C25388 a_7832_46660# a_7705_45326# 7.57e-21
C25389 a_12549_44172# a_20205_45028# 7.43e-20
C25390 a_18280_46660# a_18175_45572# 1.14e-20
C25391 a_19692_46634# a_n913_45002# 2.2e-20
C25392 a_12465_44636# a_13076_44458# 0.01224f
C25393 a_11189_46129# a_11823_42460# 1.55e-19
C25394 a_18147_46436# a_18051_46116# 1.26e-19
C25395 a_5807_45002# a_11691_44458# 0.117249f
C25396 a_13747_46662# a_22959_45036# 4.74e-20
C25397 a_13661_43548# a_19113_45348# 0.003675f
C25398 a_3483_46348# a_8791_45572# 5.57e-19
C25399 a_8270_45546# a_3232_43370# 0.020859f
C25400 a_14180_46812# a_3357_43084# 1.32e-20
C25401 a_n1613_43370# a_n1177_44458# 0.332209f
C25402 a_15009_46634# a_413_45260# 1.08e-20
C25403 a_6123_31319# comp_n 1.63e-19
C25404 a_5934_30871# a_1239_39043# 6.07e-20
C25405 a_19987_42826# VDD 0.588466f
C25406 a_18057_42282# a_18214_42558# 0.18824f
C25407 a_5342_30871# VIN_P 0.00693f
C25408 a_19164_43230# RST_Z 1.35e-21
C25409 a_n2293_45010# a_564_42282# 6.44e-21
C25410 a_2127_44172# a_n97_42460# 1.47e-19
C25411 a_18989_43940# a_4190_30871# 1.16e-19
C25412 a_15493_43940# a_22959_43948# 0.182001f
C25413 a_15433_44458# a_10341_43396# 1.5e-21
C25414 a_n1059_45260# a_n784_42308# 0.008929f
C25415 a_n913_45002# a_196_42282# 1.19e-19
C25416 a_n2017_45002# a_n327_42558# 0.005655f
C25417 a_7584_44260# a_7499_43940# 1.48e-19
C25418 a_9313_44734# a_16409_43396# 6.68e-20
C25419 en_comp COMP_P 1.92051f
C25420 a_n967_45348# a_n4318_37592# 8.19e-19
C25421 a_13925_46122# VDD 0.251868f
C25422 a_n2293_42834# a_873_42968# 1.97e-20
C25423 a_13759_46122# RST_Z 8.63e-20
C25424 a_18451_43940# a_14021_43940# 1.25e-20
C25425 a_2324_44458# a_n2661_43370# 0.082794f
C25426 a_n901_46420# a_n2661_44458# 9.89e-21
C25427 a_n2293_46098# a_n1177_44458# 1.38e-20
C25428 a_2711_45572# a_19431_45546# 2.71e-21
C25429 a_n2956_38216# a_n2840_45002# 0.01122f
C25430 a_11453_44696# a_14021_43940# 8.33e-20
C25431 a_584_46384# a_1209_43370# 0.02923f
C25432 a_n971_45724# a_n1557_42282# 0.06901f
C25433 a_n1925_42282# a_1423_45028# 0.021671f
C25434 a_11823_42460# a_11136_45572# 5.02e-20
C25435 a_11962_45724# a_11778_45572# 5.39e-20
C25436 a_n1991_46122# a_n2267_44484# 7.99e-21
C25437 a_10193_42453# a_15599_45572# 5.53e-20
C25438 a_n2438_43548# a_n3674_39768# 0.007137f
C25439 a_n2661_45546# a_n2472_45002# 0.004199f
C25440 a_8049_45260# a_11963_45334# 1.58e-20
C25441 a_12549_44172# a_15682_43940# 0.058263f
C25442 a_7754_40130# a_3726_37500# 0.021358f
C25443 a_2747_46873# a_3094_47243# 9.52e-20
C25444 a_4883_46098# a_768_44030# 0.045313f
C25445 a_18479_47436# a_5807_45002# 2.73e-19
C25446 a_16327_47482# a_16750_47204# 3.03e-19
C25447 a_6545_47178# a_2107_46812# 0.028617f
C25448 a_13258_32519# VIN_N 0.143165f
C25449 a_n3420_39072# C10_P_btm 3.37e-20
C25450 a_n4315_30879# VDD 4.0486f
C25451 a_n4209_39304# C6_P_btm 0.001067f
C25452 a_10227_46804# a_13747_46662# 0.16398f
C25453 a_18143_47464# a_13661_43548# 0.011802f
C25454 a_n237_47217# a_4651_46660# 7.27e-20
C25455 a_3160_47472# a_2959_46660# 0.00952f
C25456 a_3381_47502# a_2609_46660# 0.00165f
C25457 a_n1151_42308# a_3177_46902# 0.006126f
C25458 a_584_46384# a_1057_46660# 6.68e-21
C25459 a_2905_45572# a_3699_46634# 0.00292f
C25460 a_12861_44030# a_n2293_46634# 6.64e-19
C25461 a_9313_45822# a_n743_46660# 0.029372f
C25462 a_n2109_47186# a_5275_47026# 0.001536f
C25463 a_n1741_47186# a_6540_46812# 7e-21
C25464 a_n971_45724# a_4817_46660# 1.65e-19
C25465 a_n4209_38502# a_n1838_35608# 1.6e-19
C25466 a_12465_44636# a_12891_46348# 0.033919f
C25467 a_n3565_39304# C8_P_btm 1.15e-19
C25468 a_11967_42832# a_14635_42282# 0.018349f
C25469 a_n2293_43922# a_n4318_38216# 5.44e-19
C25470 a_18494_42460# a_18214_42558# 0.012583f
C25471 a_18184_42460# a_18220_42308# 5.62e-19
C25472 a_n2956_37592# a_n3690_37440# 0.015408f
C25473 a_15599_45572# VDD 0.390565f
C25474 a_n356_44636# a_5379_42460# 0.038779f
C25475 a_2479_44172# a_3445_43172# 1.16e-19
C25476 a_n2810_45028# a_n3420_37440# 0.009781f
C25477 a_14021_43940# a_17364_32525# 0.007637f
C25478 a_5883_43914# a_9293_42558# 2.71e-21
C25479 a_19808_44306# a_15743_43084# 5.11e-21
C25480 a_19319_43548# a_18783_43370# 9.48e-20
C25481 a_18533_43940# a_18525_43370# 7.52e-19
C25482 a_6765_43638# a_7112_43396# 0.051162f
C25483 a_15143_45578# a_11691_44458# 3.46e-19
C25484 a_10227_46804# a_10796_42968# 0.024053f
C25485 a_n971_45724# a_8483_43230# 2.48e-19
C25486 a_2711_45572# a_13076_44458# 6.99e-21
C25487 a_10180_45724# a_n2661_44458# 2.83e-19
C25488 a_2324_44458# a_2998_44172# 2.03e-19
C25489 a_413_45260# a_1667_45002# 0.00537f
C25490 a_n2017_45002# a_3232_43370# 1.68e-19
C25491 a_n1613_43370# a_n1991_42858# 0.029351f
C25492 a_n23_45546# a_n356_44636# 1.17e-20
C25493 a_13661_43548# a_21259_43561# 2.35e-20
C25494 a_5807_45002# a_4190_30871# 8.86e-22
C25495 w_1575_34946# a_n784_42308# 0.001423f
C25496 a_8667_46634# a_8492_46660# 0.233657f
C25497 a_n2497_47436# a_n1925_42282# 0.004955f
C25498 a_n971_45724# a_n722_46482# 1.89e-19
C25499 a_4915_47217# a_2324_44458# 0.022906f
C25500 a_5807_45002# a_17829_46910# 3.44e-20
C25501 a_2443_46660# a_3090_45724# 2.52e-20
C25502 a_9313_45822# a_11189_46129# 1.48e-22
C25503 a_n1435_47204# a_9823_46155# 4.27e-21
C25504 a_13747_46662# a_17339_46660# 0.015626f
C25505 a_13661_43548# a_765_45546# 1.39e-19
C25506 a_n2312_39304# a_n1991_46122# 0.00213f
C25507 a_16137_43396# a_19987_42826# 2.41e-19
C25508 a_17499_43370# a_17333_42852# 7.75e-20
C25509 a_15743_43084# a_16414_43172# 1.55e-19
C25510 a_743_42282# a_8952_43230# 3.27e-20
C25511 a_n3674_39304# a_n4318_38680# 2.92578f
C25512 a_n2129_43609# a_n961_42308# 1.71e-20
C25513 a_15493_43396# a_15051_42282# 3.6e-21
C25514 a_5649_42852# a_5755_42852# 0.089078f
C25515 a_n1853_43023# a_133_43172# 6.79e-19
C25516 a_n1991_42858# a_n1533_42852# 0.034619f
C25517 a_n4318_40392# VDD 0.573389f
C25518 a_n2267_43396# a_n1329_42308# 8.36e-21
C25519 a_n1699_43638# COMP_P 9.19e-20
C25520 a_4361_42308# a_7765_42852# 3.76e-20
C25521 a_n2293_42834# a_n699_43396# 0.00729f
C25522 a_18184_42460# a_11827_44484# 0.027981f
C25523 a_19778_44110# a_22223_45036# 6.5e-20
C25524 a_18494_42460# a_21359_45002# 4.97e-21
C25525 a_2680_45002# a_n2661_43922# 6.61e-20
C25526 a_3065_45002# a_n2661_42834# 0.022516f
C25527 a_2382_45260# a_n2293_43922# 5.18e-20
C25528 a_10193_42453# a_18326_43940# 0.130866f
C25529 a_19692_46634# a_20922_43172# 5.29e-20
C25530 a_n1925_42282# a_4181_43396# 1.15e-19
C25531 a_12861_44030# a_20107_42308# 1.45e-21
C25532 a_n2661_43370# a_n1699_44726# 0.001811f
C25533 a_5147_45002# a_5608_44484# 0.003234f
C25534 a_2437_43646# a_11967_42832# 4.65e-20
C25535 a_3090_45724# a_4156_43218# 2.05e-21
C25536 a_8191_45002# a_5891_43370# 6.65e-19
C25537 a_18587_45118# a_19113_45348# 2.02e-19
C25538 a_20567_45036# a_21101_45002# 3.03e-19
C25539 a_18315_45260# a_11691_44458# 8.2e-21
C25540 a_12427_45724# a_12429_44172# 4.6e-20
C25541 a_11823_42460# a_11750_44172# 6.71e-20
C25542 a_2324_44458# a_15681_43442# 0.006403f
C25543 a_4185_45028# a_21259_43561# 4.43e-21
C25544 a_10227_46804# a_4958_30871# 0.036177f
C25545 a_16327_47482# a_18907_42674# 0.001573f
C25546 a_12465_44636# a_11322_45546# 5.04e-19
C25547 a_4883_46098# a_11652_45724# 1.56e-19
C25548 a_n1021_46688# a_n863_45724# 5e-21
C25549 a_n2293_46634# a_310_45028# 0.020873f
C25550 a_5807_45002# a_n443_42852# 1.54e-19
C25551 a_n881_46662# a_6598_45938# 0.031336f
C25552 a_n1613_43370# a_7227_45028# 8.73e-21
C25553 a_11453_44696# a_10180_45724# 2.98e-19
C25554 a_n2438_43548# a_n2293_45546# 0.051617f
C25555 a_33_46660# a_n2661_45546# 4.08e-20
C25556 a_7715_46873# a_8034_45724# 9.01e-19
C25557 a_n743_46660# a_n1079_45724# 1.23e-19
C25558 a_12891_46348# a_2711_45572# 0.027614f
C25559 a_4791_45118# a_8696_44636# 0.097007f
C25560 a_12741_44636# a_22959_46660# 0.17409f
C25561 a_20820_30879# a_21076_30879# 8.6867f
C25562 a_765_45546# a_4185_45028# 7.51e-20
C25563 a_11735_46660# a_10809_44734# 0.030929f
C25564 a_11901_46660# a_6945_45028# 1.36e-19
C25565 a_12359_47026# a_12594_46348# 1.26e-19
C25566 a_3090_45724# a_18819_46122# 2.43e-19
C25567 a_n2661_46634# a_997_45618# 3.38e-22
C25568 a_10405_44172# CLK 6.38e-19
C25569 a_18326_43940# VDD 0.129408f
C25570 a_15743_43084# a_7174_31319# 3.05e-19
C25571 a_16823_43084# a_18057_42282# 2.44e-21
C25572 a_4361_42308# a_13657_42308# 5.57e-19
C25573 a_n2293_42282# a_n3674_38216# 0.111055f
C25574 a_7227_42852# a_6123_31319# 0.001591f
C25575 a_18989_43940# a_18753_44484# 4.75e-19
C25576 a_2779_44458# a_1414_42308# 5.89e-19
C25577 a_22612_30879# a_22459_39145# 7.31e-20
C25578 a_11823_42460# a_4361_42308# 0.056415f
C25579 a_13249_42308# a_743_42282# 0.010211f
C25580 a_n467_45028# a_n229_43646# 6.99e-21
C25581 a_12465_44636# SINGLE_ENDED 0.067716f
C25582 a_n699_43396# a_1115_44172# 6.01e-20
C25583 a_n913_45002# a_4699_43561# 8.4e-21
C25584 a_n1059_45260# a_3080_42308# 0.025424f
C25585 a_n2017_45002# a_4905_42826# 0.042734f
C25586 a_n2293_45010# a_n1557_42282# 1.08e-20
C25587 a_n357_42282# a_15279_43071# 0.007143f
C25588 a_1307_43914# a_6671_43940# 0.007083f
C25589 a_2382_45260# a_n97_42460# 0.02063f
C25590 a_949_44458# a_453_43940# 0.006129f
C25591 a_742_44458# a_2127_44172# 0.002775f
C25592 a_n2661_44458# a_5013_44260# 2.48e-20
C25593 a_9482_43914# a_10867_43940# 2.96e-19
C25594 a_22731_47423# RST_Z 4.82e-19
C25595 a_4185_45028# a_4921_42308# 0.059648f
C25596 a_n443_42852# a_10518_42984# 1.45e-19
C25597 SMPL_ON_N VDD 0.503419f
C25598 a_n2661_46634# a_13159_45002# 0.062031f
C25599 a_n743_46660# a_7705_45326# 4.03e-20
C25600 a_1176_45822# a_1260_45572# 0.00411f
C25601 a_1138_42852# a_1176_45572# 7.3e-19
C25602 a_n1151_42308# a_4223_44672# 1.31e-20
C25603 a_5894_47026# a_3357_43084# 1.88e-19
C25604 a_17957_46116# a_18051_46116# 0.062574f
C25605 a_18985_46122# a_19431_46494# 2.28e-19
C25606 a_19335_46494# a_16375_45002# 4.62e-20
C25607 a_8953_45546# a_n357_42282# 0.054106f
C25608 a_2063_45854# a_6298_44484# 5.31e-21
C25609 a_2959_46660# a_413_45260# 0.011261f
C25610 a_15227_44166# a_16115_45572# 2.6e-21
C25611 a_4646_46812# a_n1059_45260# 0.001886f
C25612 a_5257_43370# a_2437_43646# 7.48e-20
C25613 a_3090_45724# a_16223_45938# 0.002393f
C25614 a_2443_46660# a_2274_45254# 9.71e-22
C25615 a_13661_43548# a_16751_45260# 1.24e-19
C25616 a_13747_46662# a_1307_43914# 5.92e-20
C25617 a_16327_47482# a_21005_45260# 0.004367f
C25618 a_5742_30871# a_11551_42558# 0.007648f
C25619 a_5934_30871# a_9885_42308# 0.001708f
C25620 a_n4318_38216# a_n3420_39616# 0.023792f
C25621 a_5342_30871# a_11206_38545# 2.16e-20
C25622 a_22959_43396# VDD 0.303237f
C25623 a_n3674_38680# a_n4064_39616# 0.019915f
C25624 a_14209_32519# RST_Z 0.049869f
C25625 a_1606_42308# a_7174_31319# 2.41314f
C25626 a_n356_44636# a_7287_43370# 7.66e-21
C25627 a_3499_42826# a_n2661_42282# 1.48e-20
C25628 a_11691_44458# a_16867_43762# 7.88e-20
C25629 a_n2293_42834# a_n4318_38680# 0.007189f
C25630 a_1307_43914# a_10796_42968# 1.45e-20
C25631 a_2382_45260# a_3935_43218# 0.005937f
C25632 a_10057_43914# a_9145_43396# 0.121499f
C25633 a_15004_44636# a_8685_43396# 8.84e-21
C25634 a_n357_42282# a_13258_32519# 0.022774f
C25635 a_n2661_42834# a_458_43396# 0.001339f
C25636 a_7499_43078# a_9223_42460# 0.013802f
C25637 a_3065_45002# a_n2293_42282# 0.007636f
C25638 a_9482_43914# a_13635_43156# 3.22e-21
C25639 a_1423_45028# a_8387_43230# 4.08e-21
C25640 a_2698_46116# a_1423_45028# 6.57e-22
C25641 a_1823_45246# a_2903_45348# 1.47e-19
C25642 a_10355_46116# a_8953_45002# 4.75e-20
C25643 a_n2293_46098# a_5009_45028# 0.009429f
C25644 a_n2956_39304# a_n2810_45028# 0.042912f
C25645 a_3090_45724# a_949_44458# 3.71e-22
C25646 a_12549_44172# a_20512_43084# 0.002813f
C25647 a_13059_46348# a_11827_44484# 0.495367f
C25648 a_n1613_43370# a_n1331_43914# 0.16678f
C25649 a_6511_45714# a_7499_43078# 1.26e-20
C25650 a_7227_45028# a_7230_45938# 0.170618f
C25651 a_6598_45938# a_8162_45546# 9.36e-20
C25652 a_19335_46494# a_413_45260# 1.78e-21
C25653 a_2324_44458# a_4574_45260# 9.08e-20
C25654 a_8270_45546# a_8975_43940# 0.207334f
C25655 a_13747_46662# a_18579_44172# 1.11e-20
C25656 a_13661_43548# a_18681_44484# 6.47e-19
C25657 a_17339_46660# a_18911_45144# 1.25e-21
C25658 a_13351_46090# a_6171_45002# 1.13e-20
C25659 a_8016_46348# a_9482_43914# 0.293982f
C25660 a_167_45260# a_2304_45348# 6.8e-19
C25661 a_2711_45572# a_11322_45546# 0.056109f
C25662 a_2063_45854# a_10555_44260# 0.001312f
C25663 w_1575_34946# a_3080_42308# 0.001676f
C25664 a_12861_44030# a_18597_46090# 0.045766f
C25665 a_13717_47436# a_19386_47436# 8e-20
C25666 a_1431_47204# a_n881_46662# 3.11e-20
C25667 a_2124_47436# a_n1613_43370# 2.83e-20
C25668 a_n1151_42308# a_3315_47570# 0.003697f
C25669 a_4007_47204# a_2747_46873# 3.71e-20
C25670 a_n4315_30879# a_n2302_37690# 1.98e-19
C25671 a_15673_47210# a_16763_47508# 0.042509f
C25672 a_9067_47204# a_4883_46098# 1.74e-20
C25673 a_4958_30871# CAL_P 0.007236f
C25674 a_1736_39587# a_3754_38802# 1.04e-19
C25675 a_n4209_39590# a_n4334_37440# 2.73e-19
C25676 a_5742_30871# C0_dummy_N_btm 2.87e-19
C25677 a_n3565_38502# a_n2302_37984# 2.07e-19
C25678 a_2112_39137# a_2113_38308# 0.479143f
C25679 a_8337_42558# VDD 0.006426f
C25680 a_n4064_40160# a_n2946_37690# 1.87e-20
C25681 a_11599_46634# a_10227_46804# 0.60865f
C25682 a_16241_47178# a_16023_47582# 0.209641f
C25683 a_15507_47210# a_17591_47464# 1.96e-21
C25684 a_13258_32519# CAL_N 0.020535f
C25685 a_14021_43940# a_9145_43396# 0.032057f
C25686 a_5891_43370# a_7309_42852# 0.071511f
C25687 a_14539_43914# a_14853_42852# 3.54e-21
C25688 a_1307_43914# a_4958_30871# 9.67e-22
C25689 en_comp a_n4209_39304# 3.42e-19
C25690 a_n1352_43396# a_458_43396# 1.68e-20
C25691 a_19319_43548# a_3626_43646# 4.18e-20
C25692 a_n447_43370# a_n229_43646# 0.08213f
C25693 a_15682_43940# a_16977_43638# 0.003291f
C25694 a_11967_42832# a_14543_43071# 0.022161f
C25695 a_5263_45724# VDD 0.202719f
C25696 a_n2810_45028# a_n3565_39304# 0.021534f
C25697 a_17517_44484# a_18249_42858# 8.87e-22
C25698 a_18326_43940# a_16137_43396# 3.25e-22
C25699 a_3090_45724# a_11341_43940# 0.041393f
C25700 a_n357_42282# a_20193_45348# 0.006712f
C25701 a_20107_45572# a_22223_45572# 7.3e-21
C25702 a_21188_45572# a_21350_45938# 0.006453f
C25703 a_20623_45572# a_20885_45572# 0.001705f
C25704 a_20273_45572# a_2437_43646# 8.82e-20
C25705 a_16327_47482# a_16855_43396# 1.79e-19
C25706 a_10227_46804# a_15125_43396# 1.54e-19
C25707 a_10809_44734# a_10617_44484# 0.014699f
C25708 a_526_44458# a_7640_43914# 1.26e-20
C25709 a_6667_45809# a_n2661_43370# 3.11e-20
C25710 a_768_44030# a_8685_43396# 1.24e-19
C25711 a_12861_44030# a_743_42282# 6.92e-20
C25712 C0_dummy_P_btm C0_dummy_N_btm 0.033511f
C25713 C7_P_btm C7_N_btm 0.028901f
C25714 C6_P_btm C6_N_btm 0.019861f
C25715 C5_P_btm C5_N_btm 0.03705f
C25716 C4_P_btm C4_N_btm 0.02642f
C25717 C3_P_btm C3_N_btm 2.90968f
C25718 C2_P_btm C2_N_btm 0.026698f
C25719 C1_P_btm C1_N_btm 0.06624f
C25720 C0_P_btm C0_N_btm 0.044538f
C25721 a_1799_45572# a_2864_46660# 3.88e-20
C25722 a_n2661_46634# a_5257_43370# 0.005264f
C25723 a_n2497_47436# a_2698_46116# 1.45e-22
C25724 a_n2109_47186# a_167_45260# 4.41e-20
C25725 a_11453_44696# a_19692_46634# 0.05834f
C25726 a_11599_46634# a_17339_46660# 0.131185f
C25727 a_14955_47212# a_765_45546# 0.004861f
C25728 a_16763_47508# a_16388_46812# 5.51e-19
C25729 a_2107_46812# a_3877_44458# 0.070722f
C25730 a_n743_46660# a_6540_46812# 7.69e-21
C25731 a_n1741_47186# a_1823_45246# 8.12e-20
C25732 a_n881_46662# a_11735_46660# 1.34e-19
C25733 a_19864_35138# VDD 0.332629f
C25734 a_12861_44030# a_19123_46287# 0.002675f
C25735 a_n746_45260# a_376_46348# 0.010981f
C25736 a_n971_45724# a_472_46348# 5.63e-20
C25737 a_5807_45002# a_10554_47026# 0.003779f
C25738 a_2609_46660# a_2959_46660# 0.216095f
C25739 a_2443_46660# a_3699_46634# 0.043475f
C25740 a_16327_47482# a_16434_46987# 0.00105f
C25741 a_10227_46804# a_13693_46688# 0.002261f
C25742 a_n2661_42282# a_3318_42354# 1.07e-19
C25743 a_3499_42826# a_3497_42558# 1.79e-19
C25744 a_20193_45348# CAL_N 8.22e-19
C25745 a_458_43396# a_n2293_42282# 1.03e-20
C25746 a_3626_43646# a_16795_42852# 2.28e-21
C25747 a_2982_43646# a_17701_42308# 1.83e-19
C25748 a_7845_44172# a_7963_42308# 7.62e-22
C25749 a_19700_43370# a_743_42282# 0.001969f
C25750 a_15743_43084# a_21487_43396# 1.58e-19
C25751 a_18783_43370# a_19095_43396# 0.038241f
C25752 a_n2293_43922# a_1239_39587# 1.55e-20
C25753 a_2274_45254# a_949_44458# 3.92e-19
C25754 a_4927_45028# a_n2661_44458# 0.00137f
C25755 a_413_45260# a_n699_43396# 0.100762f
C25756 a_n755_45592# a_8333_44056# 1.1e-19
C25757 a_2382_45260# a_742_44458# 3.78e-19
C25758 a_n1059_45260# a_10057_43914# 6.77e-20
C25759 a_13661_43548# a_13291_42460# 7.75e-21
C25760 a_2324_44458# a_1568_43370# 0.001169f
C25761 a_13017_45260# a_11691_44458# 1.87e-20
C25762 a_2448_45028# a_n2661_43370# 2.21e-19
C25763 a_n2312_39304# a_n1329_42308# 8.42e-20
C25764 a_n2312_40392# a_n961_42308# 2.36e-20
C25765 a_n2293_42834# a_8137_45348# 0.009658f
C25766 a_13556_45296# a_11827_44484# 0.05613f
C25767 a_19692_46634# a_17364_32525# 0.001936f
C25768 a_n743_46660# a_1337_46436# 0.004605f
C25769 a_5807_45002# a_6633_46155# 1.37e-19
C25770 a_n1741_47186# a_12427_45724# 1.48e-19
C25771 a_14976_45028# a_11415_45002# 0.039578f
C25772 a_15227_46910# a_15312_46660# 1.48e-19
C25773 a_171_46873# a_518_46482# 9.21e-19
C25774 a_7715_46873# a_8016_46348# 0.009008f
C25775 a_7577_46660# a_7920_46348# 5.66e-19
C25776 a_4791_45118# a_7227_45028# 0.288276f
C25777 a_6151_47436# a_6194_45824# 0.227219f
C25778 a_19692_46634# a_17639_46660# 2.07e-22
C25779 a_15227_44166# a_19636_46660# 6.47e-19
C25780 a_10249_46116# a_3483_46348# 1.46e-20
C25781 a_7411_46660# a_8349_46414# 0.001959f
C25782 a_n901_43156# a_n4318_38216# 6.06e-21
C25783 a_12545_42858# a_12800_43218# 0.05936f
C25784 a_10341_42308# a_11136_42852# 0.003f
C25785 a_3080_42308# a_n4315_30879# 5.51e-21
C25786 a_22959_44484# VDD 0.303517f
C25787 a_n1853_43023# a_n4318_37592# 1.26e-19
C25788 a_n2157_42858# COMP_P 1.05e-19
C25789 a_n3674_39304# a_n2840_42282# 4.48e-19
C25790 a_17730_32519# RST_Z 0.049818f
C25791 a_12281_43396# a_11323_42473# 3.39e-20
C25792 a_2982_43646# a_21613_42308# 0.001693f
C25793 a_743_42282# a_2123_42473# 0.007332f
C25794 a_n1991_42858# a_n1736_42282# 0.0101f
C25795 a_3539_42460# a_7174_31319# 4.88e-21
C25796 a_n4318_39304# a_n3420_39072# 0.001411f
C25797 a_20692_30879# a_17364_32525# 0.054134f
C25798 a_3090_45724# a_10723_42308# 4.98e-22
C25799 a_n356_44636# a_n23_44458# 0.220577f
C25800 a_5518_44484# a_n2661_43922# 0.011667f
C25801 a_5343_44458# a_n2293_43922# 2.33e-20
C25802 a_10775_45002# a_10729_43914# 1.25e-21
C25803 a_20567_45036# a_20766_44850# 0.001007f
C25804 a_21005_45260# a_20835_44721# 7.06e-20
C25805 a_21101_45002# a_20679_44626# 0.001069f
C25806 a_21359_45002# a_20640_44752# 0.013689f
C25807 a_11827_44484# a_20362_44736# 0.009001f
C25808 a_n2293_42834# a_1467_44172# 9.22e-22
C25809 a_11691_44458# a_19006_44850# 0.005009f
C25810 a_2711_45572# a_16409_43396# 2.45e-19
C25811 a_4185_45028# a_13291_42460# 6.95e-20
C25812 a_n237_47217# VDD 4.05131f
C25813 a_8701_44490# a_9159_44484# 6.03e-19
C25814 a_18911_45144# a_18579_44172# 2.07e-20
C25815 a_18494_42460# a_19279_43940# 0.137363f
C25816 a_n1741_47186# DATA[2] 0.017604f
C25817 a_n2661_43370# a_n1761_44111# 1.12e-20
C25818 a_6298_44484# a_n2661_42834# 0.001263f
C25819 a_n1059_45260# a_14021_43940# 0.008971f
C25820 a_413_45260# a_22959_43948# 0.00133f
C25821 a_n1605_47204# DATA[0] 4.69e-19
C25822 a_n2312_38680# a_n4209_38502# 0.095213f
C25823 a_6419_46155# a_5066_45546# 0.038923f
C25824 a_8492_46660# a_8697_45822# 2.64e-20
C25825 a_n1151_42308# a_n2293_42834# 0.051075f
C25826 a_4791_45118# a_5009_45028# 0.007533f
C25827 a_n443_46116# a_2809_45028# 5.61e-19
C25828 a_n743_46660# a_16789_45572# 1.94e-19
C25829 a_10227_46804# a_13348_45260# 6.18e-19
C25830 a_11599_46634# a_1307_43914# 3.42e-19
C25831 a_765_45546# a_997_45618# 0.026457f
C25832 a_8270_45546# a_10193_42453# 3e-20
C25833 a_16327_47482# a_14537_43396# 3.85e-20
C25834 a_n1613_43370# a_n967_45348# 0.213625f
C25835 a_5807_45002# a_2437_43646# 0.004842f
C25836 a_19594_46812# a_19610_45572# 5.07e-20
C25837 a_3090_45724# a_1990_45572# 2.91e-20
C25838 a_5204_45822# a_5210_46155# 8.95e-19
C25839 a_5164_46348# a_5527_46155# 0.005527f
C25840 a_2324_44458# a_10809_44734# 0.026995f
C25841 a_17583_46090# a_6945_45028# 6.47e-21
C25842 a_18985_46122# a_19335_46494# 0.210876f
C25843 a_18819_46122# a_20075_46420# 0.043567f
C25844 a_1576_42282# a_6123_31319# 2.22e-20
C25845 a_2713_42308# a_3905_42558# 1.81e-21
C25846 a_3318_42354# a_3497_42558# 0.010303f
C25847 a_n1630_35242# a_5934_30871# 0.039258f
C25848 a_1606_42308# a_5932_42308# 0.111585f
C25849 a_1755_42282# a_6171_42473# 0.065035f
C25850 a_5534_30871# a_n3420_38528# 0.041746f
C25851 a_n913_45002# a_1847_42826# 0.294312f
C25852 a_526_44458# a_7174_31319# 4.88e-21
C25853 a_14815_43914# a_11341_43940# 0.001047f
C25854 a_n2661_42834# a_10555_44260# 0.003997f
C25855 a_175_44278# a_453_43940# 0.112594f
C25856 a_17061_44734# a_15682_43940# 1.68e-19
C25857 a_n2661_44458# a_4699_43561# 1.98e-20
C25858 a_1115_44172# a_1467_44172# 0.115277f
C25859 a_644_44056# a_1414_42308# 5.43e-20
C25860 a_8270_45546# VDD 1.26092f
C25861 a_5343_44458# a_n97_42460# 3.84e-19
C25862 a_13259_45724# a_13070_42354# 6.28e-20
C25863 a_n2956_39304# a_n2302_40160# 4.04e-19
C25864 a_n2956_38680# a_n4064_40160# 6.27e-19
C25865 a_n2017_45002# a_2905_42968# 7.95e-20
C25866 a_n967_45348# a_n1533_42852# 0.002483f
C25867 a_n2661_45546# a_1609_45572# 1.69e-19
C25868 a_13059_46348# a_15595_45028# 1.93e-20
C25869 SMPL_ON_P a_n4318_39768# 0.039185f
C25870 a_584_46384# a_895_43940# 0.025246f
C25871 a_n2293_46098# a_n967_45348# 2.05e-20
C25872 a_16327_47482# a_20835_44721# 0.157393f
C25873 a_n743_46660# a_14539_43914# 1.85e-19
C25874 a_11608_46482# a_11652_45724# 2.38e-19
C25875 a_n2497_47436# a_n875_44318# 9.25e-20
C25876 a_22959_46660# a_413_45260# 0.018266f
C25877 a_n1613_43370# a_9159_44484# 3.29e-21
C25878 a_4883_46098# a_17517_44484# 7.99e-22
C25879 a_12861_44030# a_19789_44512# 2.27e-19
C25880 a_n901_46420# a_n1059_45260# 2.16e-20
C25881 a_3877_44458# a_n2661_44458# 0.035165f
C25882 a_6945_45028# a_8696_44636# 4.49e-20
C25883 a_10586_45546# a_12427_45724# 2.09e-19
C25884 a_8049_45260# a_13249_42308# 0.00179f
C25885 a_n863_45724# a_n89_45572# 8.15e-19
C25886 a_n452_45724# a_n310_45572# 0.007833f
C25887 a_n755_45592# a_n443_42852# 0.469263f
C25888 a_n4064_39616# a_n2860_39866# 0.003766f
C25889 a_3160_47472# a_n1151_42308# 0.357683f
C25890 a_2905_45572# a_3381_47502# 0.208262f
C25891 a_2063_45854# a_4007_47204# 3.64e-20
C25892 a_n971_45724# a_7227_47204# 0.009537f
C25893 a_n237_47217# a_6491_46660# 0.002119f
C25894 a_n1741_47186# a_11031_47542# 0.00728f
C25895 a_2952_47436# a_3785_47178# 6.47e-19
C25896 a_n2497_47436# a_n1435_47204# 0.010029f
C25897 a_n4064_40160# a_n3690_39392# 3.42e-19
C25898 a_7174_31319# a_n4209_38502# 5.81e-22
C25899 a_14097_32519# C4_N_btm 0.030945f
C25900 a_n1630_35242# a_11530_34132# 0.029967f
C25901 a_5742_30871# VDAC_Ni 3.56e-19
C25902 a_14539_43914# a_17701_42308# 0.039977f
C25903 a_n2661_42282# a_6197_43396# 0.033187f
C25904 a_n356_44636# a_12089_42308# 5.58e-20
C25905 a_5111_44636# a_8685_42308# 3.87e-21
C25906 a_n1059_45260# a_15764_42576# 4.65e-19
C25907 a_n2017_45002# a_15803_42450# 0.005056f
C25908 a_n913_45002# a_15486_42560# 2.61e-19
C25909 a_20692_30879# a_21589_35634# 4.41e-20
C25910 a_8375_44464# a_8037_42858# 4.44e-20
C25911 a_5891_43370# a_7765_42852# 0.168516f
C25912 a_12638_46436# VDD 0.002311f
C25913 a_9165_43940# a_9420_43940# 0.005172f
C25914 a_742_44458# a_1709_42852# 0.001488f
C25915 a_n755_45592# a_375_42282# 0.366231f
C25916 a_n863_45724# a_2304_45348# 0.091195f
C25917 a_n357_42282# a_501_45348# 1.02e-19
C25918 a_n443_42852# a_13017_45260# 2.72e-20
C25919 a_12549_44172# a_21381_43940# 0.099617f
C25920 a_8049_45260# a_17613_45144# 1.7e-20
C25921 a_11415_45002# a_15433_44458# 1.94e-20
C25922 a_15765_45572# a_16147_45260# 0.005068f
C25923 a_10193_42453# a_n2017_45002# 0.081859f
C25924 a_n1613_43370# a_n1917_43396# 0.153085f
C25925 a_4915_47217# a_14579_43548# 2.85e-21
C25926 a_2324_44458# a_5883_43914# 0.002714f
C25927 a_n2661_45546# a_4185_45348# 1.35e-19
C25928 a_4099_45572# a_3232_43370# 2.19e-22
C25929 a_3483_46348# a_5205_44734# 3.63e-20
C25930 a_19692_46634# a_19237_31679# 4.44e-20
C25931 a_16115_45572# a_16377_45572# 0.001705f
C25932 a_16680_45572# a_16842_45938# 0.006453f
C25933 a_12741_44636# a_13857_44734# 0.003456f
C25934 a_3775_45552# a_3065_45002# 3.53e-20
C25935 a_2711_45572# a_6431_45366# 0.001609f
C25936 a_10903_43370# a_13720_44458# 2.88e-20
C25937 a_8128_46384# a_2107_46812# 0.028382f
C25938 a_n237_47217# a_10185_46660# 7.66e-20
C25939 a_12861_44030# a_6755_46942# 0.376009f
C25940 a_n4209_37414# C5_P_btm 1.11e-20
C25941 a_n3565_37414# C7_P_btm 1.43e-20
C25942 a_10227_46804# a_7411_46660# 2.95e-22
C25943 a_11599_46634# a_10467_46802# 0.261176f
C25944 a_n4064_37984# VIN_P 0.06139f
C25945 a_5807_45002# a_n2661_46634# 0.087532f
C25946 a_5088_37509# a_n923_35174# 7.48e-20
C25947 a_n1741_47186# a_12347_46660# 2.12e-19
C25948 a_2747_46873# a_2864_46660# 0.174836f
C25949 VDAC_Pi RST_Z 0.002358f
C25950 a_n3565_38216# VCM 0.03544f
C25951 a_4883_46098# a_5167_46660# 1.64e-20
C25952 CAL_N a_22609_37990# 4.7e-20
C25953 a_22780_40081# a_22469_39537# 1.28e-20
C25954 a_22521_40055# a_22876_39857# 4.84e-19
C25955 a_22469_40625# a_22609_38406# 0.066321f
C25956 a_22521_40599# a_22705_38406# 0.008755f
C25957 a_22521_39511# a_22821_38993# 0.112629f
C25958 a_n1613_43370# a_1110_47026# 6.37e-19
C25959 a_6151_47436# a_8601_46660# 6.03e-19
C25960 a_n1151_42308# a_13607_46688# 0.005534f
C25961 a_2952_47436# a_3090_45724# 8.88e-21
C25962 a_n881_46662# a_n935_46688# 8.8e-19
C25963 a_n3420_37984# VREF 1.33e-19
C25964 a_14021_43940# a_19987_42826# 1.06e-19
C25965 a_n1917_43396# a_n1533_42852# 1.04e-19
C25966 a_3357_43084# CLK 2.63944f
C25967 a_9313_44734# a_15890_42674# 1.49e-20
C25968 a_n1761_44111# COMP_P 2.35e-19
C25969 a_2982_43646# a_4361_42308# 0.545077f
C25970 a_n356_44636# a_18907_42674# 2.06e-20
C25971 a_n2017_45002# VDD 3.8321f
C25972 a_8685_43396# a_16759_43396# 1.34e-19
C25973 a_n1809_43762# a_n3674_39304# 9.24e-22
C25974 a_n2012_43396# a_n4318_38680# 1.79e-19
C25975 a_14579_43548# a_15681_43442# 9.87e-22
C25976 a_14358_43442# a_14621_43646# 0.011552f
C25977 a_14205_43396# a_14537_43646# 3.88e-19
C25978 a_n2293_43922# a_12563_42308# 0.015547f
C25979 a_n971_45724# a_n3674_37592# 0.022388f
C25980 a_3483_46348# a_13565_43940# 0.006953f
C25981 a_2711_45572# a_16241_44734# 0.03035f
C25982 a_5691_45260# a_5837_45348# 0.013377f
C25983 a_12549_44172# a_18249_42858# 4.15e-20
C25984 a_3090_45724# a_10341_43396# 0.07129f
C25985 a_14180_45002# a_14797_45144# 0.070624f
C25986 a_3065_45002# a_5093_45028# 1.41e-21
C25987 a_n2956_37592# a_n2661_43370# 0.044152f
C25988 a_21188_45572# a_21359_45002# 4.16e-19
C25989 a_21363_45546# a_11827_44484# 1.3e-22
C25990 a_20731_45938# a_21005_45260# 2.73e-20
C25991 a_10227_46804# a_11229_43218# 0.001903f
C25992 a_n2293_46634# a_9127_43156# 1.56e-19
C25993 a_13661_43548# a_13460_43230# 7.36e-20
C25994 a_20692_30879# a_19237_31679# 0.051625f
C25995 a_10490_45724# a_9313_44734# 4.22e-21
C25996 a_8696_44636# a_8103_44636# 1.41e-19
C25997 a_13556_45296# a_15595_45028# 1.42e-20
C25998 a_13348_45260# a_1307_43914# 3.41e-21
C25999 a_n2497_47436# a_380_45546# 9.69e-22
C26000 a_12549_44172# a_10903_43370# 0.792848f
C26001 a_12891_46348# a_12005_46116# 0.001509f
C26002 SMPL_ON_P a_n2956_38216# 0.0385f
C26003 a_n743_46660# a_1823_45246# 0.04372f
C26004 a_n1925_46634# a_167_45260# 3.51e-19
C26005 a_5807_45002# a_8199_44636# 0.001797f
C26006 a_6755_46942# a_14180_46812# 0.063843f
C26007 a_13607_46688# a_14084_46812# 0.014875f
C26008 a_n2438_43548# a_1138_42852# 0.646257f
C26009 a_n133_46660# a_1176_45822# 3.41e-19
C26010 a_n2293_46634# a_2804_46116# 1.38e-20
C26011 a_12861_44030# a_8049_45260# 0.109405f
C26012 a_n881_46662# a_2324_44458# 0.085939f
C26013 a_383_46660# a_376_46348# 3.44e-19
C26014 a_33_46660# a_805_46414# 0.001417f
C26015 a_n815_47178# a_n2661_45546# 4.98e-21
C26016 a_n2312_40392# a_n2956_39304# 0.052343f
C26017 a_5257_43370# a_765_45546# 0.002074f
C26018 a_4915_47217# a_12839_46116# 2.59e-20
C26019 a_n97_42460# a_12563_42308# 0.001953f
C26020 a_2982_43646# a_6761_42308# 3.92e-20
C26021 a_3422_30871# VDAC_N 0.480069f
C26022 a_12379_42858# a_12089_42308# 0.16885f
C26023 a_10341_42308# a_12545_42858# 9.44e-20
C26024 a_n89_44484# VDD 6.07e-19
C26025 a_3539_42460# a_5932_42308# 4.34e-21
C26026 a_3483_46348# a_5534_30871# 2.26e-20
C26027 a_11691_44458# a_18374_44850# 0.02267f
C26028 a_19113_45348# a_18989_43940# 3.13e-19
C26029 a_n2312_39304# a_n4334_39392# 3.7e-20
C26030 a_n443_42852# a_548_43396# 2.03e-19
C26031 a_n2661_44458# a_10440_44484# 0.005733f
C26032 a_16751_45260# a_11967_42832# 1.76e-21
C26033 a_18175_45572# a_18451_43940# 6.66e-21
C26034 a_n1059_45260# a_5013_44260# 2e-20
C26035 a_n2017_45002# a_5495_43940# 8.92e-22
C26036 a_8953_45546# a_8952_43230# 0.01883f
C26037 a_8199_44636# a_10518_42984# 7.84e-20
C26038 a_5257_43370# a_4921_42308# 0.002713f
C26039 a_n913_45002# a_5244_44056# 1.75e-21
C26040 a_2779_44458# a_n699_43396# 0.025176f
C26041 a_2107_46812# a_10053_45546# 1.1e-19
C26042 a_11415_45002# a_19900_46494# 1.14e-20
C26043 a_20202_43084# a_20708_46348# 0.001267f
C26044 a_765_45546# a_1337_46116# 0.011452f
C26045 a_3483_46348# a_5937_45572# 0.767636f
C26046 a_14976_45028# a_13259_45724# 0.018965f
C26047 a_21350_47026# a_10809_44734# 1.68e-19
C26048 a_4817_46660# a_2711_45572# 9.24e-20
C26049 a_n237_47217# a_5691_45260# 2.17e-21
C26050 a_n971_45724# a_6171_45002# 0.030962f
C26051 a_14180_46812# a_8049_45260# 1.24e-21
C26052 a_n1151_42308# a_413_45260# 0.135643f
C26053 a_n881_46662# a_16855_45546# 0.052296f
C26054 a_4883_46098# a_19256_45572# 1.02e-20
C26055 a_18479_47436# a_20107_45572# 0.025968f
C26056 a_16327_47482# a_20731_45938# 0.012637f
C26057 a_14311_47204# a_2437_43646# 0.00629f
C26058 a_3877_44458# a_5907_45546# 4.21e-21
C26059 a_n743_46660# a_12427_45724# 1.63e-20
C26060 a_5164_46348# a_6165_46155# 3.3e-19
C26061 a_5204_45822# a_5497_46414# 0.099282f
C26062 a_12549_44172# a_12016_45572# 7.31e-20
C26063 a_10227_46804# a_20841_45814# 3.53e-19
C26064 a_11453_44696# a_18175_45572# 0.036949f
C26065 a_13717_47436# a_3357_43084# 0.024679f
C26066 a_584_46384# a_3065_45002# 0.085314f
C26067 a_n4318_38680# a_n4064_39616# 0.021342f
C26068 a_21845_43940# VDD 0.00416f
C26069 a_17538_32519# RST_Z 0.050782f
C26070 a_4190_30871# a_n3420_38528# 0.031855f
C26071 a_526_44458# a_5932_42308# 3.79e-19
C26072 a_9290_44172# a_13657_42308# 1.07e-19
C26073 a_n2293_42834# a_n1809_43762# 0.001769f
C26074 a_19615_44636# a_18579_44172# 0.158449f
C26075 a_19006_44850# a_18753_44484# 4.61e-19
C26076 a_n743_46660# DATA[2] 1.69e-21
C26077 a_10193_42453# a_19164_43230# 0.003383f
C26078 a_5111_44636# a_9803_43646# 0.118936f
C26079 a_n133_46660# DATA[0] 1.6e-19
C26080 a_n2438_43548# DATA[1] 5.69e-20
C26081 a_1123_46634# VDD 0.469393f
C26082 a_n2661_43922# a_2127_44172# 0.007786f
C26083 a_n2661_42834# a_2479_44172# 0.027713f
C26084 a_n2293_46634# CLK 1.2e-20
C26085 a_n2017_45002# a_16137_43396# 0.63011f
C26086 a_20640_44752# a_19279_43940# 0.22152f
C26087 a_20679_44626# a_20766_44850# 0.052825f
C26088 a_375_42282# a_548_43396# 6.62e-19
C26089 a_n2661_43370# a_n2267_43396# 0.001687f
C26090 a_11387_46155# a_11652_45724# 1.9e-19
C26091 a_19321_45002# a_21359_45002# 4.39e-19
C26092 a_13747_46662# a_22223_45036# 2.35e-19
C26093 a_12549_44172# a_19929_45028# 3.72e-20
C26094 a_18597_46090# a_18287_44626# 6.68e-22
C26095 a_10903_43370# a_11525_45546# 0.040993f
C26096 a_12005_46116# a_11322_45546# 2.36e-19
C26097 a_16375_45002# a_19240_46482# 3.8e-20
C26098 a_8128_46384# a_n2661_44458# 1.73e-21
C26099 a_11453_44696# a_10440_44484# 4.13e-20
C26100 a_12465_44636# a_12883_44458# 0.017889f
C26101 a_6945_45028# a_7227_45028# 0.016808f
C26102 a_9290_44172# a_11823_42460# 0.864145f
C26103 a_2324_44458# a_8162_45546# 4.52e-20
C26104 a_6755_46942# a_11787_45002# 9.54e-22
C26105 a_11189_46129# a_12427_45724# 1.25e-19
C26106 a_12594_46348# a_10490_45724# 9.79e-19
C26107 a_5807_45002# a_19113_45348# 9.15e-19
C26108 a_3483_46348# a_8697_45572# 7.8e-19
C26109 a_14035_46660# a_3357_43084# 2.73e-20
C26110 a_n1613_43370# a_n1917_44484# 0.153277f
C26111 a_6123_31319# a_1736_39043# 6.11e-20
C26112 a_5534_30871# VIN_N 0.00357f
C26113 a_19164_43230# VDD 0.278643f
C26114 a_18727_42674# a_18907_42674# 0.185422f
C26115 a_n967_45348# a_n1736_42282# 0.001893f
C26116 a_453_43940# a_n97_42460# 2.8e-19
C26117 a_14815_43914# a_10341_43396# 8.2e-20
C26118 a_10193_42453# a_21973_42336# 3.78e-21
C26119 a_n913_45002# a_n473_42460# 7.7e-21
C26120 a_n1059_45260# a_196_42282# 4.1e-19
C26121 a_n2017_45002# a_n784_42308# 0.0226f
C26122 a_n809_44244# a_n229_43646# 0.001748f
C26123 a_9313_44734# a_16547_43609# 0.010576f
C26124 a_n699_43396# a_n13_43084# 0.001012f
C26125 a_9625_46129# CLK 2.09e-20
C26126 en_comp a_n4318_37592# 0.03345f
C26127 a_n2956_37592# COMP_P 1.39e-21
C26128 a_14539_43914# a_4361_42308# 2.29e-20
C26129 a_3422_30871# a_3626_43646# 1.22e-19
C26130 a_13759_46122# VDD 0.399995f
C26131 a_3357_43084# a_1755_42282# 4.76e-20
C26132 a_2324_44458# a_11361_45348# 1.97e-19
C26133 a_11525_45546# a_12016_45572# 0.00278f
C26134 a_n1641_46494# a_n2661_44458# 1.32e-20
C26135 a_3090_45724# a_n2293_43922# 0.02667f
C26136 SMPL_ON_N a_14021_43940# 1.94e-20
C26137 a_584_46384# a_458_43396# 0.196763f
C26138 a_12861_44030# a_15037_43940# 1.65e-19
C26139 a_n755_45592# a_2437_43646# 0.017992f
C26140 a_526_44458# a_1423_45028# 0.133656f
C26141 a_11962_45724# a_11688_45572# 2.07e-20
C26142 a_11652_45724# a_11778_45572# 0.001094f
C26143 a_n1991_46122# a_n2129_44697# 2.79e-21
C26144 a_n1853_46287# a_n2267_44484# 1.43e-21
C26145 a_n2438_43548# a_n4318_39768# 6.52e-19
C26146 a_3483_46348# a_11691_44458# 0.039125f
C26147 a_4185_45028# a_22959_45036# 0.17601f
C26148 a_12549_44172# a_14955_43940# 0.010132f
C26149 a_768_44030# a_13483_43940# 0.002743f
C26150 a_n2661_45546# a_n2661_45010# 0.014492f
C26151 a_4883_46098# a_12549_44172# 0.021771f
C26152 a_16241_47178# a_16750_47204# 2.6e-19
C26153 a_6151_47436# a_2107_46812# 0.019997f
C26154 a_7754_38636# VDAC_Ni 1.97e-19
C26155 a_n4209_39304# C7_P_btm 0.184297f
C26156 a_10227_46804# a_13661_43548# 0.072131f
C26157 a_17591_47464# a_13747_46662# 1.16e-19
C26158 a_18143_47464# a_5807_45002# 1.77e-19
C26159 a_n237_47217# a_4646_46812# 0.020773f
C26160 a_n1151_42308# a_2609_46660# 3.74e-19
C26161 a_3381_47502# a_2443_46660# 8.51e-19
C26162 a_2905_45572# a_2959_46660# 0.005466f
C26163 a_3160_47472# a_3177_46902# 0.009123f
C26164 a_2063_45854# a_2864_46660# 0.002177f
C26165 a_n971_45724# a_4955_46873# 4.2e-20
C26166 a_22465_38105# RST_Z 0.034434f
C26167 a_n3565_39304# C9_P_btm 1.64e-19
C26168 a_6197_43396# a_7112_43396# 0.118423f
C26169 a_3539_42460# a_4181_43396# 3.38e-21
C26170 a_n2661_42834# a_n2104_42282# 3.95e-21
C26171 a_11967_42832# a_13291_42460# 0.015813f
C26172 a_n2661_43922# a_n4318_38216# 5.64e-19
C26173 a_18184_42460# a_18214_42558# 0.056496f
C26174 a_18494_42460# a_19332_42282# 0.040916f
C26175 a_16922_45042# a_20712_42282# 2.62e-20
C26176 a_n2956_37592# a_n3565_37414# 0.304738f
C26177 a_9028_43914# a_8952_43230# 6.18e-20
C26178 a_9672_43914# a_9127_43156# 0.001066f
C26179 a_2479_44172# a_n2293_42282# 0.059476f
C26180 a_n356_44636# a_5267_42460# 1.4e-19
C26181 a_n2293_43922# a_n2472_42282# 1.85e-19
C26182 a_n2810_45028# a_n3690_37440# 5.77e-19
C26183 a_14021_43940# a_22959_43396# 0.191956f
C26184 a_13259_45724# a_15433_44458# 2.36e-21
C26185 a_n913_45002# a_5111_44636# 0.070773f
C26186 a_10227_46804# a_10835_43094# 0.295543f
C26187 a_n1151_42308# a_n914_42852# 1.43e-19
C26188 a_14495_45572# a_11691_44458# 2.65e-20
C26189 a_413_45260# a_327_44734# 0.195096f
C26190 a_n37_45144# a_1667_45002# 1.12e-20
C26191 a_n1613_43370# a_n1853_43023# 0.423772f
C26192 a_n356_45724# a_n356_44636# 0.001699f
C26193 a_3090_45724# a_n97_42460# 0.001209f
C26194 a_12741_44636# a_15493_43940# 2.5e-19
C26195 a_12549_44172# a_5649_42852# 9.86e-20
C26196 a_13661_43548# a_19177_43646# 0.015951f
C26197 a_3483_46348# a_8333_44056# 5.87e-19
C26198 a_7927_46660# a_8492_46660# 7.99e-20
C26199 a_n1435_47204# a_9569_46155# 2.34e-20
C26200 a_10227_46804# a_4185_45028# 3.04e-19
C26201 a_n2497_47436# a_526_44458# 0.06857f
C26202 a_n443_46116# a_2324_44458# 0.055032f
C26203 a_4646_46812# a_8270_45546# 1.8e-19
C26204 a_9313_45822# a_9290_44172# 4.81e-22
C26205 a_11031_47542# a_11189_46129# 8.25e-21
C26206 a_13661_43548# a_17339_46660# 0.599051f
C26207 a_5807_45002# a_765_45546# 0.103324f
C26208 a_n2312_39304# a_n1853_46287# 3.91e-19
C26209 a_16137_43396# a_19164_43230# 9.01e-19
C26210 a_17324_43396# a_17701_42308# 0.00643f
C26211 a_17499_43370# a_18083_42858# 0.003663f
C26212 a_743_42282# a_9127_43156# 2.23e-19
C26213 a_n1917_43396# a_n1736_42282# 7.84e-20
C26214 a_n2840_44458# VDD 0.247948f
C26215 a_5649_42852# a_5111_42852# 0.110096f
C26216 a_n1641_43230# a_n1379_43218# 0.001705f
C26217 a_n1423_42826# a_n967_43230# 4.2e-19
C26218 a_15743_43084# a_15567_42826# 0.215954f
C26219 a_19721_31679# RST_Z 0.050546f
C26220 a_n1699_43638# a_n4318_37592# 9.74e-21
C26221 a_n2267_43396# COMP_P 8.07e-20
C26222 a_4361_42308# a_7871_42858# 6.79e-20
C26223 a_n2293_42834# a_4223_44672# 0.015649f
C26224 a_6171_45002# a_9313_44734# 2.05e-20
C26225 a_19778_44110# a_11827_44484# 0.029054f
C26226 a_18494_42460# a_21101_45002# 1.76e-20
C26227 a_2680_45002# a_n2661_42834# 6.24e-21
C26228 a_2382_45260# a_n2661_43922# 0.026472f
C26229 a_10193_42453# a_18079_43940# 0.076581f
C26230 a_21188_45572# a_19279_43940# 3.06e-19
C26231 a_20731_45938# a_20835_44721# 8.44e-21
C26232 a_19692_46634# a_19987_42826# 5.42e-19
C26233 a_768_44030# a_6123_31319# 1.76e-21
C26234 a_12861_44030# a_13258_32519# 9.87e-21
C26235 a_n2661_43370# a_n2267_44484# 0.007573f
C26236 a_21513_45002# a_11967_42832# 5.76e-19
C26237 a_1823_45246# a_4361_42308# 0.11884f
C26238 a_n2293_46634# a_1755_42282# 7.99e-22
C26239 a_5837_45028# a_5518_44484# 1.43e-19
C26240 a_8191_45002# a_8375_44464# 9.04e-19
C26241 a_20567_45036# a_21005_45260# 0.015494f
C26242 a_17719_45144# a_11691_44458# 2.64e-20
C26243 a_11823_42460# a_10807_43548# 4.89e-19
C26244 a_10227_46804# a_16269_42308# 1.79e-19
C26245 a_16327_47482# a_18727_42674# 0.003774f
C26246 w_1575_34946# a_n4064_37440# 3.26e-19
C26247 a_11599_46634# a_11682_45822# 7.01e-19
C26248 a_n1925_46634# a_n863_45724# 5.47e-20
C26249 a_n2293_46634# a_n1099_45572# 0.006391f
C26250 a_12359_47026# a_12005_46116# 1.79e-19
C26251 a_n881_46662# a_6667_45809# 0.006711f
C26252 a_22591_46660# a_21076_30879# 3.06e-19
C26253 a_n1613_43370# a_6598_45938# 0.009561f
C26254 a_n743_46660# a_n2293_45546# 6.76e-20
C26255 a_171_46873# a_n2661_45546# 7.37e-21
C26256 a_n2438_43548# a_n2956_38216# 0.020852f
C26257 a_15227_44166# a_15015_46420# 1.48e-19
C26258 a_11309_47204# a_2711_45572# 1.1e-19
C26259 a_16292_46812# a_15682_46116# 0.005299f
C26260 a_20820_30879# a_22959_46660# 0.01739f
C26261 a_n1021_46688# a_n1079_45724# 4.95e-21
C26262 a_7411_46660# a_8034_45724# 6.76e-21
C26263 a_5257_43370# a_6347_46155# 2.62e-19
C26264 a_3090_45724# a_17957_46116# 1.57e-19
C26265 a_11813_46116# a_6945_45028# 1.65e-19
C26266 a_11186_47026# a_10809_44734# 3.59e-20
C26267 a_20202_43084# a_21542_46660# 7.08e-19
C26268 a_n2661_46634# a_n755_45592# 4.56e-20
C26269 a_16823_43084# a_17531_42308# 1.38e-20
C26270 a_18079_43940# VDD 0.162408f
C26271 a_19700_43370# a_13258_32519# 1.55e-20
C26272 a_15743_43084# a_20712_42282# 4.16e-20
C26273 a_4361_42308# a_11897_42308# 3.73e-19
C26274 a_n2293_42282# a_n2104_42282# 0.058363f
C26275 a_743_42282# a_17124_42282# 0.007228f
C26276 a_7227_42852# a_7227_42308# 3.59e-19
C26277 a_18374_44850# a_18753_44484# 3.16e-19
C26278 a_949_44458# a_1414_42308# 0.009641f
C26279 a_n2661_44458# a_5244_44056# 1.12e-20
C26280 a_22612_30879# a_22521_40055# 4.85e-20
C26281 a_21588_30879# a_22459_39145# 6.4e-20
C26282 a_12465_44636# START 0.065727f
C26283 a_22223_47212# RST_Z 2.25e-19
C26284 a_9313_44734# a_14673_44172# 6.42e-20
C26285 a_n699_43396# a_644_44056# 1.32e-19
C26286 a_n913_45002# a_4235_43370# 9.46e-20
C26287 a_n1059_45260# a_4699_43561# 1.87e-20
C26288 a_n2017_45002# a_3080_42308# 0.034898f
C26289 a_n357_42282# a_5534_30871# 0.04831f
C26290 a_1307_43914# a_5829_43940# 0.016223f
C26291 a_2274_45254# a_n97_42460# 6.35e-21
C26292 a_742_44458# a_453_43940# 0.001956f
C26293 a_21811_47423# SINGLE_ENDED 0.215228f
C26294 a_4185_45028# a_4933_42558# 0.001444f
C26295 a_n443_42852# a_10083_42826# 5.44e-19
C26296 a_22731_47423# VDD 0.196667f
C26297 a_5066_45546# a_5527_46155# 8.1e-19
C26298 a_n2661_46634# a_13017_45260# 0.123713f
C26299 a_n2293_46634# a_10951_45334# 3.22e-21
C26300 a_3483_46348# a_n443_42852# 1.96e-19
C26301 a_1176_45822# a_1176_45572# 0.001923f
C26302 a_765_45546# a_15143_45578# 1.48e-21
C26303 a_n2312_39304# a_n2661_43370# 1.64e-20
C26304 a_18985_46122# a_19240_46482# 0.05936f
C26305 a_18189_46348# a_18051_46116# 0.045453f
C26306 a_18819_46122# a_19431_46494# 3.82e-19
C26307 a_19553_46090# a_16375_45002# 2.34e-20
C26308 a_8199_44636# a_n755_45592# 5.59e-20
C26309 a_5937_45572# a_n357_42282# 1.32e-19
C26310 a_n1925_46634# a_8191_45002# 9.69e-19
C26311 a_n2293_46098# a_6598_45938# 8.22e-20
C26312 a_3177_46902# a_413_45260# 0.006595f
C26313 a_6151_47436# a_n2661_44458# 3.69e-21
C26314 a_15227_44166# a_16333_45814# 4.01e-21
C26315 a_4646_46812# a_n2017_45002# 5.44e-19
C26316 a_2107_46812# a_5111_44636# 7.67e-20
C26317 a_3090_45724# a_16020_45572# 0.001921f
C26318 a_12861_44030# a_20193_45348# 0.680394f
C26319 a_5807_45002# a_16751_45260# 0.001196f
C26320 a_13661_43548# a_1307_43914# 0.396211f
C26321 a_16327_47482# a_20567_45036# 0.009073f
C26322 a_22591_43396# RST_Z 3.24e-19
C26323 a_4190_30871# VIN_N 0.049977f
C26324 a_11323_42473# a_11551_42558# 0.062483f
C26325 a_5342_30871# VDAC_P 0.007514f
C26326 a_14209_32519# VDD 0.284433f
C26327 a_n3674_38216# a_n4334_39616# 9.11e-20
C26328 a_17364_32525# C10_N_btm 1.08e-19
C26329 a_5534_30871# CAL_N 0.004303f
C26330 a_n356_44636# a_6547_43396# 9.65e-22
C26331 a_5891_43370# a_2982_43646# 5.95e-19
C26332 a_1307_43914# a_10835_43094# 3.58e-20
C26333 a_n2293_42834# a_n3674_39304# 1.76e-19
C26334 a_10440_44484# a_9145_43396# 2.03e-20
C26335 a_13720_44458# a_8685_43396# 1.78e-22
C26336 a_10334_44484# a_9803_43646# 5.26e-20
C26337 a_n357_42282# a_19647_42308# 7.07e-20
C26338 a_n2661_42834# a_n229_43646# 0.001251f
C26339 a_7499_43078# a_8791_42308# 0.001313f
C26340 a_2382_45260# a_3445_43172# 1.08e-19
C26341 a_16922_45042# a_20556_43646# 0.00844f
C26342 a_1823_45246# a_2809_45348# 2.74e-19
C26343 a_9823_46155# a_8953_45002# 5.32e-19
C26344 a_n881_46662# a_n1761_44111# 6.91e-21
C26345 a_n1613_43370# a_n1899_43946# 0.038349f
C26346 a_2711_45572# a_10490_45724# 0.036939f
C26347 a_6472_45840# a_7499_43078# 2.82e-21
C26348 a_6667_45809# a_8162_45546# 1.87e-19
C26349 a_19553_46090# a_413_45260# 4.37e-21
C26350 a_2324_44458# a_3537_45260# 0.015845f
C26351 a_8270_45546# a_10057_43914# 3.3e-19
C26352 a_20916_46384# a_20640_44752# 9.21e-22
C26353 a_19321_45002# a_19279_43940# 0.019898f
C26354 a_18051_46116# a_17478_45572# 6.12e-19
C26355 a_13661_43548# a_18579_44172# 0.229269f
C26356 a_12594_46348# a_6171_45002# 4.26e-20
C26357 a_4185_45028# a_1307_43914# 0.025209f
C26358 a_13259_45724# a_13385_45572# 8.8e-20
C26359 a_17339_46660# a_18587_45118# 0.003347f
C26360 a_n1925_42282# a_3357_43084# 0.067793f
C26361 a_13717_47436# a_18597_46090# 1.1e-19
C26362 a_n237_47217# a_9804_47204# 3.49e-19
C26363 a_1239_47204# a_n881_46662# 8.4e-19
C26364 a_1431_47204# a_n1613_43370# 4.26e-19
C26365 a_3160_47472# a_3315_47570# 0.005289f
C26366 a_3815_47204# a_2747_46873# 2.57e-20
C26367 a_n4315_30879# a_n4064_37440# 0.035563f
C26368 a_15673_47210# a_16023_47582# 0.228897f
C26369 a_6575_47204# a_4883_46098# 7.51e-20
C26370 a_12861_44030# a_18780_47178# 9.61e-19
C26371 a_1343_38525# a_3754_39134# 1.67e-19
C26372 a_n4209_39590# a_n4209_37414# 0.031971f
C26373 a_5742_30871# C0_dummy_P_btm 2.87e-19
C26374 a_7174_31319# VDAC_N 0.006565f
C26375 a_n3420_38528# a_n3420_37984# 0.113087f
C26376 a_n3565_38502# a_n4064_37984# 0.028083f
C26377 a_n4064_38528# a_n3565_38216# 0.028041f
C26378 a_n4064_40160# a_n3420_37440# 0.062634f
C26379 a_16241_47178# a_16327_47482# 0.185907f
C26380 a_14955_47212# a_10227_46804# 0.175517f
C26381 a_15507_47210# a_16588_47582# 0.102325f
C26382 a_11599_46634# a_17591_47464# 1.03e-20
C26383 a_19647_42308# CAL_N 0.001755f
C26384 a_5891_43370# a_5837_42852# 0.010625f
C26385 en_comp a_1343_38525# 0.038003f
C26386 a_n2956_37592# a_n4209_39304# 0.102982f
C26387 a_n1352_43396# a_n229_43646# 2.37e-19
C26388 a_11341_43940# a_12281_43396# 0.002178f
C26389 a_15682_43940# a_16409_43396# 0.007432f
C26390 a_11967_42832# a_13460_43230# 0.038517f
C26391 a_4099_45572# VDD 0.296272f
C26392 a_15493_43396# a_15781_43660# 0.047833f
C26393 a_18079_43940# a_16137_43396# 1.32e-20
C26394 a_n357_42282# a_11691_44458# 2.63e-20
C26395 a_15227_44166# a_15493_43396# 0.046514f
C26396 a_20623_45572# a_20719_45572# 0.013793f
C26397 a_20841_45814# a_20885_45572# 3.69e-19
C26398 a_20273_45572# a_21513_45002# 2.44e-19
C26399 a_20107_45572# a_2437_43646# 3.54e-19
C26400 a_8049_45260# a_18287_44626# 1.03e-20
C26401 a_4185_45028# a_18579_44172# 1.48e-22
C26402 a_18479_45785# a_n2017_45002# 8.68e-20
C26403 a_15037_45618# a_6171_45002# 6.48e-20
C26404 a_10227_46804# a_15037_43396# 0.002187f
C26405 a_7227_45028# a_7735_45067# 1.1e-19
C26406 a_6511_45714# a_n2661_43370# 6.25e-20
C26407 a_12549_44172# a_8685_43396# 3.53e-19
C26408 C3_P_btm C2_N_btm 1.05e-19
C26409 C1_P_btm C0_N_btm 2.85e-19
C26410 C0_P_btm C0_dummy_N_btm 1.93e-19
C26411 C4_P_btm C3_N_btm 2.12e-19
C26412 a_1799_45572# a_3524_46660# 1.24e-20
C26413 a_11453_44696# a_19466_46812# 0.004642f
C26414 a_16023_47582# a_16388_46812# 0.001491f
C26415 a_16327_47482# a_16721_46634# 7.05e-19
C26416 a_n743_46660# a_5732_46660# 1.15e-21
C26417 a_2107_46812# a_3221_46660# 6.44e-19
C26418 a_19120_35138# VDD 0.318963f
C26419 a_n2109_47186# a_2202_46116# 6.76e-21
C26420 a_9804_47204# a_8270_45546# 4.96e-19
C26421 a_n881_46662# a_11186_47026# 1.85e-19
C26422 a_12861_44030# a_18285_46348# 0.247326f
C26423 a_13717_47436# a_19123_46287# 4.43e-21
C26424 a_n1741_47186# a_1138_42852# 1.21e-20
C26425 a_n746_45260# a_n1076_46494# 5.44e-19
C26426 a_5807_45002# a_10623_46897# 0.005882f
C26427 a_n1925_46634# a_5072_46660# 0.001838f
C26428 a_2443_46660# a_2959_46660# 0.110816f
C26429 a_2609_46660# a_3177_46902# 0.17072f
C26430 a_14311_47204# a_765_45546# 0.003681f
C26431 a_n2661_42282# a_2903_42308# 2.11e-19
C26432 a_15743_43084# a_20556_43646# 2.78e-21
C26433 a_19268_43646# a_743_42282# 7.11e-21
C26434 a_2982_43646# a_17595_43084# 3.45e-20
C26435 a_7845_44172# a_6123_31319# 1.02e-21
C26436 a_17324_43396# a_4361_42308# 8.49e-21
C26437 a_19692_46634# a_22959_43396# 9.22e-20
C26438 a_n2956_38680# a_n4318_39304# 0.023179f
C26439 a_15037_45618# a_14673_44172# 1.11e-21
C26440 a_n37_45144# a_n699_43396# 4.14e-19
C26441 a_5111_44636# a_n2661_44458# 0.048314f
C26442 a_n357_42282# a_8333_44056# 6.5e-22
C26443 a_n913_45002# a_10334_44484# 2.34e-21
C26444 a_n1059_45260# a_10440_44484# 7.97e-22
C26445 a_n2017_45002# a_10057_43914# 5.16e-20
C26446 a_5807_45002# a_13291_42460# 5.69e-21
C26447 a_12549_44172# a_15953_42852# 9.14e-21
C26448 a_11963_45334# a_11691_44458# 1.33e-19
C26449 a_117_45144# a_n2661_43370# 4.07e-19
C26450 a_n443_42852# a_261_44278# 2.42e-19
C26451 a_n2312_39304# COMP_P 0.00156f
C26452 a_n2312_40392# a_n1329_42308# 4e-20
C26453 a_4185_45028# a_9396_43370# 7.23e-21
C26454 a_8696_44636# a_15463_44811# 3.4e-19
C26455 a_1667_45002# a_949_44458# 0.008156f
C26456 a_9482_43914# a_11827_44484# 0.031913f
C26457 a_9290_44172# a_2982_43646# 0.001406f
C26458 a_16375_45002# a_15493_43940# 2.37e-20
C26459 w_1575_34946# a_n3420_39072# 0.023412f
C26460 a_5807_45002# a_6347_46155# 2.63e-19
C26461 a_n1741_47186# a_11962_45724# 6.79e-20
C26462 a_n971_45724# a_8746_45002# 9.8e-20
C26463 a_3090_45724# a_11415_45002# 0.16525f
C26464 a_16388_46812# a_16751_46987# 0.005265f
C26465 a_n1925_46634# a_1431_46436# 3.57e-19
C26466 a_7715_46873# a_7920_46348# 0.080253f
C26467 a_4915_47217# a_6511_45714# 2.36e-21
C26468 a_5815_47464# a_6194_45824# 2.21e-20
C26469 a_4791_45118# a_6598_45938# 3.84e-19
C26470 a_6151_47436# a_5907_45546# 0.274247f
C26471 a_2063_45854# a_6428_45938# 3.74e-19
C26472 SMPL_ON_N a_20692_30879# 0.029397f
C26473 a_11453_44696# a_20205_31679# 1.75e-20
C26474 a_18479_47436# a_n357_42282# 0.003001f
C26475 a_10554_47026# a_3483_46348# 5.06e-20
C26476 a_7411_46660# a_8016_46348# 6.73e-19
C26477 a_n2293_46634# a_n1925_42282# 0.030317f
C26478 a_n1641_43230# a_n4318_38216# 6.62e-19
C26479 a_10922_42852# a_11136_42852# 0.097745f
C26480 a_12089_42308# a_12800_43218# 0.15794f
C26481 a_12379_42858# a_12991_43230# 3.82e-19
C26482 a_17730_32519# VDD 0.289738f
C26483 a_14209_32519# a_n784_42308# 0.004411f
C26484 a_n2157_42858# a_n4318_37592# 1.43e-19
C26485 a_22591_44484# RST_Z 5.01e-19
C26486 a_14205_43396# a_14456_42282# 1.85e-20
C26487 a_19237_31679# C10_N_btm 1.19e-19
C26488 a_743_42282# a_1755_42282# 0.058846f
C26489 a_3626_43646# a_7174_31319# 0.022247f
C26490 a_n4318_39304# a_n3690_39392# 8.45e-19
C26491 a_n1853_43023# a_n1736_42282# 0.004594f
C26492 a_20205_31679# a_17364_32525# 0.053947f
C26493 a_3090_45724# a_10533_42308# 5.9e-20
C26494 a_5343_44458# a_n2661_43922# 0.094786f
C26495 a_5518_44484# a_n2661_42834# 1.65e-20
C26496 a_1307_43914# a_1241_44260# 7.06e-19
C26497 a_10775_45002# a_10405_44172# 1.45e-20
C26498 a_21005_45260# a_20679_44626# 2.52e-20
C26499 a_21101_45002# a_20640_44752# 4.25e-19
C26500 a_11827_44484# a_20159_44458# 0.012941f
C26501 a_n2293_42834# a_1115_44172# 9.47e-21
C26502 a_11691_44458# a_18588_44850# 0.00186f
C26503 a_2711_45572# a_16547_43609# 4.49e-19
C26504 a_n357_42282# a_4190_30871# 0.035963f
C26505 a_3483_46348# a_14635_42282# 1.83e-20
C26506 a_7499_43078# a_10695_43548# 0.124597f
C26507 a_n746_45260# VDD 1.41433f
C26508 a_5883_43914# a_5708_44484# 2.58e-19
C26509 a_18587_45118# a_18579_44172# 8.05e-19
C26510 a_18184_42460# a_19279_43940# 0.132218f
C26511 a_n1605_47204# CLK_DATA 1.66e-20
C26512 a_n443_42852# a_16664_43396# 2.07e-20
C26513 a_n2017_45002# a_14021_43940# 1.77e-19
C26514 a_413_45260# a_15493_43940# 0.013529f
C26515 SMPL_ON_P DATA[0] 2.42e-19
C26516 a_n1741_47186# DATA[1] 0.021536f
C26517 a_12465_44636# a_6171_45002# 0.03098f
C26518 a_6165_46155# a_5066_45546# 0.041118f
C26519 a_n1151_42308# a_7639_45394# 0.004199f
C26520 a_n443_46116# a_2448_45028# 6.56e-19
C26521 a_3315_47570# a_413_45260# 7.08e-19
C26522 a_10227_46804# a_13159_45002# 1.01e-20
C26523 a_11599_46634# a_16019_45002# 8.13e-20
C26524 a_6755_46942# a_13904_45546# 2.1e-21
C26525 a_765_45546# a_n755_45592# 0.004312f
C26526 a_12741_44636# a_16375_45002# 0.042457f
C26527 a_4883_46098# a_5205_44484# 1.69e-20
C26528 a_n1613_43370# en_comp 1.09e-19
C26529 a_19321_45002# a_19610_45572# 7.05e-19
C26530 a_2063_45854# a_10903_45394# 1.39e-19
C26531 a_5068_46348# a_5527_46155# 6.64e-19
C26532 a_5164_46348# a_5210_46155# 0.006879f
C26533 a_14840_46494# a_10809_44734# 3.79e-21
C26534 a_15682_46116# a_6945_45028# 1.56e-19
C26535 a_18985_46122# a_19553_46090# 0.16939f
C26536 a_18819_46122# a_19335_46494# 0.108964f
C26537 a_4190_30871# CAL_N 0.045535f
C26538 a_1606_42308# a_6171_42473# 1.34e-20
C26539 a_1755_42282# a_5755_42308# 4.89e-19
C26540 a_1067_42314# a_6123_31319# 9e-21
C26541 a_564_42282# a_5934_30871# 2.52e-20
C26542 a_n913_45002# a_791_42968# 0.054288f
C26543 a_n1059_45260# a_1847_42826# 0.038913f
C26544 a_n2956_38680# a_n4334_40480# 4.16e-19
C26545 a_n2661_42834# a_9895_44260# 2.38e-19
C26546 a_n699_43396# a_104_43370# 0.21575f
C26547 a_n984_44318# a_453_43940# 3.53e-20
C26548 a_16241_44734# a_15682_43940# 2.85e-19
C26549 a_6755_46942# CLK 0.031541f
C26550 a_n755_45592# a_4921_42308# 0.001431f
C26551 a_n2810_45572# a_5934_30871# 1.88e-21
C26552 a_175_44278# a_1414_42308# 1.49e-20
C26553 a_4743_44484# a_n97_42460# 1.46e-20
C26554 a_n2956_39304# a_n4064_40160# 6.96e-19
C26555 a_18479_45785# a_19164_43230# 0.001979f
C26556 a_10227_46804# a_11967_42832# 0.461417f
C26557 a_n2661_45546# a_1260_45572# 7.47e-19
C26558 a_13059_46348# a_15415_45028# 2.08e-20
C26559 a_584_46384# a_2479_44172# 0.054912f
C26560 a_2063_45854# a_2127_44172# 5.29e-20
C26561 a_n2293_46098# en_comp 0.003369f
C26562 a_12465_44636# a_14673_44172# 0.101564f
C26563 a_16327_47482# a_20679_44626# 0.318301f
C26564 a_n743_46660# a_16112_44458# 0.001708f
C26565 a_n2497_47436# a_n1287_44306# 8.39e-19
C26566 a_12741_44636# a_413_45260# 0.009139f
C26567 a_3483_46348# a_2437_43646# 4.71e-20
C26568 a_10586_45546# a_11962_45724# 0.137051f
C26569 a_8049_45260# a_13904_45546# 0.003111f
C26570 a_n863_45724# a_n310_45572# 0.002342f
C26571 a_n755_45592# a_509_45822# 2.51e-20
C26572 a_n357_42282# a_n443_42852# 0.763015f
C26573 a_n2946_39866# a_n2860_39866# 0.011479f
C26574 a_n971_45724# a_6851_47204# 0.028789f
C26575 a_2905_45572# a_n1151_42308# 0.072935f
C26576 a_2063_45854# a_3815_47204# 5.54e-20
C26577 a_n237_47217# a_6545_47178# 0.021104f
C26578 a_n1741_47186# a_9863_47436# 0.006846f
C26579 a_1239_47204# a_n443_46116# 1.76e-21
C26580 a_n2833_47464# a_n1435_47204# 2.27e-20
C26581 a_2553_47502# a_3785_47178# 7.79e-20
C26582 a_n4064_39616# a_n2302_39866# 0.239588f
C26583 a_n4064_40160# a_n3565_39304# 0.028096f
C26584 a_5932_42308# VDAC_N 0.007314f
C26585 a_6123_31319# a_3726_37500# 0.002503f
C26586 a_n1630_35242# a_n83_35174# 7.97e-19
C26587 a_17749_42852# VDD 0.00742f
C26588 a_n4209_39590# a_n3607_39616# 0.002294f
C26589 a_n4334_39616# a_n4251_39616# 0.007692f
C26590 a_n4315_30879# a_n3420_39072# 0.036979f
C26591 a_14539_43914# a_17595_43084# 0.141972f
C26592 a_n2661_42834# a_n1379_43218# 1.92e-19
C26593 a_n356_44636# a_12379_42858# 8.61e-20
C26594 a_5111_44636# a_8325_42308# 6.44e-22
C26595 a_n913_45002# a_15051_42282# 0.003302f
C26596 a_n1059_45260# a_15486_42560# 2.84e-20
C26597 a_n2017_45002# a_15764_42576# 0.014981f
C26598 a_20205_31679# a_21589_35634# 3.35e-20
C26599 a_20692_30879# a_19864_35138# 1.26e-20
C26600 a_n2661_42282# a_6293_42852# 0.16527f
C26601 a_12379_46436# VDD 0.002681f
C26602 a_742_44458# a_945_42968# 4.68e-20
C26603 a_5891_43370# a_7871_42858# 0.051552f
C26604 a_8049_45260# CLK 0.033207f
C26605 a_n357_42282# a_375_42282# 0.142311f
C26606 a_12549_44172# a_19741_43940# 0.001206f
C26607 a_5907_45546# a_5111_44636# 0.01337f
C26608 a_5263_45724# a_4927_45028# 0.001784f
C26609 a_11415_45002# a_14815_43914# 0.070306f
C26610 a_15599_45572# a_18175_45572# 4.17e-21
C26611 a_15903_45785# a_16147_45260# 0.003162f
C26612 a_15765_45572# a_17786_45822# 1.13e-19
C26613 a_n1613_43370# a_n1699_43638# 0.160308f
C26614 a_12594_46348# a_12607_44458# 1.79e-19
C26615 a_2324_44458# a_8701_44490# 0.001089f
C26616 a_n863_45724# a_2232_45348# 0.002794f
C26617 a_8049_45260# a_17023_45118# 1.03e-20
C26618 a_3483_46348# a_4181_44734# 6.14e-20
C26619 a_1823_45246# a_5891_43370# 5.34e-19
C26620 a_3260_45572# a_413_45260# 4.87e-19
C26621 a_17339_46660# a_11967_42832# 0.493072f
C26622 a_16333_45814# a_16377_45572# 3.69e-19
C26623 a_16115_45572# a_16211_45572# 0.013793f
C26624 a_12741_44636# a_13468_44734# 9.06e-19
C26625 a_2711_45572# a_6171_45002# 0.457554f
C26626 a_10903_43370# a_13076_44458# 5.54e-19
C26627 a_n1435_47204# a_6969_46634# 4e-20
C26628 a_13717_47436# a_6755_46942# 9.51e-20
C26629 a_n4209_37414# C6_P_btm 1.26e-20
C26630 a_n3565_37414# C8_P_btm 1.71e-20
C26631 a_11599_46634# a_10428_46928# 0.001591f
C26632 a_7754_39964# RST_Z 0.843939f
C26633 a_4338_37500# a_n923_35174# 1.22e-19
C26634 VDAC_Pi VDD 0.591846f
C26635 a_n3565_38216# VREF_GND 0.001975f
C26636 a_4883_46098# a_5385_46902# 6e-21
C26637 CAL_N a_22705_38406# 4.85e-21
C26638 a_22521_40055# a_22780_39857# 3.15e-19
C26639 a_22521_40599# a_22609_38406# 0.032572f
C26640 a_22469_40625# CAL_P 0.001716f
C26641 a_22459_39145# a_22469_39537# 0.351623f
C26642 a_22521_39511# a_22545_38993# 0.27533f
C26643 a_6545_47178# a_8270_45546# 4.75e-21
C26644 a_4915_47217# a_10768_47026# 4.45e-19
C26645 a_6151_47436# a_10384_47026# 2.82e-20
C26646 a_n1151_42308# a_12816_46660# 0.008712f
C26647 a_n881_46662# a_491_47026# 3.56e-21
C26648 a_768_44030# a_n2438_43548# 6.89e-19
C26649 a_14021_43940# a_19164_43230# 1.26e-20
C26650 a_9313_44734# a_15959_42545# 6.1e-20
C26651 a_n4318_40392# a_n3420_39072# 7.42e-22
C26652 a_n1761_44111# a_n4318_37592# 1.64e-20
C26653 a_9145_43396# a_13837_43396# 4.66e-20
C26654 a_3080_42308# a_14209_32519# 0.001913f
C26655 a_2982_43646# a_13467_32519# 0.006898f
C26656 a_n356_44636# a_18727_42674# 2.05e-20
C26657 a_n1899_43946# a_n1736_42282# 5.43e-21
C26658 a_n2109_45247# VDD 0.266396f
C26659 a_n97_42460# a_n1736_43218# 7.3e-22
C26660 a_n2012_43396# a_n3674_39304# 8.64e-20
C26661 a_3357_43084# EN_OFFSET_CAL 6.03e-21
C26662 a_10341_43396# a_12281_43396# 0.012652f
C26663 a_14579_43548# a_14621_43646# 8.44e-19
C26664 a_14358_43442# a_14537_43646# 0.010303f
C26665 a_n2293_46634# a_8387_43230# 4.77e-21
C26666 a_13661_43548# a_13635_43156# 0.004897f
C26667 a_2711_45572# a_14673_44172# 0.04263f
C26668 a_18953_45572# a_11691_44458# 2.11e-20
C26669 a_12549_44172# a_17333_42852# 9.44e-21
C26670 a_n971_45724# a_n327_42558# 0.01976f
C26671 a_3090_45724# a_9885_43646# 0.003881f
C26672 a_14180_45002# a_14537_43396# 0.143922f
C26673 a_3065_45002# a_5009_45028# 6.35e-21
C26674 a_20623_45572# a_11827_44484# 1.21e-20
C26675 a_21363_45546# a_21359_45002# 0.01738f
C26676 a_20731_45938# a_20567_45036# 1.28e-19
C26677 a_21188_45572# a_21101_45002# 3.83e-19
C26678 a_n2810_45028# a_n2661_43370# 0.002593f
C26679 a_20205_31679# a_19237_31679# 0.051574f
C26680 a_8746_45002# a_9313_44734# 2.85e-19
C26681 a_8953_45002# a_1423_45028# 0.011739f
C26682 a_9482_43914# a_15595_45028# 0.0011f
C26683 a_13556_45296# a_15415_45028# 1.78e-20
C26684 a_14976_45028# a_14955_43396# 6.28e-20
C26685 a_12861_44030# a_15785_43172# 4.72e-19
C26686 a_12891_46348# a_10903_43370# 0.132903f
C26687 a_n935_46688# a_n2293_46098# 2.46e-19
C26688 a_5807_45002# a_8349_46414# 2.69e-20
C26689 a_6755_46942# a_14035_46660# 0.040006f
C26690 a_12816_46660# a_14084_46812# 6.32e-20
C26691 a_n2497_47436# a_n452_45724# 5.75e-21
C26692 a_n1925_46634# a_2202_46116# 0.00159f
C26693 a_n743_46660# a_1138_42852# 0.056829f
C26694 a_n2438_43548# a_1176_45822# 0.073092f
C26695 a_n2661_46634# a_3483_46348# 0.051915f
C26696 a_n2293_46634# a_2698_46116# 3.76e-20
C26697 a_13717_47436# a_8049_45260# 5.14e-20
C26698 a_n881_46662# a_14840_46494# 4.54e-19
C26699 a_n1613_43370# a_2324_44458# 0.027159f
C26700 SMPL_ON_P a_n2472_45546# 3.24e-19
C26701 a_601_46902# a_376_46348# 8.72e-19
C26702 a_33_46660# a_472_46348# 0.003485f
C26703 a_n310_44484# VDD 7.01e-20
C26704 a_18525_43370# a_18504_43218# 6.38e-19
C26705 a_16137_43396# a_17749_42852# 0.001147f
C26706 a_9313_44734# RST_Z 0.002698f
C26707 a_n97_42460# a_11633_42558# 0.011546f
C26708 a_10341_42308# a_12089_42308# 0.003265f
C26709 a_n13_43084# a_133_42852# 0.171361f
C26710 a_3626_43646# a_5932_42308# 0.062334f
C26711 a_3080_42308# a_4169_42308# 0.001081f
C26712 a_3483_46348# a_14543_43071# 5.23e-21
C26713 a_4185_45028# a_13635_43156# 7.46e-20
C26714 a_11691_44458# a_18443_44721# 0.042634f
C26715 a_n2312_39304# a_n4209_39304# 0.19527f
C26716 a_9290_44172# a_7871_42858# 2.35e-19
C26717 a_n443_42852# a_n144_43396# 5.19e-20
C26718 a_n2661_44458# a_10334_44484# 0.009408f
C26719 a_1307_43914# a_11967_42832# 0.031135f
C26720 a_327_44734# a_644_44056# 1.79e-19
C26721 a_n2017_45002# a_5013_44260# 1.47e-20
C26722 a_8953_45546# a_9127_43156# 0.00897f
C26723 a_n1925_42282# a_743_42282# 0.052333f
C26724 a_n1059_45260# a_5244_44056# 4.98e-21
C26725 a_n913_45002# a_3905_42865# 5e-19
C26726 a_949_44458# a_n699_43396# 1.66e-19
C26727 a_13249_42308# a_13565_43940# 0.048533f
C26728 a_10227_46804# a_20273_45572# 4.14e-20
C26729 a_11415_45002# a_20075_46420# 2.53e-20
C26730 a_3483_46348# a_8199_44636# 1.81719f
C26731 a_3090_45724# a_13259_45724# 0.261789f
C26732 a_19636_46660# a_10809_44734# 3.84e-19
C26733 a_13487_47204# a_2437_43646# 0.014506f
C26734 a_4955_46873# a_2711_45572# 2.02e-20
C26735 a_2107_46812# a_9049_44484# 0.240008f
C26736 a_n971_45724# a_3232_43370# 0.058382f
C26737 a_14035_46660# a_8049_45260# 0.002246f
C26738 a_3160_47472# a_413_45260# 0.208121f
C26739 a_n1151_42308# a_n37_45144# 4.16e-19
C26740 a_n881_46662# a_16115_45572# 0.033547f
C26741 a_4883_46098# a_19431_45546# 5.31e-20
C26742 a_16327_47482# a_20528_45572# 0.011969f
C26743 a_n743_46660# a_11962_45724# 1.66e-20
C26744 a_3877_44458# a_5263_45724# 3.55e-21
C26745 a_11453_44696# a_16147_45260# 0.026325f
C26746 a_n1435_47204# a_3357_43084# 1.08491f
C26747 a_2063_45854# a_2382_45260# 5.84e-19
C26748 a_12549_44172# a_11778_45572# 1.09e-19
C26749 a_n2293_46098# a_2324_44458# 0.018455f
C26750 a_5164_46348# a_5497_46414# 0.203417f
C26751 a_12741_44636# a_18985_46122# 1.17e-19
C26752 a_n3674_39304# a_n4064_39616# 0.020873f
C26753 a_17538_32519# VDD 0.352239f
C26754 a_20974_43370# RST_Z 0.001986f
C26755 a_526_44458# a_6171_42473# 4.56e-20
C26756 a_n357_42282# a_14635_42282# 0.010701f
C26757 a_9290_44172# a_11897_42308# 7.06e-19
C26758 a_n2293_42834# a_n2012_43396# 0.001738f
C26759 a_1307_43914# a_648_43396# 6.76e-20
C26760 a_22612_30879# VCM 0.473529f
C26761 a_11967_42832# a_18579_44172# 0.158329f
C26762 a_10193_42453# a_19339_43156# 0.003128f
C26763 a_5111_44636# a_9145_43396# 0.057312f
C26764 a_n2438_43548# DATA[0] 5.04e-19
C26765 a_n743_46660# DATA[1] 1.69e-21
C26766 a_383_46660# VDD 0.198466f
C26767 a_n1925_46634# DATA[3] 4.06e-21
C26768 a_13720_44458# a_13483_43940# 0.001108f
C26769 a_n2661_43922# a_453_43940# 0.006118f
C26770 a_3363_44484# a_3600_43914# 4.63e-19
C26771 a_n2661_42834# a_2127_44172# 0.019594f
C26772 a_13249_42308# a_5534_30871# 0.215947f
C26773 a_20640_44752# a_20766_44850# 0.17072f
C26774 a_20362_44736# a_19279_43940# 0.039759f
C26775 a_20679_44626# a_20835_44721# 0.105995f
C26776 a_n2661_43370# a_n2129_43609# 3.94e-19
C26777 a_12005_46116# a_10490_45724# 6.17e-19
C26778 a_19321_45002# a_21101_45002# 0.005955f
C26779 a_7832_46660# a_7229_43940# 7.4e-21
C26780 a_13747_46662# a_11827_44484# 0.044822f
C26781 a_14513_46634# a_2437_43646# 2.95e-20
C26782 a_18597_46090# a_18248_44752# 8.18e-21
C26783 a_10903_43370# a_11322_45546# 0.313957f
C26784 a_11387_46155# a_11525_45546# 4.09e-19
C26785 a_12465_44636# a_12607_44458# 0.186652f
C26786 a_11453_44696# a_10334_44484# 0.001021f
C26787 a_6945_45028# a_6598_45938# 0.005236f
C26788 a_6755_46942# a_10951_45334# 8.67e-21
C26789 a_5257_43370# a_1307_43914# 0.020655f
C26790 a_11189_46129# a_11962_45724# 1.89e-19
C26791 a_13351_46090# a_10193_42453# 3.16e-21
C26792 a_13259_45724# a_15002_46116# 4.39e-20
C26793 a_13885_46660# a_3357_43084# 2.28e-20
C26794 a_n1613_43370# a_n1699_44726# 0.166123f
C26795 a_13607_46688# a_413_45260# 1.59e-20
C26796 a_6123_31319# a_1239_39043# 6.84e-20
C26797 a_5534_30871# VIN_P 0.00357f
C26798 a_17303_42282# a_18214_42558# 7.99e-21
C26799 a_4958_30871# a_18220_42308# 6.64e-20
C26800 a_19339_43156# VDD 0.338297f
C26801 a_18599_43230# RST_Z 8.97e-22
C26802 a_n2293_42834# a_n914_42852# 1.34e-19
C26803 en_comp a_n1736_42282# 6.61e-20
C26804 a_n967_45348# a_n3674_38216# 3.49e-20
C26805 a_n2810_45028# COMP_P 1.61e-21
C26806 a_13351_46090# VDD 0.238036f
C26807 a_18989_43940# a_19177_43646# 1.57e-19
C26808 a_18443_44721# a_4190_30871# 3.98e-20
C26809 a_11341_43940# a_22959_43948# 4.69e-19
C26810 a_22223_43948# a_15493_43940# 0.051823f
C26811 a_n2293_43922# a_12281_43396# 0.147288f
C26812 a_n913_45002# a_n961_42308# 9.71e-19
C26813 a_n1059_45260# a_n473_42460# 8.15e-19
C26814 a_n2017_45002# a_196_42282# 0.010023f
C26815 a_14955_43940# a_15301_44260# 0.013377f
C26816 a_6756_44260# a_6671_43940# 1.48e-19
C26817 a_1414_42308# a_n97_42460# 0.196768f
C26818 a_9313_44734# a_16243_43396# 1.87e-19
C26819 a_n699_43396# a_n1076_43230# 0.001631f
C26820 a_15433_44458# a_14955_43396# 1.98e-19
C26821 a_18079_43940# a_14021_43940# 4.92e-20
C26822 a_n2956_38216# a_n2216_37984# 8.63e-19
C26823 a_n2956_37592# a_n4318_37592# 0.023082f
C26824 a_8049_45260# a_10951_45334# 1.03e-20
C26825 a_n1925_42282# a_626_44172# 4.51e-21
C26826 a_2324_44458# a_8704_45028# 9.12e-20
C26827 a_11525_45546# a_11778_45572# 0.011913f
C26828 a_4185_45028# a_22223_45036# 0.002889f
C26829 a_3090_45724# a_n2661_43922# 0.044809f
C26830 a_12861_44030# a_13565_43940# 1.02e-19
C26831 a_584_46384# a_n229_43646# 3.24e-19
C26832 a_17339_46660# a_18989_43940# 0.002356f
C26833 a_6755_46942# a_17061_44484# 9.81e-19
C26834 a_n357_42282# a_2437_43646# 1.4e-19
C26835 a_11652_45724# a_11688_45572# 0.001673f
C26836 a_12549_44172# a_13483_43940# 0.007788f
C26837 a_768_44030# a_12429_44172# 0.007216f
C26838 a_n2661_45546# a_n2840_45002# 0.002083f
C26839 a_9863_47436# a_n743_46660# 1.91e-20
C26840 a_4883_46098# a_12891_46348# 0.085714f
C26841 a_16327_47482# a_19594_46812# 0.004271f
C26842 a_5815_47464# a_2107_46812# 8.74e-21
C26843 a_n3565_39304# C10_P_btm 2.44e-19
C26844 a_3754_38802# a_3754_38470# 0.02792f
C26845 a_n4209_39304# C8_P_btm 9.97e-19
C26846 a_13507_46334# a_768_44030# 0.019457f
C26847 a_10227_46804# a_5807_45002# 0.262866f
C26848 a_15673_47210# a_16750_47204# 1.46e-19
C26849 a_n237_47217# a_3877_44458# 0.059355f
C26850 a_n971_45724# a_4651_46660# 7.48e-19
C26851 a_2952_47436# a_2959_46660# 5.17e-19
C26852 a_3160_47472# a_2609_46660# 0.018687f
C26853 a_n1151_42308# a_2443_46660# 3.77e-19
C26854 a_2905_45572# a_3177_46902# 0.014554f
C26855 a_584_46384# a_2864_46660# 2.26e-19
C26856 a_n4064_37984# VDAC_P 2.99e-19
C26857 a_n1741_47186# a_5907_46634# 8.63e-20
C26858 a_n443_46116# a_491_47026# 1.47e-19
C26859 a_22465_38105# VDD 1.3089f
C26860 a_6197_43396# a_7287_43370# 0.041762f
C26861 a_n97_42460# a_12281_43396# 6.17e-19
C26862 a_3626_43646# a_4181_43396# 2.16e-20
C26863 a_n2661_42834# a_n4318_38216# 0.023647f
C26864 a_18494_42460# a_18907_42674# 0.11494f
C26865 a_18184_42460# a_19332_42282# 0.042769f
C26866 a_9028_43914# a_9127_43156# 9.19e-20
C26867 a_n356_44636# a_3823_42558# 1.46e-19
C26868 a_n2293_43922# a_n3674_38680# 2.31e-20
C26869 a_n2810_45028# a_n3565_37414# 0.135518f
C26870 a_5883_43914# a_9223_42460# 2.74e-20
C26871 a_14021_43940# a_14209_32519# 0.042544f
C26872 a_6765_43638# a_6547_43396# 0.209641f
C26873 a_6293_42852# a_7112_43396# 5.47e-21
C26874 a_3539_42460# a_3457_43396# 2.02e-20
C26875 a_6031_43396# a_8147_43396# 3.33e-21
C26876 a_20820_30879# a_15493_43940# 1.28e-20
C26877 a_19692_46634# a_21845_43940# 0.014352f
C26878 a_13259_45724# a_14815_43914# 0.001261f
C26879 a_n1059_45260# a_5111_44636# 0.038143f
C26880 a_10227_46804# a_10518_42984# 0.225803f
C26881 a_n2293_46634# a_15743_43084# 8.65e-20
C26882 a_6511_45714# a_5883_43914# 1.33e-21
C26883 a_2711_45572# a_12607_44458# 8.18e-21
C26884 a_13249_42308# a_11691_44458# 0.017891f
C26885 a_2324_44458# a_2675_43914# 7.61e-20
C26886 a_n1613_43370# a_n2157_42858# 0.303592f
C26887 a_7227_45028# a_6298_44484# 0.003074f
C26888 a_9049_44484# a_n2661_44458# 0.015549f
C26889 a_12549_44172# a_13678_32519# 0.004825f
C26890 a_5807_45002# a_17339_46660# 0.02927f
C26891 a_16131_47204# a_765_45546# 0.005958f
C26892 a_n2312_39304# a_n2157_46122# 0.00402f
C26893 a_8145_46902# a_8492_46660# 0.051162f
C26894 a_1799_45572# a_3090_45724# 1.03e-19
C26895 a_n1435_47204# a_9625_46129# 2.1e-20
C26896 a_4791_45118# a_2324_44458# 0.19212f
C26897 a_6151_47436# a_13925_46122# 5.38e-19
C26898 a_n2433_43396# a_n1329_42308# 3.94e-21
C26899 a_n2129_43609# COMP_P 2.54e-20
C26900 a_15682_43940# a_15890_42674# 1.13e-19
C26901 a_16137_43396# a_19339_43156# 2.87e-19
C26902 a_17324_43396# a_17595_43084# 6.75e-20
C26903 a_17499_43370# a_17701_42308# 8.78e-19
C26904 a_743_42282# a_8387_43230# 6e-20
C26905 a_n1076_43230# a_n4318_38680# 1.6e-20
C26906 a_n1699_43638# a_n1736_42282# 7.33e-20
C26907 a_19721_31679# VDD 0.521328f
C26908 a_n2157_42858# a_n1533_42852# 9.73e-19
C26909 a_n1641_43230# a_n1545_43230# 0.013793f
C26910 a_n1423_42826# a_n1379_43218# 3.69e-19
C26911 a_n1991_42858# a_n967_43230# 2.36e-20
C26912 a_n1853_43023# a_n722_43218# 0.001894f
C26913 a_15743_43084# a_5342_30871# 0.006894f
C26914 a_18114_32519# RST_Z 0.049686f
C26915 a_3232_43370# a_9313_44734# 0.11426f
C26916 a_18911_45144# a_11827_44484# 4.77e-20
C26917 a_16922_45042# a_16237_45028# 3.82e-19
C26918 a_18184_42460# a_21101_45002# 2.52e-36
C26919 a_19778_44110# a_21359_45002# 6.57e-19
C26920 a_18494_42460# a_21005_45260# 1.23e-20
C26921 a_526_44458# a_3457_43396# 0.002177f
C26922 a_2274_45254# a_n2661_43922# 5.45e-20
C26923 a_2382_45260# a_n2661_42834# 0.055134f
C26924 a_21363_45546# a_19279_43940# 1.63e-19
C26925 a_n2661_43370# a_n2129_44697# 0.014856f
C26926 a_n2293_42834# a_2779_44458# 7.79e-21
C26927 a_17613_45144# a_11691_44458# 5.83e-21
C26928 a_10227_46804# a_16197_42308# 0.001903f
C26929 a_10193_42453# a_17973_43940# 0.084505f
C26930 a_11823_42460# a_10949_43914# 0.002042f
C26931 a_3537_45260# a_5708_44484# 3.43e-20
C26932 a_765_45546# a_3483_46348# 1.15e-19
C26933 a_22591_46660# a_22959_46660# 7.52e-19
C26934 a_n2293_46634# a_380_45546# 6.42e-19
C26935 a_n2438_43548# a_n2472_45546# 0.008798f
C26936 a_n133_46660# a_n2661_45546# 1.33e-20
C26937 a_n881_46662# a_6511_45714# 0.149116f
C26938 a_11415_45002# a_21076_30879# 8.27e-21
C26939 a_20202_43084# a_21297_46660# 4.61e-21
C26940 a_n1613_43370# a_6667_45809# 0.007328f
C26941 a_4883_46098# a_11322_45546# 9.36e-20
C26942 a_7715_46873# a_8062_46482# 9.21e-19
C26943 a_20820_30879# a_12741_44636# 0.103478f
C26944 a_n2661_46634# a_n357_42282# 3.78e-20
C26945 a_n1925_46634# a_n1079_45724# 4.37e-19
C26946 a_n1021_46688# a_n2293_45546# 2.36e-21
C26947 a_11735_46660# a_6945_45028# 1.07e-19
C26948 a_3090_45724# a_18189_46348# 0.029136f
C26949 a_10227_46804# a_15143_45578# 0.010124f
C26950 a_17973_43940# VDD 0.265874f
C26951 a_16823_43084# a_17303_42282# 3.24e-21
C26952 a_3080_42308# VDAC_Pi 3.65e-19
C26953 a_19700_43370# a_19647_42308# 4.12e-19
C26954 a_4361_42308# a_11633_42308# 9.01e-19
C26955 a_12800_43218# a_12991_43230# 4.61e-19
C26956 a_n2293_42282# a_n4318_38216# 0.004948f
C26957 a_5342_30871# a_1606_42308# 0.023615f
C26958 a_743_42282# a_16522_42674# 0.003239f
C26959 a_15743_43084# a_20107_42308# 1.94e-20
C26960 a_7227_42852# a_6761_42308# 4.22e-19
C26961 a_18989_43940# a_18579_44172# 0.035827f
C26962 a_18443_44721# a_18753_44484# 0.013793f
C26963 a_18374_44850# a_18681_44484# 3.69e-19
C26964 a_949_44458# a_1467_44172# 0.004991f
C26965 a_n2661_44458# a_3905_42865# 2.18e-19
C26966 a_742_44458# a_1414_42308# 0.052151f
C26967 a_21588_30879# a_22521_40055# 3.72e-20
C26968 a_22223_47212# VDD 0.236555f
C26969 a_12465_44636# RST_Z 0.002855f
C26970 a_n699_43396# a_175_44278# 0.001042f
C26971 a_n1059_45260# a_4235_43370# 0.003711f
C26972 a_n2017_45002# a_4699_43561# 1.2e-20
C26973 a_n913_45002# a_4093_43548# 4.03e-21
C26974 a_n357_42282# a_14543_43071# 0.004653f
C26975 a_1307_43914# a_5745_43940# 0.001752f
C26976 a_n443_42852# a_8952_43230# 7.98e-19
C26977 a_3357_43084# a_3539_42460# 0.001767f
C26978 a_4883_46098# SINGLE_ENDED 0.1664f
C26979 a_3090_45724# a_17478_45572# 0.128299f
C26980 a_15227_44166# a_15765_45572# 2.32e-20
C26981 a_14976_45028# a_15861_45028# 1.41e-19
C26982 a_12861_44030# a_11691_44458# 0.196929f
C26983 a_18597_46090# a_16922_45042# 0.028931f
C26984 a_16327_47482# a_18494_42460# 0.083754f
C26985 a_5066_45546# a_5210_46155# 0.001301f
C26986 a_n2661_46634# a_11963_45334# 0.036874f
C26987 a_n743_46660# a_7229_43940# 6.59e-21
C26988 a_n971_45724# a_8975_43940# 7.38e-21
C26989 a_n2312_40392# a_n2661_43370# 1.34e-19
C26990 a_11599_46634# a_11827_44484# 1.7e-22
C26991 a_18819_46122# a_19240_46482# 0.089677f
C26992 a_18985_46122# a_16375_45002# 9.94e-20
C26993 a_8199_44636# a_n357_42282# 0.023438f
C26994 a_167_45260# a_2307_45899# 0.005265f
C26995 a_17715_44484# a_18051_46116# 9.64e-19
C26996 a_n1925_46634# a_7705_45326# 9.07e-21
C26997 a_n2293_46098# a_6667_45809# 1.01e-20
C26998 a_2609_46660# a_413_45260# 0.022446f
C26999 a_15368_46634# a_8696_44636# 2.65e-20
C27000 a_13747_46662# a_15595_45028# 3.1e-20
C27001 a_5807_45002# a_1307_43914# 0.007287f
C27002 a_n2293_46634# a_10775_45002# 1.79e-21
C27003 a_13661_43548# a_16019_45002# 0.001206f
C27004 a_768_44030# a_2903_45348# 0.001561f
C27005 a_2107_46812# a_5147_45002# 4.3e-20
C27006 a_13507_46334# a_13490_45067# 6.13e-20
C27007 a_13887_32519# RST_Z 0.048332f
C27008 a_4190_30871# VIN_P 0.049977f
C27009 a_11323_42473# a_5742_30871# 0.198522f
C27010 COMP_P a_n2302_40160# 4e-20
C27011 a_n3674_38680# a_n3420_39616# 0.020072f
C27012 a_10533_42308# a_11633_42558# 9.27e-21
C27013 a_17364_32525# C9_N_btm 7.29e-20
C27014 a_22591_43396# VDD 0.280354f
C27015 a_5534_30871# a_11206_38545# 2.6e-20
C27016 a_20731_47026# VDD 0.132317f
C27017 a_21188_46660# SINGLE_ENDED 4.66e-21
C27018 a_n2661_43370# a_n2840_42826# 3.35e-19
C27019 a_n2293_42834# a_n13_43084# 0.007462f
C27020 a_1307_43914# a_10518_42984# 3.51e-21
C27021 a_10157_44484# a_9803_43646# 0.001011f
C27022 a_10334_44484# a_9145_43396# 1.97e-20
C27023 a_n357_42282# a_19511_42282# 0.056757f
C27024 a_17730_32519# a_14021_43940# 9.75e-19
C27025 a_n2661_42834# a_n1655_43396# 2.44e-19
C27026 a_7499_43078# a_8685_42308# 7.11e-19
C27027 a_n863_45724# a_7174_31319# 4.84e-21
C27028 a_2382_45260# a_n2293_42282# 0.080755f
C27029 a_16922_45042# a_743_42282# 0.120316f
C27030 a_1423_45028# a_8037_42858# 1.11e-21
C27031 a_167_45260# a_1423_45028# 0.123079f
C27032 a_1823_45246# a_2304_45348# 4.41e-19
C27033 a_12005_46116# a_6171_45002# 1.39e-20
C27034 a_n1613_43370# a_n1761_44111# 0.148121f
C27035 a_2711_45572# a_8746_45002# 0.010166f
C27036 a_6511_45714# a_8162_45546# 0.004311f
C27037 a_6598_45938# a_6812_45938# 0.097745f
C27038 a_6667_45809# a_7230_45938# 0.049827f
C27039 a_6472_45840# a_8568_45546# 3.47e-20
C27040 a_18985_46122# a_413_45260# 1.46e-21
C27041 a_19321_45002# a_20766_44850# 0.004119f
C27042 a_9569_46155# a_8953_45002# 0.002046f
C27043 a_5807_45002# a_18579_44172# 0.003978f
C27044 a_8049_45260# a_19418_45938# 1.68e-19
C27045 a_n443_42852# a_13249_42308# 0.033352f
C27046 a_8199_44636# a_11963_45334# 8.83e-21
C27047 a_2324_44458# a_3429_45260# 2.54e-20
C27048 a_13259_45724# a_13297_45572# 0.003457f
C27049 a_17339_46660# a_18315_45260# 0.009833f
C27050 a_526_44458# a_3357_43084# 0.04478f
C27051 a_n237_47217# a_8128_46384# 0.113499f
C27052 a_1209_47178# a_n881_46662# 4.08e-21
C27053 a_1239_47204# a_n1613_43370# 0.001663f
C27054 a_3785_47178# a_2747_46873# 4.9e-20
C27055 a_n1151_42308# a_7_47243# 1.92e-19
C27056 a_n4315_30879# a_n2946_37690# 1.33e-19
C27057 a_14311_47204# a_10227_46804# 2.11e-19
C27058 a_15673_47210# a_16327_47482# 0.206019f
C27059 a_15811_47375# a_16023_47582# 0.003622f
C27060 a_7903_47542# a_4883_46098# 3.03e-21
C27061 a_13717_47436# a_18780_47178# 1.64e-19
C27062 a_12861_44030# a_18479_47436# 0.065796f
C27063 a_7174_31319# a_6886_37412# 4.9e-19
C27064 a_15507_47210# a_16763_47508# 0.043475f
C27065 a_5742_30871# C0_P_btm 0.014563f
C27066 a_1177_38525# a_2684_37794# 3.29e-20
C27067 a_n4334_38528# a_n4064_37984# 7.91e-19
C27068 a_n3690_38528# a_n3420_37984# 8.87e-19
C27069 a_n2946_38778# a_n3565_38216# 0.001251f
C27070 a_n2302_38778# a_n4209_38216# 0.001254f
C27071 a_n4209_38502# a_n2302_37984# 0.001417f
C27072 a_n4064_38528# a_n4334_38304# 0.001145f
C27073 a_n3420_38528# a_n3690_38304# 0.018295f
C27074 a_n3565_38502# a_n2946_37984# 0.001251f
C27075 a_n4064_40160# a_n3690_37440# 2.54e-19
C27076 a_11599_46634# a_16588_47582# 2.07e-20
C27077 a_19511_42282# CAL_N 0.001217f
C27078 a_2711_45572# RST_Z 4.2e-20
C27079 a_13565_44260# a_9145_43396# 2.31e-20
C27080 a_14539_43914# a_18695_43230# 1.08e-19
C27081 a_7499_43940# a_7112_43396# 0.001375f
C27082 a_11341_43940# a_12293_43646# 8.32e-19
C27083 a_15682_43940# a_16547_43609# 0.008948f
C27084 a_15301_44260# a_8685_43396# 1.7e-20
C27085 a_11967_42832# a_13635_43156# 0.053949f
C27086 a_15493_43396# a_15681_43442# 0.029338f
C27087 a_n2810_45028# a_n4209_39304# 0.021684f
C27088 a_3175_45822# VDD 0.193907f
C27089 a_12861_44030# a_4190_30871# 6.78e-20
C27090 a_3090_45724# a_20935_43940# 1.49e-20
C27091 a_20107_45572# a_21513_45002# 8.78e-20
C27092 a_20841_45814# a_20719_45572# 3.16e-19
C27093 a_10907_45822# a_9482_43914# 3.21e-20
C27094 a_8049_45260# a_18248_44752# 6.37e-21
C27095 a_n2293_46634# a_3539_42460# 0.003606f
C27096 a_18597_46090# a_15743_43084# 0.023066f
C27097 a_16147_45260# a_n1059_45260# 5.91e-21
C27098 a_6472_45840# a_n2661_43370# 5.95e-20
C27099 a_7227_45028# a_7418_45067# 4e-19
C27100 a_12891_46348# a_8685_43396# 3.82e-20
C27101 a_n1151_42308# a_n1076_43230# 0.00783f
C27102 C0_P_btm C0_dummy_P_btm 7.61701f
C27103 C3_P_btm C1_N_btm 5.97e-19
C27104 C1_P_btm C0_dummy_N_btm 2.22e-19
C27105 C5_P_btm C3_N_btm 2.12e-19
C27106 a_15811_47375# a_16751_46987# 1.26e-19
C27107 a_n2497_47436# a_167_45260# 0.001788f
C27108 a_13487_47204# a_765_45546# 0.006318f
C27109 a_16327_47482# a_16388_46812# 0.01513f
C27110 a_2107_46812# a_3055_46660# 0.001203f
C27111 a_18194_35068# VDD 2.17116f
C27112 a_n2109_47186# a_1823_45246# 7.36e-20
C27113 a_1239_47204# a_n2293_46098# 5.76e-21
C27114 a_8128_46384# a_8270_45546# 0.002121f
C27115 a_11453_44696# a_19333_46634# 0.026664f
C27116 a_12861_44030# a_17829_46910# 0.058114f
C27117 a_13717_47436# a_18285_46348# 1.31e-20
C27118 a_n1741_47186# a_1176_45822# 1.11e-19
C27119 a_n971_45724# a_n1076_46494# 8.23e-19
C27120 a_n746_45260# a_n901_46420# 8.55e-20
C27121 a_5807_45002# a_10467_46802# 0.007388f
C27122 a_n1925_46634# a_6540_46812# 0.008209f
C27123 a_2443_46660# a_3177_46902# 0.053479f
C27124 a_104_43370# a_133_42852# 8.41e-20
C27125 a_n2661_42282# a_2713_42308# 1.2e-19
C27126 a_15743_43084# a_743_42282# 0.029529f
C27127 a_19700_43370# a_4190_30871# 0.046581f
C27128 a_2982_43646# a_16795_42852# 1.51e-20
C27129 a_7542_44172# a_6123_31319# 8.34e-21
C27130 a_17499_43370# a_4361_42308# 6.03e-20
C27131 a_3626_43646# a_15567_42826# 2.41e-20
C27132 a_19692_46634# a_14209_32519# 9.21e-20
C27133 a_1823_45246# a_5837_43396# 3.58e-21
C27134 a_n2956_39304# a_n4318_39304# 0.023717f
C27135 a_5147_45002# a_n2661_44458# 0.024256f
C27136 a_13661_43548# a_13814_43218# 4.89e-20
C27137 a_11787_45002# a_11691_44458# 1.53e-19
C27138 a_45_45144# a_n2661_43370# 4.17e-19
C27139 a_n2312_40392# COMP_P 0.035637f
C27140 a_n2312_39304# a_n4318_37592# 0.023445f
C27141 a_4185_45028# a_8791_43396# 4.43e-22
C27142 a_16751_45260# a_17719_45144# 3.82e-19
C27143 a_13348_45260# a_11827_44484# 3.7e-22
C27144 a_5263_45724# a_5244_44056# 5.95e-21
C27145 a_8696_44636# a_15146_44811# 1.39e-19
C27146 a_327_44734# a_949_44458# 0.003334f
C27147 a_413_45260# a_2779_44458# 0.024142f
C27148 a_1667_45002# a_742_44458# 0.002122f
C27149 a_n743_46660# a_739_46482# 0.005906f
C27150 a_5807_45002# a_8034_45724# 1.95e-20
C27151 a_14513_46634# a_765_45546# 5.52e-20
C27152 a_16388_46812# a_16434_46987# 0.006879f
C27153 a_n1925_46634# a_1337_46436# 3.83e-19
C27154 a_4915_47217# a_6472_45840# 6.14e-21
C27155 a_4791_45118# a_6667_45809# 0.005119f
C27156 a_6151_47436# a_5263_45724# 3e-19
C27157 a_12861_44030# a_n443_42852# 0.015171f
C27158 SMPL_ON_N a_20205_31679# 0.029367f
C27159 a_15227_44166# a_18280_46660# 0.007923f
C27160 a_18834_46812# a_18900_46660# 0.006978f
C27161 a_10623_46897# a_3483_46348# 6.27e-20
C27162 a_6851_47204# a_2711_45572# 3.11e-21
C27163 a_5894_47026# a_5937_45572# 5.36e-21
C27164 a_7411_46660# a_7920_46348# 0.004089f
C27165 a_768_44030# a_10586_45546# 3.88e-20
C27166 a_n2442_46660# a_n1925_42282# 8.58e-20
C27167 a_n2293_46634# a_526_44458# 0.579444f
C27168 a_n1423_42826# a_n4318_38216# 3.57e-19
C27169 a_12379_42858# a_12800_43218# 0.089677f
C27170 a_n1991_42858# a_n2104_42282# 2.18e-19
C27171 a_10991_42826# a_11136_42852# 0.057222f
C27172 a_22591_44484# VDD 0.223346f
C27173 a_n2472_42826# a_n4318_37592# 2.65e-20
C27174 a_14358_43442# a_14456_42282# 1.03e-20
C27175 a_10341_43396# a_11551_42558# 3.11e-22
C27176 a_10765_43646# a_5742_30871# 3.49e-20
C27177 a_19237_31679# C9_N_btm 3.18e-20
C27178 a_3626_43646# a_20712_42282# 3.92e-19
C27179 a_2982_43646# a_21335_42336# 0.009024f
C27180 a_n4318_39304# a_n3565_39304# 3.96e-19
C27181 a_9145_43396# a_15051_42282# 0.001238f
C27182 a_22485_44484# RST_Z 4.8e-19
C27183 a_n2157_42858# a_n1736_42282# 0.001064f
C27184 a_743_42282# a_1606_42308# 0.088097f
C27185 a_6171_45002# a_15682_43940# 5.04e-19
C27186 a_8953_45546# a_9306_43218# 2.14e-19
C27187 a_4743_44484# a_n2661_43922# 0.008142f
C27188 a_5343_44458# a_n2661_42834# 0.038788f
C27189 a_20567_45036# a_20679_44626# 0.006083f
C27190 a_21005_45260# a_20640_44752# 4.55e-20
C27191 a_n2293_42834# a_644_44056# 1.25e-20
C27192 a_11691_44458# a_17325_44484# 0.0017f
C27193 a_8953_45002# a_10405_44172# 1.1e-20
C27194 a_2711_45572# a_16243_43396# 2.11e-19
C27195 a_n357_42282# a_21259_43561# 1.65e-19
C27196 a_20692_30879# a_14209_32519# 0.051612f
C27197 a_n971_45724# VDD 4.911799f
C27198 a_19778_44110# a_19279_43940# 0.020911f
C27199 a_11827_44484# a_19615_44636# 0.006593f
C27200 a_18315_45260# a_18579_44172# 1.04e-20
C27201 SMPL_ON_P CLK_DATA 0.200962f
C27202 a_n2109_47186# DATA[2] 0.05382f
C27203 a_6298_44484# a_9159_44484# 6.91e-21
C27204 a_8975_43940# a_9313_44734# 0.391938f
C27205 a_n2661_43370# a_n2472_43914# 0.00608f
C27206 a_n1741_47186# DATA[0] 0.051737f
C27207 a_7499_43078# a_9803_43646# 0.001386f
C27208 a_n2312_38680# a_n2216_39072# 3.1e-19
C27209 a_12465_44636# a_3232_43370# 1.26e-20
C27210 a_5497_46414# a_5066_45546# 0.05403f
C27211 a_n1151_42308# a_7418_45394# 1.53e-19
C27212 a_3094_47570# a_413_45260# 7.88e-19
C27213 a_10227_46804# a_13017_45260# 9.45e-19
C27214 a_11599_46634# a_15595_45028# 0.001416f
C27215 a_6755_46942# a_13527_45546# 0.001323f
C27216 a_765_45546# a_n357_42282# 0.209746f
C27217 a_16942_47570# a_2437_43646# 3.81e-19
C27218 a_13747_46662# a_21350_45938# 1.02e-20
C27219 a_20916_46384# a_21363_45546# 2.9e-19
C27220 a_5068_46348# a_5210_46155# 0.005572f
C27221 a_15015_46420# a_10809_44734# 6.69e-20
C27222 a_2324_44458# a_6945_45028# 0.183081f
C27223 a_18819_46122# a_19553_46090# 0.052547f
C27224 a_4190_30871# a_11206_38545# 1.56e-20
C27225 a_16245_42852# a_15890_42674# 0.001613f
C27226 a_n1630_35242# a_6123_31319# 0.036823f
C27227 a_1606_42308# a_5755_42308# 3.31e-20
C27228 a_n1059_45260# a_791_42968# 0.122941f
C27229 a_n913_45002# a_685_42968# 0.015577f
C27230 a_n2017_45002# a_1847_42826# 0.017915f
C27231 a_13249_42308# a_14635_42282# 1.46e-19
C27232 a_n2956_38680# a_n4315_30879# 0.024632f
C27233 a_n2956_39304# a_n4334_40480# 2.77e-19
C27234 a_n2661_42834# a_9801_44260# 2.25e-19
C27235 a_n699_43396# a_n97_42460# 0.152094f
C27236 a_14673_44172# a_15682_43940# 0.001963f
C27237 a_10249_46116# CLK 0.063525f
C27238 a_n357_42282# a_4921_42308# 3.76e-19
C27239 a_n2661_44458# a_4093_43548# 3.38e-20
C27240 a_644_44056# a_1115_44172# 0.013441f
C27241 a_n2661_43370# a_10695_43548# 6.82e-21
C27242 a_18479_45785# a_19339_43156# 0.001029f
C27243 a_n863_45724# a_5932_42308# 4.31e-21
C27244 a_n967_45348# a_n967_43230# 3.59e-19
C27245 a_13507_46334# a_17517_44484# 0.018934f
C27246 a_310_45028# a_n443_42852# 0.376934f
C27247 a_n2661_45546# a_1176_45572# 5.5e-19
C27248 a_13059_46348# a_14797_45144# 0.066603f
C27249 a_6755_46942# a_16922_45042# 6.22e-19
C27250 a_584_46384# a_2127_44172# 8.16e-20
C27251 a_n1991_46122# a_n913_45002# 2.75e-20
C27252 a_n1853_46287# a_n745_45366# 0.002206f
C27253 a_12465_44636# a_14581_44484# 5.1e-19
C27254 a_16327_47482# a_20640_44752# 0.044807f
C27255 a_12005_46436# a_10193_42453# 2.62e-20
C27256 a_n2497_47436# a_n1453_44318# 0.001884f
C27257 a_20820_30879# a_413_45260# 0.033659f
C27258 a_3147_46376# a_2437_43646# 1.06e-20
C27259 a_12861_44030# a_18753_44484# 2.16e-19
C27260 a_2324_44458# a_14127_45572# 6.43e-19
C27261 a_5066_45546# a_9241_45822# 2.98e-19
C27262 a_8049_45260# a_13527_45546# 0.001929f
C27263 a_10586_45546# a_11652_45724# 0.046802f
C27264 a_n357_42282# a_509_45822# 0.039776f
C27265 a_n3420_39616# a_n2860_39866# 0.002301f
C27266 a_n4064_40160# a_n4334_39392# 0.013157f
C27267 a_2905_45572# a_3160_47472# 0.54473f
C27268 a_n971_45724# a_6491_46660# 0.011282f
C27269 a_2952_47436# a_n1151_42308# 0.068429f
C27270 a_2063_45854# a_3785_47178# 0.001458f
C27271 a_n237_47217# a_6151_47436# 0.360224f
C27272 a_n1741_47186# a_9067_47204# 0.012401f
C27273 a_n2946_39866# a_n2302_39866# 6.68e-19
C27274 a_5932_42308# a_6886_37412# 5.75e-19
C27275 a_n1630_35242# EN_VIN_BSTR_P 0.009334f
C27276 a_17665_42852# VDD 0.006567f
C27277 a_n4209_39590# a_n4251_39616# 0.00226f
C27278 a_14539_43914# a_16795_42852# 0.037061f
C27279 a_n2293_43922# a_n4318_38680# 2.08e-19
C27280 en_comp a_14456_42282# 8.68e-21
C27281 a_17517_44484# a_21855_43396# 3.12e-22
C27282 a_n2661_42834# a_n1545_43230# 3.82e-19
C27283 a_19789_44512# a_15743_43084# 2.77e-21
C27284 a_n356_44636# a_10341_42308# 1.92e-20
C27285 a_8049_45260# EN_OFFSET_CAL 1.15e-20
C27286 a_n913_45002# a_14113_42308# 0.029759f
C27287 a_n1059_45260# a_15051_42282# 6.54e-19
C27288 a_n2017_45002# a_15486_42560# 0.005473f
C27289 a_20205_31679# a_19864_35138# 9.62e-21
C27290 a_n2661_42282# a_6031_43396# 0.036698f
C27291 a_742_44458# a_873_42968# 7.93e-21
C27292 a_5891_43370# a_7227_42852# 0.129383f
C27293 a_n2293_46634# a_3353_43940# 5.23e-19
C27294 a_5263_45724# a_5111_44636# 0.00615f
C27295 a_11415_45002# a_14112_44734# 1.45e-20
C27296 a_n881_46662# a_n2129_43609# 1.93e-21
C27297 a_15599_45572# a_16147_45260# 7.22e-19
C27298 a_n1613_43370# a_n2267_43396# 0.04778f
C27299 a_n755_45592# a_1307_43914# 0.007948f
C27300 a_n863_45724# a_1423_45028# 0.113534f
C27301 a_310_45028# a_375_42282# 0.078376f
C27302 a_n2956_39304# a_n2661_44458# 1.51e-20
C27303 a_n2956_38680# a_n4318_40392# 0.024261f
C27304 a_8049_45260# a_16922_45042# 8.87e-20
C27305 a_7499_43078# a_n913_45002# 0.548687f
C27306 a_17339_46660# a_19006_44850# 1.58e-20
C27307 a_16333_45814# a_16211_45572# 3.16e-19
C27308 a_12741_44636# a_13213_44734# 0.00239f
C27309 a_3775_45552# a_2382_45260# 2.04e-19
C27310 a_2711_45572# a_3232_43370# 0.002535f
C27311 a_n2293_45546# a_2304_45348# 0.032829f
C27312 a_10903_43370# a_12883_44458# 6.65e-20
C27313 a_n1435_47204# a_6755_46942# 0.006483f
C27314 a_7754_39964# VDD 0.848281f
C27315 a_n4209_37414# C7_P_btm 1.43e-20
C27316 a_n3565_37414# C9_P_btm 3.18e-20
C27317 a_11599_46634# a_10150_46912# 3.38e-21
C27318 a_n3420_37984# VIN_P 0.06991f
C27319 a_19594_46812# a_20843_47204# 5.41e-20
C27320 a_3726_37500# a_n923_35174# 0.029905f
C27321 a_4883_46098# a_4817_46660# 1.29e-19
C27322 a_n4209_38216# VCM 0.035453f
C27323 CAL_N a_22609_38406# 0.204621f
C27324 a_22521_40055# a_22469_39537# 0.037283f
C27325 a_22521_40599# CAL_P 6.35e-19
C27326 a_22459_39145# a_22821_38993# 0.013073f
C27327 a_n1613_43370# a_491_47026# 0.038998f
C27328 a_6575_47204# a_8035_47026# 3.94e-19
C27329 a_6151_47436# a_8270_45546# 0.142873f
C27330 a_n1151_42308# a_12991_46634# 0.013856f
C27331 a_2063_45854# a_3090_45724# 0.002495f
C27332 a_n881_46662# a_288_46660# 0.001197f
C27333 a_n3565_38216# VREF 0.057702f
C27334 a_768_44030# a_n743_46660# 0.028134f
C27335 a_n2267_43396# a_n1533_42852# 4.05e-20
C27336 a_9145_43396# a_13749_43396# 3.66e-19
C27337 a_n2293_43922# a_11551_42558# 1.93e-19
C27338 a_9313_44734# a_15803_42450# 8.69e-20
C27339 a_n2065_43946# a_n4318_37592# 2.96e-22
C27340 a_n356_44636# a_18057_42282# 0.087032f
C27341 a_n1761_44111# a_n1736_42282# 3.18e-19
C27342 a_n2293_45010# VDD 1.885f
C27343 a_8685_43396# a_16409_43396# 6.54e-20
C27344 a_19479_31679# EN_OFFSET_CAL 3.97e-20
C27345 a_8333_44056# a_8495_42852# 5.85e-22
C27346 a_3357_43084# DATA[5] 0.032568f
C27347 a_14579_43548# a_14537_43646# 0.001675f
C27348 a_3539_42460# a_743_42282# 0.054149f
C27349 a_526_44458# a_9672_43914# 1.87e-19
C27350 a_20692_30879# a_17730_32519# 0.05146f
C27351 a_18787_45572# a_11691_44458# 1.34e-19
C27352 a_12549_44172# a_18083_42858# 5.88e-21
C27353 w_11334_34010# a_1606_42308# 0.001329f
C27354 a_n971_45724# a_n784_42308# 0.006301f
C27355 a_3065_45002# a_2809_45028# 0.006555f
C27356 a_10227_46804# a_10793_43218# 2.95e-19
C27357 a_6755_46942# a_15743_43084# 7.96e-20
C27358 a_n745_45366# a_n2661_43370# 0.005292f
C27359 a_5147_45002# a_6125_45348# 1.1e-19
C27360 a_5111_44636# a_5837_45348# 0.001223f
C27361 a_4927_45028# a_5365_45348# 0.013015f
C27362 a_10193_42453# a_9313_44734# 0.078654f
C27363 a_8191_45002# a_1423_45028# 1.9e-20
C27364 a_13777_45326# a_14537_43396# 4.1e-19
C27365 a_9482_43914# a_15415_45028# 0.002812f
C27366 a_13556_45296# a_14797_45144# 2.59e-20
C27367 a_3090_45724# a_14955_43396# 0.07523f
C27368 SMPL_ON_P a_n1630_35242# 6.11548f
C27369 a_12891_46348# a_11387_46155# 1.97e-20
C27370 a_n2109_47186# a_n2293_45546# 4.56e-21
C27371 a_5807_45002# a_8016_46348# 3.22e-19
C27372 a_11309_47204# a_10903_43370# 1.95e-19
C27373 a_6755_46942# a_13885_46660# 0.078788f
C27374 a_12816_46660# a_13607_46688# 3.63e-19
C27375 a_n2497_47436# a_n863_45724# 0.337007f
C27376 a_n1925_46634# a_1823_45246# 0.001679f
C27377 a_n743_46660# a_1176_45822# 0.08607f
C27378 a_n2438_43548# a_1208_46090# 0.005695f
C27379 a_n133_46660# a_805_46414# 0.001959f
C27380 a_n2661_46634# a_3147_46376# 8.89e-20
C27381 a_22612_30879# a_4185_45028# 2.99e-19
C27382 a_n881_46662# a_15015_46420# 2.18e-20
C27383 SMPL_ON_P a_n2661_45546# 0.002242f
C27384 a_33_46660# a_376_46348# 5.66e-19
C27385 a_171_46873# a_472_46348# 0.008963f
C27386 a_9313_44734# VDD 0.389068f
C27387 a_18429_43548# a_18504_43218# 1.16e-19
C27388 a_16137_43396# a_17665_42852# 0.001078f
C27389 a_n1076_43230# a_133_42852# 1.24e-19
C27390 a_10341_42308# a_12379_42858# 2.14e-19
C27391 a_10922_42852# a_12089_42308# 8.07e-21
C27392 a_3626_43646# a_6171_42473# 0.003703f
C27393 a_3080_42308# a_3905_42308# 8.29e-20
C27394 a_n97_42460# a_11551_42558# 0.095523f
C27395 a_3483_46348# a_13460_43230# 7.53e-19
C27396 a_4185_45028# a_12895_43230# 1.02e-20
C27397 a_11691_44458# a_18287_44626# 0.032949f
C27398 a_18479_45785# a_17973_43940# 2.56e-22
C27399 a_13259_45724# a_12281_43396# 3.97e-20
C27400 SMPL_ON_P a_n3607_37440# 7.77e-21
C27401 a_n2661_44458# a_10157_44484# 0.00786f
C27402 a_16019_45002# a_11967_42832# 8.44e-20
C27403 a_327_44734# a_175_44278# 0.001132f
C27404 a_5937_45572# a_9127_43156# 5.33e-21
C27405 a_8199_44636# a_8952_43230# 1.83e-19
C27406 a_526_44458# a_743_42282# 0.042759f
C27407 a_n2017_45002# a_5244_44056# 3.28e-21
C27408 a_n1059_45260# a_3905_42865# 0.01898f
C27409 a_18494_42460# a_n356_44636# 0.003788f
C27410 a_742_44458# a_n699_43396# 0.047576f
C27411 a_10227_46804# a_20107_45572# 2.37e-20
C27412 a_4651_46660# a_2711_45572# 5.93e-20
C27413 a_11415_45002# a_19335_46494# 3.95e-20
C27414 a_3483_46348# a_8349_46414# 4.04e-20
C27415 a_n237_47217# a_5111_44636# 6.91e-20
C27416 a_15009_46634# a_13259_45724# 9.93e-20
C27417 a_14976_45028# a_15194_46482# 5.51e-19
C27418 a_21350_47026# a_6945_45028# 1.62e-19
C27419 a_18900_46660# a_10809_44734# 8.2e-19
C27420 a_12861_44030# a_2437_43646# 0.022753f
C27421 a_2107_46812# a_7499_43078# 6.63e-20
C27422 a_13885_46660# a_8049_45260# 5.7e-22
C27423 a_2905_45572# a_413_45260# 0.124898f
C27424 a_n1151_42308# a_n143_45144# 0.002247f
C27425 a_n881_46662# a_16333_45814# 0.04285f
C27426 a_16327_47482# a_21188_45572# 0.227468f
C27427 a_13381_47204# a_3357_43084# 1.79e-19
C27428 a_584_46384# a_2382_45260# 0.185451f
C27429 a_2063_45854# a_2274_45254# 2.23e-19
C27430 a_12549_44172# a_11688_45572# 6.24e-20
C27431 a_5164_46348# a_5204_45822# 0.132894f
C27432 a_12741_44636# a_18819_46122# 2.26e-20
C27433 a_3524_46660# a_3775_45552# 1.42e-20
C27434 a_3877_44458# a_4099_45572# 0.01632f
C27435 a_n743_46660# a_11652_45724# 2.53e-19
C27436 a_5342_30871# a_16104_42674# 4.45e-20
C27437 a_n4318_38680# a_n3420_39616# 0.02534f
C27438 a_20974_43370# VDD 0.550101f
C27439 a_14401_32519# RST_Z 0.048069f
C27440 a_526_44458# a_5755_42308# 3.22e-19
C27441 a_n357_42282# a_13291_42460# 0.008613f
C27442 a_9290_44172# a_11633_42308# 0.001629f
C27443 a_n2293_42834# a_104_43370# 0.003003f
C27444 a_22612_30879# VREF_GND 0.168163f
C27445 a_21588_30879# VCM 0.179761f
C27446 a_n356_44636# a_3499_42826# 1.72e-20
C27447 a_11967_42832# a_18245_44484# 1.94e-19
C27448 a_10193_42453# a_18599_43230# 0.003065f
C27449 a_n743_46660# DATA[0] 1.07e-19
C27450 a_601_46902# VDD 0.204253f
C27451 a_n2661_42834# a_453_43940# 0.04708f
C27452 a_n1925_46634# DATA[2] 9.45e-20
C27453 a_20362_44736# a_20766_44850# 0.051162f
C27454 a_n2661_43922# a_1414_42308# 0.010195f
C27455 a_20640_44752# a_20835_44721# 0.20669f
C27456 a_20159_44458# a_19279_43940# 0.06519f
C27457 a_n2661_43370# a_n2433_43396# 0.021188f
C27458 a_n913_45002# a_15781_43660# 8.25e-21
C27459 a_10903_43370# a_10490_45724# 0.057318f
C27460 a_19321_45002# a_21005_45260# 0.002433f
C27461 a_13661_43548# a_11827_44484# 0.120515f
C27462 a_13747_46662# a_21359_45002# 0.060042f
C27463 a_14180_46812# a_2437_43646# 1.36e-20
C27464 a_3877_44458# a_5365_45348# 6.25e-22
C27465 a_11387_46155# a_11322_45546# 4.47e-19
C27466 a_6755_46942# a_10775_45002# 6.89e-22
C27467 a_20916_46384# a_19778_44110# 2.1e-21
C27468 a_8270_45546# a_5111_44636# 0.035253f
C27469 a_15227_44166# a_n913_45002# 1.05e-19
C27470 a_6945_45028# a_6667_45809# 0.015851f
C27471 a_526_44458# a_2277_45546# 5.37e-21
C27472 a_12465_44636# a_8975_43940# 3.06e-19
C27473 a_n1613_43370# a_n2267_44484# 0.025052f
C27474 a_n881_46662# a_n2129_44697# 1.78e-19
C27475 a_12816_46660# a_413_45260# 4.83e-21
C27476 a_n1151_42308# a_n2293_43922# 1.39e-19
C27477 a_12594_46348# a_10193_42453# 1.09e-19
C27478 a_10249_46116# a_10951_45334# 8.11e-22
C27479 a_11189_46129# a_11652_45724# 0.00549f
C27480 a_17303_42282# a_19332_42282# 3.68e-19
C27481 a_18817_42826# RST_Z 4.49e-21
C27482 a_18057_42282# a_18727_42674# 0.003581f
C27483 a_18599_43230# VDD 0.197104f
C27484 a_n2293_42834# a_4156_43218# 6.26e-20
C27485 a_n2956_37592# a_n1736_42282# 8.96e-21
C27486 en_comp a_n3674_38216# 0.026738f
C27487 a_n2956_38216# a_n2860_37984# 0.001353f
C27488 a_n2810_45028# a_n4318_37592# 0.023097f
C27489 a_12594_46348# VDD 1.03351f
C27490 a_18287_44626# a_4190_30871# 4.63e-21
C27491 a_n2661_44458# a_685_42968# 1.08e-21
C27492 a_11341_43940# a_15493_43940# 0.216602f
C27493 a_n2661_43922# a_12281_43396# 2.21e-20
C27494 a_n2017_45002# a_n473_42460# 0.017082f
C27495 a_n1059_45260# a_n961_42308# 3.29e-21
C27496 a_n967_45348# a_n2104_42282# 4.03e-19
C27497 a_17973_43940# a_14021_43940# 4.61e-20
C27498 a_14955_43940# a_15037_44260# 0.003935f
C27499 a_n2661_42282# a_6671_43940# 0.002068f
C27500 a_1467_44172# a_n97_42460# 0.190191f
C27501 a_9313_44734# a_16137_43396# 0.044229f
C27502 a_n699_43396# a_n901_43156# 6.3e-20
C27503 a_5937_45572# CLK 1.52e-19
C27504 a_11827_44484# a_10835_43094# 8.97e-20
C27505 a_3422_30871# a_2982_43646# 0.140944f
C27506 a_11823_42460# a_7174_31319# 9.76e-21
C27507 a_15433_44458# a_15095_43370# 1.02e-20
C27508 a_526_44458# a_626_44172# 0.180416f
C27509 a_11525_45546# a_11688_45572# 0.011381f
C27510 a_n2293_46098# a_n2267_44484# 2.71e-20
C27511 a_n2157_46122# a_n2129_44697# 8.63e-21
C27512 a_18285_46348# a_18248_44752# 3.14e-21
C27513 a_4185_45028# a_11827_44484# 0.03083f
C27514 a_3090_45724# a_n2661_42834# 0.164804f
C27515 a_n1151_42308# a_n97_42460# 8.22e-19
C27516 a_n1991_46122# a_n2661_44458# 1.24e-22
C27517 a_17339_46660# a_18374_44850# 0.009147f
C27518 a_6755_46942# a_16789_44484# 2.63e-19
C27519 a_12465_44636# a_14485_44260# 0.009374f
C27520 a_8049_45260# a_10775_45002# 7.17e-20
C27521 a_12549_44172# a_12429_44172# 0.137881f
C27522 a_768_44030# a_11750_44172# 0.00229f
C27523 a_12891_46348# a_13483_43940# 0.062818f
C27524 a_n2840_45546# a_n2661_45010# 3.35e-19
C27525 a_n2810_45572# a_n2840_45002# 4.88e-19
C27526 a_10490_45724# a_12016_45572# 0.003469f
C27527 a_n1151_42308# a_n2661_46098# 0.024549f
C27528 a_4883_46098# a_11309_47204# 0.012799f
C27529 a_16327_47482# a_19321_45002# 0.925259f
C27530 a_7754_38968# a_3754_38470# 0.209356f
C27531 a_n4209_39304# C9_P_btm 3.29e-19
C27532 a_13507_46334# a_12549_44172# 0.363125f
C27533 a_17591_47464# a_5807_45002# 0.001206f
C27534 a_n971_45724# a_4646_46812# 0.303249f
C27535 a_2063_45854# a_3699_46634# 7.49e-20
C27536 a_2952_47436# a_3177_46902# 1.43e-19
C27537 a_3160_47472# a_2443_46660# 0.019074f
C27538 a_2905_45572# a_2609_46660# 0.027251f
C27539 a_584_46384# a_3524_46660# 4.24e-20
C27540 a_12861_44030# a_n2661_46634# 0.03828f
C27541 a_n1741_47186# a_5167_46660# 2.91e-20
C27542 a_n2109_47186# a_5732_46660# 0.009505f
C27543 a_n4064_39616# C0_P_btm 3.27e-20
C27544 a_22397_42558# VDD 0.006424f
C27545 a_6197_43396# a_6547_43396# 0.216095f
C27546 a_11967_42832# a_13814_43218# 0.001842f
C27547 a_18184_42460# a_18907_42674# 0.071964f
C27548 a_18494_42460# a_18727_42674# 0.031761f
C27549 a_n2956_37592# a_n4209_37414# 0.145558f
C27550 a_15037_45618# VDD 0.08759f
C27551 a_14021_43940# a_22591_43396# 0.057848f
C27552 a_n356_44636# a_3318_42354# 1.4e-19
C27553 a_n2661_42834# a_n2472_42282# 2.95e-19
C27554 a_16922_45042# a_13258_32519# 4.48e-20
C27555 a_n2810_45028# a_n4334_37440# 6.16e-20
C27556 a_6293_42852# a_7287_43370# 1.04e-20
C27557 a_3626_43646# a_3457_43396# 0.067226f
C27558 a_6031_43396# a_7112_43396# 0.101963f
C27559 a_12741_44636# a_11341_43940# 9.61e-20
C27560 a_19692_46634# a_17538_32519# 0.002f
C27561 a_13259_45724# a_14112_44734# 0.001601f
C27562 a_n1059_45260# a_5147_45002# 2.48e-21
C27563 a_n2017_45002# a_5111_44636# 0.024598f
C27564 a_10227_46804# a_10083_42826# 0.292997f
C27565 a_6472_45840# a_5883_43914# 3.93e-22
C27566 a_13904_45546# a_11691_44458# 4.03e-21
C27567 a_2324_44458# a_895_43940# 0.011941f
C27568 a_n37_45144# a_413_45260# 0.021944f
C27569 a_n1613_43370# a_n2472_42826# 6.43e-21
C27570 a_6598_45938# a_6298_44484# 0.001025f
C27571 a_2711_45572# a_8975_43940# 6.21e-21
C27572 a_12549_44172# a_21855_43396# 0.001702f
C27573 a_7499_43078# a_n2661_44458# 0.059442f
C27574 a_3877_44458# a_8189_46660# 9.93e-21
C27575 a_9313_45822# a_9823_46155# 6.69e-21
C27576 a_13747_46662# a_14226_46660# 0.001089f
C27577 a_5807_45002# a_15312_46660# 3.46e-19
C27578 a_n2312_39304# a_n2293_46098# 0.027561f
C27579 a_7577_46660# a_8492_46660# 0.118423f
C27580 a_5732_46660# a_5841_46660# 0.007416f
C27581 a_5907_46634# a_6086_46660# 0.007399f
C27582 a_6540_46812# a_6999_46987# 6.64e-19
C27583 a_n1435_47204# a_8953_45546# 5.89e-20
C27584 a_10227_46804# a_3483_46348# 0.057984f
C27585 a_6151_47436# a_13759_46122# 3.56e-19
C27586 a_4915_47217# a_14275_46494# 0.01257f
C27587 a_n2433_43396# COMP_P 0.001151f
C27588 a_15682_43940# a_15959_42545# 2.38e-19
C27589 a_16409_43396# a_17333_42852# 1.86e-19
C27590 a_17499_43370# a_17595_43084# 0.002317f
C27591 a_743_42282# a_8605_42826# 5.66e-20
C27592 a_17324_43396# a_16795_42852# 1.3e-19
C27593 a_16137_43396# a_18599_43230# 0.005055f
C27594 a_n1641_43230# a_n1736_43218# 0.049827f
C27595 a_n901_43156# a_n4318_38680# 7.68e-22
C27596 a_11341_43940# a_5742_30871# 0.0019f
C27597 a_n2267_43396# a_n1736_42282# 3.76e-21
C27598 a_18114_32519# VDD 0.550312f
C27599 a_n1423_42826# a_n1545_43230# 3.16e-19
C27600 a_n1853_43023# a_n967_43230# 8.59e-19
C27601 a_15743_43084# a_15279_43071# 1.83e-19
C27602 a_4361_42308# a_5755_42852# 2.34e-20
C27603 a_n2661_43370# a_n2433_44484# 0.018595f
C27604 a_3232_43370# a_9241_44734# 8.2e-19
C27605 a_7705_45326# a_7640_43914# 5.79e-20
C27606 a_17023_45118# a_11691_44458# 0.00304f
C27607 a_18587_45118# a_11827_44484# 5.85e-20
C27608 a_19778_44110# a_21101_45002# 0.008451f
C27609 a_18494_42460# a_20567_45036# 5.4e-19
C27610 a_16922_45042# a_20193_45348# 0.328274f
C27611 a_16501_45348# a_16237_45028# 3.62e-19
C27612 a_526_44458# a_2813_43396# 0.013054f
C27613 a_2274_45254# a_n2661_42834# 1.64e-20
C27614 a_20623_45572# a_19279_43940# 7.39e-21
C27615 a_20731_45938# a_20640_44752# 2.23e-21
C27616 a_n2438_43548# a_n1630_35242# 1.24e-19
C27617 a_20692_30879# a_17538_32519# 0.05141f
C27618 a_16327_47482# a_17531_42308# 7.43e-19
C27619 a_n1613_43370# a_9223_42460# 0.007135f
C27620 a_5093_45028# a_5343_44458# 4.13e-19
C27621 a_10227_46804# a_15761_42308# 2.95e-19
C27622 a_10193_42453# a_17737_43940# 0.02461f
C27623 a_11823_42460# a_10729_43914# 8.14e-20
C27624 a_11652_45724# a_11750_44172# 6.11e-20
C27625 a_12427_45724# a_10949_43914# 3.38e-21
C27626 a_7229_43940# a_5891_43370# 1.39e-19
C27627 a_n2293_42834# a_949_44458# 4.61e-20
C27628 w_1575_34946# a_n3420_37440# 2.64e-19
C27629 a_3090_45724# a_17715_44484# 0.108364f
C27630 a_765_45546# a_3147_46376# 2.61e-20
C27631 a_17339_46660# a_3483_46348# 7.08e-22
C27632 a_22591_46660# a_12741_44636# 0.0686f
C27633 a_11415_45002# a_22959_46660# 3.29e-19
C27634 a_4883_46098# a_10490_45724# 7.84e-20
C27635 a_10227_46804# a_14495_45572# 0.001891f
C27636 a_n2661_46634# a_310_45028# 4.45e-20
C27637 a_n2438_43548# a_n2661_45546# 0.065227f
C27638 a_12156_46660# a_10903_43370# 8.13e-19
C27639 a_n881_46662# a_6472_45840# 0.179318f
C27640 a_20202_43084# a_21076_30879# 6.04e-20
C27641 a_n1613_43370# a_6511_45714# 0.017587f
C27642 a_n2293_46634# a_n452_45724# 0.002803f
C27643 a_15559_46634# a_2324_44458# 0.012623f
C27644 a_8667_46634# a_5066_45546# 4.03e-20
C27645 a_n1925_46634# a_n2293_45546# 7.25e-20
C27646 a_11453_44696# a_7499_43078# 0.02227f
C27647 a_17737_43940# VDD 0.285511f
C27648 a_5649_42852# a_15890_42674# 5.19e-20
C27649 a_16823_43084# a_4958_30871# 5.65e-19
C27650 a_4190_30871# a_17124_42282# 7.43e-20
C27651 a_n2293_42282# a_n2472_42282# 0.163758f
C27652 a_19700_43370# a_19511_42282# 6.2e-21
C27653 a_4361_42308# a_10149_42308# 6.19e-19
C27654 a_743_42282# a_16104_42674# 0.002282f
C27655 a_15743_43084# a_13258_32519# 1.74e-19
C27656 a_9482_43914# a_9801_43940# 8.96e-19
C27657 a_13213_44734# a_13468_44734# 0.005172f
C27658 a_18374_44850# a_18579_44172# 7.6e-20
C27659 a_18443_44721# a_18681_44484# 0.001705f
C27660 a_949_44458# a_1115_44172# 0.016355f
C27661 a_742_44458# a_1467_44172# 0.018499f
C27662 a_21496_47436# SINGLE_ENDED 0.055146f
C27663 a_22612_30879# a_22469_40625# 7.32e-20
C27664 a_12465_44636# VDD 0.773277f
C27665 a_327_44734# a_n97_42460# 2.31e-20
C27666 a_n699_43396# a_n984_44318# 2.34e-20
C27667 a_n913_45002# a_1756_43548# 3.6e-21
C27668 a_n2017_45002# a_4235_43370# 2.25e-19
C27669 a_n1059_45260# a_4093_43548# 0.001865f
C27670 a_n357_42282# a_13460_43230# 0.007447f
C27671 a_4883_46098# START 2.42e-19
C27672 a_1307_43914# a_5326_44056# 0.001893f
C27673 a_21811_47423# RST_Z 5.42e-20
C27674 a_n443_42852# a_9127_43156# 0.001064f
C27675 a_3357_43084# a_3626_43646# 0.018539f
C27676 a_n2661_46098# a_327_44734# 1.48e-20
C27677 a_1799_45572# a_1667_45002# 1.16e-19
C27678 a_2905_45572# a_2779_44458# 7.14e-20
C27679 a_15227_44166# a_15903_45785# 0.005114f
C27680 a_3090_45724# a_15861_45028# 0.125763f
C27681 a_14976_45028# a_8696_44636# 2.84e-19
C27682 a_12861_44030# a_19113_45348# 0.003723f
C27683 a_12465_44636# a_14309_45348# 1.46e-20
C27684 a_16327_47482# a_18184_42460# 0.168018f
C27685 a_n2661_46634# a_11787_45002# 0.004953f
C27686 a_18819_46122# a_16375_45002# 0.002016f
C27687 a_167_45260# a_1990_45899# 0.006879f
C27688 a_17583_46090# a_18051_46116# 3.98e-20
C27689 a_n2293_46098# a_6511_45714# 7.32e-20
C27690 a_2443_46660# a_413_45260# 0.020902f
C27691 a_15368_46634# a_16680_45572# 2.35e-20
C27692 a_13747_46662# a_15415_45028# 2.47e-20
C27693 a_13661_43548# a_15595_45028# 0.214904f
C27694 a_768_44030# a_2809_45348# 0.001559f
C27695 a_2107_46812# a_4558_45348# 1.43e-21
C27696 a_2063_45854# a_4743_44484# 3.42e-21
C27697 a_n2293_46634# a_8953_45002# 4.11e-20
C27698 a_22223_43396# RST_Z 5.55e-20
C27699 a_10533_42308# a_11551_42558# 2.25e-19
C27700 a_10723_42308# a_5742_30871# 0.185564f
C27701 a_1606_42308# a_13258_32519# 0.001369f
C27702 a_5342_30871# VDAC_N 0.011613f
C27703 a_13887_32519# VDD 0.424101f
C27704 a_17364_32525# C8_N_btm 7.96e-19
C27705 a_961_42354# a_7174_31319# 4.84e-21
C27706 a_n4318_38216# a_n4334_39616# 1.11e-19
C27707 a_5534_30871# VDAC_P 0.004852f
C27708 a_20528_46660# VDD 0.077608f
C27709 a_3499_42826# a_3820_44260# 5.31e-19
C27710 a_22000_46634# RST_Z 3.42e-20
C27711 a_16922_45042# a_20301_43646# 0.00515f
C27712 a_n356_44636# a_6197_43396# 1.09e-20
C27713 a_21363_46634# SINGLE_ENDED 2.03e-20
C27714 a_11691_44458# a_19268_43646# 1.97e-21
C27715 a_20193_45348# a_15743_43084# 0.060559f
C27716 a_n2293_42834# a_n1076_43230# 0.01241f
C27717 a_1307_43914# a_10083_42826# 4.67e-20
C27718 a_9838_44484# a_9803_43646# 7.04e-22
C27719 a_10157_44484# a_9145_43396# 4.85e-21
C27720 a_20692_30879# a_22465_38105# 5.07e-19
C27721 a_n2661_42834# a_n1821_43396# 4.8e-19
C27722 a_7499_43078# a_8325_42308# 2.16e-19
C27723 a_2711_45572# a_15803_42450# 1.02e-20
C27724 a_10193_42453# a_8515_42308# 1.05e-20
C27725 a_9482_43914# a_12545_42858# 1.33e-20
C27726 a_1423_45028# a_7765_42852# 5.7e-21
C27727 a_17339_46660# a_17719_45144# 8.89e-19
C27728 a_14035_46660# a_11691_44458# 4.42e-21
C27729 a_765_45546# a_17613_45144# 1.04e-21
C27730 a_19692_46634# a_19721_31679# 5.55e-20
C27731 a_18285_46348# a_16922_45042# 4.22e-21
C27732 a_10903_43370# a_6171_45002# 0.041534f
C27733 a_n2956_38680# a_n2017_45002# 7.75e-22
C27734 a_12549_44172# a_20637_44484# 8.68e-20
C27735 a_n1613_43370# a_n2065_43946# 0.30437f
C27736 a_2711_45572# a_10193_42453# 0.218272f
C27737 a_6511_45714# a_7230_45938# 0.088127f
C27738 a_3775_45552# a_4880_45572# 1.54e-21
C27739 a_6667_45809# a_6812_45938# 0.057222f
C27740 a_6472_45840# a_8162_45546# 3.95e-19
C27741 a_167_45260# a_1145_45348# 5.7e-19
C27742 a_18819_46122# a_413_45260# 1.56e-20
C27743 a_19321_45002# a_20835_44721# 7.19e-19
C27744 a_9625_46129# a_8953_45002# 0.004507f
C27745 a_16375_45002# a_16223_45938# 3.86e-20
C27746 a_13747_46662# a_19279_43940# 0.048937f
C27747 a_8199_44636# a_11787_45002# 2.96e-20
C27748 a_3483_46348# a_1307_43914# 0.095243f
C27749 a_2324_44458# a_3065_45002# 0.017588f
C27750 a_n3690_38528# a_n3690_38304# 0.052468f
C27751 a_n3420_38528# a_n3565_38216# 0.035254f
C27752 a_n4064_38528# a_n4209_38216# 0.028013f
C27753 a_n3565_38502# a_n3420_37984# 0.028236f
C27754 a_n4209_38502# a_n4064_37984# 0.028133f
C27755 a_n4064_40160# a_n3565_37414# 4.29714f
C27756 a_n1741_47186# a_12549_44172# 9.64e-19
C27757 a_n971_45724# a_9804_47204# 1.23e-20
C27758 a_327_47204# a_n881_46662# 3.68e-20
C27759 a_1209_47178# a_n1613_43370# 0.006245f
C27760 a_3381_47502# a_2747_46873# 2.58e-20
C27761 a_2063_45854# a_2583_47243# 2.21e-19
C27762 a_n1151_42308# a_n310_47243# 3.07e-19
C27763 a_8515_42308# VDD 0.194691f
C27764 a_n4315_30879# a_n3420_37440# 0.039346f
C27765 a_15673_47210# a_16241_47178# 0.183195f
C27766 a_15811_47375# a_16327_47482# 0.038827f
C27767 a_5934_30871# RST_Z 0.003901f
C27768 a_13717_47436# a_18479_47436# 2.23e-19
C27769 a_15507_47210# a_16023_47582# 0.109156f
C27770 a_11599_46634# a_16763_47508# 4.36e-20
C27771 a_5742_30871# C1_P_btm 0.026156f
C27772 a_12861_44030# a_18143_47464# 0.394543f
C27773 a_13487_47204# a_10227_46804# 2.54e-19
C27774 a_2711_45572# VDD 1.22011f
C27775 a_14539_43914# a_18504_43218# 1.37e-19
C27776 a_7499_43940# a_7287_43370# 8.47e-19
C27777 a_15493_43940# a_10341_43396# 0.051273f
C27778 a_15682_43940# a_16243_43396# 0.013782f
C27779 a_17737_43940# a_16137_43396# 2.97e-21
C27780 a_11967_42832# a_12895_43230# 0.035759f
C27781 a_10227_46804# a_16664_43396# 5.15e-19
C27782 a_12861_44030# a_21259_43561# 3.06e-20
C27783 a_3090_45724# a_20623_43914# 4.66e-20
C27784 a_9159_45572# a_8953_45002# 0.001432f
C27785 a_20692_30879# a_19721_31679# 0.051673f
C27786 a_20841_45814# a_21350_45938# 2.6e-19
C27787 a_20273_45572# a_20719_45572# 2.28e-19
C27788 a_n2293_46634# a_3626_43646# 0.012347f
C27789 a_3483_46348# a_18579_44172# 2.2e-21
C27790 a_6194_45824# a_n2661_43370# 0.002009f
C27791 a_2711_45572# a_14309_45348# 0.002115f
C27792 a_n1151_42308# a_n901_43156# 0.01984f
C27793 C1_P_btm C0_dummy_P_btm 1.2494f
C27794 C3_P_btm C0_N_btm 3.77e-19
C27795 C6_P_btm C3_N_btm 4.24e-19
C27796 C4_P_btm C1_N_btm 1.59e-19
C27797 a_15811_47375# a_16434_46987# 8.78e-19
C27798 a_1799_45572# a_2959_46660# 3.87e-20
C27799 a_n2661_46634# a_5894_47026# 1.44e-19
C27800 a_n785_47204# a_n1853_46287# 2.37e-20
C27801 a_12861_44030# a_765_45546# 0.190301f
C27802 CAL_P VIN_N 0.001176f
C27803 a_16241_47178# a_16388_46812# 1.22e-19
C27804 a_16327_47482# a_13059_46348# 5.25e-20
C27805 a_n743_46660# a_5167_46660# 2.34e-20
C27806 a_1983_46706# a_2162_46660# 0.006978f
C27807 EN_VIN_BSTR_N VDD 1.13406f
C27808 a_8128_46384# a_8189_46660# 6.01e-19
C27809 a_11530_34132# RST_Z 0.01695f
C27810 a_n1151_42308# a_11415_45002# 2.84e-20
C27811 a_n971_45724# a_n901_46420# 0.021388f
C27812 a_n2109_47186# a_1138_42852# 1.13e-20
C27813 a_5807_45002# a_10428_46928# 0.002901f
C27814 a_n1925_46634# a_5732_46660# 0.006885f
C27815 a_2443_46660# a_2609_46660# 0.579196f
C27816 a_15673_47210# a_16721_46634# 2.97e-19
C27817 a_10227_46804# a_14513_46634# 0.004612f
C27818 a_11453_44696# a_15227_44166# 0.979188f
C27819 a_16759_43396# a_4361_42308# 7.84e-21
C27820 a_n97_42460# a_133_42852# 0.012177f
C27821 a_19700_43370# a_21259_43561# 8.8e-21
C27822 a_18783_43370# a_743_42282# 1.15e-20
C27823 a_15743_43084# a_20301_43646# 1.96e-20
C27824 a_19268_43646# a_4190_30871# 0.035721f
C27825 a_3626_43646# a_5342_30871# 0.08847f
C27826 a_327_44734# a_742_44458# 0.005551f
C27827 a_413_45260# a_949_44458# 0.018785f
C27828 a_n2312_39304# a_n1736_42282# 3.28e-20
C27829 a_12741_44636# a_10341_43396# 4.16e-20
C27830 a_4558_45348# a_n2661_44458# 0.001813f
C27831 a_n467_45028# a_n699_43396# 7.07e-21
C27832 a_18479_45785# a_9313_44734# 5.83e-19
C27833 a_19692_46634# a_22591_43396# 2.85e-19
C27834 a_3503_45724# a_3499_42826# 9.02e-22
C27835 a_n2312_40392# a_n4318_37592# 0.025292f
C27836 a_13159_45002# a_11827_44484# 9.25e-21
C27837 a_8696_44636# a_15433_44458# 0.001482f
C27838 a_16375_45002# a_11341_43940# 4.26e-20
C27839 a_10227_46804# a_n357_42282# 0.103631f
C27840 a_n743_46660# a_518_46482# 7.72e-19
C27841 a_14180_46812# a_765_45546# 4.49e-21
C27842 a_n1925_46634# a_n914_46116# 5.09e-20
C27843 a_4791_45118# a_6511_45714# 0.034343f
C27844 a_4915_47217# a_6194_45824# 1.57e-22
C27845 a_n237_47217# a_9049_44484# 0.001811f
C27846 a_3785_47178# a_3775_45552# 7.52e-20
C27847 a_11309_47204# a_11608_46482# 6.71e-19
C27848 a_19692_46634# a_20731_47026# 9.71e-20
C27849 a_16388_46812# a_16721_46634# 0.222024f
C27850 a_10467_46802# a_3483_46348# 9.89e-19
C27851 a_6491_46660# a_2711_45572# 1.46e-21
C27852 a_12549_44172# a_10586_45546# 0.003919f
C27853 a_17730_32519# C10_N_btm 7.64e-19
C27854 a_n1991_42858# a_n4318_38216# 4.7e-19
C27855 a_n1853_43023# a_n2104_42282# 2.35e-20
C27856 a_10341_42308# a_12800_43218# 5.31e-21
C27857 a_12089_42308# a_11554_42852# 8.72e-21
C27858 a_10796_42968# a_11136_42852# 0.027606f
C27859 a_3626_43646# a_20107_42308# 0.001705f
C27860 a_14579_43548# a_14456_42282# 5.92e-19
C27861 a_10341_43396# a_5742_30871# 3.28e-19
C27862 a_n4318_39304# a_n4334_39392# 0.081919f
C27863 a_22485_44484# VDD 0.258874f
C27864 a_19237_31679# C8_N_btm 1.71e-20
C27865 a_2982_43646# a_7174_31319# 0.081795f
C27866 a_20512_43084# RST_Z 4.49e-21
C27867 a_n2157_42858# a_n3674_38216# 3.67e-19
C27868 a_n2840_42826# a_n4318_37592# 2.65e-20
C27869 a_13887_32519# a_n784_42308# 0.00652f
C27870 a_8953_45546# a_9061_43230# 3.71e-19
C27871 a_4743_44484# a_n2661_42834# 9.88e-20
C27872 a_10227_46804# CAL_N 7.26e-19
C27873 a_20567_45036# a_20640_44752# 0.003077f
C27874 a_n2661_43370# a_n2840_43914# 0.008144f
C27875 a_11691_44458# a_17061_44484# 0.005038f
C27876 a_8953_45002# a_9672_43914# 0.00114f
C27877 a_2711_45572# a_16137_43396# 1.42e-19
C27878 a_20205_31679# a_14209_32519# 0.051418f
C27879 a_n452_47436# VDD 0.092189f
C27880 a_n699_43396# a_n2661_43922# 0.053529f
C27881 a_18911_45144# a_19279_43940# 3.2e-20
C27882 a_11827_44484# a_11967_42832# 0.095859f
C27883 a_18494_42460# a_20679_44626# 1.25e-20
C27884 a_n1741_47186# CLK_DATA 8.62e-20
C27885 a_10057_43914# a_9313_44734# 0.139382f
C27886 a_n1920_47178# DATA[0] 7.82e-20
C27887 a_n2109_47186# DATA[1] 0.049689f
C27888 a_7499_43078# a_9145_43396# 0.040441f
C27889 a_5204_45822# a_5066_45546# 0.402457f
C27890 a_3483_46348# a_8034_45724# 1.49e-19
C27891 a_n881_46662# a_n745_45366# 0.152998f
C27892 a_4883_46098# a_6171_45002# 0.020043f
C27893 a_10227_46804# a_11963_45334# 7.17e-21
C27894 a_11599_46634# a_15415_45028# 0.013635f
C27895 a_8953_45546# a_526_44458# 0.037032f
C27896 a_6755_46942# a_13163_45724# 6.64e-21
C27897 a_17339_46660# a_n357_42282# 1.31e-19
C27898 a_9313_45822# a_1423_45028# 1.31e-20
C27899 a_16697_47582# a_2437_43646# 1.94e-19
C27900 a_20916_46384# a_20623_45572# 0.006579f
C27901 a_765_45546# a_310_45028# 0.012232f
C27902 a_3090_45724# a_3775_45552# 0.001359f
C27903 a_8270_45546# a_9049_44484# 0.006099f
C27904 a_14275_46494# a_10809_44734# 6.38e-20
C27905 a_18189_46348# a_19335_46494# 1.11e-21
C27906 a_18819_46122# a_18985_46122# 0.749955f
C27907 a_564_42282# a_6123_31319# 2.22e-20
C27908 a_n784_42308# a_8515_42308# 1.56e-20
C27909 a_3318_42354# a_3823_42558# 1e-19
C27910 a_4190_30871# VDAC_P 0.044542f
C27911 a_16877_42852# a_15803_42450# 1.15e-19
C27912 a_961_42354# a_5932_42308# 4.31e-21
C27913 a_6755_46942# DATA[5] 2.62e-19
C27914 a_n1059_45260# a_685_42968# 0.103646f
C27915 a_13249_42308# a_13291_42460# 0.068754f
C27916 a_n2956_39304# a_n4315_30879# 0.024812f
C27917 a_n2661_43370# a_9803_43646# 6.41e-22
C27918 a_n2661_42834# a_9248_44260# 1.02e-20
C27919 a_n699_43396# a_n447_43370# 0.040315f
C27920 a_4223_44672# a_n97_42460# 1.53e-19
C27921 a_n1761_44111# a_895_43940# 7.07e-21
C27922 a_10554_47026# CLK 0.014924f
C27923 a_n443_42852# a_1755_42282# 0.055323f
C27924 a_n755_45592# a_3905_42558# 4.35e-20
C27925 a_9313_44734# a_14021_43940# 0.014591f
C27926 a_8654_47026# VDD 4.6e-19
C27927 a_n967_45348# a_n1379_43218# 3.56e-19
C27928 a_3316_45546# a_3503_45724# 0.024901f
C27929 a_310_45028# a_509_45822# 0.039722f
C27930 a_n1099_45572# a_n443_42852# 0.026572f
C27931 a_2107_46812# a_9838_44484# 5.07e-20
C27932 a_10586_45546# a_11525_45546# 0.115475f
C27933 a_n2661_45546# a_603_45572# 8.65e-19
C27934 a_768_44030# a_5891_43370# 0.050862f
C27935 a_13059_46348# a_14537_43396# 0.30244f
C27936 a_n2497_47436# a_n1644_44306# 0.008707f
C27937 a_584_46384# a_453_43940# 0.125447f
C27938 a_n1991_46122# a_n1059_45260# 3.7e-20
C27939 a_n1853_46287# a_n913_45002# 1.34e-20
C27940 a_12465_44636# a_13940_44484# 1.26e-19
C27941 a_16327_47482# a_20362_44736# 0.213851f
C27942 a_n1151_42308# a_n984_44318# 0.009157f
C27943 a_376_46348# a_n2661_45010# 7.98e-23
C27944 a_22591_46660# a_413_45260# 1.37e-20
C27945 a_12861_44030# a_18681_44484# 1.24e-19
C27946 a_2324_44458# a_14033_45572# 6.09e-19
C27947 a_5066_45546# a_8697_45822# 0.033513f
C27948 a_8049_45260# a_13163_45724# 0.008063f
C27949 a_n4064_40160# a_n4209_39304# 0.04848f
C27950 a_n784_42308# EN_VIN_BSTR_N 0.051272f
C27951 a_n971_45724# a_6545_47178# 0.295443f
C27952 a_327_47204# a_n443_46116# 1.72e-19
C27953 a_2553_47502# a_n1151_42308# 0.007448f
C27954 a_2952_47436# a_3160_47472# 0.192116f
C27955 a_n1741_47186# a_6575_47204# 0.075265f
C27956 a_2063_45854# a_3381_47502# 1.06e-19
C27957 a_584_46384# a_3785_47178# 1.58e-20
C27958 a_n2946_39866# a_n4064_39616# 0.053228f
C27959 a_n3420_39616# a_n2302_39866# 1.28e-19
C27960 a_14097_32519# C1_N_btm 5.88e-20
C27961 a_16877_42852# VDD 0.192454f
C27962 a_n4315_30879# a_n3565_39304# 0.048127f
C27963 a_n1630_35242# a_n923_35174# 0.029967f
C27964 a_7640_43914# a_7871_42858# 3.94e-21
C27965 a_14539_43914# a_16414_43172# 2.71e-20
C27966 a_n2293_43922# a_n3674_39304# 1.03e-19
C27967 a_n2661_42834# a_n1736_43218# 5.14e-19
C27968 en_comp a_13575_42558# 4.34e-21
C27969 a_20692_30879# a_18194_35068# 1.16e-19
C27970 a_n356_44636# a_10922_42852# 2.27e-20
C27971 a_1307_43914# a_2351_42308# 0.00376f
C27972 a_n1059_45260# a_14113_42308# 4.15e-19
C27973 a_n2017_45002# a_15051_42282# 0.006558f
C27974 a_10037_46155# VDD 0.001395f
C27975 a_15493_43940# a_n97_42460# 0.009021f
C27976 a_14021_43940# a_20974_43370# 0.893848f
C27977 a_5891_43370# a_5755_42852# 0.160849f
C27978 a_18597_46090# a_3626_43646# 1.01e-19
C27979 a_12549_44172# a_19478_44056# 2.21e-20
C27980 a_n2293_45546# a_2232_45348# 0.004093f
C27981 a_5263_45724# a_5147_45002# 5.54e-20
C27982 a_11415_45002# a_13857_44734# 1.47e-20
C27983 a_15765_45572# a_16211_45572# 2.28e-19
C27984 a_n1613_43370# a_n2129_43609# 0.44294f
C27985 a_n1099_45572# a_375_42282# 8.14e-19
C27986 a_n357_42282# a_1307_43914# 0.044512f
C27987 a_n2956_39304# a_n4318_40392# 0.023379f
C27988 a_n2661_45546# a_2903_45348# 4.28e-19
C27989 a_7499_43078# a_n1059_45260# 0.277353f
C27990 a_17339_46660# a_18588_44850# 0.00201f
C27991 a_16333_45814# a_16842_45938# 2.6e-19
C27992 a_12741_44636# a_n2293_43922# 0.114756f
C27993 a_2711_45572# a_5691_45260# 0.004189f
C27994 a_n863_45724# a_1145_45348# 4.99e-20
C27995 a_2324_44458# a_6298_44484# 0.315008f
C27996 a_10903_43370# a_12607_44458# 0.004073f
C27997 a_n1435_47204# a_10249_46116# 7.87e-20
C27998 a_13381_47204# a_6755_46942# 9.89e-20
C27999 a_n4209_37414# C8_P_btm 1.65e-20
C28000 a_11599_46634# a_9863_46634# 3.12e-21
C28001 a_7754_40130# RST_Z 0.022036f
C28002 a_19321_45002# a_20843_47204# 1.68e-20
C28003 a_13747_46662# a_20916_46384# 2.31e-20
C28004 a_2747_46873# a_2959_46660# 0.010672f
C28005 CAL_N CAL_P 5.91728f
C28006 a_22521_40055# a_22821_38993# 0.131339f
C28007 a_22459_39145# a_22545_38993# 0.121283f
C28008 a_22780_40081# a_22521_39511# 1.39e-19
C28009 a_4883_46098# a_4955_46873# 0.09516f
C28010 a_n4209_38216# VREF_GND 0.001997f
C28011 a_n3565_37414# C10_P_btm 1.19e-19
C28012 a_n1613_43370# a_288_46660# 0.01808f
C28013 a_6151_47436# a_8189_46660# 0.001903f
C28014 a_584_46384# a_3090_45724# 0.001068f
C28015 a_7903_47542# a_8035_47026# 9.4e-20
C28016 a_n1151_42308# a_12251_46660# 0.00985f
C28017 a_12549_44172# a_n743_46660# 0.03191f
C28018 a_14021_43940# a_18599_43230# 5.88e-20
C28019 a_9313_44734# a_15764_42576# 3.58e-20
C28020 a_n2293_43922# a_5742_30871# 0.098838f
C28021 a_n356_44636# a_17531_42308# 0.030778f
C28022 a_2982_43646# a_21487_43396# 0.169809f
C28023 a_2437_43646# CLK 0.101524f
C28024 a_n2065_43946# a_n1736_42282# 3.49e-22
C28025 a_n1761_44111# a_n3674_38216# 5.92e-21
C28026 a_n2472_45002# VDD 0.217954f
C28027 a_8685_43396# a_16547_43609# 7.59e-20
C28028 a_3357_43084# DATA[4] 0.035981f
C28029 a_10341_43396# a_10849_43646# 1.08e-20
C28030 a_3626_43646# a_743_42282# 0.147999f
C28031 a_104_43370# a_n13_43084# 7.16e-19
C28032 a_n2293_46634# a_8037_42858# 1.56e-20
C28033 a_n357_42282# a_18579_44172# 2.1e-19
C28034 a_526_44458# a_9028_43914# 3.93e-21
C28035 a_20205_31679# a_17730_32519# 0.051307f
C28036 a_12549_44172# a_17701_42308# 3.43e-21
C28037 a_12741_44636# a_n97_42460# 3.68e-21
C28038 a_2680_45002# a_2809_45028# 0.062574f
C28039 a_20623_45572# a_21101_45002# 0.00299f
C28040 a_10227_46804# a_10553_43218# 0.001965f
C28041 a_n913_45002# a_n2661_43370# 0.031604f
C28042 a_10180_45724# a_9313_44734# 6.72e-20
C28043 a_5147_45002# a_5837_45348# 2.22e-19
C28044 a_5111_44636# a_5365_45348# 0.001271f
C28045 a_4927_45028# a_5105_45348# 0.007617f
C28046 a_7705_45326# a_1423_45028# 2.06e-22
C28047 a_11963_45334# a_1307_43914# 1.89e-20
C28048 a_13556_45296# a_14537_43396# 0.590856f
C28049 a_13777_45326# a_14180_45002# 0.002746f
C28050 a_9482_43914# a_14797_45144# 0.003056f
C28051 a_14976_45028# a_14205_43396# 4.75e-21
C28052 a_3090_45724# a_15095_43370# 0.00771f
C28053 a_15227_44166# a_9145_43396# 0.001689f
C28054 a_n2288_47178# a_n2293_45546# 5.3e-21
C28055 a_n2497_47436# a_n1079_45724# 5.93e-19
C28056 a_5807_45002# a_7920_46348# 3.4e-20
C28057 a_11309_47204# a_11387_46155# 0.061891f
C28058 a_12991_46634# a_13607_46688# 0.002207f
C28059 a_n743_46660# a_1208_46090# 0.045297f
C28060 a_n133_46660# a_472_46348# 6.87e-19
C28061 a_n2438_43548# a_805_46414# 2.09e-19
C28062 a_n2293_46634# a_167_45260# 0.087596f
C28063 a_21588_30879# a_4185_45028# 2.74e-19
C28064 a_n881_46662# a_14275_46494# 0.004854f
C28065 a_22959_47212# a_10809_44734# 0.005622f
C28066 a_5894_47026# a_765_45546# 1.39e-19
C28067 a_4915_47217# a_14371_46494# 0.001038f
C28068 a_n1151_42308# a_13259_45724# 5.41e-19
C28069 a_n1925_46634# a_1138_42852# 5.27e-19
C28070 SMPL_ON_P a_n2810_45572# 0.039568f
C28071 a_12549_44172# a_11189_46129# 3.08e-20
C28072 a_768_44030# a_9290_44172# 0.189655f
C28073 a_171_46873# a_376_46348# 0.080253f
C28074 a_6031_43396# a_5379_42460# 1.01e-19
C28075 a_9241_44734# VDD 0.003445f
C28076 a_16243_43396# a_16245_42852# 5.04e-20
C28077 a_15743_43084# a_15785_43172# 3.98e-19
C28078 a_16137_43396# a_16877_42852# 0.010276f
C28079 a_n1076_43230# a_n914_42852# 0.006453f
C28080 a_10991_42826# a_12089_42308# 3.42e-21
C28081 a_10796_42968# a_12545_42858# 0.002859f
C28082 a_2982_43646# a_5932_42308# 0.073161f
C28083 a_3626_43646# a_5755_42308# 0.003368f
C28084 a_n97_42460# a_5742_30871# 0.259664f
C28085 a_3483_46348# a_13635_43156# 1.81e-20
C28086 a_4185_45028# a_13113_42826# 3.91e-21
C28087 a_16375_45002# a_10341_43396# 1.23e-20
C28088 w_11334_34010# VDAC_N 0.049022f
C28089 a_11691_44458# a_18248_44752# 0.040333f
C28090 a_n357_42282# a_9396_43370# 1.13e-19
C28091 a_n913_45002# a_2998_44172# 1.35e-20
C28092 a_n2661_44458# a_9838_44484# 0.006567f
C28093 a_11827_44484# a_18989_43940# 0.054716f
C28094 a_n2293_42834# a_n2293_43922# 0.031735f
C28095 a_949_44458# a_2779_44458# 5.8e-19
C28096 a_413_45260# a_175_44278# 1.05e-19
C28097 a_16147_45260# a_18079_43940# 2.34e-19
C28098 a_8199_44636# a_9127_43156# 0.01079f
C28099 a_8016_46348# a_10083_42826# 1.33e-19
C28100 a_8953_45546# a_8605_42826# 3.03e-19
C28101 a_n2017_45002# a_3905_42865# 5.53e-19
C28102 a_18184_42460# a_n356_44636# 0.05602f
C28103 a_n452_44636# a_n699_43396# 1.94e-21
C28104 a_13507_46334# a_19431_45546# 2.47e-20
C28105 a_n743_46660# a_11525_45546# 1.75e-21
C28106 a_4646_46812# a_2711_45572# 0.053113f
C28107 a_3483_46348# a_8016_46348# 0.019798f
C28108 a_n237_47217# a_5147_45002# 5.93e-20
C28109 a_18280_46660# a_10809_44734# 0.002977f
C28110 a_13717_47436# a_2437_43646# 0.085485f
C28111 a_12861_44030# a_21513_45002# 2.48e-20
C28112 a_2107_46812# a_8568_45546# 2.03e-20
C28113 a_2952_47436# a_413_45260# 0.026401f
C28114 a_n1151_42308# a_n467_45028# 0.406349f
C28115 a_4883_46098# a_18909_45814# 1.42e-21
C28116 a_16327_47482# a_21363_45546# 0.276554f
C28117 a_11459_47204# a_3357_43084# 5.7e-19
C28118 a_n881_46662# a_15765_45572# 0.58719f
C28119 a_584_46384# a_2274_45254# 3.31e-21
C28120 a_12549_44172# a_11136_45572# 1.78e-21
C28121 a_5068_46348# a_5204_45822# 0.20685f
C28122 a_12741_44636# a_17957_46116# 9.01e-21
C28123 a_3699_46634# a_3775_45552# 5.03e-19
C28124 a_5342_30871# a_13921_42308# 8.71e-20
C28125 a_17538_32519# C10_N_btm 2.16e-19
C28126 a_n3674_39304# a_n3420_39616# 0.152699f
C28127 a_3080_42308# EN_VIN_BSTR_N 0.04304f
C28128 a_14401_32519# VDD 0.562673f
C28129 a_21381_43940# RST_Z 3.55e-21
C28130 a_5837_42852# a_5932_42308# 4.77e-19
C28131 a_22612_30879# VREF 1.73216f
C28132 a_n2661_46634# CLK 0.032279f
C28133 a_n357_42282# a_13003_42852# 0.002208f
C28134 a_9290_44172# a_10149_42308# 0.001223f
C28135 a_1823_45246# a_7174_31319# 1.97e-20
C28136 a_n2293_42834# a_n97_42460# 0.17628f
C28137 a_21588_30879# VREF_GND 0.083908f
C28138 a_19615_44636# a_19279_43940# 1.59e-19
C28139 a_18588_44850# a_18579_44172# 9.38e-20
C28140 a_11967_42832# a_18005_44484# 2.11e-19
C28141 a_10193_42453# a_18817_42826# 0.002321f
C28142 a_n443_42852# a_9306_43218# 3.58e-20
C28143 a_33_46660# VDD 0.272723f
C28144 a_5891_43370# a_7845_44172# 0.119969f
C28145 a_13249_42308# a_13460_43230# 0.014543f
C28146 a_11823_42460# a_15567_42826# 3.26e-19
C28147 a_20362_44736# a_20835_44721# 7.99e-20
C28148 a_n2661_42834# a_1414_42308# 0.081864f
C28149 a_n2661_43922# a_1467_44172# 0.002845f
C28150 a_20640_44752# a_20679_44626# 0.582607f
C28151 a_n2661_43370# a_n4318_39304# 0.00535f
C28152 a_n1059_45260# a_15781_43660# 4.06e-20
C28153 a_18114_32519# a_14021_43940# 2.66e-19
C28154 a_n1925_46634# DATA[1] 4.06e-21
C28155 a_11387_46155# a_10490_45724# 1.07e-20
C28156 a_11189_46129# a_11525_45546# 0.085926f
C28157 a_11133_46155# a_11322_45546# 0.001455f
C28158 a_12005_46116# a_10193_42453# 0.016165f
C28159 a_10903_43370# a_8746_45002# 1.84e-19
C28160 a_19321_45002# a_20567_45036# 0.205038f
C28161 a_5807_45002# a_11827_44484# 0.022597f
C28162 a_13747_46662# a_21101_45002# 0.081818f
C28163 a_14035_46660# a_2437_43646# 1.31e-19
C28164 a_3877_44458# a_5105_45348# 9.23e-22
C28165 a_10249_46116# a_10775_45002# 1.35e-22
C28166 a_6755_46942# a_8953_45002# 6.77e-20
C28167 a_15227_44166# a_n1059_45260# 0.099892f
C28168 a_n1613_43370# a_n2129_44697# 0.026334f
C28169 a_12991_46634# a_413_45260# 4.46e-20
C28170 a_n1151_42308# a_n2661_43922# 0.056653f
C28171 a_2107_46812# a_n2661_43370# 0.02614f
C28172 a_9290_44172# a_11652_45724# 0.020364f
C28173 a_10554_47026# a_10951_45334# 2.81e-22
C28174 a_526_44458# a_1609_45822# 3.1e-20
C28175 a_n1925_42282# a_n443_42852# 0.02261f
C28176 a_6945_45028# a_6511_45714# 0.028815f
C28177 a_17303_42282# a_18907_42674# 1.62e-19
C28178 a_18249_42858# RST_Z 6.28e-21
C28179 a_18817_42826# VDD 0.204624f
C28180 a_n2293_42834# a_3935_43218# 9.69e-20
C28181 a_n2956_37592# a_n3674_38216# 0.023192f
C28182 a_n913_45002# COMP_P 1.4e-20
C28183 a_18248_44752# a_4190_30871# 2.51e-20
C28184 a_11341_43940# a_22223_43948# 0.175191f
C28185 a_21115_43940# a_15493_43940# 0.0516f
C28186 a_14673_44172# a_8685_43396# 9.41e-20
C28187 a_10193_42453# a_21421_42336# 1.05e-20
C28188 en_comp a_n2104_42282# 0.002636f
C28189 a_n2017_45002# a_n961_42308# 0.012655f
C28190 a_n967_45348# a_n4318_38216# 3e-20
C28191 a_n2810_45028# a_n1736_42282# 9.69e-21
C28192 a_12005_46116# VDD 0.518463f
C28193 a_17737_43940# a_14021_43940# 2.4e-20
C28194 a_n2661_42282# a_5829_43940# 0.002389f
C28195 a_1115_44172# a_n97_42460# 1.16e-19
C28196 a_8199_44636# CLK 0.231904f
C28197 a_n1925_42282# a_375_42282# 2.07e-19
C28198 a_11525_45546# a_11136_45572# 1.53e-19
C28199 a_n2312_38680# a_n3674_39768# 0.023176f
C28200 a_2711_45572# a_18479_45785# 0.032371f
C28201 a_n1151_42308# a_n447_43370# 1.85e-19
C28202 SMPL_ON_P a_n1557_42282# 2.98e-20
C28203 a_17339_46660# a_18443_44721# 0.006967f
C28204 a_12465_44636# a_14021_43940# 0.015806f
C28205 a_768_44030# a_10807_43548# 0.001051f
C28206 a_n863_45724# a_3357_43084# 0.003254f
C28207 a_n2840_45546# a_n2840_45002# 0.026152f
C28208 a_19692_46634# a_9313_44734# 3.49e-20
C28209 a_10490_45724# a_11778_45572# 0.004273f
C28210 a_8049_45260# a_8953_45002# 7.24e-19
C28211 a_n1741_47186# a_5385_46902# 1.59e-20
C28212 a_n2109_47186# a_5907_46634# 0.001384f
C28213 a_n1151_42308# a_1799_45572# 2.59e-19
C28214 a_6575_47204# a_n743_46660# 5.55e-20
C28215 a_n4209_39304# C10_P_btm 4.87e-19
C28216 a_4915_47217# a_2107_46812# 6.45e-20
C28217 a_3754_38802# VDAC_Ni 0.301032f
C28218 a_7754_39300# a_8530_39574# 3.17e-19
C28219 a_2113_38308# a_4338_37500# 1.76e-20
C28220 a_13507_46334# a_12891_46348# 0.076674f
C28221 a_16588_47582# a_5807_45002# 0.040789f
C28222 a_10227_46804# a_16942_47570# 0.00186f
C28223 a_n971_45724# a_3877_44458# 0.927248f
C28224 a_2063_45854# a_2959_46660# 2.88e-19
C28225 a_2952_47436# a_2609_46660# 0.006778f
C28226 a_2905_45572# a_2443_46660# 0.026052f
C28227 a_n3420_37984# VDAC_P 3.33e-19
C28228 a_n2312_40392# a_n1613_43370# 4.82e-21
C28229 a_n4064_39616# C1_P_btm 3.84e-20
C28230 a_6197_43396# a_6765_43638# 0.17072f
C28231 a_2982_43646# a_4181_43396# 1.27e-20
C28232 a_11967_42832# a_13569_43230# 8.29e-19
C28233 a_18494_42460# a_18057_42282# 0.085802f
C28234 a_18184_42460# a_18727_42674# 0.044914f
C28235 a_14033_45822# VDD 0.195067f
C28236 a_14021_43940# a_13887_32519# 0.020984f
C28237 a_8333_44056# a_8387_43230# 7.4e-22
C28238 a_n356_44636# a_2903_42308# 2.77e-19
C28239 a_n2661_42834# a_n3674_38680# 0.03399f
C28240 a_n2810_45028# a_n4209_37414# 0.09606f
C28241 a_5883_43914# a_8685_42308# 1.31e-20
C28242 a_6293_42852# a_6547_43396# 3.12e-19
C28243 a_6031_43396# a_7287_43370# 0.042271f
C28244 a_1414_42308# a_n2293_42282# 1.08e-20
C28245 a_19692_46634# a_20974_43370# 0.012779f
C28246 a_13259_45724# a_13857_44734# 0.03212f
C28247 a_8696_44636# a_8560_45348# 6.21e-19
C28248 a_20692_30879# a_9313_44734# 1.31e-20
C28249 a_n2017_45002# a_5147_45002# 4.93e-22
C28250 a_10227_46804# a_8952_43230# 7.54e-21
C28251 a_12549_44172# a_4361_42308# 8.96e-19
C28252 a_11415_45002# a_15493_43940# 1.15e-19
C28253 a_6194_45824# a_5883_43914# 1.36e-19
C28254 a_13527_45546# a_11691_44458# 2.01e-21
C28255 a_2324_44458# a_2479_44172# 0.010173f
C28256 a_n467_45028# a_327_44734# 6.38e-20
C28257 a_n2661_45010# a_3232_43370# 3.31e-19
C28258 a_13661_43548# a_16823_43084# 7.25e-19
C28259 a_4185_45028# a_n2661_42282# 0.833759f
C28260 a_8568_45546# a_n2661_44458# 4.32e-21
C28261 a_2711_45572# a_10057_43914# 7.42e-20
C28262 a_6667_45809# a_6298_44484# 0.001371f
C28263 a_3877_44458# a_8023_46660# 1.47e-20
C28264 a_6151_47436# a_13351_46090# 4.87e-21
C28265 a_5807_45002# a_14447_46660# 8.93e-19
C28266 a_n2312_40392# a_n2293_46098# 7.25e-19
C28267 a_n2312_39304# a_n2472_46090# 0.006797f
C28268 a_8145_46902# a_7927_46660# 0.209641f
C28269 a_7577_46660# a_8667_46634# 0.041879f
C28270 a_6540_46812# a_6682_46987# 0.005572f
C28271 a_7715_46873# a_8492_46660# 5.47e-21
C28272 a_9313_45822# a_9569_46155# 0.019679f
C28273 a_n1435_47204# a_5937_45572# 1.19e-20
C28274 a_7411_46660# a_9863_46634# 2.84e-21
C28275 a_4915_47217# a_14493_46090# 1.95e-19
C28276 a_n2433_43396# a_n4318_37592# 2.5e-20
C28277 a_15682_43940# a_15803_42450# 4.66e-19
C28278 a_743_42282# a_8037_42858# 5.74e-20
C28279 a_16547_43609# a_17333_42852# 2.75e-20
C28280 a_16137_43396# a_18817_42826# 8.32e-19
C28281 a_19721_31679# C10_N_btm 2.25e-20
C28282 a_n1076_43230# a_n13_43084# 3.14e-19
C28283 a_n1641_43230# a_n4318_38680# 4.97e-20
C28284 a_11341_43940# a_11323_42473# 2.29e-19
C28285 a_14401_32519# a_n784_42308# 0.003982f
C28286 a_n2129_43609# a_n1736_42282# 1.65e-20
C28287 a_20205_45028# VDD 0.005516f
C28288 a_n1991_42858# a_n1545_43230# 2.28e-19
C28289 a_n2157_42858# a_n967_43230# 2.56e-19
C28290 a_n1853_43023# a_n1379_43218# 0.002143f
C28291 a_4361_42308# a_5111_42852# 5.5e-20
C28292 a_n2661_43370# a_n2661_44458# 1.0558f
C28293 a_3232_43370# a_8855_44734# 0.001723f
C28294 a_6709_45028# a_7640_43914# 8.38e-19
C28295 a_16922_45042# a_11691_44458# 0.428229f
C28296 a_19778_44110# a_21005_45260# 0.135527f
C28297 a_16405_45348# a_16237_45028# 8.13e-19
C28298 a_18184_42460# a_20567_45036# 9.9e-21
C28299 a_18315_45260# a_11827_44484# 9.63e-19
C28300 a_11525_45546# a_11750_44172# 1.43e-21
C28301 a_11322_45546# a_12429_44172# 5.73e-21
C28302 a_20623_45572# a_20766_44850# 1.55e-20
C28303 a_21188_45572# a_20679_44626# 3.17e-20
C28304 a_2711_45572# a_14021_43940# 0.029672f
C28305 a_20205_31679# a_17538_32519# 0.051233f
C28306 a_16327_47482# a_17303_42282# 4.29e-19
C28307 a_4185_45028# a_16823_43084# 6.8e-21
C28308 a_10227_46804# a_15521_42308# 0.001965f
C28309 a_10193_42453# a_15682_43940# 0.003859f
C28310 a_327_44734# a_n2661_43922# 0.005571f
C28311 a_3537_45260# a_3363_44484# 9.26e-20
C28312 a_n2293_42834# a_742_44458# 0.039916f
C28313 a_n1613_43370# a_8791_42308# 6.28e-21
C28314 a_3090_45724# a_17583_46090# 0.003153f
C28315 a_10933_46660# a_9290_44172# 2.81e-19
C28316 a_765_45546# a_2804_46116# 1.28e-20
C28317 a_22591_46660# a_20820_30879# 0.166885f
C28318 a_11415_45002# a_12741_44636# 1.07921f
C28319 a_20202_43084# a_22959_46660# 2.07e-19
C28320 a_4883_46098# a_8746_45002# 0.032616f
C28321 a_10227_46804# a_13249_42308# 0.064815f
C28322 a_n2661_46634# a_n1099_45572# 5.05e-20
C28323 a_n743_46660# a_n2661_45546# 0.013544f
C28324 a_n2438_43548# a_n2810_45572# 4.17e-19
C28325 a_n881_46662# a_6194_45824# 0.063172f
C28326 a_n1613_43370# a_6472_45840# 0.017909f
C28327 a_n2293_46634# a_n863_45724# 0.157683f
C28328 a_9804_47204# a_2711_45572# 2.39e-19
C28329 a_15368_46634# a_2324_44458# 0.00404f
C28330 a_15682_43940# VDD 1.22657f
C28331 a_5649_42852# a_15959_42545# 1.03e-19
C28332 a_17021_43396# a_4958_30871# 5.45e-20
C28333 a_5534_30871# a_1606_42308# 0.030581f
C28334 a_4361_42308# a_9885_42308# 0.001144f
C28335 a_15743_43084# a_19647_42308# 7.14e-19
C28336 a_19268_43646# a_19511_42282# 1.08e-19
C28337 a_1823_45246# a_5932_42308# 8.68e-21
C28338 a_n967_45348# a_n1655_43396# 2.02e-19
C28339 a_18443_44721# a_18579_44172# 5.4e-19
C28340 a_18374_44850# a_18245_44484# 4.2e-19
C28341 a_18248_44752# a_18753_44484# 2.28e-19
C28342 a_742_44458# a_1115_44172# 0.001155f
C28343 a_13507_46334# SINGLE_ENDED 0.111959f
C28344 a_22612_30879# a_22521_40599# 9.6e-20
C28345 a_21588_30879# a_22469_40625# 6.62e-20
C28346 a_n37_45144# a_104_43370# 2.79e-21
C28347 a_413_45260# a_n97_42460# 1.07e-21
C28348 a_n699_43396# a_n809_44244# 1.25e-19
C28349 a_n913_45002# a_1568_43370# 0.098659f
C28350 a_n1059_45260# a_1756_43548# 6.3e-22
C28351 a_n2017_45002# a_4093_43548# 5.54e-21
C28352 a_n2661_44458# a_2998_44172# 2.23e-19
C28353 a_21811_47423# VDD 0.201359f
C28354 a_n357_42282# a_13635_43156# 0.008746f
C28355 a_1307_43914# a_5025_43940# 0.003108f
C28356 a_4883_46098# RST_Z 1.25e-19
C28357 a_21496_47436# START 3e-20
C28358 a_n443_42852# a_8387_43230# 0.006907f
C28359 a_3357_43084# a_3540_43646# 0.001122f
C28360 a_n2661_46098# a_413_45260# 1.23e-20
C28361 a_n1151_42308# a_n452_44636# 0.238824f
C28362 a_15227_44166# a_15599_45572# 4.09e-21
C28363 a_3090_45724# a_8696_44636# 0.038457f
C28364 a_n881_46662# a_6517_45366# 5.23e-19
C28365 a_11453_44696# a_n2661_43370# 0.002123f
C28366 a_16327_47482# a_19778_44110# 0.037655f
C28367 a_n2661_46634# a_10951_45334# 9.5e-21
C28368 a_n743_46660# a_5205_44484# 2.07e-20
C28369 a_167_45260# a_2277_45546# 0.214157f
C28370 a_2107_46812# a_4574_45260# 3.63e-20
C28371 a_18479_47436# a_16922_45042# 6.1e-20
C28372 a_17957_46116# a_16375_45002# 0.017118f
C28373 a_18189_46348# a_19240_46482# 1.71e-21
C28374 a_8016_46348# a_n357_42282# 3.18e-20
C28375 a_n1925_46634# a_7229_43940# 3.86e-21
C28376 a_n2293_46098# a_6472_45840# 6.84e-21
C28377 a_765_45546# a_13904_45546# 7.77e-22
C28378 a_15368_46634# a_16855_45546# 6.26e-21
C28379 a_13661_43548# a_15415_45028# 0.133591f
C28380 a_10533_42308# a_5742_30871# 0.020913f
C28381 a_10723_42308# a_11323_42473# 0.008191f
C28382 a_5649_42852# RST_Z 6.96e-19
C28383 a_n4318_37592# a_n4064_40160# 0.079413f
C28384 a_22223_43396# VDD 0.279195f
C28385 a_17364_32525# C7_N_btm 0.072179f
C28386 a_1184_42692# a_7174_31319# 6.06e-21
C28387 a_5534_30871# a_8912_37509# 3.98e-19
C28388 a_22485_44484# a_14021_43940# 1.69e-19
C28389 a_n356_44636# a_6293_42852# 2.26e-20
C28390 a_22000_46634# VDD 0.257047f
C28391 a_21188_46660# RST_Z 1.88e-21
C28392 a_16922_45042# a_4190_30871# 0.353708f
C28393 a_20623_46660# SINGLE_ENDED 2.87e-20
C28394 a_11691_44458# a_15743_43084# 3.24e-19
C28395 a_19113_45348# a_19268_43646# 1.84e-21
C28396 a_n2293_42834# a_n901_43156# 0.021108f
C28397 a_1307_43914# a_8952_43230# 1.54e-20
C28398 a_765_45546# CLK 0.0309f
C28399 a_9838_44484# a_9145_43396# 2.26e-22
C28400 a_20205_31679# a_22465_38105# 3.95e-19
C28401 a_10193_42453# a_5934_30871# 6.18e-20
C28402 a_2711_45572# a_15764_42576# 1.23e-20
C28403 a_1423_45028# a_7871_42858# 3.55e-21
C28404 a_n2661_42834# a_n1190_43762# 1.25e-19
C28405 a_n2293_43922# a_n2012_43396# 0.011692f
C28406 a_2324_44458# a_2680_45002# 9e-20
C28407 a_19692_46634# a_18114_32519# 5.21e-19
C28408 a_10903_43370# a_3232_43370# 0.114259f
C28409 a_n2956_39304# a_n2017_45002# 9.09e-22
C28410 a_12549_44172# a_20397_44484# 1.48e-19
C28411 a_n1925_42282# a_2437_43646# 2.49e-20
C28412 a_n1613_43370# a_n2472_43914# 1.2e-19
C28413 a_2711_45572# a_10180_45724# 0.01318f
C28414 a_6472_45840# a_7230_45938# 0.05936f
C28415 a_6511_45714# a_6812_45938# 9.73e-19
C28416 a_6598_45938# a_6428_45938# 2.6e-19
C28417 a_167_45260# a_626_44172# 0.04273f
C28418 a_1823_45246# a_1423_45028# 0.024089f
C28419 a_5937_45572# a_10775_45002# 1.83e-20
C28420 a_19321_45002# a_20679_44626# 0.023087f
C28421 a_8953_45546# a_8953_45002# 0.023516f
C28422 a_13661_43548# a_19279_43940# 6.72e-19
C28423 a_13747_46662# a_20766_44850# 1.67e-19
C28424 a_10809_44734# a_n913_45002# 0.0025f
C28425 a_8199_44636# a_10951_45334# 0.237774f
C28426 a_1736_39043# a_2113_38308# 0.088667f
C28427 a_n3565_38502# a_n3690_38304# 7.97e-20
C28428 a_n3690_38528# a_n3565_38216# 7.97e-20
C28429 a_n2946_38778# a_n4209_38216# 5.32e-20
C28430 a_n3420_38528# a_n4334_38304# 0.014479f
C28431 a_n4209_38502# a_n2946_37984# 5.32e-20
C28432 a_n4064_38528# a_n3607_38528# 7.1e-19
C28433 a_n4064_40160# a_n4334_37440# 0.007725f
C28434 a_13258_32519# VDAC_N 4.18e-19
C28435 a_n2109_47186# a_768_44030# 2.81e-21
C28436 a_n1741_47186# a_12891_46348# 0.107238f
C28437 a_n971_45724# a_8128_46384# 0.041637f
C28438 a_n785_47204# a_n881_46662# 6.65e-20
C28439 a_327_47204# a_n1613_43370# 0.002699f
C28440 a_n1151_42308# a_2747_46873# 0.009962f
C28441 a_2952_47436# a_3094_47570# 0.007833f
C28442 a_2063_45854# a_2266_47243# 4.14e-19
C28443 a_5934_30871# VDD 0.431204f
C28444 a_n4315_30879# a_n3690_37440# 1.35e-19
C28445 a_15811_47375# a_16241_47178# 0.003645f
C28446 a_15507_47210# a_16327_47482# 0.425757f
C28447 a_11599_46634# a_16023_47582# 1.42e-20
C28448 a_12861_44030# a_10227_46804# 0.291378f
C28449 a_13717_47436# a_18143_47464# 3.4e-19
C28450 a_4915_47217# a_11453_44696# 0.026396f
C28451 a_5742_30871# C2_P_btm 0.030783f
C28452 a_14539_43914# a_17141_43172# 0.00164f
C28453 en_comp a_1736_39587# 8.86e-19
C28454 a_n1352_43396# a_n1190_43762# 0.006453f
C28455 a_n1917_43396# a_n1655_43396# 0.001705f
C28456 a_22223_43948# a_10341_43396# 0.002507f
C28457 a_15682_43940# a_16137_43396# 0.004591f
C28458 a_7542_44172# a_4361_42308# 2.2e-21
C28459 a_11967_42832# a_13113_42826# 0.021992f
C28460 a_17517_44484# a_17595_43084# 1.18e-21
C28461 a_18479_47436# a_15743_43084# 4.35e-20
C28462 a_3090_45724# a_20365_43914# 1.09e-19
C28463 a_20205_31679# a_19721_31679# 0.052217f
C28464 a_20692_30879# a_18114_32519# 0.051555f
C28465 a_15227_44166# a_18326_43940# 5.29e-20
C28466 a_20273_45572# a_21350_45938# 1.46e-19
C28467 a_13249_42308# a_1307_43914# 0.056917f
C28468 a_11682_45822# a_11963_45334# 2.91e-20
C28469 a_8049_45260# a_17767_44458# 9.2e-21
C28470 a_n2293_46634# a_3540_43646# 0.003694f
C28471 a_n2293_46098# a_n2472_43914# 5.06e-21
C28472 a_5907_45546# a_n2661_43370# 0.007276f
C28473 a_n1925_42282# a_4181_44734# 6.6e-19
C28474 a_n1151_42308# a_n1641_43230# 9.41e-19
C28475 C2_P_btm C0_dummy_P_btm 6.66125f
C28476 C3_P_btm C0_dummy_N_btm 2.71e-19
C28477 C7_P_btm C3_N_btm 6.36e-19
C28478 C5_P_btm C1_N_btm 1.59e-19
C28479 C4_P_btm C0_N_btm 1.4e-19
C28480 C1_P_btm C0_P_btm 10.8764f
C28481 a_1799_45572# a_3177_46902# 7.67e-21
C28482 a_n2661_46098# a_2609_46660# 6e-19
C28483 a_12861_44030# a_17339_46660# 1.25428f
C28484 a_13717_47436# a_765_45546# 0.009975f
C28485 a_4883_46098# a_10425_46660# 2.44e-19
C28486 a_n743_46660# a_5385_46902# 5.02e-22
C28487 a_2107_46812# a_2162_46660# 0.002508f
C28488 a_11530_34132# VDD 0.362839f
C28489 a_n2497_47436# a_1823_45246# 0.025359f
C28490 a_327_47204# a_n2293_46098# 8.71e-21
C28491 a_8128_46384# a_8023_46660# 8e-19
C28492 a_n815_47178# a_n1076_46494# 6.69e-19
C28493 a_n2109_47186# a_1176_45822# 1.41e-19
C28494 a_5807_45002# a_10150_46912# 0.007534f
C28495 a_n1925_46634# a_5907_46634# 0.010645f
C28496 a_15811_47375# a_16721_46634# 2.3e-19
C28497 a_15673_47210# a_16388_46812# 4.51e-19
C28498 a_10227_46804# a_14180_46812# 0.008201f
C28499 a_12465_44636# a_19692_46634# 6.79e-20
C28500 a_11453_44696# a_18834_46812# 0.010577f
C28501 a_16977_43638# a_4361_42308# 4.56e-21
C28502 a_9396_43370# a_8952_43230# 6.44e-19
C28503 a_3499_42826# a_3318_42354# 4.85e-19
C28504 a_18525_43370# a_743_42282# 5.58e-21
C28505 a_7281_43914# a_7227_42308# 1.21e-20
C28506 a_11967_42832# a_18214_42558# 8.49e-19
C28507 a_16243_43396# a_5649_42852# 8.11e-21
C28508 a_15743_43084# a_4190_30871# 0.290729f
C28509 a_2982_43646# a_15567_42826# 2.67e-20
C28510 a_8696_44636# a_14815_43914# 0.002482f
C28511 a_413_45260# a_742_44458# 0.001341f
C28512 a_327_44734# a_n452_44636# 5.28e-19
C28513 a_n2312_40392# a_n1736_42282# 4.5e-20
C28514 a_n2312_39304# a_n3674_38216# 0.023615f
C28515 a_13259_45724# a_15493_43940# 0.019228f
C28516 a_16751_45260# a_17023_45118# 0.13675f
C28517 a_8953_45546# a_3626_43646# 0.005746f
C28518 a_n357_42282# a_7584_44260# 7.22e-20
C28519 a_10193_42453# a_20512_43084# 0.086337f
C28520 a_n913_45002# a_5883_43914# 1.2e-19
C28521 a_17339_46660# a_19700_43370# 3.22e-19
C28522 a_19692_46634# a_13887_32519# 2.91e-19
C28523 a_6125_45348# a_n2661_43370# 8.72e-19
C28524 a_4574_45260# a_n2661_44458# 6.04e-19
C28525 a_3483_46348# a_8791_43396# 4.38e-23
C28526 a_13017_45260# a_11827_44484# 2.91e-21
C28527 a_22223_47212# a_20205_31679# 8.22e-20
C28528 a_14035_46660# a_765_45546# 9.28e-19
C28529 a_171_46873# a_n1379_46482# 8.94e-21
C28530 a_2107_46812# a_10809_44734# 1.51e-20
C28531 a_n1741_47186# a_11322_45546# 0.003846f
C28532 a_4915_47217# a_5907_45546# 4.1e-22
C28533 a_n237_47217# a_7499_43078# 4.22e-20
C28534 a_n443_46116# a_6194_45824# 8.96e-21
C28535 a_4791_45118# a_6472_45840# 0.025301f
C28536 a_19692_46634# a_20528_46660# 0.021985f
C28537 a_17609_46634# a_18280_46660# 0.094543f
C28538 a_11309_47204# a_11387_46482# 0.006175f
C28539 a_10428_46928# a_3483_46348# 3.44e-19
C28540 a_6545_47178# a_2711_45572# 8.4e-19
C28541 a_5257_43370# a_6419_46155# 0.186651f
C28542 a_n2661_46634# a_n1925_42282# 8.9e-20
C28543 a_4883_46098# a_21167_46155# 3.61e-19
C28544 a_17730_32519# C9_N_btm 0.215899f
C28545 a_4190_30871# a_1606_42308# 0.018892f
C28546 a_n1853_43023# a_n4318_38216# 8.05e-19
C28547 a_n2157_42858# a_n2104_42282# 0.011248f
C28548 a_10835_43094# a_11136_42852# 9.73e-19
C28549 a_12379_42858# a_11554_42852# 2.33e-21
C28550 a_3626_43646# a_13258_32519# 0.006214f
C28551 a_n4318_39304# a_n4209_39304# 0.135369f
C28552 a_2982_43646# a_20712_42282# 0.003556f
C28553 a_9145_43396# a_13657_42558# 4.78e-19
C28554 a_17364_32525# COMP_P 9.77e-21
C28555 a_19237_31679# C7_N_btm 1.43e-20
C28556 a_20512_43084# VDD 0.317257f
C28557 a_6171_45002# a_13483_43940# 2.43e-21
C28558 a_n443_42852# a_15743_43084# 0.034562f
C28559 a_21076_30879# a_14097_32519# 0.054945f
C28560 a_5343_44458# a_9159_44484# 2.67e-20
C28561 a_20567_45036# a_20362_44736# 6.75e-19
C28562 a_n2293_42834# a_n984_44318# 1.22e-19
C28563 a_11691_44458# a_16789_44484# 3.16e-19
C28564 a_8953_45002# a_9028_43914# 0.001179f
C28565 a_n815_47178# VDD 0.380339f
C28566 a_4223_44672# a_n2661_43922# 0.059715f
C28567 a_n699_43396# a_n2661_42834# 0.131393f
C28568 a_21359_45002# a_11967_42832# 1.28e-19
C28569 a_19778_44110# a_20835_44721# 8.16e-19
C28570 a_18184_42460# a_20679_44626# 7.45e-21
C28571 a_11827_44484# a_19006_44850# 0.002956f
C28572 a_18494_42460# a_20640_44752# 1.1e-19
C28573 a_n1920_47178# CLK_DATA 3.9e-19
C28574 a_n2109_47186# DATA[0] 0.08202f
C28575 a_10440_44484# a_9313_44734# 0.027369f
C28576 a_7499_43078# a_8423_43396# 4.14e-19
C28577 a_n2661_45546# a_4361_42308# 1.97e-21
C28578 a_20692_30879# a_13887_32519# 0.051577f
C28579 a_n863_45724# a_743_42282# 0.05133f
C28580 a_5164_46348# a_5066_45546# 0.096188f
C28581 a_5204_45822# a_5431_46482# 0.004982f
C28582 a_12861_44030# a_1307_43914# 0.038753f
C28583 a_n881_46662# a_n913_45002# 0.00874f
C28584 a_n1613_43370# a_n745_45366# 0.012092f
C28585 a_4883_46098# a_3232_43370# 0.017979f
C28586 a_10227_46804# a_11787_45002# 1.63e-21
C28587 a_5937_45572# a_526_44458# 7.57e-20
C28588 a_19692_46634# a_2711_45572# 4.14e-20
C28589 a_20916_46384# a_20841_45814# 1.18e-19
C28590 a_19321_45002# a_20528_45572# 7.43e-20
C28591 a_16285_47570# a_2437_43646# 7.17e-19
C28592 a_11415_45002# a_16375_45002# 0.080382f
C28593 a_12741_44636# a_13259_45724# 0.113445f
C28594 a_765_45546# a_n1099_45572# 7.06e-19
C28595 a_8270_45546# a_7499_43078# 0.063428f
C28596 a_6755_46942# a_12791_45546# 4.95e-22
C28597 a_15015_46420# a_6945_45028# 4.64e-20
C28598 a_n784_42308# a_5934_30871# 0.142087f
C28599 a_1755_42282# a_4921_42308# 0.002752f
C28600 a_16245_42852# a_15803_42450# 4.81e-19
C28601 a_1184_42692# a_5932_42308# 4.31e-21
C28602 a_10249_46116# DATA[5] 3.81e-19
C28603 a_6755_46942# DATA[4] 4.06e-21
C28604 a_n2017_45002# a_685_42968# 9.17e-20
C28605 a_n2661_43370# a_9145_43396# 1.28e-20
C28606 a_n699_43396# a_n1352_43396# 0.003121f
C28607 a_6969_46634# DATA[3] 6.68e-20
C28608 a_10623_46897# CLK 0.016177f
C28609 a_n443_42852# a_1606_42308# 0.003624f
C28610 a_n755_45592# a_3581_42558# 2.25e-19
C28611 a_175_44278# a_644_44056# 0.00101f
C28612 a_2779_44458# a_n97_42460# 1.5e-20
C28613 a_n967_45348# a_n1545_43230# 5.71e-19
C28614 a_3218_45724# a_3503_45724# 0.099872f
C28615 a_n1099_45572# a_509_45822# 0.026885f
C28616 a_380_45546# a_n443_42852# 0.030032f
C28617 a_2107_46812# a_5883_43914# 0.009818f
C28618 a_10586_45546# a_11322_45546# 0.220166f
C28619 a_8049_45260# a_12791_45546# 0.005799f
C28620 a_n2661_45546# a_509_45572# 4.21e-19
C28621 a_10809_44734# a_15903_45785# 2.74e-20
C28622 a_768_44030# a_8375_44464# 0.001943f
C28623 a_13059_46348# a_14180_45002# 0.073427f
C28624 a_n2497_47436# a_n3674_39768# 5.96e-20
C28625 a_n1853_46287# a_n1059_45260# 0.006746f
C28626 a_n1991_46122# a_n2017_45002# 5.3e-19
C28627 a_12465_44636# a_13296_44484# 1.43e-19
C28628 a_16327_47482# a_20159_44458# 0.270426f
C28629 a_n863_45724# a_2277_45546# 0.00198f
C28630 a_n743_46660# a_13076_44458# 9.1e-21
C28631 a_3090_45724# a_5009_45028# 0.008714f
C28632 a_n1151_42308# a_n809_44244# 0.02481f
C28633 a_584_46384# a_1414_42308# 0.321387f
C28634 a_n1076_46494# a_n2661_45010# 1.72e-21
C28635 a_n1641_46494# a_n2293_45010# 2.7e-19
C28636 a_11415_45002# a_413_45260# 0.063143f
C28637 a_12861_44030# a_18579_44172# 0.221909f
C28638 a_2698_46116# a_2437_43646# 6.23e-21
C28639 a_5066_45546# a_8336_45822# 8.57e-20
C28640 COMP_P a_21589_35634# 7.17e-19
C28641 a_n784_42308# a_11530_34132# 0.006009f
C28642 a_2952_47436# a_2905_45572# 0.318161f
C28643 a_n971_45724# a_6151_47436# 0.29974f
C28644 a_2063_45854# a_n1151_42308# 0.425035f
C28645 a_n1741_47186# a_7903_47542# 0.00805f
C28646 a_2553_47502# a_3160_47472# 2.08e-19
C28647 a_n785_47204# a_n443_46116# 2.37e-20
C28648 a_n3420_39616# a_n4064_39616# 6.66063f
C28649 a_n3565_39590# a_n2860_39866# 2.96e-19
C28650 a_7174_31319# comp_n 1.92e-19
C28651 a_16245_42852# VDD 0.205729f
C28652 a_n1630_35242# a_n1532_35090# 0.462421f
C28653 a_18579_44172# a_19700_43370# 0.175511f
C28654 a_7640_43914# a_7227_42852# 1.75e-20
C28655 a_n2661_42834# a_n4318_38680# 0.102282f
C28656 a_n2293_43922# a_n13_43084# 4.46e-21
C28657 a_1307_43914# a_2123_42473# 0.001341f
C28658 en_comp a_13070_42354# 4.34e-21
C28659 a_20205_31679# a_18194_35068# 1.48e-19
C28660 a_20692_30879# EN_VIN_BSTR_N 2.04e-19
C28661 a_11967_42832# a_16823_43084# 0.093759f
C28662 a_14539_43914# a_15567_42826# 1.35e-20
C28663 a_n356_44636# a_10991_42826# 4.8e-20
C28664 a_n699_43396# a_n2293_42282# 5.03e-21
C28665 a_n2017_45002# a_14113_42308# 0.006853f
C28666 a_9751_46155# VDD 7.28e-19
C28667 a_14021_43940# a_14401_32519# 0.059818f
C28668 a_5205_44484# a_6761_42308# 1.57e-19
C28669 a_17517_44484# a_13467_32519# 2.74e-21
C28670 a_10903_43370# a_8975_43940# 0.043009f
C28671 a_2324_44458# a_5518_44484# 0.112753f
C28672 a_n2293_45546# a_1423_45028# 0.06244f
C28673 a_15765_45572# a_16842_45938# 1.46e-19
C28674 a_n1613_43370# a_n2433_43396# 0.299968f
C28675 a_19692_46634# a_22485_44484# 1.22e-19
C28676 a_380_45546# a_375_42282# 3.56e-19
C28677 a_9290_44172# a_13720_44458# 2.01e-19
C28678 a_n2661_45546# a_2809_45348# 9.78e-19
C28679 a_2711_45572# a_4927_45028# 0.006854f
C28680 a_5257_43370# a_n2661_42282# 0.01339f
C28681 a_7499_43078# a_n2017_45002# 0.065458f
C28682 a_12741_44636# a_n2661_43922# 0.00322f
C28683 a_10809_44734# a_n2661_44458# 0.033319f
C28684 a_n863_45724# a_626_44172# 0.097275f
C28685 a_768_44030# a_n1925_46634# 5.22e-20
C28686 a_n881_46662# a_2107_46812# 0.138703f
C28687 a_n1435_47204# a_10554_47026# 3.08e-20
C28688 a_11459_47204# a_6755_46942# 1.05e-19
C28689 a_n1613_43370# a_1983_46706# 0.020434f
C28690 a_7754_40130# VDD 13.6809f
C28691 a_n4209_37414# C9_P_btm 1.91e-20
C28692 a_n3565_38216# VIN_P 0.029343f
C28693 a_19321_45002# a_19594_46812# 0.267862f
C28694 a_n1741_47186# a_12359_47026# 8.57e-21
C28695 a_2747_46873# a_3177_46902# 3.64e-20
C28696 a_4883_46098# a_4651_46660# 2e-19
C28697 a_22521_40055# a_22545_38993# 0.004924f
C28698 a_22459_39145# a_22521_39511# 0.075012f
C28699 a_11206_38545# CAL_P 0.234643f
C28700 a_22469_40625# a_22469_39537# 0.604831f
C28701 a_6151_47436# a_8023_46660# 1.79e-19
C28702 a_n1151_42308# a_12469_46902# 0.007465f
C28703 a_n4209_38216# VREF 0.055795f
C28704 a_12891_46348# a_n743_46660# 0.044305f
C28705 a_3357_43084# DATA[3] 0.066637f
C28706 a_n2433_43396# a_n1533_42852# 1.07e-19
C28707 a_4905_42826# a_5649_42852# 0.003104f
C28708 a_n2293_43922# a_11323_42473# 3.54e-20
C28709 a_9313_44734# a_15486_42560# 8.95e-20
C28710 a_n356_44636# a_17303_42282# 0.10316f
C28711 a_2437_43646# EN_OFFSET_CAL 7.51e-19
C28712 a_19237_31679# COMP_P 1.7e-20
C28713 a_n2661_45010# VDD 0.842431f
C28714 a_8685_43396# a_16243_43396# 3.52e-19
C28715 a_n1761_44111# a_n2104_42282# 1.67e-20
C28716 a_10341_43396# a_10765_43646# 7.4e-20
C28717 a_2982_43646# a_20556_43646# 8.33e-20
C28718 a_n1352_43396# a_n4318_38680# 2.18e-20
C28719 a_n97_42460# a_n13_43084# 0.13246f
C28720 a_n2293_46634# a_7765_42852# 6.5e-21
C28721 a_13661_43548# a_12545_42858# 1.24e-19
C28722 SMPL_ON_P a_n3674_37592# 0.051746f
C28723 a_18189_46348# a_15493_43940# 1.31e-20
C28724 a_3232_43370# a_3602_45348# 7.02e-20
C28725 a_n467_45028# a_n2293_42834# 8.59e-21
C28726 a_526_44458# a_8333_44056# 1.1e-21
C28727 a_12549_44172# a_17595_43084# 2.6e-20
C28728 a_n2497_47436# a_1184_42692# 3.5e-22
C28729 a_n971_45724# a_n473_42460# 0.094491f
C28730 a_2382_45260# a_2809_45028# 0.034331f
C28731 a_20107_45572# a_11827_44484# 2.61e-21
C28732 a_20623_45572# a_21005_45260# 0.002863f
C28733 a_20273_45572# a_21359_45002# 5.74e-20
C28734 a_20841_45814# a_21101_45002# 0.001934f
C28735 a_n1059_45260# a_n2661_43370# 0.03635f
C28736 a_10053_45546# a_9313_44734# 5.63e-20
C28737 a_4558_45348# a_5837_45348# 5.43e-21
C28738 a_5147_45002# a_5365_45348# 0.001577f
C28739 a_6709_45028# a_1423_45028# 2.16e-20
C28740 a_9482_43914# a_14537_43396# 0.040878f
C28741 a_11787_45002# a_1307_43914# 1.91e-21
C28742 a_3090_45724# a_14205_43396# 0.040425f
C28743 a_12861_44030# a_13003_42852# 6.07e-20
C28744 a_n2497_47436# a_n2293_45546# 0.307373f
C28745 a_5807_45002# a_6419_46155# 0.072498f
C28746 a_12991_46634# a_12816_46660# 0.233657f
C28747 a_n743_46660# a_805_46414# 0.064413f
C28748 a_n2438_43548# a_472_46348# 4.71e-19
C28749 a_n133_46660# a_376_46348# 0.004089f
C28750 a_n2661_46634# a_2698_46116# 1.4e-20
C28751 a_11459_47204# a_8049_45260# 2.62e-22
C28752 a_9313_45822# a_9241_46436# 1.86e-19
C28753 a_n881_46662# a_14493_46090# 0.011925f
C28754 a_11453_44696# a_10809_44734# 0.274367f
C28755 a_11309_47204# a_11133_46155# 0.040357f
C28756 a_4915_47217# a_14180_46482# 4.16e-19
C28757 a_n1151_42308# a_14383_46116# 1.15e-19
C28758 a_n1925_46634# a_1176_45822# 0.001268f
C28759 SMPL_ON_P a_n2840_45546# 8.99e-19
C28760 a_12549_44172# a_9290_44172# 0.053193f
C28761 a_12891_46348# a_11189_46129# 3.11e-20
C28762 a_171_46873# a_n1076_46494# 9.82e-20
C28763 a_3080_42308# a_5934_30871# 1.27306f
C28764 a_8855_44734# VDD 4.01e-19
C28765 a_16137_43396# a_16245_42852# 0.016079f
C28766 a_10835_43094# a_12545_42858# 3.81e-19
C28767 a_10922_42852# a_10341_42308# 0.053077f
C28768 a_10796_42968# a_12089_42308# 1.05e-19
C28769 a_2982_43646# a_6171_42473# 8.09e-20
C28770 a_n97_42460# a_11323_42473# 0.003208f
C28771 a_4185_45028# a_12545_42858# 3.65e-20
C28772 a_13661_43548# a_19332_42282# 1.85e-21
C28773 a_10193_42453# a_21381_43940# 1.29e-19
C28774 a_11691_44458# a_17970_44736# 0.040435f
C28775 a_n755_45592# a_8147_43396# 0.134231f
C28776 a_n357_42282# a_8791_43396# 1.18e-21
C28777 a_n913_45002# a_2889_44172# 6.01e-22
C28778 a_16147_45260# a_17973_43940# 1.63e-19
C28779 a_n1059_45260# a_2998_44172# 3.88e-20
C28780 a_n443_42852# a_3539_42460# 0.02291f
C28781 a_n2661_44458# a_5883_43914# 0.010478f
C28782 a_742_44458# a_2779_44458# 2.48e-21
C28783 a_11827_44484# a_18374_44850# 0.004504f
C28784 a_n2293_42834# a_n2661_43922# 0.03113f
C28785 a_n37_45144# a_175_44278# 8.37e-20
C28786 a_n863_45724# a_2813_43396# 1.63e-19
C28787 a_8953_45546# a_8037_42858# 0.017317f
C28788 a_8199_44636# a_8387_43230# 9.49e-20
C28789 a_13507_46334# a_18691_45572# 6.86e-21
C28790 a_n743_46660# a_11322_45546# 3.68e-19
C28791 a_3877_44458# a_2711_45572# 0.099631f
C28792 a_11415_45002# a_18985_46122# 9.02e-21
C28793 a_3483_46348# a_7920_46348# 4.08e-21
C28794 a_4704_46090# a_5204_45822# 1.24e-19
C28795 a_n971_45724# a_5111_44636# 0.381443f
C28796 a_17639_46660# a_10809_44734# 3.03e-19
C28797 a_n1435_47204# a_2437_43646# 0.191468f
C28798 a_n2293_46634# a_11823_42460# 0.072996f
C28799 a_765_45546# a_n1925_42282# 4.84e-20
C28800 a_584_46384# a_1667_45002# 3.89e-20
C28801 a_n1151_42308# a_n955_45028# 2.98e-19
C28802 a_2553_47502# a_413_45260# 0.004176f
C28803 a_n443_46116# a_n913_45002# 0.002757f
C28804 a_4883_46098# a_18341_45572# 1.94e-20
C28805 a_9313_45822# a_3357_43084# 2.85e-19
C28806 a_n881_46662# a_15903_45785# 0.032602f
C28807 a_12741_44636# a_18189_46348# 0.00488f
C28808 a_5068_46348# a_5164_46348# 0.31819f
C28809 a_16327_47482# a_20623_45572# 0.168593f
C28810 a_5342_30871# a_13657_42308# 1.2e-20
C28811 a_17538_32519# C9_N_btm 7.08e-19
C28812 a_3080_42308# a_11530_34132# 0.001927f
C28813 a_21381_43940# VDD 0.344882f
C28814 a_n3674_39304# a_n3690_39616# 4.64e-19
C28815 a_14635_42282# a_1606_42308# 1.94e-20
C28816 a_5193_42852# a_5932_42308# 8.62e-21
C28817 a_21588_30879# VREF 0.860047f
C28818 a_3232_43370# a_8685_43396# 8.91e-20
C28819 a_4185_45028# a_19332_42282# 1.64e-19
C28820 a_n2293_42834# a_n447_43370# 0.006668f
C28821 a_11967_42832# a_19279_43940# 0.070262f
C28822 a_17517_44484# a_22315_44484# 0.063928f
C28823 a_10193_42453# a_18249_42858# 0.038446f
C28824 a_n443_42852# a_9061_43230# 1.22e-20
C28825 a_n1925_42282# a_4921_42308# 1.23e-19
C28826 a_171_46873# VDD 0.539781f
C28827 a_12883_44458# a_12429_44172# 8.45e-19
C28828 a_5891_43370# a_7542_44172# 0.002369f
C28829 a_13249_42308# a_13635_43156# 0.004017f
C28830 a_11823_42460# a_5342_30871# 0.044603f
C28831 a_n2661_42834# a_1467_44172# 0.028215f
C28832 a_n2661_43922# a_1115_44172# 0.004853f
C28833 a_20362_44736# a_20679_44626# 0.102355f
C28834 a_n2661_43370# a_n2840_43370# 0.172532f
C28835 a_n2017_45002# a_15781_43660# 2.42e-20
C28836 a_n1925_46634# DATA[0] 2.87e-19
C28837 a_3537_45260# a_9803_43646# 2.53e-19
C28838 a_22612_30879# VIN_N 0.19035f
C28839 a_9290_44172# a_11525_45546# 0.001224f
C28840 a_10903_43370# a_10193_42453# 0.402091f
C28841 a_11189_46129# a_11322_45546# 0.05577f
C28842 a_13747_46662# a_21005_45260# 0.058269f
C28843 a_13885_46660# a_2437_43646# 1.22e-20
C28844 a_4883_46098# a_8975_43940# 0.018394f
C28845 a_3877_44458# a_4640_45348# 1.44e-20
C28846 a_10554_47026# a_10775_45002# 2.81e-22
C28847 a_19321_45002# a_18494_42460# 0.084551f
C28848 a_10249_46116# a_8953_45002# 9.14e-20
C28849 a_n881_46662# a_n2661_44458# 0.001141f
C28850 a_15227_44166# a_n2017_45002# 0.005144f
C28851 a_n1613_43370# a_n2433_44484# 0.29864f
C28852 a_n1151_42308# a_n2661_42834# 0.038196f
C28853 a_13259_45724# a_16375_45002# 0.60955f
C28854 a_11133_46155# a_10490_45724# 3.4e-20
C28855 a_10623_46897# a_10951_45334# 4.99e-21
C28856 a_526_44458# a_n443_42852# 2.06448f
C28857 a_6945_45028# a_6472_45840# 0.034109f
C28858 a_n784_42308# a_7754_40130# 0.001644f
C28859 a_5932_42308# comp_n 2.3e-19
C28860 a_1606_42308# a_n3420_37984# 6.06e-20
C28861 a_17531_42308# a_18057_42282# 0.00822f
C28862 a_17303_42282# a_18727_42674# 3.04e-19
C28863 a_4958_30871# a_18907_42674# 2.39e-20
C28864 a_17333_42852# RST_Z 1.2e-21
C28865 a_18249_42858# VDD 0.250132f
C28866 a_20447_31679# a_n1630_35242# 1.81e-19
C28867 a_n2017_45002# a_n1329_42308# 0.018315f
C28868 a_742_44458# a_n13_43084# 4.27e-21
C28869 a_20935_43940# a_15493_43940# 0.037795f
C28870 a_n2293_42834# a_3445_43172# 7.71e-20
C28871 a_8953_45546# DATA[4] 7.93e-19
C28872 a_10193_42453# a_21125_42558# 8.15e-20
C28873 a_n2956_37592# a_n2104_42282# 8.96e-21
C28874 en_comp a_n4318_38216# 0.064646f
C28875 a_n2810_45028# a_n3674_38216# 0.023217f
C28876 a_10903_43370# VDD 2.60588f
C28877 a_15682_43940# a_14021_43940# 5.96e-19
C28878 a_n2661_42282# a_5745_43940# 9.04e-20
C28879 a_644_44056# a_n97_42460# 1.26e-20
C28880 a_175_44278# a_104_43370# 1.89e-21
C28881 a_14815_43914# a_14205_43396# 1.84e-19
C28882 a_526_44458# a_375_42282# 0.007075f
C28883 a_2324_44458# a_10903_45394# 3.37e-19
C28884 a_11322_45546# a_11136_45572# 0.044092f
C28885 a_2711_45572# a_18175_45572# 1.3e-21
C28886 a_n2312_38680# a_n4318_39768# 0.023285f
C28887 a_3483_46348# a_11827_44484# 0.060892f
C28888 a_17339_46660# a_18287_44626# 0.018815f
C28889 a_6755_46942# a_16241_44484# 9.75e-20
C28890 a_768_44030# a_10949_43914# 0.007821f
C28891 a_5807_45002# a_n2661_42282# 1.81e-19
C28892 a_n2293_46098# a_n2433_44484# 1.34e-21
C28893 a_10193_42453# a_12016_45572# 0.001841f
C28894 a_10490_45724# a_11688_45572# 0.003828f
C28895 a_8049_45260# a_8191_45002# 0.084237f
C28896 a_7754_38968# VDAC_Ni 1.16e-19
C28897 a_2113_38308# a_3726_37500# 1.83e-19
C28898 a_n3420_39616# C0_P_btm 1.63e-20
C28899 a_n4064_39616# C2_P_btm 4.56e-20
C28900 a_21125_42558# VDD 0.004371f
C28901 a_n2109_47186# a_5167_46660# 0.004784f
C28902 a_n1741_47186# a_4817_46660# 8.55e-20
C28903 a_3160_47472# a_1799_45572# 1.08e-20
C28904 a_7903_47542# a_n743_46660# 8.42e-22
C28905 a_16327_47482# a_13747_46662# 0.128159f
C28906 a_16763_47508# a_5807_45002# 0.127783f
C28907 a_n443_46116# a_2107_46812# 0.075963f
C28908 a_11453_44696# a_n881_46662# 4.06e-20
C28909 a_10227_46804# a_16697_47582# 8.41e-19
C28910 a_2553_47502# a_2609_46660# 0.001405f
C28911 a_2952_47436# a_2443_46660# 5.83e-19
C28912 a_584_46384# a_2959_46660# 1.91e-19
C28913 a_n1435_47204# a_n2661_46634# 0.002772f
C28914 a_18184_42460# a_18057_42282# 0.19301f
C28915 a_14021_43940# a_22223_43396# 0.028989f
C28916 a_8333_44056# a_8605_42826# 6.56e-22
C28917 a_9028_43914# a_8037_42858# 1.46e-19
C28918 a_n356_44636# a_2713_42308# 1.57e-19
C28919 a_n2661_42834# a_n2840_42282# 0.001339f
C28920 a_16922_45042# a_19511_42282# 2.37e-20
C28921 a_6293_42852# a_6765_43638# 2.33e-20
C28922 a_2982_43646# a_3457_43396# 0.074308f
C28923 a_6031_43396# a_6547_43396# 0.105995f
C28924 a_18494_42460# a_17531_42308# 1.14e-19
C28925 a_19692_46634# a_14401_32519# 4.68e-19
C28926 a_13259_45724# a_13468_44734# 0.004213f
C28927 a_20205_31679# a_9313_44734# 1.02e-20
C28928 a_12549_44172# a_13467_32519# 3.15e-20
C28929 a_20202_43084# a_15493_43940# 0.02138f
C28930 a_11415_45002# a_22223_43948# 9.62e-19
C28931 a_5907_45546# a_5883_43914# 1.52e-20
C28932 a_3775_45552# a_n699_43396# 2.51e-21
C28933 a_2324_44458# a_2127_44172# 0.00237f
C28934 a_n143_45144# a_n37_45144# 0.13675f
C28935 a_n467_45028# a_413_45260# 2.64e-19
C28936 a_n913_45002# a_3537_45260# 0.148413f
C28937 a_n1151_42308# a_n2293_42282# 3.68e-19
C28938 a_14495_45572# a_11827_44484# 1.5e-20
C28939 a_8162_45546# a_n2661_44458# 1.47e-20
C28940 a_6511_45714# a_6298_44484# 0.001903f
C28941 w_1575_34946# COMP_P 2.48e-19
C28942 a_6151_47436# a_12594_46348# 2.73e-20
C28943 a_5807_45002# a_14226_46660# 2.03e-19
C28944 a_n2312_39304# a_n2840_46090# 0.007641f
C28945 a_7577_46660# a_7927_46660# 0.206455f
C28946 a_7715_46873# a_8667_46634# 1.39e-20
C28947 a_9313_45822# a_9625_46129# 0.018694f
C28948 a_n1435_47204# a_8199_44636# 1.19e-20
C28949 a_7411_46660# a_8492_46660# 0.102325f
C28950 a_4915_47217# a_13925_46122# 0.029041f
C28951 a_n4318_39304# a_n4318_37592# 0.023243f
C28952 a_15682_43940# a_15764_42576# 3.53e-20
C28953 a_16759_43396# a_16795_42852# 9.47e-19
C28954 a_16243_43396# a_17333_42852# 4.48e-19
C28955 a_743_42282# a_7765_42852# 8.69e-20
C28956 a_16137_43396# a_18249_42858# 0.021561f
C28957 a_18114_32519# C10_N_btm 0.460005f
C28958 a_19721_31679# C9_N_btm 1.91e-20
C28959 a_n901_43156# a_n13_43084# 0.014329f
C28960 a_n1991_42858# a_n1736_43218# 0.064178f
C28961 a_n1423_42826# a_n4318_38680# 1.78e-20
C28962 a_n1641_43230# a_n3674_39304# 1.48e-21
C28963 a_n2129_43609# a_n3674_38216# 1.65e-20
C28964 a_n2433_43396# a_n1736_42282# 5.66e-21
C28965 a_19929_45028# VDD 0.005632f
C28966 a_n1853_43023# a_n1545_43230# 0.004472f
C28967 a_4361_42308# a_4520_42826# 6.25e-20
C28968 a_n2267_43396# a_n2104_42282# 4.83e-20
C28969 a_10809_44734# a_9145_43396# 4.72e-20
C28970 SMPL_ON_P a_n2302_39072# 5.6e-20
C28971 a_n2661_43370# a_n4318_40392# 0.005935f
C28972 a_7229_43940# a_7640_43914# 0.177622f
C28973 a_3232_43370# a_8783_44734# 0.001081f
C28974 a_17719_45144# a_11827_44484# 2.79e-20
C28975 a_19778_44110# a_20567_45036# 0.044967f
C28976 a_16321_45348# a_16237_45028# 9.85e-19
C28977 a_16922_45042# a_19113_45348# 0.002269f
C28978 a_11322_45546# a_11750_44172# 5.99e-21
C28979 a_20841_45814# a_20766_44850# 3.35e-20
C28980 a_20623_45572# a_20835_44721# 3.31e-20
C28981 a_21188_45572# a_20640_44752# 1.97e-20
C28982 a_21363_45546# a_20679_44626# 3.09e-22
C28983 a_20692_30879# a_14401_32519# 0.054254f
C28984 a_18184_42460# a_18494_42460# 1.31047f
C28985 a_16327_47482# a_4958_30871# 2.84e-19
C28986 a_n2438_43548# a_n3674_37592# 0.001205f
C28987 a_10227_46804# a_17124_42282# 1.7e-20
C28988 a_18479_45785# a_20512_43084# 2.57e-19
C28989 a_10490_45724# a_12429_44172# 8.84e-22
C28990 a_413_45260# a_n2661_43922# 0.031184f
C28991 a_327_44734# a_n2661_42834# 0.001646f
C28992 a_5111_44636# a_9313_44734# 6.57e-20
C28993 a_5205_44484# a_5891_43370# 7.79e-20
C28994 a_n1613_43370# a_8685_42308# 0.002002f
C28995 a_n2312_38680# a_n2956_38216# 0.044798f
C28996 a_8145_46902# a_5066_45546# 6.07e-19
C28997 a_3090_45724# a_15682_46116# 6.43e-19
C28998 a_14976_45028# a_2324_44458# 0.086305f
C28999 a_9313_45822# a_9159_45572# 0.051702f
C29000 a_765_45546# a_2698_46116# 4.07e-20
C29001 a_11415_45002# a_20820_30879# 0.056772f
C29002 a_20202_43084# a_12741_44636# 0.22243f
C29003 a_4883_46098# a_10193_42453# 0.040505f
C29004 a_10227_46804# a_13904_45546# 5.42e-19
C29005 a_n2438_43548# a_n2840_45546# 9.23e-19
C29006 a_n2293_46634# a_n1079_45724# 0.002861f
C29007 a_n881_46662# a_5907_45546# 0.070761f
C29008 a_n1613_43370# a_6194_45824# 2.79e-20
C29009 a_n1021_46688# a_n2661_45546# 5.88e-21
C29010 a_15368_46634# a_14840_46494# 2.19e-19
C29011 a_8128_46384# a_2711_45572# 1.58e-19
C29012 a_14955_43940# VDD 0.253201f
C29013 a_5649_42852# a_15803_42450# 2.29e-19
C29014 a_16855_43396# a_4958_30871# 1.08e-19
C29015 a_n2293_42282# a_n2840_42282# 2.81e-19
C29016 a_15743_43084# a_19511_42282# 1.59e-20
C29017 a_4185_45028# a_5379_42460# 0.189676f
C29018 a_9482_43914# a_9165_43940# 0.002619f
C29019 a_21496_47436# RST_Z 5.48e-20
C29020 a_n967_45348# a_n1821_43396# 3.3e-19
C29021 a_18287_44626# a_18579_44172# 0.107662f
C29022 a_18989_43940# a_19279_43940# 0.053948f
C29023 a_742_44458# a_644_44056# 7.77e-19
C29024 a_21177_47436# SINGLE_ENDED 0.057266f
C29025 a_10227_46804# CLK 0.207445f
C29026 a_21588_30879# a_22521_40599# 8.64e-20
C29027 a_10903_43370# a_n784_42308# 1.58e-20
C29028 a_8199_44636# a_1606_42308# 2.7e-20
C29029 a_n1059_45260# a_1568_43370# 0.011697f
C29030 a_11823_42460# a_743_42282# 0.147603f
C29031 a_4883_46098# VDD 1.12729f
C29032 a_n357_42282# a_12895_43230# 0.00578f
C29033 a_1307_43914# a_3992_43940# 0.005165f
C29034 a_10193_42453# a_5649_42852# 0.003188f
C29035 a_n443_42852# a_8605_42826# 0.001815f
C29036 a_13507_46334# START 4.08e-19
C29037 a_3357_43084# a_2982_43646# 0.01988f
C29038 a_13747_46662# a_14537_43396# 0.006836f
C29039 a_n2661_46634# a_10775_45002# 3.04e-22
C29040 a_13661_43548# a_14797_45144# 0.116989f
C29041 a_5807_45002# a_15415_45028# 1.7e-21
C29042 a_1823_45246# a_1990_45899# 0.001705f
C29043 a_1799_45572# a_413_45260# 7.25e-20
C29044 a_n2661_46098# a_n37_45144# 1.2e-20
C29045 a_n1151_42308# a_n1352_44484# 0.001499f
C29046 a_3090_45724# a_16680_45572# 0.009229f
C29047 a_16327_47482# a_18911_45144# 3.79e-19
C29048 a_167_45260# a_1609_45822# 0.141505f
C29049 a_2107_46812# a_3537_45260# 1.32e-20
C29050 a_2063_45854# a_4223_44672# 1.1e-20
C29051 a_584_46384# a_n699_43396# 0.632931f
C29052 a_6540_46812# a_3357_43084# 0.001035f
C29053 a_18189_46348# a_16375_45002# 0.165328f
C29054 a_17957_46116# a_18243_46436# 0.010132f
C29055 a_n1925_46634# a_7276_45260# 8.36e-22
C29056 a_n2293_46098# a_6194_45824# 2.86e-19
C29057 a_2202_46116# a_2277_45546# 0.006767f
C29058 a_765_45546# a_13527_45546# 2.42e-21
C29059 a_n443_46116# a_n2661_44458# 0.034876f
C29060 a_15368_46634# a_16115_45572# 6.95e-20
C29061 a_1576_42282# a_7174_31319# 9.76e-21
C29062 a_5534_30871# VDAC_N 0.009192f
C29063 a_n4318_37592# a_n4334_40480# 7.27e-20
C29064 COMP_P a_n4315_30879# 3.39e-19
C29065 a_5649_42852# VDD 0.438443f
C29066 a_10533_42308# a_11323_42473# 0.002638f
C29067 a_n3674_38680# a_n4334_39616# 1.39e-19
C29068 a_13678_32519# RST_Z 0.048965f
C29069 a_17364_32525# C6_N_btm 2.76e-20
C29070 a_8975_43940# a_8685_43396# 2.13e-20
C29071 a_20512_43084# a_14021_43940# 0.030282f
C29072 a_n356_44636# a_6031_43396# 1.37e-20
C29073 a_21188_46660# VDD 0.284105f
C29074 a_21363_46634# RST_Z 2.85e-20
C29075 a_16922_45042# a_21259_43561# 0.108631f
C29076 a_20841_46902# SINGLE_ENDED 3.74e-21
C29077 a_11691_44458# a_18783_43370# 7.32e-20
C29078 a_n2293_42834# a_n1641_43230# 0.014975f
C29079 a_1307_43914# a_9127_43156# 5.14e-20
C29080 a_5883_43914# a_9145_43396# 0.004333f
C29081 a_3357_43084# a_5837_42852# 2.16e-20
C29082 a_9482_43914# a_12379_42858# 3.35e-19
C29083 a_n2661_42834# a_n1809_43762# 0.003072f
C29084 a_n2293_43922# a_104_43370# 1.18e-21
C29085 a_17517_44484# a_19319_43548# 3.23e-20
C29086 a_2804_46116# a_1307_43914# 3.01e-21
C29087 a_1138_42852# a_1423_45028# 7.83e-19
C29088 a_11133_46155# a_6171_45002# 4.63e-21
C29089 a_2324_44458# a_2382_45260# 0.044897f
C29090 a_11387_46155# a_3232_43370# 3.73e-20
C29091 a_765_45546# a_16922_45042# 6.35e-21
C29092 a_526_44458# a_2437_43646# 0.005693f
C29093 a_2711_45572# a_10053_45546# 0.018932f
C29094 a_6472_45840# a_6812_45938# 0.027606f
C29095 a_8199_44636# a_10775_45002# 0.064568f
C29096 a_6755_46942# a_16979_44734# 0.00119f
C29097 a_8270_45546# a_9838_44484# 4.89e-20
C29098 a_19321_45002# a_20640_44752# 0.034599f
C29099 a_16375_45002# a_17478_45572# 0.009252f
C29100 a_5937_45572# a_8953_45002# 0.062333f
C29101 a_5807_45002# a_19279_43940# 4.49e-20
C29102 a_13747_46662# a_20835_44721# 0.006757f
C29103 a_n2497_47436# a_1443_43940# 1.71e-19
C29104 a_n1613_43370# a_n2840_43914# 6.54e-20
C29105 a_n3565_38502# a_n3565_38216# 0.0433f
C29106 a_n3420_38528# a_n4209_38216# 0.050044f
C29107 a_n4209_38502# a_n3420_37984# 0.028231f
C29108 a_n4064_38528# a_n4251_38528# 0.001077f
C29109 a_n4064_40160# a_n4209_37414# 0.055461f
C29110 a_6151_47436# a_12465_44636# 0.025929f
C29111 a_n1741_47186# a_11309_47204# 0.01734f
C29112 a_n237_47217# a_7989_47542# 5.29e-20
C29113 a_n785_47204# a_n1613_43370# 3.89e-19
C29114 a_2124_47436# a_2583_47243# 6.64e-19
C29115 a_3160_47472# a_2747_46873# 2.93e-19
C29116 a_n4315_30879# a_n3565_37414# 0.037486f
C29117 a_6491_46660# a_4883_46098# 5.95e-21
C29118 a_1343_38525# a_3754_39466# 2.99e-19
C29119 a_7963_42308# VDD 0.266057f
C29120 a_15811_47375# a_15673_47210# 0.281607f
C29121 a_15507_47210# a_16241_47178# 0.06628f
C29122 a_11599_46634# a_16327_47482# 0.526398f
C29123 a_12861_44030# a_17591_47464# 0.079093f
C29124 a_13717_47436# a_10227_46804# 3.27e-19
C29125 a_6123_31319# RST_Z 0.004252f
C29126 a_5742_30871# C3_P_btm 0.030866f
C29127 a_14539_43914# a_16877_43172# 9.62e-19
C29128 en_comp a_1239_39587# 0.003125f
C29129 a_n97_42460# a_104_43370# 0.027998f
C29130 a_n1917_43396# a_n1821_43396# 0.013793f
C29131 a_n1699_43638# a_n1655_43396# 3.69e-19
C29132 a_11341_43940# a_10341_43396# 0.289072f
C29133 a_11967_42832# a_12545_42858# 0.028062f
C29134 a_15493_43940# a_14955_43396# 0.013181f
C29135 a_5263_45724# a_n2661_43370# 8.75e-19
C29136 a_2324_44458# a_15433_44458# 0.021739f
C29137 a_11778_45572# a_3232_43370# 1.29e-19
C29138 a_3090_45724# a_20269_44172# 1.17e-19
C29139 a_20205_31679# a_18114_32519# 0.051478f
C29140 a_20623_45572# a_20731_45938# 0.057222f
C29141 a_11682_45822# a_11787_45002# 4.49e-20
C29142 a_n357_42282# a_11827_44484# 1.01e-20
C29143 a_n2293_46634# a_2982_43646# 0.015801f
C29144 C3_P_btm C0_dummy_P_btm 0.087593f
C29145 C8_P_btm C3_N_btm 0.001059f
C29146 C6_P_btm C1_N_btm 3.17e-19
C29147 C5_P_btm C0_N_btm 1.4e-19
C29148 C4_P_btm C0_dummy_N_btm 1.24e-19
C29149 C2_P_btm C0_P_btm 0.698973f
C29150 a_n2661_46098# a_2443_46660# 0.063999f
C29151 a_1799_45572# a_2609_46660# 9.48e-20
C29152 EN_VIN_BSTR_N C10_N_btm 0.320569f
C29153 a_n1435_47204# a_765_45546# 0.00799f
C29154 a_11599_46634# a_16434_46987# 8.38e-20
C29155 a_n743_46660# a_4817_46660# 7.71e-20
C29156 a_n83_35174# VDD 0.313947f
C29157 a_8128_46384# a_8654_47026# 1.16e-19
C29158 a_5807_45002# a_9863_46634# 0.009219f
C29159 a_n815_47178# a_n901_46420# 3.99e-19
C29160 a_n2497_47436# a_1138_42852# 0.144386f
C29161 a_n971_45724# a_n1423_46090# 5.47e-19
C29162 a_n1925_46634# a_5167_46660# 0.008646f
C29163 a_15811_47375# a_16388_46812# 0.010369f
C29164 a_10227_46804# a_14035_46660# 0.035412f
C29165 a_12465_44636# a_19466_46812# 3.79e-20
C29166 a_11453_44696# a_17609_46634# 0.079593f
C29167 a_16409_43396# a_4361_42308# 2.27e-20
C29168 a_3626_43646# a_5534_30871# 0.082646f
C29169 a_8791_43396# a_8952_43230# 6.83e-19
C29170 a_9396_43370# a_9127_43156# 0.00282f
C29171 a_1307_43914# CLK 8.72e-21
C29172 a_16137_43396# a_5649_42852# 5.5e-20
C29173 a_2982_43646# a_5342_30871# 0.178973f
C29174 a_19268_43646# a_19177_43646# 0.001446f
C29175 a_15743_43084# a_21259_43561# 6.3e-20
C29176 a_18783_43370# a_4190_30871# 0.044615f
C29177 a_11963_45334# a_11827_44484# 3.47e-20
C29178 a_8696_44636# a_14112_44734# 8.58e-19
C29179 a_327_44734# a_n1352_44484# 5.64e-20
C29180 a_n2312_40392# a_n3674_38216# 0.025514f
C29181 a_1823_45246# a_3457_43396# 9.91e-20
C29182 a_16751_45260# a_16922_45042# 0.12103f
C29183 a_1307_43914# a_17023_45118# 9.26e-21
C29184 a_2711_45572# a_5244_44056# 3.02e-22
C29185 a_n755_45592# a_n2661_42282# 0.025718f
C29186 a_n1059_45260# a_5883_43914# 1.35e-19
C29187 a_n2312_39304# a_n2104_42282# 3.28e-20
C29188 SMPL_ON_N COMP_P 2.13516f
C29189 a_19692_46634# a_22223_43396# 0.001051f
C29190 a_12741_44636# a_14955_43396# 6.28e-23
C29191 a_5837_45348# a_n2661_43370# 4.55e-19
C29192 a_3537_45260# a_n2661_44458# 0.056342f
C29193 a_3483_46348# a_8147_43396# 2.1e-21
C29194 a_4185_45028# a_7287_43370# 1.18e-21
C29195 a_17339_46660# a_19268_43646# 0.003554f
C29196 a_17609_46634# a_17639_46660# 0.094289f
C29197 a_13059_46348# a_16388_46812# 8.68e-20
C29198 a_12816_46660# a_11415_45002# 5.41e-22
C29199 a_13885_46660# a_765_45546# 1.88e-20
C29200 a_4883_46098# a_20850_46155# 3.81e-19
C29201 a_171_46873# a_n1545_46494# 1.06e-20
C29202 a_n1925_46634# a_518_46482# 5.09e-19
C29203 a_n971_45724# a_9049_44484# 1.51e-21
C29204 a_n237_47217# a_8568_45546# 1.04e-19
C29205 a_4791_45118# a_6194_45824# 0.004919f
C29206 a_2063_45854# a_3260_45572# 5.14e-21
C29207 a_19466_46812# a_20528_46660# 9.92e-21
C29208 a_5257_43370# a_6165_46155# 0.11382f
C29209 a_6151_47436# a_2711_45572# 0.050517f
C29210 a_11309_47204# a_10586_45546# 1.36e-19
C29211 a_n2956_39768# a_n1925_42282# 7.32e-20
C29212 a_n2661_46634# a_526_44458# 9.72e-20
C29213 a_17730_32519# C8_N_btm 0.001799f
C29214 a_5649_42852# a_n784_42308# 0.043382f
C29215 a_n2157_42858# a_n4318_38216# 0.001336f
C29216 a_10341_42308# a_11554_42852# 0.170124f
C29217 a_10922_42852# a_10752_42852# 2.6e-19
C29218 a_3626_43646# a_19647_42308# 0.170024f
C29219 a_2982_43646# a_20107_42308# 0.003276f
C29220 a_n1991_42858# a_n3674_38680# 1.73e-20
C29221 a_743_42282# a_961_42354# 0.016854f
C29222 a_19237_31679# C6_N_btm 1.26e-20
C29223 a_10334_44484# a_9313_44734# 0.018652f
C29224 a_n2661_44458# a_11541_44484# 0.053139f
C29225 a_6171_45002# a_12429_44172# 1.87e-21
C29226 a_21076_30879# a_22400_42852# 1.76e-19
C29227 a_n1809_44850# a_n356_44636# 5.9e-21
C29228 a_5518_44484# a_5708_44484# 0.045837f
C29229 a_2779_44458# a_n2661_43922# 0.013114f
C29230 a_20567_45036# a_20159_44458# 0.001074f
C29231 a_n2293_42834# a_n809_44244# 0.001759f
C29232 a_11691_44458# a_16335_44484# 2.35e-19
C29233 a_n1605_47204# VDD 0.20224f
C29234 a_19256_45572# a_19319_43548# 8.54e-21
C29235 a_4223_44672# a_n2661_42834# 0.031905f
C29236 a_5105_45348# a_3905_42865# 3.58e-20
C29237 a_21101_45002# a_11967_42832# 1.52e-19
C29238 a_18494_42460# a_20362_44736# 0.004144f
C29239 a_19778_44110# a_20679_44626# 5.45e-21
C29240 a_11827_44484# a_18588_44850# 4.54e-19
C29241 a_n2109_47186# CLK_DATA 6.42e-19
C29242 a_7499_43078# a_8317_43396# 3.9e-19
C29243 a_10193_42453# a_8685_43396# 0.024858f
C29244 a_20205_31679# a_13887_32519# 0.051379f
C29245 a_5068_46348# a_5066_45546# 0.04842f
C29246 a_5204_45822# a_5210_46482# 6.82e-19
C29247 a_n1151_42308# a_5093_45028# 1.96e-21
C29248 a_n881_46662# a_n1059_45260# 0.121542f
C29249 a_2747_46873# a_413_45260# 0.038809f
C29250 a_n1613_43370# a_n913_45002# 0.686014f
C29251 a_4883_46098# a_5691_45260# 5.88e-21
C29252 a_10227_46804# a_10951_45334# 0.001109f
C29253 a_11599_46634# a_14537_43396# 6.07e-21
C29254 a_8199_44636# a_526_44458# 0.019697f
C29255 a_n237_47217# a_n2661_43370# 3.56e-19
C29256 a_8270_45546# a_8568_45546# 0.015327f
C29257 a_765_45546# a_380_45546# 0.141908f
C29258 a_20916_46384# a_20273_45572# 9.09e-20
C29259 a_22000_46634# a_20692_30879# 4.17e-19
C29260 a_13747_46662# a_20731_45938# 2.78e-19
C29261 a_13661_43548# a_19365_45572# 9.66e-20
C29262 a_5807_45002# a_19610_45572# 7.29e-19
C29263 a_13759_47204# a_2437_43646# 8.24e-20
C29264 a_6755_46942# a_11823_42460# 3.55e-19
C29265 a_13925_46122# a_10809_44734# 6.72e-20
C29266 a_18189_46348# a_18985_46122# 3.95e-21
C29267 a_17957_46116# a_18819_46122# 4.51e-21
C29268 a_13507_46334# a_6171_45002# 5.79e-20
C29269 a_196_42282# a_5934_30871# 3.42e-20
C29270 a_1606_42308# a_4921_42308# 4.1e-20
C29271 a_8685_43396# VDD 0.261626f
C29272 a_2713_42308# a_3823_42558# 6.62e-20
C29273 a_2903_42308# a_3318_42354# 0.003549f
C29274 a_n784_42308# a_7963_42308# 1.56e-20
C29275 a_1576_42282# a_5932_42308# 8.68e-21
C29276 a_4190_30871# VDAC_N 0.048399f
C29277 a_n2293_45010# a_791_42968# 3.6e-20
C29278 a_n913_45002# a_n1533_42852# 4.76e-20
C29279 a_13249_42308# a_13814_43218# 1.82e-19
C29280 a_n2293_43922# a_11341_43940# 0.026007f
C29281 a_n699_43396# a_n1177_43370# 0.060973f
C29282 a_6755_46942# DATA[3] 6.6e-21
C29283 a_n1899_43946# a_453_43940# 7e-20
C29284 a_10467_46802# CLK 0.028547f
C29285 a_n967_45348# a_n1736_43218# 0.001166f
C29286 a_n755_45592# a_3497_42558# 2.25e-19
C29287 a_949_44458# a_n97_42460# 1.25e-19
C29288 a_742_44458# a_104_43370# 5.46e-21
C29289 a_11453_44696# a_11541_44484# 0.004713f
C29290 a_3218_45724# a_3316_45546# 0.162813f
C29291 a_n1099_45572# a_n906_45572# 0.001923f
C29292 a_380_45546# a_509_45822# 0.062574f
C29293 a_8049_45260# a_11823_42460# 0.046281f
C29294 a_n2661_45546# a_n89_45572# 4.62e-19
C29295 a_n2293_46634# a_14539_43914# 0.045317f
C29296 a_8270_45546# a_n2661_43370# 0.022558f
C29297 a_n2497_47436# a_n4318_39768# 3e-20
C29298 a_12465_44636# a_12829_44484# 3.05e-19
C29299 a_n452_45724# a_n443_42852# 0.005182f
C29300 a_n863_45724# a_1609_45822# 0.117311f
C29301 a_n2661_46098# a_949_44458# 4.97e-22
C29302 a_768_44030# a_7640_43914# 0.036222f
C29303 a_13059_46348# a_13777_45326# 0.00155f
C29304 a_n1151_42308# a_n1549_44318# 5.94e-21
C29305 a_584_46384# a_1467_44172# 0.005691f
C29306 a_n2157_46122# a_n1059_45260# 8.24e-19
C29307 a_n1613_43370# a_556_44484# 3.24e-20
C29308 a_n901_46420# a_n2661_45010# 8.48e-21
C29309 a_20202_43084# a_413_45260# 3.33e-20
C29310 a_n1423_46090# a_n2293_45010# 1.94e-19
C29311 a_1823_45246# a_3357_43084# 0.062163f
C29312 a_10586_45546# a_10490_45724# 0.235237f
C29313 a_n755_45592# a_n310_45899# 6.91e-19
C29314 a_16327_47482# a_19615_44636# 6.71e-19
C29315 a_n4064_40160# a_n3607_39616# 5.58e-20
C29316 a_5934_30871# a_n4064_37440# 0.003932f
C29317 COMP_P a_19864_35138# 3.57e-19
C29318 a_n971_45724# a_5815_47464# 7.7e-19
C29319 a_584_46384# a_n1151_42308# 0.047349f
C29320 a_2553_47502# a_2905_45572# 8.68e-19
C29321 a_n1741_47186# a_7227_47204# 0.016018f
C29322 a_n237_47217# a_4915_47217# 0.071869f
C29323 a_2063_45854# a_3160_47472# 0.005303f
C29324 a_n3420_39616# a_n2946_39866# 0.236674f
C29325 a_7174_31319# a_1736_39043# 7.24e-20
C29326 a_n4315_30879# a_n4209_39304# 0.032541f
C29327 a_15953_42852# VDD 0.005646f
C29328 a_n4209_39590# a_n2216_39866# 0.001361f
C29329 a_n3565_39590# a_n2302_39866# 0.044102f
C29330 a_n3690_39616# a_n4064_39616# 0.085414f
C29331 a_n1630_35242# a_n1386_35608# 0.019114f
C29332 a_n2661_42834# a_n3674_39304# 0.038671f
C29333 a_n2293_43922# a_n1076_43230# 1.7e-20
C29334 a_1307_43914# a_1755_42282# 1.63e-19
C29335 en_comp a_12563_42308# 8.68e-21
C29336 a_20205_31679# EN_VIN_BSTR_N 0.003421f
C29337 a_18579_44172# a_19268_43646# 6.28e-19
C29338 a_n356_44636# a_10796_42968# 4.72e-20
C29339 a_14539_43914# a_5342_30871# 2.82e-20
C29340 a_n2017_45002# a_13657_42558# 0.0086f
C29341 a_3537_45260# a_8325_42308# 3.11e-21
C29342 a_5111_44636# a_8515_42308# 5.49e-21
C29343 a_14021_43940# a_21381_43940# 0.022437f
C29344 a_11341_43940# a_n97_42460# 1.85e-19
C29345 a_18597_46090# a_2982_43646# 0.239147f
C29346 a_12549_44172# a_19319_43548# 0.024381f
C29347 a_2324_44458# a_5343_44458# 0.255488f
C29348 a_10903_43370# a_10057_43914# 0.052284f
C29349 a_15599_45572# a_16211_45572# 3.82e-19
C29350 a_n1613_43370# a_n4318_39304# 3.19e-20
C29351 a_19692_46634# a_20512_43084# 0.387138f
C29352 a_n2661_45546# a_2304_45348# 0.004487f
C29353 a_2711_45572# a_5111_44636# 0.00298f
C29354 a_12741_44636# a_n2661_42834# 5.02e-19
C29355 a_n443_42852# a_8953_45002# 2.1e-20
C29356 a_n863_45724# a_501_45348# 2.59e-19
C29357 a_n4209_37414# C10_P_btm 2.25e-20
C29358 a_22521_40055# a_22521_39511# 0.457858f
C29359 a_22469_40625# a_22821_38993# 0.002743f
C29360 VDAC_P CAL_P 6.16e-21
C29361 a_22521_40599# a_22469_39537# 0.380006f
C29362 a_n881_46662# a_948_46660# 0.002487f
C29363 a_9313_45822# a_6755_46942# 0.031706f
C29364 a_n1613_43370# a_2107_46812# 0.05377f
C29365 a_5807_45002# a_20916_46384# 3.09e-20
C29366 a_n1741_47186# a_12156_46660# 0.005703f
C29367 a_2747_46873# a_2609_46660# 0.347674f
C29368 a_4883_46098# a_4646_46812# 0.028054f
C29369 a_6545_47178# a_6903_46660# 5.61e-19
C29370 a_6151_47436# a_8654_47026# 7.05e-19
C29371 a_6491_46660# a_6682_46660# 2.88e-19
C29372 a_n1151_42308# a_11901_46660# 0.020194f
C29373 a_4915_47217# a_8270_45546# 1.62e-19
C29374 a_11309_47204# a_n743_46660# 0.001744f
C29375 a_14021_43940# a_18249_42858# 4.16e-20
C29376 a_3626_43646# a_4190_30871# 0.070713f
C29377 a_9145_43396# a_14621_43646# 0.00367f
C29378 a_2437_43646# DATA[5] 0.059749f
C29379 a_n2293_43922# a_10723_42308# 8.6e-20
C29380 a_9313_44734# a_15051_42282# 2.49e-19
C29381 a_n356_44636# a_4958_30871# 0.46356f
C29382 a_n2840_45002# VDD 0.289706f
C29383 a_8685_43396# a_16137_43396# 0.003201f
C29384 a_n2065_43946# a_n2104_42282# 2.12e-21
C29385 a_2982_43646# a_743_42282# 0.047135f
C29386 a_n97_42460# a_n1076_43230# 4.69e-19
C29387 a_n2293_46634# a_7871_42858# 6.83e-20
C29388 a_17715_44484# a_15493_43940# 0.005403f
C29389 a_13556_45296# a_13777_45326# 0.101558f
C29390 a_9049_44484# a_9313_44734# 0.034936f
C29391 a_4646_46812# a_5649_42852# 1.19e-20
C29392 a_n971_45724# a_n961_42308# 3.58e-20
C29393 a_2382_45260# a_2448_45028# 0.009378f
C29394 a_20205_31679# a_22485_44484# 2.08e-20
C29395 a_20273_45572# a_21101_45002# 0.014321f
C29396 a_20623_45572# a_20567_45036# 0.001339f
C29397 a_20841_45814# a_21005_45260# 3.92e-20
C29398 a_n2017_45002# a_n2661_43370# 0.038361f
C29399 a_5147_45002# a_5105_45348# 2.26e-21
C29400 a_4558_45348# a_5365_45348# 7.9e-20
C29401 a_7229_43940# a_1423_45028# 0.024468f
C29402 a_13348_45260# a_14537_43396# 3.8e-20
C29403 a_13017_45260# a_15415_45028# 5.39e-21
C29404 a_10951_45334# a_1307_43914# 3.62e-21
C29405 a_9482_43914# a_14180_45002# 0.022677f
C29406 a_3090_45724# a_14358_43442# 6.05e-19
C29407 a_10903_43370# a_14021_43940# 2.56e-21
C29408 a_n2497_47436# a_n2956_38216# 8.23e-20
C29409 a_5807_45002# a_6165_46155# 0.039202f
C29410 a_12251_46660# a_12816_46660# 7.99e-20
C29411 a_n743_46660# a_472_46348# 0.076758f
C29412 a_2107_46812# a_n2293_46098# 1.3e-19
C29413 a_n2661_46634# a_2521_46116# 4.54e-20
C29414 a_9313_45822# a_8049_45260# 0.086184f
C29415 a_n881_46662# a_13925_46122# 0.019683f
C29416 a_11453_44696# a_22223_46124# 1.39e-21
C29417 SMPL_ON_N a_10809_44734# 0.002895f
C29418 a_11309_47204# a_11189_46129# 0.03753f
C29419 a_4915_47217# a_12638_46436# 2.75e-20
C29420 a_n2293_46634# a_1823_45246# 0.230429f
C29421 a_n1925_46634# a_1208_46090# 0.005309f
C29422 a_n2109_47186# a_n2661_45546# 4.99e-20
C29423 a_12891_46348# a_9290_44172# 1.02e-19
C29424 a_171_46873# a_n901_46420# 2.27e-19
C29425 a_3539_42460# a_4921_42308# 3.77e-19
C29426 a_8783_44734# VDD 4.43e-19
C29427 a_16137_43396# a_15953_42852# 2.65e-19
C29428 a_10991_42826# a_10341_42308# 0.035667f
C29429 a_10835_43094# a_12089_42308# 2.32e-19
C29430 a_10796_42968# a_12379_42858# 3.81e-19
C29431 a_2982_43646# a_5755_42308# 2.01e-19
C29432 a_n97_42460# a_10723_42308# 7.44e-19
C29433 a_4185_45028# a_12089_42308# 3.84e-20
C29434 a_15861_45028# a_15493_43940# 4.14e-20
C29435 a_11691_44458# a_17767_44458# 0.060949f
C29436 a_n357_42282# a_8147_43396# 8.81e-19
C29437 a_n913_45002# a_2675_43914# 2.72e-20
C29438 a_n1059_45260# a_2889_44172# 4.48e-22
C29439 a_16147_45260# a_17737_43940# 8.05e-21
C29440 a_n2017_45002# a_2998_44172# 2.57e-20
C29441 a_n443_42852# a_3626_43646# 0.027303f
C29442 a_n2661_44458# a_8701_44490# 0.00716f
C29443 a_742_44458# a_949_44458# 0.185221f
C29444 a_16237_45028# a_14539_43914# 1.93e-19
C29445 a_11827_44484# a_18443_44721# 0.007717f
C29446 a_n2293_42834# a_n2661_42834# 0.202366f
C29447 a_15227_44166# a_17749_42852# 0.00177f
C29448 a_5257_43370# a_5379_42460# 7.23e-20
C29449 a_8953_45546# a_7765_42852# 3.74e-21
C29450 a_8199_44636# a_8605_42826# 1.4e-21
C29451 a_11415_45002# a_18819_46122# 1.5e-20
C29452 a_3483_46348# a_6419_46155# 2.02e-21
C29453 a_4704_46090# a_5164_46348# 5.86e-19
C29454 a_4419_46090# a_5204_45822# 0.001858f
C29455 a_12816_46660# a_13259_45724# 1.31e-19
C29456 a_13381_47204# a_2437_43646# 0.005327f
C29457 a_12465_44636# a_16147_45260# 2.41e-21
C29458 a_765_45546# a_526_44458# 5.75e-20
C29459 a_n237_47217# a_4574_45260# 3.04e-20
C29460 a_2063_45854# a_413_45260# 0.031952f
C29461 a_584_46384# a_327_44734# 0.040089f
C29462 a_n443_46116# a_n1059_45260# 3.62e-19
C29463 a_4791_45118# a_n913_45002# 0.254334f
C29464 a_4883_46098# a_18479_45785# 8.72e-20
C29465 a_11031_47542# a_3357_43084# 1.35e-19
C29466 a_n881_46662# a_15599_45572# 0.601034f
C29467 a_12741_44636# a_17715_44484# 0.029877f
C29468 a_n743_46660# a_10490_45724# 2.02e-20
C29469 a_16327_47482# a_20841_45814# 0.161808f
C29470 a_n4318_38680# a_n4334_39616# 1.78e-19
C29471 a_17538_32519# C8_N_btm 0.090298f
C29472 a_14401_32519# C10_N_btm 3.37e-20
C29473 a_7573_43172# a_6123_31319# 2.33e-20
C29474 a_5534_30871# a_13921_42308# 5.65e-20
C29475 a_19741_43940# VDD 0.153579f
C29476 a_13291_42460# a_1606_42308# 1.35e-20
C29477 a_5837_42852# a_5755_42308# 4.85e-19
C29478 a_17701_42308# a_15890_42674# 2.84e-21
C29479 a_11823_42460# a_15279_43071# 0.010476f
C29480 a_4185_45028# a_18907_42674# 7.14e-20
C29481 a_n133_46660# VDD 0.483405f
C29482 a_n2293_42834# a_n1352_43396# 0.006475f
C29483 a_11967_42832# a_20766_44850# 0.042853f
C29484 a_17517_44484# a_3422_30871# 0.073987f
C29485 a_18479_45785# a_5649_42852# 4.56e-21
C29486 a_10193_42453# a_17333_42852# 0.032471f
C29487 a_n443_42852# a_8649_43218# 6.31e-19
C29488 a_526_44458# a_4921_42308# 0.002257f
C29489 a_5111_44636# a_7466_43396# 0.002133f
C29490 a_12607_44458# a_12429_44172# 4.52e-19
C29491 a_5891_43370# a_7281_43914# 4.34e-19
C29492 a_n2661_46634# DATA[5] 6.56e-19
C29493 a_20159_44458# a_20679_44626# 0.043567f
C29494 a_20362_44736# a_20640_44752# 0.118759f
C29495 a_n2661_43922# a_644_44056# 1.23e-19
C29496 a_7640_43914# a_7845_44172# 0.021949f
C29497 a_n2661_42834# a_1115_44172# 0.011443f
C29498 a_n2017_45002# a_15681_43442# 1.9e-21
C29499 a_3537_45260# a_9145_43396# 0.002981f
C29500 a_21588_30879# VIN_N 0.106594f
C29501 a_13249_42308# a_12895_43230# 0.002542f
C29502 a_9290_44172# a_11322_45546# 0.077646f
C29503 a_11387_46155# a_10193_42453# 0.050391f
C29504 a_10903_43370# a_10180_45724# 7.78e-20
C29505 a_13747_46662# a_20567_45036# 0.026034f
C29506 a_4883_46098# a_10057_43914# 2.16e-19
C29507 a_3877_44458# a_4185_45348# 7.28e-19
C29508 a_10623_46897# a_10775_45002# 3.09e-22
C29509 a_19321_45002# a_18184_42460# 0.094476f
C29510 a_6969_46634# a_6709_45028# 9.02e-22
C29511 a_6755_46942# a_7705_45326# 1.11e-20
C29512 a_n1613_43370# a_n2661_44458# 0.05666f
C29513 a_12741_44636# a_15861_45028# 0.075863f
C29514 a_3483_46348# a_10907_45822# 0.140023f
C29515 a_11189_46129# a_10490_45724# 0.03271f
C29516 a_10467_46802# a_10951_45334# 2.26e-21
C29517 a_1123_46634# a_n2661_43370# 3.92e-21
C29518 a_526_44458# a_509_45822# 1.55e-20
C29519 a_5932_42308# a_1736_39043# 8.72e-20
C29520 a_17303_42282# a_18057_42282# 7.14e-19
C29521 a_4958_30871# a_18727_42674# 2.08e-20
C29522 a_18083_42858# RST_Z 1.06e-20
C29523 a_n1630_35242# a_2113_38308# 4.08e-20
C29524 a_17333_42852# VDD 0.525529f
C29525 a_5742_30871# a_n3565_39590# 7.02e-21
C29526 a_n2017_45002# COMP_P 0.012669f
C29527 a_14539_43914# a_743_42282# 3.58e-20
C29528 a_20623_43914# a_15493_43940# 0.040969f
C29529 a_21115_43940# a_11341_43940# 0.008031f
C29530 a_n2293_42834# a_n2293_42282# 0.018879f
C29531 a_5937_45572# DATA[4] 8.55e-21
C29532 a_n2293_43922# a_10341_43396# 0.022718f
C29533 a_n2956_37592# a_n4318_38216# 0.023067f
C29534 a_11387_46155# VDD 0.099732f
C29535 a_14955_43940# a_14021_43940# 1.99e-20
C29536 a_175_44278# a_n97_42460# 2.88e-20
C29537 a_n2810_45028# a_n2104_42282# 9.69e-21
C29538 en_comp a_n2472_42282# 0.018838f
C29539 a_8016_46348# CLK 0.001431f
C29540 a_2324_44458# a_8560_45348# 0.070986f
C29541 a_10586_45546# a_6171_45002# 0.001629f
C29542 a_2711_45572# a_16147_45260# 0.028186f
C29543 a_3090_45724# a_10617_44484# 0.003583f
C29544 a_n1925_42282# a_1307_43914# 0.03653f
C29545 a_n1151_42308# a_n1177_43370# 3.34e-19
C29546 a_17339_46660# a_18248_44752# 0.019889f
C29547 a_12549_44172# a_10949_43914# 0.052089f
C29548 a_768_44030# a_10729_43914# 0.004644f
C29549 a_n2293_46098# a_n2661_44458# 0.026753f
C29550 a_n2472_46090# a_n2433_44484# 5.65e-21
C29551 a_10490_45724# a_11136_45572# 0.048799f
C29552 a_10193_42453# a_11778_45572# 0.004713f
C29553 a_8049_45260# a_7705_45326# 0.032872f
C29554 a_22775_42308# RST_Z 0.001998f
C29555 a_n4064_39072# EN_VIN_BSTR_P 0.959329f
C29556 a_n2109_47186# a_5385_46902# 0.013334f
C29557 a_n1741_47186# a_4955_46873# 2.85e-19
C29558 a_2905_45572# a_1799_45572# 0.002025f
C29559 a_2747_46873# a_3094_47570# 2.88e-19
C29560 a_4883_46098# a_9804_47204# 0.020011f
C29561 a_16327_47482# a_13661_43548# 0.132061f
C29562 a_16023_47582# a_5807_45002# 0.00104f
C29563 a_4791_45118# a_2107_46812# 0.078338f
C29564 a_6575_47204# a_n1925_46634# 3.37e-19
C29565 a_7754_38968# a_7754_38636# 0.296258f
C29566 a_3754_39134# a_3754_38470# 2.48e-19
C29567 a_10227_46804# a_16285_47570# 0.002099f
C29568 a_2063_45854# a_2609_46660# 0.005947f
C29569 a_2553_47502# a_2443_46660# 0.001147f
C29570 a_584_46384# a_3177_46902# 9.68e-20
C29571 a_n3420_39616# C1_P_btm 1.92e-20
C29572 a_n4064_39616# C3_P_btm 5.52e-20
C29573 a_n1435_47204# a_n2956_39768# 1.18e-19
C29574 a_6293_42852# a_6197_43396# 0.213423f
C29575 a_n97_42460# a_10341_43396# 0.917198f
C29576 a_11967_42832# a_13157_43218# 0.002086f
C29577 en_comp a_3754_38470# 7.78e-19
C29578 a_8333_44056# a_8037_42858# 2.79e-21
C29579 a_14021_43940# a_5649_42852# 0.005268f
C29580 a_2982_43646# a_2813_43396# 0.096538f
C29581 a_6031_43396# a_6765_43638# 0.053479f
C29582 a_18184_42460# a_17531_42308# 0.001442f
C29583 a_18494_42460# a_17303_42282# 6.74e-19
C29584 a_n755_45592# a_n310_44811# 0.001544f
C29585 a_19692_46634# a_21381_43940# 0.022586f
C29586 a_13259_45724# a_13213_44734# 0.020051f
C29587 a_12861_44030# a_12895_43230# 3e-19
C29588 a_4646_46812# a_8685_43396# 7.39e-20
C29589 a_11415_45002# a_11341_43940# 6.83e-19
C29590 a_n955_45028# a_413_45260# 1.19e-20
C29591 a_n1059_45260# a_3537_45260# 0.162323f
C29592 a_13249_42308# a_11827_44484# 0.029876f
C29593 a_6472_45840# a_6298_44484# 0.002101f
C29594 a_3877_44458# a_6903_46660# 0.007019f
C29595 a_5807_45002# a_16751_46987# 0.001109f
C29596 a_13759_47204# a_765_45546# 5.9e-19
C29597 a_16327_47482# a_4185_45028# 1.37e-19
C29598 a_7577_46660# a_8145_46902# 0.170059f
C29599 a_5385_46902# a_5841_46660# 4.2e-19
C29600 a_7715_46873# a_7927_46660# 3.12e-19
C29601 a_9313_45822# a_8953_45546# 0.038855f
C29602 a_7411_46660# a_8667_46634# 0.043475f
C29603 a_6540_46812# a_6755_46942# 0.057503f
C29604 a_5732_46660# a_6969_46634# 3.02e-20
C29605 a_4915_47217# a_13759_46122# 0.024639f
C29606 a_12549_44172# a_20411_46873# 1.31e-20
C29607 a_16977_43638# a_16795_42852# 7.5e-19
C29608 a_743_42282# a_7871_42858# 9.63e-20
C29609 a_16137_43396# a_17333_42852# 0.01487f
C29610 a_18114_32519# C9_N_btm 0.003109f
C29611 a_19721_31679# C8_N_btm 1.65e-20
C29612 a_n901_43156# a_n1076_43230# 0.234322f
C29613 a_n1853_43023# a_n1736_43218# 0.183149f
C29614 a_n1991_42858# a_n4318_38680# 5.47e-19
C29615 a_n2433_43396# a_n3674_38216# 8.11e-21
C29616 a_18545_45144# VDD 3.69e-20
C29617 a_n2157_42858# a_n1545_43230# 3.82e-19
C29618 a_3626_43646# a_14635_42282# 0.002593f
C29619 a_n2129_43609# a_n2104_42282# 1.48e-19
C29620 SMPL_ON_P a_n4064_39072# 1.17e-20
C29621 a_5093_45028# a_4223_44672# 4.9e-19
C29622 a_8704_45028# a_n2661_44458# 1.59e-19
C29623 a_7229_43940# a_6109_44484# 5.71e-20
C29624 a_3232_43370# a_8333_44734# 8.77e-20
C29625 a_7276_45260# a_7640_43914# 1.59e-19
C29626 a_17613_45144# a_11827_44484# 9.36e-21
C29627 a_526_44458# a_6452_43396# 9.65e-19
C29628 a_20841_45814# a_20835_44721# 0.001113f
C29629 a_20107_45572# a_19279_43940# 1.81e-19
C29630 a_20623_45572# a_20679_44626# 6.43e-21
C29631 a_21363_45546# a_20640_44752# 9.91e-23
C29632 a_20528_45572# a_20159_44458# 2.85e-20
C29633 a_20205_31679# a_14401_32519# 0.054064f
C29634 a_19778_44110# a_18494_42460# 0.04586f
C29635 a_10227_46804# a_16522_42674# 2.46e-19
C29636 a_3483_46348# a_16823_43084# 8.97e-20
C29637 a_1823_45246# a_743_42282# 0.06422f
C29638 a_10193_42453# a_13483_43940# 2.57e-19
C29639 a_10490_45724# a_11750_44172# 1.05e-21
C29640 a_413_45260# a_n2661_42834# 0.023284f
C29641 a_n37_45144# a_n2661_43922# 4.45e-20
C29642 a_11652_45724# a_10729_43914# 5.99e-20
C29643 a_n2661_43370# a_n2840_44458# 0.011391f
C29644 a_n1613_43370# a_8325_42308# 2.95e-20
C29645 a_7577_46660# a_5066_45546# 1.32e-19
C29646 a_3090_45724# a_2324_44458# 0.684819f
C29647 a_14976_45028# a_14840_46494# 0.010576f
C29648 a_765_45546# a_2521_46116# 3.87e-20
C29649 a_20202_43084# a_20820_30879# 0.005846f
C29650 a_22365_46825# a_12741_44636# 0.062216f
C29651 a_4883_46098# a_10180_45724# 0.001751f
C29652 a_10227_46804# a_13527_45546# 6.04e-19
C29653 a_n2293_46634# a_n2293_45546# 0.065405f
C29654 a_n881_46662# a_5263_45724# 0.180025f
C29655 a_11415_45002# a_22591_46660# 0.172844f
C29656 a_n1613_43370# a_5907_45546# 2.13e-20
C29657 a_n1925_46634# a_n2661_45546# 5.29e-20
C29658 a_15368_46634# a_15015_46420# 0.012546f
C29659 a_n1151_42308# a_8696_44636# 5.67e-21
C29660 a_13483_43940# VDD 0.219591f
C29661 a_5649_42852# a_15764_42576# 1.57e-19
C29662 a_5755_42852# a_5932_42308# 0.012644f
C29663 a_4361_42308# a_15890_42674# 0.004318f
C29664 a_21177_47436# START 7.35e-20
C29665 a_4185_45028# a_5267_42460# 9.17e-19
C29666 a_13507_46334# RST_Z 0.004909f
C29667 a_n967_45348# a_n1190_43762# 1.32e-19
C29668 a_18248_44752# a_18579_44172# 0.001274f
C29669 a_18287_44626# a_18245_44484# 2.56e-19
C29670 a_20990_47178# SINGLE_ENDED 0.067698f
C29671 a_2437_43646# a_3626_43646# 6e-20
C29672 a_n143_45144# a_n97_42460# 1.93e-21
C29673 a_n913_45002# a_1209_43370# 7.74e-20
C29674 a_n2017_45002# a_1568_43370# 4.02e-19
C29675 a_n2661_44458# a_2675_43914# 9.03e-20
C29676 a_n357_42282# a_13113_42826# 0.008588f
C29677 a_1307_43914# a_3737_43940# 0.058797f
C29678 a_n443_42852# a_8037_42858# 0.007515f
C29679 a_21496_47436# VDD 0.198362f
C29680 a_3357_43084# a_2896_43646# 2.67e-19
C29681 a_17957_46116# a_18147_46436# 0.011458f
C29682 a_10809_44734# a_12638_46436# 0.003187f
C29683 a_13747_46662# a_14180_45002# 5.33e-19
C29684 a_13661_43548# a_14537_43396# 0.505634f
C29685 a_n1741_47186# a_12607_44458# 1.63e-22
C29686 a_n743_46660# a_6171_45002# 0.140224f
C29687 a_n2438_43548# a_3232_43370# 8.07e-21
C29688 a_n2661_46634# a_8953_45002# 2.39e-20
C29689 a_n2661_46098# a_n143_45144# 2.28e-22
C29690 a_n1151_42308# a_n1177_44458# 0.021669f
C29691 a_2063_45854# a_2779_44458# 1.24e-20
C29692 a_3090_45724# a_16855_45546# 0.007982f
C29693 a_16327_47482# a_18587_45118# 0.002342f
C29694 a_768_44030# a_1423_45028# 0.096238f
C29695 a_167_45260# a_n443_42852# 0.246952f
C29696 a_4419_46090# a_3503_45724# 3.27e-21
C29697 a_584_46384# a_4223_44672# 0.044788f
C29698 a_5732_46660# a_3357_43084# 0.017659f
C29699 a_12861_44030# a_11827_44484# 0.466435f
C29700 a_17715_44484# a_16375_45002# 0.026655f
C29701 a_n1925_46634# a_5205_44484# 3.1e-21
C29702 a_n2293_46098# a_5907_45546# 4.2e-19
C29703 a_1823_45246# a_2277_45546# 3.97e-20
C29704 a_2107_46812# a_3429_45260# 3.88e-21
C29705 a_15368_46634# a_16333_45814# 3.38e-20
C29706 a_4791_45118# a_n2661_44458# 0.095212f
C29707 a_765_45546# a_13163_45724# 4.54e-21
C29708 a_17364_32525# C5_N_btm 2.13e-20
C29709 a_n3674_38216# a_n4064_40160# 0.02459f
C29710 a_13678_32519# VDD 0.454512f
C29711 a_14209_32519# C7_N_btm 1.64e-19
C29712 a_10533_42308# a_10723_42308# 0.23663f
C29713 a_1067_42314# a_7174_31319# 4.88e-21
C29714 a_10057_43914# a_8685_43396# 0.007406f
C29715 a_n356_44636# a_1512_43396# 5.7e-20
C29716 a_21363_46634# VDD 0.357368f
C29717 a_20623_46660# RST_Z 2.19e-20
C29718 a_765_45546# DATA[5] 0.027477f
C29719 a_20273_46660# SINGLE_ENDED 1.13e-20
C29720 a_11691_44458# a_18525_43370# 1.92e-20
C29721 a_11827_44484# a_19700_43370# 4.41e-21
C29722 a_n2293_42834# a_n1423_42826# 0.011631f
C29723 a_1307_43914# a_8387_43230# 3.33e-20
C29724 a_n2661_42834# a_n2012_43396# 0.001847f
C29725 a_n2293_43922# a_n97_42460# 0.136247f
C29726 a_n2661_43922# a_104_43370# 7.49e-21
C29727 a_2711_45572# a_9049_44484# 0.025215f
C29728 a_2698_46116# a_1307_43914# 2.53e-20
C29729 a_3483_46348# a_15415_45028# 5.74e-21
C29730 a_1823_45246# a_626_44172# 2.16e-20
C29731 a_11189_46129# a_6171_45002# 7.06e-21
C29732 a_2324_44458# a_2274_45254# 0.007089f
C29733 a_9313_45822# a_9028_43914# 3.91e-20
C29734 a_n743_46660# a_14673_44172# 3.65e-21
C29735 a_1138_42852# a_1145_45348# 1.86e-19
C29736 a_17339_46660# a_16922_45042# 0.02918f
C29737 a_167_45260# a_375_42282# 0.017297f
C29738 a_8270_45546# a_5883_43914# 0.20967f
C29739 a_6755_46942# a_14539_43914# 0.094724f
C29740 a_19321_45002# a_20362_44736# 0.009631f
C29741 a_16375_45002# a_15861_45028# 0.029833f
C29742 a_8199_44636# a_8953_45002# 0.12099f
C29743 a_5937_45572# a_8191_45002# 0.180306f
C29744 a_17715_44484# a_413_45260# 4.56e-21
C29745 a_n2497_47436# a_1241_43940# 5.31e-20
C29746 a_12549_44172# a_3422_30871# 0.148646f
C29747 a_13747_46662# a_20679_44626# 0.030878f
C29748 a_n3690_38528# a_n4209_38216# 2.69e-19
C29749 a_n4209_38502# a_n3690_38304# 2.69e-19
C29750 a_n3420_38528# a_n3607_38528# 0.001534f
C29751 a_5934_30871# C10_N_btm 1.89e-19
C29752 a_7174_31319# a_3726_37500# 0.002891f
C29753 a_15507_47210# a_15673_47210# 0.81159f
C29754 a_n2497_47436# a_768_44030# 0.023758f
C29755 a_n1741_47186# a_11117_47542# 2.77e-19
C29756 a_n237_47217# a_n881_46662# 0.958566f
C29757 a_n23_47502# a_n1613_43370# 5.76e-20
C29758 a_2905_45572# a_2747_46873# 0.010677f
C29759 a_2124_47436# a_2266_47243# 0.005572f
C29760 a_n4315_30879# a_n4334_37440# 2.61e-19
C29761 a_6545_47178# a_4883_46098# 0.008688f
C29762 a_18214_42558# CAL_N 3.01e-20
C29763 a_12861_44030# a_16588_47582# 9.72e-20
C29764 a_13717_47436# a_17591_47464# 3.4e-19
C29765 a_n1435_47204# a_10227_46804# 0.004624f
C29766 a_5742_30871# C4_P_btm 0.03103f
C29767 a_14955_47212# a_16327_47482# 1.03e-19
C29768 a_11599_46634# a_16241_47178# 2.85e-20
C29769 a_6123_31319# VDD 0.532709f
C29770 a_5013_44260# a_5649_42852# 1.41e-20
C29771 a_n4318_40392# a_n4318_37592# 0.023213f
C29772 a_n1699_43638# a_n1821_43396# 3.16e-19
C29773 a_n447_43370# a_104_43370# 5.86e-20
C29774 a_6671_43940# a_6765_43638# 2.18e-19
C29775 a_21115_43940# a_10341_43396# 1.36e-20
C29776 a_14021_43940# a_8685_43396# 0.002318f
C29777 a_11967_42832# a_12089_42308# 0.022254f
C29778 a_10555_44260# a_10695_43548# 2.11e-20
C29779 a_15493_43940# a_15095_43370# 0.001144f
C29780 a_n984_44318# a_n1076_43230# 6.38e-21
C29781 a_4099_45572# a_n2661_43370# 0.002135f
C29782 a_8049_45260# a_14539_43914# 1.59e-36
C29783 a_2324_44458# a_14815_43914# 1.05e-20
C29784 a_11688_45572# a_3232_43370# 2.05e-19
C29785 a_15227_44166# a_17973_43940# 4.09e-19
C29786 a_n971_45724# a_685_42968# 4.15e-21
C29787 a_15143_45578# a_14797_45144# 0.001287f
C29788 a_10227_46804# a_15743_43084# 0.002448f
C29789 a_21363_45546# a_21188_45572# 0.233657f
C29790 a_20841_45814# a_20731_45938# 0.097745f
C29791 a_20623_45572# a_20528_45572# 0.049827f
C29792 a_3090_45724# a_19862_44208# 0.004983f
C29793 a_n1613_43370# a_9145_43396# 7e-20
C29794 a_n2293_46634# a_2896_43646# 7.64e-19
C29795 a_n1151_42308# a_n1991_42858# 2.39e-19
C29796 C4_P_btm C0_dummy_P_btm 0.113746f
C29797 C9_P_btm C3_N_btm 0.001271f
C29798 C7_P_btm C1_N_btm 4.76e-19
C29799 C6_P_btm C0_N_btm 2.8e-19
C29800 C5_P_btm C0_dummy_N_btm 1.24e-19
C29801 C2_P_btm C1_P_btm 5.0586f
C29802 C3_P_btm C0_P_btm 0.409996f
C29803 EN_VIN_BSTR_N C9_N_btm 0.226529f
C29804 a_22469_39537# VIN_N 2.79e-20
C29805 EN_VIN_BSTR_P VDD 0.917313f
C29806 a_n923_35174# RST_Z 0.001488f
C29807 a_12465_44636# a_19333_46634# 2.86e-20
C29808 a_4883_46098# a_19692_46634# 0.058277f
C29809 a_11599_46634# a_16721_46634# 0.00139f
C29810 a_15507_47210# a_16388_46812# 5.7e-19
C29811 a_1799_45572# a_2443_46660# 1.77e-19
C29812 a_n2661_46634# a_5275_47026# 0.003477f
C29813 a_n971_45724# a_n1991_46122# 0.010501f
C29814 a_n746_45260# a_n1853_46287# 3.3e-21
C29815 a_13381_47204# a_765_45546# 0.002617f
C29816 a_n743_46660# a_4955_46873# 0.0023f
C29817 a_n881_46662# a_8270_45546# 9.01e-20
C29818 a_n1925_46634# a_5385_46902# 0.003429f
C29819 a_5807_45002# a_8492_46660# 0.005311f
C29820 a_n2497_47436# a_1176_45822# 2.85e-20
C29821 a_15811_47375# a_13059_46348# 0.001466f
C29822 a_10227_46804# a_13885_46660# 6.78e-19
C29823 a_16547_43609# a_4361_42308# 9.06e-21
C29824 a_3626_43646# a_14543_43071# 4.05e-22
C29825 a_8791_43396# a_9127_43156# 0.007148f
C29826 a_n2661_42282# a_2351_42308# 8.86e-20
C29827 a_17324_43396# a_743_42282# 8.71e-21
C29828 a_16664_43396# a_16823_43084# 0.005264f
C29829 a_11967_42832# a_18907_42674# 4.8e-21
C29830 a_15743_43084# a_19177_43646# 4.34e-19
C29831 a_18525_43370# a_4190_30871# 0.005875f
C29832 a_11787_45002# a_11827_44484# 2.02e-20
C29833 a_8696_44636# a_13857_44734# 0.004972f
C29834 a_3429_45260# a_n2661_44458# 8.32e-19
C29835 a_n967_45348# a_n699_43396# 4.56e-20
C29836 a_327_44734# a_n1177_44458# 1.88e-21
C29837 a_1823_45246# a_2813_43396# 5.33e-20
C29838 a_13259_45724# a_11341_43940# 0.045479f
C29839 a_1307_43914# a_16922_45042# 1.8e-20
C29840 a_8199_44636# a_3626_43646# 0.001453f
C29841 a_4099_45572# a_2998_44172# 3.68e-22
C29842 a_n357_42282# a_n2661_42282# 0.055806f
C29843 a_n1059_45260# a_8701_44490# 4.94e-19
C29844 a_n2017_45002# a_5883_43914# 8.44e-20
C29845 a_n2312_40392# a_n2104_42282# 4.5e-20
C29846 a_n2312_39304# a_n4318_38216# 0.023429f
C29847 a_19692_46634# a_5649_42852# 0.01341f
C29848 a_17339_46660# a_15743_43084# 0.450316f
C29849 a_15227_44166# a_20731_47026# 1.96e-20
C29850 a_15227_46910# a_16388_46812# 1e-19
C29851 a_4883_46098# a_20692_30879# 9.38e-20
C29852 a_2107_46812# a_6945_45028# 0.028356f
C29853 a_n1925_46634# a_n1533_46116# 0.001581f
C29854 a_n1151_42308# a_7227_45028# 0.00514f
C29855 a_4791_45118# a_5907_45546# 0.02288f
C29856 a_n971_45724# a_7499_43078# 0.857375f
C29857 a_2063_45854# a_2211_45572# 0.006085f
C29858 a_19692_46634# a_21188_46660# 0.022017f
C29859 a_5257_43370# a_5497_46414# 0.002158f
C29860 a_9863_46634# a_3483_46348# 3.53e-22
C29861 a_17730_32519# C7_N_btm 1.47e-19
C29862 a_13678_32519# a_n784_42308# 0.009139f
C29863 a_14209_32519# COMP_P 7.77e-21
C29864 a_n2472_42826# a_n4318_38216# 0.006796f
C29865 a_2982_43646# a_13258_32519# 0.086314f
C29866 a_3626_43646# a_19511_42282# 0.182478f
C29867 a_n1853_43023# a_n3674_38680# 3.63e-19
C29868 a_10341_43396# a_10533_42308# 2.73e-21
C29869 a_743_42282# a_1184_42692# 0.005701f
C29870 a_19237_31679# C5_N_btm 1.11e-20
C29871 a_10157_44484# a_9313_44734# 0.026406f
C29872 a_16922_45042# a_18579_44172# 1.03e-19
C29873 a_6171_45002# a_11750_44172# 3.21e-19
C29874 a_5518_44484# a_5608_44484# 0.008441f
C29875 a_5343_44458# a_5708_44484# 0.048542f
C29876 a_949_44458# a_n2661_43922# 0.055363f
C29877 a_2779_44458# a_n2661_42834# 0.00388f
C29878 a_742_44458# a_n2293_43922# 1.56e-21
C29879 a_n2293_42834# a_n1549_44318# 7.42e-19
C29880 a_11691_44458# a_16241_44484# 2.22e-19
C29881 a_8191_45002# a_8333_44056# 4.8e-20
C29882 a_n357_42282# a_16823_43084# 0.016884f
C29883 a_20202_43084# a_20753_42852# 8.28e-19
C29884 SMPL_ON_P VDD 0.614138f
C29885 a_19431_45546# a_19319_43548# 2.72e-20
C29886 a_18494_42460# a_20159_44458# 0.024732f
C29887 a_21005_45260# a_11967_42832# 3.36e-20
C29888 a_19778_44110# a_20640_44752# 4.84e-20
C29889 a_11827_44484# a_17325_44484# 3.91e-19
C29890 a_7499_43078# a_8229_43396# 0.001513f
C29891 a_n2497_47436# DATA[0] 0.008757f
C29892 a_n1741_47186# RST_Z 7.39e-20
C29893 a_n2288_47178# CLK_DATA 6.87e-19
C29894 a_13747_46662# a_20528_45572# 2.86e-19
C29895 a_13675_47204# a_2437_43646# 6.63e-20
C29896 a_4883_46098# a_4927_45028# 2.86e-20
C29897 a_10227_46804# a_10775_45002# 0.006025f
C29898 a_584_46384# a_n2293_42834# 0.049322f
C29899 a_12861_44030# a_15595_45028# 0.012748f
C29900 a_n1613_43370# a_n1059_45260# 0.202724f
C29901 a_4704_46090# a_5066_45546# 0.002532f
C29902 a_n746_45260# a_n2661_43370# 0.060205f
C29903 a_8270_45546# a_8162_45546# 0.170838f
C29904 a_20916_46384# a_20107_45572# 6.04e-21
C29905 a_21188_46660# a_20692_30879# 3.94e-20
C29906 a_13759_46122# a_10809_44734# 6.06e-20
C29907 a_18189_46348# a_18819_46122# 1.04e-20
C29908 a_1067_42314# a_5932_42308# 4.34e-21
C29909 a_14097_32519# a_5742_30871# 0.004679f
C29910 a_2713_42308# a_3318_42354# 9.16e-19
C29911 a_n784_42308# a_6123_31319# 0.144274f
C29912 a_15597_42852# a_15803_42450# 1.45e-19
C29913 a_742_44458# a_n97_42460# 0.083982f
C29914 a_8035_47026# VDD 0.132317f
C29915 a_20193_45348# a_2982_43646# 4.86e-20
C29916 a_n2293_45010# a_685_42968# 1.26e-20
C29917 a_n2661_45010# a_1847_42826# 1.52e-22
C29918 a_n1059_45260# a_n1533_42852# 1.94e-19
C29919 a_13249_42308# a_13569_43230# 2.14e-19
C29920 a_n2661_43922# a_11341_43940# 3.15e-19
C29921 a_n699_43396# a_n1917_43396# 1.68e-20
C29922 a_10428_46928# CLK 0.032943f
C29923 a_n967_45348# a_n4318_38680# 1.38e-21
C29924 a_n755_45592# a_5379_42460# 0.038776f
C29925 a_n443_42852# a_1149_42558# 1.56e-19
C29926 a_11823_42460# a_15785_43172# 3.45e-20
C29927 a_14539_43914# a_15037_43940# 0.054182f
C29928 a_1307_43914# a_15743_43084# 1.61e-19
C29929 a_n984_44318# a_175_44278# 1.1e-19
C29930 a_167_45260# a_2437_43646# 0.025008f
C29931 a_2957_45546# a_3316_45546# 0.001625f
C29932 a_n1099_45572# a_n1013_45572# 0.00411f
C29933 a_8049_45260# a_12427_45724# 0.012343f
C29934 a_n2293_45546# a_2277_45546# 1.67e-19
C29935 a_n2661_45546# a_n310_45572# 1.2e-19
C29936 a_n971_45724# a_3600_43914# 1.64e-20
C29937 a_n1991_46122# a_n2293_45010# 4.53e-20
C29938 a_12465_44636# a_12553_44484# 3.52e-19
C29939 a_n863_45724# a_n443_42852# 0.556081f
C29940 a_n743_46660# a_12607_44458# 2.46e-22
C29941 a_1799_45572# a_949_44458# 4.76e-19
C29942 a_768_44030# a_6109_44484# 0.04198f
C29943 a_13059_46348# a_13556_45296# 0.274813f
C29944 a_584_46384# a_1115_44172# 0.174981f
C29945 a_21076_30879# en_comp 3.62e-19
C29946 a_n2293_46098# a_n1059_45260# 2.7e-19
C29947 a_n2157_46122# a_n2017_45002# 2.07e-20
C29948 a_n1613_43370# a_484_44484# 1.49e-20
C29949 a_10586_45546# a_8746_45002# 0.001538f
C29950 a_n1641_46494# a_n2661_45010# 2.26e-19
C29951 a_n755_45592# a_n23_45546# 0.001003f
C29952 a_997_45618# a_n356_45724# 2.02e-19
C29953 a_16327_47482# a_11967_42832# 0.241578f
C29954 a_n4064_40160# a_n4251_39616# 0.001069f
C29955 a_1606_42308# CAL_P 0.00911f
C29956 a_n784_42308# EN_VIN_BSTR_P 0.051272f
C29957 a_n971_45724# a_5129_47502# 3.14e-19
C29958 a_n237_47217# a_n443_46116# 0.110841f
C29959 a_2124_47436# a_n1151_42308# 0.006002f
C29960 a_2553_47502# a_2952_47436# 0.002785f
C29961 a_2063_45854# a_2905_45572# 0.037943f
C29962 a_n1741_47186# a_6851_47204# 0.030234f
C29963 a_584_46384# a_3160_47472# 2.16e-20
C29964 a_7174_31319# a_1239_39043# 7.77e-20
C29965 a_n3565_39590# a_n4064_39616# 0.231239f
C29966 a_5932_42308# a_3726_37500# 0.003378f
C29967 a_15597_42852# VDD 0.239357f
C29968 a_n1630_35242# a_n1838_35608# 0.00968f
C29969 a_n2661_42834# a_n13_43084# 6.03e-20
C29970 a_n2293_43922# a_n901_43156# 3.99e-20
C29971 a_6109_44484# a_5755_42852# 6.71e-22
C29972 a_1307_43914# a_1606_42308# 0.003969f
C29973 a_18579_44172# a_15743_43084# 0.003564f
C29974 a_n356_44636# a_10835_43094# 1.71e-20
C29975 a_n913_45002# a_14456_42282# 0.006851f
C29976 a_n2017_45002# a_13333_42558# 0.001525f
C29977 a_5111_44636# a_5934_30871# 6.55e-19
C29978 a_17517_44484# a_21487_43396# 9.64e-21
C29979 a_14673_44172# a_4361_42308# 5.89e-21
C29980 a_12549_44172# a_19808_44306# 6.88e-19
C29981 a_2324_44458# a_4743_44484# 0.042685f
C29982 a_n1613_43370# a_n2840_43370# 2.32e-21
C29983 a_n2293_45546# a_626_44172# 0.150062f
C29984 a_22959_46124# a_19721_31679# 5.11e-20
C29985 a_5263_45724# a_3537_45260# 3.44e-19
C29986 a_2711_45572# a_5147_45002# 0.003609f
C29987 a_5257_43370# a_5841_44260# 3.99e-19
C29988 a_n443_42852# a_8191_45002# 3.74e-21
C29989 a_4185_45028# a_n356_44636# 1.54308f
C29990 a_12741_44636# a_11649_44734# 3.54e-20
C29991 a_n2661_45546# a_2232_45348# 7.5e-19
C29992 a_6945_45028# a_n2661_44458# 1.65e-19
C29993 a_n863_45724# a_375_42282# 0.451905f
C29994 CAL_N a_22469_39537# 0.024229f
C29995 a_22521_40599# a_22821_38993# 0.002401f
C29996 a_22469_40625# a_22545_38993# 9.26e-21
C29997 a_8912_37509# CAL_P 0.007121f
C29998 a_22521_40055# a_22780_40081# 0.010228f
C29999 a_n881_46662# a_1123_46634# 0.004455f
C30000 a_n1435_47204# a_10467_46802# 1.8e-20
C30001 a_9313_45822# a_10249_46116# 1.36e-19
C30002 a_11031_47542# a_6755_46942# 0.001571f
C30003 a_n1613_43370# a_948_46660# 0.281392f
C30004 a_3754_39964# VDD 0.033808f
C30005 a_n4209_38216# VIN_P 0.029185f
C30006 a_13747_46662# a_19594_46812# 0.03826f
C30007 a_5807_45002# a_16750_47204# 5.29e-19
C30008 a_2747_46873# a_2443_46660# 0.129886f
C30009 a_4883_46098# a_3877_44458# 0.002191f
C30010 a_6151_47436# a_6903_46660# 4.55e-19
C30011 a_n1151_42308# a_11813_46116# 0.019835f
C30012 a_14021_43940# a_17333_42852# 4.57e-21
C30013 a_3080_42308# a_13678_32519# 0.002941f
C30014 a_2982_43646# a_20301_43646# 9.07e-21
C30015 a_9803_43646# a_10149_43396# 0.013377f
C30016 a_9145_43396# a_14537_43646# 0.003686f
C30017 a_n2293_43922# a_10533_42308# 4.97e-20
C30018 a_9313_44734# a_14113_42308# 4.32e-20
C30019 a_2437_43646# DATA[4] 0.060047f
C30020 a_n356_44636# a_16269_42308# 4.62e-19
C30021 a_3422_30871# a_n1630_35242# 0.828871f
C30022 a_17730_32519# COMP_P 1.26e-20
C30023 a_9885_43646# a_10341_43396# 0.001685f
C30024 a_n1917_43396# a_n4318_38680# 3.79e-19
C30025 a_n97_42460# a_n901_43156# 0.011039f
C30026 a_n1809_43762# a_n1991_42858# 9.16e-20
C30027 a_n1699_43638# a_n1736_43218# 1.6e-19
C30028 a_8685_43396# a_13943_43396# 5.42e-19
C30029 a_13661_43548# a_12379_42858# 1.34e-19
C30030 a_18189_46348# a_11341_43940# 2.49e-20
C30031 a_3483_46348# a_9801_43940# 0.027985f
C30032 a_9482_43914# a_13777_45326# 0.206086f
C30033 a_7499_43078# a_9313_44734# 0.0624f
C30034 a_9049_44484# a_9241_44734# 0.001498f
C30035 a_n357_42282# a_19279_43940# 3.11e-20
C30036 SMPL_ON_P a_n784_42308# 0.001291f
C30037 a_10775_45002# a_1307_43914# 2.5e-21
C30038 a_2274_45254# a_2448_45028# 5.85e-19
C30039 a_20107_45572# a_21101_45002# 0.001705f
C30040 a_20273_45572# a_21005_45260# 3.27e-19
C30041 a_4558_45348# a_5105_45348# 5.58e-20
C30042 a_5147_45002# a_4640_45348# 5.32e-21
C30043 a_n2109_45247# a_n2661_43370# 0.006863f
C30044 a_7276_45260# a_1423_45028# 2.13e-20
C30045 a_13159_45002# a_14537_43396# 3.64e-20
C30046 a_13017_45260# a_14797_45144# 1.84e-19
C30047 a_13348_45260# a_14180_45002# 5.21e-19
C30048 a_3090_45724# a_14579_43548# 0.074713f
C30049 a_11453_44696# a_6945_45028# 0.022389f
C30050 a_22731_47423# a_10809_44734# 0.005082f
C30051 a_10227_46804# a_526_44458# 5.93e-20
C30052 a_n2833_47464# a_n2956_38216# 1e-20
C30053 a_n2293_46634# a_1138_42852# 0.023262f
C30054 a_12469_46902# a_12816_46660# 0.051162f
C30055 a_n743_46660# a_376_46348# 0.076781f
C30056 a_n2438_43548# a_n1076_46494# 2.06e-20
C30057 a_n2661_46634# a_167_45260# 2.09e-19
C30058 a_n881_46662# a_13759_46122# 0.01582f
C30059 a_5275_47026# a_765_45546# 0.002883f
C30060 a_11309_47204# a_9290_44172# 4.41e-19
C30061 a_n1925_46634# a_805_46414# 9.66e-19
C30062 a_n2288_47178# a_n2661_45546# 1.03e-20
C30063 a_171_46873# a_n1641_46494# 5.78e-21
C30064 a_n13_43084# a_n2293_42282# 7.33e-21
C30065 a_3626_43646# a_4921_42308# 0.431551f
C30066 a_3539_42460# a_4933_42558# 6.41e-19
C30067 a_16137_43396# a_15597_42852# 4.88e-19
C30068 a_3080_42308# a_6123_31319# 1.45722f
C30069 a_10796_42968# a_10341_42308# 0.65943f
C30070 a_10991_42826# a_10922_42852# 0.209641f
C30071 a_10835_43094# a_12379_42858# 0.001706f
C30072 a_n1423_42826# a_n914_42852# 2.6e-19
C30073 a_n97_42460# a_10533_42308# 0.001168f
C30074 a_4185_45028# a_12379_42858# 6.62e-20
C30075 a_13661_43548# a_18727_42674# 1.61e-19
C30076 a_8696_44636# a_15493_43940# 1.53e-19
C30077 a_11823_42460# a_13565_43940# 0.046344f
C30078 a_n755_45592# a_7287_43370# 1.51e-19
C30079 a_16147_45260# a_15682_43940# 8.35e-19
C30080 a_n913_45002# a_895_43940# 3.46e-19
C30081 a_n1059_45260# a_2675_43914# 1.32e-21
C30082 a_n2017_45002# a_2889_44172# 1.5e-21
C30083 a_13259_45724# a_10341_43396# 0.08137f
C30084 a_n2661_45546# a_5565_43396# 7.68e-21
C30085 SMPL_ON_P a_n2302_37690# 3.04e-19
C30086 a_14537_43396# a_11967_42832# 7.01e-19
C30087 a_11691_44458# a_16979_44734# 0.12231f
C30088 a_11827_44484# a_18287_44626# 0.024541f
C30089 a_n2661_44458# a_8103_44636# 0.006972f
C30090 a_4646_46812# a_6123_31319# 0.004637f
C30091 a_5257_43370# a_5267_42460# 9.2e-19
C30092 a_8199_44636# a_8037_42858# 2.18e-20
C30093 a_8953_45546# a_7871_42858# 0.017048f
C30094 a_13507_46334# a_18341_45572# 7.32e-21
C30095 a_1799_45572# a_1990_45572# 2.88e-19
C30096 a_11415_45002# a_17957_46116# 4.92e-22
C30097 a_3483_46348# a_6165_46155# 1.15e-21
C30098 a_4704_46090# a_5068_46348# 5.06e-19
C30099 a_n971_45724# a_4558_45348# 1.27e-19
C30100 a_12991_46634# a_13259_45724# 6.17e-19
C30101 a_n1151_42308# a_n967_45348# 0.170453f
C30102 a_11459_47204# a_2437_43646# 0.004348f
C30103 a_18597_46090# a_18799_45938# 1.88e-19
C30104 a_11599_46634# a_20528_45572# 1.32e-20
C30105 a_765_45546# a_2981_46116# 3.97e-21
C30106 a_n237_47217# a_3537_45260# 3.39e-20
C30107 a_584_46384# a_413_45260# 0.164383f
C30108 a_n443_46116# a_n2017_45002# 1.32e-19
C30109 a_4791_45118# a_n1059_45260# 0.020789f
C30110 a_9863_47436# a_3357_43084# 1.35e-19
C30111 a_n881_46662# a_15297_45822# 0.001288f
C30112 a_12741_44636# a_17583_46090# 2.35e-20
C30113 a_n743_46660# a_8746_45002# 1.81e-19
C30114 a_16327_47482# a_20273_45572# 0.050306f
C30115 a_4883_46098# a_18175_45572# 6.22e-20
C30116 a_n3674_39304# a_n4334_39616# 4.04e-19
C30117 a_14401_32519# C9_N_btm 5.77e-20
C30118 a_17538_32519# C7_N_btm 8.17e-19
C30119 a_5534_30871# a_13657_42308# 9.47e-19
C30120 a_3080_42308# EN_VIN_BSTR_P 0.043903f
C30121 a_17701_42308# a_15959_42545# 1.03e-20
C30122 a_11823_42460# a_5534_30871# 0.511874f
C30123 a_n357_42282# a_11136_42852# 0.002171f
C30124 a_n2956_38680# a_5934_30871# 4.1e-21
C30125 a_4185_45028# a_18727_42674# 1.37e-19
C30126 a_n2438_43548# VDD 3.40589f
C30127 a_n2293_42834# a_n1177_43370# 0.007412f
C30128 a_1307_43914# a_3539_42460# 1.85e-19
C30129 a_n356_44636# a_1241_44260# 7.4e-20
C30130 a_11967_42832# a_20835_44721# 0.033569f
C30131 a_19615_44636# a_20679_44626# 1.02e-20
C30132 a_17517_44484# a_21398_44850# 0.01617f
C30133 a_n743_46660# RST_Z 1.57e-20
C30134 a_10193_42453# a_18083_42858# 0.037244f
C30135 a_n1925_42282# a_3905_42558# 8.24e-19
C30136 a_5891_43370# a_6453_43914# 3.53e-20
C30137 a_n2312_38680# CLK_DATA 1.56e-20
C30138 a_20159_44458# a_20640_44752# 0.042415f
C30139 a_n2661_43922# a_175_44278# 0.003068f
C30140 a_7640_43914# a_7542_44172# 0.20977f
C30141 a_n2293_43922# a_n984_44318# 4.06e-20
C30142 a_n2661_42834# a_644_44056# 0.005887f
C30143 en_comp a_12281_43396# 4.34e-21
C30144 a_5111_44636# a_7221_43396# 9.51e-19
C30145 a_n2661_46634# DATA[4] 7.86e-20
C30146 a_13249_42308# a_13113_42826# 0.008586f
C30147 a_10903_43370# a_10053_45546# 4.05e-19
C30148 a_11415_45002# a_16020_45572# 9.68e-19
C30149 a_4883_46098# a_10440_44484# 3.27e-21
C30150 a_3877_44458# a_3602_45348# 1.19e-19
C30151 a_10467_46802# a_10775_45002# 1.67e-22
C30152 a_19321_45002# a_19778_44110# 0.568668f
C30153 a_13747_46662# a_18494_42460# 0.004606f
C30154 a_765_45546# a_17568_45572# 2.41e-21
C30155 a_n1613_43370# a_n4318_40392# 4.23e-20
C30156 a_16327_47482# a_18989_43940# 0.100946f
C30157 a_11901_46660# a_413_45260# 4.96e-20
C30158 a_12741_44636# a_8696_44636# 2.20704f
C30159 a_8270_45546# a_3537_45260# 0.002418f
C30160 a_11189_46129# a_8746_45002# 6.97e-20
C30161 a_9290_44172# a_10490_45724# 0.022805f
C30162 a_11133_46155# a_10193_42453# 0.039441f
C30163 a_10428_46928# a_10951_45334# 1.28e-19
C30164 COMP_P VDAC_Pi 0.005217f
C30165 a_17303_42282# a_17531_42308# 0.04615f
C30166 a_5932_42308# a_1239_39043# 8.89e-20
C30167 a_4958_30871# a_18057_42282# 4.22e-19
C30168 a_17701_42308# RST_Z 1.77e-20
C30169 a_18083_42858# VDD 0.408512f
C30170 a_n2956_38216# a_n2302_37984# 0.041408f
C30171 a_n2017_45002# a_n4318_37592# 0.043579f
C30172 a_n2293_45010# a_n1329_42308# 1.37e-19
C30173 a_11133_46155# VDD 0.176249f
C30174 a_20365_43914# a_15493_43940# 0.048673f
C30175 a_20935_43940# a_11341_43940# 0.006081f
C30176 a_9313_44734# a_15781_43660# 0.00335f
C30177 a_n2661_43922# a_10341_43396# 1.08e-19
C30178 a_19963_31679# a_n1630_35242# 1.23e-19
C30179 a_13483_43940# a_14021_43940# 0.109097f
C30180 a_n2810_45028# a_n4318_38216# 0.023084f
C30181 en_comp a_n3674_38680# 0.014975f
C30182 a_n2956_37592# a_n2472_42282# 8.96e-21
C30183 a_14815_43914# a_14579_43548# 9.4e-21
C30184 a_2324_44458# a_8488_45348# 0.003185f
C30185 a_10586_45546# a_3232_43370# 8.27e-19
C30186 a_15227_44166# a_9313_44734# 0.06548f
C30187 a_n863_45724# a_2437_43646# 0.071802f
C30188 a_11453_44696# a_11173_44260# 3.43e-20
C30189 a_526_44458# a_1307_43914# 0.467539f
C30190 a_17339_46660# a_17970_44736# 0.002841f
C30191 a_n2442_46660# a_n3674_39768# 0.023663f
C30192 a_12549_44172# a_10729_43914# 4.26e-20
C30193 a_768_44030# a_10405_44172# 0.001056f
C30194 a_8746_45002# a_11136_45572# 1.91e-20
C30195 a_10490_45724# a_11064_45572# 0.001758f
C30196 a_10193_42453# a_11688_45572# 0.003765f
C30197 a_8049_45260# a_6709_45028# 4.7e-19
C30198 a_21613_42308# RST_Z 2.94e-19
C30199 a_n4064_39072# a_n923_35174# 0.007158f
C30200 a_n2109_47186# a_4817_46660# 0.028101f
C30201 a_n1151_42308# a_1110_47026# 1.25e-19
C30202 a_16327_47482# a_5807_45002# 0.451783f
C30203 a_16763_47508# a_16942_47570# 0.007399f
C30204 a_16023_47582# a_16131_47204# 0.057222f
C30205 a_4883_46098# a_8128_46384# 0.010382f
C30206 a_n443_46116# a_1123_46634# 8.72e-19
C30207 a_4700_47436# a_2107_46812# 3.8e-22
C30208 a_7903_47542# a_n1925_46634# 8.56e-21
C30209 a_7754_39300# a_3754_38470# 0.082848f
C30210 a_16588_47582# a_16697_47582# 0.007416f
C30211 a_11599_46634# a_19594_46812# 0.001035f
C30212 a_n3420_39616# C2_P_btm 2.28e-20
C30213 a_n4064_39616# C4_P_btm 6.79e-20
C30214 a_22775_42308# VDD 0.426018f
C30215 a_13717_47436# a_22612_30879# 0.00542f
C30216 a_11459_47204# a_n2661_46634# 1.65e-19
C30217 a_n971_45724# a_3686_47026# 1.68e-19
C30218 a_584_46384# a_2609_46660# 3.91e-19
C30219 a_2063_45854# a_2443_46660# 0.017518f
C30220 a_n1741_47186# a_4651_46660# 4.72e-20
C30221 a_6031_43396# a_6197_43396# 0.581047f
C30222 a_11967_42832# a_12991_43230# 0.004319f
C30223 a_9028_43914# a_7871_42858# 5.97e-19
C30224 a_14021_43940# a_13678_32519# 0.021333f
C30225 a_2982_43646# a_2437_43396# 1.82e-20
C30226 a_18494_42460# a_4958_30871# 5.63e-20
C30227 a_18184_42460# a_17303_42282# 0.027385f
C30228 a_12741_44636# a_20365_43914# 3.64e-19
C30229 a_6511_45714# a_5343_44458# 4.65e-21
C30230 a_13259_45724# a_n2293_43922# 2.67e-19
C30231 a_3357_43084# a_7229_43940# 6.23e-21
C30232 a_12549_44172# a_21487_43396# 2.13e-19
C30233 a_20202_43084# a_11341_43940# 0.033215f
C30234 a_n755_45592# a_n23_44458# 8.98e-19
C30235 a_n467_45028# a_n143_45144# 0.007343f
C30236 a_n2017_45002# a_3537_45260# 0.033622f
C30237 a_n913_45002# a_3065_45002# 0.225034f
C30238 a_2324_44458# a_1414_42308# 2.25e-19
C30239 a_11823_42460# a_11691_44458# 0.022559f
C30240 a_3877_44458# a_6682_46660# 0.002161f
C30241 a_4915_47217# a_13351_46090# 3.17e-21
C30242 a_13675_47204# a_765_45546# 7.69e-19
C30243 a_4817_46660# a_5841_46660# 2.36e-20
C30244 a_7715_46873# a_8145_46902# 2.33e-20
C30245 a_6151_47436# a_10903_43370# 6.84e-20
C30246 a_9313_45822# a_5937_45572# 0.137696f
C30247 a_n1435_47204# a_8016_46348# 1.14e-20
C30248 a_5732_46660# a_6755_46942# 1.39e-20
C30249 a_7411_46660# a_7927_46660# 0.105839f
C30250 a_17538_32519# COMP_P 1.11e-20
C30251 a_14955_43940# a_15486_42560# 2.71e-19
C30252 a_15682_43940# a_15051_42282# 2.71e-20
C30253 a_16409_43396# a_16795_42852# 0.010927f
C30254 a_16137_43396# a_18083_42858# 0.005524f
C30255 a_18114_32519# C8_N_btm 4.06e-19
C30256 a_19721_31679# C7_N_btm 1.43e-20
C30257 a_n2157_42858# a_n1736_43218# 0.089677f
C30258 a_n1853_43023# a_n4318_38680# 0.003325f
C30259 a_n1641_43230# a_n1076_43230# 7.99e-20
C30260 a_n1991_42858# a_n3674_39304# 0.002508f
C30261 a_n4318_39304# a_n3674_38216# 0.023484f
C30262 a_18450_45144# VDD 2.13e-19
C30263 a_8147_43396# a_8495_42852# 4.42e-20
C30264 a_3626_43646# a_13291_42460# 0.001564f
C30265 a_n2433_43396# a_n2104_42282# 1.29e-19
C30266 a_2809_45028# a_n699_43396# 4.51e-19
C30267 a_5205_44484# a_7640_43914# 2.61e-20
C30268 a_526_44458# a_9396_43370# 2.4e-19
C30269 a_11322_45546# a_10949_43914# 1.8e-20
C30270 a_20623_45572# a_20640_44752# 3.53e-20
C30271 a_20273_45572# a_20835_44721# 2.82e-20
C30272 a_22591_45572# a_17517_44484# 3.95e-20
C30273 a_1138_42852# a_743_42282# 8.9e-20
C30274 a_6171_45002# a_5891_43370# 9.58e-20
C30275 a_3232_43370# a_8238_44734# 2.65e-20
C30276 a_17023_45118# a_11827_44484# 3.5e-20
C30277 a_19778_44110# a_18184_42460# 0.119002f
C30278 a_n2312_38680# a_n1630_35242# 8.58e-19
C30279 a_10227_46804# a_16104_42674# 0.012196f
C30280 a_10193_42453# a_12429_44172# 9.75e-19
C30281 a_10490_45724# a_10807_43548# 2.96e-21
C30282 a_n37_45144# a_n2661_42834# 3.28e-21
C30283 a_n143_45144# a_n2661_43922# 2.71e-20
C30284 a_13259_45724# a_n97_42460# 0.182889f
C30285 a_7715_46873# a_5066_45546# 0.020181f
C30286 a_14976_45028# a_15015_46420# 0.012921f
C30287 a_3090_45724# a_14840_46494# 0.002524f
C30288 a_765_45546# a_167_45260# 0.276049f
C30289 a_22365_46825# a_20820_30879# 0.00309f
C30290 a_4883_46098# a_10053_45546# 0.008211f
C30291 a_10227_46804# a_13163_45724# 2.33e-19
C30292 a_n2293_46634# a_n2956_38216# 5.44e-19
C30293 a_n881_46662# a_4099_45572# 7.8e-20
C30294 a_20202_43084# a_22591_46660# 0.001634f
C30295 a_n1613_43370# a_5263_45724# 5.35e-21
C30296 a_13507_46334# a_10193_42453# 0.008059f
C30297 a_16327_47482# a_15143_45578# 8.76e-21
C30298 a_n2661_46634# a_n863_45724# 3.34e-20
C30299 a_n2312_38680# a_n2661_45546# 5.53e-19
C30300 a_3080_42308# a_3754_39964# 9.9e-20
C30301 a_12429_44172# VDD 0.169047f
C30302 a_5649_42852# a_15486_42560# 5.1e-20
C30303 a_5111_42852# a_5932_42308# 0.001025f
C30304 a_5755_42852# a_6171_42473# 2.22e-19
C30305 a_4361_42308# a_15959_42545# 0.008092f
C30306 a_20990_47178# START 4.18e-19
C30307 a_4185_45028# a_3823_42558# 1.01e-19
C30308 a_21177_47436# RST_Z 5.48e-20
C30309 a_n2661_43922# a_n2293_43922# 0.05908f
C30310 a_18248_44752# a_18245_44484# 2.36e-20
C30311 a_20894_47436# SINGLE_ENDED 0.044283f
C30312 a_2437_43646# a_3540_43646# 1.24e-19
C30313 a_n467_45028# a_n97_42460# 5.34e-19
C30314 a_n356_44636# a_11967_42832# 0.025796f
C30315 a_n1059_45260# a_1209_43370# 8.19e-20
C30316 a_n357_42282# a_12545_42858# 0.042417f
C30317 a_n443_42852# a_7765_42852# 0.004527f
C30318 a_13507_46334# VDD 1.4135f
C30319 a_10227_46804# DATA[5] 2.13e-20
C30320 a_1307_43914# a_3353_43940# 0.005743f
C30321 a_17957_46116# a_13259_45724# 0.011559f
C30322 a_10809_44734# a_12379_46436# 0.011204f
C30323 a_18189_46348# a_18147_46436# 9.33e-19
C30324 a_5807_45002# a_14537_43396# 0.001298f
C30325 a_13661_43548# a_14180_45002# 1.37e-19
C30326 a_n743_46660# a_3232_43370# 7.45e-20
C30327 a_479_46660# a_413_45260# 2.29e-20
C30328 a_2063_45854# a_949_44458# 9.64e-19
C30329 a_584_46384# a_2779_44458# 2.06e-20
C30330 a_n1151_42308# a_n1917_44484# 2.05e-19
C30331 a_3090_45724# a_16115_45572# 0.00765f
C30332 a_15368_46634# a_15765_45572# 3.33e-19
C30333 a_n881_46662# a_5365_45348# 2.78e-19
C30334 a_16327_47482# a_18315_45260# 4.78e-19
C30335 a_13747_46662# a_13777_45326# 1.16e-21
C30336 a_167_45260# a_509_45822# 2.36e-20
C30337 a_5907_46634# a_3357_43084# 0.013466f
C30338 a_12861_44030# a_21359_45002# 1.13e-20
C30339 a_17583_46090# a_16375_45002# 4.13e-20
C30340 a_14840_46494# a_15002_46116# 0.006453f
C30341 a_10227_46804# a_16501_45348# 4.16e-20
C30342 a_2107_46812# a_3065_45002# 2.48e-20
C30343 a_n2293_46098# a_5263_45724# 0.002594f
C30344 a_1823_45246# a_1609_45822# 0.35471f
C30345 a_17364_32525# C4_N_btm 1.7e-20
C30346 a_21855_43396# VDD 0.289066f
C30347 a_14209_32519# C6_N_btm 0.001467f
C30348 a_10545_42558# a_10723_42308# 5.98e-20
C30349 a_n1630_35242# a_7174_31319# 0.035143f
C30350 COMP_P a_22465_38105# 0.059345f
C30351 a_n3674_38216# a_n4334_40480# 8.37e-20
C30352 a_4361_42308# RST_Z 4.9e-19
C30353 a_2711_45572# a_14113_42308# 5.51e-20
C30354 a_10440_44484# a_8685_43396# 2.31e-20
C30355 a_20623_46660# VDD 0.194217f
C30356 a_20841_46902# RST_Z 1.47e-20
C30357 a_765_45546# DATA[4] 0.006502f
C30358 a_7499_43078# a_8515_42308# 1.55e-19
C30359 a_n913_45002# a_2987_42968# 1.92e-21
C30360 a_11691_44458# a_18429_43548# 1.12e-20
C30361 a_n2293_42834# a_n1991_42858# 0.02898f
C30362 a_413_45260# a_22959_42860# 7.98e-20
C30363 a_n357_42282# a_19332_42282# 1.1e-19
C30364 a_11827_44484# a_19268_43646# 1.65e-20
C30365 a_n2661_42834# a_104_43370# 0.001459f
C30366 a_n2661_43922# a_n97_42460# 6.42e-20
C30367 a_2063_45854# a_11341_43940# 0.001102f
C30368 a_2711_45572# a_7499_43078# 0.007939f
C30369 a_3483_46348# a_14797_45144# 2.2e-21
C30370 a_11189_46129# a_3232_43370# 3.91e-20
C30371 a_9290_44172# a_6171_45002# 0.028032f
C30372 a_10903_43370# a_5111_44636# 3.25e-20
C30373 a_13259_45724# a_16020_45572# 0.024851f
C30374 a_19466_46812# a_19929_45028# 0.012303f
C30375 a_n443_42852# a_11823_42460# 0.356965f
C30376 a_1138_42852# a_626_44172# 0.010739f
C30377 a_1176_45822# a_1145_45348# 5.36e-22
C30378 a_6511_45714# a_4880_45572# 8.15e-21
C30379 a_6472_45840# a_6428_45938# 1.46e-19
C30380 a_8049_45260# a_18799_45938# 0.004297f
C30381 a_13747_46662# a_20640_44752# 0.027627f
C30382 a_5937_45572# a_7705_45326# 0.070066f
C30383 a_16375_45002# a_8696_44636# 0.043034f
C30384 a_17583_46090# a_413_45260# 1.29e-21
C30385 a_8199_44636# a_8191_45002# 0.234072f
C30386 a_19321_45002# a_20159_44458# 0.065041f
C30387 a_5257_43370# a_n356_44636# 1.18e-20
C30388 a_6755_46942# a_16112_44458# 0.023983f
C30389 a_8270_45546# a_8701_44490# 0.015888f
C30390 a_n4334_38528# a_n4334_38304# 0.052468f
C30391 a_n3565_38502# a_n4209_38216# 5.84657f
C30392 a_n4209_38502# a_n3565_38216# 0.028468f
C30393 a_n2302_38778# a_n2216_38778# 0.011479f
C30394 a_n3690_38528# a_n3607_38528# 0.007692f
C30395 a_n3420_38528# a_n4251_38528# 0.001487f
C30396 a_5934_30871# C9_N_btm 1.37e-19
C30397 a_15507_47210# a_15811_47375# 0.170975f
C30398 a_11599_46634# a_15673_47210# 0.012504f
C30399 a_n1741_47186# a_10037_47542# 4.61e-19
C30400 a_n746_45260# a_n881_46662# 0.190303f
C30401 a_n971_45724# a_7989_47542# 1.99e-19
C30402 a_n237_47217# a_n1613_43370# 0.034341f
C30403 a_2952_47436# a_2747_46873# 0.078913f
C30404 a_n4315_30879# a_n4209_37414# 0.039099f
C30405 a_6151_47436# a_4883_46098# 0.032223f
C30406 a_12861_44030# a_16763_47508# 0.008377f
C30407 a_19332_42282# CAL_N 0.001755f
C30408 a_13381_47204# a_10227_46804# 7.94e-20
C30409 a_13717_47436# a_16588_47582# 6.43e-20
C30410 a_5742_30871# C5_P_btm 0.089375f
C30411 a_7227_42308# VDD 0.296912f
C30412 a_n1761_44111# a_n1736_43218# 3.37e-20
C30413 a_n809_44244# a_n1076_43230# 1.8e-20
C30414 a_n984_44318# a_n901_43156# 2.43e-19
C30415 a_19721_31679# COMP_P 2.4e-20
C30416 a_5891_43370# a_8292_43218# 0.003655f
C30417 a_1307_43914# a_16104_42674# 4.76e-21
C30418 a_n2956_37592# a_n2216_39866# 1.2e-19
C30419 a_n1352_43396# a_104_43370# 4.33e-20
C30420 a_n1917_43396# a_n1809_43762# 0.057222f
C30421 a_n1699_43638# a_n1190_43762# 2.6e-19
C30422 a_n2267_43396# a_n1821_43396# 2.28e-19
C30423 a_n447_43370# a_n97_42460# 0.00228f
C30424 a_n2129_43609# a_n1655_43396# 0.002164f
C30425 a_20935_43940# a_10341_43396# 1.76e-20
C30426 a_11967_42832# a_12379_42858# 0.492977f
C30427 a_11341_43940# a_14955_43396# 1.96e-20
C30428 a_15493_43940# a_14205_43396# 2.04e-19
C30429 a_3090_45724# a_19478_44306# 0.027139f
C30430 a_10586_45546# a_8975_43940# 2.76e-20
C30431 a_15227_44166# a_17737_43940# 0.013191f
C30432 a_12861_44030# a_16823_43084# 6.87e-21
C30433 a_7227_45028# a_n2293_42834# 3.08e-20
C30434 a_13507_46334# a_16137_43396# 1.52e-19
C30435 a_8192_45572# a_8191_45002# 0.001292f
C30436 a_20273_45572# a_20731_45938# 0.034619f
C30437 a_20623_45572# a_21188_45572# 7.99e-20
C30438 a_n2293_46634# a_1987_43646# 5.42e-20
C30439 a_n1151_42308# a_n1853_43023# 0.021207f
C30440 a_768_44030# a_3457_43396# 3.04e-20
C30441 a_16327_47482# a_16867_43762# 0.012196f
C30442 a_15928_47570# a_6755_46942# 3.42e-19
C30443 a_12465_44636# a_15227_44166# 1.22e-19
C30444 a_4883_46098# a_19466_46812# 0.028345f
C30445 C5_P_btm C0_dummy_P_btm 0.11443f
C30446 C8_P_btm C1_N_btm 7.93e-19
C30447 C7_P_btm C0_N_btm 4.2e-19
C30448 C6_P_btm C0_dummy_N_btm 2.49e-19
C30449 a_11599_46634# a_16388_46812# 0.24092f
C30450 a_15507_47210# a_13059_46348# 2.35e-19
C30451 C3_P_btm C1_P_btm 7.40325f
C30452 C4_P_btm C0_P_btm 0.138884f
C30453 a_n743_46660# a_4651_46660# 9.85e-20
C30454 a_n2661_46634# a_5072_46660# 0.002463f
C30455 EN_VIN_BSTR_N C8_N_btm 0.090252f
C30456 a_n971_45724# a_n1853_46287# 0.08556f
C30457 a_11459_47204# a_765_45546# 0.005723f
C30458 a_21496_47436# a_19692_46634# 2.68e-21
C30459 a_1799_45572# a_n2661_46098# 0.003478f
C30460 a_948_46660# a_1057_46660# 0.007416f
C30461 a_1123_46634# a_1302_46660# 0.007399f
C30462 a_n923_35174# VDD 0.340432f
C30463 a_n237_47217# a_n2293_46098# 0.044593f
C30464 a_n881_46662# a_8189_46660# 5.68e-19
C30465 a_n1925_46634# a_4817_46660# 0.008055f
C30466 a_5807_45002# a_8667_46634# 0.008461f
C30467 a_n1741_47186# a_n1076_46494# 9.46e-21
C30468 a_15811_47375# a_15227_46910# 6.58e-19
C30469 a_10227_46804# a_13170_46660# 0.003988f
C30470 a_11453_44696# a_15559_46634# 1.71e-21
C30471 C10_P_btm C3_N_btm 0.002331f
C30472 a_n1613_43370# a_8270_45546# 9.43e-20
C30473 a_n2661_42282# a_2123_42473# 8.86e-20
C30474 a_16243_43396# a_4361_42308# 7.3e-20
C30475 a_2982_43646# a_5534_30871# 0.094381f
C30476 a_8791_43396# a_8387_43230# 5.36e-19
C30477 a_17499_43370# a_743_42282# 8.79e-20
C30478 a_104_43370# a_n2293_42282# 6.62e-21
C30479 a_18429_43548# a_4190_30871# 0.001307f
C30480 a_18783_43370# a_19177_43646# 2.23e-19
C30481 a_11967_42832# a_18727_42674# 1.83e-20
C30482 a_8696_44636# a_13468_44734# 0.001421f
C30483 a_n143_45144# a_n452_44636# 6.31e-21
C30484 a_3065_45002# a_n2661_44458# 0.027917f
C30485 a_16019_45002# a_16922_45042# 7.45e-20
C30486 a_n357_42282# a_6101_44260# 4.36e-20
C30487 a_n2312_40392# a_n4318_38216# 0.025276f
C30488 a_20202_43084# a_10341_43396# 0.037863f
C30489 a_19692_46634# a_13678_32519# 0.004218f
C30490 a_17339_46660# a_18783_43370# 0.02025f
C30491 a_n2312_39304# a_n2472_42282# 3.28e-20
C30492 a_3483_46348# a_7287_43370# 3.53e-21
C30493 a_n1059_45260# a_8103_44636# 8.03e-23
C30494 a_3175_45822# a_2998_44172# 1.76e-21
C30495 a_15227_46910# a_13059_46348# 0.043664f
C30496 a_15227_44166# a_20528_46660# 4.16e-21
C30497 a_5807_45002# a_6640_46482# 9.8e-19
C30498 a_n1741_47186# a_10193_42453# 6.98e-20
C30499 a_4883_46098# a_20205_31679# 3.29e-19
C30500 a_n1925_46634# a_n722_46482# 2.37e-19
C30501 a_n971_45724# a_8568_45546# 0.009964f
C30502 a_n1151_42308# a_6598_45938# 9.17e-20
C30503 a_4791_45118# a_5263_45724# 0.021183f
C30504 a_n443_46116# a_4099_45572# 1e-20
C30505 a_19692_46634# a_21363_46634# 0.00151f
C30506 a_5257_43370# a_5204_45822# 0.005904f
C30507 a_8492_46660# a_3483_46348# 1.74e-20
C30508 a_17730_32519# C6_N_btm 1.1e-19
C30509 a_10835_43094# a_12800_43218# 2.33e-21
C30510 a_10922_42852# a_11301_43218# 3.16e-19
C30511 a_10991_42826# a_11554_42852# 0.049827f
C30512 a_10796_42968# a_10752_42852# 1.46e-19
C30513 a_2982_43646# a_19647_42308# 0.002685f
C30514 a_3626_43646# a_18548_42308# 0.001059f
C30515 a_n2840_42826# a_n4318_38216# 0.012711f
C30516 a_n2472_42826# a_n2472_42282# 0.025171f
C30517 a_n2157_42858# a_n3674_38680# 2.17e-19
C30518 a_743_42282# a_1576_42282# 0.007548f
C30519 a_19237_31679# C4_N_btm 9.91e-21
C30520 a_n913_45002# a_10555_44260# 3.18e-21
C30521 a_9838_44484# a_9313_44734# 0.037628f
C30522 a_3232_43370# a_11750_44172# 0.020452f
C30523 a_6171_45002# a_10807_43548# 3.25e-20
C30524 a_20692_30879# a_13678_32519# 0.051702f
C30525 a_2711_45572# a_15781_43660# 1.33e-19
C30526 a_3090_45724# a_9223_42460# 1.31e-21
C30527 a_4743_44484# a_5708_44484# 1.11e-19
C30528 a_5343_44458# a_5608_44484# 0.004449f
C30529 a_742_44458# a_n2661_43922# 0.066714f
C30530 a_949_44458# a_n2661_42834# 0.009741f
C30531 a_11691_44458# a_15367_44484# 0.005161f
C30532 a_n2293_42834# a_n1331_43914# 4.35e-19
C30533 a_20202_43084# a_20356_42852# 0.003203f
C30534 a_n1741_47186# VDD 0.912651f
C30535 a_7499_43078# a_7466_43396# 1.63e-19
C30536 a_20820_30879# a_14097_32519# 0.052932f
C30537 a_n2497_47436# CLK_DATA 0.026654f
C30538 a_11827_44484# a_17061_44484# 0.001186f
C30539 a_19778_44110# a_20362_44736# 1.01e-19
C30540 a_20567_45036# a_11967_42832# 2.76e-20
C30541 a_18184_42460# a_20159_44458# 0.01449f
C30542 a_19321_45002# a_20623_45572# 0.001031f
C30543 a_21363_46634# a_20692_30879# 2.83e-19
C30544 a_13747_46662# a_21188_45572# 9.45e-19
C30545 a_13569_47204# a_2437_43646# 5.26e-20
C30546 a_4883_46098# a_5111_44636# 0.048482f
C30547 a_10227_46804# a_8953_45002# 0.017713f
C30548 a_13351_46090# a_10809_44734# 5.63e-20
C30549 a_5068_46348# a_5210_46482# 0.007833f
C30550 a_4791_45118# a_5837_45348# 1.43e-20
C30551 a_765_45546# a_n863_45724# 0.00497f
C30552 a_11415_45002# a_13259_45724# 0.505354f
C30553 a_n1613_43370# a_n2017_45002# 0.015448f
C30554 a_8016_46348# a_526_44458# 0.005011f
C30555 a_4419_46090# a_5066_45546# 8.55e-19
C30556 a_768_44030# a_3357_43084# 0.09747f
C30557 a_17715_44484# a_18819_46122# 1.03e-20
C30558 a_13925_46122# a_6945_45028# 3.29e-20
C30559 a_n971_45724# a_n2661_43370# 0.064346f
C30560 a_3090_45724# a_6511_45714# 1.98e-21
C30561 a_15227_44166# a_2711_45572# 0.113396f
C30562 a_8654_47026# a_7499_43078# 5.36e-21
C30563 a_18189_46348# a_17957_46116# 0.038851f
C30564 a_11599_46634# a_13777_45326# 8.08e-19
C30565 a_n1630_35242# a_5932_42308# 0.033914f
C30566 a_2713_42308# a_2903_42308# 0.23738f
C30567 a_196_42282# a_6123_31319# 1.36e-20
C30568 a_n784_42308# a_7227_42308# 3.86e-20
C30569 a_15597_42852# a_15764_42576# 9.51e-19
C30570 a_13291_42460# a_13921_42308# 2.04e-19
C30571 a_14539_43914# a_13565_43940# 4.14e-20
C30572 a_n452_44636# a_n97_42460# 4e-21
C30573 a_7832_46660# VDD 0.077608f
C30574 a_10467_46802# DATA[5] 1.05e-19
C30575 a_n2017_45002# a_n1533_42852# 0.004733f
C30576 a_n913_45002# a_n967_43230# 8.68e-20
C30577 a_3357_43084# a_5755_42852# 8.48e-20
C30578 a_n2661_42834# a_11341_43940# 0.007026f
C30579 a_n699_43396# a_n1699_43638# 1.54e-20
C30580 a_n2065_43946# a_453_43940# 2.55e-21
C30581 a_10150_46912# CLK 0.004688f
C30582 en_comp a_n4318_38680# 0.007648f
C30583 a_n357_42282# a_5379_42460# 0.007085f
C30584 a_n443_42852# a_961_42354# 0.002615f
C30585 a_n755_45592# a_5267_42460# 1.87e-19
C30586 a_11823_42460# a_14635_42282# 0.087526f
C30587 a_n467_45028# a_n901_43156# 4.74e-20
C30588 a_5111_44636# a_5649_42852# 0.121004f
C30589 a_n809_44244# a_175_44278# 0.001854f
C30590 a_15433_44458# a_15493_43396# 1.53e-19
C30591 a_12861_44030# a_19279_43940# 0.152657f
C30592 a_10227_46804# a_16335_44484# 4.36e-20
C30593 a_2957_45546# a_3218_45724# 0.063846f
C30594 a_n1099_45572# a_7_45899# 5.1e-20
C30595 a_8049_45260# a_11962_45724# 0.019556f
C30596 a_n2293_45546# a_1609_45822# 0.159696f
C30597 a_n971_45724# a_2998_44172# 2.34e-20
C30598 a_n1853_46287# a_n2293_45010# 2.07e-20
C30599 a_2202_46116# a_2437_43646# 0.022869f
C30600 a_2107_46812# a_6298_44484# 4.34e-21
C30601 a_1799_45572# a_742_44458# 1.46e-20
C30602 a_13059_46348# a_9482_43914# 0.448068f
C30603 a_n1151_42308# a_n1899_43946# 2.4e-19
C30604 a_584_46384# a_644_44056# 0.004876f
C30605 a_n2157_46122# a_n2109_45247# 1.34e-21
C30606 a_n2293_46098# a_n2017_45002# 1.65e-19
C30607 a_n755_45592# a_n356_45724# 0.016853f
C30608 a_n743_46660# a_8975_43940# 7.99e-22
C30609 a_17957_46116# a_17478_45572# 1.77e-19
C30610 a_10586_45546# a_10193_42453# 0.380236f
C30611 a_16327_47482# a_19006_44850# 0.028858f
C30612 a_14853_42852# VDD 0.004079f
C30613 COMP_P a_18194_35068# 5.47e-19
C30614 a_n4334_39616# a_n4064_39616# 0.4504f
C30615 a_n4209_39590# a_n2302_39866# 0.406459f
C30616 a_5934_30871# a_n3420_37440# 7.32e-19
C30617 a_n784_42308# a_n923_35174# 0.003268f
C30618 a_6123_31319# a_n4064_37440# 2.49e-19
C30619 a_n3690_39616# a_n3420_39616# 0.431154f
C30620 a_n3565_39590# a_n2946_39866# 0.406088f
C30621 a_n746_45260# a_n443_46116# 0.060788f
C30622 a_n971_45724# a_4915_47217# 0.017974f
C30623 a_1431_47204# a_n1151_42308# 0.013895f
C30624 a_n237_47217# a_4791_45118# 0.10712f
C30625 a_n1741_47186# a_6491_46660# 0.023524f
C30626 a_2063_45854# a_2952_47436# 2.96e-19
C30627 a_584_46384# a_2905_45572# 1.24e-20
C30628 a_19279_43940# a_19700_43370# 8.74e-21
C30629 a_n2661_42834# a_n1076_43230# 5.44e-20
C30630 a_n2661_43922# a_n901_43156# 9.27e-21
C30631 a_n2293_43922# a_n1641_43230# 9.84e-21
C30632 a_5111_44636# a_7963_42308# 5.33e-19
C30633 a_10586_45546# VDD 0.582083f
C30634 a_18579_44172# a_18783_43370# 1.04e-19
C30635 a_n356_44636# a_10518_42984# 1.13e-20
C30636 a_15004_44636# a_5342_30871# 5.64e-20
C30637 en_comp a_11551_42558# 4.34e-21
C30638 a_n913_45002# a_13575_42558# 3.5e-19
C30639 a_n1059_45260# a_14456_42282# 7.72e-20
C30640 a_n2017_45002# a_13249_42558# 0.001525f
C30641 a_14539_43914# a_5534_30871# 1.4e-20
C30642 a_2063_45854# a_10341_43396# 1e-19
C30643 a_12549_44172# a_18797_44260# 5.67e-19
C30644 a_11415_45002# a_n2661_43922# 2.28e-19
C30645 a_2324_44458# a_n699_43396# 0.070009f
C30646 a_9290_44172# a_12607_44458# 3.67e-20
C30647 a_4099_45572# a_3537_45260# 5.2e-19
C30648 a_2711_45572# a_4558_45348# 0.001943f
C30649 a_n2661_45546# a_1423_45028# 0.020024f
C30650 a_10227_46804# a_3626_43646# 0.011826f
C30651 a_22521_40055# a_22459_39145# 0.129251f
C30652 a_22521_40599# a_22545_38993# 6.99e-20
C30653 a_22469_40625# a_22521_39511# 0.65678f
C30654 CAL_N a_22821_38993# 2.99e-19
C30655 VDAC_N CAL_P 7.22e-21
C30656 a_n881_46662# a_383_46660# 0.001801f
C30657 a_n1435_47204# a_10428_46928# 1.94e-20
C30658 a_9313_45822# a_10554_47026# 3.34e-20
C30659 a_11031_47542# a_10249_46116# 0.003514f
C30660 a_n1613_43370# a_1123_46634# 0.358475f
C30661 a_n2216_37984# VDD 0.003985f
C30662 a_13661_43548# a_19594_46812# 0.003227f
C30663 a_13747_46662# a_19321_45002# 0.080725f
C30664 a_n4064_37440# EN_VIN_BSTR_P 0.031982f
C30665 a_768_44030# a_n2293_46634# 0.26984f
C30666 a_2747_46873# a_n2661_46098# 0.004275f
C30667 a_4791_45118# a_8270_45546# 0.001618f
C30668 a_n1151_42308# a_11735_46660# 0.050593f
C30669 a_14021_43940# a_18083_42858# 1.31e-20
C30670 a_20447_31679# RST_Z 0.050985f
C30671 a_2982_43646# a_4190_30871# 0.3223f
C30672 a_14955_43396# a_10341_43396# 0.01411f
C30673 a_9803_43646# a_9885_43396# 0.003935f
C30674 a_n356_44636# a_16197_42308# 1.9e-19
C30675 a_2437_43646# DATA[3] 0.075788f
C30676 a_4905_42826# a_4361_42308# 0.005834f
C30677 a_n2472_43914# a_n4318_38216# 4.52e-19
C30678 a_n1699_43638# a_n4318_38680# 1.98e-19
C30679 a_n1917_43396# a_n3674_39304# 1.1e-19
C30680 a_n97_42460# a_n1641_43230# 3.57e-21
C30681 a_n1809_43762# a_n1853_43023# 4.91e-20
C30682 a_n447_43370# a_n901_43156# 0.008716f
C30683 a_n1352_43396# a_n1076_43230# 9.05e-19
C30684 a_8685_43396# a_13837_43396# 6.31e-19
C30685 a_n2293_45010# a_n2661_43370# 0.067876f
C30686 a_n2293_46634# a_5755_42852# 4.15e-20
C30687 a_n971_45724# COMP_P 8.93e-21
C30688 a_17715_44484# a_11341_43940# 0.001541f
C30689 a_9482_43914# a_13556_45296# 0.726155f
C30690 a_8746_45002# a_5891_43370# 1.89e-19
C30691 a_17339_46660# a_3626_43646# 3.03e-20
C30692 a_12594_46348# a_12603_44260# 1e-20
C30693 a_8953_45002# a_1307_43914# 1.41e-19
C30694 a_20273_45572# a_20567_45036# 0.005333f
C30695 a_20107_45572# a_21005_45260# 2.5e-19
C30696 a_5205_44484# a_1423_45028# 0.821456f
C30697 a_4558_45348# a_4640_45348# 0.007001f
C30698 a_n967_45348# a_n2293_42834# 0.038042f
C30699 a_13017_45260# a_14537_43396# 0.003458f
C30700 a_3090_45724# a_13667_43396# 1.98e-20
C30701 a_10903_43370# a_13565_44260# 3.14e-19
C30702 a_n2497_47436# a_n1630_35242# 2.73e-20
C30703 a_12549_44172# a_15567_42826# 1.56e-19
C30704 a_11453_44696# a_21137_46414# 7.06e-21
C30705 a_n2293_46634# a_1176_45822# 0.001481f
C30706 a_6755_46942# a_12978_47026# 3.05e-19
C30707 a_11735_46660# a_14084_46812# 3.45e-21
C30708 a_11901_46660# a_12816_46660# 0.125324f
C30709 a_22223_47212# a_10809_44734# 0.009267f
C30710 a_n743_46660# a_n1076_46494# 0.001766f
C30711 a_n2438_43548# a_n901_46420# 5.58e-20
C30712 a_1123_46634# a_n2293_46098# 4.36e-20
C30713 a_n881_46662# a_13351_46090# 5.07e-21
C30714 a_5072_46660# a_765_45546# 0.001239f
C30715 a_n1925_46634# a_472_46348# 0.002778f
C30716 a_n2497_47436# a_n2661_45546# 0.030609f
C30717 a_171_46873# a_n1423_46090# 1.51e-20
C30718 a_5649_42852# a_5837_43172# 1.5e-19
C30719 a_n1076_43230# a_n2293_42282# 3.1e-20
C30720 a_14021_43940# a_22775_42308# 1.94e-20
C30721 a_3539_42460# a_3905_42558# 0.015463f
C30722 a_4905_42826# a_6761_42308# 3.95e-20
C30723 a_10796_42968# a_10922_42852# 0.170059f
C30724 a_10835_43094# a_10341_42308# 0.541777f
C30725 a_n1991_42858# a_n914_42852# 1.46e-19
C30726 a_n1853_43023# a_133_42852# 0.001685f
C30727 a_4185_45028# a_10341_42308# 1.48e-20
C30728 a_15861_45028# a_11341_43940# 3.78e-20
C30729 a_n755_45592# a_6547_43396# 7.25e-21
C30730 a_n357_42282# a_7287_43370# 0.002031f
C30731 a_n2017_45002# a_2675_43914# 5.66e-22
C30732 a_n913_45002# a_2479_44172# 0.003813f
C30733 a_n1059_45260# a_895_43940# 2.25e-19
C30734 a_n2661_45546# a_4181_43396# 0.009936f
C30735 SMPL_ON_P a_n4064_37440# 6.21e-20
C30736 a_n443_42852# a_2982_43646# 0.037773f
C30737 a_11691_44458# a_14539_43914# 0.268287f
C30738 a_11827_44484# a_18248_44752# 0.00953f
C30739 a_n2661_43370# a_9313_44734# 3.03e-20
C30740 a_1307_43914# a_16335_44484# 8.63e-20
C30741 a_n2661_44458# a_6298_44484# 0.025865f
C30742 a_12549_44172# a_20712_42282# 3.18e-19
C30743 a_4646_46812# a_7227_42308# 1.62e-20
C30744 a_8199_44636# a_7765_42852# 1.98e-19
C30745 a_13507_46334# a_18479_45785# 8.2e-20
C30746 a_11415_45002# a_18189_46348# 0.028334f
C30747 a_4185_45028# a_5164_46348# 1.41e-19
C30748 a_3483_46348# a_5497_46414# 8.7e-21
C30749 a_4419_46090# a_5068_46348# 5.78e-21
C30750 a_20731_47026# a_10809_44734# 0.003685f
C30751 a_n1151_42308# en_comp 8.03e-21
C30752 a_9313_45822# a_2437_43646# 0.045826f
C30753 a_18597_46090# a_18596_45572# 8.84e-19
C30754 a_19386_47436# a_19256_45572# 6.77e-21
C30755 a_n2661_46634# a_11823_42460# 0.331717f
C30756 a_n2109_47186# a_6171_45002# 1.79e-19
C30757 a_765_45546# a_1431_46436# 4.27e-19
C30758 a_1823_45246# a_5937_45572# 3.25e-20
C30759 a_584_46384# a_n37_45144# 9.32e-20
C30760 a_4791_45118# a_n2017_45002# 0.023951f
C30761 a_9067_47204# a_3357_43084# 5.7e-19
C30762 a_n237_47217# a_3429_45260# 7.06e-21
C30763 a_12741_44636# a_15682_46116# 3.17e-20
C30764 a_n743_46660# a_10193_42453# 0.25279f
C30765 a_16327_47482# a_20107_45572# 0.674639f
C30766 a_18780_47178# a_18799_45938# 9.94e-22
C30767 a_n3674_39304# a_n4209_39590# 4.47e-20
C30768 a_14401_32519# C8_N_btm 8.3e-20
C30769 a_17538_32519# C6_N_btm 5.51e-20
C30770 a_5534_30871# a_11897_42308# 4.24e-20
C30771 a_3080_42308# a_n923_35174# 0.006061f
C30772 a_22400_42852# a_22765_42852# 9.38e-19
C30773 a_17701_42308# a_15803_42450# 2.65e-20
C30774 a_11823_42460# a_14543_43071# 0.028488f
C30775 a_n2956_39304# a_5934_30871# 5.05e-21
C30776 a_4185_45028# a_18057_42282# 7.92e-20
C30777 a_n743_46660# VDD 1.75634f
C30778 a_n2293_42834# a_n1917_43396# 0.006976f
C30779 a_1307_43914# a_3626_43646# 0.012223f
C30780 a_11967_42832# a_20679_44626# 0.863531f
C30781 a_17517_44484# a_20980_44850# 0.026284f
C30782 a_8953_45002# a_9396_43370# 6.95e-20
C30783 a_10193_42453# a_17701_42308# 5.98e-19
C30784 a_526_44458# a_3905_42558# 0.006254f
C30785 a_5891_43370# a_5663_43940# 1.27e-19
C30786 a_20159_44458# a_20362_44736# 0.233657f
C30787 a_n2661_43922# a_n984_44318# 0.004148f
C30788 a_n2661_42834# a_175_44278# 0.010875f
C30789 a_8975_43940# a_11750_44172# 1.78e-19
C30790 a_7640_43914# a_7281_43914# 0.003713f
C30791 a_n2293_43922# a_n809_44244# 4.38e-21
C30792 a_6109_44484# a_7542_44172# 2.12e-20
C30793 a_n2661_46634# DATA[3] 5.46e-21
C30794 a_22612_30879# EN_OFFSET_CAL 0.118817f
C30795 a_3537_45260# a_8317_43396# 7.25e-21
C30796 a_5111_44636# a_8685_43396# 0.078598f
C30797 a_13249_42308# a_12545_42858# 0.030353f
C30798 a_8199_44636# a_11823_42460# 0.00368f
C30799 a_4915_47217# a_9313_44734# 1.84e-22
C30800 a_11415_45002# a_17478_45572# 0.002665f
C30801 a_n1613_43370# a_n2840_44458# 1.2e-19
C30802 a_4883_46098# a_10334_44484# 3.73e-21
C30803 a_3877_44458# a_3495_45348# 1.26e-19
C30804 a_10903_43370# a_9049_44484# 2.44e-20
C30805 a_10428_46928# a_10775_45002# 2.17e-22
C30806 a_19321_45002# a_18911_45144# 0.050257f
C30807 a_6755_46942# a_7229_43940# 6.9e-21
C30808 a_13747_46662# a_18184_42460# 0.123281f
C30809 a_13661_43548# a_18494_42460# 0.049953f
C30810 a_11813_46116# a_413_45260# 1.63e-20
C30811 a_12741_44636# a_16680_45572# 5.61e-19
C30812 a_3483_46348# a_9241_45822# 3e-19
C30813 a_10355_46116# a_10490_45724# 0.01084f
C30814 a_9290_44172# a_8746_45002# 0.004141f
C30815 a_11189_46129# a_10193_42453# 0.123385f
C30816 a_16327_47482# a_18374_44850# 0.16003f
C30817 a_5742_30871# a_n4209_39590# 1.2e-21
C30818 a_4958_30871# a_17531_42308# 0.192941f
C30819 a_17595_43084# RST_Z 2.39e-21
C30820 a_17701_42308# VDD 0.243354f
C30821 a_5934_30871# a_n3565_39304# 5.05e-21
C30822 a_n2956_38216# a_n4064_37984# 0.054267f
C30823 a_n2810_45028# a_n2472_42282# 9.69e-21
C30824 a_11189_46129# VDD 0.944289f
C30825 a_18287_44626# a_16823_43084# 9.2e-20
C30826 a_n452_44636# a_n901_43156# 6.5e-20
C30827 a_20269_44172# a_15493_43940# 0.051355f
C30828 a_20935_43940# a_21115_43940# 0.185422f
C30829 a_20623_43914# a_11341_43940# 0.007271f
C30830 a_9313_44734# a_15681_43442# 0.001424f
C30831 a_n2661_42834# a_10341_43396# 2.59e-19
C30832 a_10193_42453# a_21613_42308# 1.95e-19
C30833 a_n2017_45002# a_n1736_42282# 0.017988f
C30834 a_13483_43940# a_13829_44260# 0.013377f
C30835 a_n1899_43946# a_n1809_43762# 8.11e-19
C30836 a_n809_44244# a_n97_42460# 3.09e-19
C30837 a_n2810_45572# a_n3607_38304# 5.7e-20
C30838 en_comp a_n2840_42282# 0.001493f
C30839 a_n2956_37592# a_n3674_38680# 0.02294f
C30840 a_14539_43914# a_4190_30871# 8.06e-21
C30841 a_2711_45572# a_16377_45572# 4.3e-19
C30842 a_13507_46334# a_14021_43940# 0.01995f
C30843 a_2324_44458# a_8137_45348# 4.79e-19
C30844 a_584_46384# a_104_43370# 0.001171f
C30845 a_n2497_47436# a_1427_43646# 8.12e-20
C30846 a_17339_46660# a_17767_44458# 9.16e-19
C30847 a_4185_45028# a_18494_42460# 2.49e-19
C30848 a_n2442_46660# a_n4318_39768# 0.023739f
C30849 a_768_44030# a_9672_43914# 0.006402f
C30850 a_n2293_46634# a_7845_44172# 3.2e-20
C30851 a_8746_45002# a_11064_45572# 9.37e-21
C30852 a_10490_45724# a_10544_45572# 0.004398f
C30853 a_8049_45260# a_7229_43940# 0.014199f
C30854 a_11599_46634# a_19321_45002# 0.091019f
C30855 a_21887_42336# RST_Z 1.97e-20
C30856 a_n4064_39072# a_n1532_35090# 9.45e-20
C30857 a_n3420_39072# EN_VIN_BSTR_P 0.772414f
C30858 a_n2109_47186# a_4955_46873# 0.001032f
C30859 a_2063_45854# a_n2661_46098# 0.021195f
C30860 a_n1151_42308# a_n935_46688# 0.001606f
C30861 a_6491_46660# a_n743_46660# 4.83e-21
C30862 a_16327_47482# a_16131_47204# 0.016621f
C30863 a_16241_47178# a_5807_45002# 0.002482f
C30864 a_4007_47204# a_2107_46812# 7.24e-20
C30865 a_n443_46116# a_383_46660# 0.001079f
C30866 a_7227_47204# a_n1925_46634# 1.2e-19
C30867 a_7754_39632# a_8530_39574# 1.05e-19
C30868 a_3754_39134# VDAC_Ni 0.00194f
C30869 a_10227_46804# a_13675_47204# 1.49e-19
C30870 a_n4064_39616# C5_P_btm 8.54e-20
C30871 a_n3420_39616# C3_P_btm 2.76e-20
C30872 a_21613_42308# VDD 0.273985f
C30873 a_13717_47436# a_21588_30879# 0.052863f
C30874 a_9313_45822# a_n2661_46634# 0.032598f
C30875 a_584_46384# a_2443_46660# 0.004099f
C30876 a_n1741_47186# a_4646_46812# 1.57e-19
C30877 a_11967_42832# a_12800_43218# 0.025258f
C30878 a_11136_45572# VDD 0.004463f
C30879 a_10907_45822# CLK 0.035046f
C30880 a_8333_44056# a_7871_42858# 5.27e-20
C30881 a_5343_44458# a_8791_42308# 3.69e-19
C30882 a_n97_42460# a_14955_43396# 2e-20
C30883 a_14021_43940# a_21855_43396# 0.025748f
C30884 a_6031_43396# a_6293_42852# 0.163953f
C30885 a_3626_43646# a_9396_43370# 2.73e-20
C30886 a_18184_42460# a_4958_30871# 0.004748f
C30887 a_12741_44636# a_20269_44172# 3.52e-20
C30888 a_n443_42852# a_14539_43914# 7.29e-19
C30889 a_n967_45348# a_413_45260# 9.61e-20
C30890 a_10227_46804# a_8037_42858# 1.91e-20
C30891 a_22612_30879# a_15743_43084# 4.17e-20
C30892 a_12861_44030# a_12545_42858# 1.63e-20
C30893 a_20202_43084# a_21115_43940# 1.71e-19
C30894 a_n755_45592# a_n356_44636# 2.42652f
C30895 a_n357_42282# a_n23_44458# 4.49e-20
C30896 a_768_44030# a_743_42282# 1.92e-19
C30897 a_12549_44172# a_20556_43646# 0.125209f
C30898 a_n1059_45260# a_3065_45002# 0.023485f
C30899 a_12427_45724# a_11691_44458# 3.08e-21
C30900 a_4646_46812# a_7832_46660# 3.69e-20
C30901 a_4915_47217# a_12594_46348# 3.27e-20
C30902 a_13569_47204# a_765_45546# 7.71e-19
C30903 a_16327_47482# a_3483_46348# 0.003076f
C30904 a_7715_46873# a_7577_46660# 0.205227f
C30905 a_4817_46660# a_6999_46987# 1.63e-20
C30906 a_9313_45822# a_8199_44636# 0.015956f
C30907 a_12549_44172# a_19551_46910# 1.88e-19
C30908 a_13661_43548# a_16388_46812# 2.4e-20
C30909 a_13747_46662# a_13059_46348# 0.273684f
C30910 a_5807_45002# a_16721_46634# 0.112018f
C30911 a_n1151_42308# a_2324_44458# 0.075066f
C30912 a_5257_43370# a_7927_46660# 7.79e-22
C30913 a_5907_46634# a_6755_46942# 5.62e-20
C30914 a_7411_46660# a_8145_46902# 0.053385f
C30915 a_n237_47217# a_6945_45028# 0.072758f
C30916 a_n2497_47436# a_n1533_46116# 0.006317f
C30917 a_14955_43940# a_15051_42282# 1.74e-20
C30918 a_15682_43940# a_14113_42308# 2.3e-19
C30919 a_16409_43396# a_16414_43172# 4.62e-21
C30920 a_743_42282# a_5755_42852# 2.61e-20
C30921 a_16137_43396# a_17701_42308# 0.025497f
C30922 a_16547_43609# a_16795_42852# 0.081093f
C30923 a_18114_32519# C7_N_btm 2.94e-19
C30924 a_19721_31679# C6_N_btm 1.26e-20
C30925 a_n2157_42858# a_n4318_38680# 9.64e-19
C30926 a_n1853_43023# a_n3674_39304# 1.5e-19
C30927 a_n1423_42826# a_n1076_43230# 0.051162f
C30928 a_2982_43646# a_14635_42282# 3.39e-19
C30929 a_n2433_43396# a_n4318_38216# 0.002497f
C30930 SMPL_ON_P a_n3420_39072# 1.03e-20
C30931 a_5205_44484# a_6109_44484# 0.029986f
C30932 a_526_44458# a_8791_43396# 1.78e-20
C30933 a_2382_45260# a_3363_44484# 9.62e-20
C30934 a_11322_45546# a_10729_43914# 3.04e-19
C30935 a_20273_45572# a_20679_44626# 3.84e-19
C30936 a_20107_45572# a_20835_44721# 6.77e-20
C30937 a_3357_43084# a_17517_44484# 0.001645f
C30938 a_17715_44484# a_10341_43396# 1.37e-19
C30939 a_6171_45002# a_8375_44464# 4.23e-20
C30940 a_3232_43370# a_5891_43370# 0.137859f
C30941 a_16922_45042# a_11827_44484# 0.032223f
C30942 a_10193_42453# a_11750_44172# 0.01114f
C30943 a_n467_45028# a_n2661_43922# 0.024697f
C30944 a_n143_45144# a_n2661_42834# 2.16e-21
C30945 a_8270_45546# a_6945_45028# 3.18e-19
C30946 a_n2293_46634# a_n2472_45546# 1.2e-19
C30947 a_15009_46634# a_14840_46494# 0.001393f
C30948 a_3090_45724# a_15015_46420# 0.019425f
C30949 a_4915_47217# a_15037_45618# 2.32e-22
C30950 a_9067_47204# a_9159_45572# 6.28e-22
C30951 a_7411_46660# a_5066_45546# 7.26e-20
C30952 a_5257_43370# a_6419_46482# 0.006417f
C30953 a_768_44030# a_2277_45546# 0.027945f
C30954 a_n2661_46634# a_n1079_45724# 4.39e-21
C30955 a_n2442_46660# a_n2956_38216# 0.048086f
C30956 a_765_45546# a_2202_46116# 4.62e-20
C30957 a_20202_43084# a_11415_45002# 0.041726f
C30958 a_n1613_43370# a_4099_45572# 1.78e-20
C30959 a_22365_46825# a_22591_46660# 0.08571f
C30960 a_4883_46098# a_9049_44484# 0.001404f
C30961 a_10227_46804# a_12791_45546# 1.59e-20
C30962 a_n2312_38680# a_n2810_45572# 0.062154f
C30963 a_11750_44172# VDD 0.131662f
C30964 a_5649_42852# a_15051_42282# 3.72e-19
C30965 a_5755_42852# a_5755_42308# 3.59e-19
C30966 a_16823_43084# a_17124_42282# 6.14e-21
C30967 a_4361_42308# a_15803_42450# 0.055869f
C30968 a_11301_43218# a_11554_42852# 4.61e-19
C30969 a_n443_42852# a_7871_42858# 0.013386f
C30970 a_21177_47436# VDD 0.179587f
C30971 a_20894_47436# START 1.67e-19
C30972 a_20990_47178# RST_Z 7.86e-20
C30973 a_18287_44626# a_19279_43940# 4.65e-20
C30974 a_18989_43940# a_20679_44626# 4.34e-21
C30975 a_n2661_42834# a_n2293_43922# 0.034793f
C30976 a_17970_44736# a_18245_44484# 0.007416f
C30977 a_2437_43646# a_2982_43646# 0.0016f
C30978 a_19787_47423# SINGLE_ENDED 2.87e-21
C30979 a_10193_42453# a_4361_42308# 0.274131f
C30980 a_15861_45028# a_10341_43396# 2.08e-20
C30981 a_n467_45028# a_n447_43370# 6.82e-20
C30982 a_n699_43396# a_n1761_44111# 0.018554f
C30983 a_n1059_45260# a_458_43396# 3e-19
C30984 a_n2017_45002# a_1209_43370# 4.18e-21
C30985 a_n2661_44458# a_2479_44172# 1.07e-19
C30986 a_n357_42282# a_12089_42308# 0.027195f
C30987 a_1307_43914# a_3052_44056# 0.001611f
C30988 a_11599_46634# a_18184_42460# 0.018223f
C30989 a_18189_46348# a_13259_45724# 0.016675f
C30990 a_5807_45002# a_14180_45002# 0.005192f
C30991 a_n743_46660# a_5691_45260# 3.07e-20
C30992 a_584_46384# a_949_44458# 0.011926f
C30993 a_n1151_42308# a_n1699_44726# 2.55e-19
C30994 a_765_45546# a_11823_42460# 2.37e-20
C30995 a_3090_45724# a_16333_45814# 0.007872f
C30996 a_15368_46634# a_15903_45785# 6.84e-19
C30997 a_15559_46634# a_15599_45572# 6.99e-21
C30998 a_16327_47482# a_17719_45144# 2.77e-19
C30999 a_13661_43548# a_13777_45326# 0.001317f
C31000 a_n971_45724# a_5883_43914# 0.027317f
C31001 a_3699_46348# a_3503_45724# 1.91e-19
C31002 a_4419_46090# a_3218_45724# 4.98e-22
C31003 a_n1925_46634# a_6171_45002# 0.005306f
C31004 a_14976_45028# a_15765_45572# 1.08e-20
C31005 a_5167_46660# a_3357_43084# 2.88e-19
C31006 a_12861_44030# a_21101_45002# 1.67e-20
C31007 a_10227_46804# a_16405_45348# 5.83e-20
C31008 a_6540_46812# a_2437_43646# 5.76e-21
C31009 a_1823_45246# a_n443_42852# 0.125287f
C31010 a_n2293_46098# a_4099_45572# 0.00692f
C31011 a_768_44030# a_626_44172# 0.186913f
C31012 a_15682_46116# a_16375_45002# 6.09e-19
C31013 a_5204_45822# a_n755_45592# 2.71e-20
C31014 a_17364_32525# C3_N_btm 1.38e-20
C31015 a_14209_32519# C5_N_btm 0.042017f
C31016 a_10545_42558# a_10533_42308# 0.011812f
C31017 a_n4318_38216# a_n4064_40160# 0.052465f
C31018 a_4361_42308# VDD 0.42717f
C31019 a_13887_32519# C7_N_btm 4.26e-20
C31020 a_13467_32519# RST_Z 0.048761f
C31021 a_564_42282# a_7174_31319# 9.76e-21
C31022 a_11827_44484# a_15743_43084# 3.38e-21
C31023 a_9482_43914# a_10991_42826# 8.72e-21
C31024 a_n967_45348# a_n914_42852# 1.98e-19
C31025 a_10334_44484# a_8685_43396# 1.89e-20
C31026 a_20841_46902# VDD 0.20446f
C31027 a_20273_46660# RST_Z 2.21e-21
C31028 a_20107_46660# SINGLE_ENDED 2.88e-21
C31029 a_7499_43078# a_5934_30871# 0.00463f
C31030 a_n913_45002# a_1793_42852# 0.00284f
C31031 a_765_45546# DATA[3] 0.004997f
C31032 a_11691_44458# a_17324_43396# 1.34e-21
C31033 a_n2293_42834# a_n1853_43023# 0.053782f
C31034 a_1307_43914# a_8037_42858# 2.06e-21
C31035 a_n2661_42834# a_n97_42460# 9.39e-19
C31036 a_20692_30879# a_22775_42308# 5.45e-21
C31037 a_n357_42282# a_18907_42674# 3.94e-20
C31038 a_2711_45572# a_8568_45546# 0.011004f
C31039 a_3483_46348# a_14537_43396# 0.087339f
C31040 a_9290_44172# a_3232_43370# 0.087744f
C31041 a_10355_46116# a_6171_45002# 3.21e-22
C31042 a_19321_45002# a_19615_44636# 0.035767f
C31043 a_13259_45724# a_17478_45572# 0.048668f
C31044 a_1799_45572# a_n2661_43922# 3.03e-20
C31045 a_1176_45822# a_626_44172# 1.95e-19
C31046 a_n2293_46098# a_5365_45348# 4.09e-19
C31047 a_n2956_39304# a_n2661_45010# 1.05e-20
C31048 a_8049_45260# a_18596_45572# 0.001924f
C31049 a_13747_46662# a_20362_44736# 5.6e-20
C31050 a_8199_44636# a_7705_45326# 8.08e-19
C31051 a_8953_45546# a_7229_43940# 7.78e-21
C31052 a_5937_45572# a_6709_45028# 0.629301f
C31053 a_8016_46348# a_8953_45002# 0.016464f
C31054 a_16375_45002# a_16680_45572# 5.99e-20
C31055 a_15682_46116# a_413_45260# 3.05e-20
C31056 a_8349_46414# a_8191_45002# 5.23e-21
C31057 a_6755_46942# a_15004_44636# 5.2e-19
C31058 a_6194_45824# a_6428_45938# 0.006453f
C31059 a_n4209_38502# a_n4334_38304# 3.3e-19
C31060 a_n4334_38528# a_n4209_38216# 3.3e-19
C31061 a_n3565_38502# a_n3607_38528# 0.001003f
C31062 a_n4064_38528# a_n2216_38778# 0.005567f
C31063 a_5934_30871# C8_N_btm 1.41e-19
C31064 a_6123_31319# C10_N_btm 1.34e-19
C31065 a_18907_42674# CAL_N 7.78e-19
C31066 a_5742_30871# C6_P_btm 0.170624f
C31067 a_6761_42308# VDD 0.259312f
C31068 a_1343_38525# VDAC_Pi 0.035744f
C31069 a_11599_46634# a_15811_47375# 0.107881f
C31070 a_14955_47212# a_15673_47210# 3.17e-19
C31071 a_4915_47217# a_12465_44636# 0.07724f
C31072 a_n1741_47186# a_9804_47204# 0.010096f
C31073 a_n971_45724# a_n881_46662# 0.236696f
C31074 a_n746_45260# a_n1613_43370# 0.146842f
C31075 a_2553_47502# a_2747_46873# 0.14563f
C31076 a_5815_47464# a_4883_46098# 4.29e-21
C31077 a_13717_47436# a_16763_47508# 2.89e-19
C31078 a_12861_44030# a_16023_47582# 2.79e-20
C31079 a_11459_47204# a_10227_46804# 6.22e-20
C31080 a_11341_43940# a_15095_43370# 4.91e-20
C31081 a_n809_44244# a_n901_43156# 0.001977f
C31082 a_n1549_44318# a_n1076_43230# 2.38e-20
C31083 a_n2293_43922# a_n2293_42282# 0.19201f
C31084 a_18114_32519# COMP_P 1.46e-20
C31085 a_509_45572# VDD 1.36e-19
C31086 a_5891_43370# a_7573_43172# 5.51e-21
C31087 a_14539_43914# a_14635_42282# 1.26e-19
C31088 a_n2956_37592# a_n2860_39866# 3.22e-20
C31089 a_n1699_43638# a_n1809_43762# 0.097745f
C31090 a_n1917_43396# a_n2012_43396# 0.049827f
C31091 a_n2267_43396# a_n1190_43762# 1.46e-19
C31092 a_n2129_43609# a_n1821_43396# 0.004509f
C31093 a_15682_43940# a_15781_43660# 0.005099f
C31094 a_20623_43914# a_10341_43396# 7.45e-20
C31095 a_3905_42865# a_5649_42852# 3.85e-20
C31096 a_11967_42832# a_10341_42308# 0.001434f
C31097 en_comp a_n2302_39866# 4.43e-20
C31098 a_n4318_40392# a_n3674_38216# 0.023361f
C31099 a_10586_45546# a_10057_43914# 1.37e-19
C31100 a_15227_44166# a_15682_43940# 0.072383f
C31101 a_n2312_38680# a_n1557_42282# 1.6e-20
C31102 a_10809_44734# a_9313_44734# 0.001335f
C31103 a_2711_45572# a_n2661_43370# 0.112998f
C31104 a_20273_45572# a_20528_45572# 0.064178f
C31105 a_20107_45572# a_20731_45938# 9.73e-19
C31106 a_20841_45814# a_21188_45572# 0.051162f
C31107 a_14495_45572# a_14537_43396# 2.49e-19
C31108 a_10907_45822# a_10951_45334# 0.002454f
C31109 a_n1151_42308# a_n2157_42858# 5.83e-19
C31110 a_3090_45724# a_15493_43396# 0.134629f
C31111 a_768_44030# a_2813_43396# 4.65e-19
C31112 a_16327_47482# a_16664_43396# 2.45e-19
C31113 a_n2293_46634# a_1891_43646# 8.05e-20
C31114 a_5807_45002# a_7927_46660# 0.004378f
C31115 a_n1741_47186# a_n901_46420# 1.81e-20
C31116 a_768_44030# a_6755_46942# 0.017611f
C31117 a_2063_45854# a_11415_45002# 5.51e-19
C31118 C6_P_btm C0_dummy_P_btm 0.120464f
C31119 C9_P_btm C1_N_btm 9.52e-19
C31120 C8_P_btm C0_N_btm 7e-19
C31121 C7_P_btm C0_dummy_N_btm 3.73e-19
C31122 a_11599_46634# a_13059_46348# 0.371555f
C31123 C3_P_btm C2_P_btm 5.64696f
C31124 C5_P_btm C0_P_btm 0.138736f
C31125 C4_P_btm C1_P_btm 0.128692f
C31126 a_n743_46660# a_4646_46812# 0.031686f
C31127 a_n2438_43548# a_3877_44458# 2.1e-20
C31128 a_n2661_46634# a_6540_46812# 0.007418f
C31129 EN_VIN_BSTR_N C7_N_btm 0.115875f
C31130 a_9313_45822# a_765_45546# 0.034184f
C31131 a_12861_44030# a_16751_46987# 7.13e-19
C31132 a_13507_46334# a_19692_46634# 0.823157f
C31133 a_4883_46098# a_19333_46634# 6.67e-20
C31134 a_2107_46812# a_2864_46660# 0.002314f
C31135 a_645_46660# a_n2661_46098# 2.43e-19
C31136 a_n1532_35090# VDD 2.19114f
C31137 a_n971_45724# a_n2157_46122# 0.001149f
C31138 a_n746_45260# a_n2293_46098# 0.027821f
C31139 a_8128_46384# a_8035_47026# 0.006018f
C31140 a_n1925_46634# a_4955_46873# 0.033508f
C31141 a_10227_46804# a_12925_46660# 0.001202f
C31142 a_11453_44696# a_15368_46634# 6.42e-20
C31143 a_n881_46662# a_8023_46660# 0.001443f
C31144 a_n2661_42282# a_1755_42282# 0.145244f
C31145 a_3422_30871# a_15890_42674# 2.49e-20
C31146 a_16137_43396# a_4361_42308# 0.019831f
C31147 a_3626_43646# a_13635_43156# 1.89e-19
C31148 a_2982_43646# a_14543_43071# 2.24e-21
C31149 a_8147_43396# a_8387_43230# 1.33e-19
C31150 a_16759_43396# a_743_42282# 1.02e-20
C31151 a_16664_43396# a_16855_43396# 4.61e-19
C31152 a_n97_42460# a_n2293_42282# 5.22e-19
C31153 a_17324_43396# a_4190_30871# 2.14e-20
C31154 a_11967_42832# a_18057_42282# 0.002498f
C31155 a_2680_45002# a_n2661_44458# 7.59e-20
C31156 a_n467_45028# a_n452_44636# 0.092885f
C31157 a_8696_44636# a_13213_44734# 0.004648f
C31158 a_15595_45028# a_16922_45042# 1.97e-20
C31159 a_16019_45002# a_16501_45348# 2.93e-19
C31160 a_8199_44636# a_2982_43646# 3.15e-19
C31161 a_17715_44484# a_n97_42460# 8.03e-20
C31162 a_4640_45348# a_n2661_43370# 4.5e-19
C31163 a_4185_45028# a_6197_43396# 7.89e-21
C31164 a_19692_46634# a_21855_43396# 0.016876f
C31165 a_17339_46660# a_18525_43370# 0.060382f
C31166 a_n2312_39304# a_n3674_38680# 0.023326f
C31167 a_n2312_40392# a_n2472_42282# 4.5e-20
C31168 a_n1059_45260# a_6298_44484# 2.2e-22
C31169 a_2711_45572# a_2998_44172# 1.79e-21
C31170 a_5257_43370# a_5164_46348# 0.02844f
C31171 a_5732_46660# a_5937_45572# 1.49e-19
C31172 a_4915_47217# a_2711_45572# 0.265557f
C31173 a_n443_46116# a_3175_45822# 0.002277f
C31174 a_8667_46634# a_3483_46348# 7.36e-19
C31175 a_15227_44166# a_22000_46634# 0.154332f
C31176 a_16292_46812# a_16434_46660# 0.007833f
C31177 a_13693_46688# a_13059_46348# 1.71e-19
C31178 a_768_44030# a_8049_45260# 0.027975f
C31179 a_13885_46660# a_14447_46660# 0.005162f
C31180 a_14035_46660# a_14226_46660# 2.88e-19
C31181 a_4883_46098# a_20062_46116# 9.7e-20
C31182 a_n1925_46634# a_n967_46494# 6.65e-20
C31183 a_5807_45002# a_6419_46482# 0.005524f
C31184 a_n1151_42308# a_6667_45809# 9.3e-20
C31185 a_n971_45724# a_8162_45546# 0.015463f
C31186 a_19692_46634# a_20623_46660# 0.03624f
C31187 a_n2438_43548# a_n1736_46482# 2.63e-20
C31188 a_16327_47482# a_n357_42282# 0.49929f
C31189 a_13507_46334# a_20692_30879# 6.68e-19
C31190 a_17730_32519# C5_N_btm 8.54e-20
C31191 a_743_42282# a_1067_42314# 0.010185f
C31192 a_10796_42968# a_11554_42852# 0.056391f
C31193 a_10991_42826# a_11301_43218# 0.013793f
C31194 a_10922_42852# a_11229_43218# 3.69e-19
C31195 a_22315_44484# RST_Z 5.65e-20
C31196 a_8685_43396# a_15051_42282# 7.21e-19
C31197 a_2982_43646# a_19511_42282# 0.014171f
C31198 a_3626_43646# a_18310_42308# 0.00142f
C31199 a_4361_42308# a_n784_42308# 2.34e-20
C31200 a_13887_32519# COMP_P 6.33e-21
C31201 a_n2472_42826# a_n3674_38680# 0.004228f
C31202 a_9145_43396# a_13575_42558# 4.11e-19
C31203 a_20820_30879# a_22400_42852# 1.3e-19
C31204 a_5883_43914# a_9313_44734# 0.124999f
C31205 a_16327_47482# CAL_N 0.001106f
C31206 a_18494_42460# a_11967_42832# 0.025796f
C31207 a_6171_45002# a_10949_43914# 9.46e-21
C31208 a_3232_43370# a_10807_43548# 0.001324f
C31209 a_n443_42852# a_17324_43396# 1.63e-21
C31210 a_20205_31679# a_13678_32519# 0.051502f
C31211 a_7499_43078# a_7221_43396# 4.61e-20
C31212 a_8975_43940# a_5891_43370# 0.021307f
C31213 a_n2012_44484# a_n1821_44484# 4.61e-19
C31214 a_n452_44636# a_n2661_43922# 0.009547f
C31215 a_742_44458# a_n2661_42834# 0.034578f
C31216 a_n2293_42834# a_n1899_43946# 0.001698f
C31217 a_20202_43084# a_20256_42852# 0.001339f
C31218 a_n1920_47178# VDD 0.229556f
C31219 a_n2833_47464# CLK_DATA 0.331592f
C31220 a_11827_44484# a_16789_44484# 2.76e-19
C31221 a_19778_44110# a_20159_44458# 2.12e-20
C31222 a_1423_45028# a_7281_43914# 0.001025f
C31223 a_18479_45785# a_19478_44056# 3.95e-19
C31224 a_2437_43646# a_2253_43940# 0.003306f
C31225 a_3090_45724# a_6472_45840# 1.07e-21
C31226 a_13747_46662# a_21363_45546# 0.001465f
C31227 a_16119_47582# a_2437_43646# 0.001405f
C31228 a_4883_46098# a_5147_45002# 5.63e-20
C31229 a_12594_46348# a_10809_44734# 0.082565f
C31230 a_4791_45118# a_5365_45348# 0.001047f
C31231 a_20202_43084# a_13259_45724# 2.57e-19
C31232 a_n881_46662# a_n2293_45010# 9.84e-21
C31233 a_4185_45028# a_5066_45546# 2.04e-20
C31234 a_12549_44172# a_3357_43084# 0.001325f
C31235 a_17583_46090# a_18819_46122# 1.6e-21
C31236 a_17715_44484# a_17957_46116# 0.005313f
C31237 a_13759_46122# a_6945_45028# 7.74e-20
C31238 a_6755_46942# a_11652_45724# 1.83e-20
C31239 a_11599_46634# a_13556_45296# 5.22e-21
C31240 a_7274_43762# VDD 4.6e-19
C31241 a_2725_42558# a_2903_42308# 5.98e-20
C31242 a_564_42282# a_5932_42308# 8.68e-21
C31243 a_n784_42308# a_6761_42308# 2.26e-20
C31244 a_13291_42460# a_13657_42308# 0.001043f
C31245 a_15004_44636# a_15037_43940# 1.72e-20
C31246 a_n452_44636# a_n447_43370# 0.001136f
C31247 a_10428_46928# DATA[5] 0.002585f
C31248 a_n2661_45010# a_685_42968# 5.86e-22
C31249 a_3357_43084# a_5111_42852# 5.76e-19
C31250 a_n699_43396# a_n2267_43396# 1.05e-19
C31251 a_9863_46634# CLK 0.001256f
C31252 a_n2956_37592# a_n4318_38680# 0.023187f
C31253 en_comp a_n3674_39304# 3.39e-19
C31254 a_n443_42852# a_1184_42692# 0.003744f
C31255 a_n357_42282# a_5267_42460# 1.81e-20
C31256 a_n755_45592# a_3823_42558# 0.001851f
C31257 a_11823_42460# a_13291_42460# 0.257506f
C31258 a_5147_45002# a_5649_42852# 2.35e-21
C31259 a_n809_44244# a_n984_44318# 0.234322f
C31260 a_12861_44030# a_20766_44850# 5.26e-19
C31261 a_10227_46804# a_16241_44484# 4.52e-20
C31262 a_310_45028# a_n23_45546# 0.022295f
C31263 a_n1099_45572# a_n310_45899# 4.53e-19
C31264 a_8049_45260# a_11652_45724# 0.002134f
C31265 a_n2293_45546# a_n443_42852# 0.084694f
C31266 a_10809_44734# a_15037_45618# 4.19e-21
C31267 a_14513_46634# a_14537_43396# 1.12e-21
C31268 a_n1991_46122# a_n2661_45010# 2.05e-19
C31269 a_1823_45246# a_2437_43646# 0.324477f
C31270 a_18597_46090# a_17517_44484# 0.021693f
C31271 a_n863_45724# a_n906_45572# 0.002589f
C31272 a_13059_46348# a_13348_45260# 0.010157f
C31273 a_584_46384# a_175_44278# 0.001131f
C31274 a_n1151_42308# a_n1761_44111# 0.642214f
C31275 a_n2157_46122# a_n2293_45010# 1.83e-20
C31276 a_n755_45592# a_3503_45724# 0.163919f
C31277 a_n357_42282# a_n356_45724# 2.1e-19
C31278 a_n743_46660# a_10057_43914# 2.57e-20
C31279 a_18189_46348# a_17478_45572# 0.002791f
C31280 a_10586_45546# a_10180_45724# 7.02e-19
C31281 a_2324_44458# a_12649_45572# 4.41e-19
C31282 a_16327_47482# a_18588_44850# 0.012252f
C31283 a_13622_42852# VDD 4.6e-19
C31284 COMP_P EN_VIN_BSTR_N 0.004364f
C31285 a_n4209_39590# a_n4064_39616# 0.269818f
C31286 a_2063_45854# a_2553_47502# 0.040297f
C31287 a_n971_45724# a_n443_46116# 0.129009f
C31288 a_1239_47204# a_n1151_42308# 0.007713f
C31289 a_n1741_47186# a_6545_47178# 0.053219f
C31290 a_1209_47178# a_3381_47502# 7.34e-20
C31291 a_n3565_39590# a_n3420_39616# 0.281955f
C31292 a_n2661_42834# a_n901_43156# 0.001144f
C31293 a_n2293_43922# a_n1423_42826# 1.71e-20
C31294 a_742_44458# a_n2293_42282# 0.006579f
C31295 a_5111_44636# a_6123_31319# 1.17e-19
C31296 a_8379_46155# VDD 2.18e-20
C31297 a_18579_44172# a_18525_43370# 0.012789f
C31298 a_19279_43940# a_19268_43646# 5.83e-21
C31299 a_n356_44636# a_10083_42826# 4.56e-20
C31300 en_comp a_5742_30871# 0.092238f
C31301 a_n913_45002# a_13070_42354# 4.84e-20
C31302 a_n1059_45260# a_13575_42558# 8.82e-21
C31303 a_n2017_45002# a_14456_42282# 0.003727f
C31304 a_375_42282# a_1184_42692# 1.26e-19
C31305 a_14539_43914# a_14543_43071# 8.67e-19
C31306 a_12549_44172# a_18533_44260# 3.67e-19
C31307 a_n863_45724# a_1307_43914# 0.050349f
C31308 a_n2661_45546# a_1145_45348# 1.22e-19
C31309 a_11415_45002# a_n2661_42834# 3.35e-20
C31310 a_n357_42282# a_14537_43396# 7.25e-21
C31311 a_2324_44458# a_4223_44672# 0.56408f
C31312 a_n2293_45546# a_375_42282# 0.104283f
C31313 a_9290_44172# a_8975_43940# 0.114958f
C31314 a_2711_45572# a_4574_45260# 8.29e-19
C31315 a_2107_46812# a_9895_44260# 6.01e-19
C31316 a_22521_40599# a_22521_39511# 0.365591f
C31317 CAL_N a_22545_38993# 0.01247f
C31318 a_6886_37412# CAL_P 0.002915f
C31319 a_n881_46662# a_601_46902# 4.24e-19
C31320 a_6575_47204# a_6969_46634# 2.23e-19
C31321 a_n1435_47204# a_10150_46912# 1.49e-20
C31322 a_9067_47204# a_6755_46942# 1.22e-19
C31323 a_11459_47204# a_10467_46802# 4.67e-19
C31324 a_n1613_43370# a_383_46660# 0.182504f
C31325 a_5807_45002# a_19594_46812# 1.59e-19
C31326 a_13661_43548# a_19321_45002# 7.35e-19
C31327 a_n4064_37440# a_n923_35174# 0.002259f
C31328 a_12549_44172# a_n2293_46634# 0.005061f
C31329 a_13747_46662# a_19452_47524# 0.003322f
C31330 a_n2860_37984# VDD 0.004232f
C31331 a_6151_47436# a_8035_47026# 0.038687f
C31332 a_n1151_42308# a_11186_47026# 4.42e-20
C31333 a_2063_45854# a_12251_46660# 2.19e-19
C31334 a_2747_46873# a_1799_45572# 5.65e-19
C31335 a_9804_47204# a_n743_46660# 0.295465f
C31336 a_20447_31679# VDD 0.665681f
C31337 a_14021_43940# a_17701_42308# 9.5e-20
C31338 a_2982_43646# a_21259_43561# 0.034927f
C31339 a_15095_43370# a_10341_43396# 0.013375f
C31340 a_13667_43396# a_12281_43396# 1.88e-20
C31341 a_n2661_42834# a_10533_42308# 4.35e-22
C31342 a_n2840_43914# a_n4318_38216# 8.56e-19
C31343 a_2437_43646# DATA[2] 0.046972f
C31344 a_3080_42308# a_4361_42308# 8.53e-19
C31345 a_22959_45572# RST_Z 0.001363f
C31346 a_8685_43396# a_13749_43396# 6.06e-19
C31347 a_n2267_43396# a_n4318_38680# 3e-19
C31348 a_n1699_43638# a_n3674_39304# 2.54e-19
C31349 a_n97_42460# a_n1423_42826# 6.33e-21
C31350 a_n1352_43396# a_n901_43156# 1.07e-20
C31351 a_n1809_43762# a_n2157_42858# 2.44e-20
C31352 a_n1177_43370# a_n1076_43230# 9.51e-21
C31353 a_9801_43940# a_9127_43156# 5.84e-20
C31354 en_comp a_n2293_42834# 0.103485f
C31355 a_n2472_45002# a_n2661_43370# 0.017331f
C31356 a_20273_45572# a_18494_42460# 0.002243f
C31357 a_n2497_47436# a_564_42282# 3.52e-21
C31358 a_2324_44458# a_15493_43940# 0.061147f
C31359 a_13348_45260# a_13556_45296# 0.189446f
C31360 a_13159_45002# a_13777_45326# 8.25e-20
C31361 a_10193_42453# a_5891_43370# 0.001973f
C31362 a_n357_42282# a_20835_44721# 8.73e-21
C31363 a_4574_45260# a_4640_45348# 0.006978f
C31364 a_3537_45260# a_5105_45348# 3.16e-19
C31365 a_n1925_42282# a_n2661_42282# 2.27741f
C31366 a_413_45260# a_2809_45028# 0.005798f
C31367 a_18799_45938# a_11691_44458# 7.04e-20
C31368 a_6431_45366# a_1423_45028# 1.36e-20
C31369 a_8049_45260# a_7845_44172# 7.46e-20
C31370 a_20107_45572# a_20567_45036# 9.82e-19
C31371 a_13017_45260# a_14180_45002# 0.079928f
C31372 a_4558_45348# a_4185_45348# 1.34e-19
C31373 a_3090_45724# a_10695_43548# 0.005861f
C31374 a_10903_43370# a_12710_44260# 0.001775f
C31375 a_12549_44172# a_5342_30871# 4.48e-20
C31376 a_n2438_43548# a_1847_42826# 3.92e-21
C31377 a_6755_46942# a_16759_43396# 5.96e-19
C31378 a_4646_46812# a_4361_42308# 9.53e-20
C31379 a_22731_47423# a_6945_45028# 8.58e-20
C31380 a_171_46873# a_n1991_46122# 7.76e-21
C31381 a_5807_45002# a_5164_46348# 5.51e-19
C31382 a_768_44030# a_8953_45546# 0.025581f
C31383 a_10249_46116# a_12978_47026# 4.67e-21
C31384 a_6755_46942# a_10933_46660# 5.53e-19
C31385 a_11735_46660# a_13607_46688# 1.3e-20
C31386 a_12469_46902# a_12251_46660# 0.209641f
C31387 a_11901_46660# a_12991_46634# 0.042415f
C31388 a_11813_46116# a_12816_46660# 5.47e-21
C31389 a_22223_47212# a_22223_46124# 8.8e-19
C31390 a_12465_44636# a_10809_44734# 0.099854f
C31391 a_n2438_43548# a_n1641_46494# 4.44e-20
C31392 a_n743_46660# a_n901_46420# 0.004763f
C31393 a_9067_47204# a_8049_45260# 1.65e-19
C31394 a_n881_46662# a_12594_46348# 1.17e-19
C31395 a_6540_46812# a_765_45546# 0.00357f
C31396 a_9804_47204# a_11189_46129# 2.45e-20
C31397 a_n2661_46634# a_1823_45246# 3e-19
C31398 a_n1021_46688# a_n1076_46494# 3.41e-20
C31399 a_n1925_46634# a_376_46348# 0.002206f
C31400 a_n2497_47436# a_n2810_45572# 1.01e-20
C31401 a_n2833_47464# a_n2661_45546# 3.61e-20
C31402 a_5649_42852# a_5457_43172# 1.97e-19
C31403 a_n901_43156# a_n2293_42282# 7.23e-20
C31404 a_2982_43646# a_4921_42308# 0.001781f
C31405 a_3539_42460# a_3581_42558# 0.002471f
C31406 a_3626_43646# a_3905_42558# 0.004928f
C31407 a_4905_42826# a_6773_42558# 8.37e-21
C31408 a_5891_43370# VDD 2.12137f
C31409 a_n97_42460# a_9885_42558# 0.011255f
C31410 a_10835_43094# a_10922_42852# 0.053385f
C31411 a_10518_42984# a_10341_42308# 0.00245f
C31412 a_10796_42968# a_10991_42826# 0.206455f
C31413 a_4185_45028# a_10922_42852# 1.72e-20
C31414 a_12549_44172# a_20107_42308# 3.8e-21
C31415 a_16855_45546# a_15493_43940# 1.91e-22
C31416 a_8696_44636# a_11341_43940# 1.44e-19
C31417 a_10193_42453# a_18533_43940# 0.007041f
C31418 a_n2661_44458# a_5518_44484# 0.01193f
C31419 a_n2661_45546# a_3457_43396# 0.030099f
C31420 a_n2312_40392# a_n2216_39866# 5.49e-20
C31421 a_n1059_45260# a_2479_44172# 0.004979f
C31422 a_n2017_45002# a_895_43940# 2.49e-20
C31423 SMPL_ON_P a_n2946_37690# 2.4e-19
C31424 a_11827_44484# a_17970_44736# 0.012326f
C31425 a_11691_44458# a_16112_44458# 0.012386f
C31426 a_1307_43914# a_16241_44484# 0.001942f
C31427 a_n467_45028# a_n809_44244# 0.010788f
C31428 a_18494_42460# a_18989_43940# 1.47e-20
C31429 a_13661_43548# a_17531_42308# 1.49e-21
C31430 a_4646_46812# a_6761_42308# 2.07e-21
C31431 a_8199_44636# a_7871_42858# 1.17e-20
C31432 a_13507_46334# a_18175_45572# 3.67e-20
C31433 a_11415_45002# a_17715_44484# 0.032854f
C31434 a_3483_46348# a_5204_45822# 2.01e-19
C31435 a_3699_46348# a_5164_46348# 1.23e-21
C31436 a_20528_46660# a_10809_44734# 0.004492f
C31437 a_11031_47542# a_2437_43646# 0.003672f
C31438 a_19386_47436# a_19431_45546# 8.77e-20
C31439 a_18597_46090# a_19256_45572# 0.001301f
C31440 a_n2661_46634# a_12427_45724# 4.09e-20
C31441 a_n2109_47186# a_3232_43370# 3.24e-19
C31442 a_n971_45724# a_3537_45260# 0.266743f
C31443 a_4419_46090# a_4704_46090# 0.016592f
C31444 a_n881_46662# a_15037_45618# 0.044816f
C31445 a_6575_47204# a_3357_43084# 8.41e-19
C31446 a_n237_47217# a_3065_45002# 2.45e-20
C31447 a_12741_44636# a_2324_44458# 0.019655f
C31448 a_n743_46660# a_10180_45724# 2.31e-19
C31449 a_16327_47482# a_18953_45572# 0.002336f
C31450 a_14401_32519# C7_N_btm 9.48e-19
C31451 a_17538_32519# C5_N_btm 4.27e-20
C31452 a_3080_42308# a_n1532_35090# 6.43e-20
C31453 a_22400_42852# a_20753_42852# 6.01e-21
C31454 a_18533_43940# VDD 0.182147f
C31455 a_17701_42308# a_15764_42576# 1.32e-20
C31456 a_n2661_43922# a_n809_44244# 0.010689f
C31457 a_n2293_43922# a_n1549_44318# 1.15e-19
C31458 a_n2661_42834# a_n984_44318# 0.012148f
C31459 a_8975_43940# a_10807_43548# 2.16e-19
C31460 a_n2661_46634# DATA[2] 1.39e-19
C31461 a_11823_42460# a_13460_43230# 0.00394f
C31462 a_n2293_42834# a_n1699_43638# 0.005603f
C31463 a_1307_43914# a_3540_43646# 0.005727f
C31464 a_19615_44636# a_20362_44736# 2.51e-19
C31465 a_11967_42832# a_20640_44752# 0.588649f
C31466 a_19006_44850# a_20679_44626# 6.41e-22
C31467 a_8953_45002# a_8791_43396# 4.51e-19
C31468 a_10193_42453# a_17595_43084# 2.47e-19
C31469 a_n2956_38680# a_6123_31319# 3.8e-21
C31470 a_10903_43370# a_14113_42308# 1.69e-20
C31471 a_n1021_46688# VDD 0.226043f
C31472 a_12607_44458# a_10949_43914# 7.79e-20
C31473 a_4185_45028# a_17531_42308# 6.87e-20
C31474 a_21588_30879# EN_OFFSET_CAL 0.047538f
C31475 a_3537_45260# a_8229_43396# 1.13e-20
C31476 a_5111_44636# a_6809_43396# 0.002123f
C31477 a_18479_45785# a_4361_42308# 5.55e-20
C31478 a_13249_42308# a_12089_42308# 0.002934f
C31479 a_10809_44734# a_2711_45572# 0.037787f
C31480 a_11415_45002# a_15861_45028# 0.041647f
C31481 a_2609_46660# a_2809_45028# 5.53e-21
C31482 a_3877_44458# a_2903_45348# 2.68e-20
C31483 a_10903_43370# a_7499_43078# 0.888628f
C31484 a_19321_45002# a_18587_45118# 2.02e-19
C31485 a_6755_46942# a_7276_45260# 4.58e-22
C31486 a_13747_46662# a_19778_44110# 0.670692f
C31487 a_13661_43548# a_18184_42460# 0.031622f
C31488 a_11735_46660# a_413_45260# 5.06e-20
C31489 a_12741_44636# a_16855_45546# 7.31e-20
C31490 a_2063_45854# a_n2661_43922# 0.033229f
C31491 a_3483_46348# a_8697_45822# 0.033264f
C31492 a_11189_46129# a_10180_45724# 4.36e-20
C31493 a_9290_44172# a_10193_42453# 1.23123f
C31494 a_10355_46116# a_8746_45002# 0.002156f
C31495 a_16327_47482# a_18443_44721# 0.1665f
C31496 a_15890_42674# a_7174_31319# 2.06e-20
C31497 a_4958_30871# a_17303_42282# 0.168656f
C31498 a_n1630_35242# a_n2302_37984# 5.02e-20
C31499 a_17595_43084# VDD 0.168112f
C31500 a_n2956_38216# a_n2946_37984# 0.150404f
C31501 a_n2810_45028# a_n3674_38680# 0.022953f
C31502 a_9290_44172# VDD 2.74561f
C31503 a_18248_44752# a_16823_43084# 1.7e-19
C31504 a_10057_43914# a_4361_42308# 3.62e-20
C31505 a_20365_43914# a_11341_43940# 0.010232f
C31506 a_8016_46348# DATA[4] 7.36e-22
C31507 a_10193_42453# a_21887_42336# 3.37e-21
C31508 a_n2017_45002# a_n3674_38216# 0.004889f
C31509 a_13483_43940# a_13565_44260# 0.003935f
C31510 a_n1761_44111# a_n1809_43762# 4.8e-19
C31511 a_n809_44244# a_n447_43370# 0.003582f
C31512 a_n984_44318# a_n1352_43396# 5.83e-20
C31513 a_n2956_37592# a_n2840_42282# 8.96e-21
C31514 a_19862_44208# a_15493_43940# 0.534481f
C31515 a_2711_45572# a_16211_45572# 0.001012f
C31516 a_n2661_45546# a_3357_43084# 0.045914f
C31517 a_2324_44458# a_n2293_42834# 0.168086f
C31518 a_584_46384# a_n97_42460# 0.526796f
C31519 a_n2497_47436# a_n1557_42282# 7.44e-20
C31520 a_6755_46942# a_17517_44484# 8.4e-20
C31521 a_4185_45028# a_18184_42460# 0.006813f
C31522 a_n2293_45546# a_2437_43646# 0.031092f
C31523 a_768_44030# a_9028_43914# 0.113848f
C31524 a_n2293_46634# a_7542_44172# 5.45e-20
C31525 a_8746_45002# a_10544_45572# 4.52e-20
C31526 a_10490_45724# a_10306_45572# 8.03e-20
C31527 a_8049_45260# a_7276_45260# 5.67e-19
C31528 a_8034_45724# a_8191_45002# 1.83e-20
C31529 a_18597_46090# a_12549_44172# 0.042681f
C31530 a_12465_44636# a_n881_46662# 0.813228f
C31531 a_n3420_39072# a_n923_35174# 0.004736f
C31532 a_2063_45854# a_1799_45572# 5.95e-19
C31533 a_584_46384# a_n2661_46098# 0.17431f
C31534 a_n1151_42308# a_491_47026# 0.002342f
C31535 a_6545_47178# a_n743_46660# 0.003782f
C31536 a_16241_47178# a_16131_47204# 0.097745f
C31537 a_16327_47482# a_16942_47570# 0.001965f
C31538 a_21335_42336# RST_Z 1.97e-20
C31539 a_3815_47204# a_2107_46812# 4.62e-20
C31540 a_6851_47204# a_n1925_46634# 6.48e-20
C31541 a_15673_47210# a_5807_45002# 0.011029f
C31542 a_21887_42336# VDD 0.210392f
C31543 a_n4064_39616# C6_P_btm 1.1e-19
C31544 a_n3420_39616# C4_P_btm 3.39e-20
C31545 a_13717_47436# a_20916_46384# 1.15e-19
C31546 a_11031_47542# a_n2661_46634# 3.8e-20
C31547 a_n746_45260# a_1057_46660# 6.69e-20
C31548 a_n2109_47186# a_4651_46660# 0.025236f
C31549 a_n1741_47186# a_3877_44458# 1.26e-19
C31550 a_14021_43940# a_4361_42308# 0.003147f
C31551 a_18533_43940# a_16137_43396# 4.77e-20
C31552 a_5883_43914# a_8515_42308# 5.6e-22
C31553 a_10210_45822# CLK 5.07e-19
C31554 a_n356_44636# a_2351_42308# 1.17e-19
C31555 a_5343_44458# a_8685_42308# 5.14e-19
C31556 a_n97_42460# a_15095_43370# 0.002411f
C31557 a_5891_43370# a_n784_42308# 6.43e-20
C31558 a_3626_43646# a_8791_43396# 1.23e-21
C31559 a_5907_45546# a_5518_44484# 2.57e-19
C31560 a_3357_43084# a_5205_44484# 0.020505f
C31561 a_21588_30879# a_15743_43084# 3.87e-20
C31562 a_4646_46812# a_7274_43762# 2.49e-19
C31563 a_n2312_39304# a_n4318_38680# 0.0235f
C31564 a_n357_42282# a_n356_44636# 0.308599f
C31565 a_12741_44636# a_19862_44208# 8.5e-21
C31566 a_12549_44172# a_743_42282# 0.119701f
C31567 a_5257_43370# a_6197_43396# 0.001674f
C31568 a_n913_45002# a_2382_45260# 0.021705f
C31569 a_n2017_45002# a_3065_45002# 0.043491f
C31570 a_310_45028# a_n23_44458# 0.002647f
C31571 a_2711_45572# a_5883_43914# 2.93e-21
C31572 a_4651_46660# a_5841_46660# 2.56e-19
C31573 a_3877_44458# a_7832_46660# 2.27e-20
C31574 SMPL_ON_P a_n2956_38680# 0.039338f
C31575 a_n1741_47186# a_n1736_46482# 1.99e-19
C31576 a_4817_46660# a_6682_46987# 4.3e-20
C31577 a_9067_47204# a_8953_45546# 0.00218f
C31578 a_12549_44172# a_19123_46287# 1.7e-19
C31579 a_13747_46662# a_15227_46910# 5.38e-22
C31580 a_5807_45002# a_16388_46812# 0.235518f
C31581 a_13661_43548# a_13059_46348# 0.267127f
C31582 a_7411_46660# a_7577_46660# 0.634781f
C31583 a_14401_32519# COMP_P 8.68e-21
C31584 a_n2433_43396# a_n2472_42282# 2.98e-20
C31585 a_16547_43609# a_16414_43172# 0.143695f
C31586 a_16243_43396# a_16795_42852# 8.18e-20
C31587 a_743_42282# a_5111_42852# 8.1e-20
C31588 a_16137_43396# a_17595_43084# 0.001749f
C31589 a_18114_32519# C6_N_btm 2.2e-19
C31590 a_19721_31679# C5_N_btm 1.11e-20
C31591 a_n2472_42826# a_n4318_38680# 0.158196f
C31592 a_n2157_42858# a_n3674_39304# 2.93e-19
C31593 a_n1991_42858# a_n1076_43230# 0.123255f
C31594 a_n1853_43023# a_n13_43084# 0.109925f
C31595 a_2982_43646# a_13291_42460# 2.6e-19
C31596 a_n4318_39304# a_n4318_38216# 0.023477f
C31597 a_n356_44636# CAL_N 5.72e-19
C31598 a_n2312_38680# a_n3674_37592# 0.026177f
C31599 a_n443_42852# a_1443_43940# 3.91e-20
C31600 a_5205_44484# a_5826_44734# 0.003766f
C31601 a_526_44458# a_8147_43396# 2.13e-19
C31602 a_3537_45260# a_9313_44734# 6.69e-20
C31603 a_20273_45572# a_20640_44752# 7.28e-19
C31604 a_20107_45572# a_20679_44626# 0.001176f
C31605 a_19479_31679# a_17517_44484# 0.002614f
C31606 a_3232_43370# a_8375_44464# 0.022129f
C31607 a_5691_45260# a_5891_43370# 3.67e-21
C31608 a_21188_45572# a_11967_42832# 2.72e-22
C31609 a_10193_42453# a_10807_43548# 0.060211f
C31610 a_10490_45724# a_10729_43914# 2.89e-21
C31611 a_8746_45002# a_10949_43914# 4.6e-20
C31612 a_n467_45028# a_n2661_42834# 0.001028f
C31613 a_6171_45002# a_7640_43914# 8.9e-20
C31614 a_6431_45366# a_6109_44484# 2.93e-19
C31615 a_2809_45028# a_2779_44458# 0.001617f
C31616 a_16751_45260# a_14539_43914# 3.77e-20
C31617 a_15227_44166# a_18249_42858# 2.56e-20
C31618 a_n2293_46634# a_n2661_45546# 0.85166f
C31619 a_n2442_46660# a_n2472_45546# 5.69e-20
C31620 a_15009_46634# a_15015_46420# 0.012232f
C31621 a_11459_47204# a_11682_45822# 6.52e-21
C31622 a_4915_47217# a_14033_45822# 0.002034f
C31623 a_21350_47026# a_12741_44636# 2.49e-19
C31624 a_5257_43370# a_5066_45546# 0.053231f
C31625 a_768_44030# a_1609_45822# 3.5e-21
C31626 a_n2661_46634# a_n2293_45546# 5.66e-20
C31627 a_n2472_46634# a_n2956_38216# 7.81e-20
C31628 a_765_45546# a_1823_45246# 0.005338f
C31629 a_22365_46825# a_11415_45002# 0.007146f
C31630 a_4883_46098# a_7499_43078# 8.38e-19
C31631 a_10227_46804# a_11823_42460# 0.428745f
C31632 a_n881_46662# a_2711_45572# 0.170524f
C31633 a_15368_46634# a_13925_46122# 7.07e-20
C31634 a_19268_43646# a_19332_42282# 2.41e-19
C31635 a_10807_43548# VDD 0.68049f
C31636 a_5649_42852# a_14113_42308# 9.77e-20
C31637 a_5342_30871# a_n1630_35242# 0.035143f
C31638 a_4361_42308# a_15764_42576# 0.009129f
C31639 a_n443_42852# a_7227_42852# 0.008558f
C31640 a_20990_47178# VDD 0.210484f
C31641 a_19787_47423# START 0.220891f
C31642 a_9290_44172# a_n784_42308# 1.07e-19
C31643 a_20894_47436# RST_Z 5.48e-20
C31644 en_comp a_n2012_43396# 4.42e-20
C31645 a_n2661_42834# a_n2661_43922# 0.841361f
C31646 a_18989_43940# a_20640_44752# 1.37e-21
C31647 a_n1352_44484# a_n984_44318# 7.43e-19
C31648 a_n452_44636# a_n809_44244# 0.002409f
C31649 a_2437_43646# a_2896_43646# 5.48e-19
C31650 a_7499_43078# a_5649_42852# 2.19e-19
C31651 a_10193_42453# a_13467_32519# 0.005873f
C31652 a_1823_45246# a_4921_42308# 4.85e-19
C31653 a_626_44172# a_726_44056# 7.66e-19
C31654 a_8696_44636# a_10341_43396# 6.7e-21
C31655 a_22612_30879# VDAC_N 0.003601f
C31656 a_n2661_45010# a_1756_43548# 2.49e-21
C31657 a_n1059_45260# a_n229_43646# 3.39e-19
C31658 a_n357_42282# a_12379_42858# 0.031137f
C31659 a_16023_47582# CLK 0.002544f
C31660 a_1307_43914# a_2455_43940# 0.047238f
C31661 a_10227_46804# a_16321_45348# 9.56e-20
C31662 a_11599_46634# a_19778_44110# 1.94e-19
C31663 a_17715_44484# a_13259_45724# 0.391904f
C31664 a_1138_42852# a_n443_42852# 0.14758f
C31665 a_n2293_46634# a_5205_44484# 2.48e-19
C31666 a_1176_45822# a_1609_45822# 0.010535f
C31667 a_n2293_46098# a_3175_45822# 0.008709f
C31668 a_491_47026# a_327_44734# 5.88e-21
C31669 a_584_46384# a_742_44458# 0.031608f
C31670 a_n1151_42308# a_n2267_44484# 2.66e-19
C31671 a_15368_46634# a_15599_45572# 0.100853f
C31672 a_16327_47482# a_17613_45144# 7.07e-20
C31673 a_13747_46662# a_9482_43914# 1.7e-20
C31674 a_5807_45002# a_13777_45326# 1.7e-21
C31675 a_13661_43548# a_13556_45296# 0.559682f
C31676 a_n971_45724# a_8701_44490# 8.96e-19
C31677 a_3483_46348# a_3503_45724# 0.009385f
C31678 a_3090_45724# a_15765_45572# 0.046838f
C31679 a_14976_45028# a_15903_45785# 1.22e-19
C31680 a_5385_46902# a_3357_43084# 0.001502f
C31681 a_12861_44030# a_21005_45260# 1.13e-21
C31682 a_13507_46334# a_13490_45394# 1.03e-19
C31683 a_2107_46812# a_2382_45260# 5.81e-22
C31684 a_n237_47217# a_6298_44484# 8.52e-20
C31685 a_17364_32525# C2_N_btm 1.14e-20
C31686 a_9885_42558# a_10533_42308# 5.68e-21
C31687 a_9803_42558# a_5742_30871# 0.002197f
C31688 a_n4318_38216# a_n4334_40480# 9.74e-20
C31689 a_13887_32519# C6_N_btm 1.01e-19
C31690 a_13467_32519# VDD 0.353373f
C31691 a_1423_45028# a_3935_42891# 2.7e-22
C31692 a_11827_44484# a_18783_43370# 1.47e-20
C31693 a_20273_46660# VDD 0.247553f
C31694 a_20411_46873# RST_Z 1.31e-20
C31695 a_n913_45002# a_1709_42852# 0.0021f
C31696 a_n1059_45260# a_1793_42852# 4.52e-19
C31697 a_765_45546# DATA[2] 0.006631f
C31698 a_11691_44458# a_17499_43370# 3.7e-20
C31699 a_n2293_42834# a_n2157_42858# 0.058852f
C31700 a_n2293_43922# a_n1177_43370# 1.47e-22
C31701 a_n2661_42834# a_n447_43370# 0.006056f
C31702 a_3357_43084# a_3863_42891# 5.79e-19
C31703 a_20205_31679# a_22775_42308# 4.58e-21
C31704 a_n357_42282# a_18727_42674# 4.23e-20
C31705 a_7499_43078# a_7963_42308# 5.61e-19
C31706 a_2711_45572# a_8162_45546# 0.019489f
C31707 a_3483_46348# a_14180_45002# 2.73e-20
C31708 a_9823_46155# a_6171_45002# 9.16e-22
C31709 a_19321_45002# a_11967_42832# 0.266816f
C31710 a_13259_45724# a_15861_45028# 0.16873f
C31711 a_1138_42852# a_375_42282# 7.22e-21
C31712 a_n2293_46098# a_5105_45348# 2.55e-19
C31713 a_16388_46812# a_18315_45260# 5e-21
C31714 a_12549_44172# a_19789_44512# 5e-19
C31715 a_8049_45260# a_19256_45572# 0.007359f
C31716 a_13661_43548# a_20362_44736# 5.77e-20
C31717 a_13747_46662# a_20159_44458# 1.78e-20
C31718 a_5937_45572# a_7229_43940# 0.126047f
C31719 a_16375_45002# a_16855_45546# 2.09e-19
C31720 a_2324_44458# a_413_45260# 0.021366f
C31721 a_8016_46348# a_8191_45002# 3.05e-20
C31722 a_4646_46812# a_5891_43370# 0.089437f
C31723 a_3775_45552# a_3733_45822# 7.47e-21
C31724 a_5263_45724# a_5437_45600# 0.006584f
C31725 a_6194_45824# a_4880_45572# 4.69e-20
C31726 a_n4209_38502# a_n4209_38216# 0.041706f
C31727 a_n4064_38528# a_n2860_38778# 0.003766f
C31728 a_5934_30871# C7_N_btm 0.007575f
C31729 a_14955_47212# a_15811_47375# 1.55e-19
C31730 a_n1151_42308# a_n2312_39304# 2.72e-19
C31731 a_n1741_47186# a_8128_46384# 0.004988f
C31732 a_n971_45724# a_n1613_43370# 0.6298f
C31733 a_2063_45854# a_2747_46873# 0.023413f
C31734 a_6123_31319# C9_N_btm 9.33e-20
C31735 a_11599_46634# a_15507_47210# 0.267808f
C31736 a_13717_47436# a_16023_47582# 1.27e-19
C31737 a_12861_44030# a_16327_47482# 0.120085f
C31738 a_9313_45822# a_10227_46804# 1.42e-19
C31739 a_18727_42674# CAL_N 0.001564f
C31740 a_6151_47436# a_13507_46334# 7.34e-21
C31741 a_5742_30871# C7_P_btm 0.04157f
C31742 a_6773_42558# VDD 0.006434f
C31743 a_11341_43940# a_14205_43396# 0.001925f
C31744 a_7542_44172# a_743_42282# 2.49e-21
C31745 a_n89_45572# VDD 0.001196f
C31746 a_5891_43370# a_7309_43172# 0.002083f
C31747 a_14539_43914# a_13291_42460# 2.89e-21
C31748 a_n1352_43396# a_n447_43370# 4.88e-19
C31749 a_n2267_43396# a_n1809_43762# 0.034619f
C31750 a_n2433_43396# a_n1821_43396# 3.82e-19
C31751 a_15682_43940# a_15681_43442# 1.6e-19
C31752 a_20365_43914# a_10341_43396# 1.17e-20
C31753 a_5013_44260# a_4361_42308# 1.27e-20
C31754 a_11967_42832# a_10922_42852# 4.37e-20
C31755 a_n2956_37592# a_n2302_39866# 0.006499f
C31756 a_11823_42460# a_1307_43914# 0.049611f
C31757 a_15227_44166# a_14955_43940# 0.134177f
C31758 a_7227_45028# a_7418_45394# 2.88e-19
C31759 a_10907_45822# a_10775_45002# 1.92e-19
C31760 a_12465_44636# a_14621_43646# 1.9e-19
C31761 a_20107_45572# a_20528_45572# 0.086377f
C31762 a_20273_45572# a_21188_45572# 0.125324f
C31763 a_3090_45724# a_19328_44172# 0.153704f
C31764 a_16327_47482# a_19700_43370# 1.38e-19
C31765 a_n2293_46634# a_1427_43646# 2.05e-21
C31766 a_10903_43370# a_12189_44484# 1.63e-19
C31767 a_13249_42308# a_14537_43396# 0.020089f
C31768 a_14495_45572# a_14180_45002# 9.07e-19
C31769 a_5807_45002# a_8145_46902# 0.003883f
C31770 a_n2109_47186# a_n1076_46494# 1.12e-20
C31771 a_12549_44172# a_6755_46942# 0.553062f
C31772 a_11453_44696# a_14976_45028# 0.014048f
C31773 C7_P_btm C0_dummy_P_btm 0.120543f
C31774 C9_P_btm C0_N_btm 8.4e-19
C31775 C8_P_btm C0_dummy_N_btm 6.22e-19
C31776 a_14955_47212# a_13059_46348# 1.12e-19
C31777 a_11599_46634# a_15227_46910# 0.006776f
C31778 C6_P_btm C0_P_btm 0.140033f
C31779 C5_P_btm C1_P_btm 0.128021f
C31780 C4_P_btm C2_P_btm 7.19288f
C31781 a_n743_46660# a_3877_44458# 0.034265f
C31782 a_n2661_46634# a_5732_46660# 0.010632f
C31783 EN_VIN_BSTR_N C6_N_btm 0.118916f
C31784 a_n815_47178# a_n1853_46287# 4.63e-19
C31785 a_11031_47542# a_765_45546# 0.003176f
C31786 a_12861_44030# a_16434_46987# 0.001423f
C31787 a_13507_46334# a_19466_46812# 0.03247f
C31788 a_4883_46098# a_15227_44166# 0.176028f
C31789 a_21177_47436# a_19692_46634# 0.001012f
C31790 a_2107_46812# a_3524_46660# 0.004383f
C31791 a_948_46660# a_2864_46660# 3.21e-21
C31792 a_479_46660# a_n2661_46098# 3.93e-19
C31793 a_n1925_46634# a_4651_46660# 0.046762f
C31794 a_n1386_35608# VDD 0.360375f
C31795 a_n971_45724# a_n2293_46098# 0.110318f
C31796 a_10227_46804# a_12513_46660# 0.004052f
C31797 a_15811_47375# a_14543_46987# 2.63e-20
C31798 C10_P_btm C1_N_btm 0.001745f
C31799 a_n2661_42282# a_1606_42308# 0.082268f
C31800 a_3422_30871# a_15959_42545# 5.29e-20
C31801 a_8147_43396# a_8605_42826# 0.003157f
C31802 a_8791_43396# a_8037_42858# 0.001631f
C31803 a_11967_42832# a_17531_42308# 0.003854f
C31804 a_2304_45348# VDD 0.004463f
C31805 a_16977_43638# a_743_42282# 1.08e-20
C31806 a_15781_43660# a_5649_42852# 4.06e-21
C31807 a_15743_43084# a_16823_43084# 0.031733f
C31808 a_17499_43370# a_4190_30871# 2.22e-19
C31809 a_2382_45260# a_n2661_44458# 0.032484f
C31810 a_n467_45028# a_n1352_44484# 1.49e-19
C31811 a_8696_44636# a_n2293_43922# 0.002811f
C31812 a_n913_45002# a_5343_44458# 0.020508f
C31813 a_19692_46634# a_4361_42308# 0.004083f
C31814 a_15227_44166# a_5649_42852# 3.43e-20
C31815 a_15415_45028# a_16922_45042# 9.08e-21
C31816 a_16019_45002# a_16405_45348# 5.59e-19
C31817 a_1307_43914# a_16321_45348# 8.2e-20
C31818 a_n755_45592# a_3499_42826# 0.003508f
C31819 a_17339_46660# a_18429_43548# 0.033468f
C31820 a_n2312_40392# a_n3674_38680# 0.025175f
C31821 a_n2312_39304# a_n2840_42282# 3.28e-20
C31822 a_4185_45028# a_6293_42852# 1.35e-20
C31823 a_4185_45348# a_n2661_43370# 1.42e-19
C31824 a_n2293_46634# a_n1533_46116# 9.21e-21
C31825 a_5907_46634# a_5937_45572# 1.19e-19
C31826 a_n443_46116# a_2711_45572# 0.060543f
C31827 a_15227_44166# a_21188_46660# 3.62e-19
C31828 a_12549_44172# a_8049_45260# 0.031115f
C31829 a_n1741_47186# a_10053_45546# 8.64e-21
C31830 a_11901_46660# a_11415_45002# 1.07e-20
C31831 a_3090_45724# a_18280_46660# 4.52e-21
C31832 a_4883_46098# a_21071_46482# 1.62e-19
C31833 a_n1925_46634# a_n1379_46482# 3.89e-19
C31834 a_5807_45002# a_5066_45546# 0.027744f
C31835 a_n1151_42308# a_6511_45714# 0.044048f
C31836 a_n2438_43548# a_n2956_38680# 0.00293f
C31837 a_13507_46334# a_20205_31679# 0.023531f
C31838 a_11453_44696# a_18051_46116# 0.00399f
C31839 a_19692_46634# a_20841_46902# 0.025536f
C31840 a_22315_44484# VDD 0.213791f
C31841 a_17730_32519# C4_N_btm 6.79e-20
C31842 a_743_42282# a_n1630_35242# 0.004023f
C31843 a_10835_43094# a_11554_42852# 0.086334f
C31844 a_10518_42984# a_10752_42852# 0.006453f
C31845 a_10991_42826# a_11229_43218# 0.001705f
C31846 a_10796_42968# a_11301_43218# 2.28e-19
C31847 a_3422_30871# RST_Z 0.0872f
C31848 a_8685_43396# a_14113_42308# 5.76e-20
C31849 a_3626_43646# a_18220_42308# 9.35e-19
C31850 a_13467_32519# a_n784_42308# 0.014901f
C31851 a_n2840_42826# a_n3674_38680# 0.019613f
C31852 a_n2293_42282# a_3445_43172# 0.009537f
C31853 a_n2312_38680# a_n2302_39072# 0.00306f
C31854 a_5883_43914# a_9241_44734# 0.010354f
C31855 a_8701_44490# a_9313_44734# 5.25e-19
C31856 a_19778_44110# a_19615_44636# 0.012379f
C31857 a_18184_42460# a_11967_42832# 0.024012f
C31858 a_16922_45042# a_19279_43940# 0.018289f
C31859 a_3232_43370# a_10949_43914# 0.093316f
C31860 a_6171_45002# a_10729_43914# 2.56e-21
C31861 a_7499_43078# a_8685_43396# 0.153217f
C31862 a_3090_45724# a_8685_42308# 3.16e-21
C31863 a_20447_31679# a_14021_43940# 1.09e-20
C31864 a_10057_43914# a_5891_43370# 0.197199f
C31865 a_8975_43940# a_8375_44464# 2.42e-20
C31866 a_n1352_44484# a_n2661_43922# 0.007747f
C31867 a_n452_44636# a_n2661_42834# 0.002825f
C31868 a_n2293_42834# a_n1761_44111# 0.03111f
C31869 a_20193_45348# a_17517_44484# 0.015762f
C31870 a_11827_44484# a_16335_44484# 7.13e-19
C31871 a_8696_44636# a_n97_42460# 9.12e-22
C31872 a_n2109_47186# VDD 2.71791f
C31873 a_765_45546# a_n2293_45546# 7.13e-22
C31874 a_19321_45002# a_20273_45572# 1.46e-20
C31875 a_13747_46662# a_20623_45572# 4.02e-19
C31876 a_15928_47570# a_2437_43646# 0.003813f
C31877 a_4883_46098# a_4558_45348# 2.08e-20
C31878 a_13351_46090# a_6945_45028# 8.55e-21
C31879 a_4791_45118# a_5105_45348# 3.48e-19
C31880 a_12861_44030# a_14537_43396# 0.015677f
C31881 a_n1613_43370# a_n2293_45010# 0.077436f
C31882 a_12005_46116# a_10809_44734# 0.029593f
C31883 a_1823_45246# a_6347_46155# 7.53e-22
C31884 a_3699_46348# a_5066_45546# 1.54e-20
C31885 a_17583_46090# a_17957_46116# 0.092344f
C31886 a_17715_44484# a_18189_46348# 0.014348f
C31887 a_11599_46634# a_9482_43914# 8.71e-21
C31888 a_12549_44172# a_19479_31679# 1.37e-20
C31889 a_12891_46348# a_3357_43084# 6.59e-20
C31890 a_1755_42282# a_5379_42460# 0.045501f
C31891 a_2725_42558# a_2713_42308# 0.01129f
C31892 COMP_P a_5934_30871# 0.028728f
C31893 a_15597_42852# a_15051_42282# 3.4e-19
C31894 a_5205_44484# a_743_42282# 2.08e-20
C31895 a_n2017_45002# a_n967_43230# 3.36e-21
C31896 a_3357_43084# a_4520_42826# 5.54e-19
C31897 a_n699_43396# a_n2129_43609# 0.062898f
C31898 a_n967_45348# a_n1076_43230# 0.019022f
C31899 a_n2956_37592# a_n3674_39304# 0.023366f
C31900 a_n443_42852# a_1576_42282# 4.39e-21
C31901 a_n755_45592# a_3318_42354# 0.152654f
C31902 a_n357_42282# a_3823_42558# 1.45e-20
C31903 a_11823_42460# a_13003_42852# 0.002475f
C31904 a_n2810_45028# a_n4318_38680# 0.023185f
C31905 a_n1899_43946# a_644_44056# 2.13e-20
C31906 a_n1549_44318# a_n984_44318# 7.99e-20
C31907 a_n2661_45546# a_2277_45546# 0.00928f
C31908 a_18189_46348# a_15861_45028# 3.09e-20
C31909 a_10586_45546# a_10053_45546# 0.024917f
C31910 a_17715_44484# a_17478_45572# 0.017416f
C31911 a_15682_46116# a_16223_45938# 5.37e-19
C31912 a_2324_44458# a_12561_45572# 4.6e-19
C31913 a_12861_44030# a_20835_44721# 3.48e-19
C31914 a_n1613_43370# a_9313_44734# 3.6e-19
C31915 a_11453_44696# a_15433_44458# 9.82e-21
C31916 a_10227_46804# a_15367_44484# 5.42e-20
C31917 a_n1099_45572# a_n23_45546# 0.042611f
C31918 a_310_45028# a_n356_45724# 0.12349f
C31919 a_n1079_45724# a_n906_45572# 0.007688f
C31920 a_14513_46634# a_14180_45002# 8.73e-22
C31921 a_n746_45260# a_895_43940# 3.56e-19
C31922 a_n1853_46287# a_n2661_45010# 1.83e-20
C31923 a_20820_30879# en_comp 3.02e-19
C31924 a_n452_45724# a_7_45899# 6.64e-19
C31925 a_n863_45724# a_n1013_45572# 0.001771f
C31926 a_8049_45260# a_11525_45546# 0.002729f
C31927 a_13059_46348# a_13159_45002# 3.4e-19
C31928 a_n1151_42308# a_n2065_43946# 1.27e-19
C31929 a_584_46384# a_n984_44318# 1.54e-20
C31930 a_n755_45592# a_3316_45546# 0.045656f
C31931 a_19321_45002# a_18989_43940# 2.21e-19
C31932 a_n2293_46098# a_n2293_45010# 5.07e-19
C31933 COMP_P a_11530_34132# 0.018284f
C31934 a_n3565_39590# a_n3690_39616# 0.246863f
C31935 a_n4334_39616# a_n3420_39616# 0.015897f
C31936 a_n4209_39590# a_n2946_39866# 0.022704f
C31937 a_n971_45724# a_4791_45118# 0.025426f
C31938 a_1209_47178# a_n1151_42308# 0.024897f
C31939 a_584_46384# a_2553_47502# 0.100103f
C31940 a_n237_47217# a_4007_47204# 2.65e-20
C31941 a_n1741_47186# a_6151_47436# 0.071065f
C31942 a_2124_47436# a_2952_47436# 5.21e-19
C31943 a_6123_31319# a_n3420_37440# 0.00105f
C31944 a_n2661_42282# a_3539_42460# 1.44e-19
C31945 a_n2661_42834# a_n1641_43230# 9.58e-19
C31946 a_n2293_43922# a_n1991_42858# 0.007113f
C31947 a_5111_44636# a_7227_42308# 1.41e-20
C31948 a_3537_45260# a_8515_42308# 3.86e-22
C31949 a_8062_46155# VDD 2.63e-20
C31950 a_19279_43940# a_15743_43084# 6.64e-19
C31951 a_18579_44172# a_18429_43548# 6.43e-20
C31952 a_16789_44484# a_16823_43084# 4.65e-20
C31953 a_n356_44636# a_8952_43230# 4.57e-21
C31954 en_comp a_11323_42473# 4.34e-21
C31955 a_n913_45002# a_12563_42308# 1.51e-19
C31956 a_n1059_45260# a_13070_42354# 2.07e-20
C31957 a_n2017_45002# a_13575_42558# 0.006408f
C31958 a_2711_45572# a_3537_45260# 0.0026f
C31959 a_4099_45572# a_3065_45002# 3.74e-19
C31960 a_15861_45028# a_17478_45572# 0.080824f
C31961 a_8696_44636# a_16020_45572# 1.4e-20
C31962 a_12549_44172# a_15037_43940# 2.39e-20
C31963 a_2324_44458# a_2779_44458# 0.092751f
C31964 a_n2661_45546# a_626_44172# 0.002437f
C31965 a_13059_46348# a_11967_42832# 2.62e-19
C31966 a_9290_44172# a_10057_43914# 0.034053f
C31967 a_2107_46812# a_9801_44260# 9.76e-19
C31968 a_10227_46804# a_2982_43646# 6.99e-19
C31969 CAL_N a_22521_39511# 0.023597f
C31970 a_22469_40625# a_22459_39145# 0.245891f
C31971 a_n881_46662# a_33_46660# 0.002482f
C31972 a_6575_47204# a_6755_46942# 1.56e-19
C31973 a_n1435_47204# a_9863_46634# 2.27e-20
C31974 a_9313_45822# a_10467_46802# 0.009777f
C31975 a_n1613_43370# a_601_46902# 0.178721f
C31976 a_5807_45002# a_19321_45002# 0.376188f
C31977 a_n3420_37440# EN_VIN_BSTR_P 0.040234f
C31978 a_12891_46348# a_n2293_46634# 5.27e-20
C31979 a_8128_46384# a_n743_46660# 0.006641f
C31980 a_6151_47436# a_7832_46660# 0.016469f
C31981 a_2113_38308# VDD 0.004903f
C31982 a_14021_43940# a_17595_43084# 2.59e-21
C31983 a_15493_43940# a_21671_42860# 2.52e-21
C31984 a_11341_43940# a_22223_42860# 4.04e-19
C31985 a_14205_43396# a_10341_43396# 0.033299f
C31986 a_10695_43548# a_12281_43396# 5.09e-20
C31987 a_3357_43084# SINGLE_ENDED 0.131897f
C31988 a_22959_45572# VDD 0.304443f
C31989 a_4699_43561# a_4361_42308# 1.18e-20
C31990 a_3080_42308# a_13467_32519# 1.61e-19
C31991 a_19963_31679# RST_Z 0.050135f
C31992 a_8685_43396# a_15781_43660# 0.001931f
C31993 a_n97_42460# a_n1991_42858# 7.96e-21
C31994 a_n2129_43609# a_n4318_38680# 7.92e-19
C31995 a_n2267_43396# a_n3674_39304# 0.001257f
C31996 a_n1352_43396# a_n1641_43230# 0.001129f
C31997 a_n2012_43396# a_n2157_42858# 4.38e-19
C31998 a_n1177_43370# a_n901_43156# 0.002573f
C31999 a_9165_43940# a_8952_43230# 7.02e-20
C32000 a_2437_43646# DATA[1] 0.014934f
C32001 a_3775_45552# a_n2661_43922# 1.64e-20
C32002 a_n2661_45010# a_n2661_43370# 0.077441f
C32003 a_20841_45814# a_19778_44110# 7.65e-21
C32004 a_20107_45572# a_18494_42460# 0.010062f
C32005 a_n2293_46634# a_4520_42826# 4.07e-20
C32006 a_n2497_47436# a_n3674_37592# 2.17e-20
C32007 a_8270_45546# a_9885_43396# 4.58e-19
C32008 a_15227_44166# a_8685_43396# 0.013522f
C32009 a_3090_45724# a_9803_43646# 0.002871f
C32010 a_14976_45028# a_9145_43396# 4.71e-20
C32011 a_3483_46348# a_8487_44056# 5.36e-21
C32012 a_13348_45260# a_9482_43914# 0.352976f
C32013 a_13017_45260# a_13777_45326# 0.195607f
C32014 a_13159_45002# a_13556_45296# 0.006136f
C32015 a_n357_42282# a_20679_44626# 3.64e-21
C32016 a_10180_45724# a_5891_43370# 2.51e-20
C32017 a_7499_43078# a_8783_44734# 1.04e-19
C32018 a_526_44458# a_n2661_42282# 0.191497f
C32019 a_413_45260# a_2448_45028# 5.27e-19
C32020 a_17339_46660# a_2982_43646# 2.08e-20
C32021 SMPL_ON_P a_n961_42308# 1.43e-19
C32022 a_9290_44172# a_14021_43940# 0.003037f
C32023 a_6171_45002# a_1423_45028# 3.32e-19
C32024 a_13249_42308# a_n356_44636# 6.2e-20
C32025 a_8049_45260# a_7542_44172# 1.33e-20
C32026 a_12861_44030# a_12991_43230# 5.91e-20
C32027 a_10903_43370# a_12603_44260# 0.004294f
C32028 w_11334_34010# a_n1630_35242# 3.10971f
C32029 a_n2438_43548# a_791_42968# 4.47e-21
C32030 a_11453_44696# a_19900_46494# 3.8e-20
C32031 a_n2661_46634# a_1138_42852# 4.66e-20
C32032 a_768_44030# a_5937_45572# 0.05116f
C32033 a_6151_47436# a_10586_45546# 1.83e-20
C32034 a_6755_46942# a_10861_46660# 2.63e-19
C32035 a_n881_46662# a_12005_46116# 1.14e-20
C32036 a_11901_46660# a_12251_46660# 0.219633f
C32037 a_11735_46660# a_12816_46660# 0.102325f
C32038 a_11813_46116# a_12991_46634# 1.29e-20
C32039 a_22223_47212# a_6945_45028# 4.85e-19
C32040 a_12465_44636# a_22223_46124# 7.35e-21
C32041 a_n2438_43548# a_n1423_46090# 9.01e-21
C32042 a_6575_47204# a_8049_45260# 0.002085f
C32043 a_5732_46660# a_765_45546# 0.003297f
C32044 a_n1021_46688# a_n901_46420# 0.001157f
C32045 a_n1925_46634# a_n1076_46494# 0.003622f
C32046 a_4883_46098# a_22959_46124# 1.36e-19
C32047 a_21811_47423# a_10809_44734# 0.005196f
C32048 a_n1641_43230# a_n2293_42282# 1.64e-20
C32049 a_14021_43940# a_21887_42336# 5.15e-21
C32050 a_3539_42460# a_3497_42558# 0.002673f
C32051 a_16547_43609# a_17141_43172# 5.08e-20
C32052 a_10341_43396# a_22400_42852# 0.004171f
C32053 a_8375_44464# VDD 0.086619f
C32054 a_4905_42826# a_6481_42558# 1.25e-20
C32055 a_10518_42984# a_10922_42852# 0.051162f
C32056 a_10835_43094# a_10991_42826# 0.105839f
C32057 a_10083_42826# a_10341_42308# 0.001156f
C32058 a_13556_45296# a_11967_42832# 1.65e-21
C32059 a_18184_42460# a_18989_43940# 2.27e-20
C32060 a_4185_45028# a_10991_42826# 3.72e-20
C32061 a_12549_44172# a_13258_32519# 1.15e-21
C32062 a_16115_45572# a_15493_43940# 3.81e-20
C32063 a_10193_42453# a_19319_43548# 1.94e-20
C32064 a_n2661_44458# a_5343_44458# 0.003787f
C32065 a_n2661_45546# a_2813_43396# 2.3e-20
C32066 a_n913_45002# a_453_43940# 2.62e-21
C32067 a_n2661_45010# a_2998_44172# 5.85e-20
C32068 a_n2017_45002# a_2479_44172# 1.51e-20
C32069 a_n755_45592# a_6197_43396# 1.2e-20
C32070 SMPL_ON_P a_n3420_37440# 0.025729f
C32071 a_n443_42852# a_1987_43646# 8.61e-20
C32072 a_n1352_44484# a_n452_44636# 1.85e-19
C32073 a_11691_44458# a_15004_44636# 0.221929f
C32074 a_11827_44484# a_17767_44458# 0.014019f
C32075 a_n2312_39304# a_n2302_39866# 0.001835f
C32076 a_13661_43548# a_17303_42282# 9.85e-21
C32077 a_5937_45572# a_5755_42852# 6.93e-21
C32078 a_10227_46804# a_16789_45572# 1.86e-22
C32079 a_11415_45002# a_17583_46090# 2.43e-20
C32080 a_3483_46348# a_5164_46348# 0.025074f
C32081 a_22000_46634# a_10809_44734# 0.012475f
C32082 a_20731_47026# a_6945_45028# 0.001536f
C32083 a_9863_47436# a_2437_43646# 0.005338f
C32084 a_18597_46090# a_19431_45546# 0.062716f
C32085 a_11599_46634# a_20623_45572# 1.32e-21
C32086 a_n2661_46634# a_11962_45724# 0.020358f
C32087 a_n2109_47186# a_5691_45260# 0.113268f
C32088 a_n971_45724# a_3429_45260# 0.171338f
C32089 a_7903_47542# a_3357_43084# 1.35e-19
C32090 a_12741_44636# a_14840_46494# 9.71e-23
C32091 a_n743_46660# a_10053_45546# 3.51e-20
C32092 a_16327_47482# a_18787_45572# 9.38e-19
C32093 a_5342_30871# a_15720_42674# 9.9e-20
C32094 a_14401_32519# C6_N_btm 0.054459f
C32095 a_17538_32519# C4_N_btm 3.39e-20
C32096 a_20836_43172# a_20753_42852# 1.48e-19
C32097 a_19319_43548# VDD 0.561461f
C32098 a_16795_42852# a_15803_42450# 6.31e-20
C32099 a_8975_43940# a_10949_43914# 2.76e-19
C32100 a_10057_43914# a_10807_43548# 0.039192f
C32101 a_6109_44484# a_6453_43914# 0.165572f
C32102 a_n2293_43922# a_n1331_43914# 1.37e-19
C32103 a_n2661_42834# a_n809_44244# 0.021917f
C32104 a_n2661_43922# a_n1549_44318# 0.004791f
C32105 a_3363_44484# a_1414_42308# 1.44e-20
C32106 a_n2442_46660# CLK_DATA 0.063913f
C32107 a_11823_42460# a_13635_43156# 0.040348f
C32108 a_n357_42282# a_12800_43218# 0.002279f
C32109 a_n2661_46634# DATA[1] 1.37e-19
C32110 a_n2293_42834# a_n2267_43396# 0.010565f
C32111 a_1307_43914# a_2982_43646# 0.028987f
C32112 a_11967_42832# a_20362_44736# 0.052989f
C32113 a_19615_44636# a_20159_44458# 0.001766f
C32114 a_17517_44484# a_20596_44850# 3.5e-19
C32115 a_10193_42453# a_16795_42852# 1.71e-19
C32116 a_n1925_42282# a_5379_42460# 2.1e-20
C32117 a_n2956_39304# a_6123_31319# 4.63e-21
C32118 a_10903_43370# a_13657_42558# 2.45e-20
C32119 a_n1925_46634# VDD 0.783093f
C32120 a_20916_46384# EN_OFFSET_CAL 8.73e-21
C32121 a_4185_45028# a_17303_42282# 0.235259f
C32122 a_n1059_45260# a_8945_43396# 0.002485f
C32123 a_3537_45260# a_7466_43396# 1.01e-19
C32124 a_5111_44636# a_6643_43396# 0.004357f
C32125 a_13249_42308# a_12379_42858# 0.029761f
C32126 a_5066_45546# a_n755_45592# 4.16e-20
C32127 a_4791_45118# a_9313_44734# 5.17e-19
C32128 a_12861_44030# a_n356_44636# 4.56e-21
C32129 a_11415_45002# a_8696_44636# 0.10924f
C32130 a_4883_46098# a_9838_44484# 0.00188f
C32131 a_10227_46804# a_14539_43914# 0.012909f
C32132 a_3877_44458# a_2809_45348# 2.21e-20
C32133 a_19321_45002# a_18315_45260# 5.84e-20
C32134 a_10150_46912# a_8953_45002# 3.4e-19
C32135 a_6755_46942# a_5205_44484# 2.7e-19
C32136 a_13747_46662# a_18911_45144# 2.43e-19
C32137 a_13661_43548# a_19778_44110# 1.55e-19
C32138 a_19692_46634# a_20447_31679# 2.89e-20
C32139 a_12741_44636# a_16115_45572# 2.27e-20
C32140 a_3090_45724# a_n913_45002# 0.039732f
C32141 a_584_46384# a_n2661_43922# 0.0255f
C32142 a_2063_45854# a_n2661_42834# 0.022984f
C32143 a_12549_44172# a_20193_45348# 0.587618f
C32144 a_768_44030# a_11691_44458# 0.029945f
C32145 a_11189_46129# a_10053_45546# 1.92e-19
C32146 a_9290_44172# a_10180_45724# 0.037823f
C32147 a_10355_46116# a_10193_42453# 0.058019f
C32148 a_16327_47482# a_18287_44626# 0.552724f
C32149 a_6123_31319# a_n3565_39304# 4.63e-21
C32150 a_15959_42545# a_7174_31319# 4.42e-20
C32151 a_5934_30871# a_n4209_39304# 5.64e-21
C32152 COMP_P a_7754_40130# 1.45e-19
C32153 a_16795_42852# VDD 0.179044f
C32154 a_18579_44172# a_2982_43646# 1.56e-20
C32155 a_19478_44306# a_15493_43940# 0.025498f
C32156 a_1307_43914# a_5837_42852# 4.88e-20
C32157 a_n2956_38216# a_n3420_37984# 0.208204f
C32158 a_19479_31679# a_n1630_35242# 8.9e-20
C32159 a_n2810_45028# a_n2840_42282# 9.69e-21
C32160 a_10355_46116# VDD 0.222751f
C32161 a_n1352_44484# a_n1641_43230# 4.5e-21
C32162 a_n1177_44458# a_n901_43156# 7.62e-22
C32163 a_20269_44172# a_11341_43940# 0.006087f
C32164 a_20623_43914# a_20935_43940# 0.040559f
C32165 a_n984_44318# a_n1177_43370# 1.43e-19
C32166 a_n2017_45002# a_n2104_42282# 0.010745f
C32167 a_n2810_45572# a_n2302_37984# 0.130495f
C32168 a_10193_42453# a_21335_42336# 3.27e-20
C32169 a_n881_46662# a_15682_43940# 8.75e-21
C32170 a_2324_44458# a_7639_45394# 0.001717f
C32171 a_n1151_42308# a_n2129_43609# 0.019226f
C32172 a_584_46384# a_n447_43370# 1.6e-19
C32173 a_n2956_39768# a_n3674_39768# 0.023472f
C32174 a_n2293_46634# a_7281_43914# 7.08e-20
C32175 a_768_44030# a_8333_44056# 0.006943f
C32176 a_20692_30879# a_20447_31679# 9.02991f
C32177 a_17339_46660# a_14539_43914# 4.86e-21
C32178 a_10490_45724# a_10216_45572# 4.26e-20
C32179 a_8746_45002# a_10306_45572# 0.007074f
C32180 a_11823_42460# a_11682_45822# 4.41e-19
C32181 a_10903_43370# a_n2661_43370# 3.63e-19
C32182 a_11599_46634# a_13747_46662# 0.25325f
C32183 a_n3565_39304# EN_VIN_BSTR_P 2.04e-19
C32184 a_584_46384# a_1799_45572# 0.179456f
C32185 a_2124_47436# a_n2661_46098# 1.36e-19
C32186 a_n1151_42308# a_288_46660# 8.13e-19
C32187 a_6151_47436# a_n743_46660# 0.03019f
C32188 a_21335_42336# VDD 0.199586f
C32189 a_16023_47582# a_16285_47570# 0.001705f
C32190 a_16327_47482# a_16697_47582# 2.95e-19
C32191 a_7174_31319# RST_Z 0.216004f
C32192 a_n443_46116# a_33_46660# 1.22e-19
C32193 a_3785_47178# a_2107_46812# 2.1e-20
C32194 a_6491_46660# a_n1925_46634# 0.003135f
C32195 a_3754_39466# a_3754_38470# 7.8e-20
C32196 VDAC_Pi a_8530_39574# 1.79e-20
C32197 a_4958_30871# VCM 0.642743f
C32198 a_10227_46804# a_16119_47582# 0.004305f
C32199 a_15811_47375# a_5807_45002# 0.004711f
C32200 a_15673_47210# a_16131_47204# 0.034619f
C32201 a_n4064_39616# C7_P_btm 1.47e-19
C32202 a_n3420_39616# C5_P_btm 4.27e-20
C32203 a_n2109_47186# a_4646_46812# 0.021783f
C32204 a_3626_43646# a_8147_43396# 1.64e-21
C32205 a_2982_43646# a_9396_43370# 2.9e-20
C32206 a_14021_43940# a_13467_32519# 0.016437f
C32207 a_5883_43914# a_5934_30871# 1.2e-20
C32208 a_n356_44636# a_2123_42473# 1.17e-19
C32209 a_11967_42832# a_11554_42852# 9.86e-20
C32210 a_5343_44458# a_8325_42308# 0.014133f
C32211 a_n97_42460# a_14205_43396# 4.02e-21
C32212 a_12549_44172# a_20301_43646# 0.008227f
C32213 a_5907_45546# a_5343_44458# 1.37e-20
C32214 a_n967_45348# a_n143_45144# 1.34e-20
C32215 a_10227_46804# a_7871_42858# 7.12e-22
C32216 a_12861_44030# a_12379_42858# 2.07e-20
C32217 a_11415_45002# a_20365_43914# 2.15e-20
C32218 a_20202_43084# a_20623_43914# 1.77e-21
C32219 a_n2312_39304# a_n3674_39304# 0.023737f
C32220 a_n2312_40392# a_n4318_38680# 0.025333f
C32221 a_6511_45714# a_4223_44672# 1.22e-21
C32222 a_5257_43370# a_6293_42852# 0.001148f
C32223 a_5937_45572# a_7845_44172# 1.02e-19
C32224 a_n659_45366# a_n467_45028# 5.76e-19
C32225 a_n1059_45260# a_2382_45260# 0.025598f
C32226 a_11652_45724# a_11691_44458# 8.35e-19
C32227 a_310_45028# a_n356_44636# 2.32e-19
C32228 a_n1099_45572# a_n23_44458# 7.95e-21
C32229 a_3877_44458# a_6086_46660# 0.002133f
C32230 a_6151_47436# a_11189_46129# 7.98e-21
C32231 a_15928_47570# a_765_45546# 0.003038f
C32232 a_22959_47212# a_21076_30879# 0.002641f
C32233 SMPL_ON_P a_n2956_39304# 0.039212f
C32234 a_4915_47217# a_10903_43370# 0.004769f
C32235 a_6575_47204# a_8953_45546# 4.65e-19
C32236 a_9313_45822# a_8016_46348# 0.02464f
C32237 a_n1435_47204# a_6165_46155# 1.3e-20
C32238 a_9067_47204# a_5937_45572# 1.6e-19
C32239 a_16131_47204# a_16388_46812# 2.48e-19
C32240 a_12549_44172# a_18285_46348# 0.008787f
C32241 a_5807_45002# a_13059_46348# 0.1145f
C32242 a_2107_46812# a_3090_45724# 0.003997f
C32243 a_5257_43370# a_7577_46660# 4.41e-20
C32244 a_4817_46660# a_6969_46634# 5.31e-20
C32245 a_7411_46660# a_7715_46873# 0.162909f
C32246 a_n971_45724# a_6945_45028# 0.247957f
C32247 a_n2497_47436# a_n967_46494# 7.99e-21
C32248 a_16243_43396# a_16414_43172# 9.71e-20
C32249 a_743_42282# a_4520_42826# 5.99e-20
C32250 a_16137_43396# a_16795_42852# 0.010001f
C32251 a_18114_32519# C5_N_btm 1.78e-19
C32252 a_19721_31679# C4_N_btm 9.91e-21
C32253 a_n1423_42826# a_n1641_43230# 0.209641f
C32254 a_n2157_42858# a_n13_43084# 9.69e-21
C32255 a_n1991_42858# a_n901_43156# 0.041762f
C32256 a_n1853_43023# a_n1076_43230# 0.040291f
C32257 a_n2472_42826# a_n3674_39304# 7.06e-19
C32258 a_10341_43396# a_22223_42860# 2.12e-20
C32259 a_3422_30871# a_n4064_39072# 0.007014f
C32260 a_17801_45144# VDD 2.88e-19
C32261 a_n2840_42826# a_n4318_38680# 0.044261f
C32262 a_n2840_43370# a_n4318_38216# 0.003324f
C32263 a_n2442_46660# a_n1630_35242# 0.02547f
C32264 SMPL_ON_P a_n3565_39304# 0.001067f
C32265 a_n443_42852# a_1241_43940# 3.12e-20
C32266 a_n1613_43370# a_8515_42308# 7.89e-20
C32267 a_5205_44484# a_5289_44734# 0.011388f
C32268 a_526_44458# a_7112_43396# 9.09e-20
C32269 a_3537_45260# a_9241_44734# 1.1e-21
C32270 a_20107_45572# a_20640_44752# 3.77e-19
C32271 a_20273_45572# a_20362_44736# 1.1e-20
C32272 a_18587_45118# a_19778_44110# 1.74e-20
C32273 a_16922_45042# a_21101_45002# 2.6e-19
C32274 a_n967_45348# a_n2293_43922# 0.001623f
C32275 a_n2312_39304# a_5742_30871# 6.2e-21
C32276 a_21363_45546# a_11967_42832# 3.52e-22
C32277 a_9290_44172# a_13943_43396# 0.003427f
C32278 a_16327_47482# a_17124_42282# 1.39e-20
C32279 a_n913_45002# a_14815_43914# 9.21e-19
C32280 a_10193_42453# a_10949_43914# 0.032349f
C32281 a_3232_43370# a_7640_43914# 1.47e-19
C32282 a_6171_45002# a_6109_44484# 1.77e-19
C32283 a_1307_43914# a_14539_43914# 0.131617f
C32284 a_15227_44166# a_17333_42852# 0.043277f
C32285 a_n2442_46660# a_n2661_45546# 6.66e-19
C32286 a_n2293_46634# a_n2810_45572# 5.41e-20
C32287 a_12816_46660# a_2324_44458# 1.64e-21
C32288 a_14976_45028# a_13925_46122# 1.92e-19
C32289 a_5257_43370# a_5431_46482# 9.25e-20
C32290 a_768_44030# a_n443_42852# 0.00732f
C32291 a_n2661_46634# a_n2956_38216# 3.93e-19
C32292 a_22365_46825# a_20202_43084# 0.115624f
C32293 a_4883_46098# a_8568_45546# 1.93e-19
C32294 a_10227_46804# a_12427_45724# 6.03e-20
C32295 a_n1613_43370# a_2711_45572# 0.028041f
C32296 a_16388_46812# a_3483_46348# 4.06e-21
C32297 a_765_45546# a_1138_42852# 0.02041f
C32298 a_15368_46634# a_13759_46122# 1.21e-20
C32299 a_743_42282# a_15720_42674# 1.14e-19
C32300 a_15743_43084# a_19332_42282# 1.97e-20
C32301 a_10949_43914# VDD 0.797824f
C32302 a_3080_42308# a_2113_38308# 1.02e-19
C32303 a_4361_42308# a_15486_42560# 0.005067f
C32304 a_n443_42852# a_5755_42852# 0.008806f
C32305 a_20894_47436# VDD 0.188358f
C32306 a_19787_47423# RST_Z 5.42e-20
C32307 a_n967_45348# a_n97_42460# 3.72e-20
C32308 a_18989_43940# a_20362_44736# 5.76e-19
C32309 a_17767_44458# a_18005_44484# 0.007399f
C32310 a_11649_44734# a_n2661_43922# 1.92e-19
C32311 a_n1177_44458# a_n984_44318# 1.7e-20
C32312 a_2437_43646# a_1987_43646# 2.32e-21
C32313 a_19386_47436# START 0.042951f
C32314 a_21588_30879# VDAC_N 0.001941f
C32315 a_9313_44734# a_10809_44484# 1.08e-19
C32316 a_14539_43914# a_18579_44172# 3.18e-21
C32317 a_n2661_45010# a_1568_43370# 5.03e-22
C32318 a_n357_42282# a_10341_42308# 0.057131f
C32319 a_1307_43914# a_2253_43940# 0.056967f
C32320 a_10227_46804# a_14309_45028# 8.79e-19
C32321 a_11599_46634# a_18911_45144# 1.61e-20
C32322 a_17583_46090# a_13259_45724# 0.191869f
C32323 a_n2293_46098# a_2711_45572# 0.530463f
C32324 a_1176_45822# a_n443_42852# 0.071187f
C32325 a_n2661_46634# a_7229_43940# 2.93e-22
C32326 a_n1151_42308# a_n2129_44697# 0.039834f
C32327 a_13059_46348# a_15143_45578# 0.262261f
C32328 a_13661_43548# a_9482_43914# 0.127225f
C32329 a_5807_45002# a_13556_45296# 0.017285f
C32330 a_3147_46376# a_3503_45724# 5.03e-19
C32331 a_3483_46348# a_3316_45546# 1.91e-21
C32332 a_n1925_46634# a_5691_45260# 1.67e-21
C32333 a_14976_45028# a_15599_45572# 5.65e-21
C32334 a_3090_45724# a_15903_45785# 0.006612f
C32335 a_4817_46660# a_3357_43084# 0.005952f
C32336 a_12861_44030# a_20567_45036# 3.84e-21
C32337 a_16327_47482# a_17023_45118# 0.006152f
C32338 a_4883_46098# a_n2661_43370# 0.022462f
C32339 a_5907_46634# a_2437_43646# 7.11e-20
C32340 a_n2661_46098# a_n967_45348# 2.74e-21
C32341 a_2107_46812# a_2274_45254# 2.87e-19
C32342 a_n743_46660# a_5111_44636# 7.53e-20
C32343 a_n971_45724# a_8103_44636# 0.003603f
C32344 a_768_44030# a_375_42282# 3.77e-19
C32345 a_14493_46090# a_15002_46116# 2.6e-19
C32346 a_17364_32525# C1_N_btm 9.59e-21
C32347 a_9223_42460# a_5742_30871# 8.72e-20
C32348 a_n3674_38680# a_n4064_40160# 0.022279f
C32349 a_13887_32519# C5_N_btm 1.01e-19
C32350 a_19095_43396# VDD 0.003529f
C32351 a_11827_44484# a_18525_43370# 8.62e-21
C32352 a_9482_43914# a_10835_43094# 1.01e-21
C32353 a_20411_46873# VDD 0.348821f
C32354 a_7845_44172# a_8333_44056# 0.065494f
C32355 a_20107_46660# RST_Z 1.12e-20
C32356 a_n913_45002# a_945_42968# 0.001032f
C32357 a_n1059_45260# a_1709_42852# 4.99e-19
C32358 a_22315_44484# a_14021_43940# 2.03e-21
C32359 a_11691_44458# a_16759_43396# 3.94e-20
C32360 a_n2293_42834# a_n2472_42826# 0.199703f
C32361 a_1307_43914# a_7871_42858# 9.1e-21
C32362 a_n2293_43922# a_n1917_43396# 3.53e-21
C32363 a_n2661_42834# a_n1352_43396# 0.005746f
C32364 a_765_45546# DATA[1] 0.009245f
C32365 a_n357_42282# a_18057_42282# 5.64e-20
C32366 a_7499_43078# a_6123_31319# 0.002947f
C32367 a_2711_45572# a_7230_45938# 0.004731f
C32368 a_19321_45002# a_19006_44850# 1.35e-20
C32369 a_13259_45724# a_8696_44636# 0.259609f
C32370 a_3090_45724# a_n2661_44458# 0.088502f
C32371 a_1823_45246# a_1307_43914# 0.013371f
C32372 a_3483_46348# a_13777_45326# 0.027519f
C32373 a_n2293_46098# a_4640_45348# 1.74e-19
C32374 a_9569_46155# a_6171_45002# 6.04e-21
C32375 a_15227_44166# a_18545_45144# 0.002275f
C32376 a_16388_46812# a_17719_45144# 5.03e-21
C32377 a_12549_44172# a_20596_44850# 2.61e-19
C32378 a_8049_45260# a_19431_45546# 0.006516f
C32379 a_13661_43548# a_20159_44458# 1.06e-19
C32380 a_7920_46348# a_8191_45002# 1.55e-20
C32381 a_8199_44636# a_7229_43940# 1.98e-19
C32382 a_5937_45572# a_7276_45260# 0.052629f
C32383 a_16375_45002# a_16115_45572# 1.66e-19
C32384 a_14840_46494# a_413_45260# 2.43e-21
C32385 a_18057_42282# CAL_N 3.79e-19
C32386 a_n4064_38528# a_n2302_38778# 0.239588f
C32387 a_n4334_38528# a_n4251_38528# 0.007692f
C32388 a_n2946_38778# a_n2860_38778# 0.011479f
C32389 a_n4209_38502# a_n3607_38528# 0.002294f
C32390 a_6481_42558# VDD 0.006426f
C32391 a_5934_30871# C6_N_btm 0.004563f
C32392 a_n1151_42308# a_n2312_40392# 1.57e-19
C32393 a_5932_42308# RST_Z 0.005263f
C32394 a_n1741_47186# a_5159_47243# 1.44e-19
C32395 a_n815_47178# a_n881_46662# 2.82e-20
C32396 a_584_46384# a_2747_46873# 2.14e-19
C32397 a_2063_45854# a_2487_47570# 0.003691f
C32398 a_1209_47178# a_3315_47570# 4.55e-20
C32399 a_6123_31319# C8_N_btm 6.73e-20
C32400 a_14955_47212# a_15507_47210# 5.87e-19
C32401 a_14311_47204# a_15811_47375# 6.14e-21
C32402 a_4915_47217# a_4883_46098# 0.024005f
C32403 a_13717_47436# a_16327_47482# 2.02e-19
C32404 a_12861_44030# a_16241_47178# 3e-20
C32405 a_17303_42282# a_22469_40625# 4.4e-19
C32406 a_11031_47542# a_10227_46804# 3.37e-19
C32407 a_5742_30871# C8_P_btm 0.003514f
C32408 a_11341_43940# a_14358_43442# 1.43e-20
C32409 a_5244_44056# a_4361_42308# 2.42e-21
C32410 a_n2472_43914# a_n4318_38680# 5.56e-21
C32411 a_n1899_43946# a_n1076_43230# 5.62e-21
C32412 a_n1549_44318# a_n1641_43230# 1.17e-21
C32413 a_n4318_40392# a_n4318_38216# 0.023287f
C32414 a_n310_45572# VDD 7.01e-20
C32415 a_n2810_45028# a_n2302_39866# 4.97e-19
C32416 a_14673_44172# a_15567_42826# 4.79e-22
C32417 a_5891_43370# a_6101_43172# 0.003606f
C32418 a_n1177_43370# a_n447_43370# 0.010921f
C32419 a_n2267_43396# a_n2012_43396# 0.064178f
C32420 a_5829_43940# a_6031_43396# 3.18e-19
C32421 a_20269_44172# a_10341_43396# 3.22e-20
C32422 a_n2956_37592# a_n4064_39616# 0.015429f
C32423 a_11967_42832# a_10991_42826# 7.44e-20
C32424 a_8049_45260# a_13076_44458# 2.05e-21
C32425 a_n357_42282# a_18494_42460# 0.033084f
C32426 a_16327_47482# a_19268_43646# 0.024286f
C32427 a_15227_44166# a_13483_43940# 1.48e-20
C32428 a_n971_45724# a_n722_43218# 3.38e-19
C32429 a_8746_45002# a_1423_45028# 2.1e-19
C32430 a_10907_45822# a_8953_45002# 1.29e-20
C32431 a_20107_45572# a_21188_45572# 0.102355f
C32432 a_20273_45572# a_21363_45546# 0.042415f
C32433 a_20841_45814# a_20623_45572# 0.209641f
C32434 a_3090_45724# a_18451_43940# 0.004024f
C32435 a_n1613_43370# a_7466_43396# 0.001965f
C32436 a_15143_45578# a_13556_45296# 9.68e-20
C32437 a_13249_42308# a_14180_45002# 0.014749f
C32438 a_6755_46942# a_15301_44260# 1.12e-19
C32439 a_5807_45002# a_7577_46660# 0.003957f
C32440 a_n2109_47186# a_n901_46420# 9.56e-21
C32441 a_12891_46348# a_6755_46942# 0.025465f
C32442 a_12861_44030# a_16721_46634# 0.070721f
C32443 a_11453_44696# a_3090_45724# 0.232756f
C32444 a_12465_44636# a_16292_46812# 2.02e-20
C32445 C8_P_btm C0_dummy_P_btm 0.236317f
C32446 C9_P_btm C0_dummy_N_btm 7.47e-19
C32447 C6_P_btm C1_P_btm 0.128559f
C32448 C7_P_btm C0_P_btm 0.142187f
C32449 C4_P_btm C3_P_btm 7.90108f
C32450 C5_P_btm C2_P_btm 0.138678f
C32451 a_n2661_46634# a_5907_46634# 0.006487f
C32452 EN_VIN_BSTR_N C5_N_btm 0.115337f
C32453 a_9863_47436# a_765_45546# 0.001205f
C32454 a_20990_47178# a_19692_46634# 1.02e-20
C32455 a_14311_47204# a_13059_46348# 7.47e-21
C32456 a_2107_46812# a_3699_46634# 0.004263f
C32457 a_601_46902# a_1057_46660# 4.2e-19
C32458 a_1110_47026# a_n2661_46098# 3.75e-20
C32459 a_n1925_46634# a_4646_46812# 0.089593f
C32460 a_n1838_35608# VDD 0.523851f
C32461 a_13507_46334# a_19333_46634# 0.009057f
C32462 a_10227_46804# a_12347_46660# 0.004629f
C32463 a_15811_47375# a_14226_46987# 2.43e-21
C32464 C10_P_btm C0_N_btm 0.00154f
C32465 a_19862_44208# a_20753_42852# 0.008633f
C32466 a_3422_30871# a_15803_42450# 1.13e-19
C32467 a_18494_42460# CAL_N 0.001361f
C32468 a_2982_43646# a_13635_43156# 1.77e-19
C32469 a_3626_43646# a_13113_42826# 5.26e-21
C32470 a_8147_43396# a_8037_42858# 3.54e-19
C32471 a_11967_42832# a_17303_42282# 0.058225f
C32472 a_16409_43396# a_743_42282# 8.5e-21
C32473 a_18783_43370# a_16823_43084# 5.12e-19
C32474 a_2274_45254# a_n2661_44458# 8.17e-20
C32475 a_8696_44636# a_n2661_43922# 0.257466f
C32476 a_327_44734# a_n2129_44697# 0.00201f
C32477 a_n467_45028# a_n1177_44458# 0.001271f
C32478 a_n1059_45260# a_5343_44458# 0.019826f
C32479 a_19692_46634# a_13467_32519# 0.015407f
C32480 a_16019_45002# a_16321_45348# 0.002468f
C32481 a_n357_42282# a_3499_42826# 0.007965f
C32482 a_n745_45366# a_n699_43396# 2.06e-22
C32483 a_17339_46660# a_17324_43396# 6.45e-20
C32484 a_3483_46348# a_6197_43396# 8.08e-22
C32485 a_n2312_40392# a_n2840_42282# 4.5e-20
C32486 a_10193_42453# a_3422_30871# 0.404849f
C32487 a_4185_45028# a_6031_43396# 4.43e-21
C32488 a_2711_45572# a_2675_43914# 1.32e-20
C32489 a_n2438_43548# a_n2956_39304# 0.014879f
C32490 a_4791_45118# a_2711_45572# 0.160646f
C32491 a_n443_46116# a_1609_45572# 2.27e-19
C32492 a_15227_44166# a_21363_46634# 1.47e-19
C32493 a_14513_46634# a_16388_46812# 2.55e-21
C32494 a_12891_46348# a_8049_45260# 0.035062f
C32495 a_11813_46116# a_11415_45002# 4.47e-21
C32496 a_3090_45724# a_17639_46660# 5.38e-20
C32497 a_4883_46098# a_20850_46482# 2.25e-19
C32498 a_n1925_46634# a_n1545_46494# 6.83e-19
C32499 a_2063_45854# a_3775_45552# 1.46e-19
C32500 a_n1151_42308# a_6472_45840# 0.01357f
C32501 a_4007_47204# a_4099_45572# 4.68e-19
C32502 a_n971_45724# a_6812_45938# 1.09e-19
C32503 a_19692_46634# a_20273_46660# 0.02419f
C32504 a_3422_30871# VDD 1.12305f
C32505 a_17730_32519# C3_N_btm 5.52e-20
C32506 a_10922_42852# a_10793_43218# 4.2e-19
C32507 a_10835_43094# a_11301_43218# 3.82e-19
C32508 a_3626_43646# a_18214_42558# 5.05e-20
C32509 a_743_42282# a_564_42282# 0.169821f
C32510 a_n2840_42826# a_n2840_42282# 0.025171f
C32511 a_19237_31679# C1_N_btm 0.001047f
C32512 a_n2312_38680# a_n4064_39072# 0.002525f
C32513 a_19778_44110# a_11967_42832# 0.024799f
C32514 a_3232_43370# a_10729_43914# 0.090148f
C32515 a_n443_42852# a_16759_43396# 1.02e-20
C32516 a_7499_43078# a_6809_43396# 1.07e-19
C32517 a_20202_43084# a_14097_32519# 7.09e-21
C32518 a_10440_44484# a_5891_43370# 0.001688f
C32519 a_8103_44636# a_9313_44734# 1.28e-19
C32520 a_n1177_44458# a_n2661_43922# 0.010791f
C32521 a_n1352_44484# a_n2661_42834# 0.002886f
C32522 a_n2293_42834# a_n2065_43946# 9.75e-19
C32523 a_11691_44458# a_17517_44484# 0.058911f
C32524 a_20692_30879# a_13467_32519# 0.051714f
C32525 a_11827_44484# a_16241_44484# 6.75e-19
C32526 a_8975_43940# a_7640_43914# 1.34e-20
C32527 a_n699_43396# a_3363_44484# 0.07346f
C32528 a_18479_45785# a_19319_43548# 0.102555f
C32529 a_18175_45572# a_18533_43940# 1.04e-21
C32530 a_n2288_47178# VDD 0.29372f
C32531 a_17583_46090# a_18189_46348# 7.78e-19
C32532 a_3090_45724# a_5907_45546# 4.4e-21
C32533 a_19321_45002# a_20107_45572# 0.006336f
C32534 a_13747_46662# a_20841_45814# 1.63e-19
C32535 a_768_44030# a_2437_43646# 0.137571f
C32536 a_12594_46348# a_6945_45028# 5.55e-20
C32537 a_2063_45854# a_5093_45028# 1.55e-21
C32538 a_n743_46660# a_16147_45260# 0.071228f
C32539 a_n881_46662# a_n2661_45010# 1.04e-19
C32540 a_10903_43370# a_10809_44734# 0.353301f
C32541 a_3483_46348# a_5066_45546# 0.081087f
C32542 a_11309_47204# a_3357_43084# 8.86e-21
C32543 a_1755_42282# a_5267_42460# 2.48e-19
C32544 a_1606_42308# a_5379_42460# 9.76e-20
C32545 a_n443_42852# a_1067_42314# 0.011239f
C32546 a_n2810_45028# a_n3674_39304# 0.023324f
C32547 a_n913_45002# a_n1736_43218# 7.53e-21
C32548 a_13720_44458# a_13565_43940# 6.18e-20
C32549 a_n1352_44484# a_n1352_43396# 1.58e-19
C32550 a_6999_46987# VDD 2.18e-20
C32551 a_5111_44636# a_4361_42308# 0.009091f
C32552 a_n2017_45002# a_n1379_43218# 2.45e-19
C32553 a_3357_43084# a_3935_42891# 0.025181f
C32554 a_n699_43396# a_n2433_43396# 1.5e-20
C32555 a_n967_45348# a_n901_43156# 0.002872f
C32556 en_comp a_n1076_43230# 4.2e-20
C32557 a_n357_42282# a_3318_42354# 1.18e-20
C32558 a_n755_45592# a_2903_42308# 0.070479f
C32559 a_10193_42453# a_18504_43218# 0.003216f
C32560 a_n1899_43946# a_175_44278# 6.25e-20
C32561 a_n1331_43914# a_n984_44318# 0.051162f
C32562 a_19321_45002# a_18374_44850# 1.39e-20
C32563 a_n2661_45546# a_1609_45822# 0.02204f
C32564 a_18189_46348# a_8696_44636# 2.18e-21
C32565 a_17715_44484# a_15861_45028# 0.184272f
C32566 a_17583_46090# a_17478_45572# 3.05e-19
C32567 a_15682_46116# a_16020_45572# 3.39e-19
C32568 a_12861_44030# a_20679_44626# 8.93e-19
C32569 a_11453_44696# a_14815_43914# 6.62e-20
C32570 a_10227_46804# a_15146_44484# 2.64e-22
C32571 a_380_45546# a_n23_45546# 0.002746f
C32572 a_n1099_45572# a_n356_45724# 0.070228f
C32573 a_n1079_45724# a_n1013_45572# 0.010598f
C32574 a_6945_45028# a_15037_45618# 3.02e-21
C32575 a_10586_45546# a_9049_44484# 0.002146f
C32576 a_14180_46812# a_14180_45002# 1.22e-20
C32577 a_12594_46348# a_14127_45572# 6.01e-19
C32578 a_n237_47217# a_2127_44172# 3.02e-21
C32579 a_8128_46384# a_5891_43370# 1.23e-21
C32580 a_n452_45724# a_n310_45899# 0.005572f
C32581 a_8049_45260# a_11322_45546# 0.004301f
C32582 a_13059_46348# a_13017_45260# 0.022433f
C32583 a_n755_45592# a_3218_45724# 0.045755f
C32584 a_18479_47436# a_17517_44484# 0.017833f
C32585 a_n2157_46122# a_n2661_45010# 4.29e-20
C32586 a_n2293_46098# a_n2472_45002# 0.001044f
C32587 a_18504_43218# VDD 0.077608f
C32588 a_n4209_39590# a_n3420_39616# 0.234699f
C32589 a_584_46384# a_2063_45854# 0.406382f
C32590 a_n971_45724# a_4700_47436# 8.66e-19
C32591 a_327_47204# a_n1151_42308# 0.013822f
C32592 a_n237_47217# a_3815_47204# 1.74e-20
C32593 a_n1741_47186# a_5815_47464# 0.021904f
C32594 a_1209_47178# a_3160_47472# 1.39e-19
C32595 a_n2302_40160# a_n2302_39866# 0.050477f
C32596 a_n4334_39616# a_n3690_39616# 8.67e-19
C32597 a_4958_30871# a_n4064_38528# 0.030901f
C32598 a_14021_43940# a_19319_43548# 0.026713f
C32599 a_n2661_42282# a_3626_43646# 0.02843f
C32600 a_n2293_43922# a_n1853_43023# 0.001113f
C32601 a_n2661_42834# a_n1423_42826# 7.48e-19
C32602 a_1307_43914# a_1184_42692# 2.31e-21
C32603 a_3537_45260# a_5934_30871# 9.2e-20
C32604 a_5111_44636# a_6761_42308# 2.87e-20
C32605 a_3065_45002# a_3905_42308# 0.001599f
C32606 a_3422_30871# a_16137_43396# 2.61e-20
C32607 a_n356_44636# a_9127_43156# 1.19e-19
C32608 a_626_44172# a_564_42282# 2.14e-19
C32609 en_comp a_10723_42308# 8.68e-21
C32610 a_n1059_45260# a_12563_42308# 5.81e-20
C32611 a_n2017_45002# a_13070_42354# 0.002239f
C32612 a_n913_45002# a_11633_42558# 1.3e-20
C32613 a_13720_44458# a_5534_30871# 6.17e-22
C32614 a_9290_44172# a_10440_44484# 5.93e-21
C32615 a_8696_44636# a_17478_45572# 0.185985f
C32616 a_12549_44172# a_13565_43940# 4.78e-21
C32617 a_2324_44458# a_949_44458# 0.323116f
C32618 a_n2661_45546# a_501_45348# 1.17e-19
C32619 a_2711_45572# a_3429_45260# 9.02e-20
C32620 a_2107_46812# a_9248_44260# 1.38e-19
C32621 a_22521_40599# a_22459_39145# 1.41583f
C32622 a_22469_40625# a_22521_40055# 0.076632f
C32623 a_n4064_38528# VCM 0.007464f
C32624 a_9804_47204# a_n1925_46634# 9.26e-22
C32625 a_n881_46662# a_171_46873# 0.018745f
C32626 a_11031_47542# a_10467_46802# 1.42e-19
C32627 a_7903_47542# a_6755_46942# 9.91e-21
C32628 a_9313_45822# a_10428_46928# 1.12e-19
C32629 a_n1613_43370# a_33_46660# 0.599895f
C32630 a_n2302_37690# a_n1838_35608# 5.27e-19
C32631 a_n3420_37440# a_n923_35174# 0.002091f
C32632 a_768_44030# a_n2661_46634# 5.84e-20
C32633 a_13661_43548# a_13747_46662# 0.095862f
C32634 a_2063_45854# a_11901_46660# 0.001041f
C32635 a_n3607_38304# VDD 2.79e-20
C32636 a_3422_30871# a_n784_42308# 0.022792f
C32637 a_3357_43084# START 0.045418f
C32638 a_15493_43940# a_21195_42852# 2.39e-21
C32639 a_11341_43940# a_22165_42308# 0.003146f
C32640 a_3626_43646# a_16823_43084# 1.31e-20
C32641 a_14358_43442# a_10341_43396# 0.00838f
C32642 a_22591_45572# RST_Z 5.34e-19
C32643 a_9313_44734# a_14456_42282# 6.48e-20
C32644 a_n356_44636# a_17124_42282# 0.025455f
C32645 a_19963_31679# VDD 0.605279f
C32646 a_4235_43370# a_4361_42308# 0.006227f
C32647 a_15095_43370# a_14955_43396# 0.130374f
C32648 a_8685_43396# a_15681_43442# 0.002304f
C32649 a_n2840_43914# a_n3674_38680# 0.001131f
C32650 a_n1557_42282# a_743_42282# 2.06e-19
C32651 a_n97_42460# a_n1853_43023# 0.151542f
C32652 a_n1177_43370# a_n1641_43230# 0.003712f
C32653 a_n2433_43396# a_n4318_38680# 0.001035f
C32654 a_n2129_43609# a_n3674_39304# 4.16e-19
C32655 a_9165_43940# a_9127_43156# 8.16e-20
C32656 a_20447_31679# C10_N_btm 2.25e-20
C32657 a_2437_43646# DATA[0] 9.16e-20
C32658 a_3775_45552# a_n2661_42834# 3.12e-21
C32659 a_n2840_45002# a_n2661_43370# 0.005868f
C32660 a_20107_45572# a_18184_42460# 0.001559f
C32661 a_20273_45572# a_19778_44110# 3.15e-20
C32662 a_n2293_46634# a_3935_42891# 4.54e-20
C32663 a_12549_44172# a_5534_30871# 2.57e-20
C32664 SMPL_ON_P a_n1329_42308# 4.56e-20
C32665 a_2324_44458# a_11341_43940# 0.007112f
C32666 a_3090_45724# a_9145_43396# 0.189557f
C32667 a_13159_45002# a_9482_43914# 0.020865f
C32668 a_13017_45260# a_13556_45296# 0.049621f
C32669 a_10053_45546# a_5891_43370# 3.54e-20
C32670 a_19256_45572# a_11691_44458# 0.001053f
C32671 a_3232_43370# a_1423_45028# 0.396815f
C32672 a_10903_43370# a_12495_44260# 0.001658f
C32673 a_6755_46942# a_16409_43396# 6.64e-20
C32674 a_11453_44696# a_20075_46420# 2.89e-20
C32675 a_768_44030# a_8199_44636# 0.026637f
C32676 a_n2293_46634# a_472_46348# 1.43e-21
C32677 a_n2661_46634# a_1176_45822# 4.24e-19
C32678 a_6755_46942# a_12359_47026# 8.58e-19
C32679 a_10554_47026# a_10933_46660# 3.16e-19
C32680 a_10249_46116# a_10861_46660# 3.67e-19
C32681 a_11735_46660# a_12991_46634# 0.043475f
C32682 a_11901_46660# a_12469_46902# 0.175891f
C32683 a_11813_46116# a_12251_46660# 3.12e-19
C32684 a_n881_46662# a_10903_43370# 3.24e-19
C32685 a_12465_44636# a_6945_45028# 0.023497f
C32686 a_171_46873# a_n2157_46122# 3.28e-21
C32687 a_33_46660# a_n2293_46098# 1.87e-20
C32688 a_13747_46662# a_4185_45028# 2.24e-20
C32689 a_7903_47542# a_8049_45260# 2.11e-20
C32690 a_n2833_47464# a_n2840_45546# 3.38e-21
C32691 a_n1925_46634# a_n901_46420# 0.004832f
C32692 a_n2438_43548# a_n1991_46122# 0.001576f
C32693 a_5907_46634# a_765_45546# 0.003106f
C32694 a_4883_46098# a_10809_44734# 0.068164f
C32695 a_7640_43914# VDD 0.196713f
C32696 a_n1423_42826# a_n2293_42282# 3.12e-20
C32697 a_2982_43646# a_3905_42558# 4.96e-19
C32698 a_16547_43609# a_16877_43172# 9.85e-19
C32699 a_16137_43396# a_18504_43218# 0.002301f
C32700 a_4905_42826# a_5932_42308# 0.058059f
C32701 a_10518_42984# a_10991_42826# 7.99e-20
C32702 a_10835_43094# a_10796_42968# 0.671797f
C32703 a_9482_43914# a_11967_42832# 3.07e-21
C32704 a_11827_44484# a_16979_44734# 0.012885f
C32705 a_19778_44110# a_18989_43940# 6.83e-20
C32706 a_3357_43084# a_6453_43914# 4.6e-20
C32707 a_4185_45028# a_10796_42968# 3.58e-20
C32708 a_n755_45592# a_6293_42852# 2.52e-20
C32709 a_n2661_44458# a_4743_44484# 0.006148f
C32710 a_n967_45348# a_n984_44318# 0.00756f
C32711 a_n1059_45260# a_453_43940# 2.04e-20
C32712 a_n2293_45010# a_895_43940# 0.283316f
C32713 a_n2661_45010# a_2889_44172# 1.48e-20
C32714 a_n357_42282# a_6197_43396# 6.51e-20
C32715 SMPL_ON_P a_n3690_37440# 1.8e-19
C32716 a_n443_42852# a_1891_43646# 1.53e-19
C32717 a_n1177_44458# a_n452_44636# 0.011059f
C32718 a_11691_44458# a_13720_44458# 0.029855f
C32719 a_13259_45724# a_14205_43396# 1.43e-20
C32720 a_13661_43548# a_4958_30871# 9.87e-21
C32721 a_15227_44166# a_15597_42852# 0.007489f
C32722 a_n913_45002# a_1414_42308# 0.021774f
C32723 a_n2312_39304# a_n4064_39616# 2.53e-19
C32724 a_n2312_40392# a_n2302_39866# 8.29e-19
C32725 a_7227_47204# a_3357_43084# 5.7e-19
C32726 a_n743_46660# a_9049_44484# 4.38e-19
C32727 a_11415_45002# a_15682_46116# 1.66e-19
C32728 a_3147_46376# a_5164_46348# 1.45e-21
C32729 a_3483_46348# a_5068_46348# 4.35e-20
C32730 a_n2109_47186# a_4927_45028# 0.00143f
C32731 a_21188_46660# a_10809_44734# 0.010814f
C32732 a_12816_46660# a_12839_46116# 1.51e-19
C32733 a_9067_47204# a_2437_43646# 0.006126f
C32734 a_18597_46090# a_18691_45572# 5.99e-19
C32735 a_n2661_46634# a_11652_45724# 1.97e-19
C32736 a_n2497_47436# a_3232_43370# 0.04813f
C32737 a_4185_45028# a_4419_46090# 0.066314f
C32738 a_1209_47178# a_413_45260# 3.61e-20
C32739 a_n443_46116# a_n2661_45010# 0.005128f
C32740 a_n1151_42308# a_n745_45366# 0.004257f
C32741 a_12741_44636# a_15015_46420# 1.62e-21
C32742 a_n971_45724# a_3065_45002# 0.220337f
C32743 a_16327_47482# a_19418_45938# 1.07e-19
C32744 a_18479_47436# a_19256_45572# 2.31e-22
C32745 a_15567_42826# a_15959_42545# 8.04e-19
C32746 a_5342_30871# a_15890_42674# 0.001531f
C32747 a_17538_32519# C3_N_btm 2.76e-20
C32748 a_14401_32519# C5_N_btm 0.001006f
C32749 a_n4318_38680# a_n4064_40160# 0.079598f
C32750 a_16414_43172# a_15803_42450# 1.98e-19
C32751 a_n2661_43922# a_n1331_43914# 0.002577f
C32752 a_6109_44484# a_5663_43940# 1.88e-19
C32753 a_n2293_43922# a_n1899_43946# 0.013114f
C32754 a_n2661_42834# a_n1549_44318# 0.011433f
C32755 a_8975_43940# a_10729_43914# 2.43e-19
C32756 a_10057_43914# a_10949_43914# 5.37e-19
C32757 a_11823_42460# a_12895_43230# 0.0142f
C32758 a_n357_42282# a_10752_42852# 1.14e-19
C32759 a_13259_45724# a_22400_42852# 0.34531f
C32760 a_3537_45260# a_7221_43396# 9.66e-20
C32761 a_n2661_46634# DATA[0] 0.012107f
C32762 a_n913_45002# a_12281_43396# 0.28203f
C32763 a_n1059_45260# a_8873_43396# 6.35e-19
C32764 a_n2293_42834# a_n2129_43609# 0.017516f
C32765 a_11967_42832# a_20159_44458# 0.056889f
C32766 a_19006_44850# a_20362_44736# 3.32e-21
C32767 a_8191_45002# a_8147_43396# 1.42e-20
C32768 a_526_44458# a_5379_42460# 1.71e-19
C32769 a_10903_43370# a_13333_42558# 0.00168f
C32770 a_n2312_38680# VDD 0.540248f
C32771 a_4185_45028# a_4958_30871# 0.121495f
C32772 a_626_44172# a_n1557_42282# 0.003837f
C32773 a_18479_45785# a_19095_43396# 0.001675f
C32774 a_3090_45724# a_n1059_45260# 0.008195f
C32775 a_6945_45028# a_2711_45572# 0.036364f
C32776 a_8199_44636# a_11652_45724# 4.91e-19
C32777 a_11133_46155# a_7499_43078# 1.49e-20
C32778 a_9625_46129# a_10490_45724# 1.99e-19
C32779 a_6969_46634# a_6171_45002# 1.08e-20
C32780 a_4791_45118# a_9241_44734# 6.15e-20
C32781 a_11415_45002# a_16680_45572# 0.003026f
C32782 a_19123_46287# a_18691_45572# 0.009086f
C32783 a_4883_46098# a_5883_43914# 0.01188f
C32784 a_10227_46804# a_16112_44458# 0.001281f
C32785 a_3877_44458# a_2304_45348# 6.26e-21
C32786 a_n133_46660# a_n2661_43370# 2.93e-22
C32787 a_19321_45002# a_17719_45144# 1.57e-20
C32788 a_13661_43548# a_18911_45144# 0.03394f
C32789 a_9863_46634# a_8953_45002# 3.37e-20
C32790 a_5807_45002# a_19778_44110# 0.032504f
C32791 a_12549_44172# a_11691_44458# 0.025825f
C32792 a_584_46384# a_n2661_42834# 0.079307f
C32793 a_12741_44636# a_16333_45814# 1.84e-20
C32794 a_9290_44172# a_10053_45546# 8.06e-21
C32795 a_9823_46155# a_10193_42453# 0.001684f
C32796 a_16327_47482# a_18248_44752# 0.050926f
C32797 a_15803_42450# a_7174_31319# 9.34e-20
C32798 a_16269_42308# a_4958_30871# 0.001757f
C32799 a_5934_30871# a_1343_38525# 1.69e-19
C32800 a_16414_43172# VDD 0.201389f
C32801 a_3422_30871# a_3080_42308# 0.022126f
C32802 a_1307_43914# a_5193_42852# 2.47e-20
C32803 a_14815_43914# a_9145_43396# 2.41e-19
C32804 a_n2956_38216# a_n3690_38304# 0.016795f
C32805 a_9823_46155# VDD 0.102474f
C32806 a_17767_44458# a_16823_43084# 7.97e-22
C32807 a_12429_44172# a_12710_44260# 0.008628f
C32808 a_n2065_43946# a_n2012_43396# 8.21e-20
C32809 a_n809_44244# a_n1177_43370# 0.002467f
C32810 a_n1549_44318# a_n1352_43396# 2.22e-19
C32811 a_10193_42453# a_7174_31319# 0.020527f
C32812 a_n2810_45572# a_n4064_37984# 0.094405f
C32813 a_n2017_45002# a_n4318_38216# 7.46e-19
C32814 a_15493_43396# a_15493_43940# 0.188034f
C32815 a_19862_44208# a_11341_43940# 0.07932f
C32816 a_14539_43914# a_17678_43396# 1.74e-19
C32817 a_2711_45572# a_14127_45572# 0.001525f
C32818 a_16388_46812# a_18443_44721# 2.06e-20
C32819 a_20692_30879# a_22959_45572# 4.31e-19
C32820 a_2324_44458# a_7418_45394# 0.00182f
C32821 a_584_46384# a_n1352_43396# 1.26e-20
C32822 a_n971_45724# a_458_43396# 1.17e-19
C32823 a_n2956_39768# a_n4318_39768# 0.023595f
C32824 a_10193_42453# a_10306_45572# 0.002653f
C32825 a_8746_45002# a_10216_45572# 0.001575f
C32826 a_n2293_46634# a_6453_43914# 6.32e-20
C32827 a_768_44030# a_8018_44260# 9.58e-19
C32828 a_20205_31679# a_20447_31679# 9.01329f
C32829 a_11387_46155# a_n2661_43370# 2.17e-21
C32830 a_n4064_39616# C8_P_btm 0.001799f
C32831 a_n3420_39616# C6_P_btm 5.51e-20
C32832 a_11599_46634# a_13661_43548# 0.078449f
C32833 a_14955_47212# a_13747_46662# 3.09e-21
C32834 a_15507_47210# a_5807_45002# 0.002062f
C32835 a_1431_47204# a_n2661_46098# 1.15e-19
C32836 a_584_46384# a_645_46660# 3.21e-21
C32837 a_7754_39964# a_8530_39574# 9.77e-19
C32838 a_7174_31319# VDD 0.669838f
C32839 a_18479_47436# a_12549_44172# 0.015281f
C32840 a_16327_47482# a_16285_47570# 0.001903f
C32841 a_16241_47178# a_16697_47582# 4.2e-19
C32842 a_4883_46098# a_n881_46662# 0.193691f
C32843 a_20712_42282# RST_Z 4.07e-20
C32844 a_n443_46116# a_171_46873# 0.029327f
C32845 a_n1151_42308# a_1983_46706# 4.68e-20
C32846 a_6545_47178# a_n1925_46634# 0.02342f
C32847 VDAC_Pi a_7754_38470# 0.008396f
C32848 a_7754_39632# a_3754_38470# 0.002634f
C32849 a_4958_30871# VREF_GND 0.054206f
C32850 a_9067_47204# a_n2661_46634# 1.36e-19
C32851 a_n237_47217# a_3524_46660# 1.32e-21
C32852 a_n2109_47186# a_3877_44458# 0.021838f
C32853 a_15811_47375# a_16131_47204# 0.002108f
C32854 a_10227_46804# a_15928_47570# 0.025137f
C32855 a_2982_43646# a_8791_43396# 1.3e-21
C32856 a_14021_43940# a_19095_43396# 1.04e-19
C32857 a_n356_44636# a_1755_42282# 0.00959f
C32858 a_11967_42832# a_11301_43218# 8.99e-21
C32859 a_10306_45572# VDD 4.3e-19
C32860 a_5883_43914# a_7963_42308# 1.91e-21
C32861 a_5343_44458# a_8337_42558# 9.56e-19
C32862 a_n97_42460# a_14358_43442# 1.05e-20
C32863 a_12549_44172# a_4190_30871# 0.270972f
C32864 a_5263_45724# a_5343_44458# 1.81e-20
C32865 a_2711_45572# a_8103_44636# 5.76e-21
C32866 a_n443_42852# a_13720_44458# 1.6e-20
C32867 a_19692_46634# a_19319_43548# 5.04e-20
C32868 a_11823_42460# a_11827_44484# 0.024482f
C32869 a_11525_45546# a_11691_44458# 4.12e-20
C32870 a_10193_42453# a_16981_45144# 0.001232f
C32871 a_n967_45348# a_n467_45028# 0.005391f
C32872 a_20202_43084# a_20365_43914# 2.68e-21
C32873 a_n2312_40392# a_n3674_39304# 0.025635f
C32874 a_5257_43370# a_6031_43396# 0.004037f
C32875 a_8199_44636# a_7845_44172# 7.26e-19
C32876 a_5937_45572# a_7542_44172# 2.83e-19
C32877 a_12741_44636# a_15493_43396# 1.11e-19
C32878 a_n2017_45002# a_2382_45260# 0.032443f
C32879 a_3357_43084# a_6171_45002# 0.003278f
C32880 a_n863_45724# a_7_44811# 7.59e-19
C32881 a_n1099_45572# a_n356_44636# 5.17e-21
C32882 a_584_46384# a_n2293_42282# 8.38e-19
C32883 a_22959_47212# a_22959_46660# 0.025171f
C32884 VREF_GND VCM 2.79113f
C32885 a_3877_44458# a_5841_46660# 9.39e-19
C32886 a_4646_46812# a_6999_46987# 4.77e-19
C32887 a_768_44030# a_765_45546# 0.033731f
C32888 a_11453_44696# a_21076_30879# 8.96e-19
C32889 a_9067_47204# a_8199_44636# 6.76e-22
C32890 a_6575_47204# a_5937_45572# 1.83e-20
C32891 a_5807_45002# a_15227_46910# 1.37e-19
C32892 a_12549_44172# a_17829_46910# 0.057751f
C32893 a_n1151_42308# a_14275_46494# 0.003302f
C32894 a_4817_46660# a_6755_46942# 5.52e-20
C32895 a_5257_43370# a_7715_46873# 1.05e-20
C32896 a_n2497_47436# a_n1379_46482# 5.68e-19
C32897 a_n4318_39304# a_n3674_38680# 0.031218f
C32898 a_13483_43940# a_13657_42558# 8.24e-21
C32899 a_16137_43396# a_16414_43172# 0.179708f
C32900 a_743_42282# a_3935_42891# 1.46e-20
C32901 a_18114_32519# C4_N_btm 1.47e-19
C32902 a_19721_31679# C3_N_btm 0.001023f
C32903 a_n1991_42858# a_n1641_43230# 0.229804f
C32904 a_n2157_42858# a_n1076_43230# 0.102325f
C32905 a_n1853_43023# a_n901_43156# 0.081949f
C32906 a_10341_43396# a_22165_42308# 3.24e-19
C32907 a_16547_43609# a_5342_30871# 1.72e-20
C32908 a_n2840_42826# a_n3674_39304# 0.16082f
C32909 a_n1613_43370# a_5934_30871# 9.62e-19
C32910 a_5205_44484# a_5205_44734# 0.015405f
C32911 a_526_44458# a_7287_43370# 5.68e-19
C32912 a_5111_44636# a_5891_43370# 0.702087f
C32913 a_7499_43078# a_12429_44172# 0.001488f
C32914 a_20107_45572# a_20362_44736# 1.08e-21
C32915 a_20273_45572# a_20159_44458# 1.49e-21
C32916 a_12465_44636# a_14456_42282# 1.36e-21
C32917 a_10809_44734# a_8685_43396# 1.08e-21
C32918 a_2324_44458# a_10341_43396# 3.06e-19
C32919 a_1423_45028# a_8975_43940# 0.331942f
C32920 a_18587_45118# a_18911_45144# 0.010993f
C32921 en_comp a_n2293_43922# 0.412872f
C32922 a_n967_45348# a_n2661_43922# 0.024232f
C32923 a_n2312_40392# a_5742_30871# 9.24e-21
C32924 a_20623_45572# a_11967_42832# 7.43e-21
C32925 a_2437_43646# a_17517_44484# 3.17e-20
C32926 a_9290_44172# a_13837_43396# 0.002072f
C32927 a_10193_42453# a_10729_43914# 0.010339f
C32928 a_8746_45002# a_10405_44172# 1.94e-20
C32929 a_n1059_45260# a_14815_43914# 2.69e-20
C32930 a_3232_43370# a_6109_44484# 0.072011f
C32931 a_1307_43914# a_16112_44458# 0.012033f
C32932 a_15227_44166# a_18083_42858# 2.37e-19
C32933 a_21076_30879# a_17364_32525# 0.057544f
C32934 w_1575_34946# a_3754_38470# 6.84e-19
C32935 a_n2442_46660# a_n2810_45572# 0.045104f
C32936 a_n2472_46634# a_n2661_45546# 0.001532f
C32937 a_14976_45028# a_13759_46122# 1.44e-20
C32938 a_3090_45724# a_13925_46122# 1.1e-19
C32939 a_12549_44172# a_n443_42852# 0.069091f
C32940 a_n2956_39768# a_n2956_38216# 0.043382f
C32941 a_20885_46660# a_20202_43084# 2.46e-21
C32942 a_10227_46804# a_11962_45724# 4.98e-21
C32943 a_765_45546# a_1176_45822# 0.241847f
C32944 a_13059_46348# a_3483_46348# 0.319214f
C32945 a_2063_45854# a_8696_44636# 0.029184f
C32946 a_18525_43370# a_18214_42558# 8.42e-21
C32947 a_15743_43084# a_18907_42674# 1.64e-20
C32948 a_743_42282# a_15890_42674# 0.010042f
C32949 a_10729_43914# VDD 0.681371f
C32950 a_4361_42308# a_15051_42282# 0.016131f
C32951 a_16137_43396# a_7174_31319# 2.14e-20
C32952 a_5755_42852# a_4921_42308# 0.002018f
C32953 a_5534_30871# a_n1630_35242# 0.033914f
C32954 a_n443_42852# a_5111_42852# 0.005368f
C32955 a_19787_47423# VDD 0.256911f
C32956 a_13259_45724# a_22223_42860# 0.007322f
C32957 en_comp a_n97_42460# 5.85e-20
C32958 a_18989_43940# a_20159_44458# 1.23e-19
C32959 a_18287_44626# a_20679_44626# 5.48e-21
C32960 a_9159_44484# a_n2661_43922# 0.004106f
C32961 a_n1177_44458# a_n809_44244# 0.00369f
C32962 a_n1352_44484# a_n1549_44318# 3.11e-20
C32963 a_18597_46090# START 0.020125f
C32964 a_1823_45246# a_3905_42558# 0.010516f
C32965 a_19386_47436# RST_Z 6.35e-20
C32966 a_n2293_45010# a_458_43396# 1.65e-19
C32967 a_n2661_45010# a_1049_43396# 1.29e-21
C32968 a_n2017_45002# a_n1655_43396# 4.3e-19
C32969 a_n2661_44458# a_1414_42308# 6.41e-20
C32970 a_8953_45002# a_9801_43940# 4.55e-20
C32971 a_8696_44636# a_14955_43396# 2.57e-23
C32972 a_1307_43914# a_1443_43940# 0.042476f
C32973 a_n357_42282# a_10922_42852# 0.006403f
C32974 a_10227_46804# a_13807_45067# 4.48e-20
C32975 a_11599_46634# a_18587_45118# 4.52e-20
C32976 a_15682_46116# a_13259_45724# 0.002706f
C32977 a_n237_47217# a_5343_44458# 0.001668f
C32978 a_1176_45822# a_509_45822# 1.26e-19
C32979 a_584_46384# a_n1352_44484# 7.22e-22
C32980 a_765_45546# a_11652_45724# 2.49e-20
C32981 a_5807_45002# a_9482_43914# 0.018229f
C32982 a_13661_43548# a_13348_45260# 1.86e-19
C32983 a_3483_46348# a_3218_45724# 1.76e-19
C32984 a_3147_46376# a_3316_45546# 0.012262f
C32985 a_13059_46348# a_14495_45572# 0.004072f
C32986 a_3090_45724# a_15599_45572# 0.022054f
C32987 a_14976_45028# a_15297_45822# 2.87e-19
C32988 a_16327_47482# a_16922_45042# 0.060018f
C32989 a_12861_44030# a_18494_42460# 0.021479f
C32990 a_n1151_42308# a_n2433_44484# 1.87e-19
C32991 a_5937_45572# a_n2661_45546# 1.02e-19
C32992 a_n2293_46634# a_6171_45002# 2.7e-21
C32993 a_n743_46660# a_5147_45002# 9.05e-20
C32994 a_13925_46122# a_15002_46116# 1.46e-19
C32995 a_17364_32525# C0_N_btm 8.17e-21
C32996 a_13678_32519# C7_N_btm 2.68e-20
C32997 a_n784_42308# a_7174_31319# 1.93626f
C32998 a_n3674_38680# a_n4334_40480# 1.51e-19
C32999 a_8791_42308# a_5742_30871# 4.57e-20
C33000 a_13887_32519# C4_N_btm 0.001746f
C33001 a_21487_43396# VDD 0.222231f
C33002 a_1423_45028# a_2905_42968# 6.76e-22
C33003 a_11827_44484# a_18429_43548# 4.78e-21
C33004 a_18494_42460# a_19700_43370# 3.28e-20
C33005 a_n2293_42834# a_n2840_42826# 9.62e-19
C33006 a_5883_43914# a_8685_43396# 3.79e-19
C33007 a_21076_30879# a_21589_35634# 5.95e-20
C33008 a_20107_46660# VDD 0.442554f
C33009 a_19123_46287# START 0.003458f
C33010 a_7845_44172# a_8018_44260# 0.007688f
C33011 a_7542_44172# a_8333_44056# 7.67e-20
C33012 a_n357_42282# a_17531_42308# 4.24e-20
C33013 a_n913_45002# a_873_42968# 7.48e-19
C33014 a_3422_30871# a_14021_43940# 0.018792f
C33015 a_11691_44458# a_16977_43638# 3.52e-19
C33016 a_16237_45028# a_16547_43609# 3.95e-21
C33017 a_n2661_42834# a_n1177_43370# 8.78e-19
C33018 a_n2661_43922# a_n1917_43396# 1.76e-20
C33019 a_765_45546# DATA[0] 6.38e-19
C33020 a_2711_45572# a_6812_45938# 0.003338f
C33021 a_4646_46812# a_7640_43914# 0.183308f
C33022 a_n2293_46634# a_14673_44172# 0.100552f
C33023 a_19321_45002# a_18588_44850# 1.03e-20
C33024 a_13259_45724# a_16680_45572# 0.038605f
C33025 a_13747_46662# a_11967_42832# 0.021948f
C33026 a_13661_43548# a_19615_44636# 1.88e-21
C33027 a_3483_46348# a_13556_45296# 0.375978f
C33028 a_8270_45546# a_5343_44458# 1.28e-19
C33029 a_9625_46129# a_6171_45002# 4.78e-21
C33030 a_15227_44166# a_18450_45144# 0.002515f
C33031 a_8049_45260# a_18691_45572# 0.006525f
C33032 a_9290_44172# a_5111_44636# 0.031975f
C33033 a_5937_45572# a_5205_44484# 0.481405f
C33034 a_15015_46420# a_413_45260# 5.92e-21
C33035 a_7920_46348# a_7705_45326# 1.67e-19
C33036 a_16375_45002# a_16333_45814# 0.001746f
C33037 a_1138_42852# a_1307_43914# 0.123153f
C33038 a_12861_44030# a_15673_47210# 5.52e-20
C33039 a_n4209_38502# a_n4251_38528# 0.00226f
C33040 a_n2946_38778# a_n2302_38778# 6.68e-19
C33041 a_n3420_38528# a_n2860_38778# 0.002301f
C33042 a_5932_42308# VDD 0.534416f
C33043 a_5934_30871# C5_N_btm 0.139996f
C33044 a_n815_47178# a_n1613_43370# 2.12e-19
C33045 a_n971_45724# a_3094_47243# 2.1e-19
C33046 a_584_46384# a_2487_47570# 0.005904f
C33047 a_1209_47178# a_3094_47570# 7.14e-20
C33048 a_6123_31319# C7_N_btm 0.005631f
C33049 a_14955_47212# a_11599_46634# 0.011007f
C33050 a_n443_46116# a_4883_46098# 0.037308f
C33051 a_13717_47436# a_16241_47178# 6.54e-20
C33052 a_17531_42308# CAL_N 7.31e-19
C33053 a_5742_30871# C9_P_btm 0.003249f
C33054 a_14311_47204# a_15507_47210# 8.1e-22
C33055 a_1736_39587# VDAC_Pi 0.009393f
C33056 a_3905_42865# a_4361_42308# 3.2e-19
C33057 a_n1899_43946# a_n901_43156# 0.001167f
C33058 a_n984_44318# a_n1853_43023# 1.28e-20
C33059 a_n1331_43914# a_n1641_43230# 1.38e-21
C33060 a_n1761_44111# a_n1076_43230# 2.91e-19
C33061 a_19862_44208# a_10341_43396# 0.028065f
C33062 a_2307_45899# VDD 7.28e-19
C33063 a_5891_43370# a_5837_43172# 4.79e-20
C33064 a_n1177_43370# a_n1352_43396# 0.233657f
C33065 a_n2129_43609# a_n2012_43396# 0.183186f
C33066 a_n2433_43396# a_n1809_43762# 9.73e-19
C33067 a_n4318_39304# a_n1190_43762# 3.5e-21
C33068 a_n2956_37592# a_n2946_39866# 3.12e-19
C33069 a_11967_42832# a_10796_42968# 0.001301f
C33070 a_n2438_43548# a_1756_43548# 2.24e-20
C33071 a_14495_45572# a_13556_45296# 1.1e-20
C33072 a_13249_42308# a_13777_45326# 2.35e-21
C33073 a_n357_42282# a_18184_42460# 0.106442f
C33074 a_n1613_43370# a_7221_43396# 2.95e-19
C33075 a_9159_45572# a_6171_45002# 0.00193f
C33076 a_16327_47482# a_15743_43084# 1.21037f
C33077 a_n971_45724# a_n967_43230# 4.78e-20
C33078 a_526_44458# a_n23_44458# 3.73e-19
C33079 a_n1925_42282# a_n356_44636# 0.020589f
C33080 a_10210_45822# a_8953_45002# 1.45e-19
C33081 a_21076_30879# a_19237_31679# 0.05495f
C33082 a_20273_45572# a_20623_45572# 0.219856f
C33083 a_20107_45572# a_21363_45546# 0.043567f
C33084 a_n2497_47436# a_2905_42968# 7.38e-22
C33085 a_3090_45724# a_18326_43940# 5.94e-19
C33086 a_n2442_46660# a_n1557_42282# 2.36e-20
C33087 a_15143_45578# a_9482_43914# 7.52e-21
C33088 a_13904_45546# a_14180_45002# 1.92e-19
C33089 a_6755_46942# a_15037_44260# 2.99e-20
C33090 a_5807_45002# a_7715_46873# 0.029268f
C33091 a_n2497_47436# a_n1076_46494# 0.001159f
C33092 a_12891_46348# a_10249_46116# 6.35e-21
C33093 a_11309_47204# a_6755_46942# 0.09972f
C33094 a_13717_47436# a_16721_46634# 6.05e-22
C33095 a_12861_44030# a_16388_46812# 0.11634f
C33096 a_13487_47204# a_13059_46348# 7.45e-20
C33097 a_12465_44636# a_15559_46634# 4.15e-21
C33098 C9_P_btm C0_dummy_P_btm 0.11363f
C33099 C6_P_btm C2_P_btm 0.138423f
C33100 C7_P_btm C1_P_btm 0.129707f
C33101 C8_P_btm C0_P_btm 0.148433f
C33102 C5_P_btm C3_P_btm 0.136119f
C33103 a_n2661_46634# a_5167_46660# 0.007924f
C33104 EN_VIN_BSTR_N C4_N_btm 0.116925f
C33105 a_n1741_47186# a_n1991_46122# 1.1e-19
C33106 SMPL_ON_P a_n1853_46287# 8.1e-21
C33107 a_9067_47204# a_765_45546# 0.007492f
C33108 a_4883_46098# a_17609_46634# 3.14e-20
C33109 a_20894_47436# a_19692_46634# 4.29e-20
C33110 a_22459_39145# VIN_N 2.29e-20
C33111 a_2107_46812# a_2959_46660# 0.003474f
C33112 a_33_46660# a_1057_46660# 2.36e-20
C33113 a_n1925_46634# a_3877_44458# 0.070082f
C33114 a_13507_46334# a_15227_44166# 0.235687f
C33115 a_15811_47375# a_14513_46634# 9.55e-20
C33116 C10_P_btm C0_dummy_N_btm 0.001369f
C33117 a_n881_46662# a_6682_46660# 3.35e-19
C33118 a_n815_47178# a_n2293_46098# 5.23e-38
C33119 a_22717_36887# VDD 1.72e-20
C33120 a_5663_43940# a_6171_42473# 3.37e-21
C33121 a_3422_30871# a_15764_42576# 7.68e-20
C33122 a_18184_42460# CAL_N 7.63e-19
C33123 a_3626_43646# a_12545_42858# 8.41e-20
C33124 a_2982_43646# a_12895_43230# 2.86e-20
C33125 a_3457_43396# a_3681_42891# 0.001119f
C33126 a_8147_43396# a_7765_42852# 7.06e-19
C33127 a_8791_43396# a_7871_42858# 1.26e-19
C33128 a_11967_42832# a_4958_30871# 0.239255f
C33129 a_16547_43609# a_743_42282# 1.93e-20
C33130 a_18525_43370# a_16823_43084# 0.009621f
C33131 a_1423_45028# VDD 4.06861f
C33132 a_n1177_43370# a_n2293_42282# 2.19e-22
C33133 a_8696_44636# a_n2661_42834# 0.004739f
C33134 a_n863_45724# a_n2661_42282# 1.84e-19
C33135 a_6171_45002# a_16237_45028# 0.05704f
C33136 a_n467_45028# a_n1917_44484# 1.34e-20
C33137 a_n1059_45260# a_4743_44484# 6.94e-22
C33138 a_n2017_45002# a_5343_44458# 0.027073f
C33139 a_4791_45118# a_5934_30871# 2.81e-20
C33140 a_n357_42282# a_2537_44260# 2.9e-20
C33141 a_n913_45002# a_n699_43396# 2.01e-19
C33142 a_16375_45002# a_15493_43396# 1.46e-20
C33143 a_17339_46660# a_17499_43370# 1.36e-19
C33144 a_327_44734# a_n2433_44484# 1.63e-21
C33145 a_1667_45002# a_n2661_44458# 1.72e-20
C33146 a_n443_42852# a_7542_44172# 1.35e-21
C33147 a_2324_44458# a_n97_42460# 5.01e-20
C33148 a_n443_46116# a_1260_45572# 0.004853f
C33149 a_7577_46660# a_3483_46348# 7.22e-22
C33150 a_9804_47204# a_10044_46482# 9.19e-19
C33151 a_15227_44166# a_20623_46660# 0.008959f
C33152 a_14513_46634# a_13059_46348# 0.006934f
C33153 a_14180_46812# a_16388_46812# 1.67e-20
C33154 a_n1925_46634# a_n1736_46482# 0.002936f
C33155 a_11309_47204# a_8049_45260# 5.06e-19
C33156 a_5257_43370# a_4419_46090# 8.58e-19
C33157 a_11735_46660# a_11415_45002# 9.22e-21
C33158 a_14976_45028# a_16434_46660# 5.98e-20
C33159 a_4883_46098# a_19443_46116# 0.002033f
C33160 a_13507_46334# a_21071_46482# 7.31e-19
C33161 a_19466_46812# a_20273_46660# 7.76e-20
C33162 a_19692_46634# a_20411_46873# 0.215749f
C33163 a_3815_47204# a_4099_45572# 1.36e-21
C33164 a_n1151_42308# a_6194_45824# 4.58e-20
C33165 a_2063_45854# a_7227_45028# 0.021063f
C33166 a_10695_43548# a_5742_30871# 3.57e-19
C33167 a_3080_42308# a_7174_31319# 0.22305f
C33168 a_21398_44850# VDD 0.077608f
C33169 a_17730_32519# C2_N_btm 4.56e-20
C33170 a_3626_43646# a_19332_42282# 0.013212f
C33171 a_4190_30871# a_n1630_35242# 0.039258f
C33172 a_743_42282# a_n3674_37592# 2.16e-19
C33173 a_10341_43396# a_9803_42558# 6.46e-20
C33174 a_13678_32519# COMP_P 2.06e-19
C33175 a_19237_31679# C0_N_btm 0.040442f
C33176 a_8701_44490# a_8855_44734# 0.008678f
C33177 a_18911_45144# a_11967_42832# 5.48e-20
C33178 a_16922_45042# a_20835_44721# 2.59e-21
C33179 a_3232_43370# a_10405_44172# 2.4e-20
C33180 a_7499_43078# a_6643_43396# 1.32e-19
C33181 a_20202_43084# a_22400_42852# 3.36e-20
C33182 a_6298_44484# a_9313_44734# 7.5e-22
C33183 a_10334_44484# a_5891_43370# 7.17e-19
C33184 a_n1917_44484# a_n2661_43922# 0.010578f
C33185 a_n1177_44458# a_n2661_42834# 0.002427f
C33186 a_n2293_42834# a_n2472_43914# 4.12e-19
C33187 a_11691_44458# a_17061_44734# 0.001749f
C33188 a_20205_31679# a_13467_32519# 0.051513f
C33189 a_5111_44636# a_10807_43548# 1.74e-20
C33190 a_11827_44484# a_15367_44484# 6.14e-19
C33191 a_1423_45028# a_5495_43940# 1.89e-20
C33192 a_n2497_47436# VDD 1.33346f
C33193 a_17583_46090# a_17715_44484# 0.22771f
C33194 SMPL_ON_P a_n2661_43370# 0.002305f
C33195 a_15559_46634# a_2711_45572# 2.74e-20
C33196 a_3090_45724# a_5263_45724# 1.96e-19
C33197 a_13747_46662# a_20273_45572# 0.002644f
C33198 a_12549_44172# a_2437_43646# 0.004577f
C33199 a_13059_46348# a_n357_42282# 1.98e-19
C33200 a_n1613_43370# a_n2661_45010# 0.223356f
C33201 a_4883_46098# a_3537_45260# 2.75e-19
C33202 a_3147_46376# a_5066_45546# 5.42e-21
C33203 a_11599_46634# a_13159_45002# 6.88e-21
C33204 a_12861_44030# a_13777_45326# 0.00239f
C33205 a_n784_42308# a_5932_42308# 0.151611f
C33206 a_1755_42282# a_3823_42558# 2.57e-19
C33207 a_1606_42308# a_5267_42460# 1.69e-20
C33208 COMP_P a_6123_31319# 0.02889f
C33209 a_2351_42308# a_2903_42308# 8.7e-20
C33210 a_n443_42852# a_n1630_35242# 6.01e-19
C33211 a_n913_45002# a_n4318_38680# 4.18e-21
C33212 a_n1059_45260# a_n1736_43218# 5.17e-20
C33213 a_n1352_44484# a_n1177_43370# 8.8e-22
C33214 a_n1177_44458# a_n1352_43396# 7.26e-20
C33215 a_6682_46987# VDD 6.34e-20
C33216 a_3537_45260# a_5649_42852# 0.048691f
C33217 a_n2017_45002# a_n1545_43230# 6.01e-19
C33218 a_3357_43084# a_3681_42891# 0.052403f
C33219 en_comp a_n901_43156# 4.8e-21
C33220 a_n967_45348# a_n1641_43230# 0.00611f
C33221 a_n357_42282# a_2903_42308# 2.49e-20
C33222 a_n755_45592# a_2713_42308# 0.243663f
C33223 a_11823_42460# a_13569_43230# 7.84e-20
C33224 a_9313_44734# a_10555_44260# 0.005264f
C33225 a_n467_45028# a_n1853_43023# 5.11e-21
C33226 a_n2065_43946# a_644_44056# 6.01e-22
C33227 a_n1899_43946# a_n984_44318# 0.118759f
C33228 a_n755_45592# a_2957_45546# 0.044162f
C33229 a_19321_45002# a_18443_44721# 6.29e-21
C33230 a_n2661_45546# a_n443_42852# 0.141363f
C33231 a_18189_46348# a_16680_45572# 6.45e-21
C33232 a_13747_46662# a_18989_43940# 0.002177f
C33233 a_17583_46090# a_15861_45028# 1.62e-19
C33234 a_17715_44484# a_8696_44636# 0.017149f
C33235 a_12861_44030# a_20640_44752# 0.001266f
C33236 a_380_45546# a_n356_45724# 0.088749f
C33237 a_n2956_38216# a_n906_45572# 1.15e-19
C33238 a_8049_45260# a_10490_45724# 0.006151f
C33239 a_10586_45546# a_7499_43078# 1.07e-19
C33240 a_10809_44734# a_11778_45572# 2.41e-19
C33241 a_14035_46660# a_14180_45002# 3.28e-19
C33242 a_12594_46348# a_14033_45572# 9.76e-19
C33243 a_8270_45546# a_8560_45348# 4.84e-20
C33244 a_8128_46384# a_8375_44464# 3.74e-20
C33245 a_11599_46634# a_11967_42832# 1.61e-22
C33246 a_1208_46090# a_2437_43646# 6.09e-20
C33247 a_n2293_46098# a_n2661_45010# 1.61e-19
C33248 COMP_P EN_VIN_BSTR_P 6.4e-19
C33249 a_n971_45724# a_4007_47204# 0.01992f
C33250 a_n785_47204# a_n1151_42308# 0.07743f
C33251 a_2124_47436# a_2063_45854# 0.074695f
C33252 a_n237_47217# a_3785_47178# 1.77e-21
C33253 a_n1741_47186# a_5129_47502# 0.012935f
C33254 a_1209_47178# a_2905_45572# 1.33e-19
C33255 a_n2109_47186# a_6151_47436# 9.88e-20
C33256 a_n4064_40160# a_n2302_39866# 2.59e-20
C33257 a_n4209_39590# a_n3690_39616# 0.045251f
C33258 a_n2302_40160# a_n4064_39616# 2.59e-20
C33259 a_n4334_39616# a_n3565_39590# 2e-19
C33260 a_3232_43370# a_6171_42473# 5.89e-23
C33261 a_n913_45002# a_11551_42558# 3.95e-19
C33262 a_14673_44172# a_743_42282# 6.85e-21
C33263 a_n2293_43922# a_n2157_42858# 0.040551f
C33264 a_n2661_43922# a_n1853_43023# 1.11e-20
C33265 a_n2661_42834# a_n1991_42858# 8.85e-19
C33266 a_375_42282# a_n1630_35242# 0.036312f
C33267 a_20835_44721# a_15743_43084# 1.25e-21
C33268 a_n356_44636# a_8387_43230# 1.68e-20
C33269 a_3537_45260# a_7963_42308# 4.5e-20
C33270 en_comp a_10533_42308# 4.34e-21
C33271 a_8049_45260# START 1.99e-20
C33272 a_n2017_45002# a_12563_42308# 0.003288f
C33273 a_n443_42852# a_5205_44484# 6.5e-20
C33274 a_16680_45572# a_17478_45572# 0.001111f
C33275 a_8696_44636# a_15861_45028# 0.26484f
C33276 a_16115_45572# a_16223_45938# 0.057222f
C33277 a_n2293_46634# a_14761_44260# 0.009374f
C33278 a_4791_45118# a_7221_43396# 2.22e-20
C33279 a_12891_46348# a_13565_43940# 0.001515f
C33280 a_2324_44458# a_742_44458# 0.00317f
C33281 a_n2661_45546# a_375_42282# 0.001753f
C33282 a_2711_45572# a_3065_45002# 0.012727f
C33283 a_14033_45822# a_14127_45572# 1.26e-19
C33284 a_19692_46634# a_3422_30871# 0.208985f
C33285 a_17339_46660# a_18204_44850# 1.39e-19
C33286 a_n237_47217# a_3090_45724# 3.45e-19
C33287 a_2063_45854# a_11813_46116# 0.093948f
C33288 a_6545_47178# a_6999_46987# 3.51e-19
C33289 a_n881_46662# a_n133_46660# 0.005885f
C33290 CAL_N a_22459_39145# 0.014789f
C33291 a_22521_40599# a_22521_40055# 0.086402f
C33292 a_22469_40625# a_22780_40945# 4.21e-20
C33293 a_n4064_38528# VREF_GND 0.034351f
C33294 a_8128_46384# a_n1925_46634# 0.21095f
C33295 a_9313_45822# a_10150_46912# 3.39e-20
C33296 a_n1435_47204# a_8667_46634# 3.08e-20
C33297 a_6851_47204# a_6969_46634# 1.59e-19
C33298 a_7227_47204# a_6755_46942# 1.17e-19
C33299 a_11031_47542# a_10428_46928# 8.15e-19
C33300 a_n1613_43370# a_171_46873# 0.11335f
C33301 a_2266_47243# a_2107_46812# 2.19e-19
C33302 a_n3565_37414# EN_VIN_BSTR_P 0.069167f
C33303 a_4338_37500# CAL_P 0.00316f
C33304 a_5807_45002# a_13747_46662# 0.103485f
C33305 a_12549_44172# a_n2661_46634# 0.024531f
C33306 a_n4251_38304# VDD 3.95e-19
C33307 a_22591_45572# VDD 0.314172f
C33308 a_14021_43940# a_16414_43172# 9.19e-22
C33309 a_15493_43940# a_21356_42826# 1.97e-20
C33310 a_11341_43940# a_21671_42860# 6.71e-21
C33311 a_14579_43548# a_10341_43396# 0.029139f
C33312 a_10695_43548# a_10849_43646# 0.010303f
C33313 a_3357_43084# RST_Z 0.031959f
C33314 a_n2293_43922# a_9803_42558# 4.58e-20
C33315 a_n356_44636# a_16522_42674# 0.001524f
C33316 a_4093_43548# a_4361_42308# 1.72e-21
C33317 a_14205_43396# a_14955_43396# 0.157423f
C33318 a_9145_43396# a_12281_43396# 0.032945f
C33319 a_n2433_43396# a_n3674_39304# 9.78e-19
C33320 a_n1917_43396# a_n1641_43230# 0.00125f
C33321 a_n1352_43396# a_n1991_42858# 0.00171f
C33322 a_n1177_43370# a_n1423_42826# 0.0016f
C33323 a_n97_42460# a_n2157_42858# 9.01e-21
C33324 a_n4318_39304# a_n4318_38680# 0.059432f
C33325 a_20447_31679# C9_N_btm 3.26e-20
C33326 a_20205_31679# a_22315_44484# 2.01e-21
C33327 a_20107_45572# a_19778_44110# 1.5e-19
C33328 a_n2293_46634# a_3681_42891# 1.32e-20
C33329 a_768_44030# a_13460_43230# 6.38e-21
C33330 SMPL_ON_P COMP_P 0.03194f
C33331 a_13159_45002# a_13348_45260# 0.105274f
C33332 a_13017_45260# a_9482_43914# 0.048717f
C33333 a_3537_45260# a_3602_45348# 2.49e-19
C33334 a_n37_45144# a_117_45144# 0.008535f
C33335 a_19431_45546# a_11691_44458# 1.76e-20
C33336 a_5691_45260# a_1423_45028# 1.19e-19
C33337 a_7229_43940# a_1307_43914# 0.004598f
C33338 a_9049_44484# a_5891_43370# 1.84e-20
C33339 a_10903_43370# a_11816_44260# 8.18e-19
C33340 a_6755_46942# a_16547_43609# 7.51e-20
C33341 a_11453_44696# a_19335_46494# 6.23e-20
C33342 a_21496_47436# a_10809_44734# 0.0112f
C33343 a_13507_46334# a_22959_46124# 5.09e-19
C33344 a_n2293_46634# a_376_46348# 2.26e-21
C33345 a_n2661_46634# a_1208_46090# 8.96e-21
C33346 a_6755_46942# a_12156_46660# 0.013732f
C33347 a_10623_46897# a_10933_46660# 0.013793f
C33348 a_10554_47026# a_10861_46660# 3.69e-19
C33349 a_10249_46116# a_12359_47026# 1.42e-19
C33350 a_11735_46660# a_12251_46660# 0.105995f
C33351 a_8270_45546# a_3090_45724# 0.046518f
C33352 a_11813_46116# a_12469_46902# 2.33e-20
C33353 a_12465_44636# a_21137_46414# 5.25e-22
C33354 a_171_46873# a_n2293_46098# 0.001626f
C33355 a_13661_43548# a_4185_45028# 2.36e-21
C33356 a_n1925_46634# a_n1641_46494# 0.005997f
C33357 a_n2438_43548# a_n1853_46287# 0.001451f
C33358 a_n1151_42308# a_14371_46494# 2.26e-19
C33359 a_9804_47204# a_9823_46155# 0.063581f
C33360 a_5167_46660# a_765_45546# 0.003506f
C33361 a_21811_47423# a_6945_45028# 4.87e-19
C33362 a_4883_46098# a_22223_46124# 0.001059f
C33363 a_n97_42460# a_9803_42558# 0.099148f
C33364 a_3080_42308# a_5932_42308# 14.0282f
C33365 a_4905_42826# a_6171_42473# 2.44e-20
C33366 a_6109_44484# VDD 0.243629f
C33367 a_3422_30871# a_n4064_37440# 0.032121f
C33368 a_n1991_42858# a_n2293_42282# 9.15e-21
C33369 a_15681_43442# a_15597_42852# 1.25e-19
C33370 a_3626_43646# a_5379_42460# 0.057009f
C33371 a_16547_43609# a_16328_43172# 1.96e-19
C33372 a_14021_43940# a_7174_31319# 9.94e-21
C33373 a_10518_42984# a_10796_42968# 0.118759f
C33374 a_18911_45144# a_18989_43940# 0.016276f
C33375 a_11827_44484# a_14539_43914# 0.044058f
C33376 a_3357_43084# a_5663_43940# 0.015908f
C33377 a_4185_45028# a_10835_43094# 1.34e-20
C33378 a_4646_46812# a_5932_42308# 2.43e-19
C33379 a_12549_44172# a_19511_42282# 5.57e-20
C33380 a_10193_42453# a_18797_44260# 0.003033f
C33381 a_n357_42282# a_6293_42852# 0.00795f
C33382 a_n755_45592# a_6031_43396# 2.22e-20
C33383 a_n2017_45002# a_453_43940# 8.57e-22
C33384 a_n2661_45010# a_2675_43914# 1.7e-19
C33385 a_n2293_45010# a_2479_44172# 1.92e-20
C33386 a_15765_45572# a_15493_43940# 2.68e-20
C33387 SMPL_ON_P a_n3565_37414# 0.016441f
C33388 a_n443_42852# a_1427_43646# 0.002947f
C33389 a_n1177_44458# a_n1352_44484# 0.233657f
C33390 a_n2661_44458# a_n699_43396# 0.002525f
C33391 a_11691_44458# a_13076_44458# 0.03093f
C33392 a_14537_43396# a_16789_44484# 2.77e-19
C33393 a_13259_45724# a_14358_43442# 1.56e-20
C33394 a_n1059_45260# a_1414_42308# 0.031011f
C33395 a_n2312_39304# a_n2946_39866# 2.85e-20
C33396 a_n2312_40392# a_n4064_39616# 9.29e-20
C33397 a_6851_47204# a_3357_43084# 2.62e-19
C33398 a_n743_46660# a_7499_43078# 1.36e-19
C33399 a_11415_45002# a_2324_44458# 0.097878f
C33400 a_n2109_47186# a_5111_44636# 0.017519f
C33401 a_22000_46634# a_6945_45028# 2.76e-19
C33402 a_21363_46634# a_10809_44734# 0.012784f
C33403 a_12991_46634# a_12839_46116# 2.15e-19
C33404 a_6575_47204# a_2437_43646# 0.029543f
C33405 a_18597_46090# a_18909_45814# 8.56e-20
C33406 a_11599_46634# a_20273_45572# 0.004992f
C33407 a_n2293_46634# a_8746_45002# 3.85e-20
C33408 a_3483_46348# a_4704_46090# 2.61e-19
C33409 a_n1151_42308# a_n913_45002# 0.395136f
C33410 a_13747_46662# a_15143_45578# 0.040557f
C33411 a_n2661_46634# a_11525_45546# 0.003942f
C33412 a_5807_45002# a_6469_45572# 4.31e-19
C33413 a_12741_44636# a_14275_46494# 1.03e-20
C33414 a_n237_47217# a_2274_45254# 3.92e-19
C33415 a_n971_45724# a_2680_45002# 0.108251f
C33416 a_16327_47482# a_17668_45572# 0.003454f
C33417 a_18780_47178# a_18691_45572# 1.83e-20
C33418 a_15567_42826# a_15803_42450# 1.29e-20
C33419 a_5342_30871# a_15959_42545# 7.85e-19
C33420 a_17538_32519# C2_N_btm 2.28e-20
C33421 a_n3674_39304# a_n4064_40160# 0.024923f
C33422 a_n4318_38680# a_n4334_40480# 1.45e-19
C33423 a_17701_42308# a_14113_42308# 4.89e-20
C33424 a_16414_43172# a_15764_42576# 0.001182f
C33425 a_n2104_46634# VDD 0.286113f
C33426 a_626_44172# a_766_43646# 9.22e-19
C33427 a_10057_43914# a_10729_43914# 0.063518f
C33428 a_n2661_43922# a_n1899_43946# 0.00455f
C33429 a_n2293_43922# a_n1761_44111# 0.005057f
C33430 a_n2661_42834# a_n1331_43914# 0.01077f
C33431 a_8975_43940# a_10405_44172# 1.35e-19
C33432 a_6109_44484# a_5495_43940# 2.63e-20
C33433 a_n2661_46634# CLK_DATA 3.38e-19
C33434 a_3232_43370# a_3457_43396# 0.131408f
C33435 a_11823_42460# a_13113_42826# 0.003218f
C33436 a_n357_42282# a_11554_42852# 0.001921f
C33437 a_3537_45260# a_8685_43396# 0.023888f
C33438 a_n1059_45260# a_12281_43396# 0.025081f
C33439 a_n2293_42834# a_n2433_43396# 0.025997f
C33440 a_1307_43914# a_1987_43646# 0.002379f
C33441 a_5205_44484# a_6655_43762# 5.14e-19
C33442 a_526_44458# a_5267_42460# 3.04e-19
C33443 a_n1925_42282# a_3823_42558# 0.010285f
C33444 a_10903_43370# a_13249_42558# 0.003601f
C33445 a_8199_44636# a_9885_42308# 0.001301f
C33446 a_5111_44636# a_5837_43396# 7.68e-19
C33447 a_10193_42453# a_15567_42826# 1.05e-20
C33448 a_11967_42832# a_19615_44636# 0.065767f
C33449 a_3090_45724# a_n2017_45002# 2.3e-19
C33450 a_19692_46634# a_19963_31679# 1.27e-19
C33451 a_11189_46129# a_7499_43078# 5.71e-20
C33452 a_9290_44172# a_9049_44484# 1.37e-20
C33453 a_9625_46129# a_8746_45002# 4.27e-19
C33454 a_6755_46942# a_6171_45002# 0.026424f
C33455 a_4791_45118# a_8855_44734# 3.24e-21
C33456 a_12741_44636# a_15765_45572# 4.82e-19
C33457 a_11415_45002# a_16855_45546# 0.004485f
C33458 a_19123_46287# a_18909_45814# 5.82e-19
C33459 a_10227_46804# a_15004_44636# 0.003988f
C33460 a_11599_46634# a_18989_43940# 7.89e-20
C33461 a_n2438_43548# a_n2661_43370# 0.147387f
C33462 a_13747_46662# a_18315_45260# 1.26e-20
C33463 a_13661_43548# a_18587_45118# 0.087703f
C33464 a_5807_45002# a_18911_45144# 2.35e-20
C33465 a_17339_46660# a_18596_45572# 0.009893f
C33466 a_4646_46812# a_1423_45028# 0.415897f
C33467 a_10355_46116# a_10053_45546# 1.96e-19
C33468 a_9823_46155# a_10180_45724# 0.002058f
C33469 a_12891_46348# a_11691_44458# 0.141379f
C33470 a_n1151_42308# a_556_44484# 9.41e-20
C33471 a_16327_47482# a_17970_44736# 0.219775f
C33472 a_15567_42826# VDD 0.163583f
C33473 a_15764_42576# a_7174_31319# 6.35e-20
C33474 a_n3674_37592# a_n4064_37984# 0.020548f
C33475 a_16197_42308# a_4958_30871# 9.31e-19
C33476 a_5342_30871# RST_Z 0.048618f
C33477 a_6123_31319# a_n4209_39304# 5.16e-21
C33478 a_19478_44306# a_11341_43940# 6.59e-19
C33479 a_1307_43914# a_4649_42852# 1.56e-19
C33480 a_n2956_38216# a_n3565_38216# 0.307285f
C33481 a_n2017_45002# a_n2472_42282# 0.001176f
C33482 a_20365_43914# a_20623_43914# 0.22264f
C33483 a_12429_44172# a_12603_44260# 0.011572f
C33484 a_3499_42826# a_3992_43940# 2.6e-19
C33485 a_9569_46155# VDD 0.19288f
C33486 a_6419_46155# DATA[3] 9.23e-21
C33487 a_n1549_44318# a_n1177_43370# 0.003012f
C33488 a_n1331_43914# a_n1352_43396# 1.74e-20
C33489 a_n1761_44111# a_n97_42460# 0.001173f
C33490 a_10193_42453# a_20712_42282# 0.157661f
C33491 a_n2810_45572# a_n2946_37984# 0.020842f
C33492 a_19328_44172# a_15493_43940# 0.062184f
C33493 a_19862_44208# a_21115_43940# 0.064973f
C33494 a_14539_43914# a_17433_43396# 1.68e-19
C33495 a_n356_44636# a_15743_43084# 2.51e-20
C33496 a_7499_43078# a_11136_45572# 1.89e-21
C33497 a_2711_45572# a_14033_45572# 6.82e-19
C33498 a_16388_46812# a_18287_44626# 4.61e-22
C33499 a_20205_31679# a_22959_45572# 0.002292f
C33500 a_20692_30879# a_19963_31679# 0.051965f
C33501 a_2324_44458# a_6945_45348# 4.69e-19
C33502 a_n971_45724# a_n229_43646# 0.059197f
C33503 a_584_46384# a_n1177_43370# 2.93e-20
C33504 a_n2497_47436# a_3080_42308# 2.97e-19
C33505 a_8049_45260# a_6171_45002# 0.048422f
C33506 a_6755_46942# a_14673_44172# 0.050772f
C33507 a_13259_45724# en_comp 0.19355f
C33508 a_n2661_45546# a_2437_43646# 0.028152f
C33509 a_11962_45724# a_11682_45822# 0.014813f
C33510 a_11823_42460# a_10907_45822# 1.3e-19
C33511 a_10193_42453# a_10216_45572# 0.003165f
C33512 a_10053_45546# a_10544_45572# 0.00278f
C33513 a_10180_45724# a_10306_45572# 9.37e-19
C33514 a_n2293_46634# a_5663_43940# 5.03e-20
C33515 a_768_44030# a_7911_44260# 0.001075f
C33516 a_n4064_39616# C9_P_btm 0.215899f
C33517 a_n3420_39616# C7_P_btm 8.17e-19
C33518 a_11599_46634# a_5807_45002# 0.303048f
C33519 a_15507_47210# a_16131_47204# 9.73e-19
C33520 a_n3565_39304# a_n1532_35090# 1.16e-19
C33521 a_1239_47204# a_n2661_46098# 0.004048f
C33522 a_1431_47204# a_1799_45572# 3.57e-19
C33523 a_584_46384# a_479_46660# 1.75e-20
C33524 a_n443_46116# a_n133_46660# 1e-19
C33525 a_7754_39964# a_7754_38470# 0.241119f
C33526 a_20712_42282# VDD 0.282526f
C33527 a_n3565_39590# C5_P_btm 1.31e-19
C33528 a_16241_47178# a_16285_47570# 3.69e-19
C33529 a_14311_47204# a_13747_46662# 2.25e-21
C33530 a_4883_46098# a_n1613_43370# 0.025959f
C33531 a_n1151_42308# a_2107_46812# 0.073605f
C33532 a_6151_47436# a_n1925_46634# 0.052327f
C33533 a_3754_39134# a_3754_38802# 0.296258f
C33534 a_3754_39466# VDAC_Ni 0.001054f
C33535 a_n3420_37984# a_n3607_37440# 2.09e-19
C33536 a_12861_44030# a_19321_45002# 0.10527f
C33537 a_6575_47204# a_n2661_46634# 6.01e-19
C33538 a_13717_47436# a_19594_46812# 3.95e-20
C33539 a_n971_45724# a_2864_46660# 1.42e-20
C33540 a_n237_47217# a_3699_46634# 1.03e-19
C33541 a_20107_42308# RST_Z 4.07e-20
C33542 a_15673_47210# a_16697_47582# 2.36e-20
C33543 a_10227_46804# a_768_44030# 0.050994f
C33544 a_18143_47464# a_12549_44172# 0.0015f
C33545 a_3626_43646# a_7287_43370# 2.15e-20
C33546 a_2982_43646# a_8147_43396# 1.75e-21
C33547 a_14021_43940# a_21487_43396# 0.023941f
C33548 a_n356_44636# a_1606_42308# 0.282657f
C33549 a_3080_42308# a_4181_43396# 2.84e-19
C33550 a_11967_42832# a_11229_43218# 3.74e-21
C33551 a_10216_45572# VDD 4.83e-19
C33552 a_n97_42460# a_14579_43548# 0.001021f
C33553 a_18494_42460# a_17124_42282# 4.91e-20
C33554 a_22959_43948# a_17364_32525# 0.005227f
C33555 a_3357_43084# a_3232_43370# 0.118744f
C33556 a_12549_44172# a_21259_43561# 0.001855f
C33557 a_n1613_43370# a_5649_42852# 2.17e-20
C33558 a_2711_45572# a_6298_44484# 6.39e-20
C33559 a_n443_42852# a_13076_44458# 4.94e-19
C33560 a_12427_45724# a_11827_44484# 3.2e-21
C33561 a_11322_45546# a_11691_44458# 1.74e-19
C33562 a_10193_42453# a_16886_45144# 0.001731f
C33563 a_n967_45348# a_n955_45028# 0.014419f
C33564 a_n2293_46634# a_16243_43396# 1.28e-22
C33565 a_20202_43084# a_20269_44172# 9.29e-21
C33566 a_5937_45572# a_7281_43914# 9.58e-19
C33567 a_n745_45366# a_413_45260# 4.33e-20
C33568 a_8049_45260# a_14673_44172# 8.94e-21
C33569 a_11415_45002# a_19862_44208# 1.39e-19
C33570 a_n863_45724# a_n310_44811# 5.09e-19
C33571 a_380_45546# a_n356_44636# 5.74e-21
C33572 a_22959_47212# a_12741_44636# 3.06e-19
C33573 a_11453_44696# a_22959_46660# 4.6e-19
C33574 a_5257_43370# a_7411_46660# 1.2e-20
C33575 a_4646_46812# a_6682_46987# 8.46e-19
C33576 a_n743_46660# a_15227_44166# 3.07e-19
C33577 a_12549_44172# a_765_45546# 0.118284f
C33578 SMPL_ON_N a_21076_30879# 0.030428f
C33579 a_4651_46660# a_6969_46634# 2.71e-21
C33580 a_n1435_47204# a_5204_45822# 1.65e-20
C33581 a_6575_47204# a_8199_44636# 1.83e-20
C33582 a_9863_47436# a_8016_46348# 8.34e-20
C33583 a_4883_46098# a_n2293_46098# 0.009323f
C33584 VREF VCM 45.073803f
C33585 a_5807_45002# a_13693_46688# 5.45e-19
C33586 a_13747_46662# a_14226_46987# 4.64e-19
C33587 a_n2497_47436# a_n1545_46494# 0.001346f
C33588 a_n2840_43370# a_n3674_38680# 0.003987f
C33589 a_743_42282# a_3681_42891# 1.37e-20
C33590 a_18114_32519# C3_N_btm 1.27e-19
C33591 a_19721_31679# C2_N_btm 0.040789f
C33592 a_n1991_42858# a_n1423_42826# 0.186387f
C33593 a_n2157_42858# a_n901_43156# 0.043475f
C33594 a_n1853_43023# a_n1641_43230# 0.036072f
C33595 a_10341_43396# a_21671_42860# 1.14e-19
C33596 a_3422_30871# a_n3420_39072# 0.096346f
C33597 a_16137_43396# a_15567_42826# 6.67e-19
C33598 a_3090_45724# a_19164_43230# 4.01e-21
C33599 a_5111_44636# a_8375_44464# 0.001962f
C33600 a_5147_45002# a_5891_43370# 0.049542f
C33601 a_7499_43078# a_11750_44172# 0.195997f
C33602 a_20107_45572# a_20159_44458# 2.4e-19
C33603 a_n2442_46660# a_n3674_37592# 0.032368f
C33604 a_9290_44172# a_13749_43396# 0.00194f
C33605 a_n1613_43370# a_7963_42308# 5.32e-20
C33606 a_n2293_42834# a_n2433_44484# 4.65e-21
C33607 a_18315_45260# a_18911_45144# 7.05e-19
C33608 a_16922_45042# a_20567_45036# 0.002083f
C33609 a_n967_45348# a_n2661_42834# 0.027185f
C33610 en_comp a_n2661_43922# 0.237031f
C33611 a_n2956_37592# a_n2293_43922# 2.05e-20
C33612 a_21513_45002# a_17517_44484# 2.37e-19
C33613 a_327_44734# a_556_44484# 0.033015f
C33614 a_1307_43914# a_15004_44636# 1.02e-20
C33615 a_16019_45002# a_16112_44458# 3.78e-19
C33616 a_n357_42282# a_7499_43940# 8.54e-20
C33617 SMPL_ON_P a_n4209_39304# 0.001361f
C33618 a_15227_44166# a_17701_42308# 0.172697f
C33619 a_n2661_46634# a_n2661_45546# 5.96e-19
C33620 a_3090_45724# a_13759_46122# 5.3e-22
C33621 a_15009_46634# a_13925_46122# 1.53e-19
C33622 a_15368_46634# a_12594_46348# 1.41e-21
C33623 a_11599_46634# a_15143_45578# 0.028879f
C33624 a_12891_46348# a_n443_42852# 7.66e-20
C33625 a_n2840_46634# a_n2956_38216# 0.001369f
C33626 a_20719_46660# a_20202_43084# 4.3e-21
C33627 a_765_45546# a_1208_46090# 0.134766f
C33628 a_10227_46804# a_11652_45724# 2.55e-20
C33629 a_15743_43084# a_18727_42674# 1.5e-19
C33630 a_743_42282# a_15959_42545# 0.006675f
C33631 a_22959_42860# a_14097_32519# 0.166017f
C33632 a_10405_44172# VDD 0.408512f
C33633 a_16867_43762# a_4958_30871# 4.18e-20
C33634 a_21195_42852# a_20753_42852# 7.65e-19
C33635 a_5111_42852# a_4921_42308# 3.76e-20
C33636 a_4361_42308# a_14113_42308# 0.075467f
C33637 a_18479_47436# SINGLE_ENDED 0.040779f
C33638 a_n443_42852# a_4520_42826# 5.33e-20
C33639 a_13259_45724# a_22165_42308# 0.001551f
C33640 a_n967_45348# a_n1352_43396# 0.010028f
C33641 a_18248_44752# a_20679_44626# 1.77e-21
C33642 a_10617_44484# a_n2661_43922# 0.004461f
C33643 a_n1177_44458# a_n1549_44318# 0.004943f
C33644 a_n1352_44484# a_n1331_43914# 7.59e-19
C33645 a_15673_47210# CLK 3.17e-19
C33646 a_19386_47436# VDD 0.121241f
C33647 a_18597_46090# RST_Z 1.14e-19
C33648 a_18989_43940# a_19615_44636# 8.51e-19
C33649 a_n2661_45010# a_1209_43370# 9.39e-22
C33650 a_n2017_45002# a_n1821_43396# 0.001012f
C33651 a_3357_43084# a_4905_42826# 0.062628f
C33652 a_1307_43914# a_1241_43940# 0.038832f
C33653 a_18780_47178# START 0.01578f
C33654 a_n357_42282# a_10991_42826# 0.005156f
C33655 a_10193_42453# a_20556_43646# 1.67e-19
C33656 a_7499_43078# a_4361_42308# 0.04291f
C33657 a_10227_46804# a_13490_45067# 6.94e-20
C33658 a_11599_46634# a_18315_45260# 2.46e-20
C33659 a_2324_44458# a_13259_45724# 0.068761f
C33660 a_768_44030# a_1307_43914# 1.13357f
C33661 a_12549_44172# a_16751_45260# 6.99e-22
C33662 a_n237_47217# a_4743_44484# 1.26e-21
C33663 a_4419_46090# a_n755_45592# 0.0037f
C33664 a_805_46414# a_n443_42852# 0.003153f
C33665 a_n2661_46634# a_5205_44484# 1.71e-21
C33666 a_288_46660# a_n37_45144# 1e-20
C33667 a_n1925_46634# a_5111_44636# 2.77e-20
C33668 a_4651_46660# a_3357_43084# 0.004361f
C33669 a_5807_45002# a_13348_45260# 9.82e-22
C33670 a_167_45260# a_n23_45546# 0.001656f
C33671 a_3147_46376# a_3218_45724# 0.0111f
C33672 a_13059_46348# a_13249_42308# 0.306398f
C33673 a_14976_45028# a_15225_45822# 5.88e-19
C33674 a_3090_45724# a_15297_45822# 8.48e-19
C33675 a_12861_44030# a_18184_42460# 0.266953f
C33676 a_5385_46902# a_2437_43646# 7.1e-20
C33677 a_n1151_42308# a_n2661_44458# 0.030695f
C33678 a_n2293_46634# a_3232_43370# 0.046281f
C33679 a_16327_47482# a_16501_45348# 5.1e-19
C33680 a_20556_43646# VDD 0.34939f
C33681 a_13678_32519# C6_N_btm 1.22e-19
C33682 a_743_42282# RST_Z 2.55e-19
C33683 a_14209_32519# C1_N_btm 4.13e-20
C33684 a_9803_42558# a_10533_42308# 5.35e-19
C33685 a_8685_42308# a_5742_30871# 4.1e-20
C33686 COMP_P a_22775_42308# 4.23e-19
C33687 a_13887_32519# C3_N_btm 0.030933f
C33688 a_11827_44484# a_17324_43396# 2.91e-21
C33689 a_18184_42460# a_19700_43370# 0.003845f
C33690 a_9482_43914# a_10083_42826# 4.71e-19
C33691 a_8701_44490# a_8685_43396# 1.11e-20
C33692 a_n356_44636# a_3539_42460# 1.86e-19
C33693 a_19551_46910# VDD 0.226848f
C33694 a_21076_30879# a_19864_35138# 5.61e-20
C33695 a_18285_46348# START 0.001916f
C33696 a_7845_44172# a_7911_44260# 0.010598f
C33697 a_7542_44172# a_8018_44260# 0.001923f
C33698 a_4185_45028# a_22469_40625# 1.54e-20
C33699 a_19123_46287# RST_Z 4.05e-21
C33700 a_18494_42460# a_19268_43646# 5.16e-21
C33701 a_n967_45348# a_n2293_42282# 5.08e-19
C33702 a_5343_44458# a_8317_43396# 1.12e-19
C33703 a_n357_42282# a_17303_42282# 4.34e-19
C33704 a_n913_45002# a_133_42852# 0.046777f
C33705 a_19237_31679# a_22959_43948# 5.09e-19
C33706 a_5708_44484# a_n97_42460# 4.19e-21
C33707 a_n2661_42834# a_n1917_43396# 0.007372f
C33708 a_n2293_43922# a_n2267_43396# 0.020404f
C33709 a_1307_43914# a_5755_42852# 2.6e-19
C33710 a_11691_44458# a_16409_43396# 6.27e-20
C33711 a_2711_45572# a_5437_45600# 5.64e-19
C33712 a_4646_46812# a_6109_44484# 0.010238f
C33713 a_16375_45002# a_15765_45572# 2.15e-19
C33714 a_13259_45724# a_16855_45546# 0.067694f
C33715 a_13661_43548# a_11967_42832# 0.165876f
C33716 a_5807_45002# a_19615_44636# 0.003455f
C33717 a_3483_46348# a_9482_43914# 0.130172f
C33718 a_8953_45546# a_6171_45002# 0.0298f
C33719 a_5937_45572# a_6431_45366# 0.129839f
C33720 a_15227_44166# a_17969_45144# 5.42e-19
C33721 a_8049_45260# a_18909_45814# 0.006015f
C33722 a_8199_44636# a_5205_44484# 1.08e-20
C33723 a_13717_47436# a_15673_47210# 1.97e-19
C33724 a_12861_44030# a_15811_47375# 0.144648f
C33725 a_n2946_38778# a_n4064_38528# 0.053228f
C33726 a_n3420_38528# a_n2302_38778# 1.28e-19
C33727 a_6171_42473# VDD 0.184622f
C33728 a_5934_30871# C4_N_btm 0.030578f
C33729 a_7174_31319# a_n4064_37440# 1.84e-19
C33730 a_n2109_47186# a_5159_47243# 0.00107f
C33731 a_n1741_47186# a_7989_47542# 4.61e-19
C33732 a_5742_30871# C10_P_btm 0.00237f
C33733 a_584_46384# a_2266_47570# 9.67e-19
C33734 a_6123_31319# C6_N_btm 6.31e-19
C33735 a_4791_45118# a_4883_46098# 0.135093f
C33736 a_17303_42282# CAL_N 0.003472f
C33737 a_n1151_42308# a_11453_44696# 2.35e-21
C33738 a_4915_47217# a_13507_46334# 0.032373f
C33739 a_14311_47204# a_11599_46634# 4.05e-22
C33740 a_11341_43940# a_13667_43396# 9.28e-19
C33741 a_5663_43940# a_743_42282# 7.52e-22
C33742 a_n1899_43946# a_n1641_43230# 3.58e-20
C33743 a_n809_44244# a_n1853_43023# 4.45e-20
C33744 a_n2065_43946# a_n1076_43230# 2.53e-21
C33745 a_n1549_44318# a_n1991_42858# 6.41e-19
C33746 a_n1761_44111# a_n901_43156# 0.013702f
C33747 a_1990_45899# VDD 0.001563f
C33748 a_n2810_45028# a_n2946_39866# 5.51e-20
C33749 a_19478_44306# a_10341_43396# 5.01e-20
C33750 a_n4318_40392# a_n3674_38680# 0.023225f
C33751 a_n2433_43396# a_n2012_43396# 0.089677f
C33752 a_n1917_43396# a_n1352_43396# 7.99e-20
C33753 a_n4318_39304# a_n1809_43762# 1.53e-19
C33754 a_n2129_43609# a_104_43370# 3.36e-19
C33755 a_n2956_37592# a_n3420_39616# 3.18e-19
C33756 a_11967_42832# a_10835_43094# 0.263495f
C33757 a_5257_43370# a_5829_43940# 0.003839f
C33758 a_n2438_43548# a_1568_43370# 4.4e-21
C33759 a_14495_45572# a_9482_43914# 2.35e-20
C33760 a_13249_42308# a_13556_45296# 0.059719f
C33761 a_13904_45546# a_13777_45326# 1.68e-19
C33762 a_13759_46122# a_14815_43914# 1.02e-21
C33763 a_8049_45260# a_12607_44458# 7.47e-21
C33764 a_2324_44458# a_n2661_43922# 0.088002f
C33765 a_n1613_43370# a_8685_43396# 0.016726f
C33766 a_8791_45572# a_6171_45002# 6.13e-19
C33767 a_4185_45028# a_11967_42832# 2.11e-19
C33768 a_16327_47482# a_18783_43370# 0.026485f
C33769 a_4791_45118# a_5649_42852# 0.075725f
C33770 a_526_44458# a_n356_44636# 0.142971f
C33771 a_20107_45572# a_20623_45572# 0.103168f
C33772 a_20273_45572# a_20841_45814# 0.175891f
C33773 a_3090_45724# a_18079_43940# 8.6e-20
C33774 a_768_44030# a_9396_43370# 0.010156f
C33775 a_n2293_46634# a_4905_42826# 0.024749f
C33776 a_6755_46942# a_14761_44260# 2.19e-20
C33777 a_10227_46804# a_10933_46660# 0.00489f
C33778 a_15811_47375# a_14180_46812# 2.14e-19
C33779 a_11309_47204# a_10249_46116# 0.033926f
C33780 a_13717_47436# a_16388_46812# 4.02e-20
C33781 a_12861_44030# a_13059_46348# 0.504219f
C33782 a_12465_44636# a_15368_46634# 7.1e-20
C33783 C6_P_btm C3_P_btm 0.134599f
C33784 C7_P_btm C2_P_btm 0.139982f
C33785 C5_P_btm C4_P_btm 15.915401f
C33786 C9_P_btm C0_P_btm 0.14782f
C33787 C8_P_btm C1_P_btm 0.131002f
C33788 a_n2661_46634# a_5385_46902# 0.007092f
C33789 a_5807_45002# a_7411_46660# 0.006898f
C33790 EN_VIN_BSTR_N C3_N_btm 0.100325f
C33791 a_n1741_47186# a_n1853_46287# 1.65e-19
C33792 a_6575_47204# a_765_45546# 0.061901f
C33793 a_4883_46098# a_16292_46812# 1.69e-20
C33794 a_19787_47423# a_19692_46634# 5.22e-20
C33795 a_2107_46812# a_3177_46902# 0.001642f
C33796 a_491_47026# a_n2661_46098# 6.63e-19
C33797 a_13507_46334# a_18834_46812# 0.004721f
C33798 a_21177_47436# a_15227_44166# 9.06e-22
C33799 C10_P_btm C0_dummy_P_btm 0.63636f
C33800 a_n1613_43370# a_6682_46660# 7.54e-19
C33801 a_n881_46662# a_8035_47026# 0.003736f
C33802 a_22717_37285# VDD 3.6e-19
C33803 a_n1925_46634# a_3221_46660# 6.56e-19
C33804 a_5013_44260# a_5932_42308# 4.06e-21
C33805 a_3499_42826# a_1755_42282# 2.38e-20
C33806 a_n2661_42282# a_961_42354# 1.35e-19
C33807 a_5663_43940# a_5755_42308# 1e-20
C33808 a_3626_43646# a_12089_42308# 0.002196f
C33809 a_2982_43646# a_13113_42826# 1.09e-20
C33810 a_8147_43396# a_7871_42858# 1.53e-19
C33811 a_11967_42832# a_16269_42308# 6.4e-20
C33812 a_16243_43396# a_743_42282# 7.51e-20
C33813 a_15781_43660# a_4361_42308# 1.85e-20
C33814 a_16409_43396# a_4190_30871# 4.44e-21
C33815 a_15743_43084# a_17486_43762# 2.49e-19
C33816 a_17499_43370# a_17678_43396# 0.007399f
C33817 a_17324_43396# a_17433_43396# 0.007416f
C33818 a_18429_43548# a_16823_43084# 0.130506f
C33819 a_n1917_43396# a_n2293_42282# 9.44e-21
C33820 a_17339_46660# a_16759_43396# 7.48e-21
C33821 a_11415_45002# a_14579_43548# 4.66e-21
C33822 a_5009_45028# a_5093_45028# 0.092725f
C33823 a_n467_45028# a_n1699_44726# 1.68e-21
C33824 a_8696_44636# a_11649_44734# 5.17e-19
C33825 a_19692_46634# a_21487_43396# 0.016698f
C33826 a_n357_42282# a_2253_44260# 1.12e-19
C33827 a_n1059_45260# a_n699_43396# 0.021143f
C33828 a_n913_45002# a_4223_44672# 6.25e-20
C33829 a_13507_46334# COMP_P 2.67e-20
C33830 a_15227_44166# a_4361_42308# 2.26e-19
C33831 a_n967_45348# a_n1352_44484# 0.007805f
C33832 a_327_44734# a_n2661_44458# 0.027103f
C33833 a_3483_46348# a_6031_43396# 5.46e-22
C33834 a_2711_45572# a_2479_44172# 9.28e-20
C33835 a_13259_45724# a_19862_44208# 1.06e-20
C33836 a_5275_47026# a_5497_46414# 7.81e-20
C33837 a_6540_46812# a_6419_46155# 7.76e-19
C33838 a_4007_47204# a_2711_45572# 9.84e-20
C33839 a_n443_46116# a_1176_45572# 0.003318f
C33840 a_9804_47204# a_9823_46482# 0.006171f
C33841 a_7715_46873# a_3483_46348# 2.08e-20
C33842 a_15227_44166# a_20841_46902# 1.43e-19
C33843 a_14180_46812# a_13059_46348# 0.074456f
C33844 a_19333_46634# a_20273_46660# 1.31e-19
C33845 a_n2312_38680# a_n1736_46482# 1.05e-19
C33846 a_768_44030# a_8034_45724# 4.91e-21
C33847 a_5257_43370# a_4185_45028# 9.55e-20
C33848 a_4883_46098# a_20254_46482# 1.42e-19
C33849 a_13507_46334# a_20850_46482# 9.11e-19
C33850 a_19466_46812# a_20411_46873# 0.001378f
C33851 a_19692_46634# a_20107_46660# 0.126737f
C33852 a_n1151_42308# a_5907_45546# 6.31e-20
C33853 a_2063_45854# a_6598_45938# 0.018518f
C33854 a_20980_44850# VDD 0.132317f
C33855 a_17730_32519# C1_N_btm 3.84e-20
C33856 a_10796_42968# a_10793_43218# 2.36e-20
C33857 a_3626_43646# a_18907_42674# 0.003037f
C33858 a_3422_30871# C10_N_btm 0.002966f
C33859 a_n913_45002# a_15493_43940# 1.64e-20
C33860 a_8701_44490# a_8783_44734# 0.004999f
C33861 a_18587_45118# a_11967_42832# 4.11e-20
C33862 a_18911_45144# a_19006_44850# 3.38e-19
C33863 a_16922_45042# a_20679_44626# 5.14e-20
C33864 a_3232_43370# a_9672_43914# 4.68e-20
C33865 a_n443_42852# a_16409_43396# 2.64e-19
C33866 a_n2442_46660# a_n2302_39072# 1.26e-19
C33867 a_6755_46942# a_15959_42545# 9.08e-38
C33868 a_10157_44484# a_5891_43370# 0.001885f
C33869 a_n1699_44726# a_n2661_43922# 0.006002f
C33870 a_n1917_44484# a_n2661_42834# 0.002676f
C33871 a_n2267_44484# a_n2293_43922# 6.94e-19
C33872 a_2779_44458# a_3363_44484# 0.020864f
C33873 a_1307_43914# a_7845_44172# 0.002954f
C33874 a_11691_44458# a_16241_44734# 4.13e-19
C33875 a_7229_43940# a_7584_44260# 0.001386f
C33876 w_11334_34010# RST_Z 0.00509f
C33877 a_11827_44484# a_15146_44484# 1.1e-19
C33878 a_1423_45028# a_5013_44260# 3.14e-20
C33879 a_n699_43396# a_484_44484# 1.33e-19
C33880 a_n2833_47464# VDD 0.461379f
C33881 a_15682_46116# a_17715_44484# 0.003258f
C33882 a_10467_46802# a_11652_45724# 4.42e-19
C33883 a_3090_45724# a_4099_45572# 0.004385f
C33884 a_15368_46634# a_2711_45572# 0.0051f
C33885 a_6755_46942# a_8746_45002# 4.26e-20
C33886 a_13747_46662# a_20107_45572# 0.012917f
C33887 a_12891_46348# a_2437_43646# 0.004901f
C33888 a_12549_44172# a_21513_45002# 0.002562f
C33889 a_n743_46660# a_16377_45572# 5.01e-19
C33890 a_10903_43370# a_6945_45028# 1.05e-19
C33891 a_22959_47212# a_413_45260# 0.024836f
C33892 a_11599_46634# a_13017_45260# 1.1e-20
C33893 a_765_45546# a_n2661_45546# 0.006374f
C33894 a_12861_44030# a_13556_45296# 0.028687f
C33895 a_6545_47178# a_1423_45028# 4.56e-21
C33896 a_5204_45822# a_526_44458# 0.001107f
C33897 a_5164_46348# a_n1925_42282# 3.73e-20
C33898 a_n784_42308# a_6171_42473# 1.56e-20
C33899 a_3457_43396# VDD 0.004013f
C33900 a_1755_42282# a_3318_42354# 2.48e-19
C33901 a_1606_42308# a_3823_42558# 1.77e-20
C33902 a_2351_42308# a_2713_42308# 0.00357f
C33903 a_n2017_45002# a_n1736_43218# 0.0083f
C33904 a_n1177_44458# a_n1177_43370# 7.08e-19
C33905 a_n443_42852# a_564_42282# 0.005734f
C33906 a_3357_43084# a_2905_42968# 0.025927f
C33907 a_6969_46634# VDD 0.154507f
C33908 a_21359_45002# a_2982_43646# 3.84e-21
C33909 a_6755_46942# RST_Z 1.33e-19
C33910 en_comp a_n1641_43230# 6.37e-21
C33911 a_n967_45348# a_n1423_42826# 0.010397f
C33912 a_3232_43370# a_743_42282# 2.67e-20
C33913 a_n1761_44111# a_n984_44318# 0.056404f
C33914 a_n1899_43946# a_n809_44244# 0.042737f
C33915 a_n2065_43946# a_175_44278# 5.71e-21
C33916 a_n1331_43914# a_n1549_44318# 0.209641f
C33917 a_8704_45028# a_8685_43396# 1.1e-21
C33918 a_n755_45592# a_1848_45724# 0.030306f
C33919 a_n743_46660# a_9838_44484# 8.79e-21
C33920 a_19321_45002# a_18287_44626# 0.00979f
C33921 a_n2661_45546# a_509_45822# 4.99e-19
C33922 a_13661_43548# a_18989_43940# 0.039099f
C33923 a_17583_46090# a_8696_44636# 7.3e-19
C33924 a_15682_46116# a_15861_45028# 0.001207f
C33925 a_17715_44484# a_16680_45572# 0.001431f
C33926 a_12861_44030# a_20362_44736# 0.004923f
C33927 a_2107_46812# a_4223_44672# 3.28e-20
C33928 a_n2956_38216# a_n1013_45572# 2.26e-19
C33929 a_n2661_46634# a_13076_44458# 7.24e-19
C33930 a_8049_45260# a_8746_45002# 0.001752f
C33931 a_8270_45546# a_8488_45348# 3.69e-19
C33932 a_n746_45260# a_453_43940# 0.004985f
C33933 a_n2312_39304# a_n2293_43922# 5.35e-20
C33934 a_n863_45724# a_n23_45546# 4.47e-19
C33935 a_n452_45724# a_n356_45724# 0.318161f
C33936 a_20202_43084# en_comp 6.61e-20
C33937 a_n237_47217# a_1414_42308# 8.74e-23
C33938 a_10903_43370# a_14127_45572# 0.003658f
C33939 a_14035_46660# a_13777_45326# 4.08e-20
C33940 a_n2293_46634# a_8975_43940# 1.9e-19
C33941 a_5932_42308# a_n4064_37440# 1.17e-19
C33942 COMP_P a_n923_35174# 0.003051f
C33943 a_n971_45724# a_3815_47204# 0.04068f
C33944 a_n23_47502# a_n1151_42308# 0.005195f
C33945 a_2124_47436# a_584_46384# 0.220021f
C33946 a_n1741_47186# a_4915_47217# 0.128899f
C33947 a_n2109_47186# a_5815_47464# 0.00257f
C33948 a_1209_47178# a_2952_47436# 4.55e-19
C33949 a_1431_47204# a_2063_45854# 1.97e-19
C33950 a_4958_30871# a_n3420_38528# 0.030871f
C33951 a_n4209_39590# a_n3565_39590# 6.15218f
C33952 a_n4064_40160# a_n4064_39616# 5.80394f
C33953 a_13720_44458# a_13460_43230# 1.78e-21
C33954 a_5745_43940# a_5829_43940# 0.092725f
C33955 a_3232_43370# a_5755_42308# 2.19e-21
C33956 a_n913_45002# a_5742_30871# 0.028271f
C33957 a_n1059_45260# a_11551_42558# 9.25e-20
C33958 a_n2661_42282# a_2982_43646# 0.076578f
C33959 a_n2293_43922# a_n2472_42826# 1.92e-19
C33960 a_n2661_42834# a_n1853_43023# 0.002855f
C33961 a_n2661_43922# a_n2157_42858# 2.6e-21
C33962 a_2382_45260# a_3905_42308# 4.58e-19
C33963 a_20679_44626# a_15743_43084# 9.47e-21
C33964 a_n356_44636# a_8605_42826# 1.43e-20
C33965 a_1307_43914# a_1067_42314# 3.75e-21
C33966 a_375_42282# a_564_42282# 0.022891f
C33967 a_8049_45260# RST_Z 0.002763f
C33968 a_n2017_45002# a_11633_42558# 0.005942f
C33969 a_3537_45260# a_6123_31319# 9.93e-19
C33970 a_3065_45002# a_5934_30871# 1.09e-20
C33971 a_19478_44306# a_n97_42460# 6.27e-19
C33972 a_167_45260# a_n23_44458# 7.57e-19
C33973 a_16333_45814# a_16223_45938# 0.097745f
C33974 a_16680_45572# a_15861_45028# 1.57e-19
C33975 a_16855_45546# a_17478_45572# 3.95e-19
C33976 a_16115_45572# a_16020_45572# 0.049827f
C33977 a_4791_45118# a_8685_43396# 4.61e-21
C33978 a_5807_45002# a_5829_43940# 8.28e-21
C33979 a_2711_45572# a_2680_45002# 2.69e-19
C33980 a_14033_45822# a_14033_45572# 6.96e-20
C33981 a_16327_47482# a_3626_43646# 3.96e-19
C33982 a_10586_45546# a_n2661_43370# 0.002741f
C33983 a_17339_46660# a_17517_44484# 0.020067f
C33984 a_n4064_38528# VREF 2.95e-20
C33985 a_2063_45854# a_11735_46660# 8.71e-19
C33986 a_6151_47436# a_6999_46987# 0.001316f
C33987 a_n881_46662# a_n2438_43548# 0.080298f
C33988 a_n1613_43370# a_n133_46660# 0.347805f
C33989 CAL_N a_22521_40055# 6.29e-19
C33990 a_22521_40599# a_22780_40945# 0.009658f
C33991 a_n3420_38528# VCM 0.00888f
C33992 a_n1435_47204# a_7927_46660# 2.14e-20
C33993 a_9313_45822# a_9863_46634# 1.77e-19
C33994 a_6851_47204# a_6755_46942# 8.96e-19
C33995 a_3726_37500# CAL_P 0.102027f
C33996 a_12891_46348# a_n2661_46634# 1.07e-19
C33997 a_5807_45002# a_13661_43548# 0.062335f
C33998 a_n2302_37984# VDD 0.350854f
C33999 a_n2312_39304# a_n2661_46098# 0.006111f
C34000 a_n2661_42282# a_5837_42852# 0.002566f
C34001 a_3357_43084# VDD 1.66202f
C34002 a_19963_31679# C10_N_btm 2.25e-20
C34003 a_15493_43940# a_20922_43172# 1.71e-21
C34004 a_11341_43940# a_21195_42852# 4.62e-21
C34005 a_2982_43646# a_16823_43084# 1.31e-20
C34006 a_13667_43396# a_10341_43396# 0.007486f
C34007 a_10695_43548# a_10765_43646# 0.011552f
C34008 a_19479_31679# RST_Z 0.049574f
C34009 a_n2293_43922# a_9223_42460# 4.38e-20
C34010 a_9313_44734# a_13070_42354# 3.27e-21
C34011 a_14021_43940# a_15567_42826# 4.16e-20
C34012 a_14205_43396# a_15095_43370# 0.086245f
C34013 a_9145_43396# a_12293_43646# 0.003544f
C34014 a_2437_43646# SINGLE_ENDED 0.117817f
C34015 a_n2840_43370# a_n4318_38680# 0.001904f
C34016 a_n1917_43396# a_n1423_42826# 0.001812f
C34017 a_n1352_43396# a_n1853_43023# 5.05e-20
C34018 a_n1177_43370# a_n1991_42858# 0.003015f
C34019 a_n2129_43609# a_n1076_43230# 3.31e-20
C34020 a_n4318_39304# a_n3674_39304# 2.9537f
C34021 a_4905_42826# a_743_42282# 0.0175f
C34022 a_20447_31679# C8_N_btm 5.41e-20
C34023 a_768_44030# a_13635_43156# 5.26e-19
C34024 SMPL_ON_P a_n4318_37592# 0.040097f
C34025 a_13017_45260# a_13348_45260# 0.044101f
C34026 a_11963_45334# a_9482_43914# 2.68e-20
C34027 a_4927_45028# a_1423_45028# 1.19e-20
C34028 a_n357_42282# a_20159_44458# 5.88e-21
C34029 a_3537_45260# a_3495_45348# 7.3e-19
C34030 a_n1925_42282# a_3499_42826# 4.47e-20
C34031 a_n37_45144# a_45_45144# 0.004937f
C34032 a_10809_44734# a_12429_44172# 2.57e-21
C34033 a_19431_45546# a_19113_45348# 0.001195f
C34034 a_n913_45002# a_n2293_42834# 0.055202f
C34035 a_18691_45572# a_11691_44458# 7.43e-20
C34036 a_20528_45572# a_16922_45042# 7.24e-19
C34037 a_n2497_47436# a_196_42282# 4.06e-22
C34038 a_9290_44172# a_12710_44260# 1.37e-19
C34039 a_10903_43370# a_11173_44260# 0.035423f
C34040 a_6755_46942# a_16243_43396# 4.46e-20
C34041 a_8034_45724# a_7845_44172# 2.09e-21
C34042 a_3429_45260# a_3602_45348# 0.007688f
C34043 a_7499_43078# a_5891_43370# 1.00892f
C34044 a_5385_46902# a_765_45546# 0.001698f
C34045 a_n881_46662# a_11133_46155# 4.96e-21
C34046 a_13507_46334# a_10809_44734# 0.603934f
C34047 a_n1021_46688# a_n1991_46122# 1.13e-19
C34048 a_n2438_43548# a_n2157_46122# 0.270054f
C34049 a_n133_46660# a_n2293_46098# 8.67e-21
C34050 a_n2293_46634# a_n1076_46494# 2.06e-20
C34051 a_768_44030# a_8016_46348# 0.034453f
C34052 a_4915_47217# a_10586_45546# 2.07e-20
C34053 a_10249_46116# a_12156_46660# 1.26e-19
C34054 a_10623_46897# a_10861_46660# 0.001705f
C34055 a_6755_46942# a_10425_46660# 2.19e-19
C34056 a_9804_47204# a_9569_46155# 0.040648f
C34057 a_11813_46116# a_11901_46660# 0.211542f
C34058 a_11735_46660# a_12469_46902# 0.053479f
C34059 a_12465_44636# a_20708_46348# 4.4e-21
C34060 a_13747_46662# a_3483_46348# 3.96e-19
C34061 a_5807_45002# a_4185_45028# 5.59e-20
C34062 a_n743_46660# a_n1853_46287# 6.94e-19
C34063 a_n1925_46634# a_n1423_46090# 0.005255f
C34064 a_n2312_38680# a_n1641_46494# 2.29e-20
C34065 a_4883_46098# a_6945_45028# 0.083863f
C34066 a_n97_42460# a_9223_42460# 0.004352f
C34067 a_4905_42826# a_5755_42308# 0.001861f
C34068 a_5826_44734# VDD 0.007376f
C34069 a_n1853_43023# a_n2293_42282# 4.92e-20
C34070 a_3539_42460# a_3823_42558# 0.07742f
C34071 a_3626_43646# a_5267_42460# 1.19e-19
C34072 a_14021_43940# a_20712_42282# 1.2e-20
C34073 a_10518_42984# a_10835_43094# 0.102355f
C34074 a_10083_42826# a_10796_42968# 0.042737f
C34075 a_11827_44484# a_16112_44458# 0.00849f
C34076 a_3357_43084# a_5495_43940# 0.004364f
C34077 a_4185_45028# a_10518_42984# 8.53e-21
C34078 a_20202_43084# a_22165_42308# 0.001287f
C34079 a_4646_46812# a_6171_42473# 2.16e-21
C34080 a_10193_42453# a_18533_44260# 0.003163f
C34081 a_n357_42282# a_6031_43396# 0.012855f
C34082 a_n967_45348# a_n1549_44318# 5.66e-19
C34083 a_n2661_45010# a_895_43940# 0.020382f
C34084 SMPL_ON_P a_n4334_37440# 4.8e-20
C34085 a_n443_42852# a_n1557_42282# 0.078868f
C34086 a_n2661_44458# a_4223_44672# 0.019953f
C34087 a_11691_44458# a_12883_44458# 0.058264f
C34088 a_n1917_44484# a_n1352_44484# 7.99e-20
C34089 a_14537_43396# a_16335_44484# 0.003972f
C34090 a_n2017_45002# a_1414_42308# 0.015426f
C34091 a_n913_45002# a_1115_44172# 1.07e-21
C34092 a_n2312_39304# a_n3420_39616# 1.17e-19
C34093 a_n2312_40392# a_n2946_39866# 2.19e-20
C34094 a_n971_45724# a_2382_45260# 0.019144f
C34095 a_6491_46660# a_3357_43084# 0.014978f
C34096 a_n743_46660# a_8568_45546# 3.92e-20
C34097 a_13747_46662# a_14495_45572# 0.288916f
C34098 a_n2109_47186# a_5147_45002# 0.05864f
C34099 a_20623_46660# a_10809_44734# 0.008272f
C34100 a_21188_46660# a_6945_45028# 0.004363f
C34101 a_7903_47542# a_2437_43646# 0.006626f
C34102 a_12861_44030# a_21363_45546# 1.6e-22
C34103 a_18597_46090# a_18341_45572# 0.010006f
C34104 a_11599_46634# a_20107_45572# 0.246047f
C34105 a_n1925_46634# a_9049_44484# 2.71e-20
C34106 a_n2293_46634# a_10193_42453# 0.037794f
C34107 a_3483_46348# a_4419_46090# 0.218073f
C34108 a_3699_46348# a_4185_45028# 0.001724f
C34109 a_n237_47217# a_1667_45002# 0.002992f
C34110 a_n1151_42308# a_n1059_45260# 0.16984f
C34111 a_3699_46634# a_4099_45572# 4.97e-20
C34112 a_n2661_46634# a_11322_45546# 0.059929f
C34113 a_5807_45002# a_6229_45572# 6.77e-19
C34114 a_16327_47482# a_17568_45572# 9.92e-19
C34115 a_18780_47178# a_18909_45814# 1.24e-20
C34116 a_15567_42826# a_15764_42576# 2.66e-20
C34117 a_5342_30871# a_15803_42450# 0.001339f
C34118 a_22400_42852# a_14097_32519# 3.83e-19
C34119 a_17538_32519# C1_N_btm 1.92e-20
C34120 a_20256_43172# a_20356_42852# 0.001534f
C34121 a_n3674_39304# a_n4334_40480# 1.8e-19
C34122 a_n2293_46634# VDD 1.52629f
C34123 a_375_42282# a_n1557_42282# 0.450989f
C34124 a_10057_43914# a_10405_44172# 0.028414f
C34125 a_n2661_43922# a_n1761_44111# 0.006596f
C34126 a_n2293_43922# a_n2065_43946# 0.02752f
C34127 a_n2661_42834# a_n1899_43946# 0.049432f
C34128 a_8975_43940# a_9672_43914# 4.08e-19
C34129 a_n2956_39768# CLK_DATA 0.015401f
C34130 a_3232_43370# a_2813_43396# 0.05929f
C34131 a_11823_42460# a_12545_42858# 0.039145f
C34132 a_9290_44172# a_14113_42308# 4.21e-20
C34133 a_3537_45260# a_6809_43396# 5.68e-19
C34134 a_n2017_45002# a_12281_43396# 0.028019f
C34135 a_1307_43914# a_1891_43646# 0.00299f
C34136 a_17517_44484# a_18579_44172# 0.031747f
C34137 a_n443_42852# a_8483_43230# 0.001379f
C34138 a_526_44458# a_3823_42558# 0.183187f
C34139 a_n1925_42282# a_3318_42354# 6.66e-20
C34140 a_10903_43370# a_14456_42282# 3.29e-21
C34141 a_1423_45028# a_4699_43561# 1.02e-20
C34142 a_5147_45002# a_5837_43396# 0.009374f
C34143 a_5111_44636# a_5565_43396# 3.27e-19
C34144 a_10193_42453# a_5342_30871# 0.151919f
C34145 a_n1243_44484# a_n4318_39768# 6.55e-21
C34146 a_15227_44166# a_20447_31679# 2.55e-19
C34147 a_1337_46116# a_997_45618# 0.001151f
C34148 a_9290_44172# a_7499_43078# 0.597117f
C34149 a_9625_46129# a_10193_42453# 0.002796f
C34150 a_5937_45572# a_10490_45724# 3.4e-20
C34151 a_8953_45546# a_8746_45002# 0.020026f
C34152 a_4791_45118# a_8783_44734# 6.39e-21
C34153 a_12741_44636# a_15903_45785# 1.65e-19
C34154 a_11415_45002# a_16115_45572# 0.004692f
C34155 a_19123_46287# a_18341_45572# 0.001192f
C34156 a_18285_46348# a_18909_45814# 1.07e-21
C34157 a_10227_46804# a_13720_44458# 0.001314f
C34158 a_n743_46660# a_n2661_43370# 7.86e-20
C34159 a_8199_44636# a_11322_45546# 8.36e-19
C34160 a_8667_46634# a_8953_45002# 8.44e-19
C34161 a_13747_46662# a_17719_45144# 3.9e-20
C34162 a_13661_43548# a_18315_45260# 0.002575f
C34163 a_5807_45002# a_18587_45118# 5.91e-22
C34164 a_526_44458# a_3503_45724# 0.06484f
C34165 a_3877_44458# a_1423_45028# 0.022537f
C34166 a_9823_46155# a_10053_45546# 8.94e-19
C34167 a_8049_45260# a_21167_46155# 3.64e-19
C34168 a_n1151_42308# a_484_44484# 2.43e-19
C34169 a_16327_47482# a_17767_44458# 0.269619f
C34170 a_5342_30871# VDD 0.496295f
C34171 a_15486_42560# a_7174_31319# 1.69e-21
C34172 a_17124_42282# a_17531_42308# 0.003716f
C34173 a_15761_42308# a_4958_30871# 1.41e-19
C34174 a_6123_31319# a_1343_38525# 1.91e-19
C34175 a_3357_43084# a_n784_42308# 4.03e-21
C34176 a_18451_43940# a_15493_43940# 0.051906f
C34177 a_15493_43396# a_11341_43940# 0.020569f
C34178 a_19279_43940# a_2982_43646# 9.07e-21
C34179 a_n4318_40392# a_n4318_38680# 0.023692f
C34180 a_1307_43914# a_4149_42891# 0.006879f
C34181 a_10193_42453# a_20107_42308# 0.007306f
C34182 a_n2956_38216# a_n4334_38304# 6.77e-20
C34183 a_n2017_45002# a_n3674_38680# 2.15e-19
C34184 a_20269_44172# a_20623_43914# 0.001885f
C34185 a_12429_44172# a_12495_44260# 0.012714f
C34186 a_3499_42826# a_3737_43940# 0.002888f
C34187 a_9625_46129# VDD 0.996485f
C34188 a_n1899_43946# a_n1352_43396# 4.29e-19
C34189 a_n1549_44318# a_n1917_43396# 9.82e-19
C34190 a_n1331_43914# a_n1177_43370# 1.74e-19
C34191 a_n1761_44111# a_n447_43370# 0.004447f
C34192 a_n2810_45572# a_n3420_37984# 6.34e-19
C34193 a_19862_44208# a_20935_43940# 0.03846f
C34194 a_14539_43914# a_16823_43084# 0.058282f
C34195 a_768_44030# a_7584_44260# 6.93e-19
C34196 a_20850_46155# a_3357_43084# 5.34e-19
C34197 a_2711_45572# a_13485_45572# 1.99e-20
C34198 a_16388_46812# a_18248_44752# 1.08e-21
C34199 a_20205_31679# a_19963_31679# 9.023429f
C34200 a_11453_44696# a_15493_43940# 5.75e-20
C34201 a_2324_44458# a_5837_45028# 0.003084f
C34202 a_n971_45724# a_n1655_43396# 2.13e-20
C34203 a_11189_46129# a_n2661_43370# 7.55e-21
C34204 a_8049_45260# a_3232_43370# 0.003961f
C34205 a_11652_45724# a_11682_45822# 0.006313f
C34206 a_12427_45724# a_10907_45822# 1.82e-21
C34207 a_10053_45546# a_10306_45572# 0.011897f
C34208 a_10180_45724# a_10216_45572# 0.002048f
C34209 a_n2293_46634# a_5495_43940# 8.7e-21
C34210 a_12741_44636# a_n2661_44458# 0.004092f
C34211 a_7174_31319# C10_N_btm 1.34e-19
C34212 a_n3420_39616# C8_P_btm 0.090298f
C34213 a_n4064_40160# C0_P_btm 3.38e-19
C34214 a_14955_47212# a_5807_45002# 2.52e-20
C34215 a_n3565_39304# a_n1386_35608# 8.05e-20
C34216 a_1209_47178# a_n2661_46098# 2.85e-19
C34217 a_n443_46116# a_n2438_43548# 0.070894f
C34218 a_4915_47217# a_n743_46660# 0.026159f
C34219 a_4958_30871# VIN_N 0.025339f
C34220 a_7754_40130# a_8530_39574# 0.013981f
C34221 a_n1151_42308# a_948_46660# 0.002412f
C34222 a_3160_47472# a_2107_46812# 0.041673f
C34223 a_5815_47464# a_n1925_46634# 5.57e-20
C34224 a_n4064_39616# C10_P_btm 7.64e-19
C34225 VDAC_Pi a_3754_38470# 0.389564f
C34226 a_n2302_37984# a_n2302_37690# 0.050477f
C34227 a_20107_42308# VDD 0.284252f
C34228 a_13487_47204# a_13747_46662# 2.35e-19
C34229 a_13717_47436# a_19321_45002# 1.59e-19
C34230 a_7903_47542# a_n2661_46634# 1.47e-20
C34231 a_n971_45724# a_3524_46660# 0.016598f
C34232 a_n237_47217# a_2959_46660# 8.83e-21
C34233 a_n2497_47436# a_3877_44458# 0.024435f
C34234 a_13258_32519# RST_Z 0.059424f
C34235 a_13507_46334# a_n881_46662# 0.019152f
C34236 a_10227_46804# a_12549_44172# 0.360691f
C34237 a_3626_43646# a_6547_43396# 1.95e-20
C34238 a_3080_42308# a_3457_43396# 1.33e-19
C34239 a_22959_43948# a_22959_43396# 0.025171f
C34240 a_n356_44636# a_1221_42558# 3.42e-19
C34241 a_9159_45572# VDD 0.004886f
C34242 a_14021_43940# a_20556_43646# 0.085306f
C34243 a_n97_42460# a_13667_43396# 2.99e-20
C34244 a_18184_42460# a_17124_42282# 9.36e-20
C34245 a_15493_43940# a_17364_32525# 9.31e-19
C34246 a_3357_43084# a_5691_45260# 0.011637f
C34247 a_13661_43548# a_16867_43762# 6.73e-22
C34248 a_n863_45724# a_n23_44458# 0.056041f
C34249 a_n452_45724# a_n356_44636# 7.27e-21
C34250 a_1823_45246# a_n2661_42282# 3.88e-19
C34251 a_19321_45002# a_19268_43646# 1.56e-20
C34252 a_n2293_46634# a_16137_43396# 4.18e-20
C34253 a_5907_45546# a_4223_44672# 3.43e-21
C34254 a_11136_45572# a_n2661_43370# 5.37e-20
C34255 a_5937_45572# a_6453_43914# 0.144397f
C34256 a_n745_45366# a_n37_45144# 6.85e-19
C34257 a_n1059_45260# a_327_44734# 1.06e-21
C34258 a_n913_45002# a_413_45260# 9.09e-20
C34259 a_20202_43084# a_19862_44208# 0.058613f
C34260 a_10193_42453# a_16237_45028# 0.049386f
C34261 a_10490_45724# a_11691_44458# 2.02e-20
C34262 a_22959_47212# a_20820_30879# 0.004677f
C34263 a_11453_44696# a_12741_44636# 1.02327f
C34264 a_11599_46634# a_3483_46348# 3.49e-19
C34265 a_4915_47217# a_11189_46129# 3.08e-22
C34266 a_6151_47436# a_9823_46155# 0.001307f
C34267 a_12891_46348# a_765_45546# 0.041192f
C34268 a_12549_44172# a_17339_46660# 0.081298f
C34269 a_22731_47423# a_21076_30879# 0.001083f
C34270 a_n2497_47436# a_n1736_46482# 0.005472f
C34271 a_4646_46812# a_6969_46634# 0.072545f
C34272 a_4651_46660# a_6755_46942# 5.05e-21
C34273 a_n1435_47204# a_5164_46348# 1.08e-20
C34274 VIN_N VCM 1.7189f
C34275 VREF VREF_GND 45.064804f
C34276 a_13747_46662# a_14513_46634# 6.82e-19
C34277 a_n1151_42308# a_13925_46122# 4.64e-19
C34278 a_2063_45854# a_2324_44458# 0.028153f
C34279 a_n1741_47186# a_10809_44734# 0.332771f
C34280 a_16237_45028# VDD 0.248452f
C34281 a_743_42282# a_2905_42968# 8.11e-20
C34282 a_18114_32519# C2_N_btm 1.17e-19
C34283 a_n2157_42858# a_n1641_43230# 0.110532f
C34284 a_n1853_43023# a_n1423_42826# 0.022091f
C34285 a_10341_43396# a_21195_42852# 1.4e-20
C34286 a_20193_45348# RST_Z 6.04e-20
C34287 a_16137_43396# a_5342_30871# 1.45e-19
C34288 a_7287_43370# a_7309_42852# 6.34e-20
C34289 a_10180_45724# a_10405_44172# 1.31e-21
C34290 a_n2810_45028# a_n2293_43922# 2.3e-20
C34291 a_21076_30879# a_14209_32519# 0.055087f
C34292 a_3090_45724# a_19339_43156# 2.9e-19
C34293 a_n2956_39768# a_n1630_35242# 0.003986f
C34294 a_3537_45260# a_8333_44734# 1.47e-20
C34295 a_7499_43078# a_10807_43548# 0.119721f
C34296 a_n1613_43370# a_6123_31319# 0.002625f
C34297 a_n2293_42834# a_n2661_44458# 0.0289f
C34298 a_18315_45260# a_18587_45118# 0.13675f
C34299 a_5111_44636# a_7640_43914# 0.001351f
C34300 en_comp a_n2661_42834# 0.080292f
C34301 a_20273_45572# a_11967_42832# 1.95e-21
C34302 a_15415_45028# a_14539_43914# 4.93e-21
C34303 a_1307_43914# a_13720_44458# 1.84e-20
C34304 a_16922_45042# a_18494_42460# 0.242236f
C34305 a_327_44734# a_484_44484# 0.004093f
C34306 a_413_45260# a_556_44484# 2.84e-19
C34307 a_n2438_43548# a_n4318_37592# 1.35e-19
C34308 a_15227_44166# a_17595_43084# 0.041195f
C34309 w_1575_34946# VDAC_Ni 7.89e-19
C34310 a_18597_46090# a_10193_42453# 0.001118f
C34311 a_n2956_39768# a_n2661_45546# 6.28e-20
C34312 a_14084_46812# a_13925_46122# 9.14e-19
C34313 a_14955_47212# a_15143_45578# 2.5e-21
C34314 a_765_45546# a_805_46414# 8.01e-20
C34315 a_11599_46634# a_14495_45572# 3.57e-19
C34316 a_18783_43370# a_18727_42674# 1.92e-19
C34317 a_743_42282# a_15803_42450# 0.037845f
C34318 a_5342_30871# a_n784_42308# 0.049079f
C34319 a_22959_42860# a_22400_42852# 8.07e-19
C34320 a_22223_42860# a_14097_32519# 5.42e-19
C34321 a_9672_43914# VDD 0.150499f
C34322 a_5649_42852# a_14456_42282# 1.31e-19
C34323 a_19700_43370# a_17303_42282# 4.48e-21
C34324 a_4190_30871# a_15890_42674# 2.93e-20
C34325 a_16664_43396# a_4958_30871# 1.61e-19
C34326 a_4520_42826# a_4921_42308# 4.91e-19
C34327 a_3357_43084# a_3080_42308# 0.233522f
C34328 a_n443_42852# a_3935_42891# 5.99e-20
C34329 a_13259_45724# a_21671_42860# 1.9e-20
C34330 a_n967_45348# a_n1177_43370# 0.013627f
C34331 a_18287_44626# a_20362_44736# 5.63e-20
C34332 a_5708_44484# a_n2661_43922# 0.004801f
C34333 a_n1917_44484# a_n1549_44318# 6.05e-19
C34334 a_n1352_44484# a_n1899_43946# 3.68e-19
C34335 a_n1177_44458# a_n1331_43914# 1.54e-19
C34336 a_n452_44636# a_n1761_44111# 4.05e-21
C34337 a_15811_47375# CLK 4.17e-19
C34338 a_18597_46090# VDD 0.930122f
C34339 a_1823_45246# a_3497_42558# 0.002234f
C34340 a_9313_44734# a_15433_44458# 1.54e-20
C34341 a_18989_43940# a_11967_42832# 0.039137f
C34342 a_18780_47178# RST_Z 1.31e-19
C34343 a_8953_45002# a_9165_43940# 4.13e-20
C34344 a_19692_46634# a_20712_42282# 1.06e-20
C34345 a_8696_44636# a_14205_43396# 8.74e-22
C34346 a_18479_47436# START 0.313639f
C34347 a_n357_42282# a_10796_42968# 0.048375f
C34348 a_10193_42453# a_743_42282# 1.1645f
C34349 a_11599_46634# a_17719_45144# 1.93e-21
C34350 a_n1925_42282# a_5066_45546# 3.2e-20
C34351 a_14840_46494# a_13259_45724# 0.002156f
C34352 a_2324_44458# a_14383_46116# 1.41e-19
C34353 a_12549_44172# a_1307_43914# 1.82879f
C34354 a_n971_45724# a_5343_44458# 0.001055f
C34355 a_4185_45028# a_n755_45592# 0.024134f
C34356 a_472_46348# a_n443_42852# 4.66e-19
C34357 a_n743_46660# a_4574_45260# 5.3e-20
C34358 a_n1925_46634# a_5147_45002# 2.49e-20
C34359 a_15368_46634# a_14033_45822# 8.96e-21
C34360 a_11813_46116# a_8696_44636# 4.79e-21
C34361 a_4646_46812# a_3357_43084# 0.024669f
C34362 a_10809_44734# a_10586_45546# 5.07e-19
C34363 a_5807_45002# a_13159_45002# 1.28e-21
C34364 a_13661_43548# a_13017_45260# 6.88e-20
C34365 a_167_45260# a_n356_45724# 9.47e-19
C34366 a_3147_46376# a_2957_45546# 8.73e-20
C34367 a_1123_46634# a_1667_45002# 3.71e-19
C34368 a_2107_46812# a_413_45260# 0.032665f
C34369 a_13059_46348# a_13904_45546# 0.001004f
C34370 a_8128_46384# a_1423_45028# 2.49e-21
C34371 a_14976_45028# a_15037_45618# 0.003888f
C34372 a_3090_45724# a_15225_45822# 7.41e-20
C34373 a_12861_44030# a_19778_44110# 0.113118f
C34374 a_4817_46660# a_2437_43646# 4.02e-20
C34375 a_743_42282# VDD 0.597869f
C34376 a_13678_32519# C5_N_btm 1.22e-19
C34377 a_8325_42308# a_5742_30871# 1.69e-20
C34378 a_9223_42460# a_10533_42308# 4.9e-20
C34379 COMP_P a_21613_42308# 1.34e-20
C34380 a_19778_44110# a_19700_43370# 0.009715f
C34381 a_11827_44484# a_17499_43370# 3.5e-20
C34382 a_n356_44636# a_3626_43646# 0.073377f
C34383 a_19123_46287# VDD 0.336379f
C34384 a_7542_44172# a_7911_44260# 0.00411f
C34385 a_4185_45028# a_22521_40599# 3.39e-20
C34386 a_18285_46348# RST_Z 1.19e-20
C34387 a_18494_42460# a_15743_43084# 0.027791f
C34388 a_18184_42460# a_19268_43646# 1.21e-21
C34389 a_13059_46348# CLK 2.07e-20
C34390 en_comp a_n2293_42282# 0.026f
C34391 a_5343_44458# a_8229_43396# 0.00134f
C34392 a_n1059_45260# a_133_42852# 0.045134f
C34393 a_n357_42282# a_4958_30871# 0.004392f
C34394 a_n913_45002# a_n914_42852# 9.04e-20
C34395 a_n2661_43922# a_n2267_43396# 1.14e-20
C34396 a_n2661_42834# a_n1699_43638# 0.00613f
C34397 a_n2293_43922# a_n2129_43609# 0.028035f
C34398 a_22959_44484# a_22959_43948# 0.026152f
C34399 a_n443_42852# a_15890_42674# 5.07e-21
C34400 a_1307_43914# a_5111_42852# 2.66e-19
C34401 a_16237_45028# a_16137_43396# 5.13e-20
C34402 a_11691_44458# a_16547_43609# 4.26e-20
C34403 a_2711_45572# a_6428_45938# 1.42e-19
C34404 a_13259_45724# a_16115_45572# 0.035684f
C34405 a_16375_45002# a_15903_45785# 0.005324f
C34406 a_5807_45002# a_11967_42832# 3.26e-19
C34407 a_22959_46124# a_20447_31679# 0.015464f
C34408 a_16388_46812# a_16922_45042# 4.23e-21
C34409 a_3483_46348# a_13348_45260# 0.041217f
C34410 a_5937_45572# a_6171_45002# 0.206948f
C34411 a_8953_45546# a_3232_43370# 0.019509f
C34412 a_12549_44172# a_18579_44172# 0.154956f
C34413 a_8049_45260# a_18341_45572# 0.021945f
C34414 a_6419_46155# a_6709_45028# 3.25e-20
C34415 a_13717_47436# a_15811_47375# 1.75e-19
C34416 a_n3420_38528# a_n4064_38528# 8.203589f
C34417 a_n4064_39072# a_n4064_37984# 0.044699f
C34418 a_n3565_38502# a_n2860_38778# 2.96e-19
C34419 a_2112_39137# a_2684_37794# 0.091415f
C34420 a_5755_42308# VDD 0.229304f
C34421 a_5934_30871# C3_N_btm 0.011274f
C34422 a_13487_47204# a_11599_46634# 9.96e-21
C34423 a_12861_44030# a_15507_47210# 2.51e-20
C34424 a_n2109_47186# a_4842_47243# 0.002652f
C34425 a_n1741_47186# a_n881_46662# 0.179671f
C34426 SMPL_ON_P a_n1613_43370# 5.27e-21
C34427 a_1343_38525# a_3754_39964# 3.37e-19
C34428 a_2124_47436# a_2266_47570# 0.007833f
C34429 a_6123_31319# C5_N_btm 0.022099f
C34430 a_4700_47436# a_4883_46098# 1.43e-19
C34431 a_14311_47204# a_14955_47212# 3.11e-20
C34432 a_5932_42308# C10_N_btm 1.34e-19
C34433 a_4958_30871# CAL_N 0.039702f
C34434 a_5495_43940# a_743_42282# 7.52e-22
C34435 a_n2065_43946# a_n901_43156# 6.54e-19
C34436 a_n1549_44318# a_n1853_43023# 7.93e-21
C34437 a_n1761_44111# a_n1641_43230# 2.7e-21
C34438 a_n1331_43914# a_n1991_42858# 3.18e-20
C34439 a_n2956_37592# a_n3690_39616# 1.91e-20
C34440 en_comp a_n3565_39590# 4.23e-19
C34441 a_15493_43396# a_10341_43396# 0.039468f
C34442 a_n2810_45028# a_n3420_39616# 2.09e-19
C34443 a_15493_43940# a_9145_43396# 3.68e-19
C34444 a_2998_44172# a_4361_42308# 9.12e-22
C34445 a_n2433_43396# a_104_43370# 2.99e-21
C34446 a_n1699_43638# a_n1352_43396# 0.051162f
C34447 a_n4318_39304# a_n2012_43396# 1.24e-19
C34448 a_n2129_43609# a_n97_42460# 3.26e-19
C34449 a_2277_45546# VDD 0.209584f
C34450 a_5111_44636# a_7174_31319# 4.88e-21
C34451 a_11967_42832# a_10518_42984# 5.09e-21
C34452 a_14673_44172# a_5534_30871# 1.22e-19
C34453 a_5257_43370# a_5745_43940# 0.005229f
C34454 a_n2438_43548# a_1049_43396# 1.79e-20
C34455 a_13904_45546# a_13556_45296# 4.14e-19
C34456 a_13249_42308# a_9482_43914# 0.061734f
C34457 a_13527_45546# a_13777_45326# 4.75e-19
C34458 a_2324_44458# a_n2661_42834# 0.004585f
C34459 a_n1613_43370# a_6809_43396# 0.001918f
C34460 a_8697_45572# a_6171_45002# 3.24e-19
C34461 a_16327_47482# a_18525_43370# 0.059008f
C34462 a_8049_45260# a_8975_43940# 6.62e-21
C34463 a_3090_45724# a_17973_43940# 0.001042f
C34464 a_20107_45572# a_20841_45814# 0.053479f
C34465 a_21076_30879# a_17730_32519# 0.054832f
C34466 a_n2293_46634# a_3080_42308# 0.039273f
C34467 a_13507_46334# a_17609_46634# 0.01055f
C34468 a_20990_47178# a_15227_44166# 4.31e-19
C34469 a_19386_47436# a_19692_46634# 2.42e-20
C34470 a_10227_46804# a_10861_46660# 0.003218f
C34471 a_n2293_46634# a_4646_46812# 0.135642f
C34472 a_n2497_47436# a_n1641_46494# 0.020605f
C34473 a_13717_47436# a_13059_46348# 5.91e-19
C34474 a_12861_44030# a_15227_46910# 0.050112f
C34475 a_11599_46634# a_14513_46634# 1.15e-20
C34476 C6_P_btm C4_P_btm 0.145942f
C34477 C7_P_btm C3_P_btm 0.136068f
C34478 C9_P_btm C1_P_btm 0.133953f
C34479 C8_P_btm C2_P_btm 0.14124f
C34480 a_n133_46660# a_1057_46660# 2.56e-19
C34481 a_n2438_43548# a_1302_46660# 5.38e-19
C34482 a_n743_46660# a_2162_46660# 3.68e-19
C34483 a_n2661_46634# a_4817_46660# 0.047477f
C34484 a_5807_45002# a_5257_43370# 0.683815f
C34485 EN_VIN_BSTR_N C2_N_btm 0.118072f
C34486 a_n2109_47186# a_n1991_46122# 8.21e-21
C34487 a_n1920_47178# a_n1853_46287# 0.001135f
C34488 a_7903_47542# a_765_45546# 0.001413f
C34489 a_12465_44636# a_14976_45028# 4.97e-20
C34490 a_4883_46098# a_15559_46634# 7.47e-20
C34491 a_19787_47423# a_19466_46812# 1.48e-19
C34492 C10_P_btm C0_P_btm 0.251079f
C34493 a_n881_46662# a_7832_46660# 7.95e-20
C34494 a_n1741_47186# a_n2157_46122# 2.78e-19
C34495 SMPL_ON_P a_n2293_46098# 7.56e-20
C34496 a_22705_37990# VDD 0.085164f
C34497 a_n1925_46634# a_3055_46660# 0.001224f
C34498 a_288_46660# a_n2661_46098# 2.31e-20
C34499 a_2107_46812# a_2609_46660# 0.003525f
C34500 a_1983_46706# a_2443_46660# 2.86e-19
C34501 a_3080_42308# a_5342_30871# 0.01896f
C34502 a_5495_43940# a_5755_42308# 4.04e-22
C34503 a_n2661_42282# a_1184_42692# 9.09e-20
C34504 a_3422_30871# a_15051_42282# 4.65e-20
C34505 a_626_44172# VDD 0.621601f
C34506 a_3626_43646# a_12379_42858# 1.5e-19
C34507 a_2982_43646# a_12545_42858# 9.98e-20
C34508 a_7287_43370# a_7765_42852# 0.002031f
C34509 a_2813_43396# a_2905_42968# 5.2e-19
C34510 a_5244_44056# a_5932_42308# 1.08e-21
C34511 a_n2293_43922# a_n2302_40160# 1.25e-19
C34512 a_11967_42832# a_16197_42308# 1.01e-20
C34513 a_16137_43396# a_743_42282# 0.183525f
C34514 a_15743_43084# a_15940_43402# 0.00103f
C34515 a_17324_43396# a_16823_43084# 0.038999f
C34516 a_17339_46660# a_16977_43638# 3.09e-20
C34517 a_12741_44636# a_9145_43396# 3.38e-20
C34518 a_6171_45002# a_11691_44458# 0.022104f
C34519 a_8696_44636# a_9159_44484# 9.98e-20
C34520 a_n467_45028# a_n2267_44484# 3.24e-21
C34521 a_n357_42282# a_1525_44260# 1.47e-19
C34522 a_n2017_45002# a_n699_43396# 4.86e-20
C34523 a_19692_46634# a_20556_43646# 0.118928f
C34524 a_n967_45348# a_n1177_44458# 0.012502f
C34525 a_413_45260# a_n2661_44458# 0.69469f
C34526 a_n443_42852# a_6453_43914# 4.9e-19
C34527 a_4791_45118# a_6123_31319# 3.81e-20
C34528 a_n2293_46634# a_n1545_46494# 1.01e-19
C34529 a_5275_47026# a_5204_45822# 4.42e-20
C34530 a_3815_47204# a_2711_45572# 3.98e-20
C34531 a_n443_46116# a_603_45572# 0.004683f
C34532 a_n881_46662# a_10586_45546# 1.46e-20
C34533 a_14035_46660# a_13059_46348# 0.072321f
C34534 a_15227_44166# a_20273_46660# 2.91e-19
C34535 a_19333_46634# a_20411_46873# 2.17e-20
C34536 a_14180_46812# a_15227_46910# 3.46e-19
C34537 a_n743_46660# a_10809_44734# 0.032324f
C34538 a_n2312_38680# a_n2956_38680# 6.25577f
C34539 a_n1925_46634# a_n2956_39304# 2.57e-19
C34540 a_7411_46660# a_3483_46348# 2.45e-19
C34541 a_9804_47204# a_9241_46436# 4.41e-20
C34542 a_12359_47026# a_765_45546# 3.39e-21
C34543 a_4883_46098# a_20009_46494# 1.23e-19
C34544 a_11453_44696# a_16375_45002# 0.104273f
C34545 a_19692_46634# a_19551_46910# 0.0536f
C34546 a_19466_46812# a_20107_46660# 1.31e-20
C34547 a_n1151_42308# a_5263_45724# 0.005089f
C34548 a_n971_45724# a_4880_45572# 2.82e-20
C34549 a_2063_45854# a_6667_45809# 0.029741f
C34550 a_n4318_39304# a_n4064_39616# 0.059009f
C34551 a_17730_32519# C0_N_btm 3.27e-20
C34552 a_10835_43094# a_10793_43218# 2.56e-19
C34553 a_8685_43396# a_14456_42282# 4.62e-21
C34554 a_9145_43396# a_5742_30871# 8.14e-20
C34555 a_3626_43646# a_18727_42674# 0.003134f
C34556 a_2982_43646# a_19332_42282# 2.01e-19
C34557 a_3422_30871# C9_N_btm 0.003737f
C34558 a_743_42282# a_n784_42308# 0.087438f
C34559 a_n1059_45260# a_15493_43940# 1.89e-19
C34560 a_n913_45002# a_22223_43948# 3.74e-21
C34561 a_1423_45028# a_5244_44056# 1.01e-20
C34562 a_16922_45042# a_20640_44752# 4.09e-19
C34563 a_18315_45260# a_11967_42832# 3.09e-19
C34564 a_3232_43370# a_9028_43914# 1.62e-19
C34565 a_n443_42852# a_16547_43609# 0.004823f
C34566 a_9838_44484# a_5891_43370# 1.24e-20
C34567 a_n2267_44484# a_n2661_43922# 0.010057f
C34568 a_n2129_44697# a_n2293_43922# 3.05e-19
C34569 a_n1699_44726# a_n2661_42834# 0.002084f
C34570 a_11691_44458# a_14673_44172# 0.371587f
C34571 a_1307_43914# a_7542_44172# 0.022371f
C34572 a_7229_43940# a_6756_44260# 5.36e-21
C34573 a_11827_44484# a_18204_44850# 1.18e-19
C34574 a_22223_45036# a_17517_44484# 1.7e-20
C34575 a_5343_44458# a_9313_44734# 6.56e-21
C34576 w_11334_34010# VDD 1.90683f
C34577 a_15682_46116# a_17583_46090# 0.013015f
C34578 a_n971_45724# a_8560_45348# 0.007243f
C34579 a_6755_46942# a_10193_42453# 0.00109f
C34580 a_10249_46116# a_8746_45002# 1.31e-20
C34581 a_17639_46660# a_16375_45002# 8.23e-20
C34582 a_11309_47204# a_2437_43646# 0.003942f
C34583 a_11189_46129# a_10809_44734# 3.89e-20
C34584 a_4646_46812# a_9159_45572# 1.29e-20
C34585 a_n443_46116# a_2903_45348# 9.86e-20
C34586 a_3090_45724# a_3175_45822# 0.008745f
C34587 a_14976_45028# a_2711_45572# 0.025742f
C34588 a_n743_46660# a_16211_45572# 8.28e-19
C34589 a_11453_44696# a_413_45260# 0.032816f
C34590 a_11599_46634# a_11963_45334# 7.4e-22
C34591 a_9804_47204# a_3357_43084# 8.68e-20
C34592 a_12861_44030# a_9482_43914# 0.021886f
C34593 a_6151_47436# a_1423_45028# 2.69e-21
C34594 a_1823_45246# a_5527_46155# 3.02e-21
C34595 a_3483_46348# a_4365_46436# 3.61e-19
C34596 a_5164_46348# a_526_44458# 2.61e-20
C34597 a_n784_42308# a_5755_42308# 3.86e-20
C34598 a_14635_42282# a_15890_42674# 7.2e-22
C34599 a_2813_43396# VDD 0.004385f
C34600 a_1755_42282# a_2903_42308# 5e-19
C34601 a_2123_42473# a_2713_42308# 6.03e-20
C34602 a_1606_42308# a_3318_42354# 1.73e-19
C34603 a_n913_45002# a_n13_43084# 0.042137f
C34604 a_n2017_45002# a_n4318_38680# 1.48e-19
C34605 a_8667_46634# DATA[4] 3.49e-19
C34606 a_n443_42852# a_n3674_37592# 6.07e-20
C34607 a_6755_46942# VDD 1.05713f
C34608 en_comp a_n1423_42826# 1.04e-20
C34609 a_n967_45348# a_n1991_42858# 0.034664f
C34610 a_n755_45592# a_n39_42308# 7.86e-19
C34611 a_n1761_44111# a_n809_44244# 0.038277f
C34612 a_n2065_43946# a_n984_44318# 0.102325f
C34613 a_n1899_43946# a_n1549_44318# 0.218775f
C34614 a_11823_42460# a_13157_43218# 5.05e-19
C34615 a_3357_43084# a_2075_43172# 8.43e-21
C34616 a_19321_45002# a_18248_44752# 0.004965f
C34617 a_2107_46812# a_2779_44458# 6.26e-21
C34618 a_n2661_45546# a_n906_45572# 6.4e-19
C34619 a_13661_43548# a_18374_44850# 0.00877f
C34620 a_5807_45002# a_18989_43940# 5.17e-20
C34621 a_15682_46116# a_8696_44636# 0.00216f
C34622 a_2324_44458# a_15861_45028# 8.69e-19
C34623 a_17715_44484# a_16855_45546# 0.001764f
C34624 a_12861_44030# a_20159_44458# 0.014378f
C34625 a_8049_45260# a_10193_42453# 0.082788f
C34626 a_n2312_39304# a_n2661_43922# 1.13e-20
C34627 a_n2312_40392# a_n2293_43922# 0.002335f
C34628 a_472_46348# a_2437_43646# 1.19e-20
C34629 a_584_46384# a_n1899_43946# 6.88e-21
C34630 a_n746_45260# a_1414_42308# 3.24e-20
C34631 a_10903_43370# a_14033_45572# 0.003863f
C34632 a_14035_46660# a_13556_45296# 1.33e-21
C34633 a_n2293_46634# a_10057_43914# 0.01757f
C34634 a_n755_45592# a_997_45618# 0.133124f
C34635 a_n863_45724# a_n356_45724# 0.003189f
C34636 a_n4334_40480# a_n4064_39616# 7.84e-19
C34637 a_n4209_39590# a_n4334_39616# 0.25243f
C34638 a_n4315_30879# a_n2302_39866# 9.79e-19
C34639 COMP_P a_n1532_35090# 4.87e-20
C34640 a_n971_45724# a_3785_47178# 0.032234f
C34641 a_n237_47217# a_n1151_42308# 0.63407f
C34642 a_1431_47204# a_584_46384# 0.005844f
C34643 a_n1741_47186# a_n443_46116# 0.053258f
C34644 a_n2109_47186# a_5129_47502# 0.021297f
C34645 a_1209_47178# a_2553_47502# 8.64e-19
C34646 a_1239_47204# a_2063_45854# 3.11e-20
C34647 a_n1630_35242# CAL_P 0.016538f
C34648 a_n4064_40160# a_n2946_39866# 1.91e-19
C34649 a_13720_44458# a_13635_43156# 5.13e-21
C34650 a_n1059_45260# a_5742_30871# 0.002047f
C34651 a_n913_45002# a_11323_42473# 6.5e-19
C34652 a_n2017_45002# a_11551_42558# 0.006777f
C34653 a_3499_42826# a_3539_42460# 0.00342f
C34654 a_n2661_42834# a_n2157_42858# 0.001323f
C34655 a_n2661_43922# a_n2472_42826# 7.7e-20
C34656 a_15493_43396# a_n97_42460# 0.002057f
C34657 a_n356_44636# a_8037_42858# 3.48e-20
C34658 a_375_42282# a_n3674_37592# 0.003119f
C34659 a_8049_45260# VDD 1.89366f
C34660 a_3537_45260# a_7227_42308# 0.001666f
C34661 a_5111_44636# a_5932_42308# 0.021257f
C34662 a_9290_44172# a_9838_44484# 6.21e-19
C34663 a_167_45260# a_n356_44636# 5.64e-19
C34664 a_16680_45572# a_8696_44636# 0.004839f
C34665 a_16855_45546# a_15861_45028# 0.001688f
C34666 a_n2293_46634# a_14021_43940# 0.202404f
C34667 a_5807_45002# a_5745_43940# 3.73e-21
C34668 a_8953_45546# a_8975_43940# 0.02155f
C34669 a_2711_45572# a_2382_45260# 1.81e-20
C34670 a_15765_45572# a_16223_45938# 0.027606f
C34671 a_19692_46634# a_20980_44850# 5.34e-20
C34672 a_n443_42852# a_6171_45002# 2.87e-20
C34673 a_n2661_45546# a_1307_43914# 0.021108f
C34674 a_2063_45854# a_11186_47026# 0.012485f
C34675 a_n971_45724# a_3090_45724# 0.071442f
C34676 a_n1151_42308# a_8270_45546# 0.01803f
C34677 a_6151_47436# a_6682_46987# 0.003543f
C34678 a_n881_46662# a_n743_46660# 0.527182f
C34679 a_n1613_43370# a_n2438_43548# 1.04064f
C34680 a_22521_40599# a_22469_40625# 1.99151f
C34681 a_n3420_38528# VREF_GND 0.047244f
C34682 a_9313_45822# a_8492_46660# 8.95e-19
C34683 a_6545_47178# a_6969_46634# 0.002934f
C34684 a_9863_47436# a_10150_46912# 4.65e-21
C34685 a_n1435_47204# a_8145_46902# 4.03e-21
C34686 a_6491_46660# a_6755_46942# 0.007927f
C34687 a_7754_38470# a_11530_34132# 7.75e-19
C34688 a_n3565_37414# a_n1532_35090# 7.27e-20
C34689 a_n4209_37414# EN_VIN_BSTR_P 0.007584f
C34690 a_11309_47204# a_n2661_46634# 0.042272f
C34691 a_n4064_37984# VDD 1.70621f
C34692 a_n2312_40392# a_n2661_46098# 1.45e-20
C34693 a_n2661_42282# a_5193_42852# 2.87e-21
C34694 a_19479_31679# VDD 0.579914f
C34695 a_19963_31679# C9_N_btm 1.91e-20
C34696 a_21115_43940# a_21195_42852# 2.21e-21
C34697 a_15493_43940# a_19987_42826# 7.44e-20
C34698 a_11341_43940# a_21356_42826# 4.25e-20
C34699 a_10695_43548# a_10341_43396# 0.008043f
C34700 a_n2293_43922# a_8791_42308# 8.6e-20
C34701 a_9313_44734# a_12563_42308# 2.09e-20
C34702 a_2437_43646# START 0.12936f
C34703 a_14021_43940# a_5342_30871# 0.001922f
C34704 a_9145_43396# a_10849_43646# 0.003354f
C34705 a_14579_43548# a_14955_43396# 4.82e-20
C34706 a_8685_43396# a_10149_43396# 7.5e-19
C34707 a_22223_45572# RST_Z 7.78e-20
C34708 a_n2840_43370# a_n3674_39304# 0.008407f
C34709 a_n1917_43396# a_n1991_42858# 1.29e-19
C34710 a_n2267_43396# a_n1641_43230# 0.00175f
C34711 a_n1352_43396# a_n2157_42858# 5.11e-19
C34712 a_n1177_43370# a_n1853_43023# 1.6e-19
C34713 a_n1699_43638# a_n1423_42826# 5.89e-19
C34714 a_n2129_43609# a_n901_43156# 0.001317f
C34715 a_3080_42308# a_743_42282# 0.069641f
C34716 a_20447_31679# C7_N_btm 7.54e-20
C34717 a_10903_43370# a_10555_44260# 0.011277f
C34718 a_21076_30879# a_17538_32519# 0.054805f
C34719 a_6511_45714# a_n2661_43922# 6.22e-21
C34720 a_n443_42852# a_14673_44172# 1.12e-19
C34721 a_9049_44484# a_7640_43914# 7.12e-20
C34722 a_4646_46812# a_743_42282# 3.55e-19
C34723 a_12891_46348# a_13460_43230# 1.83e-20
C34724 a_12549_44172# a_13635_43156# 2.09e-20
C34725 a_13017_45260# a_13159_45002# 0.160415f
C34726 a_11787_45002# a_9482_43914# 8.24e-21
C34727 a_2711_45572# a_15433_44458# 2.54e-20
C34728 a_5111_44636# a_1423_45028# 0.028542f
C34729 a_526_44458# a_3499_42826# 0.089844f
C34730 a_n143_45144# a_45_45144# 7.47e-21
C34731 a_10809_44734# a_11750_44172# 6e-21
C34732 a_18909_45814# a_11691_44458# 7.74e-19
C34733 a_18691_45572# a_19113_45348# 0.001513f
C34734 a_n1059_45260# a_n2293_42834# 0.035031f
C34735 w_11334_34010# a_n784_42308# 0.001604f
C34736 SMPL_ON_P a_n1736_42282# 5.11e-20
C34737 a_6755_46942# a_16137_43396# 1.16e-19
C34738 a_8034_45724# a_7542_44172# 7e-22
C34739 a_3065_45002# a_3602_45348# 5.93e-19
C34740 a_3429_45260# a_3495_45348# 0.010598f
C34741 a_7499_43078# a_8375_44464# 2.35e-19
C34742 a_8568_45546# a_5891_43370# 4.55e-19
C34743 a_5205_44484# a_1307_43914# 0.006798f
C34744 w_1575_34946# a_5742_30871# 0.032598f
C34745 a_4817_46660# a_765_45546# 0.010165f
C34746 a_6755_46942# a_10185_46660# 3.5e-19
C34747 a_n881_46662# a_11189_46129# 2.91e-19
C34748 a_11453_44696# a_18985_46122# 9.23e-20
C34749 a_13507_46334# a_22223_46124# 0.024274f
C34750 a_21496_47436# a_6945_45028# 0.001335f
C34751 a_21177_47436# a_10809_44734# 0.009997f
C34752 a_n1021_46688# a_n1853_46287# 2.81e-20
C34753 a_n2438_43548# a_n2293_46098# 0.409291f
C34754 a_n1925_46634# a_n1991_46122# 0.008581f
C34755 a_n2293_46634# a_n901_46420# 3.18e-20
C34756 a_n2661_46634# a_472_46348# 1.17e-20
C34757 a_10428_46928# a_10933_46660# 2.28e-19
C34758 a_10249_46116# a_10425_46660# 3.17e-19
C34759 a_9804_47204# a_9625_46129# 0.037672f
C34760 a_11735_46660# a_11901_46660# 0.579036f
C34761 a_8128_46384# a_9569_46155# 3.31e-20
C34762 a_13661_43548# a_3483_46348# 0.381471f
C34763 a_6575_47204# a_8034_45724# 2.35e-20
C34764 a_4883_46098# a_21137_46414# 0.010468f
C34765 a_14021_43940# a_20107_42308# 2.15e-20
C34766 a_n97_42460# a_8791_42308# 4.89e-19
C34767 a_4905_42826# a_5421_42558# 0.002476f
C34768 a_6293_42852# a_1755_42282# 1.75e-19
C34769 a_5289_44734# VDD 5.21e-19
C34770 a_3422_30871# a_n3420_37440# 0.0344f
C34771 a_n2157_42858# a_n2293_42282# 5.22e-20
C34772 a_3539_42460# a_3318_42354# 0.161793f
C34773 a_3626_43646# a_3823_42558# 0.017529f
C34774 a_2982_43646# a_5379_42460# 0.068435f
C34775 a_16137_43396# a_16328_43172# 5.93e-19
C34776 a_8952_43230# a_10796_42968# 2e-20
C34777 a_10083_42826# a_10835_43094# 0.043619f
C34778 a_13259_45724# a_13667_43396# 0.160676f
C34779 a_18587_45118# a_18374_44850# 9.02e-19
C34780 a_n2661_43370# a_5891_43370# 3.67e-19
C34781 a_11827_44484# a_15004_44636# 0.007895f
C34782 a_19778_44110# a_18287_44626# 5.65e-21
C34783 a_413_45260# a_19237_31679# 0.119197f
C34784 a_3357_43084# a_5013_44260# 2.89e-19
C34785 a_4185_45028# a_10083_42826# 3.49e-20
C34786 a_20202_43084# a_21671_42860# 0.002893f
C34787 a_n2661_44458# a_2779_44458# 0.011596f
C34788 a_n967_45348# a_n1331_43914# 0.003919f
C34789 a_n2293_45010# a_453_43940# 0.181603f
C34790 a_n2661_45010# a_2479_44172# 7.5e-19
C34791 SMPL_ON_P a_n4209_37414# 8.3e-19
C34792 a_n443_42852# a_766_43646# 8.62e-19
C34793 a_n1059_45260# a_1115_44172# 2.41e-21
C34794 a_n2312_40392# a_n3420_39616# 6.3e-21
C34795 a_14537_43396# a_16241_44484# 0.003767f
C34796 a_n1699_44726# a_n1352_44484# 0.051162f
C34797 a_11691_44458# a_12607_44458# 0.042423f
C34798 w_1575_34946# C0_dummy_P_btm 3.87e-21
C34799 a_12741_44636# a_13925_46122# 7.71e-21
C34800 a_n971_45724# a_2274_45254# 0.002827f
C34801 a_6545_47178# a_3357_43084# 0.005247f
C34802 a_n743_46660# a_8162_45546# 2.28e-21
C34803 a_13747_46662# a_13249_42308# 0.134714f
C34804 a_11415_45002# a_15015_46420# 4.21e-20
C34805 a_n2109_47186# a_4558_45348# 5.21e-20
C34806 a_n2497_47436# a_5111_44636# 8.27e-21
C34807 a_21188_46660# a_21137_46414# 4.35e-19
C34808 a_21363_46634# a_6945_45028# 1.28e-19
C34809 a_20841_46902# a_10809_44734# 0.006187f
C34810 a_7227_47204# a_2437_43646# 0.006315f
C34811 a_12861_44030# a_20623_45572# 7.98e-22
C34812 a_18597_46090# a_18479_45785# 0.009071f
C34813 a_2107_46812# a_2211_45572# 3.18e-20
C34814 a_n1925_46634# a_7499_43078# 9.19e-20
C34815 a_n2661_46634# a_10490_45724# 0.01771f
C34816 a_1823_45246# a_6165_46155# 3.85e-21
C34817 a_3483_46348# a_4185_45028# 0.430982f
C34818 a_n746_45260# a_1667_45002# 2.7e-22
C34819 a_n1151_42308# a_n2017_45002# 0.058036f
C34820 a_16327_47482# a_17034_45572# 0.002231f
C34821 a_5257_43370# a_n755_45592# 2.64e-20
C34822 a_5807_45002# a_15143_45578# 3.06e-21
C34823 a_18780_47178# a_18341_45572# 1.16e-20
C34824 a_15567_42826# a_15486_42560# 1.56e-19
C34825 a_5342_30871# a_15764_42576# 0.002004f
C34826 a_5837_42852# a_5379_42460# 4.94e-19
C34827 a_17538_32519# C0_N_btm 1.63e-20
C34828 a_20256_43172# a_20256_42852# 9.31e-19
C34829 a_5837_43172# a_5932_42308# 3.37e-21
C34830 a_15037_43940# VDD 0.190221f
C34831 a_5147_45002# a_5565_43396# 2.01e-22
C34832 a_n2442_46660# VDD 0.693209f
C34833 a_10440_44484# a_10405_44172# 0.001304f
C34834 a_n2293_43922# a_n2472_43914# 0.189122f
C34835 a_n2661_43922# a_n2065_43946# 0.013023f
C34836 a_n2661_42834# a_n1761_44111# 0.073205f
C34837 a_8975_43940# a_9028_43914# 0.184602f
C34838 a_10057_43914# a_9672_43914# 0.143523f
C34839 a_n2840_46634# CLK_DATA 9e-19
C34840 a_11823_42460# a_12089_42308# 0.335983f
C34841 a_18479_45785# a_743_42282# 7.51e-20
C34842 a_9290_44172# a_13657_42558# 4.35e-20
C34843 a_3537_45260# a_6643_43396# 0.001481f
C34844 a_21076_30879# a_22465_38105# 6.77e-19
C34845 a_1307_43914# a_1427_43646# 2.4e-19
C34846 a_7705_45326# a_7287_43370# 9.03e-21
C34847 a_n443_42852# a_8292_43218# 0.002007f
C34848 a_526_44458# a_3318_42354# 3.31e-19
C34849 a_n1925_42282# a_2903_42308# 1.31e-19
C34850 a_10903_43370# a_13575_42558# 8.65e-20
C34851 a_19006_44850# a_11967_42832# 0.013801f
C34852 a_n1151_42308# a_n89_44484# 0.007033f
C34853 a_6151_47436# a_6109_44484# 1.83e-20
C34854 a_16327_47482# a_16979_44734# 4.27e-19
C34855 a_1337_46116# a_n755_45592# 8.94e-20
C34856 a_8199_44636# a_10490_45724# 0.019372f
C34857 a_5937_45572# a_8746_45002# 0.121678f
C34858 a_9625_46129# a_10180_45724# 0.00231f
C34859 a_8953_45546# a_10193_42453# 6e-19
C34860 a_768_44030# a_11827_44484# 0.831344f
C34861 a_12549_44172# a_22223_45036# 8.25e-20
C34862 a_4791_45118# a_8333_44734# 4.95e-19
C34863 a_12741_44636# a_15599_45572# 3.13e-19
C34864 a_11415_45002# a_16333_45814# 0.00197f
C34865 a_18285_46348# a_18341_45572# 2.47e-21
C34866 a_19123_46287# a_18479_45785# 3.74e-20
C34867 a_10227_46804# a_13076_44458# 1.5e-19
C34868 a_11599_46634# a_18443_44721# 1.76e-20
C34869 a_8049_45260# a_20850_46155# 3.79e-19
C34870 a_13747_46662# a_17613_45144# 1.85e-20
C34871 a_5807_45002# a_18315_45260# 5.54e-21
C34872 a_13661_43548# a_17719_45144# 2.08e-20
C34873 a_526_44458# a_3316_45546# 0.128261f
C34874 a_2324_44458# a_3775_45552# 6.98e-21
C34875 a_n1021_46688# a_n2661_43370# 1.67e-22
C34876 a_19321_45002# a_16922_45042# 0.493823f
C34877 a_4883_46098# a_6298_44484# 9.77e-21
C34878 a_19692_46634# a_3357_43084# 0.046179f
C34879 a_15051_42282# a_7174_31319# 6.09e-20
C34880 a_n3674_37592# a_n3420_37984# 0.172946f
C34881 a_17124_42282# a_17303_42282# 0.172579f
C34882 a_15521_42308# a_4958_30871# 1.44e-19
C34883 a_5934_30871# a_1736_39587# 8.81e-20
C34884 a_15279_43071# VDD 0.189193f
C34885 a_n784_42308# a_n4064_37984# 0.00652f
C34886 a_n1630_35242# a_n3565_38216# 1.42e-19
C34887 a_5742_30871# a_n4315_30879# 9.24e-21
C34888 a_5534_30871# RST_Z 0.031803f
C34889 a_n2810_45572# a_n3690_38304# 4.13e-19
C34890 a_18326_43940# a_15493_43940# 0.075033f
C34891 a_19328_44172# a_11341_43940# 0.004787f
C34892 a_n4318_40392# a_n3674_39304# 0.024125f
C34893 a_1307_43914# a_3863_42891# 0.005265f
C34894 a_10193_42453# a_13258_32519# 0.061618f
C34895 a_n2956_38216# a_n4209_38216# 0.232905f
C34896 a_n2017_45002# a_n2840_42282# 7.53e-19
C34897 a_5883_43914# a_4361_42308# 2.27e-20
C34898 a_n2267_44484# a_n1641_43230# 7.05e-22
C34899 a_n2129_44697# a_n901_43156# 3.52e-20
C34900 a_20269_44172# a_20365_43914# 0.419086f
C34901 en_comp a_14097_32519# 5.98e-20
C34902 a_20447_31679# COMP_P 4.66e-20
C34903 a_10949_43914# a_12710_44260# 0.001055f
C34904 a_8953_45546# VDD 1.32809f
C34905 a_19862_44208# a_20623_43914# 0.023134f
C34906 a_14539_43914# a_17021_43396# 5.66e-19
C34907 a_10057_43914# a_743_42282# 4.3e-20
C34908 a_n1761_44111# a_n1352_43396# 1.05e-20
C34909 a_n984_44318# a_n2129_43609# 5.84e-20
C34910 a_n1899_43946# a_n1177_43370# 0.001333f
C34911 a_n2293_46634# a_5013_44260# 3.03e-20
C34912 a_21076_30879# a_19721_31679# 0.05488f
C34913 a_768_44030# a_6756_44260# 3.81e-19
C34914 a_11525_45546# a_11682_45822# 0.18824f
C34915 a_2711_45572# a_13385_45572# 6.27e-20
C34916 SMPL_ON_N a_15493_43940# 1.94e-20
C34917 a_10227_46804# a_15301_44260# 2.48e-19
C34918 w_11334_34010# a_3080_42308# 0.001073f
C34919 a_n971_45724# a_n1821_43396# 2.41e-20
C34920 a_9290_44172# a_n2661_43370# 0.185465f
C34921 a_3090_45724# a_9313_44734# 2.43867f
C34922 a_16375_45002# a_n1059_45260# 0.001787f
C34923 a_11962_45724# a_10907_45822# 2.36e-20
C34924 a_10053_45546# a_10216_45572# 0.011381f
C34925 a_18597_46090# a_14021_43940# 0.0185f
C34926 a_7174_31319# C9_N_btm 9.33e-20
C34927 a_n3420_39616# C9_P_btm 7.08e-19
C34928 a_n4064_40160# C1_P_btm 1.21e-19
C34929 a_15507_47210# a_16697_47582# 2.56e-19
C34930 a_n3565_39304# a_n1838_35608# 1.81e-19
C34931 a_4958_30871# VIN_P 0.025339f
C34932 a_1209_47178# a_1799_45572# 1.57e-19
C34933 a_327_47204# a_n2661_46098# 2.08e-20
C34934 a_n443_46116# a_n743_46660# 0.532861f
C34935 a_7754_40130# a_7754_38470# 0.111791f
C34936 a_7754_39964# a_3754_38470# 0.081868f
C34937 a_n3565_39590# C7_P_btm 0.00198f
C34938 a_16023_47582# a_16119_47582# 0.013793f
C34939 a_14311_47204# a_5807_45002# 3.38e-19
C34940 a_n1151_42308# a_1123_46634# 0.002563f
C34941 a_2905_45572# a_2107_46812# 0.031826f
C34942 a_7754_39300# a_7754_38968# 0.296258f
C34943 a_n4064_37984# a_n2302_37690# 2.59e-20
C34944 a_n2302_37984# a_n4064_37440# 2.59e-20
C34945 a_13258_32519# VDD 3.19231f
C34946 a_7227_47204# a_n2661_46634# 1.7e-19
C34947 a_12861_44030# a_13747_46662# 0.139424f
C34948 a_n971_45724# a_3699_46634# 0.024384f
C34949 a_n4209_39304# a_n1532_35090# 1.52e-19
C34950 a_19647_42308# RST_Z 4.07e-20
C34951 a_17591_47464# a_12549_44172# 0.001606f
C34952 a_10227_46804# a_12891_46348# 0.058451f
C34953 a_n4209_39590# C5_P_btm 5.07e-20
C34954 a_548_43396# a_648_43396# 0.005294f
C34955 a_4699_43561# a_3457_43396# 9.15e-20
C34956 a_2982_43646# a_7287_43370# 6.68e-21
C34957 a_3080_42308# a_2813_43396# 9.02e-20
C34958 a_15493_43940# a_22959_43396# 3.06e-19
C34959 a_3539_42460# a_6197_43396# 4.71e-21
C34960 a_n356_44636# a_1149_42558# 2.72e-19
C34961 a_14673_44172# a_14635_42282# 0.002024f
C34962 a_11967_42832# a_10793_43218# 1.94e-21
C34963 a_14021_43940# a_743_42282# 0.002697f
C34964 a_5343_44458# a_8515_42308# 9e-19
C34965 a_n1761_44111# a_n2293_42282# 8.68e-20
C34966 a_22223_43948# a_17364_32525# 6.31e-19
C34967 a_10193_42453# a_20193_45348# 0.305022f
C34968 a_8746_45002# a_11691_44458# 4.34e-20
C34969 a_11415_45002# a_15493_43396# 1.63e-20
C34970 a_n443_42852# a_12607_44458# 4.46e-20
C34971 a_n863_45724# a_n356_44636# 0.301674f
C34972 a_3877_44458# a_3457_43396# 3.97e-22
C34973 a_19321_45002# a_15743_43084# 6.69e-20
C34974 a_n2312_40392# a_n901_43156# 1.65e-20
C34975 a_5263_45724# a_4223_44672# 7.35e-19
C34976 a_4099_45572# a_n699_43396# 9.59e-21
C34977 a_2711_45572# a_5343_44458# 3.61e-20
C34978 a_5937_45572# a_5663_43940# 0.177912f
C34979 a_1138_42852# a_n2661_42282# 1.46e-20
C34980 a_n745_45366# a_n143_45144# 8.24e-19
C34981 a_n1059_45260# a_413_45260# 1.08e-19
C34982 a_11453_44696# a_20820_30879# 0.002153f
C34983 SMPL_ON_N a_12741_44636# 8.39e-20
C34984 a_5429_46660# a_5257_43370# 2.57e-20
C34985 a_4915_47217# a_9290_44172# 0.002979f
C34986 a_12549_44172# a_15312_46660# 5.76e-20
C34987 a_11309_47204# a_765_45546# 0.03506f
C34988 a_n2497_47436# a_n2956_38680# 2.47e-20
C34989 a_4646_46812# a_6755_46942# 0.362783f
C34990 a_3877_44458# a_6969_46634# 0.101189f
C34991 a_6151_47436# a_9569_46155# 2.49e-19
C34992 a_6575_47204# a_8016_46348# 5.51e-20
C34993 a_n1435_47204# a_5068_46348# 3.74e-21
C34994 VIN_P VCM 1.7189f
C34995 VIN_N VREF_GND 16.4969f
C34996 a_13747_46662# a_14180_46812# 0.021289f
C34997 a_n2661_46634# a_12156_46660# 0.009815f
C34998 a_584_46384# a_2324_44458# 2.7e-19
C34999 a_n1151_42308# a_13759_46122# 2.36e-19
C35000 a_22223_47212# a_21076_30879# 7.91e-19
C35001 a_16137_43396# a_15279_43071# 2.14e-19
C35002 a_20193_45348# VDD 0.793111f
C35003 a_18114_32519# C1_N_btm 1.21e-19
C35004 a_n1853_43023# a_n1991_42858# 0.237526f
C35005 a_n2157_42858# a_n1423_42826# 0.07009f
C35006 a_10341_43396# a_21356_42826# 8.92e-20
C35007 a_16922_45042# a_18184_42460# 0.028064f
C35008 a_10180_45724# a_9672_43914# 9.13e-20
C35009 a_10227_46804# a_15720_42674# 1.7e-19
C35010 a_7499_43078# a_10949_43914# 0.152939f
C35011 a_19431_45546# a_18579_44172# 2.71e-21
C35012 a_20820_30879# a_17364_32525# 0.055604f
C35013 a_526_44458# a_6197_43396# 5.62e-19
C35014 a_n1613_43370# a_7227_42308# 0.001156f
C35015 a_5111_44636# a_6109_44484# 0.003573f
C35016 a_3537_45260# a_8238_44734# 0.001272f
C35017 a_20107_45572# a_11967_42832# 6.49e-21
C35018 a_14797_45144# a_14539_43914# 1.54e-19
C35019 a_n357_42282# a_5829_43940# 3.11e-19
C35020 a_2324_44458# a_15095_43370# 5.95e-19
C35021 a_n2442_46660# a_n784_42308# 3.54e-19
C35022 a_15227_44166# a_16795_42852# 3.87e-19
C35023 a_10227_46804# a_11322_45546# 6.46e-22
C35024 a_13661_43548# a_n357_42282# 2.24e-19
C35025 a_n2956_39768# a_n2810_45572# 0.043168f
C35026 a_n2840_46634# a_n2661_45546# 6.53e-19
C35027 a_14084_46812# a_13759_46122# 0.001243f
C35028 a_11901_46660# a_2324_44458# 9.43e-21
C35029 a_9313_45822# a_9241_45822# 7.24e-19
C35030 a_16327_47482# a_11823_42460# 1.03e-20
C35031 a_15368_46634# a_10903_43370# 4.05e-21
C35032 a_765_45546# a_472_46348# 6.08e-19
C35033 a_4646_46812# a_8049_45260# 0.001749f
C35034 a_11599_46634# a_13249_42308# 4.64e-20
C35035 a_743_42282# a_15764_42576# 0.054445f
C35036 a_22223_42860# a_22400_42852# 0.154104f
C35037 a_22165_42308# a_14097_32519# 1.3e-19
C35038 a_9028_43914# VDD 0.17194f
C35039 a_5649_42852# a_13575_42558# 6.94e-20
C35040 a_4190_30871# a_15959_42545# 6.15e-20
C35041 a_20922_43172# a_20753_42852# 0.08213f
C35042 a_15743_43084# a_17531_42308# 2.2e-21
C35043 a_19268_43646# a_17303_42282# 2.14e-21
C35044 a_n2661_44458# a_644_44056# 6.99e-20
C35045 a_3357_43084# a_4699_43561# 0.002313f
C35046 a_n443_42852# a_3681_42891# 1.37e-20
C35047 a_10193_42453# a_20301_43646# 2.72e-19
C35048 a_13259_45724# a_21195_42852# 1.73e-20
C35049 a_18143_47464# START 0.006044f
C35050 a_n967_45348# a_n1917_43396# 9.47e-19
C35051 a_18287_44626# a_20159_44458# 5.37e-21
C35052 a_18248_44752# a_20362_44736# 2.99e-20
C35053 a_5608_44484# a_n2661_43922# 0.001386f
C35054 a_n1352_44484# a_n1761_44111# 1.85e-21
C35055 a_n1177_44458# a_n1899_43946# 7.1e-19
C35056 a_n2129_44697# a_n984_44318# 1.03e-20
C35057 a_10227_46804# SINGLE_ENDED 1.93e-19
C35058 a_1823_45246# a_5379_42460# 1.01e-20
C35059 a_9313_44734# a_14815_43914# 1.48e-20
C35060 a_18374_44850# a_11967_42832# 0.053726f
C35061 a_18989_43940# a_19006_44850# 0.168452f
C35062 a_n913_45002# a_104_43370# 2.19e-20
C35063 a_n2017_45002# a_n1809_43762# 0.003534f
C35064 a_n2661_43370# a_10807_43548# 7.36e-20
C35065 a_15507_47210# CLK 6.68e-19
C35066 a_18479_47436# RST_Z 1.77e-19
C35067 a_18780_47178# VDD 0.245515f
C35068 a_n357_42282# a_10835_43094# 0.02434f
C35069 a_10227_46804# a_15060_45348# 3.31e-19
C35070 a_11599_46634# a_17613_45144# 4.99e-21
C35071 a_526_44458# a_5066_45546# 0.009401f
C35072 a_15015_46420# a_13259_45724# 0.001291f
C35073 a_12891_46348# a_1307_43914# 0.008663f
C35074 a_12549_44172# a_16019_45002# 8.08e-21
C35075 a_3699_46348# a_n755_45592# 0.003336f
C35076 a_472_46348# a_509_45822# 2.66e-19
C35077 a_376_46348# a_n443_42852# 7.22e-19
C35078 a_4185_45028# a_n357_42282# 0.023019f
C35079 a_n743_46660# a_3537_45260# 4.3e-20
C35080 a_3877_44458# a_3357_43084# 0.02473f
C35081 a_5807_45002# a_13017_45260# 4.58e-19
C35082 a_167_45260# a_3503_45724# 1.15e-19
C35083 a_2804_46116# a_2957_45546# 0.009196f
C35084 a_n746_45260# a_n699_43396# 0.002245f
C35085 a_n237_47217# a_4223_44672# 2.68e-21
C35086 a_13059_46348# a_13527_45546# 0.017655f
C35087 a_3090_45724# a_15037_45618# 8.98e-19
C35088 a_4955_46873# a_2437_43646# 1.65e-19
C35089 a_12861_44030# a_18911_45144# 0.169f
C35090 a_n2661_46634# a_6171_45002# 0.042529f
C35091 a_13678_32519# C4_N_btm 1.42e-19
C35092 a_5342_30871# a_n4064_37440# 0.028573f
C35093 a_20301_43646# VDD 0.296691f
C35094 a_9803_42558# a_9885_42558# 0.171361f
C35095 a_13467_32519# C7_N_btm 1.83e-20
C35096 a_n784_42308# a_13258_32519# 0.140549f
C35097 a_4190_30871# RST_Z 0.087843f
C35098 a_13887_32519# C1_N_btm 8.65e-20
C35099 a_9482_43914# a_9127_43156# 4.2e-19
C35100 a_18285_46348# VDD 0.259614f
C35101 a_7542_44172# a_7584_44260# 0.009099f
C35102 a_4185_45028# CAL_N 0.002972f
C35103 a_18184_42460# a_15743_43084# 0.182123f
C35104 a_18494_42460# a_18783_43370# 4.06e-21
C35105 en_comp a_22959_42860# 1.14e-21
C35106 a_n2956_37592# a_n2293_42282# 1.77e-20
C35107 a_n2017_45002# a_133_42852# 0.001378f
C35108 a_n1059_45260# a_n914_42852# 6.52e-20
C35109 a_n2293_43922# a_n2433_43396# 0.028793f
C35110 a_n2661_42834# a_n2267_43396# 0.014077f
C35111 a_n2661_43922# a_n2129_43609# 1.04e-20
C35112 a_20820_30879# a_21589_35634# 5.09e-20
C35113 a_17730_32519# a_22959_43948# 0.00961f
C35114 a_22959_44484# a_15493_43940# 3.35e-19
C35115 a_n443_42852# a_15959_42545# 1.56e-19
C35116 a_1307_43914# a_4520_42826# 6.56e-19
C35117 a_11691_44458# a_16243_43396# 4.28e-20
C35118 a_2711_45572# a_4880_45572# 0.006167f
C35119 a_13259_45724# a_16333_45814# 0.02201f
C35120 a_16375_45002# a_15599_45572# 1.1e-19
C35121 a_13661_43548# a_18588_44850# 0.005669f
C35122 a_10809_44734# a_20447_31679# 0.005556f
C35123 a_3483_46348# a_13159_45002# 0.017316f
C35124 a_5937_45572# a_3232_43370# 0.662525f
C35125 a_8199_44636# a_6171_45002# 0.163434f
C35126 a_22959_46124# a_22959_45572# 0.025171f
C35127 a_15227_44166# a_17801_45144# 8.12e-20
C35128 a_8049_45260# a_18479_45785# 0.0037f
C35129 a_8270_45546# a_4223_44672# 1.84e-19
C35130 a_13925_46122# a_413_45260# 9.96e-21
C35131 a_6598_45938# a_7227_45028# 1.78e-20
C35132 a_n3420_38528# a_n2946_38778# 0.236674f
C35133 a_2112_39137# a_1177_38525# 3.38e-19
C35134 a_n3690_38528# a_n4064_38528# 0.085414f
C35135 a_n3565_38502# a_n2302_38778# 0.044367f
C35136 a_n4209_38502# a_n2216_38778# 0.001361f
C35137 a_5421_42558# VDD 0.007373f
C35138 a_5934_30871# C2_N_btm 0.011047f
C35139 a_7174_31319# a_n3420_37440# 0.002179f
C35140 a_13717_47436# a_15507_47210# 2.86e-19
C35141 a_12861_44030# a_11599_46634# 0.169929f
C35142 a_n1741_47186# a_n1613_43370# 0.018791f
C35143 a_n971_45724# a_2583_47243# 0.006608f
C35144 a_n785_47204# a_7_47243# 7.85e-19
C35145 a_1209_47178# a_2747_46873# 2.14e-19
C35146 a_6123_31319# C4_N_btm 0.132906f
C35147 a_5932_42308# C9_N_btm 9.33e-20
C35148 a_4958_30871# a_11206_38545# 1.83e-20
C35149 a_5013_44260# a_743_42282# 1.7e-20
C35150 a_n2065_43946# a_n1641_43230# 6.4e-21
C35151 a_n1899_43946# a_n1991_42858# 6.45e-19
C35152 a_n1549_44318# a_n2157_42858# 2.53e-21
C35153 a_n1331_43914# a_n1853_43023# 6.71e-22
C35154 a_n2956_37592# a_n3565_39590# 0.023811f
C35155 a_n2267_43396# a_n1352_43396# 0.124988f
C35156 a_n2129_43609# a_n447_43370# 0.119518f
C35157 a_1609_45822# VDD 0.270106f
C35158 a_14673_44172# a_14543_43071# 2.46e-19
C35159 a_n2438_43548# a_1209_43370# 8.21e-21
C35160 a_13904_45546# a_9482_43914# 0.002673f
C35161 a_13527_45546# a_13556_45296# 0.006724f
C35162 a_13759_46122# a_13857_44734# 2.43e-22
C35163 a_13249_42308# a_13348_45260# 3.41e-20
C35164 a_11823_42460# a_14537_43396# 0.001649f
C35165 a_n1613_43370# a_6643_43396# 2.72e-19
C35166 a_8192_45572# a_6171_45002# 0.00429f
C35167 a_3483_46348# a_11967_42832# 0.264293f
C35168 a_16327_47482# a_18429_43548# 0.057366f
C35169 a_20820_30879# a_19237_31679# 0.053048f
C35170 a_n2497_47436# a_791_42968# 2.18e-21
C35171 a_11322_45546# a_1307_43914# 3.56e-20
C35172 a_8049_45260# a_10057_43914# 5.59e-20
C35173 a_2711_45572# a_8560_45348# 0.002436f
C35174 a_10227_46804# a_16409_43396# 6.95e-19
C35175 a_3090_45724# a_17737_43940# 3.24e-20
C35176 a_20107_45572# a_20273_45572# 0.667378f
C35177 a_768_44030# a_8147_43396# 2.39e-22
C35178 a_n2442_46660# a_3080_42308# 4.94e-21
C35179 a_n2956_39768# a_n1557_42282# 2.12e-20
C35180 a_n2293_46634# a_4699_43561# 0.006722f
C35181 a_9049_44484# a_1423_45028# 0.024539f
C35182 a_6755_46942# a_14021_43940# 2.04e-19
C35183 C10_P_btm C1_P_btm 0.204172f
C35184 a_13507_46334# a_16292_46812# 3.92e-19
C35185 a_20894_47436# a_15227_44166# 9.3e-22
C35186 a_18597_46090# a_19692_46634# 0.019861f
C35187 a_10227_46804# a_12359_47026# 0.012196f
C35188 a_19386_47436# a_19466_46812# 2.89e-19
C35189 a_15811_47375# a_13885_46660# 0.0013f
C35190 a_1983_46706# a_n2661_46098# 0.147223f
C35191 a_n2293_46634# a_3877_44458# 1.3e-21
C35192 a_n2497_47436# a_n1423_46090# 0.008067f
C35193 a_9804_47204# a_6755_46942# 0.028571f
C35194 a_n1435_47204# a_13059_46348# 2.88e-21
C35195 a_12861_44030# a_13693_46688# 5.48e-19
C35196 a_11453_44696# a_12816_46660# 8.81e-22
C35197 a_11599_46634# a_14180_46812# 2.26e-20
C35198 C6_P_btm C5_P_btm 18.2841f
C35199 C7_P_btm C4_P_btm 0.148546f
C35200 C9_P_btm C2_P_btm 0.144261f
C35201 C8_P_btm C3_P_btm 0.13616f
C35202 a_n743_46660# a_1302_46660# 0.002121f
C35203 a_n2661_46634# a_4955_46873# 0.03751f
C35204 a_5807_45002# a_5429_46660# 1.03e-19
C35205 EN_VIN_BSTR_N C1_N_btm 0.110046f
C35206 a_n2109_47186# a_n1853_46287# 3.06e-20
C35207 a_7227_47204# a_765_45546# 0.005844f
C35208 a_12465_44636# a_3090_45724# 1.51e-19
C35209 a_4883_46098# a_15368_46634# 0.023335f
C35210 a_22469_40625# VIN_N 2.79e-20
C35211 a_n1741_47186# a_n2293_46098# 2.17e-20
C35212 SMPL_ON_P a_n2472_46090# 2.92e-19
C35213 a_n1920_47178# a_n2157_46122# 7.93e-21
C35214 a_22609_37990# VDD 0.079488f
C35215 a_288_46660# a_1799_45572# 7.3e-22
C35216 a_948_46660# a_2609_46660# 2.98e-20
C35217 a_2107_46812# a_2443_46660# 0.013591f
C35218 a_9482_43914# CLK 3.96e-20
C35219 a_10341_43396# a_20749_43396# 0.003778f
C35220 a_n2661_42282# a_1576_42282# 2.11e-19
C35221 a_3422_30871# a_14113_42308# 5.01e-20
C35222 a_3626_43646# a_10341_42308# 0.001954f
C35223 a_2982_43646# a_12089_42308# 1.34e-19
C35224 a_7112_43396# a_7227_42852# 3.34e-19
C35225 a_7287_43370# a_7871_42858# 0.003663f
C35226 a_3905_42865# a_5932_42308# 0.003844f
C35227 a_15743_43084# a_15868_43402# 4.12e-21
C35228 a_17499_43370# a_16823_43084# 0.064861f
C35229 a_16243_43396# a_4190_30871# 1.24e-20
C35230 a_n2267_43396# a_n2293_42282# 6.24e-21
C35231 a_17339_46660# a_16409_43396# 4.94e-20
C35232 a_3232_43370# a_11691_44458# 0.251483f
C35233 a_3175_45822# a_1414_42308# 7.59e-22
C35234 a_n467_45028# a_n2129_44697# 0.007241f
C35235 a_8696_44636# a_10617_44484# 0.002097f
C35236 a_n913_45002# a_949_44458# 7.6e-21
C35237 a_n1059_45260# a_2779_44458# 8.54e-22
C35238 a_n357_42282# a_1241_44260# 3.97e-19
C35239 a_19692_46634# a_743_42282# 0.150479f
C35240 a_13259_45724# a_15493_43396# 0.021264f
C35241 a_n2956_38216# a_n2661_42282# 3.02e-20
C35242 a_n37_45144# a_n2661_44458# 8.09e-19
C35243 a_n443_42852# a_5663_43940# 3.4e-21
C35244 a_2304_45348# a_n2661_43370# 1.44e-19
C35245 w_1575_34946# a_n4064_39616# 0.027505f
C35246 a_18479_47436# a_21167_46155# 5.49e-19
C35247 a_5732_46660# a_6165_46155# 0.001142f
C35248 a_3785_47178# a_2711_45572# 1.05e-20
C35249 a_n443_46116# a_509_45572# 0.003835f
C35250 a_19333_46634# a_20107_46660# 1.09e-20
C35251 a_15227_44166# a_20411_46873# 0.041968f
C35252 a_13885_46660# a_13059_46348# 9.73e-19
C35253 a_18834_46812# a_20273_46660# 4.32e-20
C35254 a_n2312_38680# a_n2956_39304# 5.96956f
C35255 a_5257_43370# a_3483_46348# 0.028522f
C35256 a_9804_47204# a_8049_45260# 8.45e-19
C35257 a_8128_46384# a_9241_46436# 1.58e-20
C35258 a_12156_46660# a_765_45546# 0.001818f
C35259 a_4883_46098# a_19597_46482# 1.2e-19
C35260 a_11453_44696# a_18243_46436# 1.02e-19
C35261 a_13507_46334# a_20254_46482# 3.81e-19
C35262 a_19692_46634# a_19123_46287# 0.00443f
C35263 a_19466_46812# a_19551_46910# 0.008633f
C35264 a_4646_46812# a_8953_45546# 2.27e-20
C35265 a_n237_47217# a_3260_45572# 6.54e-22
C35266 a_n1151_42308# a_4099_45572# 9.09e-21
C35267 a_2063_45854# a_6511_45714# 0.037319f
C35268 a_n2293_46634# a_n1736_46482# 0.004173f
C35269 a_743_42282# a_196_42282# 7.61e-19
C35270 a_22165_42308# a_22959_42860# 6.47e-20
C35271 a_10695_43548# a_10533_42308# 9.55e-22
C35272 a_20596_44850# VDD 4.6e-19
C35273 a_13467_32519# COMP_P 5.83e-19
C35274 a_10518_42984# a_10793_43218# 0.007416f
C35275 a_3626_43646# a_18057_42282# 0.01061f
C35276 a_2982_43646# a_18907_42674# 8.43e-20
C35277 a_3080_42308# a_13258_32519# 7.3e-19
C35278 a_3422_30871# C8_N_btm 4.06e-19
C35279 a_8945_43396# a_5934_30871# 1.73e-20
C35280 a_n2312_38680# a_n3565_39304# 0.418567f
C35281 a_n913_45002# a_11341_43940# 0.001663f
C35282 a_n2017_45002# a_15493_43940# 9.45e-20
C35283 a_n2433_44484# a_n2293_43922# 0.010009f
C35284 a_1423_45028# a_3905_42865# 9.59e-20
C35285 a_17719_45144# a_11967_42832# 2.77e-21
C35286 a_18587_45118# a_18588_44850# 3.44e-19
C35287 a_16922_45042# a_20362_44736# 0.00806f
C35288 a_3232_43370# a_8333_44056# 2.98e-19
C35289 a_n443_42852# a_16243_43396# 0.001298f
C35290 a_20202_43084# a_20256_43172# 0.006261f
C35291 a_5883_43914# a_5891_43370# 0.216958f
C35292 a_8103_44636# a_8333_44734# 0.004937f
C35293 a_18374_44850# a_18989_43940# 3.56e-21
C35294 a_n2129_44697# a_n2661_43922# 0.00767f
C35295 a_n2267_44484# a_n2661_42834# 0.002133f
C35296 a_949_44458# a_556_44484# 0.001921f
C35297 a_1307_43914# a_7281_43914# 0.004629f
C35298 a_7229_43940# a_n2661_42282# 2.13e-19
C35299 a_526_44458# a_10922_42852# 2.42e-20
C35300 a_11827_44484# a_17517_44484# 0.05115f
C35301 a_3090_45724# a_8515_42308# 1.5e-21
C35302 a_11599_46634# a_11787_45002# 1.65e-20
C35303 a_n2109_47186# a_n2661_43370# 0.008032f
C35304 a_n971_45724# a_8488_45348# 0.001106f
C35305 a_4704_46090# a_n1925_42282# 2.45e-19
C35306 a_6755_46942# a_10180_45724# 4.84e-20
C35307 a_10249_46116# a_10193_42453# 0.034764f
C35308 a_10623_46897# a_10490_45724# 3.15e-20
C35309 a_20411_46873# a_21071_46482# 2.24e-19
C35310 a_5807_45002# a_20107_45572# 4.31e-21
C35311 a_13661_43548# a_18953_45572# 5.68e-19
C35312 a_11117_47542# a_2437_43646# 5.27e-19
C35313 a_9290_44172# a_10809_44734# 0.239594f
C35314 a_n443_46116# a_2809_45348# 0.001393f
C35315 a_n237_47217# a_n2293_42834# 0.002403f
C35316 a_3090_45724# a_2711_45572# 0.555348f
C35317 a_n743_46660# a_16842_45938# 1.64e-19
C35318 SMPL_ON_N a_413_45260# 0.199669f
C35319 a_8128_46384# a_3357_43084# 5.77e-20
C35320 a_12861_44030# a_13348_45260# 2.51e-20
C35321 a_1823_45246# a_5210_46155# 1.93e-20
C35322 a_1755_42282# a_2713_42308# 9.85e-19
C35323 a_1606_42308# a_2903_42308# 0.001317f
C35324 a_5342_30871# a_n3420_39072# 0.062032f
C35325 a_n1059_45260# a_n13_43084# 0.027848f
C35326 a_n913_45002# a_n1076_43230# 0.05439f
C35327 a_n2017_45002# a_n3674_39304# 6.29e-20
C35328 a_n2956_39304# a_7174_31319# 4.27e-21
C35329 a_n1917_44484# a_n1917_43396# 9.63e-19
C35330 a_n2267_44484# a_n1352_43396# 6.41e-21
C35331 a_n1352_44484# a_n2267_43396# 2.85e-20
C35332 a_10249_46116# VDD 1.03004f
C35333 a_11541_44484# a_11750_44172# 2.79e-19
C35334 a_3537_45260# a_4361_42308# 0.017454f
C35335 a_413_45260# a_22959_43396# 2.15e-19
C35336 en_comp a_n1991_42858# 2.41e-19
C35337 a_n967_45348# a_n1853_43023# 0.021497f
C35338 a_n1761_44111# a_n1549_44318# 0.033724f
C35339 a_n2065_43946# a_n809_44244# 0.043475f
C35340 a_n1899_43946# a_n1331_43914# 0.171939f
C35341 a_18494_42460# a_3626_43646# 0.066461f
C35342 a_n2661_44458# a_104_43370# 8.68e-21
C35343 a_11823_42460# a_12991_43230# 0.001129f
C35344 a_3357_43084# a_1847_42826# 0.010588f
C35345 a_n755_45592# a_n327_42308# 7.83e-20
C35346 a_n357_42282# a_n39_42308# 0.001655f
C35347 a_19321_45002# a_17970_44736# 1.04e-21
C35348 a_2107_46812# a_949_44458# 8.97e-21
C35349 a_n2661_45546# a_n1013_45572# 0.001202f
C35350 a_13661_43548# a_18443_44721# 0.011774f
C35351 a_13747_46662# a_18287_44626# 1.75e-20
C35352 a_15682_46116# a_16680_45572# 0.006985f
C35353 a_2324_44458# a_8696_44636# 0.033373f
C35354 a_17715_44484# a_16115_45572# 6.11e-20
C35355 a_10227_46804# a_16241_44734# 4.02e-19
C35356 a_n1079_45724# a_n356_45724# 9.52e-19
C35357 a_n2661_46634# a_12607_44458# 1.26e-19
C35358 a_8049_45260# a_10180_45724# 0.002472f
C35359 a_n2661_46098# a_n2433_44484# 5.13e-22
C35360 a_12861_44030# a_19615_44636# 0.094785f
C35361 a_n2312_40392# a_n2661_43922# 1.45e-20
C35362 a_n2312_39304# a_n2661_42834# 6.52e-20
C35363 a_12465_44636# a_14815_43914# 3.16e-19
C35364 a_584_46384# a_n1761_44111# 1.76e-20
C35365 a_n971_45724# a_1414_42308# 4.43e-21
C35366 a_n746_45260# a_1467_44172# 9.96e-21
C35367 a_8270_45546# a_n2293_42834# 1.57e-20
C35368 a_10903_43370# a_13485_45572# 0.001122f
C35369 a_14035_46660# a_9482_43914# 8.69e-20
C35370 a_n2293_46634# a_10440_44484# 3.4e-20
C35371 a_n357_42282# a_997_45618# 0.023595f
C35372 a_n4315_30879# a_n4064_39616# 0.034877f
C35373 a_5932_42308# a_n3420_37440# 5.13e-19
C35374 a_1209_47178# a_2063_45854# 0.00786f
C35375 a_1431_47204# a_2124_47436# 0.010942f
C35376 a_n971_45724# a_3381_47502# 0.008848f
C35377 a_n746_45260# a_n1151_42308# 0.116939f
C35378 a_1239_47204# a_584_46384# 1.75e-19
C35379 a_n1741_47186# a_4791_45118# 0.024211f
C35380 a_n2109_47186# a_4915_47217# 0.352259f
C35381 a_n237_47217# a_3160_47472# 0.037234f
C35382 a_7174_31319# a_n3565_39304# 4.27e-21
C35383 a_n4064_40160# a_n3420_39616# 0.05705f
C35384 a_375_42282# a_n327_42558# 7.38e-21
C35385 a_22959_43948# a_17538_32519# 0.168682f
C35386 a_15493_43940# a_21845_43940# 5.9e-19
C35387 a_3065_45002# a_6123_31319# 9.58e-21
C35388 a_n913_45002# a_10723_42308# 0.006785f
C35389 a_n1059_45260# a_11323_42473# 6.13e-20
C35390 a_n2017_45002# a_5742_30871# 0.007608f
C35391 a_3499_42826# a_3626_43646# 0.001049f
C35392 a_6453_43914# a_6452_43396# 8.84e-19
C35393 a_n2661_42834# a_n2472_42826# 0.03087f
C35394 a_19328_44172# a_n97_42460# 9.4e-21
C35395 a_19615_44636# a_19700_43370# 1.17e-20
C35396 a_11967_42832# a_16664_43396# 1.34e-19
C35397 a_n356_44636# a_7765_42852# 1.83e-20
C35398 a_3537_45260# a_6761_42308# 0.057884f
C35399 a_2382_45260# a_5934_30871# 1.02e-20
C35400 a_5111_44636# a_6171_42473# 2.14e-20
C35401 a_9290_44172# a_5883_43914# 0.026946f
C35402 a_16855_45546# a_8696_44636# 0.112262f
C35403 a_15227_44166# a_3422_30871# 2.1e-20
C35404 a_5937_45572# a_8975_43940# 6.52e-19
C35405 a_8953_45546# a_10057_43914# 1.06e-19
C35406 a_15765_45572# a_16020_45572# 0.056391f
C35407 a_16327_47482# a_2982_43646# 0.030062f
C35408 a_21076_30879# a_9313_44734# 1.55e-20
C35409 a_n443_42852# a_3232_43370# 0.02112f
C35410 a_n3420_38528# VREF 2.43e-19
C35411 a_2063_45854# a_10768_47026# 0.005084f
C35412 a_n1613_43370# a_n743_46660# 0.521102f
C35413 CAL_N a_22469_40625# 0.007453f
C35414 a_n3565_38502# VCM 0.035399f
C35415 a_n1435_47204# a_7577_46660# 5.91e-21
C35416 a_6151_47436# a_6969_46634# 0.030417f
C35417 a_6545_47178# a_6755_46942# 0.022995f
C35418 a_9863_47436# a_9863_46634# 0.003636f
C35419 a_9313_45822# a_8667_46634# 0.004188f
C35420 a_n881_46662# a_n1021_46688# 0.15991f
C35421 a_n4064_38528# VIN_P 0.044919f
C35422 a_16131_47204# a_5807_45002# 6.5e-19
C35423 a_n2946_37984# VDD 0.38275f
C35424 a_n1699_43638# a_n1991_42858# 4.92e-20
C35425 a_n1917_43396# a_n1853_43023# 0.001737f
C35426 a_n2267_43396# a_n1423_42826# 0.001766f
C35427 a_n1177_43370# a_n2157_42858# 6.59e-19
C35428 a_n2129_43609# a_n1641_43230# 1.1e-19
C35429 a_4699_43561# a_743_42282# 1.35e-20
C35430 a_19963_31679# C8_N_btm 1.65e-20
C35431 a_15493_43940# a_19164_43230# 3.58e-20
C35432 a_11341_43940# a_20922_43172# 7.6e-21
C35433 a_n2661_42834# a_9223_42460# 8.65e-22
C35434 a_n2293_43922# a_8685_42308# 3.58e-20
C35435 a_n4318_40392# a_n4064_39616# 6.39e-21
C35436 a_22223_45572# VDD 0.287831f
C35437 a_14358_43442# a_14205_43396# 0.163543f
C35438 a_9803_43646# a_10341_43396# 0.11445f
C35439 a_14579_43548# a_15095_43370# 0.109081f
C35440 a_9145_43396# a_10765_43646# 0.00303f
C35441 a_8685_43396# a_9885_43396# 4.64e-19
C35442 a_2437_43646# RST_Z 0.082469f
C35443 a_14021_43940# a_15279_43071# 5.5e-21
C35444 a_20447_31679# C6_N_btm 0.001141f
C35445 a_6511_45714# a_n2661_42834# 6.91e-21
C35446 a_11823_42460# a_n356_44636# 5.09e-19
C35447 a_7499_43078# a_7640_43914# 0.021219f
C35448 a_3090_45724# a_7466_43396# 9.39e-20
C35449 a_10951_45334# a_9482_43914# 5.58e-21
C35450 a_2711_45572# a_14815_43914# 9.7e-21
C35451 a_6171_45002# a_16751_45260# 0.104212f
C35452 a_5147_45002# a_1423_45028# 0.017515f
C35453 a_n2312_39304# a_n2293_42282# 4.65e-20
C35454 a_10809_44734# a_10807_43548# 1.71e-19
C35455 a_18341_45572# a_11691_44458# 4.3e-20
C35456 a_n2017_45002# a_n2293_42834# 0.28698f
C35457 a_18479_45785# a_20193_45348# 1.42e-21
C35458 a_n2497_47436# a_n961_42308# 1.14e-20
C35459 SMPL_ON_P a_n3674_38216# 0.044338f
C35460 a_18189_46348# a_15493_43396# 4.56e-21
C35461 a_3065_45002# a_3495_45348# 0.001093f
C35462 a_n357_42282# a_11967_42832# 0.153035f
C35463 a_8162_45546# a_5891_43370# 4.81e-19
C35464 a_4955_46873# a_765_45546# 0.008652f
C35465 a_10249_46116# a_10185_46660# 7.29e-19
C35466 a_11453_44696# a_18819_46122# 7.1e-20
C35467 a_13507_46334# a_6945_45028# 0.187229f
C35468 a_20990_47178# a_10809_44734# 0.00204f
C35469 a_n743_46660# a_n2293_46098# 0.213418f
C35470 a_n2438_43548# a_n2472_46090# 0.020059f
C35471 a_n1925_46634# a_n1853_46287# 0.012373f
C35472 a_n2312_38680# a_n1991_46122# 2.37e-19
C35473 a_n2293_46634# a_n1641_46494# 0.002502f
C35474 a_10554_47026# a_10425_46660# 4.2e-19
C35475 a_9804_47204# a_8953_45546# 3.84e-19
C35476 a_11735_46660# a_11813_46116# 0.162547f
C35477 a_8128_46384# a_9625_46129# 3.11e-20
C35478 a_12465_44636# a_20075_46420# 5.91e-21
C35479 a_n1021_46688# a_n2157_46122# 0.00108f
C35480 a_5807_45002# a_3483_46348# 0.018693f
C35481 a_7903_47542# a_8034_45724# 8.49e-21
C35482 a_4883_46098# a_20708_46348# 0.014516f
C35483 a_n97_42460# a_8685_42308# 2.19e-19
C35484 a_6031_43396# a_1755_42282# 3.75e-21
C35485 a_5205_44734# VDD 0.001314f
C35486 a_n2472_42826# a_n2293_42282# 3.06e-19
C35487 a_2982_43646# a_5267_42460# 1.03e-19
C35488 a_4905_42826# a_5337_42558# 0.005481f
C35489 a_3539_42460# a_2903_42308# 6.02e-19
C35490 a_11967_42832# CAL_N 0.001103f
C35491 a_9127_43156# a_10796_42968# 1.62e-19
C35492 a_10083_42826# a_10518_42984# 0.234322f
C35493 a_18587_45118# a_18443_44721# 7.68e-20
C35494 a_18911_45144# a_18287_44626# 3.74e-19
C35495 a_n2661_43370# a_8375_44464# 9.68e-20
C35496 a_11691_44458# a_8975_43940# 0.048259f
C35497 a_11827_44484# a_13720_44458# 0.00996f
C35498 a_n2312_39304# a_n3565_39590# 0.491833f
C35499 a_4185_45028# a_8952_43230# 3.54e-21
C35500 a_20202_43084# a_21195_42852# 0.018373f
C35501 a_n357_42282# a_648_43396# 0.003365f
C35502 a_n2661_44458# a_949_44458# 0.041721f
C35503 a_413_45260# a_22959_44484# 0.202222f
C35504 a_n967_45348# a_n1899_43946# 0.025102f
C35505 a_n2661_45010# a_2127_44172# 0.096614f
C35506 a_3357_43084# a_5244_44056# 1.59e-20
C35507 a_n2293_45010# a_1414_42308# 3e-19
C35508 a_n2017_45002# a_1115_44172# 3.58e-21
C35509 a_n1059_45260# a_644_44056# 6.29e-19
C35510 a_n745_45366# a_n984_44318# 1.8e-20
C35511 a_14537_43396# a_15367_44484# 0.001966f
C35512 a_n2129_44697# a_n452_44636# 0.079904f
C35513 a_n2267_44484# a_n1352_44484# 0.118759f
C35514 a_1307_43914# a_16241_44734# 0.010259f
C35515 a_n443_42852# a_4905_42826# 0.037419f
C35516 a_5257_43370# a_n357_42282# 3.28e-19
C35517 a_12741_44636# a_13759_46122# 1e-20
C35518 a_768_44030# a_10907_45822# 7.18e-20
C35519 a_6151_47436# a_3357_43084# 0.025786f
C35520 a_3699_46634# a_2711_45572# 0.001403f
C35521 a_n743_46660# a_7230_45938# 8.13e-19
C35522 a_13661_43548# a_13249_42308# 0.486588f
C35523 a_5807_45002# a_14495_45572# 0.012666f
C35524 a_13747_46662# a_13904_45546# 0.031534f
C35525 a_11415_45002# a_14275_46494# 1.84e-19
C35526 a_20528_46660# a_20075_46420# 4.61e-19
C35527 a_18280_46660# a_17957_46116# 1.49e-19
C35528 a_21363_46634# a_21137_46414# 0.001902f
C35529 a_19692_46634# a_8049_45260# 0.045516f
C35530 a_20623_46660# a_6945_45028# 0.004994f
C35531 a_20273_46660# a_10809_44734# 0.027345f
C35532 a_11901_46660# a_12839_46116# 3.72e-20
C35533 a_6851_47204# a_2437_43646# 0.003764f
C35534 a_18597_46090# a_18175_45572# 0.002203f
C35535 a_n2661_46634# a_8746_45002# 3.38e-20
C35536 a_1823_45246# a_5497_46414# 1.22e-20
C35537 a_3483_46348# a_3699_46348# 0.06281f
C35538 a_n237_47217# a_413_45260# 0.030002f
C35539 a_n746_45260# a_327_44734# 0.256943f
C35540 a_n971_45724# a_1667_45002# 1.51e-19
C35541 a_18780_47178# a_18479_45785# 1.02e-21
C35542 a_18479_47436# a_18341_45572# 3.11e-21
C35543 a_16327_47482# a_16789_45572# 4.55e-19
C35544 a_15567_42826# a_15051_42282# 0.001656f
C35545 a_5342_30871# a_15486_42560# 0.006845f
C35546 a_5193_42852# a_5379_42460# 3.15e-19
C35547 a_14401_32519# C1_N_btm 6.64e-20
C35548 a_12089_42308# a_11897_42308# 1.97e-19
C35549 a_16414_43172# a_14113_42308# 0.004427f
C35550 a_4190_30871# a_n4064_39072# 1.46e-20
C35551 a_13565_43940# VDD 0.175245f
C35552 a_n2472_46634# VDD 0.287589f
C35553 a_10334_44484# a_10405_44172# 0.002711f
C35554 a_n2661_43922# a_n2472_43914# 0.068474f
C35555 a_n2661_42834# a_n2065_43946# 0.035267f
C35556 a_8975_43940# a_8333_44056# 7.34e-19
C35557 a_11823_42460# a_12379_42858# 0.033971f
C35558 a_13747_46662# CLK 3.82e-20
C35559 a_10193_42453# a_5534_30871# 0.136243f
C35560 a_n357_42282# a_9114_42852# 1.14e-19
C35561 a_13259_45724# a_18707_42852# 1.69e-20
C35562 a_n2661_44458# a_11341_43940# 0.001405f
C35563 a_3537_45260# a_7274_43762# 4.26e-19
C35564 a_n913_45002# a_10341_43396# 0.032712f
C35565 a_1307_43914# a_n1557_42282# 6.39e-20
C35566 a_n2293_43922# a_n2840_43914# 0.001304f
C35567 a_n443_42852# a_7573_43172# 4.79e-19
C35568 a_n1925_42282# a_2713_42308# 7.52e-20
C35569 a_526_44458# a_2903_42308# 5.08e-21
C35570 a_10903_43370# a_13070_42354# 0.04369f
C35571 a_20193_45348# a_14021_43940# 0.118757f
C35572 a_n2956_39304# a_5932_42308# 3.95e-21
C35573 a_18588_44850# a_11967_42832# 8.49e-19
C35574 a_1423_45028# a_4093_43548# 1.31e-20
C35575 a_n1925_46634# a_n2661_43370# 1.37e-20
C35576 a_3483_46348# a_15143_45578# 1.45e-21
C35577 a_16327_47482# a_14539_43914# 0.031714f
C35578 a_9625_46129# a_10053_45546# 0.086776f
C35579 a_8199_44636# a_8746_45002# 0.680077f
C35580 a_5937_45572# a_10193_42453# 4.34e-20
C35581 a_4185_45028# a_13249_42308# 3.74e-20
C35582 a_12549_44172# a_11827_44484# 1.40268f
C35583 a_10623_46897# a_6171_45002# 1.49e-20
C35584 a_n1151_42308# a_n310_44484# 0.00221f
C35585 a_19123_46287# a_18175_45572# 7.15e-20
C35586 a_18285_46348# a_18479_45785# 2.17e-20
C35587 a_11599_46634# a_18287_44626# 3.51e-19
C35588 a_8049_45260# a_20692_30879# 5.54e-20
C35589 a_5807_45002# a_17719_45144# 4.18e-21
C35590 a_13661_43548# a_17613_45144# 1.21e-20
C35591 a_4791_45118# a_8238_44734# 0.001045f
C35592 a_11415_45002# a_15765_45572# 0.003223f
C35593 a_526_44458# a_3218_45724# 0.032949f
C35594 a_2324_44458# a_7227_45028# 0.035814f
C35595 a_19692_46634# a_19479_31679# 5.21e-19
C35596 a_19466_46812# a_3357_43084# 0.006916f
C35597 a_5342_30871# C10_N_btm 2.16e-19
C35598 a_14113_42308# a_7174_31319# 4.19e-20
C35599 a_17124_42282# a_4958_30871# 0.20224f
C35600 a_16522_42674# a_17303_42282# 2.42e-20
C35601 COMP_P a_2113_38308# 1.33e-19
C35602 a_5934_30871# a_1239_39587# 1.67e-19
C35603 a_5932_42308# a_n3565_39304# 3.95e-21
C35604 a_5534_30871# VDD 0.513761f
C35605 a_n2661_43922# a_10695_43548# 1.39e-20
C35606 a_9313_44734# a_12281_43396# 0.027032f
C35607 a_n2810_45572# a_n3565_38216# 0.104999f
C35608 a_18079_43940# a_15493_43940# 0.040279f
C35609 a_18451_43940# a_11341_43940# 0.004129f
C35610 a_10193_42453# a_19647_42308# 0.004706f
C35611 a_7499_43078# a_7174_31319# 9.76e-21
C35612 a_n1917_44484# a_n1853_43023# 1.77e-20
C35613 en_comp a_22400_42852# 0.730145f
C35614 a_11750_44172# a_11816_44260# 0.006978f
C35615 a_10949_43914# a_12603_44260# 0.001915f
C35616 a_19862_44208# a_20365_43914# 0.075162f
C35617 a_14539_43914# a_16855_43396# 9.74e-19
C35618 a_n1761_44111# a_n1177_43370# 1.22e-19
C35619 a_n1549_44318# a_n2267_43396# 9.07e-20
C35620 a_n1331_43914# a_n1699_43638# 1.55e-19
C35621 a_n2065_43946# a_n1352_43396# 0.009873f
C35622 a_n809_44244# a_n2129_43609# 3.98e-20
C35623 a_n1899_43946# a_n1917_43396# 4.39e-19
C35624 a_5937_45572# VDD 2.20055f
C35625 a_11652_45724# a_10907_45822# 1.68e-19
C35626 a_21076_30879# a_18114_32519# 0.054909f
C35627 a_768_44030# a_n2661_42282# 0.002669f
C35628 a_20205_31679# a_3357_43084# 3.97e-19
C35629 a_20692_30879# a_19479_31679# 0.051569f
C35630 a_11322_45546# a_11682_45822# 0.034435f
C35631 a_5066_45546# a_8953_45002# 0.013782f
C35632 a_2711_45572# a_13297_45572# 8.55e-20
C35633 a_n2293_46634# a_5244_44056# 1.54e-20
C35634 a_11453_44696# a_11341_43940# 0.006646f
C35635 a_10227_46804# a_15037_44260# 2.81e-19
C35636 a_14495_45572# a_15143_45578# 8.73e-19
C35637 a_n971_45724# a_n1190_43762# 3.04e-20
C35638 a_9290_44172# a_11361_45348# 4.93e-19
C35639 a_7174_31319# C8_N_btm 7.53e-20
C35640 a_n4064_40160# C2_P_btm 1.17e-19
C35641 a_584_46384# a_491_47026# 5.54e-20
C35642 a_n785_47204# a_n2661_46098# 3.17e-20
C35643 a_4791_45118# a_n743_46660# 0.080217f
C35644 a_n3565_39590# C8_P_btm 0.384801f
C35645 a_16327_47482# a_16119_47582# 1.79e-19
C35646 a_16023_47582# a_15928_47570# 0.049827f
C35647 a_4883_46098# a_5063_47570# 2.16e-22
C35648 a_n1151_42308# a_383_46660# 0.002404f
C35649 a_4915_47217# a_n1925_46634# 1.12e-19
C35650 a_n3420_39616# C10_P_btm 2.16e-19
C35651 VDAC_Pi VDAC_Ni 3.18068f
C35652 a_n4064_37984# a_n4064_37440# 0.061238f
C35653 a_6851_47204# a_n2661_46634# 9.8e-20
C35654 a_12861_44030# a_13661_43548# 0.8566f
C35655 a_13717_47436# a_13747_46662# 0.003701f
C35656 a_13487_47204# a_5807_45002# 5.04e-20
C35657 a_n237_47217# a_2609_46660# 4.06e-20
C35658 a_n971_45724# a_2959_46660# 2.33e-19
C35659 a_n4209_39304# a_n1386_35608# 9.16e-20
C35660 a_19511_42282# RST_Z 2.38e-20
C35661 a_10227_46804# a_11309_47204# 0.026748f
C35662 a_16588_47582# a_12549_44172# 2.25e-20
C35663 a_19647_42308# VDD 0.227331f
C35664 a_4699_43561# a_2813_43396# 1.26e-20
C35665 a_2982_43646# a_6547_43396# 4.43e-21
C35666 a_15493_43940# a_14209_32519# 3.85e-21
C35667 a_3626_43646# a_6197_43396# 3.15e-20
C35668 a_n356_44636# a_961_42354# 0.005209f
C35669 a_4093_43548# a_4181_43396# 2.48e-19
C35670 a_16922_45042# a_17303_42282# 1.31e-20
C35671 a_n2661_42282# a_5755_42852# 0.006322f
C35672 a_5343_44458# a_5934_30871# 7.67e-19
C35673 a_n97_42460# a_9803_43646# 1.56e-20
C35674 a_14021_43940# a_20301_43646# 0.024612f
C35675 a_11341_43940# a_17364_32525# 0.005541f
C35676 a_10193_42453# a_11691_44458# 0.046462f
C35677 en_comp a_n967_45348# 0.001993f
C35678 a_13661_43548# a_19700_43370# 0.042923f
C35679 a_1823_45246# a_5841_44260# 1.17e-20
C35680 a_2437_43646# a_3232_43370# 2.01e-19
C35681 a_n1613_43370# a_4361_42308# 1.74e-19
C35682 a_4099_45572# a_4223_44672# 3.68e-19
C35683 a_2711_45572# a_4743_44484# 4.71e-21
C35684 a_n443_42852# a_8975_43940# 0.001317f
C35685 a_n357_42282# a_18989_43940# 6.13e-20
C35686 a_5937_45572# a_5495_43940# 3.03e-19
C35687 a_n745_45366# a_n467_45028# 0.110406f
C35688 a_3357_43084# a_5111_44636# 0.318002f
C35689 SMPL_ON_N a_20820_30879# 0.029764f
C35690 a_5263_46660# a_5257_43370# 2.87e-20
C35691 a_n1151_42308# a_13351_46090# 5.07e-20
C35692 a_n743_46660# a_16292_46812# 0.064277f
C35693 a_12549_44172# a_14447_46660# 9.1e-20
C35694 a_11453_44696# a_22591_46660# 7.09e-19
C35695 VIN_N VREF 0.775904f
C35696 a_n2833_47464# a_n2956_38680# 1.71e-20
C35697 a_n2497_47436# a_n2956_39304# 2.52e-20
C35698 a_3877_44458# a_6755_46942# 0.388535f
C35699 a_6151_47436# a_9625_46129# 2.77e-19
C35700 a_7903_47542# a_8016_46348# 1.87e-20
C35701 a_6575_47204# a_7920_46348# 3.65e-19
C35702 VIN_P VREF_GND 16.4969f
C35703 a_5807_45002# a_14513_46634# 0.006821f
C35704 a_13747_46662# a_14035_46660# 0.040628f
C35705 a_13759_47204# a_13059_46348# 1.99e-19
C35706 a_12861_44030# a_4185_45028# 2.17e-20
C35707 a_n1741_47186# a_6945_45028# 2.51584f
C35708 a_4883_46098# a_21542_46660# 5.31e-19
C35709 a_12465_44636# a_21076_30879# 2.7e-19
C35710 a_13483_43940# a_13575_42558# 1.75e-21
C35711 a_11691_44458# VDD 3.25709f
C35712 a_18114_32519# C0_N_btm 3.38e-19
C35713 a_n2157_42858# a_n1991_42858# 0.905962f
C35714 a_10341_43396# a_20922_43172# 8.95e-20
C35715 a_n97_42460# a_19518_43218# 3.81e-19
C35716 a_743_42282# a_1847_42826# 0.004285f
C35717 a_16922_45042# a_19778_44110# 0.026041f
C35718 a_n745_45366# a_n2661_43922# 2.34e-20
C35719 a_n913_45002# a_n2293_43922# 0.019153f
C35720 a_10227_46804# a_15890_42674# 0.159412f
C35721 a_4185_45028# a_19700_43370# 1.48e-22
C35722 a_n2438_43548# a_n3674_38216# 5.26e-20
C35723 a_526_44458# a_6293_42852# 0.029694f
C35724 a_7499_43078# a_10729_43914# 0.23002f
C35725 a_21076_30879# a_13887_32519# 0.055154f
C35726 a_n2956_39768# a_n3674_37592# 0.031375f
C35727 a_1423_45028# a_10157_44484# 5.42e-19
C35728 a_n1613_43370# a_6761_42308# 4.15e-20
C35729 a_17719_45144# a_18315_45260# 0.017382f
C35730 a_3537_45260# a_5891_43370# 0.359819f
C35731 a_5147_45002# a_6109_44484# 7.39e-19
C35732 a_14537_43396# a_14539_43914# 0.135541f
C35733 a_1307_43914# a_12883_44458# 2.26e-21
C35734 a_5807_45002# a_n357_42282# 6.44e-20
C35735 a_n2956_39768# a_n2840_45546# 7e-20
C35736 a_13607_46688# a_13759_46122# 0.004856f
C35737 a_11813_46116# a_2324_44458# 1.71e-20
C35738 a_18479_47436# a_10193_42453# 8.24e-21
C35739 a_765_45546# a_376_46348# 1.21e-19
C35740 a_10227_46804# a_10490_45724# 0.031f
C35741 a_11599_46634# a_13904_45546# 6.03e-20
C35742 a_14209_32519# a_5742_30871# 0.005505f
C35743 a_18525_43370# a_18057_42282# 6.86e-21
C35744 a_743_42282# a_15486_42560# 0.010882f
C35745 a_22165_42308# a_22400_42852# 0.005425f
C35746 a_21671_42860# a_14097_32519# 8.99e-20
C35747 a_8333_44056# VDD 0.124235f
C35748 a_5649_42852# a_13070_42354# 6.66e-20
C35749 a_4190_30871# a_15803_42450# 1.32e-19
C35750 a_5534_30871# a_n784_42308# 9.92256f
C35751 a_19987_42826# a_20753_42852# 0.07365f
C35752 a_15743_43084# a_17303_42282# 1.95e-20
C35753 a_4361_42308# a_13249_42558# 7.13e-20
C35754 a_n2661_44458# a_175_44278# 5.37e-21
C35755 a_3357_43084# a_4235_43370# 0.00216f
C35756 a_n443_42852# a_2905_42968# 3.32e-21
C35757 a_10193_42453# a_4190_30871# 0.305842f
C35758 a_13259_45724# a_21356_42826# 1.24e-20
C35759 a_10227_46804# START 0.088203f
C35760 a_19692_46634# a_13258_32519# 1.9e-20
C35761 a_15227_44166# a_7174_31319# 5.34e-21
C35762 a_18143_47464# RST_Z 2.7e-19
C35763 a_n967_45348# a_n1699_43638# 0.001377f
C35764 a_3363_44484# a_n2661_43922# 0.005466f
C35765 a_n1917_44484# a_n1899_43946# 0.012479f
C35766 a_n2267_44484# a_n1549_44318# 5.88e-19
C35767 a_n1352_44484# a_n2065_43946# 0.00236f
C35768 a_n1177_44458# a_n1761_44111# 4.25e-20
C35769 a_n2129_44697# a_n809_44244# 3.14e-20
C35770 a_18443_44721# a_11967_42832# 0.035979f
C35771 a_18287_44626# a_19615_44636# 9.28e-19
C35772 a_n2017_45002# a_n2012_43396# 0.009581f
C35773 a_n913_45002# a_n97_42460# 0.109647f
C35774 a_n1059_45260# a_104_43370# 1.35e-20
C35775 a_n2293_45010# a_n1190_43762# 4.42e-20
C35776 a_n2661_43370# a_10949_43914# 2.82e-20
C35777 a_8696_44636# a_14579_43548# 5.14e-23
C35778 a_18479_47436# VDD 1.47669f
C35779 a_n357_42282# a_10518_42984# 0.010947f
C35780 a_11599_46634# CLK 6.41e-19
C35781 a_10227_46804# a_14976_45348# 7.06e-20
C35782 a_14275_46494# a_13259_45724# 2.55e-19
C35783 a_12549_44172# a_15595_45028# 6.29e-22
C35784 a_3483_46348# a_n755_45592# 5.99e-19
C35785 a_n237_47217# a_2779_44458# 8.08e-21
C35786 a_765_45546# a_8746_45002# 2.27e-20
C35787 a_11599_46634# a_17023_45118# 3.91e-20
C35788 a_6945_45028# a_10586_45546# 3.78e-20
C35789 a_n971_45724# a_n699_43396# 0.139047f
C35790 a_383_46660# a_327_44734# 1.22e-20
C35791 a_n743_46660# a_3429_45260# 1.28e-20
C35792 a_n1925_46634# a_4574_45260# 2.53e-20
C35793 a_n2293_46634# a_5111_44636# 0.130609f
C35794 a_13059_46348# a_13163_45724# 0.00596f
C35795 a_15009_46634# a_15037_45618# 1.9e-20
C35796 a_4651_46660# a_2437_43646# 7.1e-21
C35797 a_12861_44030# a_18587_45118# 0.011009f
C35798 a_n2661_46634# a_3232_43370# 3e-21
C35799 a_n1853_46287# a_n310_45572# 2.88e-19
C35800 a_13678_32519# C3_N_btm 0.001771f
C35801 a_4190_30871# VDD 1.36846f
C35802 a_8685_42308# a_10533_42308# 4.55e-21
C35803 a_13467_32519# C6_N_btm 1.49e-19
C35804 a_20820_30879# a_19864_35138# 1.44e-20
C35805 a_n356_44636# a_2982_43646# 0.434193f
C35806 a_17829_46910# VDD 0.37446f
C35807 a_7281_43914# a_7584_44260# 0.001377f
C35808 a_18911_45144# a_19268_43646# 5.23e-21
C35809 a_18494_42460# a_18525_43370# 4.73e-19
C35810 a_18184_42460# a_18783_43370# 2.81e-21
C35811 a_19778_44110# a_15743_43084# 0.00304f
C35812 en_comp a_22223_42860# 4.89e-22
C35813 a_n2017_45002# a_n914_42852# 1.25e-19
C35814 a_n2661_44458# a_10341_43396# 7.76e-20
C35815 a_20692_30879# a_13258_32519# 0.055049f
C35816 a_17339_46660# START 0.00197f
C35817 a_17730_32519# a_15493_43940# 0.006052f
C35818 a_n2661_43922# a_n2433_43396# 0.001232f
C35819 a_n2661_42834# a_n2129_43609# 0.009349f
C35820 a_n2293_43922# a_n4318_39304# 5.19e-19
C35821 a_n2810_45028# a_n2293_42282# 1.93e-20
C35822 a_n443_42852# a_15803_42450# 6.37e-21
C35823 a_1307_43914# a_3935_42891# 0.318189f
C35824 a_11691_44458# a_16137_43396# 5.49e-20
C35825 a_765_45546# RST_Z 0.002113f
C35826 a_2711_45572# a_4808_45572# 9.57e-19
C35827 a_9290_44172# a_3537_45260# 2.24e-20
C35828 a_22223_46124# a_20447_31679# 9.73e-19
C35829 a_n443_42852# a_10193_42453# 0.026599f
C35830 a_3483_46348# a_13017_45260# 0.51131f
C35831 a_13259_45724# a_15765_45572# 0.025388f
C35832 a_8199_44636# a_3232_43370# 0.32342f
C35833 a_8349_46414# a_6171_45002# 1.52e-21
C35834 a_5937_45572# a_5691_45260# 0.061637f
C35835 a_22959_46124# a_19963_31679# 3.42e-20
C35836 a_10809_44734# a_22959_45572# 3.06e-19
C35837 a_8049_45260# a_18175_45572# 0.014402f
C35838 a_19692_46634# a_20193_45348# 0.060606f
C35839 a_13759_46122# a_413_45260# 1.21e-20
C35840 a_6667_45809# a_7227_45028# 4.77e-19
C35841 a_n3565_38502# a_n4064_38528# 0.228245f
C35842 a_n4064_39072# a_n3420_37984# 0.045543f
C35843 a_n3420_39072# a_n4064_37984# 0.045827f
C35844 a_5934_30871# C1_N_btm 0.011025f
C35845 a_13717_47436# a_11599_46634# 3.05e-19
C35846 a_12861_44030# a_14955_47212# 6.92e-20
C35847 a_n2109_47186# a_n881_46662# 0.023562f
C35848 a_n971_45724# a_2266_47243# 0.00941f
C35849 a_n785_47204# a_n310_47243# 0.001173f
C35850 a_1209_47178# a_2487_47570# 2.94e-19
C35851 a_5337_42558# VDD 0.008564f
C35852 a_6123_31319# C3_N_btm 0.011333f
C35853 a_5932_42308# C8_N_btm 1.4e-19
C35854 a_4958_30871# VDAC_P 0.01779f
C35855 a_13487_47204# a_14311_47204# 0.00114f
C35856 a_n1761_44111# a_n1991_42858# 1.58e-21
C35857 a_n1899_43946# a_n1853_43023# 4.54e-20
C35858 a_n1331_43914# a_n2157_42858# 3.92e-20
C35859 a_18451_43940# a_10341_43396# 1.01e-20
C35860 a_11341_43940# a_9145_43396# 0.017582f
C35861 a_5244_44056# a_743_42282# 1.87e-21
C35862 a_1307_43914# a_15890_42674# 3.24e-21
C35863 en_comp a_n4209_39590# 7.54e-19
C35864 a_n2267_43396# a_n1177_43370# 0.041762f
C35865 a_n1699_43638# a_n1917_43396# 0.209641f
C35866 a_n2129_43609# a_n1352_43396# 0.041828f
C35867 a_n2433_43396# a_n447_43370# 1.32e-20
C35868 a_15493_43396# a_14955_43396# 0.076347f
C35869 a_n2810_45028# a_n3565_39590# 0.021277f
C35870 a_n443_42852# VDD 3.69394f
C35871 a_n2438_43548# a_458_43396# 8.26e-20
C35872 a_13527_45546# a_9482_43914# 7.42e-19
C35873 a_13163_45724# a_13556_45296# 0.001027f
C35874 a_11823_42460# a_14180_45002# 6.93e-21
C35875 a_2324_44458# a_9159_44484# 1.37e-20
C35876 a_n1613_43370# a_7274_43762# 2.77e-19
C35877 a_8192_45572# a_3232_43370# 5.95e-19
C35878 a_8120_45572# a_6171_45002# 6.76e-19
C35879 a_16327_47482# a_17324_43396# 0.216094f
C35880 a_n2497_47436# a_685_42968# 9.26e-22
C35881 a_2711_45572# a_8488_45348# 5.77e-19
C35882 a_9290_44172# a_11541_44484# 0.001162f
C35883 a_10227_46804# a_16547_43609# 8.56e-19
C35884 a_3090_45724# a_15682_43940# 0.001971f
C35885 a_14976_45028# a_14955_43940# 2.22e-19
C35886 a_11453_44696# a_10341_43396# 1.84e-21
C35887 a_768_44030# a_7112_43396# 4.37e-21
C35888 a_n2293_46634# a_4235_43370# 0.012147f
C35889 a_7499_43078# a_1423_45028# 0.020575f
C35890 a_4791_45118# a_4361_42308# 0.111224f
C35891 C10_P_btm C2_P_btm 0.215144f
C35892 VDAC_P VCM 10.716001f
C35893 C7_P_btm C5_P_btm 0.15419f
C35894 C9_P_btm C3_P_btm 0.138859f
C35895 C8_P_btm C4_P_btm 0.149948f
C35896 EN_VIN_BSTR_N C0_N_btm 0.12803f
C35897 a_22705_38406# VDD 0.085998f
C35898 a_4883_46098# a_14976_45028# 0.019383f
C35899 a_13507_46334# a_15559_46634# 0.216791f
C35900 a_18597_46090# a_19466_46812# 0.074092f
C35901 a_10227_46804# a_12156_46660# 0.025653f
C35902 a_2107_46812# a_n2661_46098# 0.037509f
C35903 a_1983_46706# a_1799_45572# 0.089984f
C35904 a_n2661_46634# a_4651_46660# 0.020633f
C35905 a_n2293_46634# a_3221_46660# 2.47e-21
C35906 a_11309_47204# a_10467_46802# 0.023291f
C35907 a_9804_47204# a_10249_46116# 0.034717f
C35908 a_8128_46384# a_6755_46942# 0.01823f
C35909 a_13381_47204# a_13059_46348# 3.39e-21
C35910 a_12861_44030# a_14543_46987# 6.49e-19
C35911 a_19386_47436# a_19333_46634# 0.001224f
C35912 a_11599_46634# a_14035_46660# 0.021792f
C35913 a_n743_46660# a_1057_46660# 9.22e-19
C35914 a_5807_45002# a_5263_46660# 1.75e-19
C35915 a_n2497_47436# a_n1991_46122# 0.037858f
C35916 a_6851_47204# a_765_45546# 0.006814f
C35917 a_12465_44636# a_15009_46634# 2.01e-20
C35918 a_n1613_43370# a_6086_46660# 0.001965f
C35919 SMPL_ON_P a_n2840_46090# 7.81e-19
C35920 a_n2109_47186# a_n2157_46122# 1.26e-21
C35921 a_n1925_46634# a_2162_46660# 4.85e-19
C35922 a_1123_46634# a_2609_46660# 3.37e-20
C35923 a_948_46660# a_2443_46660# 4.94e-20
C35924 a_10341_43396# a_17364_32525# 5.25e-19
C35925 a_375_42282# VDD 0.591443f
C35926 a_3626_43646# a_10922_42852# 4.54e-20
C35927 a_2982_43646# a_12379_42858# 1.63e-19
C35928 a_3080_42308# a_5534_30871# 0.019853f
C35929 a_7287_43370# a_7227_42852# 0.008095f
C35930 a_n2661_42282# a_1067_42314# 8.97e-20
C35931 a_16759_43396# a_16823_43084# 0.038761f
C35932 a_16137_43396# a_4190_30871# 0.113768f
C35933 a_16977_43638# a_17433_43396# 4.2e-19
C35934 a_19862_44208# a_22400_42852# 5.55e-21
C35935 a_2813_43396# a_1847_42826# 2.9e-19
C35936 a_19692_46634# a_20301_43646# 0.110092f
C35937 a_2711_45572# a_1414_42308# 1.75e-21
C35938 a_n863_45724# a_3499_42826# 9.47e-19
C35939 a_n745_45366# a_n452_44636# 0.001046f
C35940 a_n913_45002# a_742_44458# 0.302053f
C35941 a_n1059_45260# a_949_44458# 2.96e-19
C35942 a_15595_45028# a_15685_45394# 0.004764f
C35943 a_14537_43396# a_14309_45028# 0.006215f
C35944 a_n2293_45010# a_n699_43396# 0.005002f
C35945 a_n467_45028# a_n2433_44484# 2.79e-19
C35946 a_n143_45144# a_n2661_44458# 4.34e-20
C35947 a_n443_42852# a_5495_43940# 1.65e-21
C35948 a_13249_42308# a_11967_42832# 0.023012f
C35949 a_4791_45118# a_6761_42308# 0.001495f
C35950 a_13507_46334# a_20009_46494# 1.94e-19
C35951 a_5907_46634# a_6165_46155# 0.003895f
C35952 a_n443_46116# a_n89_45572# 0.006092f
C35953 a_n1151_42308# a_3175_45822# 2.87e-20
C35954 a_n881_46662# a_8062_46155# 1.93e-19
C35955 a_15227_44166# a_20107_46660# 4.52e-19
C35956 a_18834_46812# a_20411_46873# 4.86e-22
C35957 a_14180_46812# a_14543_46987# 0.005265f
C35958 a_19333_46634# a_19551_46910# 0.08213f
C35959 a_13885_46660# a_15227_46910# 1.69e-19
C35960 a_17609_46634# a_20273_46660# 3.59e-21
C35961 a_n743_46660# a_6945_45028# 0.029165f
C35962 a_9804_47204# a_8781_46436# 1.48e-20
C35963 a_8128_46384# a_8049_45260# 0.00208f
C35964 a_4883_46098# a_18051_46116# 0.003099f
C35965 a_18479_47436# a_20850_46155# 0.003424f
C35966 a_19692_46634# a_18285_46348# 5.98e-20
C35967 a_19466_46812# a_19123_46287# 0.007907f
C35968 a_4646_46812# a_5937_45572# 0.105447f
C35969 a_n237_47217# a_2211_45572# 0.005215f
C35970 a_2063_45854# a_6472_45840# 0.545607f
C35971 a_n2104_46634# a_n2956_39304# 6.41e-19
C35972 a_n2293_46634# a_n2956_38680# 1.99e-19
C35973 a_743_42282# a_n473_42460# 1.85e-19
C35974 a_22165_42308# a_22223_42860# 0.171681f
C35975 a_8873_43396# a_5934_30871# 4.31e-21
C35976 a_n4318_39304# a_n3420_39616# 0.256393f
C35977 a_3626_43646# a_17531_42308# 0.003944f
C35978 a_4190_30871# a_n784_42308# 0.019472f
C35979 a_14209_32519# a_22765_42852# 4.61e-20
C35980 a_8952_43230# a_9114_42852# 0.006453f
C35981 a_2982_43646# a_18727_42674# 1.36e-19
C35982 a_3422_30871# C7_N_btm 2.94e-19
C35983 a_n1059_45260# a_11341_43940# 4.96e-19
C35984 a_n2433_44484# a_n2661_43922# 0.075698f
C35985 a_n2661_44458# a_n2293_43922# 1.21e-19
C35986 a_17613_45144# a_11967_42832# 8.83e-21
C35987 a_16922_45042# a_20159_44458# 0.012027f
C35988 a_n443_42852# a_16137_43396# 0.020044f
C35989 a_8701_44490# a_5891_43370# 0.001099f
C35990 a_18443_44721# a_18989_43940# 0.0016f
C35991 a_n2129_44697# a_n2661_42834# 0.001254f
C35992 a_742_44458# a_556_44484# 0.044092f
C35993 a_1307_43914# a_6453_43914# 0.006717f
C35994 a_5205_44484# a_6756_44260# 1.27e-19
C35995 a_n357_42282# a_16867_43762# 8.18e-21
C35996 a_526_44458# a_10991_42826# 2.56e-21
C35997 a_5111_44636# a_9672_43914# 0.001516f
C35998 a_11827_44484# a_17061_44734# 0.0048f
C35999 a_21359_45002# a_17517_44484# 9.2e-20
C36000 a_8103_44636# a_8238_44734# 0.008535f
C36001 a_3090_45724# a_5934_30871# 2.22e-20
C36002 a_22731_47423# a_413_45260# 0.005286f
C36003 a_10227_46804# a_6171_45002# 0.087616f
C36004 a_2324_44458# a_15682_46116# 0.343876f
C36005 a_4704_46090# a_526_44458# 2.04e-19
C36006 a_4419_46090# a_n1925_42282# 0.056546f
C36007 a_6755_46942# a_10053_45546# 1.29e-20
C36008 a_10467_46802# a_10490_45724# 2.95e-19
C36009 a_20411_46873# a_20850_46482# 9.61e-19
C36010 a_13747_46662# a_19418_45938# 6.02e-19
C36011 a_13661_43548# a_18787_45572# 0.001493f
C36012 a_10037_47542# a_2437_43646# 9.04e-19
C36013 a_11189_46129# a_6945_45028# 9.57e-21
C36014 a_n746_45260# a_n2293_42834# 1.39e-21
C36015 a_n443_46116# a_2304_45348# 0.008048f
C36016 a_n971_45724# a_8137_45348# 7.49e-20
C36017 a_3090_45724# a_1609_45572# 1.86e-20
C36018 a_12861_44030# a_13159_45002# 0.008506f
C36019 a_6655_43762# VDD 0.132357f
C36020 a_1606_42308# a_2713_42308# 0.002318f
C36021 a_n2293_42282# a_n2302_40160# 3.05e-20
C36022 a_n913_45002# a_n901_43156# 0.075029f
C36023 a_n1059_45260# a_n1076_43230# 0.001392f
C36024 a_n2017_45002# a_n13_43084# 8.63e-19
C36025 a_n1917_44484# a_n1699_43638# 2.44e-20
C36026 a_n1177_44458# a_n2267_43396# 2.68e-21
C36027 a_n1699_44726# a_n1917_43396# 8.81e-20
C36028 a_n863_45724# a_3318_42354# 9.94e-19
C36029 a_10554_47026# VDD 0.205847f
C36030 a_15433_44458# a_14955_43940# 0.005438f
C36031 a_5111_44636# a_743_42282# 0.024053f
C36032 a_413_45260# a_14209_32519# 3.38e-20
C36033 a_n2065_43946# a_n1549_44318# 0.110816f
C36034 a_n1761_44111# a_n1331_43914# 0.043168f
C36035 a_18184_42460# a_3626_43646# 0.052679f
C36036 a_n2661_44458# a_n97_42460# 3.24e-21
C36037 a_9313_44734# a_22959_43948# 5.71e-19
C36038 a_10193_42453# a_14635_42282# 0.00461f
C36039 a_11823_42460# a_12800_43218# 0.00522f
C36040 a_n443_42852# a_n784_42308# 0.005038f
C36041 a_n357_42282# a_n327_42308# 0.00216f
C36042 a_n755_45592# a_2351_42308# 0.057532f
C36043 en_comp a_n1853_43023# 2.91e-19
C36044 a_n967_45348# a_n2157_42858# 0.02564f
C36045 a_4883_46098# a_15433_44458# 2.94e-21
C36046 a_310_45028# a_997_45618# 3.77e-20
C36047 a_19321_45002# a_17767_44458# 1.52e-37
C36048 a_13661_43548# a_18287_44626# 0.021421f
C36049 a_13747_46662# a_18248_44752# 2.31e-20
C36050 a_14840_46494# a_8696_44636# 1.02e-21
C36051 a_15682_46116# a_16855_45546# 0.011741f
C36052 a_17715_44484# a_16333_45814# 2.81e-19
C36053 a_11415_45002# a_n913_45002# 4.59e-20
C36054 a_11453_44696# a_n2293_43922# 1.93e-20
C36055 a_10227_46804# a_14673_44172# 0.012944f
C36056 a_n2293_45546# a_n356_45724# 6.95e-20
C36057 a_8049_45260# a_10053_45546# 0.002369f
C36058 a_18189_46348# a_15765_45572# 7.83e-21
C36059 a_12861_44030# a_11967_42832# 0.209245f
C36060 a_n1613_43370# a_5891_43370# 0.064769f
C36061 a_n2312_40392# a_n2661_42834# 8.33e-20
C36062 a_n746_45260# a_1115_44172# 2.04e-19
C36063 a_584_46384# a_n2065_43946# 2.03e-21
C36064 a_3090_45724# a_4185_45348# 1.98e-19
C36065 a_10903_43370# a_13385_45572# 0.006432f
C36066 a_13885_46660# a_9482_43914# 3.2e-20
C36067 a_n2293_46634# a_10334_44484# 2.78e-20
C36068 a_n2661_46634# a_8975_43940# 1.39e-19
C36069 a_n863_45724# a_3316_45546# 8.84e-21
C36070 a_n357_42282# a_n755_45592# 0.664842f
C36071 a_n4315_30879# a_n2946_39866# 4.06e-20
C36072 a_5742_30871# VDAC_Pi 1.57e-19
C36073 a_n4064_40160# a_n3690_39616# 2.54e-19
C36074 a_14635_42282# VDD 0.369964f
C36075 a_5934_30871# a_3754_38470# 1.86e-19
C36076 a_n2109_47186# a_n443_46116# 0.080373f
C36077 a_n1741_47186# a_4700_47436# 0.008526f
C36078 a_n237_47217# a_2905_45572# 0.025329f
C36079 a_1209_47178# a_584_46384# 0.104123f
C36080 a_n971_45724# a_n1151_42308# 0.682801f
C36081 a_375_42282# a_n784_42308# 0.004284f
C36082 a_15493_43940# a_17538_32519# 0.013565f
C36083 a_14021_43940# a_13565_43940# 0.001756f
C36084 a_22959_43948# a_20974_43370# 0.005835f
C36085 a_n913_45002# a_10533_42308# 0.246621f
C36086 a_n1059_45260# a_10723_42308# 5.28e-20
C36087 a_n2017_45002# a_11323_42473# 0.003882f
C36088 a_3499_42826# a_3540_43646# 0.007239f
C36089 a_3905_42865# a_3457_43396# 5.36e-20
C36090 a_20692_30879# a_22609_37990# 1.07e-20
C36091 a_11967_42832# a_19700_43370# 1.03e-21
C36092 a_n2661_42834# a_n2840_42826# 0.174935f
C36093 a_n356_44636# a_7871_42858# 2.26e-20
C36094 a_6633_46155# VDD 6.34e-20
C36095 a_3537_45260# a_6773_42558# 0.001736f
C36096 a_5111_44636# a_5755_42308# 6.35e-19
C36097 a_3483_46348# a_18374_44850# 1.41e-21
C36098 a_16855_45546# a_16680_45572# 0.233657f
C36099 a_16115_45572# a_8696_44636# 7.81e-20
C36100 a_10193_42453# a_2437_43646# 2.74e-20
C36101 a_8199_44636# a_8975_43940# 0.028334f
C36102 a_1823_45246# a_n356_44636# 4.79e-19
C36103 a_15599_45572# a_16223_45938# 9.73e-19
C36104 a_15903_45785# a_16020_45572# 0.157972f
C36105 a_15765_45572# a_17478_45572# 2.62e-19
C36106 a_2063_45854# a_10695_43548# 3.18e-19
C36107 CAL_N a_22521_40599# 0.006786f
C36108 a_n3565_38502# VREF_GND 0.001993f
C36109 a_n1435_47204# a_7715_46873# 8.51e-20
C36110 a_6151_47436# a_6755_46942# 0.361724f
C36111 a_9313_45822# a_7927_46660# 9.18e-20
C36112 a_n881_46662# a_n1925_46634# 0.467945f
C36113 a_n1613_43370# a_n1021_46688# 0.006304f
C36114 a_2747_46873# a_1983_46706# 3.11e-19
C36115 a_n3565_37414# a_n1838_35608# 1.2e-19
C36116 a_n4209_37414# a_n1532_35090# 8.48e-20
C36117 a_n3420_37984# VDD 0.930532f
C36118 a_14021_43940# a_5534_30871# 1.65e-19
C36119 a_n1699_43638# a_n1853_43023# 7.66e-20
C36120 a_n2267_43396# a_n1991_42858# 3.69e-20
C36121 a_n1917_43396# a_n2157_42858# 1.43e-19
C36122 a_n2433_43396# a_n1641_43230# 0.001096f
C36123 a_n2129_43609# a_n1423_42826# 1.14e-19
C36124 a_4235_43370# a_743_42282# 1.55e-19
C36125 a_19963_31679# C7_N_btm 1.43e-20
C36126 a_11341_43940# a_19987_42826# 1.11e-19
C36127 a_21115_43940# a_20922_43172# 6.4e-20
C36128 a_15493_43940# a_19339_43156# 2.37e-20
C36129 a_3080_42308# a_4190_30871# 0.01835f
C36130 a_n2293_43922# a_8325_42308# 4.97e-20
C36131 a_2437_43646# VDD 1.17411f
C36132 a_14579_43548# a_14205_43396# 0.066243f
C36133 a_9145_43396# a_10341_43396# 0.085699f
C36134 a_9803_43646# a_9885_43646# 0.171361f
C36135 a_8685_43396# a_8945_43396# 3.33e-19
C36136 a_19479_31679# C10_N_btm 2.25e-20
C36137 a_20447_31679# C5_N_btm 0.040445f
C36138 a_3422_30871# COMP_P 0.208163f
C36139 a_9313_44734# a_11551_42558# 8.33e-20
C36140 SMPL_ON_P a_n2104_42282# 5.11e-20
C36141 a_21076_30879# a_14401_32519# 0.057698f
C36142 a_768_44030# a_12545_42858# 2.24e-19
C36143 a_11963_45334# a_13017_45260# 3.97e-20
C36144 a_4558_45348# a_1423_45028# 1.71e-19
C36145 a_6171_45002# a_1307_43914# 0.037515f
C36146 a_n2312_40392# a_n2293_42282# 0.001844f
C36147 a_10809_44734# a_10949_43914# 0.002017f
C36148 a_18341_45572# a_19113_45348# 5.8e-19
C36149 a_18479_45785# a_11691_44458# 0.025645f
C36150 a_16147_45260# a_16237_45028# 0.005426f
C36151 a_19431_45546# a_11827_44484# 1.24e-20
C36152 a_17715_44484# a_15493_43396# 3.2e-19
C36153 a_8162_45546# a_8375_44464# 1.5e-21
C36154 a_n1151_42308# a_12005_46436# 1.31e-20
C36155 a_2063_45854# a_11315_46155# 2.18e-19
C36156 a_n1613_43370# a_9290_44172# 0.003987f
C36157 a_11453_44696# a_17957_46116# 0.0084f
C36158 a_13507_46334# a_21137_46414# 0.007257f
C36159 a_21177_47436# a_6945_45028# 0.008435f
C36160 a_20894_47436# a_10809_44734# 0.003478f
C36161 a_n2438_43548# a_n2840_46090# 0.002055f
C36162 a_n2312_38680# a_n1853_46287# 3.4e-19
C36163 a_n2661_46634# a_n1076_46494# 1.61e-20
C36164 a_10467_46802# a_12156_46660# 3.88e-21
C36165 a_9804_47204# a_5937_45572# 5.55e-20
C36166 a_11186_47026# a_11813_46116# 2.23e-20
C36167 a_8128_46384# a_8953_45546# 5.55e-20
C36168 a_12465_44636# a_19335_46494# 6.74e-21
C36169 a_n1021_46688# a_n2293_46098# 6.25e-19
C36170 a_n1925_46634# a_n2157_46122# 0.00977f
C36171 a_n2104_46634# a_n1991_46122# 2.68e-19
C36172 a_4883_46098# a_19900_46494# 0.008904f
C36173 a_4651_46660# a_765_45546# 0.004164f
C36174 a_6151_47436# a_8049_45260# 1.58e-19
C36175 a_14021_43940# a_19647_42308# 1.51e-21
C36176 a_n97_42460# a_8325_42308# 3e-19
C36177 a_4181_44734# VDD 0.004392f
C36178 a_4905_42826# a_4921_42308# 0.046918f
C36179 a_3539_42460# a_2713_42308# 8.99e-20
C36180 a_2982_43646# a_3823_42558# 0.006269f
C36181 a_9127_43156# a_10835_43094# 4.52e-21
C36182 a_8952_43230# a_10518_42984# 0.002305f
C36183 a_15227_44166# a_17141_43172# 4.12e-20
C36184 a_18587_45118# a_18287_44626# 3.25e-20
C36185 a_18911_45144# a_18248_44752# 3.13e-19
C36186 a_18315_45260# a_18443_44721# 4.68e-19
C36187 a_11827_44484# a_13076_44458# 0.007928f
C36188 a_11691_44458# a_10057_43914# 1.34e-20
C36189 a_13556_45296# a_16335_44484# 1.13e-19
C36190 a_4185_45028# a_9127_43156# 9.18e-20
C36191 a_20202_43084# a_21356_42826# 0.011854f
C36192 a_10193_42453# a_11257_43940# 2.15e-19
C36193 a_n357_42282# a_548_43396# 0.001387f
C36194 a_n2433_44484# a_n452_44636# 1.17e-20
C36195 a_n2661_44458# a_742_44458# 0.026794f
C36196 a_n2661_43370# a_7640_43914# 1.31e-19
C36197 a_413_45260# a_17730_32519# 0.026007f
C36198 a_n967_45348# a_n1761_44111# 0.015839f
C36199 a_n2661_45010# a_453_43940# 0.004674f
C36200 a_3357_43084# a_3905_42865# 0.125186f
C36201 a_n2293_45010# a_1467_44172# 1.84e-19
C36202 a_n745_45366# a_n809_44244# 1.57e-19
C36203 a_n913_45002# a_n984_44318# 0.013973f
C36204 a_15861_45028# a_15493_43396# 1.31e-20
C36205 a_14537_43396# a_15146_44484# 0.002264f
C36206 a_1307_43914# a_14673_44172# 0.012594f
C36207 a_n2129_44697# a_n1352_44484# 0.048248f
C36208 a_n1699_44726# a_n1917_44484# 0.209641f
C36209 a_n2267_44484# a_n1177_44458# 0.042415f
C36210 a_n443_42852# a_3080_42308# 0.029846f
C36211 a_4646_46812# a_n443_42852# 0.038263f
C36212 a_12549_44172# a_10907_45822# 9.26e-20
C36213 a_5815_47464# a_3357_43084# 0.029103f
C36214 a_2959_46660# a_2711_45572# 2.89e-21
C36215 a_n743_46660# a_6812_45938# 0.002228f
C36216 a_5807_45002# a_13249_42308# 0.725941f
C36217 a_13747_46662# a_13527_45546# 5.21e-20
C36218 a_13661_43548# a_13904_45546# 9.04e-21
C36219 a_11415_45002# a_14493_46090# 2.96e-20
C36220 a_12741_44636# a_13351_46090# 5.89e-22
C36221 a_20623_46660# a_21137_46414# 0.001102f
C36222 a_19466_46812# a_8049_45260# 0.061209f
C36223 a_20841_46902# a_6945_45028# 0.013693f
C36224 a_20411_46873# a_10809_44734# 0.010692f
C36225 a_6491_46660# a_2437_43646# 0.002468f
C36226 a_11599_46634# a_19418_45938# 1.59e-19
C36227 a_n1925_46634# a_8162_45546# 0.104508f
C36228 a_n2661_46634# a_10193_42453# 0.351509f
C36229 a_1823_45246# a_5204_45822# 1.73e-19
C36230 a_n2109_47186# a_3537_45260# 5.89e-19
C36231 a_18780_47178# a_18175_45572# 2.7e-19
C36232 a_18479_47436# a_18479_45785# 2.68e-19
C36233 a_16327_47482# a_18799_45938# 0.013823f
C36234 a_n1151_42308# a_n2293_45010# 0.020357f
C36235 a_n746_45260# a_413_45260# 0.031693f
C36236 a_3147_46376# a_3699_46348# 0.001175f
C36237 a_14635_42282# a_n784_42308# 2.26e-20
C36238 a_5342_30871# a_15051_42282# 0.029795f
C36239 a_15567_42826# a_14113_42308# 1.63e-20
C36240 a_5193_42852# a_5267_42460# 3.13e-19
C36241 a_5193_43172# a_5932_42308# 1.9e-21
C36242 a_11257_43940# VDD 9.66e-19
C36243 a_4185_45028# a_17124_42282# 1.64e-19
C36244 a_11827_44484# a_15301_44260# 4.18e-19
C36245 a_n2661_46634# VDD 2.23057f
C36246 a_n2661_42834# a_n2472_43914# 0.012267f
C36247 a_10193_42453# a_14543_43071# 1.03e-21
C36248 a_n1059_45260# a_10341_43396# 0.037338f
C36249 a_17517_44484# a_19279_43940# 0.020718f
C36250 a_n2661_43922# a_n2840_43914# 0.171265f
C36251 a_7229_43940# a_7287_43370# 8.37e-20
C36252 a_18479_45785# a_4190_30871# 0.123942f
C36253 a_n443_42852# a_7309_43172# 0.00116f
C36254 a_526_44458# a_2713_42308# 6.21e-21
C36255 a_10903_43370# a_12563_42308# 0.002814f
C36256 a_11691_44458# a_14021_43940# 3.38e-19
C36257 a_526_44458# a_2957_45546# 1.97e-19
C36258 a_2324_44458# a_6598_45938# 2.88e-20
C36259 a_n2312_38680# a_n2661_43370# 1.32e-20
C36260 a_13661_43548# a_17023_45118# 1.73e-20
C36261 a_13747_46662# a_16922_45042# 0.00477f
C36262 a_19333_46634# a_3357_43084# 2.08e-20
C36263 a_19692_46634# a_22223_45572# 1.03e-19
C36264 a_4883_46098# a_5343_44458# 6.41e-22
C36265 a_16327_47482# a_16112_44458# 3.69e-19
C36266 a_8199_44636# a_10193_42453# 0.236934f
C36267 a_5937_45572# a_10180_45724# 8.62e-20
C36268 a_3483_46348# a_14495_45572# 9.37e-21
C36269 a_8016_46348# a_10490_45724# 2.74e-21
C36270 a_12891_46348# a_11827_44484# 0.020579f
C36271 a_10467_46802# a_6171_45002# 4.36e-22
C36272 a_12549_44172# a_21359_45002# 9.07e-19
C36273 a_12861_44030# a_18989_43940# 0.047422f
C36274 a_18285_46348# a_18175_45572# 0.010439f
C36275 a_10227_46804# a_12607_44458# 3.68e-19
C36276 a_11599_46634# a_18248_44752# 2.26e-19
C36277 a_8049_45260# a_20205_31679# 0.301209f
C36278 a_5807_45002# a_17613_45144# 8.23e-21
C36279 a_9625_46129# a_9049_44484# 0.00226f
C36280 a_4791_45118# a_5891_43370# 0.066388f
C36281 a_11415_45002# a_15903_45785# 0.02962f
C36282 a_6123_31319# a_1736_39587# 1.03e-19
C36283 a_n1630_35242# a_n4209_38216# 2.41e-19
C36284 a_5342_30871# C9_N_btm 5.28e-19
C36285 a_n3674_37592# a_n3565_38216# 1.57e-19
C36286 a_16522_42674# a_4958_30871# 0.020415f
C36287 a_14543_43071# VDD 0.18866f
C36288 a_n784_42308# a_n3420_37984# 0.009139f
C36289 a_n2661_42834# a_10695_43548# 2.95e-20
C36290 a_n2810_45572# a_n4334_38304# 3.54e-20
C36291 a_19963_31679# COMP_P 2.93e-20
C36292 a_18326_43940# a_11341_43940# 0.003644f
C36293 a_n2661_44458# a_n901_43156# 5.46e-22
C36294 a_n2661_43922# a_9803_43646# 1.71e-20
C36295 a_n2293_43922# a_9145_43396# 0.019866f
C36296 a_10193_42453# a_19511_42282# 0.133376f
C36297 a_n2017_45002# a_20753_42852# 3.3e-20
C36298 a_n1917_44484# a_n2157_42858# 1.66e-21
C36299 a_19862_44208# a_20269_44172# 0.049487f
C36300 a_14539_43914# a_17486_43762# 1.39e-19
C36301 a_5343_44458# a_5649_42852# 3.17e-20
C36302 a_n356_44636# a_17324_43396# 2.85e-21
C36303 a_n1331_43914# a_n2267_43396# 0.001024f
C36304 a_n1549_44318# a_n2129_43609# 1.85e-20
C36305 a_n2065_43946# a_n1177_43370# 2.42e-19
C36306 a_n1761_44111# a_n1917_43396# 2.84e-19
C36307 a_n1899_43946# a_n1699_43638# 2.25e-19
C36308 a_8199_44636# VDD 1.43837f
C36309 a_10949_43914# a_12495_44260# 0.002649f
C36310 a_17973_43940# a_15493_43940# 0.028173f
C36311 a_526_44458# a_9482_43914# 0.001072f
C36312 a_10490_45724# a_11682_45822# 0.014138f
C36313 a_768_44030# a_6101_44260# 4.28e-19
C36314 a_13259_45724# a_n913_45002# 0.142601f
C36315 a_20205_31679# a_19479_31679# 0.06173f
C36316 a_4883_46098# a_9801_44260# 1.5e-19
C36317 a_18479_47436# a_14021_43940# 1.76e-19
C36318 a_5066_45546# a_8191_45002# 7.35e-19
C36319 a_11525_45546# a_10907_45822# 4.14e-19
C36320 a_8049_45260# a_5111_44636# 0.00103f
C36321 a_9049_44484# a_9159_45572# 0.007938f
C36322 a_11415_45002# a_n2661_44458# 2.26e-19
C36323 a_n2293_46634# a_3905_42865# 0.039006f
C36324 a_10227_46804# a_14761_44260# 6.06e-20
C36325 a_584_46384# a_n2129_43609# 6.92e-20
C36326 a_n971_45724# a_n1809_43762# 8.16e-19
C36327 a_8034_45724# a_6171_45002# 0.002969f
C36328 a_7174_31319# C7_N_btm 9.97e-20
C36329 a_n4064_40160# C3_P_btm 1.27e-19
C36330 a_n4064_38528# VDAC_P 2.4e-19
C36331 a_584_46384# a_288_46660# 1.99e-21
C36332 a_7754_39964# VDAC_Ni 0.207118f
C36333 a_7754_40130# a_3754_38470# 0.191861f
C36334 a_n3565_39590# C9_P_btm 0.001137f
C36335 a_16241_47178# a_16119_47582# 3.16e-19
C36336 a_16763_47508# a_12549_44172# 2.49e-19
C36337 a_16327_47482# a_15928_47570# 0.001167f
C36338 a_2063_45854# a_1983_46706# 0.001595f
C36339 a_n1151_42308# a_601_46902# 0.001897f
C36340 a_2553_47502# a_2107_46812# 1.02e-21
C36341 a_n443_46116# a_n1925_46634# 0.080855f
C36342 a_n237_47217# a_2443_46660# 6.7e-20
C36343 a_n971_45724# a_3177_46902# 0.001193f
C36344 a_6491_46660# a_n2661_46634# 0.013828f
C36345 a_13717_47436# a_13661_43548# 2.13e-20
C36346 a_12861_44030# a_5807_45002# 0.214011f
C36347 a_n4209_39304# a_n1838_35608# 2.06e-19
C36348 a_10227_46804# a_11117_47542# 5.57e-20
C36349 a_19511_42282# VDD 0.244902f
C36350 a_n3565_38216# a_n2216_37690# 1e-19
C36351 a_n4064_37984# a_n2946_37690# 3.78e-20
C36352 a_n2946_37984# a_n4064_37440# 3.78e-20
C36353 VDAC_Pi a_7754_38636# 1.59e-19
C36354 a_5883_43914# a_6481_42558# 9.74e-21
C36355 a_n97_42460# a_9145_43396# 4.77e-19
C36356 a_20935_43940# a_20749_43396# 1.23e-20
C36357 a_3626_43646# a_6293_42852# 6.33e-20
C36358 a_4093_43548# a_3457_43396# 7.01e-20
C36359 a_n356_44636# a_1184_42692# 0.03675f
C36360 a_5343_44458# a_7963_42308# 0.108654f
C36361 a_8192_45572# VDD 0.004463f
C36362 a_15493_43940# a_22591_43396# 1.85e-20
C36363 a_n2661_42282# a_5111_42852# 4.21e-20
C36364 a_14021_43940# a_4190_30871# 0.086029f
C36365 a_2711_45572# a_n699_43396# 1.83e-20
C36366 a_n2293_45546# a_n356_44636# 1.65e-19
C36367 a_12549_44172# a_16823_43084# 8.9e-20
C36368 a_4646_46812# a_6655_43762# 8.82e-19
C36369 a_1823_45246# a_3820_44260# 7.74e-19
C36370 a_12741_44636# a_17973_43940# 1.04e-20
C36371 a_13747_46662# a_15743_43084# 6.22e-21
C36372 a_13661_43548# a_19268_43646# 0.136251f
C36373 a_n2312_40392# a_n1423_42826# 4.82e-21
C36374 a_n443_42852# a_10057_43914# 0.06562f
C36375 a_11322_45546# a_11827_44484# 8.07e-20
C36376 a_5937_45572# a_5013_44260# 4.74e-20
C36377 a_n913_45002# a_n467_45028# 1.15e-19
C36378 a_3357_43084# a_5147_45002# 0.09352f
C36379 a_n2293_45010# a_327_44734# 6.84e-21
C36380 a_n1059_45260# a_n143_45144# 4.32e-20
C36381 VIN_P VREF 0.775904f
C36382 a_n1435_47204# a_4419_46090# 1.69e-20
C36383 a_13487_47204# a_3483_46348# 4.28e-19
C36384 a_22731_47423# a_20820_30879# 0.001051f
C36385 a_4883_46098# a_21297_46660# 1.2e-19
C36386 a_21811_47423# a_21076_30879# 1.63e-19
C36387 a_n1151_42308# a_12594_46348# 4.07e-19
C36388 a_n743_46660# a_15559_46634# 2.71e-19
C36389 a_4915_47217# a_9823_46155# 1.19e-20
C36390 a_11453_44696# a_11415_45002# 0.123733f
C36391 SMPL_ON_N a_22591_46660# 0.011048f
C36392 a_22223_47212# a_12741_44636# 7.08e-20
C36393 a_6151_47436# a_8953_45546# 8.27e-19
C36394 a_7903_47542# a_7920_46348# 2.96e-21
C36395 a_6545_47178# a_5937_45572# 1.49e-20
C36396 a_5807_45002# a_14180_46812# 0.007999f
C36397 a_13747_46662# a_13885_46660# 0.028801f
C36398 a_13675_47204# a_13059_46348# 8.27e-20
C36399 a_n97_42460# a_19273_43230# 4.33e-20
C36400 a_19113_45348# VDD 9.31e-19
C36401 a_n2157_42858# a_n1853_43023# 0.290902f
C36402 a_n2472_42826# a_n1991_42858# 9.31e-19
C36403 a_15781_43660# a_15567_42826# 2.55e-19
C36404 a_10341_43396# a_19987_42826# 2.55e-19
C36405 a_22959_45036# RST_Z 0.001356f
C36406 a_743_42282# a_791_42968# 5.89e-19
C36407 a_14797_45144# a_15004_44636# 2.66e-19
C36408 a_1307_43914# a_12607_44458# 4.31e-20
C36409 a_14537_43396# a_16112_44458# 0.093722f
C36410 a_14180_45002# a_14539_43914# 4.34e-20
C36411 a_16922_45042# a_18911_45144# 0.042178f
C36412 a_n913_45002# a_n2661_43922# 0.024256f
C36413 a_n745_45366# a_n2661_42834# 3.35e-21
C36414 a_n1059_45260# a_n2293_43922# 0.02309f
C36415 a_10227_46804# a_15959_42545# 0.152289f
C36416 a_15227_44166# a_15567_42826# 0.075768f
C36417 a_3090_45724# a_18249_42858# 1.21e-20
C36418 a_n2312_38680# COMP_P 4.95e-19
C36419 a_n443_42852# a_14021_43940# 0.05804f
C36420 a_526_44458# a_6031_43396# 0.002054f
C36421 a_7499_43078# a_10405_44172# 0.132405f
C36422 a_n2438_43548# a_n2104_42282# 0.009764f
C36423 a_1423_45028# a_9838_44484# 0.254741f
C36424 a_n1613_43370# a_6773_42558# 1.71e-19
C36425 a_3537_45260# a_8375_44464# 0.10437f
C36426 a_5111_44636# a_5289_44734# 0.001056f
C36427 a_5147_45002# a_5826_44734# 7.2e-19
C36428 a_20820_30879# a_14209_32519# 0.053104f
C36429 a_14311_47204# a_13249_42308# 1.62e-21
C36430 a_11735_46660# a_2324_44458# 1.17e-20
C36431 a_12861_44030# a_15143_45578# 4.39e-20
C36432 a_21363_46634# a_21542_46660# 0.007399f
C36433 a_20731_47026# a_12741_44636# 8.49e-19
C36434 a_5072_46660# a_5066_45546# 3.51e-21
C36435 a_21188_46660# a_21297_46660# 0.007416f
C36436 a_3090_45724# a_10903_43370# 0.031245f
C36437 a_10227_46804# a_8746_45002# 0.117547f
C36438 a_11599_46634# a_13527_45546# 5.7e-19
C36439 a_4883_46098# a_4880_45572# 7.06e-20
C36440 a_743_42282# a_15051_42282# 0.011096f
C36441 a_16137_43396# a_19511_42282# 0.002509f
C36442 a_21195_42852# a_14097_32519# 2.56e-20
C36443 a_21671_42860# a_22400_42852# 8.4e-20
C36444 a_5649_42852# a_12563_42308# 1.31e-19
C36445 a_4190_30871# a_15764_42576# 9.01e-20
C36446 a_19164_43230# a_20753_42852# 9.53e-20
C36447 a_19987_42826# a_20356_42852# 0.014848f
C36448 a_3080_42308# a_n3420_37984# 0.002941f
C36449 a_15743_43084# a_4958_30871# 3.06e-20
C36450 a_18783_43370# a_17303_42282# 2.56e-21
C36451 a_4361_42308# a_14456_42282# 0.007582f
C36452 a_n2661_44458# a_n984_44318# 1.3e-20
C36453 a_3357_43084# a_4093_43548# 0.031759f
C36454 a_18143_47464# VDD 0.388551f
C36455 a_13259_45724# a_20922_43172# 7.71e-21
C36456 a_17591_47464# START 5.79e-19
C36457 a_10227_46804# RST_Z 7.13e-19
C36458 a_n967_45348# a_n2267_43396# 0.001133f
C36459 a_556_44484# a_n2661_43922# 0.00482f
C36460 a_3363_44484# a_n2661_42834# 0.003152f
C36461 a_n1917_44484# a_n1761_44111# 3.33e-19
C36462 a_n2267_44484# a_n1331_43914# 7.69e-19
C36463 a_n1177_44458# a_n2065_43946# 0.001595f
C36464 a_n1699_44726# a_n1899_43946# 1.33e-19
C36465 a_n2129_44697# a_n1549_44318# 7.49e-21
C36466 a_n443_42852# a_2075_43172# 1.18e-20
C36467 a_1823_45246# a_3823_42558# 0.137565f
C36468 a_8199_44636# a_n784_42308# 3.13e-20
C36469 a_18287_44626# a_11967_42832# 0.789765f
C36470 a_18374_44850# a_18588_44850# 0.097745f
C36471 a_18443_44721# a_19006_44850# 0.049827f
C36472 a_18248_44752# a_19615_44636# 2.73e-19
C36473 a_n1059_45260# a_n97_42460# 0.869353f
C36474 a_n2017_45002# a_104_43370# 7.08e-21
C36475 a_n2661_43370# a_10729_43914# 4.79e-19
C36476 a_4185_45028# a_1755_42282# 0.023564f
C36477 a_n357_42282# a_10083_42826# 0.017324f
C36478 a_14955_47212# CLK 3.68e-19
C36479 a_10227_46804# a_14403_45348# 1.32e-19
C36480 a_n1925_42282# a_4365_46436# 0.009374f
C36481 a_14493_46090# a_13259_45724# 7.12e-20
C36482 a_14840_46494# a_14949_46494# 0.007416f
C36483 a_15015_46420# a_15194_46482# 0.007399f
C36484 a_14275_46494# a_14383_46116# 0.057222f
C36485 a_2324_44458# a_14537_46482# 2.56e-21
C36486 a_12549_44172# a_15415_45028# 1.12e-20
C36487 a_1138_42852# a_n356_45724# 1.67e-20
C36488 a_3147_46376# a_n755_45592# 1.44e-19
C36489 a_3483_46348# a_n357_42282# 5.91e-21
C36490 a_n237_47217# a_949_44458# 0.002359f
C36491 a_584_46384# a_n2129_44697# 1.52e-20
C36492 a_765_45546# a_10193_42453# 1.36e-19
C36493 a_11599_46634# a_16922_45042# 1.05e-19
C36494 a_5807_45002# a_11787_45002# 1.03e-21
C36495 a_167_45260# a_3218_45724# 1.73e-19
C36496 a_n971_45724# a_4223_44672# 0.006952f
C36497 a_n743_46660# a_3065_45002# 4.32e-20
C36498 a_n1925_46634# a_3537_45260# 4.08e-19
C36499 a_383_46660# a_413_45260# 1.7e-20
C36500 a_601_46902# a_327_44734# 6.92e-20
C36501 a_n2293_46634# a_5147_45002# 0.009806f
C36502 a_14513_46634# a_14495_45572# 1.75e-20
C36503 a_6755_46942# a_16147_45260# 0.001071f
C36504 a_4646_46812# a_2437_43646# 9.69e-20
C36505 a_1823_45246# a_3503_45724# 0.295715f
C36506 a_12861_44030# a_18315_45260# 0.009909f
C36507 a_13678_32519# C2_N_btm 0.03058f
C36508 a_5342_30871# a_n3420_37440# 0.030303f
C36509 a_1606_42308# a_4958_30871# 0.019472f
C36510 a_21259_43561# VDD 0.192954f
C36511 a_9223_42460# a_9377_42558# 0.010303f
C36512 a_13467_32519# C5_N_btm 1.49e-19
C36513 a_5534_30871# a_n4064_37440# 0.041703f
C36514 COMP_P a_7174_31319# 0.029185f
C36515 a_11827_44484# a_16409_43396# 1.18e-21
C36516 a_22485_44484# a_22959_43948# 8.19e-19
C36517 a_7542_44172# a_n2661_42282# 1.24e-20
C36518 a_18911_45144# a_15743_43084# 1.13e-21
C36519 a_18184_42460# a_18525_43370# 6.19e-21
C36520 a_18494_42460# a_18429_43548# 2.84e-20
C36521 en_comp a_22165_42308# 4.83e-21
C36522 a_20205_31679# a_13258_32519# 0.054848f
C36523 a_765_45546# VDD 2.19953f
C36524 a_22591_44484# a_15493_43940# 2.12e-21
C36525 a_n2661_43922# a_n4318_39304# 8.01e-19
C36526 a_n2661_42834# a_n2433_43396# 0.02044f
C36527 a_5343_44458# a_8685_43396# 2.44e-19
C36528 a_n443_42852# a_15764_42576# 1.17e-20
C36529 a_1307_43914# a_3681_42891# 0.236785f
C36530 a_3175_45822# a_3260_45572# 1.48e-19
C36531 a_2711_45572# a_5024_45822# 3.69e-19
C36532 a_20916_46384# a_17517_44484# 4.81e-21
C36533 a_13351_46090# a_413_45260# 3.41e-21
C36534 a_5937_45572# a_4927_45028# 2.22e-19
C36535 a_8953_45546# a_5111_44636# 0.181796f
C36536 a_6945_45028# a_20447_31679# 5.49e-19
C36537 a_3483_46348# a_11963_45334# 0.016005f
C36538 a_13259_45724# a_15903_45785# 0.064252f
C36539 a_8016_46348# a_6171_45002# 0.022961f
C36540 a_10809_44734# a_19963_31679# 1.75e-20
C36541 a_6419_46155# a_5205_44484# 1.38e-21
C36542 a_8049_45260# a_16147_45260# 0.005281f
C36543 a_12549_44172# a_19279_43940# 0.062614f
C36544 a_19466_46812# a_20193_45348# 0.00748f
C36545 a_2107_46812# a_n2661_43922# 0.027806f
C36546 a_6511_45714# a_7227_45028# 0.213161f
C36547 a_6667_45809# a_6598_45938# 0.209641f
C36548 a_n4334_38528# a_n4064_38528# 0.449049f
C36549 a_n3690_38528# a_n3420_38528# 0.431104f
C36550 a_n3565_38502# a_n2946_38778# 0.406164f
C36551 a_n4209_38502# a_n2302_38778# 0.406492f
C36552 a_n3565_39304# a_n2302_37984# 1.31e-19
C36553 a_5934_30871# C0_N_btm 0.015126f
C36554 a_n1151_42308# a_12465_44636# 0.02014f
C36555 a_n1435_47204# a_11599_46634# 3.32e-20
C36556 a_13717_47436# a_14955_47212# 1.64e-19
C36557 a_n2109_47186# a_n1613_43370# 0.054203f
C36558 a_1209_47178# a_2266_47570# 9.52e-19
C36559 a_n971_45724# a_3315_47570# 3.15e-19
C36560 a_4921_42308# VDD 0.214995f
C36561 a_6123_31319# C2_N_btm 0.01106f
C36562 a_1606_42308# VCM 0.152876f
C36563 a_1343_38525# a_2113_38308# 0.325474f
C36564 a_5932_42308# C7_N_btm 0.003981f
C36565 a_12861_44030# a_14311_47204# 0.037394f
C36566 a_n2065_43946# a_n1991_42858# 1.27e-20
C36567 a_n1761_44111# a_n1853_43023# 0.019636f
C36568 a_n1899_43946# a_n2157_42858# 4.17e-19
C36569 a_3905_42865# a_743_42282# 3.39e-19
C36570 a_1307_43914# a_15959_42545# 1.52e-21
C36571 a_n2956_37592# a_n4209_39590# 0.090416f
C36572 a_n2433_43396# a_n1352_43396# 0.102325f
C36573 a_n2267_43396# a_n1917_43396# 0.227165f
C36574 a_n2129_43609# a_n1177_43370# 0.08445f
C36575 a_15493_43396# a_15095_43370# 1.04e-20
C36576 a_509_45822# VDD 0.190119f
C36577 a_n746_45260# a_n13_43084# 7.03e-21
C36578 a_13527_45546# a_13348_45260# 0.002161f
C36579 a_13163_45724# a_9482_43914# 8.82e-21
C36580 a_13249_42308# a_13017_45260# 1.91e-19
C36581 a_8746_45002# a_1307_43914# 9.72e-20
C36582 a_10193_42453# a_16751_45260# 0.048213f
C36583 a_16327_47482# a_17499_43370# 0.34052f
C36584 a_11823_42460# a_13777_45326# 5.57e-20
C36585 a_10227_46804# a_16243_43396# 0.001446f
C36586 a_20820_30879# a_17730_32519# 0.052913f
C36587 a_3090_45724# a_14955_43940# 0.018423f
C36588 SMPL_ON_N a_10341_43396# 4.16e-20
C36589 a_768_44030# a_7287_43370# 6.62e-20
C36590 a_n2293_46634# a_4093_43548# 0.007782f
C36591 a_2711_45572# a_8137_45348# 7.99e-20
C36592 C10_P_btm C3_P_btm 0.208539f
C36593 a_13507_46334# a_15368_46634# 0.023781f
C36594 a_4883_46098# a_3090_45724# 0.052016f
C36595 a_10227_46804# a_10425_46660# 6.24e-19
C36596 a_2107_46812# a_1799_45572# 0.079386f
C36597 a_948_46660# a_n2661_46098# 0.018472f
C36598 a_n2661_46634# a_4646_46812# 0.087334f
C36599 a_11309_47204# a_10428_46928# 0.025525f
C36600 VDAC_P VREF_GND 0.327446f
C36601 a_n1435_47204# a_13693_46688# 1.97e-20
C36602 a_12861_44030# a_14226_46987# 2.1e-19
C36603 a_18479_47436# a_19692_46634# 0.078022f
C36604 a_18597_46090# a_19333_46634# 1.8e-19
C36605 a_19386_47436# a_15227_44166# 2.72e-20
C36606 a_11599_46634# a_13885_46660# 1.52e-20
C36607 C7_P_btm C6_P_btm 20.5296f
C36608 C8_P_btm C5_P_btm 0.148944f
C36609 C9_P_btm C4_P_btm 0.1579f
C36610 a_n2438_43548# a_2864_46660# 3.97e-20
C36611 EN_VIN_BSTR_N C0_dummy_N_btm 0.026355f
C36612 a_n2497_47436# a_n1853_46287# 0.029452f
C36613 a_6491_46660# a_765_45546# 0.042766f
C36614 a_12465_44636# a_14084_46812# 2.03e-19
C36615 CAL_P RST_Z 0.551895f
C36616 a_n1613_43370# a_5841_46660# 2.95e-19
C36617 a_n2109_47186# a_n2293_46098# 1.23e-19
C36618 a_n2288_47178# a_n2157_46122# 1.61e-20
C36619 a_22609_38406# VDD 0.317066f
C36620 a_n1925_46634# a_1302_46660# 1.88e-19
C36621 a_288_46660# a_479_46660# 4.61e-19
C36622 a_1123_46634# a_2443_46660# 2.91e-21
C36623 a_14311_47204# a_14180_46812# 5.09e-19
C36624 a_10341_43396# a_22959_43396# 0.001295f
C36625 a_20365_43914# a_20256_43172# 4.57e-20
C36626 a_14021_43940# a_14635_42282# 6.42e-20
C36627 a_3626_43646# a_10991_42826# 1e-19
C36628 a_2982_43646# a_10341_42308# 4.06e-20
C36629 a_n2661_42282# a_n1630_35242# 0.093522f
C36630 a_11967_42832# a_17124_42282# 0.067231f
C36631 a_16751_45260# VDD 0.121848f
C36632 a_n2293_43922# a_n4315_30879# 2.47e-20
C36633 a_16977_43638# a_16823_43084# 0.022663f
C36634 a_17324_43396# a_17486_43762# 0.006453f
C36635 a_16759_43396# a_17021_43396# 0.001705f
C36636 a_16409_43396# a_17433_43396# 2.36e-20
C36637 a_19862_44208# a_20836_43172# 8.42e-20
C36638 a_n2433_43396# a_n2293_42282# 7.51e-20
C36639 a_19692_46634# a_4190_30871# 0.013919f
C36640 a_1423_45028# a_n2661_43370# 0.027675f
C36641 a_n1059_45260# a_742_44458# 0.030569f
C36642 a_16375_45002# a_17973_43940# 8.39e-19
C36643 a_11415_45002# a_9145_43396# 8.88e-21
C36644 a_14180_45002# a_14309_45028# 0.062574f
C36645 a_n357_42282# a_261_44278# 1.78e-19
C36646 a_413_45260# a_19721_31679# 0.116395f
C36647 a_n443_42852# a_5013_44260# 6.73e-20
C36648 a_n467_45028# a_n2661_44458# 0.031118f
C36649 a_n967_45348# a_n2267_44484# 1.92e-19
C36650 a_10586_45546# a_10555_44260# 3.3e-20
C36651 a_3090_45724# a_5649_42852# 4.39e-22
C36652 w_1575_34946# a_n3420_39616# 0.036508f
C36653 a_13507_46334# a_19597_46482# 7.17e-19
C36654 a_5072_46660# a_5068_46348# 5.86e-19
C36655 a_n1151_42308# a_2711_45572# 0.039506f
C36656 a_3160_47472# a_3175_45822# 7.95e-19
C36657 a_18834_46812# a_20107_46660# 2.51e-21
C36658 a_19333_46634# a_19123_46287# 0.113955f
C36659 a_14180_46812# a_14226_46987# 0.006879f
C36660 a_13885_46660# a_13693_46688# 5.76e-19
C36661 a_15227_44166# a_19551_46910# 0.018691f
C36662 a_11453_44696# a_13259_45724# 0.251534f
C36663 a_8128_46384# a_8781_46436# 4.93e-20
C36664 a_19466_46812# a_18285_46348# 7.08e-22
C36665 a_3877_44458# a_5937_45572# 2.07e-20
C36666 a_4646_46812# a_8199_44636# 9.29e-19
C36667 a_n237_47217# a_1990_45572# 2.46e-19
C36668 a_2905_45572# a_4099_45572# 1.64e-20
C36669 a_2063_45854# a_6194_45824# 0.041827f
C36670 a_n2293_46634# a_n2956_39304# 3.78e-19
C36671 a_n2442_46660# a_n2956_38680# 0.047296f
C36672 a_3422_30871# C6_N_btm 2.2e-19
C36673 a_743_42282# a_n961_42308# 1.36e-19
C36674 a_21671_42860# a_22223_42860# 3.81e-19
C36675 a_3626_43646# a_17303_42282# 0.037411f
C36676 a_10083_42826# a_10553_43218# 0.007399f
C36677 a_2982_43646# a_18057_42282# 9.61e-20
C36678 a_3090_45724# a_7963_42308# 4e-21
C36679 a_n2017_45002# a_11341_43940# 9e-20
C36680 en_comp a_19862_44208# 4.89e-21
C36681 a_n2661_44458# a_n2661_43922# 6.64988f
C36682 a_n2433_44484# a_n2661_42834# 0.002352f
C36683 a_18287_44626# a_18989_43940# 0.193279f
C36684 a_8701_44490# a_8375_44464# 0.001158f
C36685 a_18443_44721# a_18374_44850# 0.209641f
C36686 a_1423_45028# a_2998_44172# 0.006884f
C36687 a_1307_43914# a_5663_43940# 0.11718f
C36688 a_17023_45118# a_11967_42832# 5.47e-20
C36689 a_5205_44484# a_n2661_42282# 2.56e-19
C36690 a_21101_45002# a_17517_44484# 1.93e-19
C36691 a_5111_44636# a_9028_43914# 3.72e-19
C36692 a_5883_43914# a_7640_43914# 0.003384f
C36693 a_8103_44636# a_5891_43370# 0.029956f
C36694 a_n2312_38680# a_n4209_39304# 0.062228f
C36695 a_526_44458# a_10796_42968# 1.9e-20
C36696 a_10227_46804# a_3232_43370# 0.028168f
C36697 a_14840_46494# a_15682_46116# 3.86e-19
C36698 a_n2497_47436# a_n2661_43370# 0.031125f
C36699 a_4419_46090# a_526_44458# 0.099848f
C36700 a_4185_45028# a_n1925_42282# 0.638728f
C36701 a_10623_46897# a_10193_42453# 5.98e-20
C36702 a_10428_46928# a_10490_45724# 1.87e-20
C36703 a_13747_46662# a_17668_45572# 2.27e-19
C36704 a_9804_47204# a_2437_43646# 0.005678f
C36705 a_22223_47212# a_413_45260# 0.001872f
C36706 a_4646_46812# a_8192_45572# 1.94e-19
C36707 a_n971_45724# a_n2293_42834# 0.088674f
C36708 a_6755_46942# a_9049_44484# 5.93e-20
C36709 a_14084_46812# a_2711_45572# 1.95e-20
C36710 a_17639_46660# a_13259_45724# 5.11e-19
C36711 a_12861_44030# a_13017_45260# 0.032265f
C36712 a_n443_46116# a_2232_45348# 8.27e-19
C36713 a_3699_46348# a_3873_46454# 0.006584f
C36714 a_5534_30871# a_n3420_39072# 0.339008f
C36715 a_14635_42282# a_15764_42576# 9.01e-21
C36716 a_6452_43396# VDD 0.083252f
C36717 a_4190_30871# a_n4064_37440# 0.032722f
C36718 a_n784_42308# a_4921_42308# 4.81e-20
C36719 COMP_P a_5932_42308# 0.029797f
C36720 a_1307_43914# a_16243_43396# 0.001611f
C36721 a_3065_45002# a_4361_42308# 8.6e-19
C36722 a_n1059_45260# a_n901_43156# 0.021049f
C36723 a_n2017_45002# a_n1076_43230# 0.006096f
C36724 a_n913_45002# a_n1641_43230# 3.71e-20
C36725 a_n2267_44484# a_n1917_43396# 2.3e-19
C36726 a_n1917_44484# a_n2267_43396# 5.62e-21
C36727 a_n1352_44484# a_n2433_43396# 1.79e-21
C36728 a_n863_45724# a_2903_42308# 0.007352f
C36729 a_n755_45592# a_2123_42473# 0.022891f
C36730 a_10623_46897# VDD 0.189083f
C36731 a_14815_43914# a_14955_43940# 3.05e-19
C36732 a_n1761_44111# a_n1899_43946# 0.737653f
C36733 a_n2065_43946# a_n1331_43914# 0.053479f
C36734 a_18494_42460# a_2982_43646# 8.78e-19
C36735 a_n2433_44484# a_n1352_43396# 3.97e-20
C36736 a_9313_44734# a_15493_43940# 4.02e-19
C36737 a_10193_42453# a_13291_42460# 0.050019f
C36738 a_n443_42852# a_196_42282# 3.14e-19
C36739 en_comp a_n2157_42858# 0.005749f
C36740 a_16327_47482# a_18204_44850# 1.7e-19
C36741 a_310_45028# a_n755_45592# 0.02846f
C36742 a_n1099_45572# a_997_45618# 5.02e-19
C36743 a_13661_43548# a_18248_44752# 0.019034f
C36744 a_15682_46116# a_16115_45572# 0.008647f
C36745 a_15015_46420# a_8696_44636# 5.75e-21
C36746 a_20202_43084# a_n913_45002# 0.322116f
C36747 a_11453_44696# a_n2661_43922# 0.009016f
C36748 a_10227_46804# a_14581_44484# 1.42e-20
C36749 a_n743_46660# a_6298_44484# 1.32e-20
C36750 a_8034_45724# a_8746_45002# 2.6e-20
C36751 a_1799_45572# a_n2661_44458# 3.78e-20
C36752 a_17715_44484# a_15765_45572# 4.5e-19
C36753 a_12594_46348# a_12649_45572# 2.33e-19
C36754 a_n2497_47436# a_2998_44172# 1.03e-19
C36755 a_12861_44030# a_19006_44850# 0.008813f
C36756 a_n746_45260# a_644_44056# 9.68e-19
C36757 a_3090_45724# a_3602_45348# 4.94e-19
C36758 a_10903_43370# a_13297_45572# 0.00546f
C36759 a_8049_45260# a_9049_44484# 0.002717f
C36760 a_n2293_46634# a_10157_44484# 5.67e-21
C36761 a_n4315_30879# a_n3420_39616# 0.03477f
C36762 a_n4064_40160# a_n3565_39590# 0.031111f
C36763 a_13291_42460# VDD 0.546706f
C36764 COMP_P a_22717_36887# 0.001989f
C36765 a_7174_31319# a_n4209_39304# 4.73e-21
C36766 a_n2109_47186# a_4791_45118# 0.34446f
C36767 a_n1741_47186# a_4007_47204# 0.012359f
C36768 a_1209_47178# a_2124_47436# 0.095065f
C36769 a_327_47204# a_584_46384# 6.38e-19
C36770 a_n452_47436# a_n1151_42308# 0.0065f
C36771 a_n971_45724# a_3160_47472# 0.011577f
C36772 a_1239_47204# a_1431_47204# 0.219138f
C36773 a_n357_42282# CAL_N 0.001017f
C36774 a_11967_42832# a_19268_43646# 4.72e-19
C36775 a_19615_44636# a_15743_43084# 9.04e-21
C36776 a_375_42282# a_196_42282# 0.165785f
C36777 a_15493_43940# a_20974_43370# 0.069596f
C36778 a_22959_43948# a_14401_32519# 0.006409f
C36779 a_22223_43948# a_17538_32519# 0.001143f
C36780 a_11341_43940# a_21845_43940# 4.76e-19
C36781 a_2382_45260# a_6123_31319# 9e-21
C36782 a_n1059_45260# a_10533_42308# 6.69e-21
C36783 a_n2017_45002# a_10723_42308# 0.003736f
C36784 a_n913_45002# a_10545_42558# 0.001151f
C36785 a_5066_45546# DATA[3] 7.36e-22
C36786 a_3499_42826# a_2982_43646# 0.018486f
C36787 a_7542_44172# a_7112_43396# 0.001277f
C36788 a_7845_44172# a_7287_43370# 0.011834f
C36789 a_18326_43940# a_n97_42460# 7.83e-21
C36790 a_20205_31679# a_22609_37990# 9e-21
C36791 a_6347_46155# VDD 2.18e-20
C36792 a_18479_45785# a_19511_42282# 5.07e-20
C36793 en_comp a_9803_42558# 4.34e-21
C36794 a_5111_44636# a_5421_42558# 0.003313f
C36795 a_5147_45002# a_5755_42308# 1.29e-20
C36796 a_18681_44484# a_16137_43396# 5.5e-22
C36797 a_3483_46348# a_18443_44721# 1.15e-20
C36798 a_3175_45822# a_413_45260# 0.011644f
C36799 a_16333_45814# a_8696_44636# 5.96e-20
C36800 a_16115_45572# a_16680_45572# 7.99e-20
C36801 a_15227_44166# a_20980_44850# 7.56e-21
C36802 a_768_44030# a_9420_43940# 0.001442f
C36803 a_8199_44636# a_10057_43914# 0.113262f
C36804 a_12741_44636# a_9313_44734# 1.82e-21
C36805 a_15599_45572# a_16020_45572# 0.086708f
C36806 a_15765_45572# a_15861_45028# 9.85e-20
C36807 a_1138_42852# a_n356_44636# 0.29814f
C36808 a_n3565_38502# VREF 0.056031f
C36809 a_n4209_38502# VCM 0.035344f
C36810 a_6151_47436# a_10249_46116# 0.056387f
C36811 a_9313_45822# a_8145_46902# 3.14e-19
C36812 a_n881_46662# a_n2312_38680# 4.41e-20
C36813 a_n1613_43370# a_n1925_46634# 0.33524f
C36814 a_2747_46873# a_2107_46812# 0.0019f
C36815 a_n3420_38528# VIN_P 0.053985f
C36816 a_n3690_38304# VDD 0.363068f
C36817 a_n1435_47204# a_7411_46660# 3.15e-20
C36818 a_9804_47204# a_n2661_46634# 0.02862f
C36819 a_16697_47582# a_5807_45002# 1.37e-19
C36820 a_n4209_37414# a_n1386_35608# 6.24e-22
C36821 a_14021_43940# a_14543_43071# 4.97e-20
C36822 a_n1699_43638# a_n2157_42858# 0.008327f
C36823 a_n2267_43396# a_n1853_43023# 0.003945f
C36824 a_n2433_43396# a_n1423_42826# 1.44e-19
C36825 a_n2129_43609# a_n1991_42858# 2.81e-19
C36826 a_4093_43548# a_743_42282# 4.56e-21
C36827 a_8685_43396# a_8873_43396# 0.001422f
C36828 a_19963_31679# C6_N_btm 1.26e-20
C36829 a_20935_43940# a_20922_43172# 4.63e-19
C36830 a_15493_43940# a_18599_43230# 1.61e-20
C36831 a_11341_43940# a_19164_43230# 1.25e-20
C36832 a_n4318_40392# a_n3420_39616# 4.98e-21
C36833 a_21513_45002# VDD 0.416919f
C36834 a_14579_43548# a_14358_43442# 0.142377f
C36835 a_13667_43396# a_14205_43396# 0.076384f
C36836 a_9145_43396# a_9885_43646# 0.052876f
C36837 a_19479_31679# C9_N_btm 1.91e-20
C36838 a_9313_44734# a_5742_30871# 9.25e-19
C36839 SMPL_ON_P a_n4318_38216# 0.037528f
C36840 a_5907_45546# a_n2661_43922# 2.29e-20
C36841 a_8953_45002# a_9482_43914# 0.010057f
C36842 a_12549_44172# a_12545_42858# 3.73e-20
C36843 a_n2497_47436# COMP_P 1.63e-20
C36844 a_11787_45002# a_13017_45260# 4.5e-20
C36845 a_3232_43370# a_1307_43914# 0.14252f
C36846 a_6171_45002# a_16019_45002# 0.01229f
C36847 a_10809_44734# a_10729_43914# 6.71e-21
C36848 a_18175_45572# a_11691_44458# 7.13e-20
C36849 a_18479_45785# a_19113_45348# 0.013845f
C36850 a_n2293_45010# a_n2293_42834# 0.001084f
C36851 a_2680_45002# a_2903_45348# 0.011458f
C36852 a_4574_45260# a_1423_45028# 1.58e-19
C36853 a_20820_30879# a_17538_32519# 0.052874f
C36854 a_3090_45724# a_8685_43396# 2.11639f
C36855 a_8270_45546# a_10341_43396# 5.91e-19
C36856 a_9290_44172# a_11173_44260# 0.0082f
C36857 a_9313_45822# a_5066_45546# 0.019449f
C36858 a_n881_46662# a_9823_46155# 1.37e-20
C36859 a_11453_44696# a_18189_46348# 0.534507f
C36860 a_13507_46334# a_20708_46348# 0.007683f
C36861 a_21177_47436# a_21137_46414# 1.13e-19
C36862 a_20990_47178# a_6945_45028# 0.026188f
C36863 a_19787_47423# a_10809_44734# 0.002525f
C36864 a_n2661_46634# a_n901_46420# 9.25e-21
C36865 a_10467_46802# a_10425_46660# 2.56e-19
C36866 a_9804_47204# a_8199_44636# 8.66e-19
C36867 a_11186_47026# a_11735_46660# 3.88e-21
C36868 a_8128_46384# a_5937_45572# 1.99e-19
C36869 a_12465_44636# a_19553_46090# 6.8e-21
C36870 a_4883_46098# a_20075_46420# 0.014562f
C36871 a_4646_46812# a_765_45546# 0.001856f
C36872 a_n2104_46634# a_n1853_46287# 1.31e-20
C36873 a_n2293_46634# a_n1991_46122# 0.0181f
C36874 a_n1925_46634# a_n2293_46098# 0.077794f
C36875 a_n2312_38680# a_n2157_46122# 0.001134f
C36876 a_14021_43940# a_19511_42282# 1.9e-21
C36877 a_1512_43396# a_1606_42308# 9.64e-21
C36878 a_700_44734# VDD 0.004666f
C36879 a_3626_43646# a_2713_42308# 2.32e-20
C36880 a_2982_43646# a_3318_42354# 9.73e-19
C36881 a_3080_42308# a_4921_42308# 1e-19
C36882 a_4905_42826# a_4933_42558# 4.27e-19
C36883 a_9127_43156# a_10518_42984# 6.11e-20
C36884 a_8952_43230# a_10083_42826# 6.11e-20
C36885 a_15037_43940# a_15051_42282# 2.46e-20
C36886 a_n2293_46634# a_14113_42308# 1.19e-21
C36887 a_15227_44166# a_16877_43172# 1.05e-20
C36888 a_18315_45260# a_18287_44626# 0.005579f
C36889 a_18587_45118# a_18248_44752# 6.46e-20
C36890 a_11827_44484# a_12883_44458# 0.003401f
C36891 a_11691_44458# a_10440_44484# 2.28e-20
C36892 a_13556_45296# a_16241_44484# 1.49e-19
C36893 a_4185_45028# a_8387_43230# 1.29e-20
C36894 a_20202_43084# a_20922_43172# 2.39e-19
C36895 a_13259_45724# a_9145_43396# 0.155949f
C36896 a_10193_42453# a_11173_43940# 2.8e-20
C36897 a_n357_42282# a_n144_43396# 5.4e-19
C36898 a_n2433_44484# a_n1352_44484# 0.102355f
C36899 a_n2661_44458# a_n452_44636# 0.006933f
C36900 a_n2661_43370# a_6109_44484# 1.34e-19
C36901 a_413_45260# a_22591_44484# 0.024147f
C36902 a_n967_45348# a_n2065_43946# 0.02253f
C36903 en_comp a_n1761_44111# 2.29e-21
C36904 a_n2312_39304# a_n4209_39590# 0.065703f
C36905 a_5257_43370# a_1755_42282# 2.9e-20
C36906 a_n2293_45010# a_1115_44172# 0.09282f
C36907 a_n2661_45010# a_1414_42308# 0.059385f
C36908 a_n913_45002# a_n809_44244# 0.002076f
C36909 a_n1059_45260# a_n984_44318# 0.001489f
C36910 a_8696_44636# a_15493_43396# 4.65e-20
C36911 a_n2129_44697# a_n1177_44458# 0.027646f
C36912 a_n2267_44484# a_n1917_44484# 0.212549f
C36913 a_16019_45002# a_14673_44172# 5.98e-19
C36914 a_n443_42852# a_4699_43561# 0.004673f
C36915 a_3877_44458# a_n443_42852# 2.84e-23
C36916 a_n2293_46634# a_7499_43078# 0.14773f
C36917 a_5129_47502# a_3357_43084# 0.001711f
C36918 a_11453_44696# a_17478_45572# 5.17e-21
C36919 a_13507_46334# a_13485_45572# 1.11e-19
C36920 a_18143_47464# a_18479_45785# 2.32e-21
C36921 a_5807_45002# a_13904_45546# 0.009766f
C36922 a_13747_46662# a_13163_45724# 8.69e-21
C36923 a_13661_43548# a_13527_45546# 5.13e-20
C36924 a_11415_45002# a_13925_46122# 3.85e-20
C36925 a_20841_46902# a_21137_46414# 2.33e-19
C36926 a_20623_46660# a_20708_46348# 6.62e-19
C36927 a_20273_46660# a_6945_45028# 0.02808f
C36928 a_20107_46660# a_10809_44734# 0.026612f
C36929 a_12991_46634# a_12638_46436# 2.6e-19
C36930 a_11735_46660# a_12839_46116# 3.01e-20
C36931 a_6545_47178# a_2437_43646# 0.010642f
C36932 a_12861_44030# a_20107_45572# 2.65e-22
C36933 a_11599_46634# a_17668_45572# 5.66e-19
C36934 a_18479_47436# a_18175_45572# 1.22e-21
C36935 a_16327_47482# a_18596_45572# 0.00301f
C36936 a_2063_45854# a_n913_45002# 2.32e-21
C36937 a_n746_45260# a_n37_45144# 0.031257f
C36938 a_n971_45724# a_413_45260# 0.937818f
C36939 a_3147_46376# a_3483_46348# 0.207919f
C36940 a_2698_46116# a_4185_45028# 5.29e-21
C36941 a_1823_45246# a_5164_46348# 3.04e-19
C36942 a_n2661_46634# a_10180_45724# 3.78e-20
C36943 a_13291_42460# a_n784_42308# 1.58e-20
C36944 a_5342_30871# a_14113_42308# 0.203397f
C36945 a_15279_43071# a_15051_42282# 0.006313f
C36946 a_4190_30871# a_n3420_39072# 0.10848f
C36947 a_11173_43940# VDD 0.004114f
C36948 a_18114_32519# a_15493_43940# 0.001192f
C36949 a_11827_44484# a_15037_44260# 4.08e-19
C36950 a_20820_30879# a_22465_38105# 5.82e-19
C36951 a_n2956_39768# VDD 0.697168f
C36952 a_5883_43914# a_10729_43914# 5.61e-21
C36953 a_3232_43370# a_9396_43370# 5.79e-19
C36954 a_21588_30879# SINGLE_ENDED 0.001491f
C36955 a_5807_45002# CLK 0.033646f
C36956 a_n755_45592# a_8495_42852# 0.001078f
C36957 a_9290_44172# a_14456_42282# 1.41e-20
C36958 a_n1059_45260# a_9885_43646# 7.13e-20
C36959 a_n2017_45002# a_10341_43396# 2.51e-19
C36960 a_1307_43914# a_4905_42826# 7.98e-19
C36961 a_17517_44484# a_20766_44850# 0.018462f
C36962 a_n2661_42834# a_n2840_43914# 0.014735f
C36963 a_n443_42852# a_6101_43172# 7.15e-19
C36964 a_10903_43370# a_11633_42558# 9.37e-21
C36965 a_n913_45002# a_14955_43396# 6.71e-21
C36966 a_2981_46116# a_2957_45546# 6.65e-19
C36967 a_2324_44458# a_6667_45809# 4.9e-20
C36968 a_13661_43548# a_16922_45042# 0.080391f
C36969 a_5807_45002# a_17023_45118# 1.36e-21
C36970 a_584_46384# a_3363_44484# 2.51e-20
C36971 a_19692_46634# a_2437_43646# 0.293918f
C36972 a_15227_44166# a_3357_43084# 0.026794f
C36973 a_4883_46098# a_4743_44484# 5.83e-20
C36974 a_3483_46348# a_13249_42308# 0.338396f
C36975 a_8199_44636# a_10180_45724# 0.216999f
C36976 a_8016_46348# a_8746_45002# 0.078716f
C36977 a_5937_45572# a_10053_45546# 1.28e-19
C36978 a_12549_44172# a_21101_45002# 0.00335f
C36979 a_12861_44030# a_18374_44850# 0.004423f
C36980 a_12741_44636# a_15037_45618# 1.47e-21
C36981 a_17639_46660# a_17478_45572# 2.83e-21
C36982 a_11599_46634# a_17970_44736# 1.08e-19
C36983 a_8049_45260# a_20062_46116# 1.01e-19
C36984 a_10227_46804# a_8975_43940# 0.037352f
C36985 a_17339_46660# a_18341_45572# 0.015732f
C36986 a_11415_45002# a_15599_45572# 0.007945f
C36987 a_4791_45118# a_8375_44464# 0.010645f
C36988 a_8953_45546# a_9049_44484# 0.03092f
C36989 a_7577_46660# a_8191_45002# 7.23e-22
C36990 a_6123_31319# a_1239_39587# 1.95e-19
C36991 a_5342_30871# C8_N_btm 0.093874f
C36992 a_5932_42308# a_n4209_39304# 4.36e-21
C36993 a_n3674_37592# a_n4334_38304# 7.84e-20
C36994 a_5534_30871# C10_N_btm 1.08e-19
C36995 a_16104_42674# a_4958_30871# 0.029272f
C36996 a_16522_42674# a_16269_42308# 4.61e-19
C36997 a_1606_42308# a_n4064_38528# 1.87e-20
C36998 a_13460_43230# VDD 0.276534f
C36999 a_5891_43370# a_10149_43396# 3.71e-19
C37000 a_n2810_45572# a_n4209_38216# 0.195791f
C37001 a_18079_43940# a_11341_43940# 0.00423f
C37002 a_4185_45028# EN_OFFSET_CAL 4.56e-21
C37003 a_20640_44752# a_2982_43646# 1.2e-20
C37004 a_n2661_44458# a_n1641_43230# 2.46e-22
C37005 a_n2661_42834# a_9803_43646# 5.53e-20
C37006 a_n2661_43922# a_9145_43396# 3.97e-20
C37007 a_10193_42453# a_18548_42308# 5.7e-19
C37008 a_n2017_45002# a_20356_42852# 5.14e-20
C37009 a_n2267_44484# a_n1853_43023# 7.38e-22
C37010 a_14815_43914# a_8685_43396# 3.62e-20
C37011 a_n356_44636# a_17499_43370# 2.72e-19
C37012 a_n1549_44318# a_n2433_43396# 3.69e-20
C37013 a_n1331_43914# a_n2129_43609# 3.76e-21
C37014 a_n1761_44111# a_n1699_43638# 0.003713f
C37015 a_n2065_43946# a_n1917_43396# 0.003538f
C37016 a_n1899_43946# a_n2267_43396# 1.93e-19
C37017 a_8349_46414# VDD 0.209819f
C37018 a_17737_43940# a_15493_43940# 0.037029f
C37019 a_10807_43548# a_11173_44260# 0.05223f
C37020 a_10809_44734# a_1423_45028# 3.48e-20
C37021 a_13249_42308# a_14495_45572# 0.027073f
C37022 a_n2438_43548# a_2127_44172# 1.46e-19
C37023 a_4185_45028# a_16922_45042# 9.87e-21
C37024 a_768_44030# a_5841_44260# 1.86e-19
C37025 a_13259_45724# a_n1059_45260# 0.390886f
C37026 a_11322_45546# a_10907_45822# 0.012408f
C37027 a_5066_45546# a_7705_45326# 3.84e-20
C37028 a_2711_45572# a_12649_45572# 4.51e-19
C37029 a_20205_31679# a_22223_45572# 9.5e-19
C37030 a_20692_30879# a_2437_43646# 4.72e-20
C37031 a_10227_46804# a_14485_44260# 1.37e-20
C37032 a_n746_45260# a_104_43370# 9.55e-19
C37033 a_n971_45724# a_n2012_43396# 1.54e-19
C37034 a_8034_45724# a_3232_43370# 7.93e-21
C37035 a_20820_30879# a_19721_31679# 0.052985f
C37036 a_n2293_46634# a_3600_43914# 2.97e-20
C37037 a_6545_47178# a_n2661_46634# 0.022455f
C37038 a_13717_47436# a_5807_45002# 2.74e-19
C37039 a_n3565_39590# C10_P_btm 9.75e-19
C37040 a_7174_31319# C6_N_btm 2.51e-19
C37041 a_n4064_40160# C4_P_btm 1.47e-19
C37042 a_n237_47217# a_n2661_46098# 0.01906f
C37043 a_4007_47204# a_n743_46660# 4.48e-20
C37044 a_7754_39964# a_7754_38636# 0.005394f
C37045 a_16023_47582# a_12549_44172# 7.14e-20
C37046 a_584_46384# a_1983_46706# 0.062968f
C37047 a_n1151_42308# a_33_46660# 0.005251f
C37048 a_2063_45854# a_2107_46812# 0.214026f
C37049 a_4791_45118# a_n1925_46634# 0.026798f
C37050 a_n971_45724# a_2609_46660# 0.004485f
C37051 a_15673_47210# a_16119_47582# 2.28e-19
C37052 a_n4209_39590# C8_P_btm 0.002806f
C37053 a_n4064_37984# a_n3420_37440# 0.053897f
C37054 a_n2946_37984# a_n2946_37690# 0.050477f
C37055 a_n3420_37984# a_n4064_37440# 7.43287f
C37056 a_9313_44734# a_22765_42852# 2.97e-19
C37057 a_3626_43646# a_6031_43396# 3.24e-20
C37058 a_2982_43646# a_6197_43396# 7.06e-21
C37059 a_n356_44636# a_1576_42282# 0.003861f
C37060 a_5343_44458# a_6123_31319# 0.003724f
C37061 a_8120_45572# VDD 3.83e-19
C37062 a_n2661_42282# a_4520_42826# 1.86e-20
C37063 a_14021_43940# a_21259_43561# 0.021338f
C37064 a_2711_45572# a_4223_44672# 1.51e-20
C37065 a_5937_45572# a_5244_44056# 2.04e-20
C37066 a_n2956_37592# en_comp 0.013325f
C37067 a_n2293_46634# a_15781_43660# 3.39e-19
C37068 a_22223_46124# a_3422_30871# 3.23e-21
C37069 a_4646_46812# a_6452_43396# 0.013786f
C37070 a_1823_45246# a_3499_42826# 0.003055f
C37071 a_12741_44636# a_17737_43940# 2.79e-21
C37072 a_13661_43548# a_15743_43084# 0.092364f
C37073 a_n443_42852# a_10440_44484# 1.3e-20
C37074 a_n913_45002# a_n955_45028# 6.28e-19
C37075 a_3357_43084# a_4558_45348# 2.13e-21
C37076 a_n745_45366# a_n659_45366# 0.006584f
C37077 a_n1059_45260# a_n467_45028# 0.229142f
C37078 a_n2293_45010# a_413_45260# 9.42e-22
C37079 a_5807_45002# a_14035_46660# 0.025174f
C37080 a_n2293_46634# a_15227_44166# 3.53e-19
C37081 a_12861_44030# a_3483_46348# 0.06952f
C37082 a_13507_46334# a_21542_46660# 0.001196f
C37083 a_4883_46098# a_21076_30879# 2.94e-20
C37084 a_n743_46660# a_15368_46634# 0.026392f
C37085 a_12549_44172# a_16751_46987# 3.29e-19
C37086 a_9804_47204# a_765_45546# 0.028432f
C37087 a_22731_47423# a_22591_46660# 0.011433f
C37088 a_12465_44636# a_12741_44636# 0.914049f
C37089 a_11453_44696# a_20202_43084# 0.002113f
C37090 SMPL_ON_N a_11415_45002# 4.16e-20
C37091 a_n1151_42308# a_12005_46116# 3.22e-19
C37092 a_4915_47217# a_9569_46155# 1.77e-20
C37093 a_6151_47436# a_5937_45572# 0.008183f
C37094 a_n97_42460# a_18861_43218# 0.001021f
C37095 a_22959_45036# VDD 0.30999f
C37096 a_n2472_42826# a_n1853_43023# 0.00154f
C37097 a_15681_43442# a_15567_42826# 3.35e-19
C37098 a_10341_43396# a_19164_43230# 1.41e-20
C37099 a_22223_45036# RST_Z 1.13e-19
C37100 a_n2840_42826# a_n1991_42858# 1.88e-19
C37101 a_743_42282# a_685_42968# 0.001652f
C37102 a_14537_43396# a_15004_44636# 0.047224f
C37103 a_16922_45042# a_18587_45118# 0.021516f
C37104 a_3537_45260# a_7640_43914# 0.006345f
C37105 a_n1059_45260# a_n2661_43922# 0.034597f
C37106 a_n913_45002# a_n2661_42834# 0.027216f
C37107 a_n2017_45002# a_n2293_43922# 0.654835f
C37108 a_10227_46804# a_15803_42450# 0.296174f
C37109 a_15227_44166# a_5342_30871# 0.01169f
C37110 a_n2312_38680# a_n4318_37592# 0.02327f
C37111 a_10903_43370# a_12281_43396# 1.87e-19
C37112 a_12861_44030# a_15761_42308# 2.44e-20
C37113 a_1307_43914# a_8975_43940# 0.00588f
C37114 a_526_44458# a_1512_43396# 3.44e-19
C37115 a_413_45260# a_9313_44734# 4.55e-20
C37116 a_9049_44484# a_9028_43914# 7.44e-19
C37117 a_19431_45546# a_19279_43940# 1.77e-21
C37118 a_4185_45028# a_15743_43084# 0.061074f
C37119 a_n2438_43548# a_n4318_38216# 0.00199f
C37120 a_2711_45572# a_15493_43940# 0.128282f
C37121 a_9290_44172# a_10149_43396# 4.47e-19
C37122 a_1423_45028# a_5883_43914# 0.067915f
C37123 a_17613_45144# a_17719_45144# 0.080654f
C37124 a_5111_44636# a_5205_44734# 1.91e-19
C37125 a_n2956_39768# a_n784_42308# 8.06e-21
C37126 a_20528_46660# a_12741_44636# 0.018376f
C37127 a_12861_44030# a_14495_45572# 2.03e-19
C37128 a_21188_46660# a_21076_30879# 9.43e-21
C37129 a_5257_43370# a_n1925_42282# 1.27e-20
C37130 a_10227_46804# a_10193_42453# 0.039217f
C37131 a_11599_46634# a_13163_45724# 3.12e-20
C37132 a_743_42282# a_14113_42308# 0.015227f
C37133 a_21356_42826# a_14097_32519# 2.8e-20
C37134 a_21195_42852# a_22400_42852# 4.89e-20
C37135 a_13887_32519# a_5742_30871# 0.004679f
C37136 a_4190_30871# a_15486_42560# 2.48e-19
C37137 a_16867_43762# a_17124_42282# 8.78e-22
C37138 a_19987_42826# a_20256_42852# 0.015204f
C37139 a_5111_42852# a_5379_42460# 1.62e-19
C37140 a_4361_42308# a_13575_42558# 0.006929f
C37141 a_n2433_44484# a_n1549_44318# 1.09e-19
C37142 a_n2661_44458# a_n809_44244# 8.95e-20
C37143 a_14311_47204# CLK 1.56e-19
C37144 a_7499_43078# a_743_42282# 0.087933f
C37145 a_10227_46804# VDD 2.77567f
C37146 a_13259_45724# a_19987_42826# 2.7e-20
C37147 a_19692_46634# a_19511_42282# 1.1e-20
C37148 a_17591_47464# RST_Z 2.7e-19
C37149 a_n967_45348# a_n2129_43609# 0.021282f
C37150 en_comp a_n2267_43396# 0.028399f
C37151 a_484_44484# a_n2661_43922# 6.52e-19
C37152 a_556_44484# a_n2661_42834# 2.49e-19
C37153 a_11599_46634# DATA[5] 9.31e-19
C37154 a_n1699_44726# a_n1761_44111# 0.008854f
C37155 a_n2267_44484# a_n1899_43946# 5.37e-19
C37156 a_n1917_44484# a_n2065_43946# 6.49e-19
C37157 a_n2129_44697# a_n1331_43914# 1.13e-20
C37158 a_n443_42852# a_1847_42826# 9.74e-19
C37159 a_1823_45246# a_3318_42354# 0.055532f
C37160 a_18248_44752# a_11967_42832# 0.500539f
C37161 a_18287_44626# a_19006_44850# 0.086658f
C37162 a_18443_44721# a_18588_44850# 0.057222f
C37163 a_n913_45002# a_n1352_43396# 0.002153f
C37164 a_n1059_45260# a_n447_43370# 0.018401f
C37165 a_n2017_45002# a_n97_42460# 0.169401f
C37166 a_4185_45028# a_1606_42308# 5.4e-20
C37167 a_8696_44636# a_10695_43548# 6.31e-21
C37168 a_n357_42282# a_8952_43230# 0.011989f
C37169 a_n2661_43370# a_10405_44172# 2.85e-21
C37170 a_12861_44030# a_17719_45144# 2.48e-19
C37171 a_10227_46804# a_14309_45348# 1.15e-19
C37172 a_14493_46090# a_14383_46116# 0.097745f
C37173 a_13925_46122# a_13259_45724# 0.003795f
C37174 a_12549_44172# a_14797_45144# 1.61e-20
C37175 a_768_44030# a_14537_43396# 9.19e-20
C37176 a_1176_45822# a_n356_45724# 1.67e-19
C37177 a_2804_46116# a_n755_45592# 2.12e-20
C37178 a_n971_45724# a_2779_44458# 0.009966f
C37179 a_n746_45260# a_949_44458# 0.00147f
C37180 a_n237_47217# a_742_44458# 0.002559f
C37181 a_12741_44636# a_2711_45572# 0.044854f
C37182 a_17339_46660# a_10193_42453# 0.023481f
C37183 a_n2661_46098# a_n2017_45002# 1.63e-20
C37184 a_765_45546# a_10180_45724# 2.49e-20
C37185 a_5807_45002# a_10951_45334# 1.45e-20
C37186 a_167_45260# a_2957_45546# 7.72e-19
C37187 a_n2438_43548# a_2382_45260# 4.79e-21
C37188 a_33_46660# a_327_44734# 1.67e-20
C37189 a_14180_46812# a_14495_45572# 3.41e-19
C37190 a_n881_46662# a_1423_45028# 1.63e-19
C37191 a_3877_44458# a_2437_43646# 9.39e-20
C37192 a_1823_45246# a_3316_45546# 0.099099f
C37193 a_n1925_46634# a_3429_45260# 2.79e-22
C37194 a_2063_45854# a_n2661_44458# 0.029811f
C37195 a_13059_46348# a_11823_42460# 0.256727f
C37196 a_13678_32519# C1_N_btm 1.26e-19
C37197 a_4190_30871# C10_N_btm 0.446355f
C37198 a_19177_43646# VDD 0.004534f
C37199 a_9223_42460# a_9293_42558# 0.011552f
C37200 a_13467_32519# C4_N_btm 1.74e-19
C37201 a_8515_42308# a_5742_30871# 1.16e-20
C37202 a_n2661_43922# a_n2840_43370# 3.06e-19
C37203 a_n2661_42834# a_n4318_39304# 0.041301f
C37204 a_8975_43940# a_9396_43370# 1.2e-20
C37205 a_11827_44484# a_16547_43609# 5.55e-20
C37206 a_22485_44484# a_15493_43940# 0.087012f
C37207 a_6453_43914# a_6756_44260# 0.001377f
C37208 a_7281_43914# a_n2661_42282# 8.78e-20
C37209 en_comp a_21671_42860# 4.89e-21
C37210 a_n2956_38680# a_n2946_37984# 0.004795f
C37211 a_17339_46660# VDD 0.555596f
C37212 a_n443_42852# a_15486_42560# 3.9e-21
C37213 a_n913_45002# a_n2293_42282# 0.028018f
C37214 a_1307_43914# a_2905_42968# 0.003188f
C37215 a_626_44172# a_685_42968# 9.72e-19
C37216 a_20820_30879# a_18194_35068# 1.52e-19
C37217 a_2711_45572# a_3260_45572# 3.63e-19
C37218 a_12594_46348# a_413_45260# 4.56e-21
C37219 a_5937_45572# a_5111_44636# 0.06133f
C37220 a_15227_44166# a_16237_45028# 8.33e-19
C37221 a_3483_46348# a_11787_45002# 0.019413f
C37222 a_13259_45724# a_15599_45572# 0.205417f
C37223 a_8016_46348# a_3232_43370# 0.025981f
C37224 a_7920_46348# a_6171_45002# 8.34e-21
C37225 a_6472_45840# a_7227_45028# 0.208286f
C37226 a_6511_45714# a_6598_45938# 0.06628f
C37227 a_n357_42282# a_13249_42308# 0.024753f
C37228 a_2107_46812# a_n2661_42834# 0.028012f
C37229 a_6165_46155# a_5205_44484# 3.92e-22
C37230 a_18189_46348# a_n1059_45260# 7.59e-21
C37231 a_8049_45260# a_17786_45822# 0.001566f
C37232 a_12549_44172# a_20766_44850# 1.16e-19
C37233 a_19466_46812# a_11691_44458# 0.008122f
C37234 a_3090_45724# a_18545_45144# 2.17e-19
C37235 a_5932_42308# C6_N_btm 3.73e-19
C37236 a_4958_30871# VDAC_N 0.021935f
C37237 a_5742_30871# EN_VIN_BSTR_N 0.643089f
C37238 a_1736_39043# a_2684_37794# 0.193802f
C37239 comp_n a_1177_38525# 0.003093f
C37240 a_n4209_38502# a_n4064_38528# 0.265711f
C37241 a_n3565_38502# a_n3420_38528# 0.278952f
C37242 a_n3565_39304# a_n4064_37984# 0.028081f
C37243 a_n4064_39072# a_n3565_38216# 0.030681f
C37244 a_n3420_39072# a_n3420_37984# 0.046468f
C37245 a_5934_30871# C0_dummy_N_btm 1.48e-19
C37246 a_4933_42558# VDD 0.004279f
C37247 a_6123_31319# C1_N_btm 0.011005f
C37248 a_1606_42308# VREF_GND 9e-19
C37249 a_2063_45854# a_11453_44696# 6.07e-19
C37250 a_12861_44030# a_13487_47204# 0.127147f
C37251 a_13381_47204# a_11599_46634# 2.3e-21
C37252 a_n2497_47436# a_n881_46662# 2.87e-19
C37253 a_n2109_47186# a_3411_47243# 0.001394f
C37254 a_n1741_47186# a_5063_47570# 2.13e-19
C37255 a_n746_45260# a_7_47243# 1.85e-19
C37256 a_n971_45724# a_3094_47570# 5.15e-19
C37257 a_13717_47436# a_14311_47204# 0.00371f
C37258 a_n2810_45028# a_n4209_39590# 0.021994f
C37259 a_n2065_43946# a_n1853_43023# 2.64e-21
C37260 a_n1761_44111# a_n2157_42858# 2.98e-19
C37261 a_3537_45260# a_7174_31319# 4.88e-21
C37262 a_18079_43940# a_10341_43396# 3.24e-20
C37263 a_1307_43914# a_15803_42450# 7.31e-22
C37264 a_n2956_37592# a_n2216_40160# 1.2e-19
C37265 a_n2267_43396# a_n1699_43638# 0.179796f
C37266 a_n2129_43609# a_n1917_43396# 0.036131f
C37267 a_n2433_43396# a_n1177_43370# 0.043475f
C37268 a_n4318_39304# a_n1352_43396# 4.15e-20
C37269 a_15493_43396# a_14205_43396# 5.22e-20
C37270 a_n906_45572# VDD 2.32e-19
C37271 a_11453_44696# a_14955_43396# 3.7e-22
C37272 a_n971_45724# a_n13_43084# 1.75e-19
C37273 a_n746_45260# a_n1076_43230# 8.81e-21
C37274 a_13904_45546# a_13017_45260# 1.12e-19
C37275 a_13163_45724# a_13348_45260# 8.77e-21
C37276 a_10193_42453# a_1307_43914# 0.054328f
C37277 a_2324_44458# a_5708_44484# 7.43e-19
C37278 a_11682_45822# a_3232_43370# 1.34e-19
C37279 a_3483_46348# a_17325_44484# 0.001497f
C37280 a_16327_47482# a_16759_43396# 0.152273f
C37281 a_12861_44030# a_16664_43396# 2.54e-20
C37282 a_11823_42460# a_13556_45296# 0.001625f
C37283 a_5907_45546# a_5837_45028# 9.32e-20
C37284 a_13351_46090# a_13213_44734# 1.41e-20
C37285 a_10227_46804# a_16137_43396# 0.001438f
C37286 a_20202_43084# a_19237_31679# 2.47e-20
C37287 a_3090_45724# a_13483_43940# 2.45e-20
C37288 a_18175_45572# a_2437_43646# 1.98e-21
C37289 a_19256_45572# a_19365_45572# 0.007416f
C37290 a_19431_45546# a_19610_45572# 0.007399f
C37291 a_8162_45546# a_1423_45028# 5.61e-21
C37292 a_2711_45572# a_n2293_42834# 0.002511f
C37293 a_n2956_39768# a_3080_42308# 4.45e-21
C37294 a_n2293_46634# a_1756_43548# 3.05e-19
C37295 a_768_44030# a_6547_43396# 8.31e-20
C37296 C10_P_btm C4_P_btm 0.348092f
C37297 VDAC_P VREF 0.254986f
C37298 a_948_46660# a_1799_45572# 5.85e-19
C37299 a_1123_46634# a_n2661_46098# 0.041919f
C37300 a_n2661_46634# a_3877_44458# 0.010452f
C37301 a_12861_44030# a_14513_46634# 0.036912f
C37302 a_13487_47204# a_14180_46812# 0.001914f
C37303 VDAC_N VCM 10.717099f
C37304 a_13507_46334# a_14976_45028# 0.020647f
C37305 a_18479_47436# a_19466_46812# 0.007963f
C37306 a_18597_46090# a_15227_44166# 0.150202f
C37307 C9_P_btm C5_P_btm 0.153949f
C37308 C8_P_btm C6_P_btm 0.170091f
C37309 a_n2438_43548# a_3524_46660# 7.85e-21
C37310 a_6545_47178# a_765_45546# 0.035873f
C37311 a_n881_46662# a_6682_46987# 1.68e-19
C37312 a_n2288_47178# a_n2293_46098# 1.13e-19
C37313 a_n2497_47436# a_n2157_46122# 0.034181f
C37314 CAL_P VDD 22.4716f
C37315 a_n1925_46634# a_1057_46660# 1.6e-19
C37316 a_10227_46804# a_10185_46660# 0.002879f
C37317 a_12281_43396# a_5649_42852# 1.3e-19
C37318 a_10341_43396# a_14209_32519# 0.006519f
C37319 a_15781_43660# a_743_42282# 1.91e-20
C37320 a_20269_44172# a_20256_43172# 5.7e-20
C37321 a_14021_43940# a_13291_42460# 3.77e-20
C37322 a_3626_43646# a_10796_42968# 8.42e-20
C37323 a_2982_43646# a_10922_42852# 4.62e-20
C37324 a_5013_44260# a_4921_42308# 7.51e-21
C37325 a_11967_42832# a_16522_42674# 5.62e-19
C37326 a_1307_43914# VDD 3.92807f
C37327 a_n2661_42282# a_564_42282# 2.77e-19
C37328 a_16409_43396# a_16823_43084# 0.020816f
C37329 a_16759_43396# a_16855_43396# 0.013793f
C37330 a_16977_43638# a_17021_43396# 3.69e-19
C37331 a_n97_42460# a_19164_43230# 0.005382f
C37332 a_10227_46804# a_n784_42308# 8.64e-21
C37333 a_17339_46660# a_16137_43396# 1.34e-19
C37334 a_15227_44166# a_743_42282# 3.95e-19
C37335 a_19692_46634# a_21259_43561# 0.014184f
C37336 a_n443_42852# a_5244_44056# 5.78e-21
C37337 a_16375_45002# a_17737_43940# 0.001093f
C37338 a_n913_45002# a_n1352_44484# 0.003041f
C37339 a_n1059_45260# a_n452_44636# 0.010366f
C37340 a_n745_45366# a_n1177_44458# 1.89e-21
C37341 a_n2017_45002# a_742_44458# 2.47e-19
C37342 a_1823_45246# a_6197_43396# 5.44e-21
C37343 a_6171_45002# a_11827_44484# 0.09294f
C37344 a_413_45260# a_18114_32519# 0.053981f
C37345 a_n2661_45010# a_n699_43396# 3.08e-20
C37346 a_n2810_45572# a_n2661_42282# 3.31e-20
C37347 a_310_45028# a_261_44278# 6.05e-20
C37348 a_4185_45028# a_3539_42460# 0.065262f
C37349 a_10193_42453# a_18579_44172# 0.12582f
C37350 en_comp a_n2267_44484# 0.029536f
C37351 a_n967_45348# a_n2129_44697# 0.017689f
C37352 a_n955_45028# a_n2661_44458# 2.09e-19
C37353 a_13259_45724# a_18326_43940# 8.21e-19
C37354 a_10227_46804# a_20850_46155# 2.21e-19
C37355 a_5167_46660# a_5497_46414# 0.003426f
C37356 a_2905_45572# a_3175_45822# 0.046585f
C37357 a_n443_46116# a_2307_45899# 0.001194f
C37358 a_15227_44166# a_19123_46287# 0.069758f
C37359 a_14180_46812# a_14513_46634# 0.253235f
C37360 a_13885_46660# a_14543_46987# 7.87e-19
C37361 a_14035_46660# a_14226_46987# 3.26e-19
C37362 a_12465_44636# a_16375_45002# 4.56e-21
C37363 a_12861_44030# a_n357_42282# 2.04e-19
C37364 a_4883_46098# a_19431_46494# 2.01e-19
C37365 a_2063_45854# a_5907_45546# 0.023999f
C37366 a_n2442_46660# a_n2956_39304# 0.046604f
C37367 a_n2472_46634# a_n2956_38680# 4.88e-19
C37368 a_n1925_46634# a_6945_45028# 0.028603f
C37369 a_18479_47436# a_20205_31679# 0.001643f
C37370 a_3422_30871# C5_N_btm 1.71e-19
C37371 a_21671_42860# a_22165_42308# 0.009789f
C37372 a_21195_42852# a_22223_42860# 1.88e-19
C37373 a_3626_43646# a_4958_30871# 0.087921f
C37374 a_2982_43646# a_17531_42308# 1.21e-19
C37375 a_18579_44172# VDD 0.38178f
C37376 a_13887_32519# a_22765_42852# 8.08e-19
C37377 a_3090_45724# a_6123_31319# 3.25e-20
C37378 a_n2661_44458# a_n2661_42834# 0.008313f
C37379 a_n4318_40392# a_n2661_43922# 3.97e-19
C37380 a_n2956_39768# a_n2946_39072# 0.004795f
C37381 a_18287_44626# a_18374_44850# 0.053385f
C37382 a_18248_44752# a_18989_43940# 0.207562f
C37383 a_1307_43914# a_5495_43940# 0.024105f
C37384 a_1423_45028# a_2889_44172# 4.49e-19
C37385 a_16922_45042# a_11967_42832# 0.019919f
C37386 a_21005_45260# a_17517_44484# 5.11e-20
C37387 a_11827_44484# a_14673_44172# 0.150125f
C37388 a_8746_45002# a_8791_43396# 6.27e-21
C37389 a_5111_44636# a_8333_44056# 0.280148f
C37390 a_8701_44490# a_7640_43914# 2.97e-19
C37391 a_5883_43914# a_6109_44484# 0.078113f
C37392 a_6298_44484# a_5891_43370# 1.52e-21
C37393 a_8103_44636# a_8375_44464# 0.13675f
C37394 a_526_44458# a_10835_43094# 1.38e-20
C37395 a_n357_42282# a_19700_43370# 6.27e-20
C37396 a_n2312_40392# a_n967_45348# 4.63e-20
C37397 a_n2312_39304# en_comp 0.001599f
C37398 a_14840_46494# a_2324_44458# 0.002377f
C37399 a_4185_45028# a_526_44458# 0.162857f
C37400 a_3699_46348# a_n1925_42282# 0.011511f
C37401 a_1823_45246# a_5066_45546# 5.66e-19
C37402 a_10150_46912# a_10490_45724# 5.77e-22
C37403 a_10623_46897# a_10180_45724# 5.76e-20
C37404 a_10467_46802# a_10193_42453# 5.21e-20
C37405 a_8128_46384# a_2437_43646# 0.005098f
C37406 a_12465_44636# a_413_45260# 0.28925f
C37407 a_6755_46942# a_7499_43078# 4.83e-20
C37408 a_n443_46116# a_1423_45028# 0.022652f
C37409 a_3483_46348# a_3873_46454# 6.61e-19
C37410 a_14635_42282# a_15486_42560# 0.002155f
C37411 a_9396_43370# VDD 0.288403f
C37412 a_2123_42473# a_2351_42308# 0.084895f
C37413 a_1307_43914# a_16137_43396# 4.75e-21
C37414 a_n2293_45010# a_n13_43084# 3.54e-20
C37415 a_n2017_45002# a_n901_43156# 0.005917f
C37416 a_n913_45002# a_n1423_42826# 2.51e-19
C37417 a_n1059_45260# a_n1641_43230# 1.74e-19
C37418 a_2437_43646# a_1847_42826# 1.57e-20
C37419 a_5891_43370# a_10555_44260# 0.015358f
C37420 a_n2267_44484# a_n1699_43638# 6.29e-20
C37421 a_n863_45724# a_2713_42308# 0.044499f
C37422 a_n755_45592# a_1755_42282# 1.52791f
C37423 a_n357_42282# a_2123_42473# 1.65e-20
C37424 a_10467_46802# VDD 0.401016f
C37425 a_18184_42460# a_2982_43646# 0.020575f
C37426 a_n2065_43946# a_n1899_43946# 0.614122f
C37427 a_n443_42852# a_n473_42460# 0.001248f
C37428 en_comp a_n2472_42826# 0.019667f
C37429 a_16327_47482# a_17517_44484# 0.090308f
C37430 a_n1099_45572# a_n755_45592# 0.193775f
C37431 a_310_45028# a_n357_42282# 0.113929f
C37432 a_380_45546# a_997_45618# 0.070624f
C37433 a_n2661_45546# a_n23_45546# 0.006975f
C37434 a_16375_45002# a_2711_45572# 0.00407f
C37435 a_5807_45002# a_18248_44752# 4.21e-21
C37436 a_13661_43548# a_17970_44736# 2.76e-21
C37437 a_13747_46662# a_17767_44458# 5.22e-21
C37438 a_15682_46116# a_16333_45814# 0.011944f
C37439 a_14275_46494# a_8696_44636# 9.68e-21
C37440 a_768_44030# a_n356_44636# 0.098499f
C37441 a_11453_44696# a_n2661_42834# 4.17e-19
C37442 a_10227_46804# a_13940_44484# 1.36e-20
C37443 a_n2293_45546# a_3316_45546# 1.26e-20
C37444 a_18189_46348# a_15599_45572# 2.91e-37
C37445 a_12861_44030# a_18588_44850# 0.006708f
C37446 a_12465_44636# a_13468_44734# 1.06e-20
C37447 a_n1613_43370# a_7640_43914# 2.1e-20
C37448 a_n881_46662# a_6109_44484# 0.001229f
C37449 a_n746_45260# a_175_44278# 0.159759f
C37450 a_3090_45724# a_3495_45348# 6.6e-19
C37451 a_10903_43370# a_12749_45572# 1.89e-20
C37452 a_6969_46634# a_n2661_43370# 5.75e-22
C37453 a_14035_46660# a_13017_45260# 1.07e-19
C37454 a_8049_45260# a_7499_43078# 0.00119f
C37455 a_n2293_46634# a_9838_44484# 2.45e-22
C37456 a_n1925_46634# a_8103_44636# 5.79e-21
C37457 a_13003_42852# VDD 0.132655f
C37458 a_n2302_40160# a_n4209_39590# 9.15e-19
C37459 a_n4064_40160# a_n4334_39616# 0.014656f
C37460 a_7174_31319# a_1343_38525# 2.49e-19
C37461 a_5934_30871# VDAC_Ni 3.94e-19
C37462 a_n784_42308# CAL_P 0.006719f
C37463 a_6123_31319# a_3754_38470# 2.11e-19
C37464 a_n785_47204# a_584_46384# 0.002399f
C37465 a_n2109_47186# a_4700_47436# 0.038955f
C37466 a_n1741_47186# a_3815_47204# 0.023296f
C37467 a_n237_47217# a_2553_47502# 4.45e-21
C37468 a_1209_47178# a_1431_47204# 0.095209f
C37469 a_n815_47178# a_n1151_42308# 0.011772f
C37470 a_n971_45724# a_2905_45572# 0.118495f
C37471 a_n2497_47436# a_n443_46116# 0.026321f
C37472 a_11967_42832# a_15743_43084# 0.180938f
C37473 a_13076_44458# a_12545_42858# 1.33e-20
C37474 a_375_42282# a_n473_42460# 8.64e-19
C37475 a_15493_43940# a_14401_32519# 0.052433f
C37476 a_22223_43948# a_20974_43370# 7.69e-19
C37477 a_11341_43940# a_17538_32519# 4.23e-19
C37478 a_3537_45260# a_5932_42308# 0.008724f
C37479 a_n2017_45002# a_10533_42308# 0.003333f
C37480 a_n913_45002# a_9885_42558# 0.001674f
C37481 a_n2661_42282# a_n1557_42282# 4.93e-19
C37482 a_7281_43914# a_7112_43396# 0.001258f
C37483 a_7542_44172# a_7287_43370# 0.003428f
C37484 a_1307_43914# a_n784_42308# 2.99e-19
C37485 a_18079_43940# a_n97_42460# 3.05e-20
C37486 a_8034_45724# VDD 0.812726f
C37487 en_comp a_9223_42460# 4.34e-21
C37488 a_n356_44636# a_5755_42852# 5.65e-21
C37489 a_18579_44172# a_16137_43396# 9.57e-20
C37490 a_20692_30879# a_22609_38406# 4.83e-21
C37491 a_2063_45854# a_9145_43396# 1.47e-19
C37492 a_3483_46348# a_18287_44626# 2.49e-19
C37493 a_2711_45572# a_413_45260# 0.022324f
C37494 a_16333_45814# a_16680_45572# 0.051162f
C37495 a_10053_45546# a_2437_43646# 8.54e-21
C37496 a_768_44030# a_9165_43940# 0.00651f
C37497 a_8199_44636# a_10440_44484# 8.12e-19
C37498 a_8016_46348# a_8975_43940# 0.01976f
C37499 a_n443_42852# a_5111_44636# 0.584506f
C37500 a_20820_30879# a_9313_44734# 1.42e-20
C37501 a_15903_45785# a_15861_45028# 0.232345f
C37502 a_15765_45572# a_8696_44636# 6.07e-19
C37503 a_15599_45572# a_17478_45572# 1.88e-20
C37504 a_4646_46812# a_7911_44260# 2.43e-21
C37505 a_2063_45854# a_10384_47026# 1.72e-19
C37506 a_11206_38545# CAL_N 0.050483f
C37507 a_n4209_38502# VREF_GND 0.00199f
C37508 a_4915_47217# a_6969_46634# 1.7e-19
C37509 a_6151_47436# a_10554_47026# 1.71e-19
C37510 a_9067_47204# a_8667_46634# 0.005569f
C37511 a_9313_45822# a_7577_46660# 3.38e-19
C37512 a_n1613_43370# a_n2312_38680# 4.23e-21
C37513 a_2747_46873# a_948_46660# 4.23e-19
C37514 a_n3565_38216# VDD 0.901259f
C37515 a_8128_46384# a_n2661_46634# 0.029397f
C37516 a_n1435_47204# a_5257_43370# 2.43e-20
C37517 a_n4209_37414# a_n1838_35608# 1.81e-19
C37518 a_n2433_43396# a_n1991_42858# 6.51e-19
C37519 a_n2267_43396# a_n2157_42858# 6.7e-20
C37520 a_n2129_43609# a_n1853_43023# 1.06e-19
C37521 a_9145_43396# a_14955_43396# 0.06858f
C37522 a_8685_43396# a_12281_43396# 0.038443f
C37523 a_19963_31679# C5_N_btm 1.11e-20
C37524 a_11341_43940# a_19339_43156# 1.47e-20
C37525 a_19479_31679# C8_N_btm 1.65e-20
C37526 a_14539_43914# a_17531_42308# 5.33e-20
C37527 a_9313_44734# a_11323_42473# 5.36e-20
C37528 a_13667_43396# a_14358_43442# 0.001448f
C37529 a_5907_45546# a_n2661_42834# 1.65e-20
C37530 a_11682_45822# a_8975_43940# 1.53e-20
C37531 a_768_44030# a_12379_42858# 1.38e-20
C37532 a_12891_46348# a_12545_42858# 1.12e-20
C37533 a_12549_44172# a_12089_42308# 1.47e-19
C37534 SMPL_ON_P a_n2472_42282# 2.48e-19
C37535 a_11787_45002# a_11963_45334# 0.185422f
C37536 a_5691_45260# a_1307_43914# 1.36e-19
C37537 a_6171_45002# a_15595_45028# 0.012742f
C37538 a_18175_45572# a_19113_45348# 3.29e-19
C37539 a_16147_45260# a_11691_44458# 7.44e-20
C37540 a_3357_43084# a_n2661_43370# 0.030835f
C37541 a_20273_45572# a_16922_45042# 4.48e-20
C37542 a_2680_45002# a_2809_45348# 0.010132f
C37543 a_3537_45260# a_1423_45028# 0.046355f
C37544 a_8270_45546# a_9885_43646# 0.002107f
C37545 a_6755_46942# a_15781_43660# 1.89e-20
C37546 a_9290_44172# a_10555_44260# 3.43e-21
C37547 a_n2104_46634# a_n2157_46122# 0.013135f
C37548 a_11453_44696# a_17715_44484# 0.036977f
C37549 a_13507_46334# a_19900_46494# 0.005187f
C37550 a_20894_47436# a_6945_45028# 0.016564f
C37551 a_n2661_46634# a_n1641_46494# 6.71e-19
C37552 a_10428_46928# a_10425_46660# 2.36e-20
C37553 a_9804_47204# a_8349_46414# 3.47e-20
C37554 a_10037_47542# a_8016_46348# 3.96e-20
C37555 a_6755_46942# a_15227_44166# 0.288173f
C37556 a_8128_46384# a_8199_44636# 3.12e-19
C37557 a_n881_46662# a_9569_46155# 2.93e-20
C37558 a_12465_44636# a_18985_46122# 7.56e-21
C37559 a_19386_47436# a_10809_44734# 9.09e-19
C37560 a_4883_46098# a_19335_46494# 0.007327f
C37561 a_3877_44458# a_765_45546# 0.001935f
C37562 a_n2293_46634# a_n1853_46287# 0.014216f
C37563 a_n2312_38680# a_n2293_46098# 0.003636f
C37564 a_14401_32519# a_5742_30871# 0.005978f
C37565 a_n998_44484# VDD 1.32e-19
C37566 a_2982_43646# a_2903_42308# 4.44e-21
C37567 a_4905_42826# a_3905_42558# 3.25e-20
C37568 a_9127_43156# a_10083_42826# 0.011187f
C37569 a_18315_45260# a_18248_44752# 3.25e-19
C37570 a_11691_44458# a_10334_44484# 2.3e-20
C37571 a_11827_44484# a_12607_44458# 0.023193f
C37572 a_13556_45296# a_15367_44484# 0.003919f
C37573 a_3483_46348# a_9127_43156# 0.001097f
C37574 a_4185_45028# a_8605_42826# 1.07e-20
C37575 a_20202_43084# a_19987_42826# 0.177726f
C37576 a_n2661_44458# a_n1352_44484# 0.00782f
C37577 a_16922_45042# a_18989_43940# 3.37e-19
C37578 a_n2433_44484# a_n1177_44458# 0.043567f
C37579 en_comp a_n2065_43946# 2.47e-19
C37580 a_n2312_40392# a_n4209_39590# 1.62e-19
C37581 a_3357_43084# a_2998_44172# 0.119142f
C37582 a_n2293_45010# a_644_44056# 0.014621f
C37583 a_n2017_45002# a_n984_44318# 3.14e-21
C37584 a_n2661_45010# a_1467_44172# 0.001683f
C37585 a_n1059_45260# a_n809_44244# 0.021842f
C37586 a_413_45260# a_22485_44484# 6.37e-21
C37587 a_14537_43396# a_17517_44484# 6.26e-21
C37588 a_n2129_44697# a_n1917_44484# 0.030172f
C37589 a_n2267_44484# a_n1699_44726# 0.172319f
C37590 a_15595_45028# a_14673_44172# 2.84e-20
C37591 a_n443_42852# a_4235_43370# 0.026532f
C37592 a_16327_47482# a_19256_45572# 0.235006f
C37593 a_8128_46384# a_8192_45572# 2.19e-19
C37594 a_4915_47217# a_3357_43084# 0.028255f
C37595 a_11453_44696# a_15861_45028# 0.044605f
C37596 a_10227_46804# a_18479_45785# 6.39e-22
C37597 a_2609_46660# a_2711_45572# 7.29e-21
C37598 a_n743_46660# a_6428_45938# 1.23e-19
C37599 a_5807_45002# a_13527_45546# 2.96e-20
C37600 a_11415_45002# a_13759_46122# 7.28e-21
C37601 a_20411_46873# a_6945_45028# 1.76e-19
C37602 a_20273_46660# a_21137_46414# 0.007288f
C37603 a_20841_46902# a_20708_46348# 3.45e-19
C37604 a_12251_46660# a_12638_46436# 2.72e-19
C37605 a_19551_46910# a_10809_44734# 0.006863f
C37606 a_17639_46660# a_17715_44484# 3.97e-19
C37607 a_6151_47436# a_2437_43646# 0.017593f
C37608 a_2063_45854# a_n1059_45260# 1.14e-20
C37609 a_584_46384# a_n913_45002# 7.62e-20
C37610 a_n1151_42308# a_n2661_45010# 0.155007f
C37611 a_n746_45260# a_n143_45144# 0.043399f
C37612 a_2804_46116# a_3483_46348# 4.05e-19
C37613 a_2698_46116# a_3699_46348# 6.47e-20
C37614 a_15227_44166# a_8049_45260# 0.036339f
C37615 a_n2497_47436# a_3537_45260# 7.77e-19
C37616 a_1823_45246# a_5068_46348# 9.64e-20
C37617 a_n2661_46634# a_10053_45546# 2.08e-20
C37618 a_5534_30871# a_15051_42282# 2e-19
C37619 a_10867_43940# VDD 0.008055f
C37620 a_10903_43370# a_11551_42558# 9.18e-20
C37621 a_18114_32519# a_22223_43948# 0.003272f
C37622 a_11827_44484# a_14761_44260# 1.07e-19
C37623 a_n2840_46634# VDD 0.306342f
C37624 a_9838_44484# a_9672_43914# 7.43e-19
C37625 a_5883_43914# a_10405_44172# 6.88e-21
C37626 a_n1655_44484# a_n4318_39768# 1.21e-19
C37627 a_3232_43370# a_8791_43396# 1.36e-20
C37628 a_22612_30879# RST_Z 0.058603f
C37629 a_20916_46384# SINGLE_ENDED 0.020511f
C37630 a_16131_47204# CLK 3.58e-19
C37631 a_10193_42453# a_13635_43156# 0.001112f
C37632 a_n357_42282# a_8495_42852# 0.002316f
C37633 a_9290_44172# a_13575_42558# 0.001995f
C37634 a_1307_43914# a_3080_42308# 0.01819f
C37635 a_17517_44484# a_20835_44721# 0.029603f
C37636 a_n443_42852# a_5837_43172# 2.77e-19
C37637 a_n913_45002# a_15095_43370# 0.00588f
C37638 a_n1059_45260# a_14955_43396# 4.49e-20
C37639 a_2324_44458# a_6511_45714# 0.001394f
C37640 a_5807_45002# a_16922_45042# 0.030945f
C37641 a_n237_47217# a_n2661_43922# 1.49e-20
C37642 a_584_46384# a_556_44484# 0.004299f
C37643 a_4791_45118# a_7640_43914# 0.027432f
C37644 a_19466_46812# a_2437_43646# 1.21e-19
C37645 a_19692_46634# a_21513_45002# 0.098725f
C37646 a_n2293_46634# a_n2661_43370# 2.59564f
C37647 a_8016_46348# a_10193_42453# 0.125497f
C37648 a_8199_44636# a_10053_45546# 0.014322f
C37649 a_3483_46348# a_13904_45546# 0.125708f
C37650 a_12549_44172# a_21005_45260# 0.002789f
C37651 a_12861_44030# a_18443_44721# 0.007707f
C37652 a_17639_46660# a_15861_45028# 4.98e-21
C37653 a_11599_46634# a_17767_44458# 0.001378f
C37654 a_n1925_42282# a_n755_45592# 0.020368f
C37655 a_10227_46804# a_10057_43914# 0.054198f
C37656 a_17339_46660# a_18479_45785# 0.027772f
C37657 a_8953_45546# a_7499_43078# 0.108436f
C37658 a_5937_45572# a_9049_44484# 0.311862f
C37659 a_7577_46660# a_7705_45326# 3.37e-20
C37660 a_4646_46812# a_1307_43914# 0.031289f
C37661 a_5342_30871# C7_N_btm 5.39e-19
C37662 a_5932_42308# a_1343_38525# 2.86e-19
C37663 a_n3674_37592# a_n4209_38216# 1.31e-19
C37664 a_5534_30871# C9_N_btm 7.29e-20
C37665 a_13635_43156# VDD 0.463701f
C37666 a_5891_43370# a_9885_43396# 7.85e-20
C37667 a_3483_46348# CLK 0.408122f
C37668 a_n2661_42834# a_9145_43396# 1.09e-19
C37669 a_10193_42453# a_18310_42308# 0.004586f
C37670 a_n2017_45002# a_20256_42852# 4.86e-19
C37671 a_n2129_44697# a_n1853_43023# 6.76e-22
C37672 a_19478_44306# a_19862_44208# 0.001187f
C37673 a_18989_43940# a_15743_43084# 3.46e-19
C37674 a_n356_44636# a_16759_43396# 3.62e-21
C37675 a_n1549_44318# a_n4318_39304# 1.68e-19
C37676 a_n1331_43914# a_n2433_43396# 0.003897f
C37677 a_n1899_43946# a_n2129_43609# 4.63e-20
C37678 a_n1761_44111# a_n2267_43396# 1.9e-19
C37679 a_n2065_43946# a_n1699_43638# 1.48e-19
C37680 a_8016_46348# VDD 1.42798f
C37681 a_10729_43914# a_11816_44260# 0.003322f
C37682 a_10949_43914# a_11173_44260# 6.19e-19
C37683 a_10807_43548# a_10555_44260# 9.97e-20
C37684 a_17973_43940# a_11341_43940# 0.005348f
C37685 a_15682_43940# a_15493_43940# 0.067033f
C37686 a_13904_45546# a_14495_45572# 0.092344f
C37687 a_10193_42453# a_11682_45822# 0.032292f
C37688 a_10490_45724# a_10907_45822# 0.229517f
C37689 a_n2438_43548# a_453_43940# 0.001215f
C37690 a_768_44030# a_3820_44260# 3.84e-19
C37691 a_13259_45724# a_n2017_45002# 0.065062f
C37692 a_20850_46482# a_3357_43084# 7.81e-19
C37693 a_7499_43078# a_8791_45572# 0.004777f
C37694 a_8568_45546# a_9159_45572# 0.011449f
C37695 a_2711_45572# a_12561_45572# 4.68e-19
C37696 a_8270_45546# a_n2661_43922# 0.025118f
C37697 a_20205_31679# a_2437_43646# 3.32e-19
C37698 a_10227_46804# a_14021_43940# 0.062062f
C37699 a_n746_45260# a_n97_42460# 2.64e-19
C37700 a_n2497_47436# a_1049_43396# 3.45e-20
C37701 a_n971_45724# a_104_43370# 0.156156f
C37702 a_12741_44636# a_20205_45028# 0.001258f
C37703 a_20820_30879# a_18114_32519# 0.053f
C37704 a_n2293_46634# a_2998_44172# 0.06774f
C37705 a_13059_46348# a_14539_43914# 0.05997f
C37706 a_7174_31319# C5_N_btm 3.27e-20
C37707 a_n4064_40160# C5_P_btm 1.78e-19
C37708 a_n3420_38528# VDAC_P 2.69e-19
C37709 a_n4209_39590# C9_P_btm 0.786375f
C37710 a_n2946_37984# a_n3420_37440# 2.59e-20
C37711 a_n4064_37984# a_n3690_37440# 6.81e-20
C37712 a_n3565_38216# a_n2302_37690# 0.002384f
C37713 a_n3420_37984# a_n2946_37690# 2.59e-20
C37714 a_n3690_38304# a_n4064_37440# 6.81e-20
C37715 a_6151_47436# a_n2661_46634# 0.140541f
C37716 a_4915_47217# a_n2293_46634# 5.93e-19
C37717 a_n1435_47204# a_5807_45002# 3.71e-20
C37718 a_n237_47217# a_1799_45572# 0.417887f
C37719 a_n746_45260# a_n2661_46098# 0.049386f
C37720 a_3815_47204# a_n743_46660# 3.77e-20
C37721 a_16327_47482# a_12549_44172# 0.123271f
C37722 a_2063_45854# a_948_46660# 4.3e-21
C37723 a_n1151_42308# a_171_46873# 6.23e-19
C37724 a_2124_47436# a_1983_46706# 5.47e-20
C37725 a_584_46384# a_2107_46812# 0.007756f
C37726 a_4700_47436# a_n1925_46634# 7e-21
C37727 a_n1741_47186# a_3524_46660# 1.63e-20
C37728 a_n971_45724# a_2443_46660# 0.004065f
C37729 a_10227_46804# a_9804_47204# 4.77e-19
C37730 a_15673_47210# a_15928_47570# 0.064178f
C37731 a_5883_43914# a_6171_42473# 6.43e-23
C37732 a_9313_44734# a_20753_42852# 4.13e-19
C37733 a_2982_43646# a_6293_42852# 5.06e-20
C37734 a_4223_44672# a_5934_30871# 1.39e-21
C37735 a_5343_44458# a_7227_42308# 2.39e-19
C37736 a_11682_45822# VDD 0.316586f
C37737 a_22223_43948# a_13887_32519# 4.31e-19
C37738 a_15493_43940# a_22223_43396# 2.09e-20
C37739 a_n2661_42282# a_3935_42891# 2.51e-22
C37740 a_n356_44636# a_1067_42314# 0.019369f
C37741 a_14021_43940# a_19177_43646# 8.27e-19
C37742 a_17339_46660# a_14021_43940# 0.037923f
C37743 a_3775_45552# a_n2661_44458# 6.23e-21
C37744 a_5937_45572# a_3905_42865# 6.25e-21
C37745 a_3357_43084# a_4574_45260# 2.55e-21
C37746 a_n2293_46634# a_15681_43442# 1.89e-19
C37747 a_8746_45002# a_11827_44484# 1.23e-19
C37748 a_12741_44636# a_15682_43940# 0.003137f
C37749 a_n745_45366# a_n967_45348# 0.010748f
C37750 a_n2810_45028# en_comp 4.45e-19
C37751 a_13661_43548# a_18783_43370# 0.057336f
C37752 a_n2312_40392# a_n1853_43023# 2.89e-21
C37753 a_n443_42852# a_10334_44484# 1.29e-20
C37754 a_n357_42282# a_18287_44626# 1.16e-21
C37755 a_15227_44166# a_15037_43940# 0.010516f
C37756 a_2711_45572# a_2779_44458# 2.23e-20
C37757 a_n1059_45260# a_n955_45028# 4.12e-19
C37758 a_n2661_45010# a_327_44734# 0.04375f
C37759 a_n2293_45010# a_n37_45144# 7.8e-21
C37760 a_n2017_45002# a_n467_45028# 8.92e-22
C37761 a_5257_43370# a_3539_42460# 5.78e-20
C37762 a_5807_45002# a_13885_46660# 0.014137f
C37763 a_12549_44172# a_16434_46987# 6.15e-19
C37764 a_8128_46384# a_765_45546# 0.03129f
C37765 a_11453_44696# a_22365_46825# 0.001094f
C37766 a_13507_46334# a_21297_46660# 5.92e-19
C37767 a_21496_47436# a_21076_30879# 1.39e-19
C37768 a_n1151_42308# a_10903_43370# 7.29e-19
C37769 a_n743_46660# a_14976_45028# 0.024461f
C37770 a_4915_47217# a_9625_46129# 5.76e-20
C37771 a_6151_47436# a_8199_44636# 0.0013f
C37772 a_6540_46812# a_7577_46660# 3.44e-19
C37773 a_21811_47423# a_12741_44636# 1.79e-20
C37774 a_6293_42852# a_5837_42852# 0.001685f
C37775 a_20974_43370# a_20753_42852# 2.74e-20
C37776 a_n2472_42826# a_n2157_42858# 0.080495f
C37777 a_10341_43396# a_19339_43156# 9.56e-19
C37778 a_n2840_42826# a_n1853_43023# 3.22e-19
C37779 a_22223_45036# VDD 0.300162f
C37780 a_16922_45042# a_18315_45260# 0.065907f
C37781 a_3537_45260# a_6109_44484# 1.75e-19
C37782 a_n467_45028# a_n89_44484# 0.003687f
C37783 a_n2017_45002# a_n2661_43922# 0.034672f
C37784 a_n1059_45260# a_n2661_42834# 0.029616f
C37785 a_n2109_45247# a_n2293_43922# 7.56e-20
C37786 a_10227_46804# a_15764_42576# 0.024352f
C37787 a_20820_30879# a_13887_32519# 0.053104f
C37788 a_3090_45724# a_18083_42858# 9.89e-21
C37789 a_4791_45118# a_7174_31319# 9.47e-21
C37790 a_1307_43914# a_10057_43914# 0.03199f
C37791 a_9482_43914# a_16979_44734# 5.28e-20
C37792 a_13556_45296# a_14539_43914# 0.025347f
C37793 a_526_44458# a_648_43396# 0.04105f
C37794 a_7499_43078# a_9028_43914# 5.08e-20
C37795 a_18479_45785# a_18579_44172# 0.045071f
C37796 a_4185_45028# a_18783_43370# 1.92e-21
C37797 a_15227_44166# a_15279_43071# 0.002075f
C37798 a_n2312_38680# a_n1736_42282# 2.73e-20
C37799 a_n2442_46660# a_n1329_42308# 3.57e-20
C37800 a_1423_45028# a_8701_44490# 0.063232f
C37801 a_5093_45028# a_n2661_44458# 0.002375f
C37802 a_21076_30879# a_13678_32519# 0.05537f
C37803 a_14084_46812# a_10903_43370# 1.67e-21
C37804 a_14035_46660# a_3483_46348# 0.007996f
C37805 a_11599_46634# a_12791_45546# 5.33e-20
C37806 a_n743_46660# a_18051_46116# 1.36e-19
C37807 a_22000_46634# a_12741_44636# 0.044691f
C37808 a_21188_46660# a_22959_46660# 8.11e-21
C37809 a_5732_46660# a_5066_45546# 3.6e-22
C37810 a_768_44030# a_3503_45724# 1.76e-21
C37811 a_12991_46634# a_13351_46090# 0.011685f
C37812 a_12816_46660# a_12594_46348# 1.63e-20
C37813 a_12861_44030# a_13249_42308# 4.25e-19
C37814 a_13487_47204# a_13904_45546# 3e-19
C37815 a_4646_46812# a_8034_45724# 0.014576f
C37816 a_5257_43370# a_526_44458# 0.003403f
C37817 a_10227_46804# a_10180_45724# 0.03118f
C37818 a_17499_43370# a_18057_42282# 4.45e-19
C37819 a_743_42282# a_13657_42558# 0.007754f
C37820 a_21356_42826# a_22400_42852# 3.91e-20
C37821 a_4190_30871# a_15051_42282# 5.46e-20
C37822 a_13635_43156# a_n784_42308# 1.68e-20
C37823 a_5342_30871# COMP_P 0.027184f
C37824 a_17324_43396# a_17531_42308# 2.3e-21
C37825 a_5111_42852# a_5267_42460# 6.12e-19
C37826 a_4361_42308# a_13070_42354# 0.007985f
C37827 a_5649_42852# a_11551_42558# 6.94e-20
C37828 a_n2433_44484# a_n1331_43914# 0.001693f
C37829 a_n2661_44458# a_n1549_44318# 1.29e-20
C37830 a_17591_47464# VDD 0.421992f
C37831 a_13259_45724# a_19164_43230# 4.12e-20
C37832 a_n2293_46098# a_5932_42308# 1.61e-20
C37833 a_8696_44636# a_9803_43646# 5.08e-21
C37834 a_16588_47582# RST_Z 5.09e-20
C37835 a_n967_45348# a_n2433_43396# 0.00115f
C37836 en_comp a_n2129_43609# 0.008951f
C37837 a_n89_44484# a_n2661_43922# 3.35e-19
C37838 a_484_44484# a_n2661_42834# 4.92e-19
C37839 a_n1699_44726# a_n2065_43946# 7.01e-20
C37840 a_n2267_44484# a_n1761_44111# 1.89e-19
C37841 a_n2129_44697# a_n1899_43946# 2.08e-20
C37842 a_n443_42852# a_791_42968# 0.04806f
C37843 a_13487_47204# CLK 7.51e-19
C37844 a_1823_45246# a_2903_42308# 0.002746f
C37845 a_413_45260# a_14401_32519# 5.55e-20
C37846 a_1307_43914# a_14021_43940# 0.017312f
C37847 a_n755_45592# a_8387_43230# 0.010497f
C37848 a_n357_42282# a_9127_43156# 0.021342f
C37849 a_n2661_43370# a_9672_43914# 1.19e-37
C37850 a_n2661_45010# a_n1809_43762# 9.47e-20
C37851 a_n1059_45260# a_n1352_43396# 3.37e-20
C37852 a_n2293_45010# a_104_43370# 2.23e-19
C37853 a_n913_45002# a_n1177_43370# 0.014185f
C37854 a_18248_44752# a_19006_44850# 0.056391f
C37855 a_18287_44626# a_18588_44850# 9.73e-19
C37856 a_17970_44736# a_11967_42832# 0.00733f
C37857 a_584_46384# a_n2661_44458# 0.031143f
C37858 a_n2293_46634# a_4574_45260# 1.72e-21
C37859 a_15227_46910# a_11823_42460# 9.32e-22
C37860 a_10227_46804# a_13711_45394# 2.22e-20
C37861 a_13759_46122# a_13259_45724# 7.02e-19
C37862 a_13925_46122# a_14383_46116# 0.027606f
C37863 a_768_44030# a_14180_45002# 0.003277f
C37864 a_12549_44172# a_14537_43396# 0.037266f
C37865 a_2698_46116# a_n755_45592# 1.12e-19
C37866 a_n2293_46098# a_2307_45899# 3.74e-19
C37867 a_n746_45260# a_742_44458# 0.0971f
C37868 a_765_45546# a_10053_45546# 1.49e-20
C37869 a_167_45260# a_1848_45724# 0.359783f
C37870 a_n2438_43548# a_2274_45254# 1.51e-21
C37871 a_33_46660# a_413_45260# 4.39e-19
C37872 a_n1613_43370# a_1423_45028# 0.023846f
C37873 a_22959_46124# a_8049_45260# 0.003236f
C37874 a_1823_45246# a_3218_45724# 0.002867f
C37875 a_n1925_46634# a_3065_45002# 1.56e-20
C37876 a_4190_30871# C9_N_btm 0.002182f
C37877 a_8325_42308# a_9885_42558# 1.55e-21
C37878 a_8685_42308# a_9377_42558# 0.003285f
C37879 a_9223_42460# a_9803_42558# 0.001368f
C37880 a_13467_32519# C3_N_btm 1.74e-19
C37881 a_5534_30871# a_n3420_37440# 0.04166f
C37882 a_5934_30871# a_5742_30871# 16.7261f
C37883 a_n2661_42834# a_n2840_43370# 0.026572f
C37884 a_8975_43940# a_8791_43396# 4e-20
C37885 a_10057_43914# a_9396_43370# 1.26e-19
C37886 a_11827_44484# a_16243_43396# 1.51e-20
C37887 a_1307_43914# a_2075_43172# 0.077359f
C37888 a_13259_45724# a_21973_42336# 5.32e-20
C37889 a_22485_44484# a_22223_43948# 0.016889f
C37890 a_20512_43084# a_15493_43940# 0.021257f
C37891 a_6453_43914# a_n2661_42282# 0.122766f
C37892 a_14513_46634# CLK 2.54e-20
C37893 en_comp a_21195_42852# 4.83e-21
C37894 a_n357_42282# a_17124_42282# 0.011823f
C37895 a_n2956_38680# a_n3420_37984# 8.07e-19
C37896 a_18579_44172# a_14021_43940# 0.033047f
C37897 a_n443_42852# a_15051_42282# 9.06e-21
C37898 a_n1059_45260# a_n2293_42282# 0.033257f
C37899 a_12549_44172# a_20835_44721# 0.002438f
C37900 a_17715_44484# a_n1059_45260# 2.97e-20
C37901 a_19466_46812# a_19113_45348# 6.36e-19
C37902 a_13661_43548# a_16335_44484# 0.002382f
C37903 a_5937_45572# a_5147_45002# 8.8e-19
C37904 a_8199_44636# a_5111_44636# 0.024227f
C37905 a_13059_46348# a_14309_45028# 0.050896f
C37906 a_10809_44734# a_3357_43084# 0.035293f
C37907 a_15227_44166# a_20193_45348# 1.63e-20
C37908 a_n743_46660# a_15433_44458# 1.16e-21
C37909 a_3483_46348# a_10951_45334# 0.027449f
C37910 a_12005_46116# a_413_45260# 5.61e-21
C37911 a_6419_46155# a_6171_45002# 1.62e-19
C37912 a_13259_45724# a_15297_45822# 1.06e-19
C37913 a_6472_45840# a_6598_45938# 0.178024f
C37914 a_6511_45714# a_6667_45809# 0.113977f
C37915 a_n2293_46098# a_1423_45028# 0.017396f
C37916 a_5497_46414# a_5205_44484# 6.8e-22
C37917 a_5932_42308# C5_N_btm 5.59e-19
C37918 a_5742_30871# a_11530_34132# 7.08e-19
C37919 a_13717_47436# a_13487_47204# 0.061247f
C37920 a_n3565_38502# a_n3690_38528# 0.246863f
C37921 a_1736_39043# a_1177_38525# 1.72e-19
C37922 a_n4334_38528# a_n3420_38528# 0.015595f
C37923 a_n4209_38502# a_n2946_38778# 0.022704f
C37924 a_n4064_39072# a_n4334_38304# 3.17e-19
C37925 a_5934_30871# C0_dummy_P_btm 1.48e-19
C37926 a_11459_47204# a_11599_46634# 0.019787f
C37927 a_n2497_47436# a_n1613_43370# 0.402561f
C37928 a_n2109_47186# a_3094_47243# 0.003449f
C37929 a_n1741_47186# a_4842_47570# 2.25e-19
C37930 a_n237_47217# a_2747_46873# 5.93e-20
C37931 a_n971_45724# a_7_47243# 0.005756f
C37932 a_3905_42558# VDD 0.176395f
C37933 a_6123_31319# C0_N_btm 0.018968f
C37934 a_n4209_39304# a_n2302_37984# 1.04e-19
C37935 a_17124_42282# CAL_N 0.001755f
C37936 a_n1151_42308# a_4883_46098# 0.407909f
C37937 en_comp a_n2302_40160# 2.07e-19
C37938 a_n1013_45572# VDD 4.04e-19
C37939 a_17973_43940# a_10341_43396# 1.83e-20
C37940 a_n2065_43946# a_n2157_42858# 6.86e-21
C37941 a_1307_43914# a_15764_42576# 8.77e-22
C37942 a_n2433_43396# a_n1917_43396# 0.108815f
C37943 a_n2129_43609# a_n1699_43638# 0.022218f
C37944 a_2998_44172# a_743_42282# 1.28e-20
C37945 a_768_44030# a_6765_43638# 1.04e-20
C37946 a_8696_44636# a_n913_45002# 2.6e-20
C37947 a_n971_45724# a_n1076_43230# 0.003103f
C37948 a_13527_45546# a_13017_45260# 9.04e-20
C37949 a_13163_45724# a_13159_45002# 0.010135f
C37950 a_2277_45546# a_n2661_43370# 5.63e-21
C37951 a_10193_42453# a_16019_45002# 6.67e-19
C37952 a_10907_45822# a_6171_45002# 0.024408f
C37953 a_16327_47482# a_16977_43638# 0.15941f
C37954 a_n2497_47436# a_n1533_42852# 2.22e-19
C37955 a_12861_44030# a_19700_43370# 1.67e-20
C37956 a_11823_42460# a_9482_43914# 0.033152f
C37957 a_10227_46804# a_13943_43396# 2.15e-20
C37958 a_3090_45724# a_12429_44172# 1.23e-21
C37959 a_n443_42852# a_13105_45348# 1.05e-20
C37960 a_2711_45572# a_7639_45394# 2.87e-19
C37961 a_n2293_46634# a_1568_43370# 2.04e-19
C37962 a_13661_43548# a_3626_43646# 2.98e-20
C37963 C10_P_btm C5_P_btm 0.285351f
C37964 a_4883_46098# a_14084_46812# 4.58e-20
C37965 a_1123_46634# a_1799_45572# 0.037438f
C37966 a_383_46660# a_n2661_46098# 0.002826f
C37967 a_9804_47204# a_10467_46802# 3.93e-21
C37968 a_n881_46662# a_6969_46634# 1.79e-19
C37969 a_13717_47436# a_14513_46634# 1.71e-20
C37970 a_12861_44030# a_14180_46812# 0.238709f
C37971 a_13487_47204# a_14035_46660# 0.002982f
C37972 a_11453_44696# a_11901_46660# 2.64e-21
C37973 VDAC_N VREF_GND 0.327524f
C37974 a_13507_46334# a_3090_45724# 0.020036f
C37975 a_18597_46090# a_18834_46812# 0.010699f
C37976 C9_P_btm C6_P_btm 0.169882f
C37977 C8_P_btm C7_P_btm 23.7884f
C37978 a_6151_47436# a_765_45546# 0.191559f
C37979 a_n1613_43370# a_6682_46987# 1.74e-19
C37980 a_n2497_47436# a_n2293_46098# 0.039224f
C37981 a_22876_39857# VDD 3.12e-19
C37982 a_14311_47204# a_13885_46660# 2.65e-19
C37983 a_18780_47178# a_15227_44166# 2.49e-19
C37984 a_18479_47436# a_19333_46634# 5.75e-19
C37985 a_10227_46804# a_19692_46634# 0.239326f
C37986 a_12465_44636# a_12816_46660# 4.51e-21
C37987 a_16547_43609# a_16823_43084# 0.08061f
C37988 a_15743_43084# a_16867_43762# 8.49e-19
C37989 a_16977_43638# a_16855_43396# 3.16e-19
C37990 a_16243_43396# a_17433_43396# 2.56e-19
C37991 a_2982_43646# a_10991_42826# 1.03e-19
C37992 a_3626_43646# a_10835_43094# 2.04e-20
C37993 a_11967_42832# a_16104_42674# 4.18e-19
C37994 a_16019_45002# VDD 0.174085f
C37995 a_5244_44056# a_4921_42308# 1.76e-21
C37996 a_n2661_42282# a_n3674_37592# 0.12829f
C37997 a_n97_42460# a_19339_43156# 0.012502f
C37998 a_10341_43396# a_22591_43396# 0.172197f
C37999 a_6197_43396# a_7227_42852# 3.42e-20
C38000 a_3357_43084# a_5883_43914# 0.046158f
C38001 a_13259_45724# a_18079_43940# 0.007888f
C38002 a_19692_46634# a_19177_43646# 8.77e-21
C38003 a_4791_45118# a_5932_42308# 0.212275f
C38004 a_n443_42852# a_3905_42865# 0.043488f
C38005 a_n863_45724# a_1525_44260# 2.55e-19
C38006 a_n1059_45260# a_n1352_44484# 2.66e-19
C38007 a_n913_45002# a_n1177_44458# 0.017911f
C38008 a_16375_45002# a_15682_43940# 5.84e-19
C38009 a_n2293_45010# a_949_44458# 0.001253f
C38010 a_626_44172# a_n2661_43370# 0.008858f
C38011 a_14797_45144# a_15060_45348# 0.010598f
C38012 a_3232_43370# a_11827_44484# 0.094278f
C38013 a_n967_45348# a_n2433_44484# 3.53e-20
C38014 a_4185_45028# a_3626_43646# 0.035503f
C38015 en_comp a_n2129_44697# 0.00879f
C38016 a_10193_42453# a_18245_44484# 1.51e-19
C38017 a_10227_46804# a_20692_30879# 1.56e-20
C38018 a_n2293_46634# a_10809_44734# 7.76e-20
C38019 a_5385_46902# a_5497_46414# 5.03e-20
C38020 a_5167_46660# a_5204_45822# 0.002145f
C38021 a_2905_45572# a_2711_45572# 0.041827f
C38022 a_n443_46116# a_1990_45899# 0.002313f
C38023 a_18834_46812# a_19123_46287# 0.039405f
C38024 a_15227_44166# a_18285_46348# 0.097182f
C38025 a_13885_46660# a_14226_46987# 0.003464f
C38026 a_19692_46634# a_17339_46660# 8.51e-21
C38027 a_9804_47204# a_8034_45724# 1.12e-19
C38028 a_4646_46812# a_8016_46348# 4.3e-21
C38029 a_2063_45854# a_5263_45724# 0.030969f
C38030 a_n2472_46634# a_n2956_39304# 8.55e-19
C38031 a_4883_46098# a_19240_46482# 0.002371f
C38032 a_3422_30871# C4_N_btm 1.36e-19
C38033 a_21195_42852# a_22165_42308# 0.007883f
C38034 a_2982_43646# a_17303_42282# 0.139588f
C38035 a_3626_43646# a_16269_42308# 0.001405f
C38036 a_8605_42826# a_9114_42852# 2.6e-19
C38037 a_n4318_39304# a_n4334_39616# 7.95e-19
C38038 a_17364_32525# a_14097_32519# 0.059348f
C38039 a_5111_44636# a_8018_44260# 4.54e-19
C38040 a_n357_42282# a_19268_43646# 1.71e-20
C38041 a_3090_45724# a_7227_42308# 4.26e-20
C38042 a_8103_44636# a_7640_43914# 0.101633f
C38043 a_5518_44484# a_5891_43370# 2.14e-20
C38044 a_5343_44458# a_8238_44734# 1.98e-21
C38045 a_n2661_44458# a_11649_44734# 8.36e-19
C38046 a_3232_43370# a_6756_44260# 6.17e-21
C38047 a_n2956_39768# a_n3420_39072# 8.07e-19
C38048 a_18287_44626# a_18443_44721# 0.10279f
C38049 a_18248_44752# a_18374_44850# 0.170059f
C38050 a_17970_44736# a_18989_43940# 1.91e-21
C38051 a_1423_45028# a_2675_43914# 4.85e-20
C38052 a_1307_43914# a_5013_44260# 0.358053f
C38053 a_6298_44484# a_8375_44464# 8.94e-21
C38054 a_20567_45036# a_17517_44484# 7.16e-20
C38055 a_n2840_44458# a_n2661_43922# 0.001534f
C38056 a_11827_44484# a_14581_44484# 1.34e-19
C38057 a_526_44458# a_10518_42984# 1.06e-19
C38058 a_n2312_40392# en_comp 0.036842f
C38059 a_n2312_39304# a_n2956_37592# 0.047801f
C38060 a_15015_46420# a_2324_44458# 0.027704f
C38061 a_3699_46348# a_526_44458# 0.00137f
C38062 a_3483_46348# a_n1925_42282# 0.536704f
C38063 a_10428_46928# a_10193_42453# 3.41e-20
C38064 a_10150_46912# a_8746_45002# 1.91e-19
C38065 a_9823_46155# a_6945_45028# 1.27e-20
C38066 a_12816_46660# a_2711_45572# 2.6e-20
C38067 a_n881_46662# a_3357_43084# 0.028875f
C38068 a_4791_45118# a_1423_45028# 0.721318f
C38069 a_2107_46812# a_8696_44636# 0.025973f
C38070 a_21811_47423# a_413_45260# 8.86e-20
C38071 a_14635_42282# a_15051_42282# 0.007421f
C38072 a_8791_43396# VDD 0.191045f
C38073 a_4190_30871# a_n3420_37440# 0.034998f
C38074 a_1755_42282# a_2351_42308# 3.31e-19
C38075 a_n2293_42282# a_n4315_30879# 3.44e-21
C38076 a_n2065_43946# a_n1761_44111# 0.617556f
C38077 a_2382_45260# a_4361_42308# 3.26e-20
C38078 en_comp a_n2840_42826# 0.002468f
C38079 a_n2293_45010# a_n1076_43230# 3.21e-21
C38080 a_n2017_45002# a_n1641_43230# 0.011397f
C38081 a_n913_45002# a_n1991_42858# 0.024791f
C38082 a_n1059_45260# a_n1423_42826# 2.7e-19
C38083 a_n2267_44484# a_n2267_43396# 0.001024f
C38084 a_n1917_44484# a_n2433_43396# 2.16e-20
C38085 a_n357_42282# a_1755_42282# 2.68e-19
C38086 a_n755_45592# a_1606_42308# 0.104938f
C38087 a_n863_45724# a_2725_42558# 0.003172f
C38088 a_10428_46928# VDD 0.278873f
C38089 a_7715_46873# DATA[3] 7.9e-19
C38090 a_n2433_44484# a_n1917_43396# 2.93e-20
C38091 a_9313_44734# a_11341_43940# 1.41e-19
C38092 a_380_45546# a_n755_45592# 4.05e-19
C38093 a_n1099_45572# a_n357_42282# 0.013419f
C38094 a_n2661_45546# a_n356_45724# 0.008001f
C38095 a_13661_43548# a_17767_44458# 5.86e-21
C38096 a_22000_46634# a_413_45260# 4.39e-20
C38097 a_20202_43084# a_n2017_45002# 0.005245f
C38098 a_11453_44696# a_11649_44734# 3.12e-19
C38099 a_15682_46116# a_15765_45572# 0.015911f
C38100 a_17715_44484# a_15599_45572# 1.85e-19
C38101 a_n2497_47436# a_2675_43914# 6.16e-20
C38102 a_12465_44636# a_13213_44734# 1.97e-20
C38103 a_n1613_43370# a_6109_44484# 0.099934f
C38104 a_n746_45260# a_n984_44318# 4.22e-20
C38105 a_10903_43370# a_12649_45572# 0.006357f
C38106 a_8049_45260# a_8568_45546# 0.003997f
C38107 a_n2293_46634# a_5883_43914# 0.00136f
C38108 a_n743_46660# a_5343_44458# 5.3e-23
C38109 a_n863_45724# a_1848_45724# 5.68e-20
C38110 a_n4064_40160# a_n4209_39590# 0.059936f
C38111 a_n2302_40160# a_n2216_40160# 0.011479f
C38112 a_n4315_30879# a_n3565_39590# 0.027163f
C38113 a_5742_30871# a_7754_40130# 0.005581f
C38114 a_n4334_40480# a_n4334_39616# 0.050585f
C38115 a_n2109_47186# a_4007_47204# 0.047269f
C38116 a_n1741_47186# a_3785_47178# 0.047034f
C38117 a_n237_47217# a_2063_45854# 0.947844f
C38118 a_327_47204# a_1431_47204# 1.62e-20
C38119 a_n1605_47204# a_n1151_42308# 0.001389f
C38120 a_n971_45724# a_2952_47436# 0.019506f
C38121 a_1209_47178# a_1239_47204# 0.264529f
C38122 a_2998_44172# a_2813_43396# 2e-19
C38123 a_11967_42832# a_18783_43370# 0.001091f
C38124 a_375_42282# a_n961_42308# 3.02e-20
C38125 a_11341_43940# a_20974_43370# 0.013722f
C38126 a_22223_43948# a_14401_32519# 0.157135f
C38127 a_15493_43940# a_21381_43940# 0.02116f
C38128 a_5111_44636# a_4921_42308# 0.004461f
C38129 a_3537_45260# a_6171_42473# 3.79e-20
C38130 a_22591_44484# a_10341_43396# 3.21e-19
C38131 a_n913_45002# a_9377_42558# 2.17e-19
C38132 a_n2017_45002# a_10545_42558# 9.16e-19
C38133 a_17973_43940# a_n97_42460# 1.1e-21
C38134 a_7281_43914# a_7287_43370# 0.003639f
C38135 a_3232_43370# a_3581_42558# 7.4e-20
C38136 a_n356_44636# a_5111_42852# 1.83e-20
C38137 a_20205_31679# a_22609_38406# 4.1e-21
C38138 a_8049_45260# a_n2661_43370# 0.013528f
C38139 a_3483_46348# a_18248_44752# 2.73e-21
C38140 a_n2293_46098# a_6109_44484# 2.32e-19
C38141 a_n443_46116# a_3457_43396# 3.38e-20
C38142 a_8953_45546# a_9838_44484# 9.26e-20
C38143 a_8199_44636# a_10334_44484# 6.58e-19
C38144 a_8016_46348# a_10057_43914# 0.09388f
C38145 a_n443_42852# a_5147_45002# 0.004185f
C38146 a_15599_45572# a_15861_45028# 1.72e-20
C38147 a_15903_45785# a_8696_44636# 1.89e-19
C38148 a_15765_45572# a_16680_45572# 0.118759f
C38149 a_4646_46812# a_7584_44260# 5.27e-19
C38150 a_19692_46634# a_18579_44172# 3.19e-19
C38151 a_n4209_38502# VREF 0.059621f
C38152 VDAC_P CAL_N 2.76e-19
C38153 a_n4334_38304# VDD 0.385989f
C38154 a_3754_38470# a_n923_35174# 0.002509f
C38155 a_n3565_38502# VIN_P 0.029053f
C38156 a_2063_45854# a_8270_45546# 0.017994f
C38157 a_6575_47204# a_8667_46634# 0.01088f
C38158 a_4915_47217# a_6755_46942# 0.260675f
C38159 a_6151_47436# a_10623_46897# 4.99e-20
C38160 a_2747_46873# a_1123_46634# 2.46e-20
C38161 a_2266_47570# a_2107_46812# 2.38e-19
C38162 a_n881_46662# a_n2293_46634# 0.026189f
C38163 a_14021_43940# a_13635_43156# 0.001414f
C38164 a_n2129_43609# a_n2157_42858# 0.007212f
C38165 a_n2433_43396# a_n1853_43023# 4.61e-19
C38166 a_1568_43370# a_743_42282# 2.22e-19
C38167 a_9145_43396# a_15095_43370# 0.213415f
C38168 a_19963_31679# C4_N_btm 0.001041f
C38169 a_20623_43914# a_19987_42826# 1.37e-19
C38170 a_15493_43940# a_18249_42858# 2.89e-20
C38171 a_11341_43940# a_18599_43230# 3.88e-20
C38172 a_19237_31679# a_14097_32519# 0.052198f
C38173 a_19479_31679# C7_N_btm 1.43e-20
C38174 a_9313_44734# a_10723_42308# 1.32e-20
C38175 a_13667_43396# a_14579_43548# 5.78e-19
C38176 a_19862_44208# a_21195_42852# 0.002065f
C38177 a_4099_45572# a_n2661_43922# 2.36e-20
C38178 a_4927_45028# a_1307_43914# 8.94e-21
C38179 a_8696_44636# a_n2661_44458# 1.37553f
C38180 a_12549_44172# a_12379_42858# 3.65e-20
C38181 w_11334_34010# COMP_P 0.004781f
C38182 SMPL_ON_P a_n3674_38680# 0.038963f
C38183 a_6171_45002# a_15415_45028# 0.008633f
C38184 a_n2661_45010# a_n2293_42834# 2.08e-20
C38185 a_20107_45572# a_16922_45042# 1.06e-19
C38186 a_n2438_43548# a_n1736_43218# 2.63e-20
C38187 a_18341_45572# a_11827_44484# 6.05e-21
C38188 a_17715_44484# a_18326_43940# 0.003424f
C38189 a_2324_44458# a_15493_43396# 4.05e-19
C38190 a_18189_46348# a_18079_43940# 1.25e-19
C38191 a_2274_45254# a_2903_45348# 6.01e-19
C38192 a_2680_45002# a_2304_45348# 1.96e-19
C38193 a_20820_30879# a_14401_32519# 0.055735f
C38194 a_9290_44172# a_9895_44260# 3.38e-19
C38195 a_n2497_47436# a_n1736_42282# 3.98e-19
C38196 a_n1151_42308# a_11608_46482# 7.22e-19
C38197 a_n2293_46634# a_n2157_46122# 0.04308f
C38198 a_n2104_46634# a_n2293_46098# 0.002261f
C38199 a_11453_44696# a_17583_46090# 1.99e-20
C38200 a_13507_46334# a_20075_46420# 0.006404f
C38201 a_20990_47178# a_20708_46348# 2.85e-21
C38202 a_19787_47423# a_6945_45028# 0.009959f
C38203 a_768_44030# a_5164_46348# 4.84e-20
C38204 a_10150_46912# a_10425_46660# 0.007416f
C38205 a_9804_47204# a_8016_46348# 0.009763f
C38206 a_8128_46384# a_8349_46414# 0.101217f
C38207 a_n881_46662# a_9625_46129# 3.67e-20
C38208 a_12465_44636# a_18819_46122# 2.8e-20
C38209 a_18597_46090# a_10809_44734# 0.036294f
C38210 a_4883_46098# a_19553_46090# 0.005361f
C38211 a_4915_47217# a_8049_45260# 0.022494f
C38212 a_n2312_38680# a_n2472_46090# 0.001445f
C38213 a_n1243_44484# VDD 7.26e-20
C38214 a_3422_30871# a_8530_39574# 1.13e-19
C38215 a_2982_43646# a_2713_42308# 1.35e-21
C38216 a_2896_43646# a_2903_42308# 7.11e-21
C38217 a_3080_42308# a_3905_42558# 0.008414f
C38218 a_4905_42826# a_3581_42558# 8.56e-21
C38219 a_17364_32525# a_22959_42860# 5e-19
C38220 a_9127_43156# a_8952_43230# 0.234322f
C38221 a_15227_44166# a_15785_43172# 9.28e-19
C38222 a_n863_45724# a_1512_43396# 1.35e-19
C38223 a_18315_45260# a_17970_44736# 6.02e-19
C38224 a_11691_44458# a_10157_44484# 1.48e-20
C38225 a_13556_45296# a_15146_44484# 4.94e-20
C38226 a_4185_45028# a_8037_42858# 2.64e-20
C38227 a_3483_46348# a_8387_43230# 7.21e-22
C38228 a_20202_43084# a_19164_43230# 1.12e-19
C38229 a_12549_44172# a_18727_42674# 1.47e-21
C38230 a_3090_45724# a_14853_42852# 4.1e-19
C38231 a_n755_45592# a_3539_42460# 0.008691f
C38232 a_n2433_44484# a_n1917_44484# 0.113784f
C38233 a_16922_45042# a_18374_44850# 9.15e-20
C38234 a_n2661_44458# a_n1177_44458# 0.006328f
C38235 a_11827_44484# a_8975_43940# 0.076327f
C38236 a_n2661_43370# a_5289_44734# 3.39e-19
C38237 en_comp a_n2472_43914# 0.014244f
C38238 a_n2312_40392# a_n2216_40160# 0.001083f
C38239 a_n913_45002# a_n1331_43914# 3.47e-19
C38240 a_n2293_45010# a_175_44278# 0.030523f
C38241 a_n2017_45002# a_n809_44244# 1.63e-21
C38242 a_n2661_45010# a_1115_44172# 0.003124f
C38243 a_n1059_45260# a_n1549_44318# 3.77e-19
C38244 a_n2129_44697# a_n1699_44726# 0.018607f
C38245 a_15415_45028# a_14673_44172# 9.28e-20
C38246 a_n443_42852# a_4093_43548# 0.028988f
C38247 a_15037_45618# a_11341_43940# 2.21e-21
C38248 a_16327_47482# a_19431_45546# 0.344862f
C38249 a_n2661_46634# a_9049_44484# 4.26e-20
C38250 a_1823_45246# a_4704_46090# 0.164557f
C38251 a_n443_46116# a_3357_43084# 0.006081f
C38252 a_11453_44696# a_8696_44636# 2.67247f
C38253 a_10227_46804# a_18175_45572# 1.6e-21
C38254 a_2443_46660# a_2711_45572# 5.4e-21
C38255 a_5807_45002# a_13163_45724# 7.62e-21
C38256 a_19123_46287# a_10809_44734# 0.009463f
C38257 a_20273_46660# a_20708_46348# 0.004461f
C38258 a_20107_46660# a_6945_45028# 0.024966f
C38259 a_12251_46660# a_12379_46436# 4.35e-19
C38260 a_20411_46873# a_21137_46414# 2.11e-20
C38261 a_17639_46660# a_17583_46090# 3.95e-19
C38262 a_5815_47464# a_2437_43646# 0.00818f
C38263 a_12861_44030# a_18787_45572# 1.98e-19
C38264 a_2063_45854# a_n2017_45002# 1.9e-20
C38265 a_584_46384# a_n1059_45260# 6.25e-20
C38266 a_n746_45260# a_n467_45028# 0.054826f
C38267 a_2804_46116# a_3147_46376# 0.017019f
C38268 a_2698_46116# a_3483_46348# 1.66e-19
C38269 a_3090_45724# a_10586_45546# 0.002067f
C38270 a_11415_45002# a_13351_46090# 4.86e-21
C38271 a_12741_44636# a_10903_43370# 4.89e-19
C38272 a_13747_46662# a_11823_42460# 0.521845f
C38273 a_2107_46812# a_7227_45028# 7.51e-20
C38274 a_20256_43172# a_20573_43172# 0.001295f
C38275 a_10341_42308# a_10149_42308# 1.97e-19
C38276 a_5534_30871# a_14113_42308# 5.72e-21
C38277 a_10651_43940# VDD 0.003431f
C38278 a_10903_43370# a_5742_30871# 5.9e-20
C38279 a_22612_30879# VDD 3.2377f
C38280 a_626_44172# a_1568_43370# 1.82e-21
C38281 a_5883_43914# a_9672_43914# 4.69e-19
C38282 a_n1821_44484# a_n4318_39768# 3.01e-19
C38283 a_3232_43370# a_8147_43396# 1.83e-19
C38284 a_3537_45260# a_3457_43396# 3.07e-20
C38285 a_21588_30879# RST_Z 0.052092f
C38286 a_11823_42460# a_10796_42968# 5.88e-19
C38287 a_10193_42453# a_12895_43230# 1.15e-20
C38288 a_n357_42282# a_9306_43218# 1.74e-19
C38289 a_9290_44172# a_13070_42354# 0.140007f
C38290 a_13259_45724# a_17749_42852# 0.001312f
C38291 a_21076_30879# a_22775_42308# 6.58e-21
C38292 a_1307_43914# a_4699_43561# 1.54e-19
C38293 a_17517_44484# a_20679_44626# 0.031895f
C38294 a_5205_44484# a_6547_43396# 1.82e-19
C38295 a_7229_43940# a_6197_43396# 0.001981f
C38296 a_n443_42852# a_5457_43172# 2.37e-19
C38297 a_n1925_42282# a_2351_42308# 5.44e-20
C38298 a_5807_45002# DATA[5] 3.78e-20
C38299 a_5111_44636# a_6452_43396# 0.024938f
C38300 a_n1059_45260# a_15095_43370# 0.108103f
C38301 a_n913_45002# a_14205_43396# 3.11e-19
C38302 a_2324_44458# a_6472_45840# 2.1e-19
C38303 a_n2661_46634# a_13105_45348# 0.009374f
C38304 a_7411_46660# a_8191_45002# 2.65e-23
C38305 a_n746_45260# a_n2661_43922# 0.037244f
C38306 a_n971_45724# a_n2293_43922# 2.81e-19
C38307 a_584_46384# a_484_44484# 0.001797f
C38308 a_4791_45118# a_6109_44484# 3.61e-20
C38309 a_n2442_46660# a_n2661_43370# 1.23e-19
C38310 a_3483_46348# a_13527_45546# 4.96e-19
C38311 a_8016_46348# a_10180_45724# 0.259851f
C38312 a_9863_46634# a_6171_45002# 1.59e-22
C38313 a_12549_44172# a_20567_45036# 0.176249f
C38314 a_12861_44030# a_18287_44626# 0.029719f
C38315 a_19333_46634# a_2437_43646# 3.78e-21
C38316 a_10227_46804# a_10440_44484# 0.025362f
C38317 a_17339_46660# a_18175_45572# 0.019286f
C38318 a_5937_45572# a_7499_43078# 0.033831f
C38319 a_8199_44636# a_9049_44484# 0.029722f
C38320 a_8953_45546# a_8568_45546# 0.136365f
C38321 a_7715_46873# a_7705_45326# 0.001207f
C38322 a_3877_44458# a_1307_43914# 4.73e-20
C38323 a_n1925_42282# a_n357_42282# 0.023161f
C38324 a_526_44458# a_n755_45592# 0.065199f
C38325 a_5342_30871# C6_N_btm 0.012f
C38326 a_14456_42282# a_7174_31319# 9.76e-21
C38327 a_5534_30871# C8_N_btm 5.29e-19
C38328 a_12895_43230# VDD 0.212352f
C38329 a_1606_42308# a_n3420_38528# 2.3e-20
C38330 a_9313_44734# a_10341_43396# 0.175125f
C38331 a_5891_43370# a_8945_43396# 2.41e-19
C38332 a_11823_42460# a_4958_30871# 4.65e-19
C38333 a_n2017_45002# a_19326_42852# 3.73e-19
C38334 a_n913_45002# a_22400_42852# 0.002067f
C38335 a_5343_44458# a_4361_42308# 0.004068f
C38336 a_n2433_44484# a_n1853_43023# 2.06e-21
C38337 a_10193_42453# a_18220_42308# 0.004148f
C38338 a_15493_43396# a_19862_44208# 8.78e-19
C38339 a_11967_42832# a_3626_43646# 0.001552f
C38340 a_n356_44636# a_16977_43638# 1.19e-21
C38341 a_5883_43914# a_743_42282# 3.05e-20
C38342 a_18989_43940# a_18783_43370# 4.79e-19
C38343 a_n1899_43946# a_n2433_43396# 6.91e-19
C38344 a_n1761_44111# a_n2129_43609# 0.029483f
C38345 a_n2065_43946# a_n2267_43396# 0.009359f
C38346 a_7920_46348# VDD 0.100184f
C38347 a_17737_43940# a_11341_43940# 0.004705f
C38348 a_14955_43940# a_15493_43940# 0.110232f
C38349 a_10949_43914# a_10555_44260# 0.034175f
C38350 a_10729_43914# a_11173_44260# 0.057346f
C38351 a_19479_31679# COMP_P 2e-20
C38352 a_6945_45028# a_1423_45028# 1.15e-19
C38353 a_13904_45546# a_13249_42308# 0.13587f
C38354 a_10490_45724# a_10210_45822# 0.014252f
C38355 a_8746_45002# a_10907_45822# 1.47e-19
C38356 a_8953_45546# a_n2661_43370# 0.02624f
C38357 a_3483_46348# a_16922_45042# 3.56e-19
C38358 a_768_44030# a_3499_42826# 0.034429f
C38359 a_11415_45002# a_19721_31679# 0.001159f
C38360 a_5066_45546# a_7229_43940# 4.19e-21
C38361 a_8568_45546# a_8791_45572# 0.011458f
C38362 a_7499_43078# a_8697_45572# 0.004673f
C38363 a_n2438_43548# a_1414_42308# 0.001019f
C38364 a_8270_45546# a_n2661_42834# 0.034362f
C38365 a_10227_46804# a_13829_44260# 1.01e-19
C38366 a_12465_44636# a_11341_43940# 0.002963f
C38367 a_12741_44636# a_19929_45028# 0.001258f
C38368 a_n2293_46634# a_2889_44172# 1.86e-19
C38369 a_n2497_47436# a_1209_43370# 1.74e-20
C38370 a_n971_45724# a_n97_42460# 0.581616f
C38371 a_n1741_47186# a_3699_46634# 1.51e-19
C38372 a_n443_46116# a_n2293_46634# 0.050675f
C38373 a_5815_47464# a_n2661_46634# 1.29e-19
C38374 a_13381_47204# a_5807_45002# 5.2e-20
C38375 a_7174_31319# C4_N_btm 2.64e-20
C38376 a_n4064_40160# C6_P_btm 2.2e-19
C38377 a_15507_47210# a_16119_47582# 3.82e-19
C38378 a_n971_45724# a_n2661_46098# 0.023255f
C38379 a_n746_45260# a_1799_45572# 4.63e-22
C38380 a_n1151_42308# a_n133_46660# 0.002432f
C38381 a_3785_47178# a_n743_46660# 2.74e-21
C38382 a_n4209_39590# C10_P_btm 0.002325f
C38383 a_13258_32519# C7_N_btm 1.33e-20
C38384 a_584_46384# a_948_46660# 0.002817f
C38385 a_2124_47436# a_2107_46812# 0.010665f
C38386 a_4007_47204# a_n1925_46634# 8.66e-20
C38387 a_15673_47210# a_768_44030# 2.86e-20
C38388 a_15811_47375# a_15928_47570# 0.161235f
C38389 a_n4064_37984# a_n3565_37414# 0.029309f
C38390 a_n3420_37984# a_n3420_37440# 0.132162f
C38391 a_n3565_38216# a_n4064_37440# 0.032797f
C38392 VDAC_Pi a_3754_38802# 0.00191f
C38393 a_5883_43914# a_5755_42308# 4.69e-21
C38394 a_2982_43646# a_6031_43396# 8.49e-21
C38395 a_1568_43370# a_2813_43396# 4.85e-19
C38396 a_20974_43370# a_10341_43396# 0.08579f
C38397 a_5343_44458# a_6761_42308# 1.34e-19
C38398 a_11280_45822# VDD 0.004437f
C38399 a_22223_43948# a_22223_43396# 0.025171f
C38400 a_n2661_42282# a_3681_42891# 1.24e-20
C38401 a_15493_43940# a_5649_42852# 3.25e-20
C38402 a_n356_44636# a_n1630_35242# 5.72e-21
C38403 a_4223_44672# a_7963_42308# 2.12e-21
C38404 a_3090_45724# a_19478_44056# 0.002976f
C38405 a_3357_43084# a_3537_45260# 0.026461f
C38406 a_n2293_46634# a_14621_43646# 0.002737f
C38407 a_10193_42453# a_11827_44484# 0.121679f
C38408 a_7499_43078# a_11691_44458# 0.007969f
C38409 a_n913_45002# a_n967_45348# 1.00127f
C38410 a_n2810_45028# a_n2956_37592# 6.13705f
C38411 a_13661_43548# a_18525_43370# 0.031188f
C38412 a_n2312_40392# a_n2157_42858# 5.78e-21
C38413 a_n1059_45260# a_n659_45366# 0.001645f
C38414 a_n2661_45010# a_413_45260# 0.003446f
C38415 a_n2293_45010# a_n143_45144# 7.12e-21
C38416 a_16147_45260# a_16751_45260# 0.054632f
C38417 a_n2661_45546# a_n356_44636# 3.08e-21
C38418 a_5257_43370# a_3626_43646# 5.37e-20
C38419 a_n357_42282# a_18248_44752# 9.12e-22
C38420 a_n443_42852# a_10157_44484# 1.48e-20
C38421 a_5732_46660# a_7577_46660# 3.52e-20
C38422 a_6540_46812# a_7715_46873# 1.3e-19
C38423 a_5807_45002# a_13170_46660# 3.81e-19
C38424 a_12549_44172# a_16721_46634# 0.013883f
C38425 a_n1435_47204# a_3483_46348# 1.31e-20
C38426 a_5159_47243# a_765_45546# 2e-19
C38427 a_n1151_42308# a_11387_46155# 0.195225f
C38428 a_n743_46660# a_3090_45724# 0.050883f
C38429 a_6545_47178# a_8016_46348# 4.25e-20
C38430 a_4915_47217# a_8953_45546# 1.73e-19
C38431 a_6151_47436# a_8349_46414# 1.15e-19
C38432 a_4883_46098# a_12741_44636# 0.076276f
C38433 a_6031_43396# a_5837_42852# 5.29e-20
C38434 a_10341_43396# a_18599_43230# 1.21e-19
C38435 a_n2840_42826# a_n2157_42858# 7.58e-21
C38436 a_11827_44484# VDD 0.615802f
C38437 a_n2438_43548# a_n3674_38680# 8.18e-20
C38438 a_14180_45002# a_13720_44458# 4.96e-19
C38439 a_1423_45028# a_8103_44636# 0.064947f
C38440 a_16922_45042# a_17719_45144# 0.22253f
C38441 a_17023_45118# a_17613_45144# 0.001643f
C38442 a_n2293_45010# a_n2293_43922# 0.00103f
C38443 a_n2017_45002# a_n2661_42834# 0.037965f
C38444 a_10227_46804# a_15486_42560# 0.227612f
C38445 a_10903_43370# a_10849_43646# 0.003042f
C38446 a_1307_43914# a_10440_44484# 5.64e-20
C38447 a_9482_43914# a_14539_43914# 2.22e-19
C38448 a_13556_45296# a_16112_44458# 0.001671f
C38449 a_526_44458# a_548_43396# 0.002535f
C38450 a_n467_45028# a_n310_44484# 2.23e-19
C38451 a_7499_43078# a_8333_44056# 0.005667f
C38452 a_18175_45572# a_18579_44172# 5.04e-22
C38453 a_3483_46348# a_15743_43084# 8.98e-20
C38454 a_11415_45002# a_22591_43396# 1.64e-20
C38455 a_n2312_38680# a_n3674_38216# 0.023419f
C38456 a_n2442_46660# COMP_P 0.024155f
C38457 a_2711_45572# a_11341_43940# 1.54309f
C38458 a_5009_45028# a_n2661_44458# 0.002424f
C38459 a_13885_46660# a_3483_46348# 2.24e-19
C38460 a_11599_46634# a_11823_42460# 5.18e-19
C38461 a_n743_46660# a_15002_46116# 1.44e-19
C38462 a_21188_46660# a_12741_44636# 0.052893f
C38463 a_22000_46634# a_20820_30879# 0.001417f
C38464 a_5907_46634# a_5066_45546# 9.12e-19
C38465 a_768_44030# a_3316_45546# 5.1e-21
C38466 a_6755_46942# a_10809_44734# 0.042402f
C38467 a_12991_46634# a_12594_46348# 7.99e-21
C38468 a_12861_44030# a_13904_45546# 0.027907f
C38469 a_n881_46662# a_2277_45546# 1.72e-20
C38470 a_20841_46902# a_21297_46660# 4.2e-19
C38471 a_10227_46804# a_10053_45546# 0.009863f
C38472 a_743_42282# a_13333_42558# 0.001019f
C38473 a_19164_43230# a_19326_42852# 0.006453f
C38474 a_20922_43172# a_22400_42852# 1.28e-20
C38475 a_4190_30871# a_14113_42308# 6.14e-20
C38476 a_17499_43370# a_17531_42308# 9.86e-20
C38477 a_17324_43396# a_17303_42282# 2.04e-20
C38478 a_4361_42308# a_12563_42308# 0.009982f
C38479 a_5649_42852# a_5742_30871# 0.059614f
C38480 a_14537_43396# a_15301_44260# 2.79e-19
C38481 a_16763_47508# RST_Z 2.3e-19
C38482 a_n2433_44484# a_n1899_43946# 2.69e-19
C38483 a_n2661_44458# a_n1331_43914# 8.46e-21
C38484 a_16588_47582# VDD 0.282243f
C38485 a_13259_45724# a_19339_43156# 7.95e-21
C38486 a_n2293_46098# a_6171_42473# 1.9e-21
C38487 a_8696_44636# a_9145_43396# 2.59e-20
C38488 en_comp a_n2433_43396# 0.036527f
C38489 a_5608_44484# a_5708_44484# 0.005294f
C38490 a_n89_44484# a_n2661_42834# 2.61e-19
C38491 a_n2267_44484# a_n2065_43946# 1.98e-19
C38492 a_n2129_44697# a_n1761_44111# 5.53e-19
C38493 a_n443_42852# a_685_42968# 0.104532f
C38494 a_12861_44030# CLK 4.17e-19
C38495 a_1823_45246# a_2713_42308# 2.25e-19
C38496 a_n755_45592# a_8605_42826# 0.003535f
C38497 a_n357_42282# a_8387_43230# 0.009479f
C38498 a_n2661_43370# a_9028_43914# 5.67e-21
C38499 a_n2017_45002# a_n1352_43396# 8.78e-19
C38500 a_n2293_45010# a_n97_42460# 4.81e-19
C38501 a_n310_44484# a_n2661_43922# 1.2e-19
C38502 a_9313_44734# a_n2293_43922# 0.026681f
C38503 a_18248_44752# a_18588_44850# 0.027606f
C38504 a_17767_44458# a_11967_42832# 0.003339f
C38505 a_5204_45822# a_n2661_45546# 5.48e-19
C38506 a_n2293_46634# a_3537_45260# 0.155982f
C38507 a_13059_46348# a_11962_45724# 0.001121f
C38508 a_10227_46804# a_13490_45394# 1.9e-20
C38509 a_13759_46122# a_14383_46116# 9.73e-19
C38510 a_14275_46494# a_14537_46482# 0.001705f
C38511 a_14493_46090# a_14949_46494# 4.2e-19
C38512 a_12891_46348# a_14537_43396# 5.09e-20
C38513 a_167_45260# a_997_45618# 0.052039f
C38514 a_2521_46116# a_n755_45592# 3.63e-20
C38515 a_n2293_46098# a_1990_45899# 6.77e-19
C38516 a_n746_45260# a_n452_44636# 0.042999f
C38517 a_5807_45002# a_8953_45002# 7.32e-20
C38518 a_n133_46660# a_327_44734# 9.06e-21
C38519 a_n2438_43548# a_1667_45002# 0.001763f
C38520 a_n2661_46098# a_n2293_45010# 1.46e-20
C38521 a_4883_46098# a_n2293_42834# 2.72e-20
C38522 a_13351_46090# a_13259_45724# 7.81e-20
C38523 a_768_44030# a_13777_45326# 0.011242f
C38524 a_33_46660# a_n37_45144# 3.74e-22
C38525 a_n2661_46634# a_5147_45002# 2.08e-20
C38526 a_14180_46812# a_13904_45546# 2.21e-22
C38527 a_13885_46660# a_14495_45572# 1.27e-20
C38528 a_765_45546# a_9049_44484# 2.74e-20
C38529 a_10809_44734# a_8049_45260# 0.059599f
C38530 a_1823_45246# a_2957_45546# 0.009473f
C38531 a_7963_42308# a_5742_30871# 1.16e-20
C38532 a_4190_30871# C8_N_btm 4.06e-19
C38533 COMP_P a_13258_32519# 0.010297f
C38534 a_8685_42308# a_9293_42558# 0.003228f
C38535 a_13467_32519# C2_N_btm 0.001797f
C38536 a_16823_43084# RST_Z 5.98e-22
C38537 a_3357_43084# a_4649_43172# 1.01e-20
C38538 a_10057_43914# a_8791_43396# 2.04e-20
C38539 a_n2293_42834# a_5649_42852# 0.002922f
C38540 a_11827_44484# a_16137_43396# 8.22e-20
C38541 a_1307_43914# a_1847_42826# 0.428505f
C38542 a_18114_32519# a_10341_43396# 4.67e-19
C38543 a_13259_45724# a_22465_38105# 1.69e-19
C38544 a_22485_44484# a_11341_43940# 0.006131f
C38545 a_20512_43084# a_22223_43948# 0.001071f
C38546 a_9313_44734# a_n97_42460# 1.76217f
C38547 a_n356_44636# a_1427_43646# 0.00321f
C38548 a_5663_43940# a_n2661_42282# 0.00715f
C38549 a_18587_45118# a_18525_43370# 1.2e-22
C38550 a_18184_42460# a_17499_43370# 2.47e-20
C38551 a_14180_46812# CLK 1.54e-20
C38552 en_comp a_21356_42826# 4.89e-21
C38553 a_n443_42852# a_14113_42308# 3.7e-20
C38554 a_n913_45002# a_22223_42860# 0.011179f
C38555 a_n2017_45002# a_n2293_42282# 0.095773f
C38556 a_375_42282# a_685_42968# 2.44e-19
C38557 a_5204_45822# a_5205_44484# 2.74e-21
C38558 a_12549_44172# a_20679_44626# 0.006058f
C38559 a_17715_44484# a_n2017_45002# 7.39e-21
C38560 a_3483_46348# a_10775_45002# 0.025931f
C38561 a_13661_43548# a_16241_44484# 5.03e-19
C38562 a_5937_45572# a_4558_45348# 1.53e-20
C38563 a_22223_46124# a_3357_43084# 2.09e-20
C38564 a_15227_44166# a_11691_44458# 0.443265f
C38565 a_19692_46634# a_22223_45036# 8.92e-20
C38566 a_6165_46155# a_6171_45002# 9.99e-20
C38567 a_10903_43370# a_413_45260# 4.56e-21
C38568 a_13259_45724# a_15225_45822# 7.2e-20
C38569 a_6472_45840# a_6667_45809# 0.215953f
C38570 a_6194_45824# a_6598_45938# 0.051162f
C38571 a_n443_42852# a_7499_43078# 0.375366f
C38572 a_2107_46812# a_9159_44484# 5.96e-19
C38573 a_1736_39587# a_2113_38308# 0.100626f
C38574 a_n4209_39304# a_n4064_37984# 0.029462f
C38575 a_5932_42308# C4_N_btm 0.032349f
C38576 a_6151_47436# a_10227_46804# 0.032659f
C38577 a_1606_42308# VIN_N 0.014401f
C38578 a_13717_47436# a_12861_44030# 0.319645f
C38579 a_n1435_47204# a_13487_47204# 0.135076f
C38580 a_1239_39043# a_1177_38525# 0.031327f
C38581 a_n4209_38502# a_n3420_38528# 0.230544f
C38582 a_n3565_39304# a_n3420_37984# 0.028129f
C38583 a_n4064_39072# a_n4209_38216# 0.03057f
C38584 a_n3420_39072# a_n3565_38216# 0.030682f
C38585 a_n4334_38528# a_n3690_38528# 8.67e-19
C38586 a_5934_30871# C0_P_btm 0.015126f
C38587 a_n971_45724# a_n310_47243# 0.007307f
C38588 a_n452_47436# a_7_47243# 6.64e-19
C38589 a_3581_42558# VDD 0.006789f
C38590 a_6123_31319# C0_dummy_N_btm 1.31e-19
C38591 a_16522_42674# CAL_N 2.6e-20
C38592 a_3160_47472# a_4883_46098# 1.62e-19
C38593 en_comp a_n4064_40160# 1.93e-20
C38594 a_n2956_37592# a_n2302_40160# 0.006106f
C38595 a_7_45899# VDD 0.001958f
C38596 a_12429_44172# a_12281_43396# 1.87e-20
C38597 a_17737_43940# a_10341_43396# 4.05e-20
C38598 a_n2293_42834# a_7963_42308# 7.42e-19
C38599 a_1307_43914# a_15486_42560# 9.69e-21
C38600 a_3065_45002# a_7174_31319# 4.88e-21
C38601 a_n2433_43396# a_n1699_43638# 0.062578f
C38602 a_n2129_43609# a_n2267_43396# 0.230013f
C38603 a_n4318_39304# a_n1917_43396# 1.69e-19
C38604 a_15493_43940# a_8685_43396# 6.24e-19
C38605 a_13747_46662# a_2982_43646# 0.010585f
C38606 a_5807_45002# a_3626_43646# 2.2e-22
C38607 a_11415_45002# a_22591_44484# 6.11e-19
C38608 a_8696_44636# a_n1059_45260# 2.7e-21
C38609 a_12465_44636# a_10341_43396# 8.52e-20
C38610 a_11453_44696# a_14205_43396# 1.6e-22
C38611 a_n971_45724# a_n901_43156# 0.019025f
C38612 SMPL_ON_P a_n4318_38680# 0.039103f
C38613 a_n443_46116# a_743_42282# 1.1e-19
C38614 a_768_44030# a_6197_43396# 4.37e-20
C38615 a_13163_45724# a_13017_45260# 2.76e-20
C38616 a_1609_45822# a_n2661_43370# 0.008983f
C38617 a_2324_44458# a_3363_44484# 0.004792f
C38618 a_10907_45822# a_3232_43370# 4.17e-19
C38619 a_16327_47482# a_16409_43396# 0.022593f
C38620 a_5263_45724# a_5093_45028# 4.44e-20
C38621 a_11823_42460# a_13348_45260# 4.52e-20
C38622 a_8049_45260# a_5883_43914# 3.03e-20
C38623 a_n357_42282# a_16922_45042# 9.6e-19
C38624 a_10227_46804# a_13837_43396# 1.96e-20
C38625 a_3090_45724# a_11750_44172# 3.43e-21
C38626 a_2711_45572# a_7418_45394# 9.37e-20
C38627 a_12861_44030# a_19268_43646# 9.01e-21
C38628 a_19256_45572# a_20528_45572# 1.03e-20
C38629 C10_P_btm C6_P_btm 0.421276f
C38630 a_383_46660# a_1799_45572# 2.74e-20
C38631 a_601_46902# a_n2661_46098# 0.003957f
C38632 a_9804_47204# a_10428_46928# 3.61e-20
C38633 VDAC_N VREF 0.254986f
C38634 a_n881_46662# a_6755_46942# 0.063288f
C38635 a_12861_44030# a_14035_46660# 0.153051f
C38636 a_13717_47436# a_14180_46812# 1e-20
C38637 a_13487_47204# a_13885_46660# 0.002202f
C38638 a_n1613_43370# a_6969_46634# 3.94e-19
C38639 a_11453_44696# a_11813_46116# 5.74e-21
C38640 a_13507_46334# a_15009_46634# 7.3e-20
C38641 a_18597_46090# a_17609_46634# 8.28e-19
C38642 C9_P_btm C7_P_btm 0.227839f
C38643 a_n743_46660# a_3699_46634# 1.08e-19
C38644 a_n2438_43548# a_2959_46660# 3.53e-20
C38645 a_5815_47464# a_765_45546# 0.01398f
C38646 VDAC_P VIN_P 0.252066f
C38647 a_22780_39857# VDD 2.73e-20
C38648 a_n1925_46634# a_2864_46660# 0.004284f
C38649 a_18780_47178# a_18834_46812# 0.010748f
C38650 a_18479_47436# a_15227_44166# 0.199537f
C38651 a_10227_46804# a_19466_46812# 1.18e-19
C38652 a_3905_42865# a_4921_42308# 1.92e-19
C38653 a_19268_43646# a_19700_43370# 0.017165f
C38654 a_16243_43396# a_16823_43084# 0.05964f
C38655 a_15743_43084# a_16664_43396# 0.01372f
C38656 a_16977_43638# a_17486_43762# 2.6e-19
C38657 a_16409_43396# a_16855_43396# 2.28e-19
C38658 a_3626_43646# a_10518_42984# 2.25e-20
C38659 a_2982_43646# a_10796_42968# 8.58e-20
C38660 a_15595_45028# VDD 0.156299f
C38661 a_n97_42460# a_18599_43230# 0.006824f
C38662 a_10341_43396# a_13887_32519# 0.030175f
C38663 a_6197_43396# a_5755_42852# 4.26e-20
C38664 a_3090_45724# a_4361_42308# 1.2e-19
C38665 a_4791_45118# a_6171_42473# 5.34e-19
C38666 a_n863_45724# a_1241_44260# 1.7e-19
C38667 a_1823_45246# a_6031_43396# 3.31e-19
C38668 a_n1059_45260# a_n1177_44458# 9.59e-19
C38669 a_n2293_45010# a_742_44458# 3.27e-20
C38670 a_n2661_45010# a_2779_44458# 4.72e-20
C38671 SMPL_ON_N a_14097_32519# 0.029158f
C38672 a_15227_44166# a_4190_30871# 2.91e-20
C38673 a_12741_44636# a_8685_43396# 5.43e-21
C38674 a_14797_45144# a_14976_45348# 0.007688f
C38675 a_14537_43396# a_15060_45348# 0.001339f
C38676 en_comp a_n2433_44484# 0.029809f
C38677 a_n967_45348# a_n2661_44458# 0.0255f
C38678 a_13259_45724# a_17973_43940# 0.025372f
C38679 a_9482_43914# a_14309_45028# 3.6e-19
C38680 a_13556_45296# a_13807_45067# 2.63e-19
C38681 a_13507_46334# a_19431_46494# 0.001128f
C38682 a_4817_46660# a_5497_46414# 0.001967f
C38683 a_5167_46660# a_5164_46348# 0.003259f
C38684 a_5385_46902# a_5204_45822# 1.84e-20
C38685 a_18834_46812# a_18285_46348# 0.144972f
C38686 a_13885_46660# a_14513_46634# 0.101344f
C38687 a_14035_46660# a_14180_46812# 0.00994f
C38688 a_15227_44166# a_17829_46910# 1.41e-19
C38689 a_17609_46634# a_19123_46287# 1.84e-20
C38690 a_19466_46812# a_17339_46660# 1.16e-20
C38691 a_9804_47204# a_8283_46482# 3.67e-21
C38692 a_8128_46384# a_8034_45724# 0.003967f
C38693 a_n881_46662# a_8049_45260# 0.025172f
C38694 a_n443_46116# a_2277_45546# 0.048113f
C38695 a_4646_46812# a_7920_46348# 2.09e-20
C38696 a_n971_45724# a_3733_45822# 3.4e-19
C38697 a_2063_45854# a_4099_45572# 1.09e-19
C38698 a_n237_47217# a_3775_45552# 1.02e-19
C38699 a_768_44030# a_5066_45546# 2.81e-20
C38700 a_n2661_46634# a_n2956_39304# 4.64e-19
C38701 a_n2956_39768# a_n2956_38680# 0.043291f
C38702 a_18479_47436# a_21071_46482# 5.89e-19
C38703 a_4883_46098# a_16375_45002# 0.01007f
C38704 a_3422_30871# C3_N_btm 1.1e-19
C38705 a_21195_42852# a_21671_42860# 0.177876f
C38706 a_21356_42826# a_22165_42308# 5.1e-21
C38707 a_22959_43396# a_14097_32519# 0.00104f
C38708 a_2982_43646# a_4958_30871# 0.136637f
C38709 a_3626_43646# a_16197_42308# 7.17e-19
C38710 a_8037_42858# a_9114_42852# 1.46e-19
C38711 a_8685_43396# a_5742_30871# 4.78e-19
C38712 a_17364_32525# a_22400_42852# 1.05e-20
C38713 a_1307_43914# a_5244_44056# 0.025291f
C38714 a_n2840_44458# a_n2661_42834# 8.29e-19
C38715 a_11827_44484# a_13940_44484# 4.46e-19
C38716 a_n357_42282# a_15743_43084# 0.055032f
C38717 a_n443_42852# a_15781_43660# 0.22553f
C38718 a_n2442_46660# a_n4209_39304# 2.66e-20
C38719 a_6298_44484# a_7640_43914# 0.031665f
C38720 a_5343_44458# a_5891_43370# 1.06553f
C38721 a_n2661_44458# a_9159_44484# 1.56e-19
C38722 a_18494_42460# a_17517_44484# 0.022635f
C38723 a_3232_43370# a_n2661_42282# 0.005579f
C38724 a_18248_44752# a_18443_44721# 0.206455f
C38725 a_17970_44736# a_18374_44850# 0.051162f
C38726 a_17767_44458# a_18989_43940# 3.82e-21
C38727 a_n452_44636# a_n310_44484# 0.007833f
C38728 a_2711_45572# a_10341_43396# 0.03441f
C38729 a_526_44458# a_10083_42826# 0.012145f
C38730 a_n1613_43370# a_3357_43084# 0.228593f
C38731 a_n2312_40392# a_n2956_37592# 0.060336f
C38732 a_14275_46494# a_2324_44458# 5.45e-20
C38733 a_15015_46420# a_14840_46494# 0.233657f
C38734 a_3483_46348# a_526_44458# 0.134907f
C38735 a_10150_46912# a_10193_42453# 1.25e-20
C38736 a_9863_46634# a_8746_45002# 5.88e-19
C38737 a_10467_46802# a_10053_45546# 1.61e-20
C38738 a_n443_46116# a_626_44172# 2.44e-20
C38739 a_19594_46812# a_19256_45572# 2.98e-19
C38740 a_12549_44172# a_20528_45572# 1.17e-19
C38741 a_n2312_39304# a_n2810_45028# 0.043636f
C38742 a_15227_44166# a_n443_42852# 0.023429f
C38743 a_167_45260# a_1337_46116# 2.67e-20
C38744 a_9569_46155# a_6945_45028# 3.28e-20
C38745 a_10227_46804# a_5111_44636# 7.06e-20
C38746 a_4883_46098# a_413_45260# 2.47e-19
C38747 a_1755_42282# a_2123_42473# 0.014573f
C38748 a_14635_42282# a_14113_42308# 0.052122f
C38749 a_8147_43396# VDD 0.393534f
C38750 a_1184_42692# a_2713_42308# 4.61e-20
C38751 a_1606_42308# a_2351_42308# 0.191324f
C38752 a_n2472_43914# a_n1761_44111# 1.8e-19
C38753 a_3537_45260# a_743_42282# 0.033447f
C38754 a_n2293_45010# a_n901_43156# 2.97e-20
C38755 a_n2661_45010# a_n13_43084# 4.49e-21
C38756 a_n2017_45002# a_n1423_42826# 0.008318f
C38757 a_n913_45002# a_n1853_43023# 0.094845f
C38758 a_n1059_45260# a_n1991_42858# 8.68e-20
C38759 a_n2293_42834# a_8685_43396# 1.23e-19
C38760 a_n2129_44697# a_n2267_43396# 1.8e-20
C38761 a_n357_42282# a_1606_42308# 0.001349f
C38762 a_10057_43914# a_10651_43940# 0.003719f
C38763 a_10150_46912# VDD 0.284144f
C38764 a_13857_44734# a_13483_43940# 3.4e-20
C38765 a_7411_46660# DATA[3] 7.26e-20
C38766 a_9313_44734# a_21115_43940# 9.92e-21
C38767 a_n2661_45546# a_3823_42558# 7.7e-21
C38768 a_16327_47482# a_16241_44734# 4.54e-20
C38769 a_380_45546# a_n357_42282# 0.071576f
C38770 a_n2661_45546# a_3503_45724# 0.006856f
C38771 a_5807_45002# a_17767_44458# 1.7e-21
C38772 a_13925_46122# a_8696_44636# 7.96e-21
C38773 a_21188_46660# a_413_45260# 4.93e-21
C38774 a_n2293_46098# a_3357_43084# 0.16657f
C38775 a_n452_45724# a_n755_45592# 0.03904f
C38776 a_n1099_45572# a_310_45028# 0.333219f
C38777 a_n863_45724# a_997_45618# 3.46e-19
C38778 a_13747_46662# a_14539_43914# 1.14e-20
C38779 a_13661_43548# a_16979_44734# 5.5e-20
C38780 a_15682_46116# a_15903_45785# 0.011633f
C38781 a_2324_44458# a_15765_45572# 0.005634f
C38782 a_n2497_47436# a_895_43940# 0.0309f
C38783 a_n971_45724# a_n984_44318# 0.003098f
C38784 a_n746_45260# a_n809_44244# 1.75e-19
C38785 a_10903_43370# a_12561_45572# 0.002063f
C38786 a_8049_45260# a_8162_45546# 0.057007f
C38787 a_n743_46660# a_4743_44484# 1.08e-21
C38788 a_12465_44636# a_n2293_43922# 0.025736f
C38789 COMP_P a_22609_37990# 0.010152f
C38790 a_n4064_40160# a_n2216_40160# 0.005638f
C38791 a_6123_31319# VDAC_Ni 4.39e-19
C38792 a_n4334_40480# a_n4209_39590# 6.38e-20
C38793 a_n4315_30879# a_n4334_39616# 6.38e-20
C38794 SMPL_ON_P a_n1151_42308# 2.27e-19
C38795 a_n785_47204# a_1431_47204# 6.54e-19
C38796 a_n2109_47186# a_3815_47204# 0.045952f
C38797 a_n1741_47186# a_3381_47502# 0.011573f
C38798 a_327_47204# a_1239_47204# 6.56e-19
C38799 a_n971_45724# a_2553_47502# 0.23907f
C38800 a_n237_47217# a_584_46384# 0.645142f
C38801 a_1606_42308# CAL_N 0.006757f
C38802 a_2889_44172# a_2813_43396# 4.01e-20
C38803 a_11967_42832# a_18525_43370# 0.010117f
C38804 a_13076_44458# a_12379_42858# 1.36e-20
C38805 a_12607_44458# a_12545_42858# 5.22e-21
C38806 a_21115_43940# a_20974_43370# 2.85e-19
C38807 a_11341_43940# a_14401_32519# 0.008534f
C38808 a_15493_43940# a_19741_43940# 0.027038f
C38809 a_3537_45260# a_5755_42308# 0.002651f
C38810 a_5147_45002# a_4921_42308# 2e-19
C38811 a_n2017_45002# a_9885_42558# 0.006803f
C38812 a_n913_45002# a_9293_42558# 2.08e-19
C38813 a_17737_43940# a_n97_42460# 1.26e-20
C38814 a_n2661_42282# a_4905_42826# 5.42e-20
C38815 a_3232_43370# a_3497_42558# 7.4e-20
C38816 a_3065_45002# a_5932_42308# 4.34e-21
C38817 a_22485_44484# a_10341_43396# 4.73e-20
C38818 en_comp a_8685_42308# 4.34e-21
C38819 a_n356_44636# a_4520_42826# 2.14e-20
C38820 a_3483_46348# a_17970_44736# 1.12e-19
C38821 a_16333_45814# a_16115_45572# 0.209641f
C38822 a_n443_46116# a_2813_43396# 0.124521f
C38823 a_n971_45724# a_9885_43646# 9.07e-21
C38824 a_22612_30879# a_14021_43940# 1.68e-20
C38825 a_8199_44636# a_10157_44484# 5.53e-20
C38826 a_8953_45546# a_5883_43914# 0.262126f
C38827 a_8016_46348# a_10440_44484# 0.001273f
C38828 a_15599_45572# a_8696_44636# 5.37e-19
C38829 a_15765_45572# a_16855_45546# 0.042415f
C38830 a_15903_45785# a_16680_45572# 5.47e-21
C38831 a_19466_46812# a_18579_44172# 0.003312f
C38832 a_n1151_42308# a_8035_47026# 6.49e-20
C38833 VDAC_P a_11206_38545# 0.101449f
C38834 a_8912_37509# CAL_N 0.017398f
C38835 a_6575_47204# a_7927_46660# 1.99e-19
C38836 a_4791_45118# a_6969_46634# 0.001756f
C38837 a_6151_47436# a_10467_46802# 2.6e-19
C38838 a_4915_47217# a_10249_46116# 0.001348f
C38839 a_n4209_38216# VDD 0.833976f
C38840 a_n1613_43370# a_n2293_46634# 0.103089f
C38841 a_n881_46662# a_n2442_46660# 1.71e-20
C38842 a_9313_45822# a_7411_46660# 1.38e-19
C38843 a_12549_44172# a_19594_46812# 7.14e-20
C38844 a_19479_31679# C6_N_btm 1.26e-20
C38845 a_n2433_43396# a_n2157_42858# 2.73e-19
C38846 a_9145_43396# a_14205_43396# 0.13322f
C38847 a_19963_31679# C3_N_btm 0.041776f
C38848 a_20365_43914# a_19987_42826# 4.65e-20
C38849 a_15493_43940# a_17333_42852# 1.29e-20
C38850 a_19237_31679# a_22400_42852# 2.13e-20
C38851 a_21350_45938# VDD 7.19e-19
C38852 a_14539_43914# a_4958_30871# 0.00214f
C38853 a_n2293_43922# a_8515_42308# 3.54e-20
C38854 a_9313_44734# a_10533_42308# 8.54e-19
C38855 a_19862_44208# a_21356_42826# 0.001265f
C38856 a_4099_45572# a_n2661_42834# 4.28e-22
C38857 a_10907_45822# a_8975_43940# 1.46e-19
C38858 a_20202_43084# a_17538_32519# 2.29e-20
C38859 a_3065_45002# a_1423_45028# 0.017813f
C38860 a_5111_44636# a_1307_43914# 0.114933f
C38861 a_12891_46348# a_12379_42858# 0.001173f
C38862 SMPL_ON_P a_n2840_42282# 6.32e-19
C38863 a_6171_45002# a_14797_45144# 0.00824f
C38864 a_18189_46348# a_17973_43940# 4.22e-19
C38865 a_n2438_43548# a_n4318_38680# 0.001622f
C38866 a_18479_45785# a_11827_44484# 0.03055f
C38867 a_17715_44484# a_18079_43940# 4.31e-19
C38868 a_2274_45254# a_2809_45348# 9.76e-19
C38869 a_2382_45260# a_2304_45348# 0.045704f
C38870 a_3090_45724# a_7274_43762# 1.37e-19
C38871 a_18780_47178# a_10809_44734# 0.002996f
C38872 a_n2293_46634# a_n2293_46098# 0.062583f
C38873 a_11453_44696# a_15682_46116# 1.17e-20
C38874 a_13507_46334# a_19335_46494# 0.004216f
C38875 a_20894_47436# a_20708_46348# 1.02e-19
C38876 a_n1151_42308# a_11387_46482# 0.005536f
C38877 a_8128_46384# a_8016_46348# 0.09182f
C38878 a_n881_46662# a_8953_45546# 1.01e-19
C38879 a_19386_47436# a_6945_45028# 0.008586f
C38880 a_4883_46098# a_18985_46122# 0.027089f
C38881 a_6151_47436# a_8034_45724# 9.18e-19
C38882 a_n2661_46634# a_n1991_46122# 9.31e-19
C38883 a_n2312_38680# a_n2840_46090# 0.003997f
C38884 a_7_44811# VDD 0.001865f
C38885 a_3422_30871# a_7754_38470# 6.77e-20
C38886 a_22959_43948# a_22775_42308# 3.38e-21
C38887 a_n97_42460# a_8515_42308# 2.07e-19
C38888 a_3080_42308# a_3581_42558# 3.31e-19
C38889 a_22959_43396# a_22959_42860# 0.026152f
C38890 a_8387_43230# a_8952_43230# 7.99e-20
C38891 a_8037_42858# a_10518_42984# 2e-20
C38892 a_2711_45572# a_n97_42460# 0.137121f
C38893 a_n863_45724# a_648_43396# 6.1e-19
C38894 a_17719_45144# a_17970_44736# 4.66e-19
C38895 a_8560_45348# a_5891_43370# 7.06e-20
C38896 a_4185_45028# a_7765_42852# 1.44e-20
C38897 a_20202_43084# a_19339_43156# 2.42e-20
C38898 a_n357_42282# a_3539_42460# 0.019382f
C38899 a_n755_45592# a_3626_43646# 0.095572f
C38900 a_n2661_44458# a_n1917_44484# 0.008101f
C38901 a_n2433_44484# a_n1699_44726# 0.058433f
C38902 a_16922_45042# a_18443_44721# 6.14e-20
C38903 a_n2661_43370# a_5205_44734# 1.1e-19
C38904 a_11827_44484# a_10057_43914# 2.12e-19
C38905 a_n2956_37592# a_n2472_43914# 9.42e-21
C38906 a_n2312_39304# a_n2302_40160# 3.32e-19
C38907 a_n1059_45260# a_n1331_43914# 4.5e-20
C38908 a_n913_45002# a_n1899_43946# 0.017336f
C38909 a_n745_45366# a_n1761_44111# 5.25e-20
C38910 a_n2661_45010# a_644_44056# 8.47e-20
C38911 a_n2017_45002# a_n1549_44318# 9.31e-19
C38912 a_n2293_45010# a_n984_44318# 0.048428f
C38913 a_n2129_44697# a_n2267_44484# 0.698671f
C38914 a_14797_45144# a_14673_44172# 9.74e-20
C38915 a_n443_42852# a_1756_43548# 0.006388f
C38916 a_7499_43078# a_11257_43940# 6.52e-20
C38917 a_16327_47482# a_18691_45572# 0.162157f
C38918 a_n2661_46634# a_7499_43078# 3.96e-20
C38919 a_n2497_47436# a_3065_45002# 0.022803f
C38920 a_1823_45246# a_4419_46090# 0.340207f
C38921 a_4791_45118# a_3357_43084# 0.144996f
C38922 a_11453_44696# a_16680_45572# 2.06e-21
C38923 a_10227_46804# a_16147_45260# 0.001138f
C38924 a_20411_46873# a_20708_46348# 0.081063f
C38925 a_20273_46660# a_19900_46494# 3.92e-19
C38926 a_20107_46660# a_21137_46414# 0.001469f
C38927 a_11901_46660# a_12638_46436# 4.56e-19
C38928 a_12469_46902# a_12379_46436# 5.5e-19
C38929 a_18285_46348# a_10809_44734# 0.014976f
C38930 a_5129_47502# a_2437_43646# 0.004f
C38931 a_584_46384# a_n2017_45002# 4e-20
C38932 a_n746_45260# a_n955_45028# 2.13e-20
C38933 a_n971_45724# a_n467_45028# 2.65e-20
C38934 a_167_45260# a_3699_46348# 4.42e-20
C38935 a_2521_46116# a_3483_46348# 1.75e-19
C38936 a_2698_46116# a_3147_46376# 0.003074f
C38937 a_17609_46634# a_8049_45260# 1.64e-21
C38938 a_11415_45002# a_12594_46348# 1.51e-20
C38939 a_5807_45002# a_12791_45546# 7.66e-21
C38940 a_13661_43548# a_11823_42460# 0.116839f
C38941 a_1799_45572# a_3175_45822# 6.77e-21
C38942 a_2107_46812# a_6598_45938# 1.55e-20
C38943 a_5534_30871# a_13657_42558# 1.73e-19
C38944 a_10555_43940# VDD 0.002652f
C38945 a_5807_45002# DATA[4] 3.14e-21
C38946 a_11827_44484# a_14021_43940# 3.51e-19
C38947 a_21588_30879# VDD 1.78413f
C38948 a_626_44172# a_1049_43396# 2.99e-19
C38949 a_5883_43914# a_9028_43914# 0.05428f
C38950 a_20916_46384# RST_Z 3.17e-20
C38951 a_11823_42460# a_10835_43094# 0.006753f
C38952 a_20843_47204# SINGLE_ENDED 0.007105f
C38953 a_10193_42453# a_13113_42826# 4.41e-21
C38954 a_n357_42282# a_9061_43230# 7.05e-20
C38955 a_n755_45592# a_8649_43218# 1.17e-19
C38956 a_n1925_42282# a_2123_42473# 5.44e-20
C38957 a_9290_44172# a_12563_42308# 0.052279f
C38958 a_20202_43084# a_22465_38105# 1.3e-19
C38959 a_1307_43914# a_4235_43370# 0.016608f
C38960 a_17517_44484# a_20640_44752# 0.54753f
C38961 a_5205_44484# a_6765_43638# 8.52e-19
C38962 a_5147_45002# a_6452_43396# 2.05e-19
C38963 a_5111_44636# a_9396_43370# 0.203348f
C38964 a_n2017_45002# a_15095_43370# 0.002423f
C38965 a_n1059_45260# a_14205_43396# 4.2e-20
C38966 a_n913_45002# a_14358_43442# 3.05e-20
C38967 a_526_44458# a_2351_42308# 8.58e-19
C38968 a_n443_42852# a_5193_43172# 4.01e-19
C38969 a_10227_46804# a_10334_44484# 0.020432f
C38970 a_11599_46634# a_14539_43914# 5.29e-21
C38971 a_2324_44458# a_6194_45824# 0.001699f
C38972 a_13747_46662# a_14309_45028# 1.11e-19
C38973 a_7411_46660# a_7705_45326# 2.02e-20
C38974 a_13661_43548# a_16321_45348# 3.11e-19
C38975 a_n746_45260# a_n2661_42834# 0.01463f
C38976 a_n971_45724# a_n2661_43922# 0.052944f
C38977 a_4791_45118# a_5826_44734# 3.51e-20
C38978 a_16292_46812# a_3357_43084# 1.44e-20
C38979 a_3483_46348# a_13163_45724# 5.34e-20
C38980 a_8016_46348# a_10053_45546# 0.017312f
C38981 a_12861_44030# a_18248_44752# 0.072535f
C38982 a_15227_44166# a_2437_43646# 0.167451f
C38983 a_17339_46660# a_16147_45260# 0.006901f
C38984 a_11415_45002# a_15037_45618# 5.65e-19
C38985 a_12549_44172# a_18494_42460# 0.331306f
C38986 a_4185_45028# a_11823_42460# 3.07e-19
C38987 a_8199_44636# a_7499_43078# 0.859274f
C38988 a_5937_45572# a_8568_45546# 0.028968f
C38989 a_7715_46873# a_6709_45028# 3.14e-19
C38990 a_7577_46660# a_7229_43940# 1.48e-22
C38991 a_8049_45260# a_19443_46116# 0.001302f
C38992 a_526_44458# a_n357_42282# 0.220537f
C38993 a_5342_30871# C5_N_btm 9.85e-20
C38994 a_13575_42558# a_7174_31319# 4.88e-21
C38995 a_5534_30871# C7_N_btm 0.060228f
C38996 a_n4318_37592# a_n4064_37984# 0.050508f
C38997 a_n3674_38216# a_n4251_38304# 8.42e-19
C38998 a_13113_42826# VDD 0.217254f
C38999 a_18443_44721# a_15743_43084# 1.36e-21
C39000 a_18287_44626# a_19268_43646# 6.61e-20
C39001 a_n356_44636# a_16409_43396# 3.54e-20
C39002 a_4419_46090# DATA[2] 2.81e-19
C39003 a_n2661_44458# a_n1853_43023# 1.84e-21
C39004 a_n2433_44484# a_n2157_42858# 1.17e-21
C39005 a_5891_43370# a_8873_43396# 0.001547f
C39006 a_10193_42453# a_18214_42558# 0.028997f
C39007 a_19328_44172# a_19862_44208# 0.002604f
C39008 a_n1899_43946# a_n4318_39304# 2.93e-19
C39009 a_n1761_44111# a_n2433_43396# 5.56e-19
C39010 a_n2065_43946# a_n2129_43609# 7.7e-19
C39011 a_7542_44172# a_8487_44056# 2.54e-20
C39012 a_7845_44172# a_8415_44056# 9.13e-21
C39013 a_6419_46155# VDD 0.094119f
C39014 a_15493_43396# a_19478_44306# 0.154347f
C39015 a_15682_43940# a_11341_43940# 0.021147f
C39016 a_10729_43914# a_10555_44260# 0.038445f
C39017 a_8746_45002# a_10210_45822# 0.013725f
C39018 a_10193_42453# a_10907_45822# 6.45e-20
C39019 a_5937_45572# a_n2661_43370# 0.202031f
C39020 a_3090_45724# a_5891_43370# 0.166094f
C39021 a_11415_45002# a_18114_32519# 0.002006f
C39022 a_20202_43084# a_19721_31679# 3.09e-20
C39023 a_768_44030# a_2537_44260# 1.56e-20
C39024 a_8034_45724# a_5111_44636# 9.19e-22
C39025 a_8568_45546# a_8697_45572# 0.010132f
C39026 a_8162_45546# a_8791_45572# 6.1e-19
C39027 a_2711_45572# a_16020_45572# 0.006155f
C39028 a_7499_43078# a_8192_45572# 9.59e-19
C39029 a_n2438_43548# a_1467_44172# 9.81e-19
C39030 a_10227_46804# a_13565_44260# 8.58e-20
C39031 a_12741_44636# a_18545_45144# 2.26e-19
C39032 a_n2293_46634# a_2675_43914# 0.026226f
C39033 a_13059_46348# a_15004_44636# 2.9e-20
C39034 a_8049_45260# a_3537_45260# 7.55e-20
C39035 a_n2497_47436# a_458_43396# 4.17e-20
C39036 a_n971_45724# a_n447_43370# 0.113797f
C39037 a_2324_44458# a_6517_45366# 0.002583f
C39038 a_n2109_47186# a_3524_46660# 6.67e-20
C39039 a_n1741_47186# a_2959_46660# 3.8e-20
C39040 a_5129_47502# a_n2661_46634# 5.07e-21
C39041 a_4791_45118# a_n2293_46634# 0.030843f
C39042 a_11459_47204# a_5807_45002# 5.3e-20
C39043 a_13487_47204# a_13759_47204# 0.001672f
C39044 a_7174_31319# C3_N_btm 3.5e-20
C39045 a_n4064_40160# C7_P_btm 2.94e-19
C39046 a_15507_47210# a_15928_47570# 0.089677f
C39047 a_n971_45724# a_1799_45572# 2.58e-19
C39048 a_327_47204# a_491_47026# 0.001941f
C39049 a_n746_45260# a_645_46660# 4.3e-19
C39050 a_n1151_42308# a_n2438_43548# 0.093859f
C39051 a_3754_39964# VDAC_Ni 7.07e-21
C39052 a_13258_32519# C6_N_btm 1.87e-19
C39053 a_584_46384# a_1123_46634# 0.370049f
C39054 a_3815_47204# a_n1925_46634# 2.59e-20
C39055 a_15673_47210# a_12549_44172# 3.81e-20
C39056 a_15811_47375# a_768_44030# 9.22e-21
C39057 a_n2312_40392# a_n2312_39304# 0.057374f
C39058 a_19332_42282# RST_Z 4.07e-20
C39059 a_18214_42558# VDD 0.295211f
C39060 a_n3565_38216# a_n2946_37690# 0.001566f
C39061 a_n4064_37984# a_n4334_37440# 9.42e-19
C39062 a_n4209_38216# a_n2302_37690# 0.001686f
C39063 a_n3420_37984# a_n3690_37440# 0.017537f
C39064 a_n2302_37984# a_n4209_37414# 9.15e-19
C39065 a_n2946_37984# a_n3565_37414# 9.15e-19
C39066 a_n3690_38304# a_n3420_37440# 7.84e-19
C39067 a_n4334_38304# a_n4064_37440# 7.84e-19
C39068 VDAC_Pi a_7754_38968# 8.23e-20
C39069 a_3754_39466# a_3754_39134# 0.296258f
C39070 a_n356_44636# a_564_42282# 9.95e-19
C39071 a_1568_43370# a_2437_43396# 7.56e-20
C39072 a_14401_32519# a_10341_43396# 0.133035f
C39073 a_5343_44458# a_6773_42558# 4.65e-20
C39074 a_19862_44208# a_20749_43396# 0.008749f
C39075 a_10907_45822# VDD 0.352181f
C39076 a_11341_43940# a_22223_43396# 0.00507f
C39077 a_n2661_42282# a_2905_42968# 1.83e-20
C39078 a_22223_43948# a_5649_42852# 3.06e-19
C39079 a_15493_43940# a_13678_32519# 7.99e-22
C39080 a_4223_44672# a_6123_31319# 4.56e-21
C39081 a_n1613_43370# a_743_42282# 2.11e-19
C39082 a_3090_45724# a_18533_43940# 5.95e-19
C39083 a_6598_45938# a_n2661_44458# 5.14e-21
C39084 a_12549_44172# a_15940_43402# 1.28e-20
C39085 a_n2293_46634# a_14537_43646# 0.00342f
C39086 a_4646_46812# a_8147_43396# 5.39e-20
C39087 a_12741_44636# a_13483_43940# 9.28e-21
C39088 a_n1059_45260# a_n967_45348# 0.081574f
C39089 a_n913_45002# en_comp 7.44e-20
C39090 a_13661_43548# a_18429_43548# 0.010678f
C39091 a_4915_47217# a_5534_30871# 5.12e-19
C39092 a_n2293_45010# a_n467_45028# 5.33e-20
C39093 a_n2661_45010# a_n37_45144# 6.21e-20
C39094 a_16147_45260# a_1307_43914# 0.150161f
C39095 a_13259_45724# a_9313_44734# 0.048952f
C39096 a_5732_46660# a_7715_46873# 1.03e-20
C39097 a_5907_46634# a_7577_46660# 5.36e-20
C39098 a_5807_45002# a_12925_46660# 9.54e-20
C39099 a_12549_44172# a_16388_46812# 0.03419f
C39100 a_768_44030# a_13059_46348# 0.062321f
C39101 a_n1435_47204# a_3147_46376# 6.37e-21
C39102 a_21496_47436# a_12741_44636# 4.23e-20
C39103 a_6540_46812# a_7411_46660# 5.06e-21
C39104 a_5072_46660# a_5257_43370# 1.51e-20
C39105 a_n1151_42308# a_11133_46155# 0.162011f
C39106 a_4842_47243# a_765_45546# 4.26e-19
C39107 a_n743_46660# a_15009_46634# 1.24e-21
C39108 a_4883_46098# a_20820_30879# 1.84e-19
C39109 a_12465_44636# a_11415_45002# 0.375509f
C39110 a_22223_47212# a_20202_43084# 1.25e-19
C39111 a_6151_47436# a_8016_46348# 1.03e-19
C39112 a_4915_47217# a_5937_45572# 2.78e-20
C39113 a_n97_42460# a_16877_42852# 0.011527f
C39114 a_21381_43940# a_20753_42852# 2.35e-19
C39115 a_11750_44172# a_11633_42558# 6.73e-22
C39116 a_10807_43548# a_12563_42308# 4.73e-21
C39117 a_n2840_42826# a_n2472_42826# 7.52e-19
C39118 a_21359_45002# VDD 0.319372f
C39119 a_n2312_38680# a_n2104_42282# 2.73e-20
C39120 a_13259_45724# a_20974_43370# 2.3e-20
C39121 a_1423_45028# a_6298_44484# 0.103777f
C39122 a_16922_45042# a_17613_45144# 0.10967f
C39123 a_n2293_45010# a_n2661_43922# 0.030818f
C39124 a_n2472_45002# a_n2293_43922# 7.11e-20
C39125 a_10227_46804# a_15051_42282# 0.361922f
C39126 a_768_44030# a_2903_42308# 2.31e-19
C39127 SMPL_ON_P a_n2302_39866# 5.6e-20
C39128 a_13777_45326# a_13720_44458# 1.97e-19
C39129 a_1307_43914# a_10334_44484# 3.55e-20
C39130 a_9482_43914# a_16112_44458# 3.24e-19
C39131 a_13556_45296# a_15004_44636# 0.127354f
C39132 a_7499_43078# a_8018_44260# 9.13e-21
C39133 a_18341_45572# a_19279_43940# 1.85e-20
C39134 a_n2442_46660# a_n4318_37592# 0.023729f
C39135 a_2711_45572# a_21115_43940# 7.44e-20
C39136 a_22612_30879# a_20692_30879# 0.07827f
C39137 a_12816_46660# a_10903_43370# 3.28e-19
C39138 a_n237_47217# a_8696_44636# 4e-22
C39139 a_10227_46804# a_9049_44484# 1.51e-20
C39140 a_11599_46634# a_12427_45724# 1.84e-20
C39141 a_14955_47212# a_11823_42460# 8.49e-21
C39142 a_21188_46660# a_20820_30879# 3.56e-19
C39143 a_21363_46634# a_12741_44636# 0.053741f
C39144 a_5167_46660# a_5066_45546# 1.61e-20
C39145 a_768_44030# a_3218_45724# 3.61e-19
C39146 a_6969_46634# a_6945_45028# 0.017662f
C39147 a_10249_46116# a_10809_44734# 4.78e-19
C39148 a_12251_46660# a_12594_46348# 0.011817f
C39149 a_3090_45724# a_9290_44172# 0.196232f
C39150 a_13717_47436# a_13904_45546# 8.89e-22
C39151 a_12861_44030# a_13527_45546# 0.274077f
C39152 a_n1613_43370# a_2277_45546# 3.18e-21
C39153 a_20273_46660# a_21297_46660# 2.36e-20
C39154 a_16137_43396# a_18214_42558# 0.0459f
C39155 a_743_42282# a_13249_42558# 0.001357f
C39156 a_1847_42826# a_3905_42558# 1.42e-20
C39157 a_5534_30871# COMP_P 0.027557f
C39158 a_20922_43172# a_20836_43172# 0.001377f
C39159 a_n2661_42282# VDD 0.406474f
C39160 a_16823_43084# a_15803_42450# 0.008769f
C39161 a_17499_43370# a_17303_42282# 4.37e-20
C39162 a_13678_32519# a_5742_30871# 0.004679f
C39163 a_5649_42852# a_11323_42473# 5.44e-20
C39164 a_4361_42308# a_11633_42558# 4.09e-20
C39165 a_16327_47482# START 4.67e-19
C39166 a_14537_43396# a_15037_44260# 0.001968f
C39167 a_7229_43940# a_7499_43940# 6.92e-19
C39168 a_16023_47582# RST_Z 1.03e-19
C39169 a_16979_44734# a_11967_42832# 3.65e-19
C39170 a_n2433_44484# a_n1761_44111# 7.96e-20
C39171 a_n2661_44458# a_n1899_43946# 3.15e-20
C39172 a_10193_42453# a_16823_43084# 0.03411f
C39173 a_13259_45724# a_18599_43230# 1.09e-19
C39174 en_comp a_n4318_39304# 1.82e-19
C39175 a_n2129_44697# a_n2065_43946# 7.26e-19
C39176 a_2437_43646# a_1756_43548# 8.79e-19
C39177 a_n443_42852# a_421_43172# 4.81e-19
C39178 a_13717_47436# CLK 0.057477f
C39179 a_n755_45592# a_8037_42858# 0.033004f
C39180 a_n357_42282# a_8605_42826# 0.011429f
C39181 a_16763_47508# VDD 0.392885f
C39182 a_n2661_43370# a_8333_44056# 5.2e-21
C39183 a_n2017_45002# a_n1177_43370# 4.91e-19
C39184 a_n2661_45010# a_104_43370# 1.69e-20
C39185 a_n2293_45010# a_n447_43370# 1.3e-19
C39186 a_n310_44484# a_n2661_42834# 9.37e-20
C39187 a_9313_44734# a_n2661_43922# 0.028486f
C39188 a_22223_46124# a_8049_45260# 0.007569f
C39189 a_1823_45246# a_1848_45724# 0.028459f
C39190 a_n2293_46098# a_2277_45546# 0.005746f
C39191 a_5164_46348# a_n2661_45546# 8.06e-20
C39192 a_n1925_46634# a_2382_45260# 8.42e-21
C39193 a_n1613_43370# a_626_44172# 0.001807f
C39194 a_1431_46436# a_1337_46116# 1.26e-19
C39195 a_14493_46090# a_14537_46482# 3.69e-19
C39196 a_13925_46122# a_14949_46494# 2.36e-20
C39197 a_12891_46348# a_14180_45002# 2.92e-20
C39198 a_167_45260# a_n755_45592# 1.02724f
C39199 a_n746_45260# a_n1352_44484# 0.001882f
C39200 a_n971_45724# a_n452_44636# 1.31e-21
C39201 a_n2438_43548# a_327_44734# 0.013318f
C39202 a_n743_46660# a_1667_45002# 2.23e-20
C39203 a_n133_46660# a_413_45260# 3.34e-21
C39204 a_n2293_46634# a_3429_45260# 0.001376f
C39205 a_8270_45546# a_8696_44636# 0.023406f
C39206 a_4915_47217# a_11691_44458# 0.020788f
C39207 a_12861_44030# a_16922_45042# 0.120012f
C39208 a_12594_46348# a_13259_45724# 0.012487f
C39209 a_12549_44172# a_13777_45326# 1.49e-20
C39210 a_768_44030# a_13556_45296# 0.267809f
C39211 a_n1853_46287# a_n443_42852# 0.003661f
C39212 a_171_46873# a_n37_45144# 2.73e-19
C39213 a_11415_45002# a_2711_45572# 0.337384f
C39214 a_14035_46660# a_13904_45546# 8.04e-20
C39215 a_765_45546# a_7499_43078# 2.08e-20
C39216 a_6123_31319# a_5742_30871# 0.106954f
C39217 a_4190_30871# C7_N_btm 2.94e-19
C39218 a_16823_43084# VDD 0.159922f
C39219 a_8791_42308# a_9223_42460# 0.014257f
C39220 a_8325_42308# a_9293_42558# 7.62e-20
C39221 a_13467_32519# C1_N_btm 0.031032f
C39222 a_n913_45002# a_22165_42308# 0.074472f
C39223 a_20512_43084# a_11341_43940# 0.02996f
C39224 a_n356_44636# a_n1557_42282# 0.017569f
C39225 a_5663_43940# a_6101_44260# 0.013015f
C39226 a_5495_43940# a_n2661_42282# 0.003301f
C39227 a_17613_45144# a_15743_43084# 1.82e-22
C39228 a_18587_45118# a_18429_43548# 1.57e-21
C39229 a_14035_46660# CLK 3.17e-20
C39230 en_comp a_20922_43172# 3.26e-22
C39231 a_13249_42308# a_1606_42308# 1.12e-20
C39232 a_n2956_38680# a_n3565_38216# 0.003389f
C39233 a_375_42282# a_421_43172# 0.00164f
C39234 a_4099_45572# a_3775_45552# 0.003943f
C39235 a_6472_45840# a_6511_45714# 0.781352f
C39236 a_6194_45824# a_6667_45809# 7.99e-20
C39237 a_5164_46348# a_5205_44484# 7.43e-20
C39238 a_8049_45260# a_16842_45938# 1.72e-19
C39239 a_12549_44172# a_20640_44752# 0.004896f
C39240 a_2324_44458# a_n913_45002# 1.92e-20
C39241 a_19321_45002# a_17517_44484# 0.264473f
C39242 a_3483_46348# a_8953_45002# 0.121322f
C39243 a_8016_46348# a_5111_44636# 0.001121f
C39244 a_22223_46124# a_19479_31679# 4.31e-19
C39245 a_6945_45028# a_3357_43084# 0.033591f
C39246 a_19692_46634# a_11827_44484# 0.04136f
C39247 a_13259_45724# a_15037_45618# 0.098143f
C39248 a_6165_46155# a_3232_43370# 9.41e-20
C39249 a_8953_45546# a_3537_45260# 0.009809f
C39250 a_5937_45572# a_4574_45260# 7.5e-21
C39251 a_5932_42308# C3_N_btm 0.121156f
C39252 a_n1151_42308# a_13507_46334# 0.001912f
C39253 a_1606_42308# VIN_P 0.014401f
C39254 a_5742_30871# EN_VIN_BSTR_P 0.645417f
C39255 a_n1435_47204# a_12861_44030# 0.036547f
C39256 a_13381_47204# a_13487_47204# 0.152045f
C39257 a_n4209_38502# a_n3690_38528# 0.045251f
C39258 a_n3420_39072# a_n4334_38304# 2.34e-19
C39259 a_n4334_38528# a_n3565_38502# 2e-19
C39260 a_5934_30871# C1_P_btm 0.011025f
C39261 a_n971_45724# a_2747_46873# 0.047519f
C39262 a_n452_47436# a_n310_47243# 0.005572f
C39263 a_3497_42558# VDD 0.007751f
C39264 a_6123_31319# C0_dummy_P_btm 1.31e-19
C39265 a_16104_42674# CAL_N 1.8e-20
C39266 a_2905_45572# a_4883_46098# 3.03e-20
C39267 a_n2956_37592# a_n4064_40160# 0.012264f
C39268 a_n310_45899# VDD 0.002211f
C39269 a_15682_43940# a_10341_43396# 3.89e-19
C39270 a_n2472_43914# a_n2472_42826# 0.001034f
C39271 a_n2810_45028# a_n2302_40160# 0.001344f
C39272 a_n2293_42834# a_6123_31319# 4.85e-19
C39273 a_1307_43914# a_15051_42282# 1.26e-20
C39274 a_n2433_43396# a_n2267_43396# 0.756435f
C39275 a_n4318_39304# a_n1699_43638# 8.9e-20
C39276 a_2711_45572# a_6945_45348# 9.26e-20
C39277 a_10903_43370# a_13213_44734# 4.28e-19
C39278 a_13661_43548# a_2982_43646# 2.6e-20
C39279 a_768_44030# a_6293_42852# 5.95e-20
C39280 SMPL_ON_P a_n3674_39304# 0.040131f
C39281 a_4791_45118# a_743_42282# 0.053017f
C39282 a_n443_42852# a_n2661_43370# 0.082119f
C39283 a_16327_47482# a_16547_43609# 0.00506f
C39284 a_11415_45002# a_22485_44484# 3.2e-20
C39285 a_10227_46804# a_13749_43396# 3.64e-19
C39286 a_11823_42460# a_13159_45002# 7.87e-19
C39287 a_12791_45546# a_13017_45260# 3.34e-19
C39288 a_20205_31679# a_22223_45036# 2.02e-20
C39289 a_12861_44030# a_15743_43084# 0.01437f
C39290 a_18909_45814# a_19365_45572# 4.2e-19
C39291 a_3090_45724# a_10807_43548# 0.031941f
C39292 VDAC_N VIN_N 0.253278f
C39293 a_22821_38993# RST_Z 1.55e-20
C39294 C10_P_btm C7_P_btm 0.680974f
C39295 a_4883_46098# a_12816_46660# 3.12e-20
C39296 a_10227_46804# a_19333_46634# 8.89e-20
C39297 a_18143_47464# a_15227_44166# 1.06e-19
C39298 a_601_46902# a_1799_45572# 1.3e-20
C39299 a_33_46660# a_n2661_46098# 0.007289f
C39300 a_948_46660# a_1110_47026# 0.006453f
C39301 a_383_46660# a_645_46660# 0.001705f
C39302 a_n2661_46634# a_3686_47026# 1.44e-19
C39303 a_9804_47204# a_10150_46912# 3.14e-19
C39304 a_n881_46662# a_10249_46116# 3.58e-19
C39305 a_12861_44030# a_13885_46660# 0.042236f
C39306 a_13717_47436# a_14035_46660# 2.07e-20
C39307 a_n1613_43370# a_6755_46942# 0.006199f
C39308 a_11453_44696# a_11735_46660# 5.11e-21
C39309 a_13507_46334# a_14084_46812# 4.22e-20
C39310 C9_P_btm C8_P_btm 29.256199f
C39311 a_n743_46660# a_2959_46660# 1.5e-20
C39312 a_n133_46660# a_2609_46660# 1.38e-21
C39313 a_n2438_43548# a_3177_46902# 2.59e-20
C39314 a_5807_45002# a_5072_46660# 7.94e-20
C39315 EN_VIN_BSTR_P C0_dummy_P_btm 0.026355f
C39316 a_5129_47502# a_765_45546# 0.004549f
C39317 a_22469_39537# VDD 0.356405f
C39318 a_n1925_46634# a_3524_46660# 0.008296f
C39319 a_15743_43084# a_19700_43370# 0.004331f
C39320 a_16137_43396# a_16823_43084# 0.038492f
C39321 a_16409_43396# a_17486_43762# 1.46e-19
C39322 a_10951_45334# CLK 0.005907f
C39323 a_n2661_42282# a_n784_42308# 0.062364f
C39324 a_12281_43396# a_4361_42308# 0.021275f
C39325 a_6031_43396# a_7227_42852# 1.51e-19
C39326 a_6293_42852# a_5755_42852# 0.114235f
C39327 a_3626_43646# a_10083_42826# 9.29e-20
C39328 a_2982_43646# a_10835_43094# 2.09e-20
C39329 a_15415_45028# VDD 0.191729f
C39330 a_n97_42460# a_18817_42826# 0.003814f
C39331 a_10341_43396# a_22223_43396# 0.038582f
C39332 a_9482_43914# a_13807_45067# 0.00608f
C39333 a_4185_45028# a_2982_43646# 0.243496f
C39334 a_10193_42453# a_19279_43940# 4.41e-19
C39335 a_4791_45118# a_5755_42308# 0.003736f
C39336 a_11823_42460# a_11967_42832# 0.573139f
C39337 a_n2293_45010# a_n452_44636# 3.23e-20
C39338 a_n2661_45010# a_949_44458# 0.071688f
C39339 SMPL_ON_N a_22400_42852# 3.97e-19
C39340 a_375_42282# a_n2661_43370# 0.012518f
C39341 a_14537_43396# a_14976_45348# 9.13e-19
C39342 a_n443_42852# a_2998_44172# 1.29e-19
C39343 en_comp a_n2661_44458# 0.030481f
C39344 a_n2661_45546# a_3499_42826# 5.13e-21
C39345 a_13259_45724# a_17737_43940# 0.016944f
C39346 a_526_44458# a_5025_43940# 1.8e-20
C39347 a_13507_46334# a_19240_46482# 0.002125f
C39348 a_5385_46902# a_5164_46348# 0.001231f
C39349 a_4817_46660# a_5204_45822# 0.001084f
C39350 a_2063_45854# a_3175_45822# 0.002195f
C39351 a_13885_46660# a_14180_46812# 0.150851f
C39352 a_17609_46634# a_18285_46348# 0.115413f
C39353 a_18597_46090# a_20254_46482# 0.002021f
C39354 a_8128_46384# a_8283_46482# 0.007532f
C39355 a_15227_44166# a_765_45546# 3.46e-20
C39356 a_n1613_43370# a_8049_45260# 2.61e-20
C39357 a_4646_46812# a_6419_46155# 6.54e-20
C39358 a_n443_46116# a_1609_45822# 0.096281f
C39359 a_4915_47217# a_n443_42852# 1.15e-20
C39360 a_n237_47217# a_7227_45028# 1.15e-19
C39361 a_n971_45724# a_3638_45822# 2.91e-19
C39362 a_n2956_39768# a_n2956_39304# 0.098523f
C39363 a_2107_46812# a_2324_44458# 0.051531f
C39364 a_18479_47436# a_20850_46482# 7.88e-19
C39365 a_4883_46098# a_18243_46436# 1.03e-19
C39366 a_12465_44636# a_13259_45724# 0.096616f
C39367 a_3422_30871# C2_N_btm 9.13e-20
C39368 a_21356_42826# a_21671_42860# 0.084365f
C39369 a_14209_32519# a_14097_32519# 10.7606f
C39370 a_4190_30871# COMP_P 0.027242f
C39371 a_3626_43646# a_15761_42308# 1.94e-19
C39372 a_19279_43940# VDD 0.302681f
C39373 a_8952_43230# a_9061_43230# 0.007416f
C39374 a_9127_43156# a_9306_43218# 0.007399f
C39375 a_8387_43230# a_8495_42852# 0.057222f
C39376 a_1307_43914# a_3905_42865# 0.224019f
C39377 a_11827_44484# a_13296_44484# 6.45e-19
C39378 a_n357_42282# a_18783_43370# 5.79e-20
C39379 a_n443_42852# a_15681_43442# 0.035093f
C39380 a_6298_44484# a_6109_44484# 0.068396f
C39381 a_5343_44458# a_8375_44464# 0.007376f
C39382 a_n2661_44458# a_10617_44484# 0.003557f
C39383 a_18184_42460# a_17517_44484# 0.020871f
C39384 a_7499_43078# a_6452_43396# 1.51e-20
C39385 a_3232_43370# a_6101_44260# 0.001648f
C39386 a_3537_45260# a_9028_43914# 1.3e-19
C39387 a_13259_45724# a_13887_32519# 0.002751f
C39388 a_n2956_39768# a_n3565_39304# 0.003389f
C39389 a_18248_44752# a_18287_44626# 0.633819f
C39390 a_17970_44736# a_18443_44721# 7.99e-20
C39391 a_n913_45002# a_19862_44208# 3.9e-20
C39392 a_1423_45028# a_2479_44172# 3.74e-20
C39393 a_526_44458# a_8952_43230# 0.039329f
C39394 a_21496_47436# a_413_45260# 8.97e-20
C39395 a_14493_46090# a_2324_44458# 6.29e-20
C39396 a_14275_46494# a_14840_46494# 7.99e-20
C39397 a_3147_46376# a_526_44458# 0.352f
C39398 a_3483_46348# a_2981_46116# 2.44e-19
C39399 a_8270_45546# a_7227_45028# 1.35e-20
C39400 a_9863_46634# a_10193_42453# 1.87e-19
C39401 a_10428_46928# a_10053_45546# 2.44e-21
C39402 a_10150_46912# a_10180_45724# 7.45e-19
C39403 a_n443_46116# a_501_45348# 1.62e-19
C39404 a_19594_46812# a_19431_45546# 2.2e-19
C39405 a_19321_45002# a_19256_45572# 0.004884f
C39406 a_13747_46662# a_18799_45938# 0.028671f
C39407 a_12549_44172# a_21188_45572# 4.02e-21
C39408 a_7989_47542# a_2437_43646# 9.04e-19
C39409 a_n2312_40392# a_n2810_45028# 0.055228f
C39410 SMPL_ON_P a_n2293_42834# 1.07e-19
C39411 a_6969_46634# a_6812_45938# 4.71e-20
C39412 a_5937_45572# a_10809_44734# 0.001476f
C39413 a_9625_46129# a_6945_45028# 1.2e-19
C39414 a_16327_47482# a_6171_45002# 0.001024f
C39415 a_1606_42308# a_2123_42473# 0.011716f
C39416 a_14635_42282# a_13657_42558# 4.38e-21
C39417 a_13291_42460# a_14113_42308# 0.025652f
C39418 a_7112_43396# VDD 0.273193f
C39419 a_1576_42282# a_2713_42308# 1.15e-20
C39420 a_1184_42692# a_2725_42558# 1.23e-20
C39421 a_n2472_43914# a_n2065_43946# 0.039807f
C39422 a_14537_43396# a_16547_43609# 2.37e-20
C39423 en_comp a_17364_32525# 8.05e-20
C39424 a_n2017_45002# a_n1991_42858# 0.053113f
C39425 a_n913_45002# a_n2157_42858# 0.00135f
C39426 a_n1059_45260# a_n1853_43023# 0.03561f
C39427 a_n2293_45010# a_n1641_43230# 2.03e-19
C39428 a_n2129_44697# a_n2129_43609# 9.9e-19
C39429 a_n2267_44484# a_n2433_43396# 0.00138f
C39430 a_n2840_43914# a_n1761_44111# 1.61e-20
C39431 a_10057_43914# a_10555_43940# 0.001842f
C39432 a_9863_46634# VDD 0.411318f
C39433 a_n2433_44484# a_n2267_43396# 2.4e-19
C39434 a_5257_43370# DATA[3] 9.23e-21
C39435 a_n2661_45546# a_3316_45546# 0.027868f
C39436 a_n2293_46634# a_8103_44636# 7.43e-21
C39437 a_13759_46122# a_8696_44636# 1.49e-20
C39438 a_21363_46634# a_413_45260# 3.6e-20
C39439 a_11453_44696# a_10617_44484# 3.76e-20
C39440 a_380_45546# a_310_45028# 0.057269f
C39441 a_n863_45724# a_n755_45592# 1.76733f
C39442 a_13259_45724# a_2711_45572# 1.26722f
C39443 a_13661_43548# a_14539_43914# 0.193767f
C39444 a_15682_46116# a_15599_45572# 0.009928f
C39445 a_2324_44458# a_15903_45785# 0.017867f
C39446 a_15227_44166# a_16751_45260# 1.7e-20
C39447 a_n2497_47436# a_2479_44172# 4.48e-20
C39448 a_21076_30879# a_20447_31679# 0.055814f
C39449 a_n971_45724# a_n809_44244# 0.002895f
C39450 a_8049_45260# a_7230_45938# 1.18e-19
C39451 a_8034_45724# a_9049_44484# 2.06e-20
C39452 a_12465_44636# a_n2661_43922# 0.17969f
C39453 a_11136_42852# VDD 0.132515f
C39454 a_7174_31319# a_1736_39587# 1.22e-19
C39455 a_n4064_40160# a_n4251_40480# 0.00119f
C39456 a_n4315_30879# a_n4209_39590# 4.31257f
C39457 a_1606_42308# a_11206_38545# 3.98e-20
C39458 a_n785_47204# a_1239_47204# 4.16e-19
C39459 a_n746_45260# a_584_46384# 0.491308f
C39460 a_n2109_47186# a_3785_47178# 0.190973f
C39461 a_n971_45724# a_2063_45854# 0.164981f
C39462 a_n237_47217# a_2124_47436# 0.001177f
C39463 a_n1741_47186# a_n1151_42308# 2.98024f
C39464 a_11967_42832# a_18429_43548# 0.019775f
C39465 a_18588_44850# a_18783_43370# 7.03e-21
C39466 a_20935_43940# a_20974_43370# 0.005283f
C39467 a_11341_43940# a_21381_43940# 0.034147f
C39468 a_3737_43940# a_3992_43940# 0.005172f
C39469 a_n913_45002# a_9803_42558# 0.001906f
C39470 a_n2017_45002# a_9377_42558# 0.001128f
C39471 a_15682_43940# a_n97_42460# 0.002081f
C39472 a_n2661_42282# a_3080_42308# 0.161683f
C39473 a_20512_43084# a_10341_43396# 0.758407f
C39474 a_5527_46155# VDD 2.18e-20
C39475 a_n356_44636# a_3935_42891# 2.82e-22
C39476 a_2324_44458# a_n2661_44458# 0.134417f
C39477 a_3483_46348# a_17767_44458# 8.35e-19
C39478 a_n443_46116# a_2437_43396# 7.55e-19
C39479 a_21588_30879# a_14021_43940# 1.53e-20
C39480 a_768_44030# a_7499_43940# 1.16e-19
C39481 a_5937_45572# a_5883_43914# 0.454323f
C39482 a_8953_45546# a_8701_44490# 0.005445f
C39483 a_8199_44636# a_9838_44484# 0.024921f
C39484 a_10809_44734# a_11691_44458# 0.354084f
C39485 a_8016_46348# a_10334_44484# 0.007545f
C39486 a_15765_45572# a_16115_45572# 0.20669f
C39487 a_15599_45572# a_16680_45572# 0.102355f
C39488 a_4646_46812# a_n2661_42282# 0.025072f
C39489 a_15903_45785# a_16855_45546# 9.79e-21
C39490 a_20202_43084# a_9313_44734# 0.044152f
C39491 a_1609_45822# a_3537_45260# 1.84e-20
C39492 a_n443_42852# a_4574_45260# 1.14e-21
C39493 a_n2109_47186# a_3090_45724# 2.79e-20
C39494 a_8912_37509# a_11206_38545# 1.26605f
C39495 VDAC_N CAL_N 2.77e-19
C39496 a_4791_45118# a_6755_46942# 2.99e-19
C39497 a_6151_47436# a_10428_46928# 0.001405f
C39498 a_6575_47204# a_8145_46902# 0.001541f
C39499 a_7903_47542# a_7927_46660# 1.47e-20
C39500 a_n3607_38528# VDD 2.79e-20
C39501 a_n1613_43370# a_n2442_46660# 4.46e-21
C39502 a_12549_44172# a_19321_45002# 0.238866f
C39503 VDAC_Ni a_n923_35174# 7.46e-19
C39504 a_n4209_38502# VIN_P 0.028945f
C39505 a_19479_31679# C5_N_btm 1.11e-20
C39506 a_n2433_43396# a_n2472_42826# 9.53e-19
C39507 a_1209_43370# a_743_42282# 3.61e-21
C39508 a_9145_43396# a_14358_43442# 0.053427f
C39509 a_20269_44172# a_19987_42826# 8.09e-21
C39510 a_15493_43940# a_18083_42858# 1.12e-20
C39511 a_11341_43940# a_18249_42858# 4.65e-20
C39512 a_n356_44636# a_15890_42674# 2.92e-19
C39513 a_17730_32519# a_14097_32519# 0.053763f
C39514 a_9313_44734# a_10545_42558# 6.42e-19
C39515 a_n2293_43922# a_5934_30871# 0.079987f
C39516 a_19862_44208# a_20922_43172# 0.164553f
C39517 a_10903_43370# a_11341_43940# 0.061205f
C39518 a_20202_43084# a_20974_43370# 0.026132f
C39519 a_2680_45002# a_1423_45028# 0.003069f
C39520 a_5147_45002# a_1307_43914# 0.032106f
C39521 a_17668_45572# a_17613_45144# 5.67e-19
C39522 a_18799_45938# a_18911_45144# 4.07e-20
C39523 a_768_44030# a_10991_42826# 1.43e-20
C39524 a_6171_45002# a_14537_43396# 0.054973f
C39525 a_2711_45572# a_n2661_43922# 4.93e-20
C39526 a_17715_44484# a_17973_43940# 0.00355f
C39527 a_18175_45572# a_11827_44484# 1.29e-20
C39528 a_2437_43646# a_n2661_43370# 0.033415f
C39529 a_2274_45254# a_2304_45348# 0.062682f
C39530 a_1823_45246# a_5829_43940# 1.54e-19
C39531 a_9290_44172# a_9248_44260# 5.95e-19
C39532 a_n2438_43548# a_n3674_39304# 0.001617f
C39533 a_18479_47436# a_10809_44734# 0.04504f
C39534 a_n2293_46634# a_n2472_46090# 3.35e-19
C39535 a_6575_47204# a_5066_45546# 2.37e-20
C39536 a_9863_46634# a_10185_46660# 0.007399f
C39537 a_11453_44696# a_2324_44458# 0.023884f
C39538 a_13507_46334# a_19553_46090# 0.002559f
C39539 a_n1151_42308# a_10586_45546# 0.02493f
C39540 a_8128_46384# a_7920_46348# 0.197919f
C39541 a_n881_46662# a_5937_45572# 0.195456f
C39542 a_n1613_43370# a_8953_45546# 0.024821f
C39543 a_12465_44636# a_18189_46348# 1.08e-20
C39544 a_18597_46090# a_6945_45028# 0.049383f
C39545 a_4883_46098# a_18819_46122# 0.054304f
C39546 a_3686_47026# a_765_45546# 1.39e-19
C39547 a_4791_45118# a_8049_45260# 3.69e-19
C39548 a_n2661_46634# a_n1853_46287# 2.3e-19
C39549 a_14209_32519# a_22959_42860# 0.007868f
C39550 a_8605_42826# a_8952_43230# 0.051162f
C39551 a_8037_42858# a_10083_42826# 1.62e-19
C39552 a_n310_44811# VDD 0.001779f
C39553 a_15493_43940# a_22775_42308# 6.96e-21
C39554 a_n97_42460# a_5934_30871# 0.221607f
C39555 a_4905_42826# a_5379_42460# 0.077171f
C39556 a_3080_42308# a_3497_42558# 4.3e-19
C39557 a_n2293_46634# a_14456_42282# 3e-20
C39558 a_12549_44172# a_17531_42308# 1.47e-21
C39559 a_n863_45724# a_548_43396# 0.001035f
C39560 a_17719_45144# a_17767_44458# 0.001046f
C39561 a_2437_43646# a_2998_44172# 1.59e-20
C39562 a_4185_45028# a_7871_42858# 1.73e-20
C39563 a_20202_43084# a_18599_43230# 5.72e-21
C39564 a_n357_42282# a_3626_43646# 0.020238f
C39565 a_n2661_44458# a_n1699_44726# 0.009008f
C39566 a_n2433_44484# a_n2267_44484# 0.730194f
C39567 a_16922_45042# a_18287_44626# 1.76e-19
C39568 a_n4318_40392# a_n1917_44484# 3.81e-20
C39569 a_n2661_43370# a_4181_44734# 4.39e-19
C39570 a_11827_44484# a_10440_44484# 1.55e-19
C39571 a_17478_45572# a_17737_43940# 7.33e-21
C39572 en_comp a_19237_31679# 1.18e-19
C39573 a_n2312_39304# a_n4064_40160# 5.41e-19
C39574 a_n2312_40392# a_n2302_40160# 0.151095f
C39575 a_n913_45002# a_n1761_44111# 0.036392f
C39576 a_n1059_45260# a_n1899_43946# 5.95e-19
C39577 a_n2661_45010# a_175_44278# 6.99e-20
C39578 a_n2293_45010# a_n809_44244# 0.041966f
C39579 a_14537_43396# a_14673_44172# 0.044194f
C39580 a_n443_42852# a_1568_43370# 0.038016f
C39581 a_7499_43078# a_11173_43940# 5.28e-20
C39582 a_n2661_45546# a_6197_43396# 1.24e-21
C39583 a_16327_47482# a_18909_45814# 0.16767f
C39584 a_11415_45002# a_12005_46116# 1.53e-20
C39585 a_n2497_47436# a_2680_45002# 1.29e-19
C39586 a_1823_45246# a_4185_45028# 0.081652f
C39587 a_4700_47436# a_3357_43084# 6.56e-19
C39588 a_11453_44696# a_16855_45546# 3.46e-20
C39589 a_20411_46873# a_19900_46494# 6.79e-19
C39590 a_20107_46660# a_20708_46348# 2.61e-20
C39591 a_20273_46660# a_20075_46420# 5.46e-21
C39592 a_19123_46287# a_6945_45028# 1.85e-19
C39593 a_17829_46910# a_10809_44734# 0.02024f
C39594 a_11813_46116# a_12638_46436# 3.97e-19
C39595 a_4915_47217# a_2437_43646# 0.114772f
C39596 a_n971_45724# a_n955_45028# 5.28e-19
C39597 a_167_45260# a_3483_46348# 1.26e-19
C39598 a_2698_46116# a_2804_46116# 0.313533f
C39599 a_5807_45002# a_11823_42460# 0.022934f
C39600 a_1799_45572# a_2711_45572# 7.16e-20
C39601 a_2107_46812# a_6667_45809# 4.38e-20
C39602 a_11599_46634# a_18799_45938# 0.001679f
C39603 a_5342_30871# a_14456_42282# 0.160195f
C39604 a_9801_43940# VDD 0.19512f
C39605 a_3626_43646# CAL_N 0.00204f
C39606 a_5534_30871# a_13333_42558# 0.002157f
C39607 a_10903_43370# a_10723_42308# 1.71e-19
C39608 a_21359_45002# a_14021_43940# 5.71e-21
C39609 a_20916_46384# VDD 0.302226f
C39610 a_375_42282# a_1568_43370# 3.7e-21
C39611 a_5807_45002# DATA[3] 4.68e-21
C39612 a_20843_47204# START 1.11e-19
C39613 a_8701_44490# a_9028_43914# 0.008509f
C39614 a_5883_43914# a_8333_44056# 0.152643f
C39615 a_10193_42453# a_12545_42858# 8.12e-20
C39616 a_n357_42282# a_8649_43218# 3.99e-19
C39617 a_526_44458# a_2123_42473# 0.012631f
C39618 a_n1925_42282# a_1755_42282# 0.019802f
C39619 a_9290_44172# a_11633_42558# 0.014294f
C39620 a_13259_45724# a_16877_42852# 3.34e-20
C39621 a_20202_43084# a_22397_42558# 1.54e-19
C39622 a_1307_43914# a_4093_43548# 0.002897f
C39623 a_7229_43940# a_6031_43396# 1.49e-19
C39624 a_17517_44484# a_20362_44736# 0.047565f
C39625 a_3065_45002# a_3457_43396# 0.005043f
C39626 a_5111_44636# a_8791_43396# 0.05316f
C39627 a_22612_30879# C10_N_btm 1.5848f
C39628 a_n2017_45002# a_14205_43396# 6.74e-21
C39629 a_n1059_45260# a_14358_43442# 1.98e-20
C39630 a_n913_45002# a_14579_43548# 0.239851f
C39631 a_5205_44484# a_6197_43396# 1.83e-19
C39632 a_10227_46804# a_10157_44484# 0.008568f
C39633 a_2324_44458# a_5907_45546# 0.002504f
C39634 a_526_44458# a_310_45028# 1.77e-21
C39635 a_10809_44734# a_n443_42852# 3.02e-20
C39636 a_n2438_43548# a_n2293_42834# 0.138621f
C39637 a_13661_43548# a_14309_45028# 1.43e-19
C39638 a_n971_45724# a_n2661_42834# 0.165951f
C39639 a_4791_45118# a_5289_44734# 7.66e-19
C39640 a_n881_46662# a_11691_44458# 4.5e-20
C39641 a_15559_46634# a_3357_43084# 2.61e-21
C39642 a_18189_46348# a_2711_45572# 3.03e-20
C39643 a_5066_45546# a_n2661_45546# 9.86e-19
C39644 a_n2661_46634# a_n2661_43370# 7.12e-19
C39645 a_8667_46634# a_6171_45002# 7.94e-23
C39646 a_2063_45854# a_9313_44734# 3.29e-20
C39647 a_12861_44030# a_17970_44736# 0.001384f
C39648 a_12549_44172# a_18184_42460# 0.03123f
C39649 a_8199_44636# a_8568_45546# 0.141772f
C39650 a_8016_46348# a_9049_44484# 4.89e-19
C39651 a_7715_46873# a_7229_43940# 2.31e-19
C39652 a_5342_30871# C4_N_btm 8.98e-20
C39653 a_n4318_38216# a_n3607_38304# 7.49e-20
C39654 a_5932_42308# a_1736_39587# 1.46e-19
C39655 a_13070_42354# a_7174_31319# 4.88e-21
C39656 a_5534_30871# C6_N_btm 0.01116f
C39657 a_12545_42858# VDD 0.285703f
C39658 a_18287_44626# a_15743_43084# 3.79e-20
C39659 a_18374_44850# a_18525_43370# 8.44e-21
C39660 a_18443_44721# a_18783_43370# 1.12e-19
C39661 a_n356_44636# a_16547_43609# 3.88e-21
C39662 a_14539_43914# a_15037_43396# 8.32e-22
C39663 a_4185_45028# DATA[2] 0.002615f
C39664 a_9313_44734# a_14955_43396# 0.001014f
C39665 a_10193_42453# a_19332_42282# 0.004163f
C39666 a_n2956_38216# a_n2302_38778# 4.36e-19
C39667 a_11967_42832# a_2982_43646# 5.64e-19
C39668 a_20512_43084# a_n97_42460# 2.54e-19
C39669 a_n1761_44111# a_n4318_39304# 3.05e-19
C39670 a_n2065_43946# a_n2433_43396# 6.16e-19
C39671 a_7542_44172# a_8415_44056# 2.49e-20
C39672 a_6165_46155# VDD 0.204296f
C39673 a_19328_44172# a_19478_44306# 0.188181f
C39674 a_10405_44172# a_10555_44260# 0.085098f
C39675 a_14955_43940# a_11341_43940# 0.005859f
C39676 a_11823_42460# a_15143_45578# 0.120787f
C39677 a_13527_45546# a_13904_45546# 3.21e-19
C39678 a_10193_42453# a_10210_45822# 0.026406f
C39679 a_10180_45724# a_10907_45822# 6.72e-20
C39680 a_8199_44636# a_n2661_43370# 0.126664f
C39681 a_3090_45724# a_8375_44464# 9.88e-21
C39682 a_20202_43084# a_18114_32519# 1.27e-19
C39683 a_n1613_43370# a_9028_43914# 2.5e-20
C39684 a_5066_45546# a_5205_44484# 1.52e-20
C39685 a_8568_45546# a_8192_45572# 1.96e-19
C39686 a_8162_45546# a_8697_45572# 0.001108f
C39687 a_7499_43078# a_8120_45572# 1.34e-20
C39688 a_n2438_43548# a_1115_44172# 5.77e-19
C39689 a_8270_45546# a_9159_44484# 4.45e-19
C39690 a_13507_46334# a_15493_43940# 0.021188f
C39691 a_12741_44636# a_18450_45144# 4.86e-19
C39692 a_13059_46348# a_13720_44458# 0.008849f
C39693 a_n2497_47436# a_n229_43646# 0.022782f
C39694 a_n971_45724# a_n1352_43396# 0.005968f
C39695 a_2324_44458# a_6125_45348# 0.001467f
C39696 a_18907_42674# RST_Z 1.72e-20
C39697 a_n2109_47186# a_3699_46634# 6.42e-20
C39698 a_4915_47217# a_n2661_46634# 9.46e-19
C39699 a_9313_45822# a_5807_45002# 0.031627f
C39700 a_13487_47204# a_13675_47204# 0.001217f
C39701 a_12861_44030# a_13759_47204# 0.001988f
C39702 a_7174_31319# C2_N_btm 1.86e-20
C39703 a_n4064_40160# C8_P_btm 4.06e-19
C39704 a_15507_47210# a_768_44030# 5.43e-20
C39705 a_n4064_39616# EN_VIN_BSTR_P 0.072552f
C39706 a_n815_47178# a_n2661_46098# 3.57e-20
C39707 a_n746_45260# a_479_46660# 0.001012f
C39708 a_n1151_42308# a_n743_46660# 0.195953f
C39709 a_3160_47472# a_n2438_43548# 3.61e-21
C39710 a_7754_39964# a_7754_38968# 1.48e-20
C39711 a_13258_32519# C5_N_btm 1.87e-19
C39712 a_584_46384# a_383_46660# 0.001651f
C39713 a_15811_47375# a_12549_44172# 0.024519f
C39714 a_19332_42282# VDD 0.227361f
C39715 a_n4209_38216# a_n4064_37440# 0.028219f
C39716 a_n3565_38216# a_n3420_37440# 0.038559f
C39717 a_n4064_37984# a_n4209_37414# 0.027993f
C39718 a_2113_38308# a_3754_38470# 2.91e-19
C39719 a_n3420_37984# a_n3565_37414# 0.032929f
C39720 a_n3690_38304# a_n3690_37440# 0.050585f
C39721 a_3785_47178# a_n1925_46634# 3.96e-20
C39722 a_n356_44636# a_n3674_37592# 4.6e-21
C39723 a_21381_43940# a_10341_43396# 0.03047f
C39724 a_n97_42460# a_7221_43396# 1.23e-19
C39725 a_10210_45822# VDD 0.323342f
C39726 a_11341_43940# a_5649_42852# 0.01232f
C39727 a_15493_43940# a_21855_43396# 2.4e-19
C39728 a_14021_43940# a_16823_43084# 0.005626f
C39729 a_4223_44672# a_7227_42308# 3.26e-37
C39730 a_n971_45724# a_n2293_42282# 6.84e-19
C39731 a_3090_45724# a_19319_43548# 1.22e-19
C39732 a_6667_45809# a_n2661_44458# 6.66e-21
C39733 a_n2293_46634# a_10149_43396# 4e-19
C39734 a_4646_46812# a_7112_43396# 0.07278f
C39735 a_12741_44636# a_12429_44172# 3.86e-19
C39736 a_n2017_45002# a_n967_45348# 0.095287f
C39737 a_3357_43084# a_3065_45002# 0.316449f
C39738 a_n1059_45260# en_comp 8.56e-20
C39739 a_13661_43548# a_17324_43396# 9.28e-20
C39740 a_4915_47217# a_14543_43071# 1.12e-21
C39741 a_11415_45002# a_15682_43940# 6.37e-20
C39742 a_n2293_45010# a_n955_45028# 8.22e-21
C39743 a_n2661_45010# a_n143_45144# 5.24e-21
C39744 a_1138_42852# a_1525_44260# 2.28e-20
C39745 a_16147_45260# a_16019_45002# 0.186254f
C39746 a_5257_43370# a_2982_43646# 2.26e-20
C39747 a_n443_42852# a_5883_43914# 8.2e-19
C39748 a_5907_46634# a_7715_46873# 8.55e-21
C39749 a_n1925_46634# a_3090_45724# 8.91e-20
C39750 a_5807_45002# a_12513_46660# 7.17e-19
C39751 a_12549_44172# a_13059_46348# 0.808395f
C39752 a_13507_46334# a_12741_44636# 0.137731f
C39753 a_6540_46812# a_5257_43370# 0.00507f
C39754 a_5732_46660# a_7411_46660# 1.96e-20
C39755 a_n1151_42308# a_11189_46129# 0.12414f
C39756 a_11453_44696# a_21350_47026# 3.86e-19
C39757 a_22223_47212# a_22365_46825# 0.011422f
C39758 a_12465_44636# a_20202_43084# 8.04e-20
C39759 a_4915_47217# a_8199_44636# 2.73e-20
C39760 a_n443_46116# a_5937_45572# 4.89e-20
C39761 a_4791_45118# a_8953_45546# 1.45e-19
C39762 a_6545_47178# a_6419_46155# 0.080336f
C39763 a_n97_42460# a_16245_42852# 0.088473f
C39764 a_17538_32519# a_14097_32519# 0.050981f
C39765 a_10807_43548# a_11633_42558# 8.38e-19
C39766 a_10341_43396# a_18249_42858# 9.84e-20
C39767 a_21101_45002# VDD 0.2903f
C39768 a_n2293_43922# a_7754_40130# 6.5e-19
C39769 a_11750_44172# a_11551_42558# 8.92e-22
C39770 a_n2312_38680# a_n4318_38216# 0.023247f
C39771 a_n2442_46660# a_n1736_42282# 4.03e-20
C39772 a_9290_44172# a_12281_43396# 0.36475f
C39773 a_13259_45724# a_14401_32519# 4.2e-20
C39774 a_14537_43396# a_12607_44458# 1.38e-21
C39775 a_3537_45260# a_5205_44734# 6.62e-22
C39776 a_n2472_45002# a_n2661_43922# 6.45e-19
C39777 a_n2661_45010# a_n2293_43922# 2.75e-20
C39778 a_n2293_45010# a_n2661_42834# 0.083461f
C39779 a_10227_46804# a_14113_42308# 0.627404f
C39780 a_21076_30879# a_13467_32519# 0.055522f
C39781 a_768_44030# a_2713_42308# 5.49e-20
C39782 a_2324_44458# a_9145_43396# 9.23e-23
C39783 a_10903_43370# a_10341_43396# 0.042836f
C39784 SMPL_ON_P a_n4064_39616# 1.56e-20
C39785 a_13556_45296# a_13720_44458# 0.212774f
C39786 a_1423_45028# a_5518_44484# 0.047243f
C39787 a_1307_43914# a_10157_44484# 6.43e-20
C39788 a_9482_43914# a_15004_44636# 0.34299f
C39789 a_16922_45042# a_17023_45118# 0.099834f
C39790 a_7499_43078# a_7911_44260# 7.28e-19
C39791 a_18479_45785# a_19279_43940# 0.019159f
C39792 a_4185_45028# a_17324_43396# 1.18e-21
C39793 a_20820_30879# a_13678_32519# 0.053259f
C39794 a_11415_45002# a_22223_43396# 2.17e-20
C39795 a_5257_43370# a_5837_42852# 4.04e-20
C39796 a_n2956_39768# a_n1329_42308# 3.21e-20
C39797 a_2711_45572# a_20935_43940# 1.09e-19
C39798 a_22612_30879# a_20205_31679# 0.111294f
C39799 a_21588_30879# a_20692_30879# 0.056225f
C39800 a_12251_46660# a_12005_46116# 8.94e-19
C39801 a_12991_46634# a_10903_43370# 1.94e-19
C39802 a_2747_46873# a_2711_45572# 3.81e-20
C39803 a_11599_46634# a_11962_45724# 1.79e-20
C39804 a_10227_46804# a_7499_43078# 0.033512f
C39805 a_n1151_42308# a_11136_45572# 3.27e-20
C39806 a_20623_46660# a_12741_44636# 0.034292f
C39807 a_21363_46634# a_20820_30879# 2.73e-19
C39808 a_14311_47204# a_11823_42460# 2.5e-21
C39809 a_768_44030# a_2957_45546# 0.027276f
C39810 a_6755_46942# a_6945_45028# 0.024014f
C39811 a_12469_46902# a_12594_46348# 4.31e-19
C39812 a_21188_46660# a_22591_46660# 1.52e-20
C39813 a_22000_46634# a_11415_45002# 1.58e-19
C39814 a_n881_46662# a_n443_42852# 0.005862f
C39815 a_13717_47436# a_13527_45546# 3.58e-22
C39816 a_12861_44030# a_13163_45724# 0.098707f
C39817 a_4361_42308# a_11551_42558# 0.011423f
C39818 a_743_42282# a_14456_42282# 0.006738f
C39819 a_16137_43396# a_19332_42282# 2.66e-19
C39820 a_1847_42826# a_3581_42558# 2.17e-20
C39821 a_19987_42826# a_20836_43172# 1.48e-20
C39822 a_16823_43084# a_15764_42576# 0.0016f
C39823 a_12545_42858# a_n784_42308# 5.9e-21
C39824 a_5649_42852# a_10723_42308# 1.31e-19
C39825 a_3935_42891# a_3823_42558# 0.012124f
C39826 a_17499_43370# a_4958_30871# 0.001145f
C39827 a_15743_43084# a_17124_42282# 1.95e-21
C39828 a_16023_47582# VDD 0.201413f
C39829 a_15415_45028# a_14021_43940# 6.12e-21
C39830 a_16327_47482# RST_Z 1.85e-19
C39831 a_14539_43914# a_11967_42832# 0.512158f
C39832 a_n2433_44484# a_n2065_43946# 0.008496f
C39833 a_n2661_44458# a_n1761_44111# 1.08e-19
C39834 a_13259_45724# a_18817_42826# 2.9e-20
C39835 a_13717_47436# EN_OFFSET_CAL 0.002392f
C39836 en_comp a_n2840_43370# 7.28e-20
C39837 a_n2956_37592# a_n4318_39304# 0.023222f
C39838 a_2437_43646# a_1568_43370# 0.058471f
C39839 a_n1435_47204# CLK 1.41989f
C39840 a_n755_45592# a_7765_42852# 0.00466f
C39841 a_n357_42282# a_8037_42858# 0.048934f
C39842 a_n2017_45002# a_n1917_43396# 0.01343f
C39843 a_n2661_45010# a_n97_42460# 8.74e-21
C39844 a_n2293_45010# a_n1352_43396# 0.002774f
C39845 a_n745_45366# a_n2129_43609# 6.64e-20
C39846 a_9241_44734# a_n2661_43922# 1.54e-35
C39847 a_9313_44734# a_n2661_42834# 0.02321f
C39848 a_6945_45028# a_8049_45260# 0.009745f
C39849 a_n2293_46098# a_1609_45822# 0.002761f
C39850 a_n2661_46634# a_4574_45260# 1.32e-20
C39851 a_n881_46662# a_375_42282# 5.71e-20
C39852 a_1337_46436# a_1337_46116# 6.96e-20
C39853 a_13759_46122# a_14949_46494# 2.56e-19
C39854 a_167_45260# a_n357_42282# 0.148401f
C39855 a_376_46348# a_n356_45724# 7.46e-20
C39856 a_n971_45724# a_n1352_44484# 0.005662f
C39857 a_n746_45260# a_n1177_44458# 0.064145f
C39858 a_5807_45002# a_7705_45326# 8.49e-21
C39859 a_n743_46660# a_327_44734# 4e-19
C39860 a_n133_46660# a_n37_45144# 4.9e-21
C39861 a_n2438_43548# a_413_45260# 0.032468f
C39862 a_n2293_46634# a_3065_45002# 0.102991f
C39863 a_n2661_46098# a_n2661_45010# 1.31e-20
C39864 a_12549_44172# a_13556_45296# 0.030045f
C39865 a_12891_46348# a_13777_45326# 0.03955f
C39866 a_768_44030# a_9482_43914# 0.77718f
C39867 a_2202_46116# a_n755_45592# 2.03e-20
C39868 a_20202_43084# a_2711_45572# 1.42e-19
C39869 a_2162_46660# a_2437_43646# 0.002257f
C39870 a_13885_46660# a_13904_45546# 8.51e-20
C39871 a_5934_30871# a_10533_42308# 7.8e-20
C39872 a_7227_42308# a_5742_30871# 2.87e-20
C39873 a_5342_30871# a_8530_39574# 1.55e-19
C39874 a_4190_30871# C6_N_btm 0.005085f
C39875 a_14097_32519# a_22465_38105# 0.002065f
C39876 a_8325_42308# a_9803_42558# 5.62e-20
C39877 a_8685_42308# a_9223_42460# 0.166964f
C39878 a_n913_45002# a_21671_42860# 8.31e-20
C39879 a_20512_43084# a_21115_43940# 1.49e-21
C39880 a_n356_44636# a_766_43646# 9.89e-19
C39881 a_5663_43940# a_5841_44260# 0.007617f
C39882 a_5013_44260# a_n2661_42282# 1.85e-20
C39883 a_13885_46660# CLK 2.64e-20
C39884 en_comp a_19987_42826# 9.77e-21
C39885 a_375_42282# a_133_43172# 7.97e-20
C39886 a_16922_45042# a_19268_43646# 1.77e-21
C39887 a_16751_46987# VDD 8.63e-19
C39888 a_19279_43940# a_14021_43940# 2.21e-19
C39889 a_6194_45824# a_6511_45714# 0.102325f
C39890 a_12549_44172# a_20362_44736# 0.015111f
C39891 a_765_45546# a_n2661_43370# 6.55e-22
C39892 a_2324_44458# a_n1059_45260# 4.3e-20
C39893 a_3090_45724# a_17801_45144# 7.84e-20
C39894 a_11133_46155# a_413_45260# 1.62e-21
C39895 a_3483_46348# a_8191_45002# 0.081038f
C39896 a_21137_46414# a_3357_43084# 1.6e-20
C39897 a_19466_46812# a_11827_44484# 1.45e-20
C39898 a_19692_46634# a_21359_45002# 7.78e-21
C39899 a_13259_45724# a_14033_45822# 0.004141f
C39900 a_10586_45546# a_12649_45572# 6.62e-20
C39901 a_10809_44734# a_2437_43646# 0.13907f
C39902 a_22223_46124# a_22223_45572# 0.025171f
C39903 a_5937_45572# a_3537_45260# 9.77e-19
C39904 a_n4209_39304# a_n3420_37984# 0.029539f
C39905 a_5932_42308# C2_N_btm 0.011289f
C39906 a_5742_30871# a_n923_35174# 0.099784f
C39907 a_n1435_47204# a_13717_47436# 0.196889f
C39908 a_13381_47204# a_12861_44030# 4.15e-20
C39909 a_n4209_38502# a_n3565_38502# 6.84323f
C39910 a_n3565_39304# a_n3565_38216# 0.02823f
C39911 a_n3420_39072# a_n4209_38216# 0.030577f
C39912 a_n785_47204# a_n2312_39304# 9.48e-20
C39913 a_5934_30871# C2_P_btm 0.011047f
C39914 a_n2109_47186# a_2583_47243# 8.31e-19
C39915 a_n971_45724# a_2487_47570# 6.45e-19
C39916 a_n1741_47186# a_3315_47570# 2.13e-19
C39917 a_6123_31319# C0_P_btm 0.018968f
C39918 a_n237_47217# a_n89_47570# 0.005668f
C39919 a_5379_42460# VDD 0.213136f
C39920 a_19721_31679# a_14097_32519# 0.051111f
C39921 a_n23_45546# VDD 0.150941f
C39922 a_14955_43940# a_10341_43396# 6.65e-21
C39923 a_10807_43548# a_12281_43396# 7.83e-20
C39924 a_1848_45724# DATA[1] 9.34e-21
C39925 a_n2956_37592# a_n4334_40480# 0.0011f
C39926 en_comp a_n4315_30879# 0.001378f
C39927 a_n2810_45028# a_n4064_40160# 0.001122f
C39928 a_n2293_42834# a_7227_42308# 7.22e-20
C39929 a_2382_45260# a_7174_31319# 4.88e-21
C39930 a_n2433_43396# a_n2129_43609# 0.283605f
C39931 a_n4318_39304# a_n2267_43396# 4.55e-19
C39932 a_11341_43940# a_8685_43396# 2.48e-19
C39933 a_895_43940# a_743_42282# 2.08e-20
C39934 a_8049_45260# a_8103_44636# 0.012205f
C39935 a_11322_45546# a_13777_45326# 2.22e-21
C39936 a_10903_43370# a_n2293_43922# 0.029114f
C39937 a_12005_46116# a_n2661_43922# 2.87e-22
C39938 a_768_44030# a_6031_43396# 3.88e-20
C39939 a_11453_44696# a_14579_43548# 1.66e-22
C39940 a_n881_46662# a_6655_43762# 2.11e-20
C39941 a_n971_45724# a_n1423_42826# 1.4e-20
C39942 a_n2438_43548# a_n2012_43396# 0.003029f
C39943 a_16327_47482# a_16243_43396# 0.295263f
C39944 a_11415_45002# a_20512_43084# 0.001234f
C39945 a_4883_46098# a_10341_43396# 4.87e-19
C39946 a_10227_46804# a_15781_43660# 0.002214f
C39947 a_11823_42460# a_13017_45260# 0.030503f
C39948 a_7499_43078# a_1307_43914# 0.109806f
C39949 a_17715_44484# a_9313_44734# 6.46e-20
C39950 a_12861_44030# a_18783_43370# 2.29e-20
C39951 a_18479_45785# a_19610_45572# 8.18e-19
C39952 a_18341_45572# a_19365_45572# 2.36e-20
C39953 a_3090_45724# a_10949_43914# 0.001234f
C39954 a_22545_38993# RST_Z 1.94e-21
C39955 C10_P_btm C8_P_btm 0.878696f
C39956 a_4883_46098# a_12991_46634# 8.79e-20
C39957 a_10227_46804# a_15227_44166# 0.013242f
C39958 a_171_46873# a_n2661_46098# 0.168482f
C39959 a_383_46660# a_479_46660# 0.013793f
C39960 a_601_46902# a_645_46660# 3.69e-19
C39961 a_33_46660# a_1799_45572# 3.91e-21
C39962 a_9804_47204# a_9863_46634# 0.017882f
C39963 a_13717_47436# a_13885_46660# 0.003475f
C39964 a_12861_44030# a_13170_46660# 9.11e-20
C39965 a_n133_46660# a_2443_46660# 4.17e-21
C39966 a_n2438_43548# a_2609_46660# 8.62e-19
C39967 a_5807_45002# a_6540_46812# 0.007069f
C39968 a_4915_47217# a_765_45546# 0.169406f
C39969 EN_VIN_BSTR_P C0_P_btm 0.12803f
C39970 a_n1925_46634# a_3699_46634# 0.014429f
C39971 a_22821_38993# VDD 0.431879f
C39972 a_n2833_47464# a_n2840_46090# 2.94e-20
C39973 a_18479_47436# a_17609_46634# 3.14e-19
C39974 a_3905_42865# a_3905_42558# 2.95e-19
C39975 a_16243_43396# a_16855_43396# 3.82e-19
C39976 a_10341_43396# a_5649_42852# 0.049047f
C39977 a_n2661_42282# a_196_42282# 2.77e-19
C39978 a_15743_43084# a_19268_43646# 0.010228f
C39979 a_6031_43396# a_5755_42852# 4.17e-19
C39980 a_3626_43646# a_8952_43230# 9.54e-21
C39981 a_2982_43646# a_10518_42984# 2.29e-20
C39982 a_10775_45002# CLK 0.058141f
C39983 a_n97_42460# a_18249_42858# 0.003512f
C39984 a_14797_45144# VDD 0.124624f
C39985 a_9482_43914# a_13490_45067# 0.007606f
C39986 a_13348_45260# a_13807_45067# 6.64e-19
C39987 a_4791_45118# a_5421_42558# 0.00311f
C39988 a_n863_45724# a_261_44278# 9.97e-19
C39989 a_n745_45366# a_n2129_44697# 0.00194f
C39990 a_n2293_45010# a_n1352_44484# 0.020183f
C39991 a_n2661_45010# a_742_44458# 0.694478f
C39992 a_n2017_45002# a_n1917_44484# 0.012037f
C39993 a_n913_45002# a_n2267_44484# 1.1e-19
C39994 a_3357_43084# a_6298_44484# 3.5e-19
C39995 a_10903_43370# a_n97_42460# 0.021999f
C39996 a_14537_43396# a_14403_45348# 2.86e-19
C39997 a_n443_42852# a_2889_44172# 1.05e-20
C39998 a_n2956_37592# a_n2661_44458# 0.003435f
C39999 en_comp a_n4318_40392# 3.37e-20
C40000 a_13507_46334# a_22765_42852# 0.003797f
C40001 a_13259_45724# a_15682_43940# 9.31e-21
C40002 a_13507_46334# a_16375_45002# 0.002576f
C40003 a_4883_46098# a_18147_46436# 2.8e-19
C40004 a_n2661_46634# a_10809_44734# 0.023983f
C40005 a_4817_46660# a_5164_46348# 5.41e-19
C40006 a_4955_46873# a_5204_45822# 3.57e-19
C40007 a_2063_45854# a_2711_45572# 0.185507f
C40008 a_13885_46660# a_14035_46660# 0.25868f
C40009 a_17609_46634# a_17829_46910# 0.111805f
C40010 a_18597_46090# a_20009_46494# 8.96e-19
C40011 a_8128_46384# a_8062_46482# 7.91e-19
C40012 a_n881_46662# a_6633_46155# 8.73e-19
C40013 a_15227_44166# a_17339_46660# 0.524034f
C40014 a_n2840_46634# a_n2956_39304# 0.001899f
C40015 a_n971_45724# a_3775_45552# 0.091275f
C40016 a_n237_47217# a_6598_45938# 2.15e-19
C40017 a_4646_46812# a_6165_46155# 3.41e-20
C40018 a_3877_44458# a_6419_46155# 0.002843f
C40019 a_4651_46660# a_5497_46414# 2.21e-19
C40020 a_n443_46116# a_n443_42852# 0.145452f
C40021 a_5257_43370# a_1823_45246# 0.003231f
C40022 a_18479_47436# a_19443_46116# 3.9e-22
C40023 a_12465_44636# a_14383_46116# 0.00348f
C40024 a_3422_30871# C1_N_btm 7.67e-20
C40025 a_21356_42826# a_21195_42852# 0.03853f
C40026 a_14209_32519# a_22400_42852# 8.65e-21
C40027 a_3626_43646# a_15521_42308# 3.81e-19
C40028 a_20766_44850# VDD 0.197657f
C40029 a_8605_42826# a_8495_42852# 0.097745f
C40030 a_626_44172# a_895_43940# 0.038336f
C40031 a_9482_43914# a_7845_44172# 5.64e-21
C40032 a_11827_44484# a_12829_44484# 2.53e-19
C40033 a_n357_42282# a_18525_43370# 3.71e-20
C40034 a_n443_42852# a_14621_43646# 0.001398f
C40035 a_19778_44110# a_17517_44484# 0.018823f
C40036 a_1307_43914# a_3600_43914# 0.153686f
C40037 a_9049_44484# a_8791_43396# 1.63e-20
C40038 a_7499_43078# a_9396_43370# 2.11e-19
C40039 a_3232_43370# a_5841_44260# 5.8e-19
C40040 a_3537_45260# a_8333_44056# 0.012371f
C40041 a_17970_44736# a_18287_44626# 0.102355f
C40042 a_13249_42308# a_3626_43646# 0.007551f
C40043 a_5518_44484# a_6109_44484# 0.050093f
C40044 a_5343_44458# a_7640_43914# 0.152634f
C40045 a_11691_44458# a_11541_44484# 0.037586f
C40046 a_4185_45028# a_5193_42852# 2.2e-19
C40047 a_526_44458# a_9127_43156# 0.054699f
C40048 a_13507_46334# a_413_45260# 3.41e-19
C40049 a_13759_46122# a_15682_46116# 1.44e-20
C40050 a_13925_46122# a_2324_44458# 4.65e-20
C40051 a_14493_46090# a_14840_46494# 0.051162f
C40052 a_2698_46116# a_n1925_42282# 1.04e-20
C40053 a_1823_45246# a_1337_46116# 1.69e-19
C40054 a_3147_46376# a_2981_46116# 0.003565f
C40055 a_2804_46116# a_526_44458# 0.00297f
C40056 a_9863_46634# a_10180_45724# 1.87e-19
C40057 a_10150_46912# a_10053_45546# 1.88e-20
C40058 a_8667_46634# a_8746_45002# 4.9e-22
C40059 a_n443_46116# a_375_42282# 0.001544f
C40060 a_19321_45002# a_19431_45546# 0.029441f
C40061 a_13661_43548# a_18799_45938# 0.004963f
C40062 a_13747_46662# a_18596_45572# 0.01625f
C40063 a_5807_45002# a_16789_45572# 1.08e-19
C40064 a_n881_46662# a_2437_43646# 0.084076f
C40065 a_2905_45572# a_3495_45348# 3.62e-20
C40066 a_6755_46942# a_6812_45938# 2.21e-20
C40067 a_8953_45546# a_6945_45028# 2.77e-19
C40068 a_8199_44636# a_10809_44734# 0.022266f
C40069 SMPL_ON_N en_comp 8.94e-19
C40070 a_22959_42860# a_22465_38105# 9e-19
C40071 a_1606_42308# a_1755_42282# 0.278431f
C40072 a_13291_42460# a_13657_42558# 0.026223f
C40073 a_7287_43370# VDD 0.457521f
C40074 a_n784_42308# a_5379_42460# 1.36e-19
C40075 a_n2433_44484# a_n2129_43609# 4.74e-21
C40076 a_n2017_45002# a_n1853_43023# 0.03086f
C40077 a_n2661_45010# a_n901_43156# 1.36e-21
C40078 a_n1059_45260# a_n2157_42858# 1.41e-19
C40079 a_n913_45002# a_n2472_42826# 7.39e-21
C40080 a_n2293_45010# a_n1423_42826# 4.06e-19
C40081 a_n2840_43914# a_n2065_43946# 6.33e-21
C40082 a_3065_45002# a_743_42282# 0.040577f
C40083 a_n863_45724# a_2351_42308# 0.038802f
C40084 a_n755_45592# a_961_42354# 0.01273f
C40085 a_2711_45572# a_19326_42852# 1.2e-19
C40086 a_8975_43940# a_9420_43940# 2.6e-19
C40087 a_10057_43914# a_9801_43940# 0.006215f
C40088 a_8492_46660# VDD 0.273866f
C40089 a_9313_44734# a_20623_43914# 4.63e-20
C40090 a_1307_43914# a_15781_43660# 2.51e-20
C40091 a_n2661_45546# a_3218_45724# 0.010947f
C40092 a_n1079_45724# a_n755_45592# 0.109544f
C40093 a_n2293_46634# a_6298_44484# 1.21e-19
C40094 a_20623_46660# a_413_45260# 2.82e-20
C40095 a_22959_46660# a_20447_31679# 3.72e-20
C40096 a_13507_46334# a_13468_44734# 1.04e-19
C40097 a_n863_45724# a_n357_42282# 0.172013f
C40098 a_380_45546# a_n1099_45572# 0.148825f
C40099 a_5807_45002# a_14539_43914# 0.066683f
C40100 a_13661_43548# a_16112_44458# 0.053099f
C40101 a_2324_44458# a_15599_45572# 0.042604f
C40102 a_13351_46090# a_8696_44636# 5.82e-22
C40103 a_15227_44166# a_1307_43914# 0.059667f
C40104 a_8034_45724# a_7499_43078# 0.001227f
C40105 a_8049_45260# a_6812_45938# 2.61e-19
C40106 a_10623_46897# a_n2661_43370# 6.28e-21
C40107 a_n971_45724# a_n1549_44318# 0.00442f
C40108 a_n452_45724# a_310_45028# 5.77e-21
C40109 a_12465_44636# a_n2661_42834# 7.41e-19
C40110 COMP_P a_22609_38406# 0.00369f
C40111 a_7174_31319# a_1239_39587# 2.3e-19
C40112 a_n4064_40160# a_n2302_40160# 0.249627f
C40113 a_n4334_40480# a_n4251_40480# 0.007692f
C40114 a_n4315_30879# a_n2216_40160# 0.001403f
C40115 a_n1920_47178# a_n1151_42308# 8.17e-19
C40116 a_n785_47204# a_1209_47178# 3.43e-19
C40117 a_n23_47502# a_1239_47204# 8.7e-21
C40118 a_n2109_47186# a_3381_47502# 0.035813f
C40119 a_n1741_47186# a_3160_47472# 0.012286f
C40120 a_n237_47217# a_1431_47204# 0.045044f
C40121 a_n971_45724# a_584_46384# 0.152617f
C40122 a_1606_42308# VDAC_P 0.006306f
C40123 a_11967_42832# a_17324_43396# 8.32e-19
C40124 a_12607_44458# a_12379_42858# 3.9e-21
C40125 a_21115_43940# a_21381_43940# 0.073198f
C40126 a_11341_43940# a_19741_43940# 0.003328f
C40127 a_15493_43940# a_19478_44056# 6.87e-19
C40128 a_n913_45002# a_9223_42460# 8.58e-19
C40129 a_n1059_45260# a_9803_42558# 8.94e-21
C40130 a_n2017_45002# a_9293_42558# 0.001147f
C40131 a_14955_43940# a_n97_42460# 6.16e-22
C40132 a_n2661_42282# a_4699_43561# 1.76e-21
C40133 a_7281_43914# a_6197_43396# 3.25e-19
C40134 a_2382_45260# a_5932_42308# 4.34e-21
C40135 a_18479_45785# a_19332_42282# 2.44e-19
C40136 a_5210_46155# VDD 6.34e-20
C40137 a_n356_44636# a_3681_42891# 1.42e-20
C40138 a_n2293_43922# a_5649_42852# 1.78418f
C40139 a_20692_30879# a_22469_39537# 6.23e-20
C40140 a_n2293_46098# a_5205_44734# 5.05e-20
C40141 a_12861_44030# a_3626_43646# 3.03e-20
C40142 a_15227_44166# a_18579_44172# 9.13e-21
C40143 a_n2312_39304# a_n4318_39304# 0.023404f
C40144 a_768_44030# a_6671_43940# 1.23e-19
C40145 a_8199_44636# a_5883_43914# 7.86e-19
C40146 a_5937_45572# a_8701_44490# 0.022661f
C40147 a_8016_46348# a_10157_44484# 0.016596f
C40148 a_3483_46348# a_16979_44734# 0.173123f
C40149 a_15765_45572# a_16333_45814# 0.17072f
C40150 a_15599_45572# a_16855_45546# 0.043567f
C40151 a_15903_45785# a_16115_45572# 3.12e-19
C40152 a_n443_42852# a_3537_45260# 0.567413f
C40153 a_376_46348# a_n356_44636# 3.01e-22
C40154 a_19692_46634# a_19279_43940# 8.61e-20
C40155 a_4883_46098# a_n97_42460# 1.42e-20
C40156 a_n4251_38528# VDD 3.95e-19
C40157 a_2063_45854# a_8654_47026# 1.72e-19
C40158 a_8912_37509# VDAC_P 3.15325f
C40159 VDAC_N a_11206_38545# 0.15219f
C40160 a_6886_37412# CAL_N 1.24e-19
C40161 a_6151_47436# a_10150_46912# 0.006237f
C40162 a_6575_47204# a_7577_46660# 3.98e-19
C40163 a_7903_47542# a_8145_46902# 0.010369f
C40164 a_4915_47217# a_10623_46897# 0.002626f
C40165 a_n881_46662# a_n2661_46634# 0.035376f
C40166 a_768_44030# a_13747_46662# 0.434325f
C40167 a_19479_31679# C4_N_btm 9.91e-21
C40168 a_458_43396# a_743_42282# 3.19e-21
C40169 a_9145_43396# a_14579_43548# 0.024497f
C40170 a_8685_43396# a_10341_43396# 2.41562f
C40171 a_n2293_43922# a_7963_42308# 3.54e-20
C40172 a_n2661_42282# a_6101_43172# 7.12e-20
C40173 a_15493_43940# a_17701_42308# 2.87e-20
C40174 a_11341_43940# a_17333_42852# 1.63e-20
C40175 a_n97_42460# a_5649_42852# 0.008438f
C40176 a_3626_43646# a_19700_43370# 7.81e-19
C40177 a_n356_44636# a_15959_42545# 0.001149f
C40178 a_17730_32519# a_22400_42852# 1.31e-20
C40179 a_19862_44208# a_19987_42826# 2.09e-19
C40180 a_10775_45002# a_10951_45334# 0.185422f
C40181 a_20202_43084# a_14401_32519# 9.39e-20
C40182 a_2382_45260# a_1423_45028# 0.036767f
C40183 a_4558_45348# a_1307_43914# 1.16e-20
C40184 a_2274_45254# a_2232_45348# 0.002765f
C40185 a_13259_45724# a_20512_43084# 1.37e-20
C40186 a_768_44030# a_10796_42968# 2.7e-22
C40187 a_6171_45002# a_14180_45002# 0.012672f
C40188 a_2711_45572# a_n2661_42834# 2.44e-21
C40189 a_413_45260# a_2903_45348# 4.7e-19
C40190 a_17715_44484# a_17737_43940# 0.289085f
C40191 a_16147_45260# a_11827_44484# 7.51e-20
C40192 a_1823_45246# a_5745_43940# 9.33e-20
C40193 a_4883_46098# a_17957_46116# 0.013641f
C40194 a_18780_47178# a_6945_45028# 0.013003f
C40195 a_18479_47436# a_22223_46124# 5.82e-20
C40196 a_n2661_46634# a_n2157_46122# 1.89e-19
C40197 a_n2472_46634# a_n2293_46098# 0.00197f
C40198 a_n2442_46660# a_n2472_46090# 6.07e-19
C40199 a_11453_44696# a_14840_46494# 7.84e-22
C40200 a_13507_46334# a_18985_46122# 0.002665f
C40201 a_18143_47464# a_10809_44734# 0.006426f
C40202 a_n743_46660# a_12741_44636# 9.6e-19
C40203 a_n1435_47204# a_n1925_42282# 4.56e-21
C40204 a_6755_46942# a_15559_46634# 1.64e-19
C40205 a_n881_46662# a_8199_44636# 2.26e-20
C40206 a_n1613_43370# a_5937_45572# 0.117604f
C40207 a_12465_44636# a_17715_44484# 1.19e-20
C40208 a_768_44030# a_4419_46090# 2.08e-20
C40209 a_8037_42858# a_8952_43230# 0.118759f
C40210 a_3539_42460# a_1755_42282# 3.25e-19
C40211 a_14621_43646# a_14635_42282# 1.99e-20
C40212 a_4905_42826# a_5267_42460# 0.146764f
C40213 a_4093_43548# a_3905_42558# 4.12e-21
C40214 a_3080_42308# a_5379_42460# 1.73e-20
C40215 a_n23_44458# VDD 0.169093f
C40216 a_n97_42460# a_7963_42308# 0.002153f
C40217 a_n356_44636# RST_Z 2.99e-19
C40218 a_3357_43084# a_2479_44172# 0.0305f
C40219 a_12549_44172# a_17303_42282# 4.74e-21
C40220 a_n863_45724# a_n144_43396# 1.49e-19
C40221 a_17613_45144# a_17767_44458# 0.003f
C40222 a_n2312_39304# a_n4334_40480# 2.31e-19
C40223 a_20202_43084# a_18817_42826# 1.4e-20
C40224 a_n755_45592# a_2982_43646# 0.221452f
C40225 a_n2661_44458# a_n2267_44484# 0.046548f
C40226 a_n2433_44484# a_n2129_44697# 0.130072f
C40227 a_16922_45042# a_18248_44752# 7.57e-20
C40228 a_11827_44484# a_10334_44484# 1.87e-19
C40229 a_n4318_40392# a_n1699_44726# 2.56e-21
C40230 a_n2293_42834# a_8238_44734# 2.49e-21
C40231 a_8137_45348# a_5891_43370# 4.09e-20
C40232 a_n2312_40392# a_n4064_40160# 0.103899f
C40233 a_n913_45002# a_n2065_43946# 0.018244f
C40234 a_n2293_45010# a_n1549_44318# 0.014826f
C40235 a_n2661_45010# a_n984_44318# 2.17e-20
C40236 a_n2017_45002# a_n1899_43946# 0.017371f
C40237 a_n1059_45260# a_n1761_44111# 0.535535f
C40238 a_n443_42852# a_1049_43396# 0.047375f
C40239 a_7499_43078# a_10867_43940# 0.004845f
C40240 w_11334_34010# a_8530_39574# 2.13e-19
C40241 a_4646_46812# a_5379_42460# 1.84e-21
C40242 a_16327_47482# a_18341_45572# 0.04767f
C40243 a_11415_45002# a_10903_43370# 0.085164f
C40244 a_n2497_47436# a_2382_45260# 0.042349f
C40245 a_1823_45246# a_3699_46348# 2.62e-19
C40246 a_2202_46116# a_3483_46348# 9.66e-20
C40247 a_4007_47204# a_3357_43084# 1.6e-20
C40248 a_11453_44696# a_16115_45572# 1.16e-20
C40249 a_10227_46804# a_16377_45572# 1.61e-19
C40250 a_20107_46660# a_19900_46494# 1.04e-19
C40251 a_20411_46873# a_20075_46420# 0.007002f
C40252 a_11735_46660# a_12638_46436# 1.61e-19
C40253 a_11813_46116# a_12379_46436# 0.001157f
C40254 a_18285_46348# a_6945_45028# 1.31e-19
C40255 a_n746_45260# a_n967_45348# 0.028689f
C40256 a_n443_46116# a_2437_43646# 0.410719f
C40257 a_584_46384# a_n2293_45010# 0.02901f
C40258 a_n971_45724# a_n659_45366# 3.11e-21
C40259 a_n1741_47186# a_413_45260# 0.026099f
C40260 a_167_45260# a_3147_46376# 3.32e-19
C40261 a_n2293_46098# a_5937_45572# 0.078393f
C40262 a_15559_46634# a_8049_45260# 3.55e-20
C40263 a_765_45546# a_10809_44734# 2.52248f
C40264 a_2107_46812# a_6511_45714# 3.47e-20
C40265 a_11599_46634# a_18596_45572# 0.01377f
C40266 a_5342_30871# a_13575_42558# 4.35e-19
C40267 a_9420_43940# VDD 0.0046f
C40268 a_5534_30871# a_13249_42558# 0.002316f
C40269 a_13460_43230# a_13657_42558# 2.98e-19
C40270 a_13635_43156# a_14113_42308# 0.002123f
C40271 a_11827_44484# a_13565_44260# 4.08e-19
C40272 a_20820_30879# a_22775_42308# 5.97e-21
C40273 a_16750_47204# VDD 6.26e-19
C40274 a_626_44172# a_458_43396# 0.065365f
C40275 a_19594_46812# START 0.020669f
C40276 a_5883_43914# a_8018_44260# 2.21e-19
C40277 a_n2012_44484# a_n4318_39768# 4.36e-19
C40278 a_3537_45260# a_6655_43762# 0.031868f
C40279 a_19321_45002# SINGLE_ENDED 1.12e-19
C40280 a_10193_42453# a_12089_42308# 0.005996f
C40281 a_6431_45366# a_6197_43396# 9.15e-21
C40282 a_n357_42282# a_7309_42852# 0.016177f
C40283 a_526_44458# a_1755_42282# 0.006616f
C40284 a_n1925_42282# a_1606_42308# 0.065478f
C40285 a_13259_45724# a_16245_42852# 2.29e-20
C40286 a_1307_43914# a_1756_43548# 0.267667f
C40287 a_17517_44484# a_20159_44458# 0.026718f
C40288 a_3065_45002# a_2813_43396# 3.35e-21
C40289 a_5111_44636# a_8147_43396# 0.08322f
C40290 a_22612_30879# C9_N_btm 0.003123f
C40291 a_21588_30879# C10_N_btm 0.002325f
C40292 a_n2017_45002# a_14358_43442# 2.42e-20
C40293 a_n1059_45260# a_14579_43548# 0.250544f
C40294 a_9290_44172# a_11551_42558# 0.123803f
C40295 a_526_44458# a_n1099_45572# 1.36e-19
C40296 a_n743_46660# a_n2293_42834# 6.42e-20
C40297 a_7411_46660# a_7229_43940# 3.82e-19
C40298 a_5807_45002# a_14309_45028# 0.003656f
C40299 a_13661_43548# a_13807_45067# 4.93e-20
C40300 a_4791_45118# a_5205_44734# 0.001884f
C40301 a_15368_46634# a_3357_43084# 5.03e-20
C40302 a_17715_44484# a_2711_45572# 0.009119f
C40303 a_n2956_39768# a_n2661_43370# 1.14e-19
C40304 a_12861_44030# a_17767_44458# 2.43e-19
C40305 a_n2312_39304# a_n2661_44458# 1.84e-20
C40306 a_n1151_42308# a_5891_43370# 9.29e-22
C40307 a_12549_44172# a_19778_44110# 0.294084f
C40308 a_5937_45572# a_7230_45938# 7.84e-20
C40309 a_8349_46414# a_8568_45546# 0.001282f
C40310 a_8016_46348# a_7499_43078# 7.22e-19
C40311 a_3483_46348# a_11823_42460# 0.377948f
C40312 a_8199_44636# a_8162_45546# 0.119979f
C40313 a_7715_46873# a_7276_45260# 4.09e-20
C40314 a_5342_30871# C3_N_btm 8.34e-20
C40315 a_n4318_38216# a_n4251_38304# 2.47e-19
C40316 a_5932_42308# a_1239_39587# 2.77e-19
C40317 a_12563_42308# a_7174_31319# 9.76e-21
C40318 a_5534_30871# C5_N_btm 8.45e-20
C40319 a_n4318_37592# a_n3420_37984# 0.404896f
C40320 a_n3674_38216# a_n4064_37984# 0.65176f
C40321 a_14113_42308# a_18310_42308# 4.09e-21
C40322 a_12089_42308# VDD 0.807892f
C40323 a_18248_44752# a_15743_43084# 8.41e-20
C40324 a_18443_44721# a_18525_43370# 0.001063f
C40325 a_18287_44626# a_18783_43370# 4.14e-20
C40326 a_18374_44850# a_18429_43548# 2e-20
C40327 a_n356_44636# a_16243_43396# 4.44e-20
C40328 a_14539_43914# a_16867_43762# 0.004505f
C40329 a_9313_44734# a_15095_43370# 0.039448f
C40330 a_10193_42453# a_18907_42674# 0.002509f
C40331 a_n2956_38216# a_n4064_38528# 3.3e-20
C40332 a_19328_44172# a_15493_43396# 0.019584f
C40333 a_4223_44672# a_4361_42308# 7.99e-22
C40334 a_n2065_43946# a_n4318_39304# 3.62e-19
C40335 a_n2472_43914# a_n2433_43396# 7.88e-19
C40336 a_7542_44172# a_7499_43940# 0.157633f
C40337 a_5497_46414# VDD 0.200657f
C40338 a_18451_43940# a_19478_44306# 1.92e-19
C40339 a_13483_43940# a_11341_43940# 0.005417f
C40340 a_n2293_43922# a_8685_43396# 0.026511f
C40341 a_10180_45724# a_10210_45822# 0.006836f
C40342 a_8746_45002# a_8697_45822# 3e-20
C40343 a_10053_45546# a_10907_45822# 0.003363f
C40344 a_5937_45572# a_8704_45028# 0.010036f
C40345 a_n1613_43370# a_8333_44056# 1.05e-20
C40346 a_11823_42460# a_14495_45572# 0.023559f
C40347 a_8162_45546# a_8192_45572# 0.134163f
C40348 a_2711_45572# a_15861_45028# 0.02395f
C40349 a_n2438_43548# a_644_44056# 4.81e-19
C40350 a_3090_45724# a_7640_43914# 0.020595f
C40351 a_13507_46334# a_22223_43948# 0.00424f
C40352 a_12741_44636# a_17969_45144# 3.55e-19
C40353 a_n2293_46634# a_2479_44172# 0.00465f
C40354 a_13059_46348# a_13076_44458# 7.55e-19
C40355 a_n971_45724# a_n1177_43370# 0.014733f
C40356 a_2324_44458# a_5837_45348# 3.04e-19
C40357 a_18727_42674# RST_Z 3.5e-20
C40358 a_n2109_47186# a_2959_46660# 1.8e-19
C40359 a_n1741_47186# a_2609_46660# 8.05e-20
C40360 a_n443_46116# a_n2661_46634# 0.121882f
C40361 a_13487_47204# a_13569_47204# 0.014524f
C40362 a_13717_47436# a_13759_47204# 0.013673f
C40363 a_12861_44030# a_13675_47204# 0.001416f
C40364 a_7174_31319# C1_N_btm 5.34e-20
C40365 a_n4064_40160# C9_P_btm 0.003109f
C40366 a_15507_47210# a_12549_44172# 7.15e-20
C40367 a_11599_46634# a_768_44030# 0.018831f
C40368 a_n746_45260# a_1110_47026# 5.54e-20
C40369 a_3160_47472# a_n743_46660# 0.011563f
C40370 a_2905_45572# a_n2438_43548# 2.97e-21
C40371 a_13258_32519# C4_N_btm 2.18e-19
C40372 a_18907_42674# VDD 0.148872f
C40373 a_n4209_38216# a_n2946_37690# 5.11e-19
C40374 a_n3690_38304# a_n3565_37414# 6.38e-20
C40375 a_n3420_37984# a_n4334_37440# 0.008459f
C40376 a_n3565_38216# a_n3690_37440# 7.25e-19
C40377 a_7754_39632# a_7754_39300# 0.296258f
C40378 a_3381_47502# a_n1925_46634# 2.29e-21
C40379 a_n1151_42308# a_n1021_46688# 0.105326f
C40380 a_1431_47204# a_1123_46634# 0.012069f
C40381 a_1239_47204# a_948_46660# 1.6e-20
C40382 a_584_46384# a_601_46902# 0.00376f
C40383 a_1209_47178# a_2107_46812# 2.05e-19
C40384 a_n2661_42282# a_1847_42826# 2.73e-20
C40385 a_15493_43940# a_4361_42308# 7.71e-20
C40386 a_n97_42460# a_8685_43396# 1.81e-19
C40387 a_9241_45822# VDD 0.003665f
C40388 a_11341_43940# a_13678_32519# 0.001425f
C40389 a_9313_44734# a_14097_32519# 0.053061f
C40390 a_3499_42826# a_3935_42891# 7.16e-19
C40391 a_n357_42282# a_16979_44734# 5e-21
C40392 a_6511_45714# a_n2661_44458# 1.46e-20
C40393 a_n2293_46634# a_9885_43396# 1.99e-19
C40394 a_4646_46812# a_7287_43370# 0.07176f
C40395 a_n2017_45002# en_comp 0.004677f
C40396 a_n1059_45260# a_n2956_37592# 2.56e-20
C40397 a_2437_43646# a_3537_45260# 2.74e-21
C40398 a_n2109_45247# a_n967_45348# 1e-19
C40399 a_13661_43548# a_17499_43370# 8.74e-19
C40400 a_n2661_45010# a_n467_45028# 0.227953f
C40401 a_1138_42852# a_1241_44260# 6.56e-19
C40402 a_16147_45260# a_15595_45028# 0.00203f
C40403 a_n443_42852# a_8701_44490# 2.96e-20
C40404 a_13059_46348# a_15301_44260# 1e-19
C40405 a_n237_47217# a_2324_44458# 1.65e-19
C40406 a_5807_45002# a_12347_46660# 0.001248f
C40407 a_12891_46348# a_13059_46348# 0.372745f
C40408 a_12549_44172# a_15227_46910# 0.008471f
C40409 a_n1435_47204# a_2698_46116# 2.19e-21
C40410 a_9313_45822# a_3483_46348# 0.087132f
C40411 a_21811_47423# a_20202_43084# 1.66e-20
C40412 a_21177_47436# a_12741_44636# 4.05e-21
C40413 a_4883_46098# a_11415_45002# 1.14e-19
C40414 a_13507_46334# a_20820_30879# 3.67e-19
C40415 a_5732_46660# a_5257_43370# 0.001523f
C40416 a_5072_46660# a_5263_46660# 4.61e-19
C40417 a_n1151_42308# a_9290_44172# 0.10853f
C40418 a_n881_46662# a_765_45546# 0.333008f
C40419 DATA[5] CLK 0.059607f
C40420 a_6151_47436# a_6419_46155# 0.004367f
C40421 a_4791_45118# a_5937_45572# 0.151145f
C40422 a_20916_46384# a_19692_46634# 0.117693f
C40423 a_2063_45854# a_12005_46116# 0.051126f
C40424 a_4646_46812# a_8492_46660# 2.79e-21
C40425 a_n97_42460# a_15953_42852# 0.001782f
C40426 a_17538_32519# a_22400_42852# 1.17e-20
C40427 a_10341_43396# a_17333_42852# 3.64e-20
C40428 a_21005_45260# VDD 0.184261f
C40429 a_10807_43548# a_11551_42558# 0.001883f
C40430 a_11415_45002# a_5649_42852# 2.71e-20
C40431 a_n2442_46660# a_n3674_38216# 0.023932f
C40432 a_9290_44172# a_12293_43646# 9.78e-19
C40433 a_13259_45724# a_21381_43940# 9.63e-21
C40434 a_n2661_45010# a_n2661_43922# 0.111071f
C40435 a_10227_46804# a_13657_42558# 8.38e-19
C40436 a_n2312_38680# a_n2472_42282# 2.73e-20
C40437 SMPL_ON_P a_n2946_39866# 1.96e-20
C40438 a_13556_45296# a_13076_44458# 8.16e-20
C40439 a_9482_43914# a_13720_44458# 0.188323f
C40440 a_1423_45028# a_5343_44458# 0.128331f
C40441 a_1307_43914# a_9838_44484# 5.82e-22
C40442 a_n1925_42282# a_3539_42460# 0.024736f
C40443 a_3232_43370# a_n356_44636# 1.34e-20
C40444 a_18175_45572# a_19279_43940# 9.28e-21
C40445 a_4185_45028# a_17499_43370# 9.45e-21
C40446 a_5257_43370# a_5193_42852# 1.09e-19
C40447 a_n2956_39768# COMP_P 0.003427f
C40448 a_2711_45572# a_20623_43914# 2.17e-19
C40449 a_20623_45572# a_17517_44484# 1.02e-20
C40450 a_20916_46384# a_20692_30879# 0.001701f
C40451 a_21588_30879# a_20205_31679# 0.058932f
C40452 a_12251_46660# a_10903_43370# 5.76e-22
C40453 a_12469_46902# a_12005_46116# 0.003112f
C40454 a_n971_45724# a_8696_44636# 0.003003f
C40455 a_12861_44030# a_12791_45546# 0.248928f
C40456 a_13487_47204# a_11823_42460# 3.88e-21
C40457 a_11599_46634# a_11652_45724# 5.18e-19
C40458 a_n743_46660# a_16375_45002# 0.03035f
C40459 a_8270_45546# a_2324_44458# 0.039817f
C40460 a_20841_46902# a_12741_44636# 0.043075f
C40461 a_20623_46660# a_20820_30879# 8.87e-21
C40462 a_16327_47482# a_10193_42453# 0.163668f
C40463 a_4817_46660# a_5066_45546# 7.24e-20
C40464 a_768_44030# a_1848_45724# 5.61e-19
C40465 a_22000_46634# a_20202_43084# 0.154237f
C40466 a_n1613_43370# a_n443_42852# 0.062474f
C40467 a_20107_46660# a_21297_46660# 2.56e-19
C40468 a_n881_46662# a_509_45822# 0.001201f
C40469 a_11901_46660# a_12594_46348# 1.15e-19
C40470 a_11813_46116# a_13351_46090# 7.95e-20
C40471 a_10249_46116# a_6945_45028# 6.69e-19
C40472 a_4361_42308# a_5742_30871# 0.071684f
C40473 a_743_42282# a_13575_42558# 0.009742f
C40474 a_16137_43396# a_18907_42674# 0.001947f
C40475 a_1847_42826# a_3497_42558# 2.53e-20
C40476 a_19987_42826# a_20573_43172# 0.006947f
C40477 a_18817_42826# a_19326_42852# 2.6e-19
C40478 a_5649_42852# a_10533_42308# 7.52e-20
C40479 a_3681_42891# a_3823_42558# 0.001239f
C40480 a_16759_43396# a_4958_30871# 1.9e-19
C40481 a_16327_47482# VDD 2.81451f
C40482 a_1307_43914# a_12603_44260# 2.49e-19
C40483 a_16241_47178# RST_Z 5.18e-20
C40484 a_16112_44458# a_11967_42832# 2.42e-19
C40485 a_n2433_44484# a_n2472_43914# 9.53e-19
C40486 a_n2661_44458# a_n2065_43946# 8.48e-20
C40487 a_13259_45724# a_18249_42858# 2.6e-19
C40488 a_526_44458# a_9306_43218# 0.001865f
C40489 a_13381_47204# CLK 2.37e-19
C40490 a_n755_45592# a_7871_42858# 0.033537f
C40491 a_n357_42282# a_7765_42852# 0.042157f
C40492 a_n913_45002# a_n2129_43609# 0.023791f
C40493 a_n2810_45028# a_n4318_39304# 0.023142f
C40494 a_n2661_45010# a_n447_43370# 3.19e-22
C40495 a_n2017_45002# a_n1699_43638# 0.004053f
C40496 a_n2293_45010# a_n1177_43370# 0.001252f
C40497 a_8855_44734# a_n2661_43922# 1.87e-20
C40498 a_21137_46414# a_8049_45260# 0.004656f
C40499 a_10903_43370# a_13259_45724# 0.600111f
C40500 a_n2293_46098# a_n443_42852# 0.086171f
C40501 a_1138_42852# a_997_45618# 0.005258f
C40502 a_n2661_46634# a_3537_45260# 9.12e-22
C40503 a_n1613_43370# a_375_42282# 3.94e-20
C40504 a_n2497_47436# a_5343_44458# 7.63e-21
C40505 a_n971_45724# a_n1177_44458# 0.007865f
C40506 a_5807_45002# a_6709_45028# 8.09e-19
C40507 a_n743_46660# a_413_45260# 0.031499f
C40508 a_n2438_43548# a_n37_45144# 2.58e-21
C40509 a_n133_46660# a_n143_45144# 1.25e-21
C40510 a_n2293_46634# a_2680_45002# 0.017731f
C40511 a_13059_46348# a_11322_45546# 2.64e-21
C40512 a_1799_45572# a_n2661_45010# 1.31e-20
C40513 a_10227_46804# a_n2661_43370# 0.033611f
C40514 a_526_44458# a_n1925_42282# 0.213917f
C40515 a_12549_44172# a_9482_43914# 0.06308f
C40516 a_12891_46348# a_13556_45296# 0.29495f
C40517 a_768_44030# a_13348_45260# 1.76e-19
C40518 a_n1925_46634# a_1667_45002# 4.73e-21
C40519 a_1823_45246# a_n755_45592# 0.390511f
C40520 a_167_45260# a_310_45028# 0.035247f
C40521 a_6761_42308# a_5742_30871# 1.69e-20
C40522 a_5342_30871# a_7754_38470# 1.06e-19
C40523 a_4190_30871# C5_N_btm 1.71e-19
C40524 a_22400_42852# a_22465_38105# 0.199207f
C40525 a_8325_42308# a_9223_42460# 8.85e-19
C40526 a_8685_42308# a_8791_42308# 0.147376f
C40527 a_n913_45002# a_21195_42852# 0.002742f
C40528 a_5883_43914# a_6452_43396# 0.001768f
C40529 a_20512_43084# a_20935_43940# 1.43e-20
C40530 a_n356_44636# a_4905_42826# 6.1e-20
C40531 a_16721_46634# RST_Z 5.46e-22
C40532 a_n2293_42834# a_4361_42308# 2.59e-19
C40533 en_comp a_19164_43230# 1.47e-21
C40534 a_n2956_38680# a_n4209_38216# 0.001636f
C40535 a_16922_45042# a_15743_43084# 0.00548f
C40536 a_5244_44056# a_n2661_42282# 1.4e-20
C40537 a_16434_46987# VDD 0.001765f
C40538 a_6194_45824# a_6472_45840# 0.118423f
C40539 a_5907_45546# a_6511_45714# 0.043475f
C40540 a_12549_44172# a_20159_44458# 0.005504f
C40541 a_2324_44458# a_n2017_45002# 5.73e-20
C40542 a_2711_45572# a_3775_45552# 0.044123f
C40543 a_n357_42282# a_11823_42460# 0.063073f
C40544 a_n2293_46098# a_375_42282# 2.05e-20
C40545 a_13747_46662# a_17517_44484# 0.022087f
C40546 a_3483_46348# a_7705_45326# 8.97e-19
C40547 a_20708_46348# a_3357_43084# 0.017189f
C40548 a_13059_46348# a_15060_45348# 0.001051f
C40549 a_19692_46634# a_21101_45002# 2.38e-19
C40550 a_4791_45118# a_8333_44056# 4.81e-20
C40551 a_22223_46124# a_2437_43646# 3.38e-19
C40552 a_6945_45028# a_22223_45572# 3.06e-19
C40553 a_8199_44636# a_3537_45260# 0.199536f
C40554 a_5164_46348# a_6171_45002# 1.28e-19
C40555 a_10586_45546# a_12561_45572# 8.99e-20
C40556 a_5497_46414# a_5691_45260# 1.88e-19
C40557 a_5932_42308# C1_N_btm 0.011049f
C40558 a_4915_47217# a_10227_46804# 0.062269f
C40559 a_5742_30871# a_n1532_35090# 1.92e-19
C40560 a_13381_47204# a_13717_47436# 4.77e-21
C40561 a_n4209_38502# a_n4334_38528# 0.25243f
C40562 a_n3420_39072# a_n3607_38528# 2.09e-19
C40563 a_7174_31319# a_3754_38470# 2.41e-19
C40564 a_n237_47217# a_n310_47570# 6.1e-19
C40565 a_n785_47204# a_n2312_40392# 2.56e-20
C40566 a_5934_30871# C3_P_btm 0.011274f
C40567 a_6123_31319# C1_P_btm 0.011005f
C40568 a_n746_45260# a_n89_47570# 0.004982f
C40569 a_5267_42460# VDD 0.170631f
C40570 a_n1741_47186# a_3094_47570# 2.25e-19
C40571 a_n971_45724# a_2266_47570# 4.39e-19
C40572 a_n2109_47186# a_2266_47243# 0.001164f
C40573 a_18114_32519# a_14097_32519# 0.054468f
C40574 a_19721_31679# a_22400_42852# 3.49e-20
C40575 a_n356_45724# VDD 0.719282f
C40576 a_13483_43940# a_10341_43396# 3.72e-20
C40577 a_10949_43914# a_12281_43396# 5.57e-19
C40578 a_n2956_37592# a_n4315_30879# 0.107228f
C40579 a_15433_44458# a_15567_42826# 4.21e-21
C40580 a_9313_44734# a_22959_42860# 0.174475f
C40581 a_n2293_42834# a_6761_42308# 3.63e-21
C40582 a_2479_44172# a_743_42282# 2.08e-20
C40583 a_n2810_45028# a_n4334_40480# 8.59e-19
C40584 a_n2840_43370# a_n2267_43396# 6.1e-19
C40585 a_n4318_39304# a_n2129_43609# 5.32e-19
C40586 a_11322_45546# a_13556_45296# 1.25e-20
C40587 a_10903_43370# a_n2661_43922# 0.039051f
C40588 a_13259_45724# a_19929_45028# 2.15e-20
C40589 a_12741_44636# a_20397_44484# 1.18e-19
C40590 a_n1613_43370# a_6655_43762# 0.013792f
C40591 a_n971_45724# a_n1991_42858# 8.17e-20
C40592 a_10193_42453# a_14537_43396# 1.09e-19
C40593 a_8192_45572# a_3537_45260# 2.88e-19
C40594 a_16327_47482# a_16137_43396# 2.72e-19
C40595 a_20202_43084# a_20512_43084# 0.130366f
C40596 a_11415_45002# a_21145_44484# 9.18e-20
C40597 a_4883_46098# a_9885_43646# 1.07e-20
C40598 a_10227_46804# a_15681_43442# 0.001396f
C40599 a_n2497_47436# a_n1545_43230# 1.72e-19
C40600 a_11823_42460# a_11963_45334# 0.110904f
C40601 a_11962_45724# a_13159_45002# 2.65e-19
C40602 a_9290_44172# a_13857_44734# 1.78e-19
C40603 a_16375_45002# a_17969_45144# 5.89e-19
C40604 a_12861_44030# a_18525_43370# 1.13e-19
C40605 a_18479_45785# a_19365_45572# 0.001158f
C40606 a_3090_45724# a_10729_43914# 0.135702f
C40607 C10_P_btm C9_P_btm 37.815998f
C40608 a_4883_46098# a_12251_46660# 1.41e-19
C40609 a_10227_46804# a_18834_46812# 2.09e-20
C40610 a_18143_47464# a_17609_46634# 0.001435f
C40611 a_601_46902# a_479_46660# 3.16e-19
C40612 a_171_46873# a_1799_45572# 2.16e-21
C40613 a_9804_47204# a_8492_46660# 8.56e-22
C40614 a_n743_46660# a_2609_46660# 6.69e-20
C40615 a_n2438_43548# a_2443_46660# 0.237765f
C40616 a_5807_45002# a_5732_46660# 9.62e-19
C40617 a_n443_46116# a_765_45546# 0.297346f
C40618 EN_VIN_BSTR_P C1_P_btm 0.110046f
C40619 a_n1925_46634# a_2959_46660# 0.009513f
C40620 a_n133_46660# a_n2661_46098# 0.005588f
C40621 a_22545_38993# VDD 0.536989f
C40622 a_15493_43396# a_19518_43218# 8.64e-20
C40623 a_10341_43396# a_13678_32519# 0.011962f
C40624 a_n2661_42282# a_n473_42460# 1.46e-19
C40625 a_18783_43370# a_19268_43646# 0.001296f
C40626 a_3626_43646# a_9127_43156# 2.22e-19
C40627 a_2982_43646# a_10083_42826# 9.5e-20
C40628 a_n97_42460# a_17333_42852# 0.003266f
C40629 a_8953_45002# CLK 0.310391f
C40630 a_14537_43396# VDD 0.779752f
C40631 a_1307_43914# a_n2661_43370# 1.06e-19
C40632 a_13348_45260# a_13490_45067# 0.005572f
C40633 a_10193_42453# a_20835_44721# 2.06e-19
C40634 a_n863_45724# a_n1441_43940# 4.78e-21
C40635 a_n913_45002# a_n2129_44697# 0.017685f
C40636 a_n2293_45010# a_n1177_44458# 0.00518f
C40637 a_n2661_45010# a_n452_44636# 0.020671f
C40638 a_n2017_45002# a_n1699_44726# 0.002575f
C40639 a_15227_44166# a_17678_43396# 3.54e-19
C40640 a_4791_45118# a_5337_42558# 0.003599f
C40641 a_14180_45002# a_14403_45348# 0.011458f
C40642 a_14537_43396# a_14309_45348# 2.07e-19
C40643 a_13507_46334# a_20753_42852# 7.33e-21
C40644 a_13259_45724# a_14955_43940# 8.97e-22
C40645 a_3357_43084# a_5518_44484# 0.009558f
C40646 a_18799_45938# a_18989_43940# 1.13e-19
C40647 a_n2956_37592# a_n4318_40392# 2.71462f
C40648 a_8696_44636# a_9313_44734# 0.003528f
C40649 a_n443_42852# a_2675_43914# 6.34e-20
C40650 a_4883_46098# a_13259_45724# 0.011246f
C40651 a_13507_46334# a_18243_46436# 6.14e-19
C40652 a_10227_46804# a_20850_46482# 6.4e-19
C40653 a_4955_46873# a_5164_46348# 0.009022f
C40654 a_4817_46660# a_5068_46348# 0.001467f
C40655 a_584_46384# a_2711_45572# 1.02e-20
C40656 a_16292_46812# a_17829_46910# 1.46e-19
C40657 a_18597_46090# a_19597_46482# 0.002198f
C40658 a_17609_46634# a_765_45546# 0.256159f
C40659 a_n971_45724# a_7227_45028# 1.87e-20
C40660 a_n237_47217# a_6667_45809# 2.43e-19
C40661 a_3877_44458# a_6165_46155# 1.87e-19
C40662 a_4646_46812# a_5497_46414# 2.5e-20
C40663 a_4651_46660# a_5204_45822# 2.21e-19
C40664 a_4791_45118# a_n443_42852# 0.02747f
C40665 a_n443_46116# a_509_45822# 0.006202f
C40666 a_16327_47482# a_20850_46155# 2.49e-19
C40667 a_3422_30871# C0_N_btm 6.53e-20
C40668 a_20922_43172# a_21195_42852# 0.119168f
C40669 a_3626_43646# a_17124_42282# 0.004372f
C40670 a_20835_44721# VDD 0.198384f
C40671 a_8037_42858# a_8495_42852# 0.027317f
C40672 a_13887_32519# a_14097_32519# 10.5943f
C40673 a_22591_43396# a_22400_42852# 5.76e-19
C40674 a_9145_43396# a_9223_42460# 1.05e-20
C40675 a_8685_43396# a_10533_42308# 6.52e-23
C40676 a_14539_43914# a_18374_44850# 9.06e-21
C40677 a_626_44172# a_2479_44172# 1.03e-20
C40678 a_11827_44484# a_12553_44484# 2.82e-19
C40679 a_5111_44636# a_n2661_42282# 0.025961f
C40680 a_n443_42852# a_14537_43646# 0.001647f
C40681 a_n2956_39768# a_n4209_39304# 0.001636f
C40682 a_18911_45144# a_17517_44484# 2.31e-19
C40683 a_1307_43914# a_2998_44172# 0.233292f
C40684 a_7499_43078# a_8791_43396# 0.04623f
C40685 a_3232_43370# a_3820_44260# 0.003566f
C40686 a_8270_45546# a_9803_42558# 2.56e-20
C40687 a_3090_45724# a_5932_42308# 2.53e-20
C40688 a_20447_31679# a_15493_43940# 1.09e-20
C40689 a_17767_44458# a_18287_44626# 0.043567f
C40690 a_17970_44736# a_18248_44752# 0.117156f
C40691 a_5343_44458# a_6109_44484# 0.285594f
C40692 a_4223_44672# a_5891_43370# 0.020744f
C40693 a_5518_44484# a_5826_44734# 0.017351f
C40694 a_n2017_45002# a_19862_44208# 1e-20
C40695 a_4185_45028# a_4649_42852# 0.00531f
C40696 a_526_44458# a_8387_43230# 0.032585f
C40697 a_13259_45724# a_5649_42852# 1.92021f
C40698 a_5063_47570# a_3357_43084# 1.58e-19
C40699 a_21177_47436# a_413_45260# 8.97e-20
C40700 a_13925_46122# a_14840_46494# 0.118759f
C40701 a_13759_46122# a_2324_44458# 8.3e-20
C40702 a_2804_46116# a_2981_46116# 0.134298f
C40703 a_2698_46116# a_526_44458# 0.002083f
C40704 a_9863_46634# a_10053_45546# 1.27e-19
C40705 a_13747_46662# a_19256_45572# 0.040187f
C40706 a_13661_43548# a_18596_45572# 7.95e-20
C40707 a_12549_44172# a_20623_45572# 1.26e-21
C40708 a_n1613_43370# a_2437_43646# 0.027497f
C40709 a_n2312_40392# a_n913_45002# 7.85e-21
C40710 a_1138_42852# a_1337_46116# 0.039951f
C40711 a_11901_46660# a_2711_45572# 4.34e-20
C40712 a_4915_47217# a_1307_43914# 5.85e-20
C40713 a_5937_45572# a_6945_45028# 0.22046f
C40714 a_22165_42308# a_21973_42336# 5.76e-19
C40715 a_13291_42460# a_13333_42558# 0.001565f
C40716 a_6547_43396# VDD 0.219105f
C40717 a_n784_42308# a_5267_42460# 1.96e-20
C40718 a_n2433_44484# a_n2433_43396# 0.001566f
C40719 a_14537_43396# a_16137_43396# 2.96e-20
C40720 a_n2017_45002# a_n2157_42858# 0.040763f
C40721 a_n2661_45010# a_n1641_43230# 4.2e-20
C40722 a_n2293_45010# a_n1991_42858# 7.5e-20
C40723 a_n863_45724# a_2123_42473# 0.036254f
C40724 a_n2840_43914# a_n2472_43914# 7.52e-19
C40725 en_comp a_14209_32519# 6.81e-20
C40726 a_n755_45592# a_1184_42692# 0.016193f
C40727 a_n357_42282# a_961_42354# 3.8e-19
C40728 a_8975_43940# a_9165_43940# 0.004776f
C40729 a_8667_46634# VDD 0.39254f
C40730 a_1307_43914# a_15681_43442# 2.36e-20
C40731 a_9313_44734# a_20365_43914# 1.7e-20
C40732 a_21076_30879# a_19963_31679# 0.055082f
C40733 a_4883_46098# a_n2661_43922# 0.022558f
C40734 a_n2661_45546# a_2957_45546# 0.008098f
C40735 a_n2293_45546# a_n755_45592# 0.061822f
C40736 a_3090_45724# a_1423_45028# 0.450367f
C40737 a_20841_46902# a_413_45260# 1.91e-20
C40738 a_13661_43548# a_15004_44636# 0.012894f
C40739 a_12594_46348# a_8696_44636# 1.12e-20
C40740 a_15227_44166# a_16019_45002# 4.44e-19
C40741 a_n2497_47436# a_453_43940# 0.09742f
C40742 a_n2293_46098# a_2437_43646# 0.027185f
C40743 a_n863_45724# a_310_45028# 0.033427f
C40744 a_n452_45724# a_n1099_45572# 0.053931f
C40745 a_n2438_43548# a_949_44458# 1.62911f
C40746 a_n743_46660# a_2779_44458# 1.72e-20
C40747 a_n971_45724# a_n1331_43914# 0.015263f
C40748 a_n746_45260# a_n1899_43946# 2.35e-20
C40749 a_11599_46634# a_17517_44484# 1.5e-21
C40750 a_14097_32519# EN_VIN_BSTR_N 0.031973f
C40751 a_5932_42308# a_3754_38470# 2.78e-19
C40752 COMP_P CAL_P 0.037476f
C40753 a_n4315_30879# a_n4251_40480# 0.00226f
C40754 a_n746_45260# a_1431_47204# 2.26e-19
C40755 a_n2109_47186# a_n1151_42308# 0.235661f
C40756 a_n1741_47186# a_2905_45572# 0.012244f
C40757 a_n237_47217# a_1239_47204# 0.203126f
C40758 a_n971_45724# a_2124_47436# 0.352461f
C40759 a_n785_47204# a_327_47204# 0.237391f
C40760 a_2479_44172# a_2813_43396# 0.115852f
C40761 a_11967_42832# a_17499_43370# 0.006642f
C40762 a_15493_43940# a_18533_43940# 0.052096f
C40763 a_20935_43940# a_21381_43940# 1.53e-19
C40764 a_11341_43940# a_21205_44306# 3.95e-19
C40765 a_n913_45002# a_8791_42308# 0.005212f
C40766 a_n1059_45260# a_9223_42460# 1.29e-20
C40767 a_n2017_45002# a_9803_42558# 0.003827f
C40768 a_n2661_42282# a_4235_43370# 3.96e-21
C40769 a_13483_43940# a_n97_42460# 1.05e-21
C40770 a_6453_43914# a_6197_43396# 0.001638f
C40771 a_3537_45260# a_4921_42308# 0.01091f
C40772 a_19862_44208# a_21845_43940# 7.54e-21
C40773 a_n356_44636# a_2905_42968# 2.11e-20
C40774 a_20205_31679# a_22469_39537# 4.7e-20
C40775 a_20692_30879# a_22821_38993# 8.99e-20
C40776 a_19692_46634# a_20766_44850# 1.17e-21
C40777 a_19466_46812# a_19279_43940# 4.38e-20
C40778 a_8034_45724# a_n2661_43370# 1.49e-20
C40779 a_9290_44172# a_4223_44672# 7.92e-21
C40780 a_1609_45822# a_3065_45002# 3.61e-21
C40781 a_509_45572# a_413_45260# 3.88e-19
C40782 a_n2312_40392# a_n4318_39304# 0.025248f
C40783 a_768_44030# a_5829_43940# 2.06e-19
C40784 a_8199_44636# a_8701_44490# 0.25266f
C40785 a_8016_46348# a_9838_44484# 0.004677f
C40786 a_3483_46348# a_14539_43914# 1.24006f
C40787 a_15037_45618# a_8696_44636# 3.1e-21
C40788 a_15599_45572# a_16115_45572# 0.105995f
C40789 a_15903_45785# a_16333_45814# 2.33e-20
C40790 a_3503_45724# a_3232_43370# 1.73e-19
C40791 a_5937_45572# a_8103_44636# 5.28e-21
C40792 a_2684_37794# VDD 0.286898f
C40793 a_n2497_47436# a_3090_45724# 0.16041f
C40794 VDAC_N VDAC_P 4.74149f
C40795 a_6151_47436# a_9863_46634# 0.0481f
C40796 a_6575_47204# a_7715_46873# 4.64e-19
C40797 a_7903_47542# a_7577_46660# 4e-20
C40798 a_4915_47217# a_10467_46802# 0.003258f
C40799 a_n1613_43370# a_n2661_46634# 0.279652f
C40800 a_15928_47570# a_5807_45002# 1.22e-19
C40801 a_768_44030# a_13661_43548# 0.175469f
C40802 a_12549_44172# a_13747_46662# 0.072812f
C40803 a_9803_43646# a_10695_43548# 0.007519f
C40804 a_9145_43396# a_13667_43396# 0.074541f
C40805 a_n2293_43922# a_6123_31319# 0.080985f
C40806 a_5891_43370# a_5742_30871# 1.08e-19
C40807 a_n2661_42282# a_5837_43172# 7.96e-20
C40808 a_n4318_40392# a_n4251_40480# 0.001483f
C40809 a_15493_43940# a_17595_43084# 1.73e-20
C40810 a_11341_43940# a_18083_42858# 7.11e-21
C40811 a_n4318_39304# a_n2840_42826# 4.88e-19
C40812 a_n356_44636# a_15803_42450# 0.078793f
C40813 a_20731_45938# VDD 0.142103f
C40814 a_n2661_42834# a_5934_30871# 1.84e-21
C40815 a_19862_44208# a_19164_43230# 1.82e-21
C40816 a_3626_43646# a_19268_43646# 7.05e-22
C40817 a_14495_45572# a_14539_43914# 9.15e-22
C40818 a_20202_43084# a_21381_43940# 0.108097f
C40819 a_2274_45254# a_1423_45028# 8.25e-20
C40820 a_10193_42453# a_n356_44636# 2.49128f
C40821 a_n2956_38680# a_n2661_42282# 3.65e-20
C40822 a_19431_45546# a_19778_44110# 0.010264f
C40823 a_18596_45572# a_18587_45118# 4.99e-19
C40824 a_19256_45572# a_18911_45144# 3.16e-19
C40825 a_4574_45260# a_1307_43914# 1.78e-21
C40826 a_17715_44484# a_15682_43940# 0.007815f
C40827 a_17668_45572# a_16922_45042# 4.77e-19
C40828 a_6171_45002# a_13777_45326# 0.010994f
C40829 a_1823_45246# a_5326_44056# 7.22e-20
C40830 a_3090_45724# a_4181_43396# 2.49e-22
C40831 a_n2438_43548# a_n1076_43230# 2.79e-21
C40832 a_4883_46098# a_18189_46348# 0.012818f
C40833 a_18479_47436# a_6945_45028# 0.348097f
C40834 a_n2472_46634# a_n2472_46090# 0.026152f
C40835 a_n2661_46634# a_n2293_46098# 2.67e-19
C40836 a_13507_46334# a_18819_46122# 0.004962f
C40837 a_10227_46804# a_10809_44734# 0.17883f
C40838 a_n1435_47204# a_526_44458# 4.56e-21
C40839 a_6755_46942# a_15368_46634# 0.033754f
C40840 a_n881_46662# a_8349_46414# 7.22e-20
C40841 a_n1613_43370# a_8199_44636# 5.93e-20
C40842 a_12465_44636# a_17583_46090# 1.75e-21
C40843 a_768_44030# a_4185_45028# 0.022613f
C40844 a_4791_45118# a_6633_46155# 0.006879f
C40845 a_4915_47217# a_8034_45724# 7.21e-21
C40846 a_18597_46090# a_20708_46348# 0.003878f
C40847 a_8605_42826# a_8387_43230# 0.209641f
C40848 a_7871_42858# a_10083_42826# 4.52e-21
C40849 a_8037_42858# a_9127_43156# 0.042737f
C40850 a_7765_42852# a_8952_43230# 3.38e-20
C40851 a_3539_42460# a_1606_42308# 2.57e-20
C40852 a_3626_43646# a_1755_42282# 0.119352f
C40853 a_13887_32519# a_22959_42860# 0.012735f
C40854 a_15493_43940# a_21887_42336# 6.82e-21
C40855 a_4905_42826# a_3823_42558# 3.67e-20
C40856 a_n356_44636# VDD 1.17667f
C40857 a_n97_42460# a_6123_31319# 0.182488f
C40858 a_n1059_45260# a_n2065_43946# 7.97e-21
C40859 a_n2661_45010# a_n809_44244# 2.22e-19
C40860 a_n2017_45002# a_n1761_44111# 0.02974f
C40861 a_n2293_45010# a_n1331_43914# 0.02919f
C40862 a_9482_43914# a_17061_44734# 2.21e-21
C40863 en_comp a_17730_32519# 9.67e-20
C40864 a_n2312_40392# a_n4334_40480# 3.26e-19
C40865 a_n2312_39304# a_n4315_30879# 0.033437f
C40866 a_2437_43646# a_2675_43914# 3.12e-21
C40867 a_3483_46348# a_7871_42858# 5.12e-21
C40868 a_4185_45028# a_5755_42852# 4.48e-21
C40869 a_20202_43084# a_18249_42858# 2.75e-20
C40870 a_n357_42282# a_2982_43646# 0.04908f
C40871 a_n2661_44458# a_n2129_44697# 0.035428f
C40872 a_16922_45042# a_17970_44736# 2.81e-20
C40873 a_n2293_42834# a_5891_43370# 0.669411f
C40874 a_n4318_40392# a_n2267_44484# 0.004061f
C40875 a_11827_44484# a_10157_44484# 6.15e-20
C40876 a_15861_45028# a_15682_43940# 8.44e-19
C40877 a_n443_42852# a_1209_43370# 0.010053f
C40878 w_11334_34010# a_7754_38470# 2.62e-19
C40879 a_13259_45724# a_8685_43396# 0.031693f
C40880 a_4883_46098# a_17478_45572# 3.85e-20
C40881 a_16327_47482# a_18479_45785# 0.841261f
C40882 a_11415_45002# a_11387_46155# 3.86e-20
C40883 a_n2497_47436# a_2274_45254# 3.04e-20
C40884 a_1823_45246# a_3483_46348# 0.070929f
C40885 a_11453_44696# a_16333_45814# 2.89e-21
C40886 a_10227_46804# a_16211_45572# 3.48e-19
C40887 a_20107_46660# a_20075_46420# 0.001101f
C40888 a_11813_46116# a_12005_46436# 6.29e-19
C40889 a_12741_44636# a_9290_44172# 0.004434f
C40890 a_n971_45724# a_n967_45348# 0.581053f
C40891 a_n746_45260# en_comp 2.06e-20
C40892 a_4791_45118# a_2437_43646# 0.00511f
C40893 a_12465_44636# a_8696_44636# 0.038471f
C40894 a_2521_46116# a_2698_46116# 0.159555f
C40895 a_167_45260# a_2804_46116# 0.003847f
C40896 a_17339_46660# a_10809_44734# 0.003677f
C40897 a_15368_46634# a_8049_45260# 0.032468f
C40898 a_5807_45002# a_11962_45724# 6.78e-21
C40899 a_2107_46812# a_6472_45840# 4.62e-20
C40900 a_11599_46634# a_19256_45572# 0.051691f
C40901 a_5342_30871# a_13070_42354# 2.82e-21
C40902 a_9165_43940# VDD 0.192035f
C40903 a_2982_43646# CAL_N 0.181412f
C40904 a_5534_30871# a_14456_42282# 4.39e-19
C40905 a_13635_43156# a_13657_42558# 4.38e-19
C40906 a_20843_47204# VDD 0.188032f
C40907 a_19321_45002# START 0.10793f
C40908 a_5883_43914# a_7911_44260# 2.82e-19
C40909 a_3537_45260# a_6452_43396# 0.00408f
C40910 a_19594_46812# RST_Z 3.35e-20
C40911 a_10193_42453# a_12379_42858# 7.83e-20
C40912 a_6171_45002# a_6197_43396# 1.3e-20
C40913 a_n357_42282# a_5837_42852# 0.01329f
C40914 a_526_44458# a_1606_42308# 0.011179f
C40915 a_20202_43084# a_21125_42558# 0.002691f
C40916 a_1307_43914# a_1568_43370# 0.182552f
C40917 a_5205_44484# a_6031_43396# 9.87e-20
C40918 a_2382_45260# a_3457_43396# 0.004922f
C40919 a_17517_44484# a_19615_44636# 0.018532f
C40920 a_5111_44636# a_7112_43396# 0.041581f
C40921 a_21588_30879# C9_N_btm 0.786375f
C40922 a_n2017_45002# a_14579_43548# 0.003714f
C40923 a_9290_44172# a_5742_30871# 0.118117f
C40924 a_10227_46804# a_5883_43914# 2.83e-21
C40925 a_2324_44458# a_4099_45572# 1.48e-20
C40926 a_526_44458# a_380_45546# 8.89e-21
C40927 a_5257_43370# a_7229_43940# 4.91e-22
C40928 SMPL_ON_P a_n2293_43922# 2.28e-19
C40929 a_12638_46436# a_12839_46116# 0.005425f
C40930 a_16292_46812# a_2437_43646# 3.48e-20
C40931 a_14976_45028# a_3357_43084# 3.74e-20
C40932 a_n2312_40392# a_n2661_44458# 2.36e-20
C40933 a_n2312_39304# a_n4318_40392# 0.023465f
C40934 a_12861_44030# a_16979_44734# 5.79e-19
C40935 a_12549_44172# a_18911_45144# 6.77e-20
C40936 a_8199_44636# a_7230_45938# 8.25e-21
C40937 a_5937_45572# a_6812_45938# 3.01e-19
C40938 a_8349_46414# a_8162_45546# 3.15e-21
C40939 a_8016_46348# a_8568_45546# 3.81e-20
C40940 a_3483_46348# a_12427_45724# 1.97e-20
C40941 a_n1630_35242# a_n2302_38778# 5.02e-20
C40942 a_5342_30871# C2_N_btm 7.86e-20
C40943 a_5934_30871# a_n3565_39590# 6.35e-21
C40944 a_5534_30871# C4_N_btm 8.01e-20
C40945 a_n3674_38216# a_n2946_37984# 4.03e-21
C40946 a_14113_42308# a_18220_42308# 1.46e-20
C40947 a_12379_42858# VDD 0.484153f
C40948 a_18443_44721# a_18429_43548# 4.83e-19
C40949 a_18248_44752# a_18783_43370# 4.75e-20
C40950 a_n356_44636# a_16137_43396# 0.001161f
C40951 a_14539_43914# a_16664_43396# 0.001335f
C40952 a_n2017_45002# a_20573_43172# 1.71e-20
C40953 a_3483_46348# DATA[2] 6.68e-19
C40954 a_9313_44734# a_14205_43396# 9.81e-20
C40955 a_10193_42453# a_18727_42674# 0.003839f
C40956 a_n2956_38216# a_n2946_38778# 0.004751f
C40957 a_18451_43940# a_15493_43396# 2.04e-20
C40958 a_n2472_43914# a_n4318_39304# 0.001031f
C40959 a_7281_43914# a_7499_43940# 0.08213f
C40960 a_5204_45822# VDD 0.359177f
C40961 a_18326_43940# a_19478_44306# 3.31e-20
C40962 a_9672_43914# a_9895_44260# 0.011458f
C40963 a_12429_44172# a_11341_43940# 0.001958f
C40964 a_n2661_43922# a_8685_43396# 4.82e-20
C40965 a_13249_42308# a_13657_42308# 1.5e-19
C40966 a_11453_44696# a_15493_43396# 1.19e-21
C40967 a_13163_45724# a_13527_45546# 0.124682f
C40968 a_5066_45546# a_6171_45002# 0.002485f
C40969 a_10053_45546# a_10210_45822# 0.18824f
C40970 a_8016_46348# a_n2661_43370# 0.028709f
C40971 a_5937_45572# a_7735_45067# 6.35e-19
C40972 a_8199_44636# a_8704_45028# 3.64e-19
C40973 a_11415_45002# a_18545_45144# 1.83e-20
C40974 a_16327_47482# a_14021_43940# 0.061511f
C40975 a_11823_42460# a_13249_42308# 0.360411f
C40976 a_9049_44484# a_10907_45822# 9.64e-21
C40977 a_2711_45572# a_8696_44636# 0.02621f
C40978 a_8162_45546# a_8120_45572# 0.005491f
C40979 a_3090_45724# a_6109_44484# 0.001946f
C40980 a_13507_46334# a_11341_43940# 0.162723f
C40981 a_12741_44636# a_17896_45144# 1.01e-19
C40982 a_n971_45724# a_n1917_43396# 0.001021f
C40983 a_10809_44734# a_1307_43914# 2.22e-19
C40984 a_18057_42282# RST_Z 1.94e-20
C40985 a_10227_46804# a_n881_46662# 0.146883f
C40986 a_n2109_47186# a_3177_46902# 1.13e-19
C40987 a_n1741_47186# a_2443_46660# 1.18e-19
C40988 a_4791_45118# a_n2661_46634# 0.026643f
C40989 a_13717_47436# a_13675_47204# 0.006407f
C40990 a_12861_44030# a_13569_47204# 6.43e-19
C40991 a_n1435_47204# a_13759_47204# 5.48e-19
C40992 a_7174_31319# C0_N_btm 0.050478f
C40993 a_11599_46634# a_12549_44172# 0.075725f
C40994 a_14955_47212# a_768_44030# 1.84e-19
C40995 a_n4064_39616# a_n1532_35090# 1.21e-19
C40996 a_n3420_39616# EN_VIN_BSTR_P 0.06758f
C40997 SMPL_ON_P a_n2661_46098# 0.004205f
C40998 a_2905_45572# a_n743_46660# 0.03492f
C40999 a_13258_32519# C3_N_btm 2.18e-19
C41000 a_18727_42674# VDD 0.181095f
C41001 a_n4209_38216# a_n3420_37440# 0.035706f
C41002 a_2113_38308# VDAC_Ni 0.315941f
C41003 a_n3420_37984# a_n4209_37414# 0.03f
C41004 a_n3565_38216# a_n3565_37414# 0.046412f
C41005 VDAC_Pi a_3754_39134# 0.012307f
C41006 a_n4064_40160# C10_P_btm 0.460005f
C41007 a_n1151_42308# a_n1925_46634# 0.105874f
C41008 a_1239_47204# a_1123_46634# 2.42e-19
C41009 a_1209_47178# a_948_46660# 0.002172f
C41010 a_584_46384# a_33_46660# 8.87e-19
C41011 a_11341_43940# a_21855_43396# 0.005468f
C41012 a_15493_43940# a_13467_32519# 1.32e-20
C41013 a_n356_44636# a_n784_42308# 0.084978f
C41014 a_8697_45822# VDD 0.189893f
C41015 a_9313_44734# a_22400_42852# 0.007141f
C41016 a_3499_42826# a_3681_42891# 0.033957f
C41017 a_n443_42852# a_8103_44636# 2.86e-19
C41018 a_n357_42282# a_14539_43914# 0.028064f
C41019 a_3090_45724# a_18797_44260# 9.33e-20
C41020 a_6472_45840# a_n2661_44458# 1.35e-20
C41021 a_20447_31679# a_413_45260# 0.226658f
C41022 a_4646_46812# a_6547_43396# 0.03374f
C41023 a_n2293_45010# a_n967_45348# 0.018659f
C41024 a_n2109_45247# en_comp 0.108653f
C41025 a_3357_43084# a_2382_45260# 0.219664f
C41026 a_n2017_45002# a_n2956_37592# 2.81e-19
C41027 a_13661_43548# a_16759_43396# 9.73e-21
C41028 a_4915_47217# a_13635_43156# 1.83e-20
C41029 a_n913_45002# a_n745_45366# 0.002509f
C41030 a_11415_45002# a_13483_43940# 2.17e-21
C41031 a_16211_45572# a_1307_43914# 1.74e-19
C41032 a_16147_45260# a_15415_45028# 6.7e-19
C41033 a_7499_43078# a_11827_44484# 0.104754f
C41034 a_13059_46348# a_15037_44260# 7.67e-20
C41035 a_12549_44172# a_13693_46688# 1.21e-19
C41036 a_768_44030# a_14543_46987# 3.15e-19
C41037 a_n1435_47204# a_2521_46116# 3.94e-21
C41038 a_4883_46098# a_20202_43084# 0.135688f
C41039 a_20990_47178# a_12741_44636# 5.68e-20
C41040 a_5907_46634# a_5257_43370# 0.070316f
C41041 a_n1151_42308# a_10355_46116# 0.043227f
C41042 a_n881_46662# a_17339_46660# 7.38e-21
C41043 a_n1613_43370# a_765_45546# 0.205521f
C41044 a_13507_46334# a_22591_46660# 1.58e-19
C41045 DATA[4] CLK 1.11e-19
C41046 a_6151_47436# a_6165_46155# 0.00218f
C41047 a_4915_47217# a_8016_46348# 2.37e-20
C41048 a_4791_45118# a_8199_44636# 0.14611f
C41049 a_n743_46660# a_12816_46660# 4.05e-20
C41050 a_2063_45854# a_10903_43370# 0.277624f
C41051 a_3877_44458# a_8492_46660# 1.48e-21
C41052 a_4646_46812# a_8667_46634# 3.58e-21
C41053 a_14401_32519# a_14097_32519# 0.051264f
C41054 a_n97_42460# a_15597_42852# 0.004581f
C41055 a_18494_42460# RST_Z 5.9e-20
C41056 a_10341_43396# a_18083_42858# 5.86e-20
C41057 a_20567_45036# VDD 0.237324f
C41058 a_10807_43548# a_5742_30871# 0.020937f
C41059 a_20202_43084# a_5649_42852# 0.011671f
C41060 a_8953_45546# a_9885_43396# 0.002213f
C41061 a_n2661_45010# a_n2661_42834# 0.01412f
C41062 a_n2312_38680# a_n3674_38680# 0.023204f
C41063 a_n2442_46660# a_n2104_42282# 4.03e-20
C41064 SMPL_ON_P a_n3420_39616# 1.92e-20
C41065 a_9482_43914# a_13076_44458# 0.103066f
C41066 a_13348_45260# a_13720_44458# 2.46e-19
C41067 a_1423_45028# a_4743_44484# 0.022983f
C41068 a_1307_43914# a_5883_43914# 0.289388f
C41069 a_13556_45296# a_12883_44458# 8.08e-20
C41070 a_526_44458# a_3539_42460# 0.213772f
C41071 a_n1925_42282# a_3626_43646# 0.031012f
C41072 a_3483_46348# a_17324_43396# 1.78e-19
C41073 a_20841_45814# a_17517_44484# 4.23e-21
C41074 a_2711_45572# a_20365_43914# 7.09e-19
C41075 a_n2956_39768# a_n4318_37592# 0.02357f
C41076 a_20916_46384# a_20205_31679# 2.22e-19
C41077 a_11901_46660# a_12005_46116# 1.13e-19
C41078 a_12469_46902# a_10903_43370# 1.97e-19
C41079 a_12861_44030# a_11823_42460# 1.2465f
C41080 a_20273_46660# a_12741_44636# 0.540506f
C41081 a_20841_46902# a_20820_30879# 4.77e-20
C41082 a_11599_46634# a_11525_45546# 1.45e-19
C41083 a_22000_46634# a_22365_46825# 0.001038f
C41084 a_21188_46660# a_20202_43084# 0.002416f
C41085 a_765_45546# a_n2293_46098# 0.054689f
C41086 a_n881_46662# a_n906_45572# 3.16e-20
C41087 a_11813_46116# a_12594_46348# 1.68e-19
C41088 a_10467_46802# a_10809_44734# 4.91e-19
C41089 a_4955_46873# a_5066_45546# 0.006456f
C41090 a_12281_43396# a_7174_31319# 4.88e-21
C41091 a_4361_42308# a_11323_42473# 0.009186f
C41092 a_743_42282# a_13070_42354# 0.007989f
C41093 a_13467_32519# a_5742_30871# 0.004687f
C41094 a_16137_43396# a_18727_42674# 0.007994f
C41095 a_18249_42858# a_19326_42852# 1.46e-19
C41096 a_19987_42826# a_20256_43172# 0.043356f
C41097 a_12379_42858# a_n784_42308# 1.29e-20
C41098 a_3681_42891# a_3318_42354# 0.001606f
C41099 a_16977_43638# a_4958_30871# 7.21e-20
C41100 a_16409_43396# a_17303_42282# 7.54e-20
C41101 a_n357_42282# a_7871_42858# 0.035744f
C41102 a_16241_47178# VDD 0.208959f
C41103 a_14537_43396# a_14021_43940# 0.048774f
C41104 a_1307_43914# a_12495_44260# 3.12e-19
C41105 a_5205_44484# a_6671_43940# 0.049504f
C41106 a_15004_44636# a_11967_42832# 3.52e-21
C41107 a_16979_44734# a_17325_44484# 0.013377f
C41108 a_n2661_44458# a_n2472_43914# 0.002397f
C41109 a_n1435_47204# DATA[5] 0.031859f
C41110 a_13259_45724# a_17333_42852# 0.077331f
C41111 a_526_44458# a_9061_43230# 8.29e-19
C41112 a_13556_45296# a_15037_44260# 0.001318f
C41113 a_5111_44636# a_9801_43940# 2.57e-20
C41114 en_comp a_17538_32519# 8.81e-20
C41115 a_15673_47210# RST_Z 1.57e-19
C41116 a_11459_47204# CLK 7.93e-19
C41117 a_n1059_45260# a_n2129_43609# 0.005575f
C41118 a_n2661_45010# a_n1352_43396# 8.59e-22
C41119 a_n913_45002# a_n2433_43396# 5.3e-22
C41120 a_n2017_45002# a_n2267_43396# 0.033995f
C41121 a_8783_44734# a_n2661_43922# 5.11e-21
C41122 a_9313_44734# a_9159_44484# 0.056359f
C41123 a_20708_46348# a_8049_45260# 0.006053f
C41124 a_10903_43370# a_14383_46116# 2.99e-20
C41125 a_1138_42852# a_n755_45592# 0.062548f
C41126 a_1176_45822# a_997_45618# 0.140567f
C41127 a_n2293_46098# a_509_45822# 0.003882f
C41128 a_14180_46812# a_11823_42460# 8.14e-22
C41129 a_14275_46494# a_14371_46494# 0.013793f
C41130 a_n2497_47436# a_4743_44484# 0.003104f
C41131 a_n901_46420# a_n356_45724# 0.003091f
C41132 a_5807_45002# a_7229_43940# 3.1e-20
C41133 a_n2438_43548# a_n143_45144# 1.67e-20
C41134 a_n743_46660# a_n37_45144# 5.42e-20
C41135 a_4419_46090# a_n2661_45546# 0.019708f
C41136 a_n2293_46634# a_2382_45260# 0.046113f
C41137 a_n881_46662# a_1307_43914# 1.96e-19
C41138 a_n1925_46634# a_327_44734# 2.4e-20
C41139 a_1823_45246# a_n357_42282# 0.031648f
C41140 a_167_45260# a_n1099_45572# 2.69e-19
C41141 a_12891_46348# a_9482_43914# 0.314487f
C41142 a_12549_44172# a_13348_45260# 0.001434f
C41143 a_4190_30871# C4_N_btm 1.36e-19
C41144 a_22400_42852# a_22397_42558# 0.001581f
C41145 a_17486_43762# VDD 4.6e-19
C41146 a_8325_42308# a_8791_42308# 0.173196f
C41147 a_5534_30871# a_8530_39574# 1.75e-19
C41148 a_n1630_35242# a_4958_30871# 0.036823f
C41149 a_n443_42852# a_14456_42282# 7.8e-21
C41150 a_n913_45002# a_21356_42826# 7.3e-21
C41151 a_n2661_44458# a_10695_43548# 9.47e-21
C41152 a_20512_43084# a_20623_43914# 2.29e-20
C41153 a_n356_44636# a_3080_42308# 0.072716f
C41154 a_16721_46634# VDD 0.186443f
C41155 a_16388_46812# RST_Z 3.56e-20
C41156 a_17719_45144# a_17324_43396# 1.66e-20
C41157 a_3232_43370# a_10341_42308# 2.53e-19
C41158 a_16922_45042# a_18783_43370# 1.97e-21
C41159 a_3905_42865# a_n2661_42282# 3.49e-20
C41160 a_22315_44484# a_15493_43940# 6.3e-21
C41161 a_20835_44721# a_14021_43940# 6.15e-21
C41162 a_5263_45724# a_6511_45714# 6.81e-21
C41163 a_5907_45546# a_6472_45840# 0.041762f
C41164 a_2711_45572# a_7227_45028# 0.014767f
C41165 a_13661_43548# a_17517_44484# 0.01824f
C41166 a_9290_44172# a_413_45260# 3.87e-22
C41167 a_3483_46348# a_6709_45028# 0.002873f
C41168 a_768_44030# a_11967_42832# 1.22e-21
C41169 a_12549_44172# a_19615_44636# 0.157395f
C41170 a_19900_46494# a_3357_43084# 7.4e-21
C41171 a_19692_46634# a_21005_45260# 4.64e-19
C41172 a_19466_46812# a_21101_45002# 2.51e-20
C41173 a_13059_46348# a_14976_45348# 0.001245f
C41174 a_15227_44166# a_11827_44484# 0.084637f
C41175 a_6945_45028# a_2437_43646# 2.26888f
C41176 a_5164_46348# a_3232_43370# 5.59e-20
C41177 a_4646_46812# a_n356_44636# 1.8e-20
C41178 a_n2438_43548# a_n2293_43922# 0.575621f
C41179 a_n4209_39304# a_n3565_38216# 0.02945f
C41180 a_5932_42308# C0_N_btm 0.015561f
C41181 a_13381_47204# a_n1435_47204# 0.050056f
C41182 a_n3565_39304# a_n4209_38216# 0.02863f
C41183 a_5934_30871# C4_P_btm 0.030578f
C41184 a_6151_47436# a_16023_47582# 6.16e-20
C41185 a_2063_45854# a_4883_46098# 0.116597f
C41186 a_6123_31319# C2_P_btm 0.01106f
C41187 a_n971_45724# a_n89_47570# 4.31e-19
C41188 a_3823_42558# VDD 0.170296f
C41189 a_n2109_47186# a_3315_47570# 3.55e-19
C41190 a_18114_32519# a_22400_42852# 1.47e-20
C41191 a_3503_45724# VDD 0.129733f
C41192 a_12429_44172# a_10341_43396# 9.54e-20
C41193 a_10807_43548# a_10849_43646# 0.003445f
C41194 a_15493_43396# a_9145_43396# 1.4e-20
C41195 a_14955_43940# a_14955_43396# 0.012141f
C41196 a_9313_44734# a_22223_42860# 0.012144f
C41197 a_n2810_45028# a_n4315_30879# 0.02588f
C41198 en_comp a_22465_38105# 0.533581f
C41199 a_3737_43940# a_3626_43646# 7.51e-19
C41200 a_n4318_39304# a_n2433_43396# 6.19e-19
C41201 a_n2840_43370# a_n2129_43609# 0.001183f
C41202 a_11322_45546# a_9482_43914# 8.92e-20
C41203 a_10903_43370# a_n2661_42834# 0.269313f
C41204 a_13259_45724# a_18545_45144# 2.48e-21
C41205 a_768_44030# a_648_43396# 5.84e-19
C41206 a_n1613_43370# a_6452_43396# 3.31e-19
C41207 a_n971_45724# a_n1853_43023# 0.02483f
C41208 SMPL_ON_P a_n901_43156# 4.04e-21
C41209 a_6977_45572# a_6171_45002# 0.001188f
C41210 a_4185_45028# a_17517_44484# 0.006178f
C41211 a_11415_45002# a_21073_44484# 4.79e-20
C41212 a_12465_44636# a_14205_43396# 8.42e-21
C41213 a_10227_46804# a_14621_43646# 3.58e-19
C41214 a_11823_42460# a_11787_45002# 0.217891f
C41215 a_11962_45724# a_13017_45260# 6.79e-20
C41216 a_12861_44030# a_18429_43548# 3.85e-19
C41217 a_13507_46334# a_10341_43396# 0.030637f
C41218 a_18175_45572# a_19365_45572# 2.56e-19
C41219 a_3090_45724# a_10405_44172# 0.126512f
C41220 a_16375_45002# a_17896_45144# 3.43e-20
C41221 a_22521_39511# VDD 0.910209f
C41222 a_10227_46804# a_17609_46634# 1.17e-19
C41223 a_601_46902# a_1110_47026# 2.6e-19
C41224 a_33_46660# a_479_46660# 2.28e-19
C41225 a_8128_46384# a_8492_46660# 0.002286f
C41226 a_n881_46662# a_10467_46802# 5.33e-19
C41227 a_16327_47482# a_19692_46634# 0.023298f
C41228 a_n743_46660# a_2443_46660# 7.25e-20
C41229 a_2107_46812# a_1983_46706# 0.212212f
C41230 a_5807_45002# a_5907_46634# 0.00171f
C41231 a_768_44030# a_5257_43370# 0.028882f
C41232 a_4791_45118# a_765_45546# 0.052444f
C41233 EN_VIN_BSTR_P C2_P_btm 0.118072f
C41234 a_n1925_46634# a_3177_46902# 0.003436f
C41235 a_n133_46660# a_1799_45572# 3.14e-19
C41236 a_n2438_43548# a_n2661_46098# 0.391488f
C41237 a_10341_43396# a_21855_43396# 0.011519f
C41238 a_n2661_42282# a_n961_42308# 2.77e-19
C41239 a_18783_43370# a_15743_43084# 0.303966f
C41240 a_14955_43396# a_5649_42852# 3.11e-21
C41241 a_3626_43646# a_8387_43230# 3.45e-20
C41242 a_2982_43646# a_8952_43230# 9.76e-21
C41243 a_n97_42460# a_18083_42858# 0.010531f
C41244 a_14180_45002# VDD 0.151315f
C41245 a_5013_44260# a_5267_42460# 1.11e-21
C41246 a_526_44458# a_3353_43940# 0.002743f
C41247 a_13159_45002# a_13490_45067# 2.82e-19
C41248 a_10193_42453# a_20679_44626# 1.62e-21
C41249 a_n745_45366# a_n2661_44458# 9.14e-19
C41250 a_n913_45002# a_n2433_44484# 1.25e-20
C41251 a_n2810_45028# a_n4318_40392# 0.026026f
C41252 a_5257_43370# a_5755_42852# 7.53e-19
C41253 a_n2017_45002# a_n2267_44484# 0.034473f
C41254 a_n1059_45260# a_n2129_44697# 0.032443f
C41255 a_n2956_37592# a_n2840_44458# 1.36e-20
C41256 a_n2661_45010# a_n1352_44484# 0.051998f
C41257 a_n2293_45010# a_n1917_44484# 0.00169f
C41258 en_comp a_19721_31679# 1.48e-19
C41259 a_15227_44166# a_17433_43396# 1.76e-19
C41260 a_4791_45118# a_4921_42308# 0.172224f
C41261 a_14180_45002# a_14309_45348# 0.010132f
C41262 a_13259_45724# a_13483_43940# 0.002807f
C41263 a_3357_43084# a_5343_44458# 0.02588f
C41264 a_8696_44636# a_9241_44734# 4.73e-19
C41265 a_n443_42852# a_895_43940# 6.44e-19
C41266 a_n2661_46634# a_6945_45028# 0.03015f
C41267 a_4955_46873# a_5068_46348# 0.081759f
C41268 a_13507_46334# a_18147_46436# 0.001182f
C41269 a_4817_46660# a_4704_46090# 2.68e-19
C41270 a_n881_46662# a_8034_45724# 0.020183f
C41271 a_17609_46634# a_17339_46660# 0.010277f
C41272 a_16292_46812# a_765_45546# 2.99e-38
C41273 a_n237_47217# a_6511_45714# 3.49e-19
C41274 a_n971_45724# a_6598_45938# 2.89e-20
C41275 a_3877_44458# a_5497_46414# 1.88e-19
C41276 a_4646_46812# a_5204_45822# 1.32e-19
C41277 a_4651_46660# a_5164_46348# 0.002696f
C41278 a_3422_30871# C0_dummy_N_btm 1.28e-20
C41279 a_20922_43172# a_21356_42826# 0.017093f
C41280 a_19987_42826# a_21195_42852# 4.49e-20
C41281 a_n4318_39304# a_n4064_40160# 0.062069f
C41282 a_3626_43646# a_16522_42674# 0.002817f
C41283 a_20679_44626# VDD 0.439119f
C41284 a_8387_43230# a_8649_43218# 0.001705f
C41285 a_8605_42826# a_9061_43230# 4.2e-19
C41286 a_4361_42308# a_20753_42852# 7.12e-19
C41287 a_13887_32519# a_22400_42852# 0.098244f
C41288 a_n2017_45002# a_19478_44306# 1.53e-20
C41289 a_16979_44734# a_18287_44626# 2.91e-20
C41290 a_14539_43914# a_18443_44721# 2.14e-20
C41291 a_1423_45028# a_1414_42308# 0.005518f
C41292 a_626_44172# a_2127_44172# 3.19e-20
C41293 a_375_42282# a_895_43940# 5.29e-20
C41294 a_11827_44484# a_12189_44484# 1.28e-19
C41295 a_5147_45002# a_n2661_42282# 3.8e-19
C41296 a_n357_42282# a_17324_43396# 1.48e-20
C41297 a_n443_42852# a_10149_43396# 8.96e-19
C41298 a_18587_45118# a_17517_44484# 5.57e-20
C41299 a_1307_43914# a_2889_44172# 0.02756f
C41300 a_7499_43078# a_8147_43396# 0.227361f
C41301 a_3232_43370# a_3499_42826# 0.339727f
C41302 a_8270_45546# a_9223_42460# 2.21e-19
C41303 a_17767_44458# a_18248_44752# 0.041822f
C41304 a_13249_42308# a_2982_43646# 1.48e-19
C41305 a_4743_44484# a_6109_44484# 2.06e-20
C41306 a_4223_44672# a_8375_44464# 0.001207f
C41307 a_5518_44484# a_5289_44734# 6.46e-20
C41308 a_526_44458# a_8605_42826# 0.021896f
C41309 a_13259_45724# a_13678_32519# 0.013938f
C41310 a_n1059_45260# a_15493_43396# 0.044794f
C41311 a_11691_44458# a_15463_44811# 7.26e-19
C41312 a_4842_47570# a_3357_43084# 1.16e-19
C41313 a_20990_47178# a_413_45260# 1.26e-19
C41314 a_10227_46804# a_3537_45260# 2.05e-20
C41315 a_13925_46122# a_15015_46420# 0.042415f
C41316 a_13759_46122# a_14840_46494# 0.102325f
C41317 a_14493_46090# a_14275_46494# 0.209641f
C41318 a_2698_46116# a_2981_46116# 0.003683f
C41319 a_2521_46116# a_526_44458# 3.89e-20
C41320 a_19123_46287# a_18051_46116# 8.02e-20
C41321 a_13747_46662# a_19431_45546# 0.02276f
C41322 a_13661_43548# a_19256_45572# 0.00171f
C41323 a_n2312_39304# a_n2017_45002# 9.89e-22
C41324 a_13351_46090# a_2324_44458# 1.29e-20
C41325 a_n971_45724# a_2809_45028# 0.037351f
C41326 a_1176_45822# a_1337_46116# 0.026848f
C41327 a_11813_46116# a_2711_45572# 1.5e-19
C41328 a_n743_46660# a_16223_45938# 1.43e-19
C41329 a_n443_46116# a_1307_43914# 0.442637f
C41330 a_8199_44636# a_6945_45028# 5.83e-20
C41331 a_8016_46348# a_10809_44734# 6.66e-20
C41332 a_22165_42308# a_22465_38105# 1.77e-19
C41333 a_14635_42282# a_14456_42282# 0.172313f
C41334 a_13291_42460# a_13249_42558# 0.002309f
C41335 a_6765_43638# VDD 0.218204f
C41336 a_4190_30871# a_8530_39574# 1.25e-19
C41337 a_1184_42692# a_2351_42308# 4.23e-20
C41338 a_n784_42308# a_3823_42558# 2.06e-20
C41339 a_14097_32519# a_5934_30871# 2.14e-19
C41340 a_n2293_45010# a_n1853_43023# 4.48e-20
C41341 a_n863_45724# a_1755_42282# 0.050501f
C41342 a_2382_45260# a_743_42282# 0.023665f
C41343 a_n357_42282# a_1184_42692# 2.11e-19
C41344 a_n755_45592# a_1576_42282# 0.025747f
C41345 a_7927_46660# VDD 0.187888f
C41346 a_9313_44734# a_20269_44172# 1.88e-20
C41347 a_n2293_43922# a_12429_44172# 0.006182f
C41348 a_n2661_43370# a_8791_43396# 2.79e-21
C41349 a_n746_45260# a_n1761_44111# 2.69e-20
C41350 a_n971_45724# a_n1899_43946# 0.021838f
C41351 a_n2497_47436# a_1414_42308# 0.005579f
C41352 a_4883_46098# a_n2661_42834# 0.019268f
C41353 a_n2293_45546# a_n357_42282# 0.032623f
C41354 a_n2661_45546# a_1848_45724# 0.005986f
C41355 a_13059_46348# a_6171_45002# 0.070496f
C41356 a_20273_46660# a_413_45260# 2.73e-21
C41357 a_20820_30879# a_20447_31679# 0.053904f
C41358 a_11415_45002# a_21542_45572# 5.19e-19
C41359 a_n2293_46634# a_5343_44458# 0.026475f
C41360 a_13661_43548# a_13720_44458# 0.122691f
C41361 a_15227_44166# a_15595_45028# 0.007902f
C41362 a_n863_45724# a_n1099_45572# 0.172847f
C41363 a_n452_45724# a_380_45546# 5.21e-19
C41364 a_8034_45724# a_8162_45546# 0.14162f
C41365 a_5066_45546# a_8746_45002# 1.34e-19
C41366 a_n743_46660# a_949_44458# 3.73e-20
C41367 a_n2438_43548# a_742_44458# 0.171623f
C41368 a_12005_46116# a_8696_44636# 7.73e-21
C41369 a_10428_46928# a_n2661_43370# 2.58e-21
C41370 a_1606_42308# VDAC_N 0.01093f
C41371 a_14097_32519# a_11530_34132# 0.002965f
C41372 a_n4334_40480# a_n4064_40160# 0.43652f
C41373 a_n4315_30879# a_n2302_40160# 0.407166f
C41374 a_5742_30871# a_2113_38308# 6.13e-20
C41375 a_12800_43218# VDD 0.078978f
C41376 a_n2288_47178# a_n1151_42308# 6.07e-19
C41377 a_n746_45260# a_1239_47204# 2.56e-19
C41378 a_n23_47502# a_327_47204# 0.140943f
C41379 a_n2109_47186# a_3160_47472# 0.054333f
C41380 a_n1741_47186# a_2952_47436# 0.010669f
C41381 a_n237_47217# a_1209_47178# 0.206644f
C41382 a_n971_45724# a_1431_47204# 0.030942f
C41383 a_2479_44172# a_2437_43396# 5.86e-20
C41384 a_11967_42832# a_16759_43396# 0.001677f
C41385 a_15493_43940# a_19319_43548# 0.36082f
C41386 a_21115_43940# a_21205_44306# 0.004764f
C41387 a_11173_44260# a_11257_43940# 0.002303f
C41388 a_20623_43914# a_21381_43940# 1.02e-19
C41389 a_11341_43940# a_19478_44056# 2.7e-20
C41390 a_5111_44636# a_5379_42460# 0.118194f
C41391 a_n1059_45260# a_8791_42308# 8.01e-19
C41392 a_n2017_45002# a_9223_42460# 0.003774f
C41393 a_n913_45002# a_8685_42308# 0.007967f
C41394 a_n2661_42282# a_4093_43548# 9.71e-22
C41395 a_6453_43914# a_6293_42852# 0.00419f
C41396 a_5663_43940# a_6197_43396# 1.2e-19
C41397 a_3232_43370# a_3318_42354# 1.69e-19
C41398 a_19862_44208# a_17538_32519# 7.43e-20
C41399 a_20205_31679# a_22821_38993# 5.5e-20
C41400 a_15903_45785# a_15765_45572# 0.205788f
C41401 a_19692_46634# a_20835_44721# 1.53e-19
C41402 a_13507_46334# a_n97_42460# 1.31e-19
C41403 a_2277_45546# a_2382_45260# 0.00187f
C41404 a_n443_42852# a_3065_45002# 0.022494f
C41405 a_1609_45822# a_2680_45002# 1.31e-20
C41406 a_12861_44030# a_2982_43646# 2.08e-20
C41407 a_2063_45854# a_8685_43396# 9.17e-20
C41408 a_768_44030# a_5745_43940# 9.71e-20
C41409 a_8016_46348# a_5883_43914# 2.29e-20
C41410 a_15599_45572# a_16333_45814# 0.053479f
C41411 a_13059_46348# a_14673_44172# 0.108306f
C41412 a_3316_45546# a_3232_43370# 2.28e-19
C41413 a_5937_45572# a_6298_44484# 0.036004f
C41414 a_8199_44636# a_8103_44636# 0.256009f
C41415 a_n901_46420# a_n356_44636# 9.91e-21
C41416 a_1177_38525# VDD 0.373535f
C41417 VDAC_N a_8912_37509# 3.43288f
C41418 a_6886_37412# VDAC_P 0.062773f
C41419 a_6151_47436# a_8492_46660# 0.302615f
C41420 a_7227_47204# a_7577_46660# 5.88e-19
C41421 a_4915_47217# a_10428_46928# 7.56e-19
C41422 a_6575_47204# a_7411_46660# 2.14e-19
C41423 a_n1613_43370# a_n2956_39768# 3.32e-21
C41424 a_12891_46348# a_13747_46662# 6.08e-22
C41425 a_768_44030# a_5807_45002# 0.025167f
C41426 a_12549_44172# a_13661_43548# 0.149087f
C41427 a_5700_37509# a_11206_38545# 4.96e-20
C41428 a_19479_31679# C2_N_btm 0.001057f
C41429 a_19478_44306# a_19164_43230# 4.47e-20
C41430 a_9145_43396# a_10695_43548# 0.053202f
C41431 a_n2661_42834# a_7963_42308# 2.63e-21
C41432 a_n2293_43922# a_7227_42308# 8.6e-20
C41433 a_11341_43940# a_17701_42308# 7.35e-20
C41434 a_n2840_43370# a_n2840_42826# 0.026152f
C41435 a_2982_43646# a_19700_43370# 3.31e-20
C41436 a_8685_43396# a_14955_43396# 0.111211f
C41437 a_n356_44636# a_15764_42576# 0.012586f
C41438 a_3626_43646# a_15743_43084# 2.37e-19
C41439 a_20528_45572# VDD 0.08228f
C41440 a_n2312_38680# a_n4318_38680# 0.023332f
C41441 a_13249_42308# a_14539_43914# 0.032256f
C41442 a_n2956_39304# a_n2661_42282# 5.57e-20
C41443 a_3537_45260# a_1307_43914# 0.290878f
C41444 a_413_45260# a_2304_45348# 9.35e-20
C41445 a_1823_45246# a_5025_43940# 8.65e-20
C41446 a_12741_44636# a_19319_43548# 3.83e-20
C41447 a_6171_45002# a_13556_45296# 0.017156f
C41448 a_1667_45002# a_1423_45028# 0.0017f
C41449 a_n2438_43548# a_n901_43156# 3.58e-21
C41450 a_4883_46098# a_17715_44484# 0.024632f
C41451 a_18479_47436# a_21137_46414# 0.002071f
C41452 a_2063_45854# a_11608_46482# 0.001173f
C41453 a_11453_44696# a_14275_46494# 6.78e-21
C41454 a_13507_46334# a_17957_46116# 0.007078f
C41455 a_19787_47423# a_19335_46494# 0.001054f
C41456 a_17591_47464# a_10809_44734# 0.007346f
C41457 a_18143_47464# a_6945_45028# 0.023139f
C41458 a_n1151_42308# a_10044_46482# 0.001342f
C41459 a_n881_46662# a_8016_46348# 0.024184f
C41460 a_12465_44636# a_15682_46116# 4.04e-20
C41461 a_6755_46942# a_14976_45028# 0.029836f
C41462 a_12549_44172# a_4185_45028# 3.66e-21
C41463 a_6545_47178# a_6640_46482# 9.37e-19
C41464 a_4791_45118# a_6347_46155# 0.005265f
C41465 a_18597_46090# a_19900_46494# 0.039688f
C41466 a_8037_42858# a_8387_43230# 0.225358f
C41467 a_7871_42858# a_8952_43230# 0.102355f
C41468 a_3626_43646# a_1606_42308# 2.02e-20
C41469 a_13887_32519# a_22223_42860# 0.013362f
C41470 a_11341_43940# a_21613_42308# 4e-22
C41471 a_3080_42308# a_3823_42558# 0.016209f
C41472 a_4905_42826# a_3318_42354# 4.93e-21
C41473 a_n1655_44484# VDD 1.27e-19
C41474 a_n97_42460# a_7227_42308# 0.032716f
C41475 a_20749_43396# a_20922_43172# 3.92e-19
C41476 a_n2017_45002# a_n2065_43946# 0.045593f
C41477 a_n2293_45010# a_n1899_43946# 0.18948f
C41478 a_n2661_45010# a_n1549_44318# 2.9e-20
C41479 a_9482_43914# a_16241_44734# 9.38e-20
C41480 a_13556_45296# a_14673_44172# 0.137701f
C41481 a_n2661_44458# a_n2433_44484# 0.039874f
C41482 a_n2840_44458# a_n2267_44484# 4.89e-19
C41483 a_413_45260# a_22315_44484# 1.08e-20
C41484 a_n2312_40392# a_n4315_30879# 0.389397f
C41485 a_2437_43646# a_895_43940# 0.025092f
C41486 a_4185_45028# a_5111_42852# 0.001197f
C41487 a_16922_45042# a_17767_44458# 2.79e-19
C41488 a_n4318_40392# a_n2129_44697# 4.04e-19
C41489 a_8696_44636# a_15682_43940# 0.001466f
C41490 a_n443_42852# a_458_43396# 0.023429f
C41491 a_17023_45118# a_16979_44734# 1.26e-19
C41492 a_4883_46098# a_15861_45028# 3.69e-21
C41493 a_16327_47482# a_18175_45572# 0.346603f
C41494 a_14976_45028# a_8049_45260# 0.025611f
C41495 a_1823_45246# a_3147_46376# 1.55e-20
C41496 a_3785_47178# a_3357_43084# 9.76e-20
C41497 a_n971_45724# en_comp 5.07e-20
C41498 a_4700_47436# a_2437_43646# 0.007905f
C41499 a_584_46384# a_n2661_45010# 0.017317f
C41500 a_n2109_47186# a_413_45260# 0.027314f
C41501 a_n2497_47436# a_1667_45002# 9.11e-20
C41502 a_167_45260# a_2698_46116# 0.019127f
C41503 a_765_45546# a_6945_45028# 4.99804f
C41504 a_5807_45002# a_11652_45724# 7.11e-20
C41505 a_2107_46812# a_6194_45824# 1.15e-20
C41506 a_11599_46634# a_19431_45546# 0.056971f
C41507 a_11453_44696# a_15765_45572# 5.36e-20
C41508 a_5534_30871# a_13575_42558# 0.002235f
C41509 a_14543_43071# a_14456_42282# 0.009977f
C41510 a_5111_44636# a_7287_43370# 0.104641f
C41511 a_20567_45036# a_14021_43940# 3.06e-22
C41512 a_19594_46812# VDD 0.349555f
C41513 a_375_42282# a_458_43396# 0.014454f
C41514 a_19452_47524# START 0.003297f
C41515 a_5883_43914# a_7584_44260# 1.86e-20
C41516 a_3537_45260# a_9396_43370# 5.47e-19
C41517 a_19321_45002# RST_Z 1.28e-19
C41518 a_10193_42453# a_10341_42308# 0.061874f
C41519 a_3232_43370# a_6197_43396# 6.79e-20
C41520 a_n357_42282# a_5193_42852# 0.00356f
C41521 a_1307_43914# a_1049_43396# 0.001373f
C41522 a_21588_30879# C8_N_btm 0.002806f
C41523 a_17517_44484# a_11967_42832# 0.342031f
C41524 a_9290_44172# a_11323_42473# 0.006277f
C41525 a_11599_46634# a_13076_44458# 8.18e-23
C41526 a_13661_43548# a_15685_45394# 4.18e-20
C41527 SMPL_ON_P a_n2661_43922# 0.002089f
C41528 a_19692_46634# a_20731_45938# 3.6e-19
C41529 a_15682_46116# a_2711_45572# 0.001308f
C41530 a_n1925_42282# a_n863_45724# 1.17e-19
C41531 a_n1925_46634# a_n2293_42834# 0.004172f
C41532 a_7577_46660# a_6171_45002# 3.93e-21
C41533 a_3090_45724# a_3357_43084# 0.546562f
C41534 a_n2312_40392# a_n4318_40392# 0.025284f
C41535 a_12861_44030# a_14539_43914# 0.02276f
C41536 a_12549_44172# a_18587_45118# 5.24e-21
C41537 a_5937_45572# a_5437_45600# 3.8e-19
C41538 a_8016_46348# a_8162_45546# 0.001995f
C41539 a_5342_30871# C1_N_btm 9.04e-20
C41540 a_n4318_38216# a_n4064_37984# 0.017009f
C41541 a_5534_30871# C3_N_btm 7.69e-20
C41542 a_15890_42674# a_17303_42282# 1.66e-20
C41543 a_n4318_37592# a_n3565_38216# 5.63e-19
C41544 a_n3674_38216# a_n3420_37984# 0.064303f
C41545 a_11551_42558# a_7174_31319# 4.88e-21
C41546 a_10341_42308# VDD 0.931019f
C41547 a_18287_44626# a_18429_43548# 8.45e-21
C41548 a_n2810_45572# a_n2302_38778# 0.001992f
C41549 a_n1059_45260# a_18707_42852# 8.57e-19
C41550 a_n2017_45002# a_20256_43172# 3.49e-19
C41551 a_n2840_43914# a_n4318_39304# 0.002229f
C41552 a_9313_44734# a_14358_43442# 5.8e-20
C41553 a_10193_42453# a_18057_42282# 0.099046f
C41554 a_n2956_38216# a_n3420_38528# 8.07e-19
C41555 a_18451_43940# a_19328_44172# 0.008311f
C41556 a_18326_43940# a_15493_43396# 3.68e-20
C41557 a_18079_43940# a_19478_44306# 2.26e-20
C41558 a_5164_46348# VDD 0.717083f
C41559 a_9672_43914# a_9801_44260# 0.010132f
C41560 a_11750_44172# a_11341_43940# 0.002015f
C41561 a_n2661_42834# a_8685_43396# 9.54e-20
C41562 a_5343_44458# a_743_42282# 0.010119f
C41563 a_5066_45546# a_3232_43370# 0.00301f
C41564 a_7920_46348# a_n2661_43370# 1.68e-20
C41565 a_5937_45572# a_7418_45067# 9.73e-20
C41566 a_3483_46348# a_13807_45067# 2.62e-19
C41567 a_11823_42460# a_13904_45546# 0.067334f
C41568 a_7499_43078# a_10907_45822# 5.14e-19
C41569 a_9049_44484# a_10210_45822# 1.6e-20
C41570 a_n2438_43548# a_n984_44318# 2.41e-21
C41571 a_12741_44636# a_17801_45144# 3.91e-19
C41572 a_13059_46348# a_12607_44458# 0.033056f
C41573 a_6755_46942# a_15433_44458# 0.006016f
C41574 a_8034_45724# a_3537_45260# 1.54e-20
C41575 a_526_44458# a_8953_45002# 1.35e-19
C41576 a_n971_45724# a_n1699_43638# 0.001253f
C41577 a_n2497_47436# a_n1190_43762# 4.44e-19
C41578 a_n2109_47186# a_2609_46660# 5.01e-20
C41579 a_4700_47436# a_n2661_46634# 1.58e-20
C41580 a_9067_47204# a_5807_45002# 7.49e-20
C41581 a_n1435_47204# a_13675_47204# 0.012767f
C41582 a_13381_47204# a_13759_47204# 8.62e-21
C41583 a_7174_31319# C0_dummy_N_btm 0.029132f
C41584 a_11599_46634# a_12891_46348# 0.150715f
C41585 a_14955_47212# a_12549_44172# 7.05e-20
C41586 a_n3420_39616# a_n923_35174# 0.002953f
C41587 a_n1741_47186# a_n2661_46098# 3.12e-19
C41588 a_n746_45260# a_491_47026# 0.002692f
C41589 a_11453_44696# a_22959_47212# 0.182671f
C41590 a_13258_32519# C2_N_btm 2.75e-19
C41591 a_n4315_30879# C9_P_btm 0.003123f
C41592 a_14311_47204# a_768_44030# 0.033509f
C41593 a_18057_42282# VDD 0.130308f
C41594 a_n4209_38216# a_n3690_37440# 5.18e-19
C41595 a_n3565_38216# a_n4334_37440# 6.61e-19
C41596 a_3160_47472# a_n1925_46634# 0.026425f
C41597 a_n1151_42308# a_n2312_38680# 6.25e-20
C41598 a_584_46384# a_171_46873# 0.007683f
C41599 a_1209_47178# a_1123_46634# 0.001301f
C41600 a_17531_42308# RST_Z 1.65e-20
C41601 a_14021_43940# a_17486_43762# 1.72e-19
C41602 a_n2661_42282# a_685_42968# 1.62e-20
C41603 a_18494_42460# a_15803_42450# 1.58e-20
C41604 a_1427_43646# a_1512_43396# 1.48e-19
C41605 a_3626_43646# a_3539_42460# 0.017877f
C41606 a_11341_43940# a_4361_42308# 0.001978f
C41607 a_11823_42460# CLK 3.11e-20
C41608 a_4905_42826# a_6197_43396# 1.53e-20
C41609 a_8336_45822# VDD 0.004437f
C41610 a_9313_44734# a_20836_43172# 9.15e-20
C41611 a_3499_42826# a_2905_42968# 0.00265f
C41612 a_n443_42852# a_6298_44484# 2.15e-20
C41613 a_14976_45028# a_15037_43940# 3.42e-20
C41614 a_8049_45260# a_15433_44458# 4.08e-21
C41615 a_4646_46812# a_6765_43638# 0.043651f
C41616 a_12741_44636# a_10949_43914# 7.98e-20
C41617 a_22959_45572# a_413_45260# 0.021231f
C41618 a_n2293_45010# en_comp 0.066194f
C41619 a_n2109_45247# a_n2956_37592# 3.33e-19
C41620 a_13661_43548# a_16977_43638# 1.71e-20
C41621 a_11415_45002# a_12429_44172# 1.15e-21
C41622 a_n1059_45260# a_n745_45366# 0.0613f
C41623 a_n2017_45002# a_n2810_45028# 1.6e-19
C41624 a_5164_46348# a_5495_43940# 9.57e-20
C41625 a_16147_45260# a_14797_45144# 1.1e-19
C41626 a_10193_42453# a_18494_42460# 0.074751f
C41627 a_13249_42308# a_14309_45028# 0.008249f
C41628 a_13059_46348# a_14761_44260# 8.03e-20
C41629 a_n971_45724# a_2324_44458# 0.021839f
C41630 a_5807_45002# a_10933_46660# 0.001833f
C41631 a_768_44030# a_14226_46987# 5.35e-19
C41632 a_12549_44172# a_14543_46987# 3.29e-19
C41633 a_n1435_47204# a_167_45260# 1.15e-20
C41634 a_20894_47436# a_12741_44636# 4.32e-20
C41635 a_5167_46660# a_5257_43370# 6.3e-20
C41636 a_n1151_42308# a_9823_46155# 0.061688f
C41637 a_n2293_46634# a_3090_45724# 1.2853f
C41638 a_3411_47243# a_765_45546# 2.63e-19
C41639 a_11453_44696# a_18280_46660# 0.005332f
C41640 a_13507_46334# a_11415_45002# 0.160889f
C41641 a_21496_47436# a_20202_43084# 0.00124f
C41642 a_20843_47204# a_19692_46634# 4.52e-20
C41643 a_n743_46660# a_12991_46634# 1.55e-20
C41644 a_2063_45854# a_11387_46155# 0.079443f
C41645 a_4646_46812# a_7927_46660# 7.75e-20
C41646 a_21381_43940# a_14097_32519# 1.99e-20
C41647 a_14401_32519# a_22400_42852# 8.97e-20
C41648 a_18494_42460# VDD 0.73193f
C41649 a_18184_42460# RST_Z 0.001648f
C41650 a_10341_43396# a_17701_42308# 2.12e-19
C41651 a_10807_43548# a_11323_42473# 0.109765f
C41652 a_20202_43084# a_13678_32519# 0.027425f
C41653 a_20820_30879# a_13467_32519# 0.053319f
C41654 a_n2956_39768# a_n1736_42282# 3.63e-20
C41655 a_n755_45592# a_1241_43940# 3.29e-21
C41656 a_n2312_38680# a_n2840_42282# 2.73e-20
C41657 a_n2442_46660# a_n4318_38216# 0.023718f
C41658 a_13348_45260# a_13076_44458# 4.88e-20
C41659 a_1307_43914# a_8701_44490# 7.15e-21
C41660 a_9482_43914# a_12883_44458# 7.92e-20
C41661 a_13556_45296# a_12607_44458# 0.01896f
C41662 a_526_44458# a_3626_43646# 0.022127f
C41663 a_3065_45002# a_4181_44734# 3.66e-20
C41664 a_7499_43078# a_n2661_42282# 5.53e-21
C41665 a_1423_45028# a_n699_43396# 0.008455f
C41666 a_2711_45572# a_20269_44172# 8.26e-19
C41667 a_22612_30879# COMP_P 3.57e-19
C41668 a_3090_45724# a_5342_30871# 0.001809f
C41669 a_11901_46660# a_10903_43370# 5.8e-19
C41670 a_11813_46116# a_12005_46116# 0.038046f
C41671 a_12861_44030# a_12427_45724# 0.002445f
C41672 a_13717_47436# a_11823_42460# 1.19e-20
C41673 a_4651_46660# a_5066_45546# 4.76e-19
C41674 a_768_44030# a_n755_45592# 0.202175f
C41675 a_20411_46873# a_12741_44636# 0.095741f
C41676 a_20273_46660# a_20820_30879# 2.63e-19
C41677 a_11599_46634# a_11322_45546# 1.09e-19
C41678 a_20528_46660# a_20719_46660# 4.61e-19
C41679 a_21188_46660# a_22365_46825# 2e-20
C41680 a_n1613_43370# a_n906_45572# 2.51e-19
C41681 a_21363_46634# a_20202_43084# 0.048242f
C41682 a_13381_47204# a_13163_45724# 4.49e-21
C41683 a_11735_46660# a_12594_46348# 1.94e-19
C41684 a_10428_46928# a_10809_44734# 1.88e-19
C41685 a_16409_43396# a_4958_30871# 5.65e-20
C41686 a_4361_42308# a_10723_42308# 0.010334f
C41687 a_743_42282# a_12563_42308# 0.00803f
C41688 a_16137_43396# a_18057_42282# 0.01884f
C41689 a_19164_43230# a_20256_43172# 1.29e-19
C41690 a_3499_42826# VDD 0.333472f
C41691 a_10341_42308# a_n784_42308# 1.87e-21
C41692 a_3080_42308# a_1177_38525# 2.16e-19
C41693 a_10341_43396# a_21613_42308# 2.29e-20
C41694 a_n357_42282# a_7227_42852# 0.185359f
C41695 a_n755_45592# a_5755_42852# 6.41e-21
C41696 a_14180_45002# a_14021_43940# 2.49e-20
C41697 a_13720_44458# a_11967_42832# 1.06e-21
C41698 a_16979_44734# a_17061_44484# 0.003935f
C41699 a_14539_43914# a_17325_44484# 2.02e-20
C41700 a_13259_45724# a_18083_42858# 0.002348f
C41701 a_15673_47210# VDD 0.569224f
C41702 a_526_44458# a_8649_43218# 0.002066f
C41703 a_n1435_47204# DATA[4] 0.033859f
C41704 a_15811_47375# RST_Z 1.42e-19
C41705 a_n2661_44458# a_n2840_43914# 0.002411f
C41706 a_n1059_45260# a_n2433_43396# 3.64e-21
C41707 a_n2017_45002# a_n2129_43609# 0.024338f
C41708 a_8333_44734# a_n2661_43922# 1.54e-35
C41709 a_18374_44850# a_18204_44850# 2.6e-19
C41710 a_9313_44734# a_10617_44484# 0.006463f
C41711 a_9241_44734# a_9159_44484# 5.37e-19
C41712 a_18989_43940# a_17517_44484# 0.021791f
C41713 a_3232_43370# a_8415_44056# 1.41e-19
C41714 a_9313_45822# CLK 0.027301f
C41715 a_19900_46494# a_8049_45260# 0.005334f
C41716 a_1208_46090# a_997_45618# 6.64e-20
C41717 a_1176_45822# a_n755_45592# 0.091892f
C41718 a_1138_42852# a_n357_42282# 0.325445f
C41719 a_14035_46660# a_11823_42460# 0.003215f
C41720 a_14275_46494# a_14180_46482# 0.049827f
C41721 a_14493_46090# a_14371_46494# 3.16e-19
C41722 a_n746_45260# a_n2267_44484# 0.003717f
C41723 a_5807_45002# a_7276_45260# 1.33e-20
C41724 a_n743_46660# a_n143_45144# 0.00133f
C41725 a_4185_45028# a_n2661_45546# 0.047991f
C41726 a_n2661_46634# a_3065_45002# 3.58e-21
C41727 a_n2293_46634# a_2274_45254# 0.018017f
C41728 a_n881_46662# a_16019_45002# 5.4e-20
C41729 a_n1613_43370# a_1307_43914# 0.056988f
C41730 a_4915_47217# a_11827_44484# 0.002572f
C41731 a_n1925_46634# a_413_45260# 0.02974f
C41732 a_n1853_46287# a_7_45899# 1.33e-19
C41733 a_167_45260# a_380_45546# 6.63e-19
C41734 a_n2497_47436# a_n699_43396# 0.355158f
C41735 a_768_44030# a_13017_45260# 0.031385f
C41736 a_12891_46348# a_13348_45260# 0.097519f
C41737 a_12549_44172# a_13159_45002# 4.23e-20
C41738 a_13351_46090# a_12839_46116# 7.06e-19
C41739 a_2981_46116# a_526_44458# 0.077706f
C41740 a_5934_30871# a_9377_42558# 0.001873f
C41741 a_4190_30871# C3_N_btm 1.1e-19
C41742 a_8325_42308# a_8685_42308# 0.141819f
C41743 a_5534_30871# a_7754_38470# 1.19e-19
C41744 a_n443_42852# a_13575_42558# 2.2e-21
C41745 a_n913_45002# a_20922_43172# 0.010679f
C41746 a_n2017_45002# a_21195_42852# 8.32e-21
C41747 a_5883_43914# a_8791_43396# 1.82e-19
C41748 a_n2661_44458# a_9803_43646# 6.14e-21
C41749 a_13259_45724# a_22775_42308# 0.007982f
C41750 a_20512_43084# a_20365_43914# 1.4e-19
C41751 a_n356_44636# a_4699_43561# 2.33e-21
C41752 a_16388_46812# VDD 0.797417f
C41753 a_6298_44484# a_6655_43762# 5.21e-20
C41754 a_13059_46348# RST_Z 0.002761f
C41755 a_17613_45144# a_17324_43396# 4.37e-19
C41756 a_17719_45144# a_17499_43370# 2.73e-21
C41757 a_18494_42460# a_16137_43396# 0.115144f
C41758 a_22315_44484# a_22223_43948# 0.012307f
C41759 a_3422_30871# a_15493_43940# 0.014587f
C41760 a_20679_44626# a_14021_43940# 2.62e-20
C41761 en_comp a_18599_43230# 9.77e-22
C41762 a_5907_45546# a_6194_45824# 0.233657f
C41763 a_2711_45572# a_6598_45938# 0.011792f
C41764 a_n2293_46634# a_14815_43914# 0.057388f
C41765 a_5807_45002# a_17517_44484# 1.9e-19
C41766 a_5204_45822# a_4927_45028# 4.9e-19
C41767 a_5497_46414# a_5111_44636# 3.91e-19
C41768 a_3483_46348# a_7229_43940# 0.03702f
C41769 a_12549_44172# a_11967_42832# 0.193926f
C41770 a_19692_46634# a_20567_45036# 5.15e-19
C41771 a_20075_46420# a_3357_43084# 4.81e-21
C41772 a_15368_46634# a_11691_44458# 0.002402f
C41773 a_6945_45028# a_21513_45002# 1.8e-20
C41774 a_21137_46414# a_2437_43646# 3.15e-23
C41775 a_8016_46348# a_3537_45260# 5.67e-20
C41776 a_5164_46348# a_5691_45260# 0.00167f
C41777 a_n2293_46098# a_1307_43914# 0.107603f
C41778 a_n2438_43548# a_n2661_43922# 0.06887f
C41779 a_5932_42308# C0_dummy_N_btm 1.2e-19
C41780 a_11459_47204# a_n1435_47204# 0.001005f
C41781 a_7174_31319# VDAC_Ni 4.91e-19
C41782 a_5934_30871# C5_P_btm 0.139996f
C41783 a_6151_47436# a_16327_47482# 3.69e-20
C41784 a_6123_31319# C3_P_btm 0.011333f
C41785 a_3318_42354# VDD 0.203036f
C41786 a_n2109_47186# a_3094_47570# 6.18e-19
C41787 a_453_43940# a_743_42282# 8.67e-23
C41788 a_n755_45592# DATA[0] 1.08e-20
C41789 a_3316_45546# VDD 0.428912f
C41790 a_11750_44172# a_10341_43396# 2.18e-21
C41791 a_10807_43548# a_10765_43646# 9.53e-19
C41792 a_14955_43940# a_15095_43370# 1.49e-19
C41793 a_9313_44734# a_22165_42308# 0.028818f
C41794 a_n2840_43370# a_n2433_43396# 0.039807f
C41795 a_11322_45546# a_13348_45260# 4.97e-20
C41796 a_13259_45724# a_18450_45144# 3.75e-19
C41797 a_n971_45724# a_n2157_42858# 2.88e-19
C41798 a_8049_45260# a_5343_44458# 3.51e-20
C41799 a_6905_45572# a_6171_45002# 5.84e-19
C41800 a_11415_45002# a_20637_44484# 2.19e-20
C41801 a_12465_44636# a_14358_43442# 3.52e-20
C41802 a_10227_46804# a_14537_43646# 2.7e-19
C41803 a_18479_45785# a_20528_45572# 7.66e-21
C41804 a_17568_45572# a_17668_45572# 0.005294f
C41805 a_19256_45572# a_20273_45572# 1.1e-19
C41806 a_3090_45724# a_9672_43914# 0.004104f
C41807 a_2324_44458# a_9313_44734# 0.001086f
C41808 a_11652_45724# a_13017_45260# 8.37e-21
C41809 a_11823_42460# a_10951_45334# 8.18e-20
C41810 a_11962_45724# a_11963_45334# 0.006674f
C41811 a_n743_46660# a_n2661_46098# 0.414618f
C41812 a_n1925_46634# a_2609_46660# 0.009041f
C41813 a_n2438_43548# a_1799_45572# 0.137623f
C41814 a_22780_40081# VDD 2.4e-19
C41815 a_4883_46098# a_11901_46660# 2.38e-19
C41816 a_10227_46804# a_16292_46812# 3.76e-20
C41817 a_17591_47464# a_17609_46634# 0.014668f
C41818 a_383_46660# a_491_47026# 0.057222f
C41819 a_33_46660# a_1110_47026# 1.46e-19
C41820 a_n2661_46634# a_3067_47026# 0.003055f
C41821 a_8128_46384# a_8667_46634# 0.001141f
C41822 a_n881_46662# a_10428_46928# 0.004039f
C41823 a_16327_47482# a_19466_46812# 0.203994f
C41824 a_948_46660# a_1983_46706# 3.51e-19
C41825 a_5807_45002# a_5167_46660# 3.94e-19
C41826 a_18597_46090# a_3090_45724# 4.27e-20
C41827 EN_VIN_BSTR_P C3_P_btm 0.100325f
C41828 a_4915_47217# a_14447_46660# 3.78e-19
C41829 a_4700_47436# a_765_45546# 0.004317f
C41830 a_n97_42460# a_17701_42308# 0.001768f
C41831 a_20974_43370# a_22165_42308# 8.68e-20
C41832 a_14401_32519# a_22223_42860# 8.04e-20
C41833 a_5244_44056# a_5267_42460# 1.4e-21
C41834 a_3905_42865# a_5379_42460# 1.34e-20
C41835 a_n2661_42282# a_n1329_42308# 2.6e-19
C41836 a_16759_43396# a_16867_43762# 0.057222f
C41837 a_16137_43396# a_15940_43402# 4.65e-19
C41838 a_13777_45326# VDD 0.145151f
C41839 a_3499_42826# a_n784_42308# 4.32e-21
C41840 a_18525_43370# a_15743_43084# 0.058072f
C41841 a_10341_43396# a_4361_42308# 0.027045f
C41842 a_2982_43646# a_9127_43156# 2.28e-19
C41843 a_3626_43646# a_8605_42826# 2.77e-20
C41844 a_3422_30871# a_5742_30871# 0.029732f
C41845 a_n2293_45546# a_n1441_43940# 1.11e-19
C41846 a_n913_45002# a_n2661_44458# 0.024357f
C41847 a_n1059_45260# a_n2433_44484# 3e-21
C41848 a_5257_43370# a_5111_42852# 0.013892f
C41849 a_n2109_45247# a_n2267_44484# 3.19e-19
C41850 a_n2017_45002# a_n2129_44697# 0.033299f
C41851 a_n2661_45010# a_n1177_44458# 0.052759f
C41852 a_n2293_45010# a_n1699_44726# 0.005129f
C41853 en_comp a_18114_32519# 1.07e-19
C41854 a_3090_45724# a_743_42282# 1.62e-19
C41855 a_15227_44166# a_16823_43084# 0.022136f
C41856 a_4791_45118# a_4933_42558# 0.001758f
C41857 a_n2810_45028# a_n2840_44458# 4.31e-19
C41858 a_3357_43084# a_4743_44484# 2.98e-20
C41859 a_17668_45572# a_17767_44458# 7.33e-21
C41860 a_8696_44636# a_8855_44734# 2.74e-19
C41861 a_n443_42852# a_2479_44172# 0.035023f
C41862 w_1575_34946# a_n4064_40160# 9.7e-19
C41863 a_n237_47217# a_6472_45840# 4e-19
C41864 a_n971_45724# a_6667_45809# 9.13e-19
C41865 a_3877_44458# a_5204_45822# 3.25e-19
C41866 a_4651_46660# a_5068_46348# 8.9e-19
C41867 a_4646_46812# a_5164_46348# 6.79e-20
C41868 a_4883_46098# a_15194_46482# 1.02e-19
C41869 a_22612_30879# a_10809_44734# 7.79e-20
C41870 a_13507_46334# a_13259_45724# 0.023413f
C41871 a_n743_46660# a_17957_46116# 1.41e-19
C41872 a_4955_46873# a_4704_46090# 0.109136f
C41873 a_12465_44636# a_14537_46482# 5.66e-19
C41874 a_3090_45724# a_19123_46287# 2.83e-19
C41875 a_16292_46812# a_17339_46660# 1.37e-19
C41876 a_3422_30871# C0_dummy_P_btm 1.28e-20
C41877 a_19164_43230# a_21195_42852# 3.2e-21
C41878 a_2982_43646# a_17124_42282# 3.02e-19
C41879 a_20640_44752# VDD 0.246486f
C41880 a_7871_42858# a_8495_42852# 9.73e-19
C41881 a_8605_42826# a_8649_43218# 3.69e-19
C41882 a_8037_42858# a_9061_43230# 2.36e-20
C41883 a_13467_32519# a_20753_42852# 1.97e-19
C41884 a_22223_43396# a_22400_42852# 4.88e-19
C41885 a_5649_42852# a_14097_32519# 1.23e-20
C41886 a_n4318_39304# a_n4334_40480# 3.36e-19
C41887 a_14539_43914# a_18287_44626# 3.64e-20
C41888 a_4223_44672# a_7640_43914# 0.002847f
C41889 a_626_44172# a_453_43940# 0.163589f
C41890 a_11827_44484# a_11909_44484# 0.00995f
C41891 a_5147_45002# a_6101_44260# 3.6e-20
C41892 a_n357_42282# a_17499_43370# 1.53e-19
C41893 a_2711_45572# a_14358_43442# 1.67e-21
C41894 a_n443_42852# a_9885_43396# 0.001051f
C41895 a_n2312_38680# a_n2302_39866# 1.63e-19
C41896 a_n2661_44458# a_556_44484# 1.56e-19
C41897 a_1307_43914# a_2675_43914# 0.453622f
C41898 a_7499_43078# a_7112_43396# 0.012965f
C41899 a_3090_45724# a_5755_42308# 1.13e-20
C41900 a_526_44458# a_8037_42858# 0.01672f
C41901 a_n2017_45002# a_15493_43396# 6.52e-20
C41902 a_11691_44458# a_15146_44811# 0.002578f
C41903 a_5518_44484# a_5205_44734# 3.77e-20
C41904 a_17767_44458# a_17970_44736# 0.233657f
C41905 a_n1151_42308# a_1423_45028# 1.11e-19
C41906 a_11415_45002# a_10586_45546# 9.19e-19
C41907 a_11453_44696# a_n913_45002# 1.71e-20
C41908 a_20894_47436# a_413_45260# 8.97e-20
C41909 a_13759_46122# a_15015_46420# 0.043475f
C41910 a_13925_46122# a_14275_46494# 0.20669f
C41911 a_167_45260# a_526_44458# 0.003875f
C41912 a_8270_45546# a_6472_45840# 1.23e-19
C41913 a_3090_45724# a_2277_45546# 4.31e-19
C41914 a_19321_45002# a_18341_45572# 0.001456f
C41915 a_18285_46348# a_18051_46116# 0.028958f
C41916 a_13747_46662# a_18691_45572# 0.030666f
C41917 a_5807_45002# a_19256_45572# 0.015716f
C41918 a_13661_43548# a_19431_45546# 4.64e-19
C41919 a_12549_44172# a_20273_45572# 1.54e-20
C41920 a_n2312_40392# a_n2017_45002# 1.3e-21
C41921 a_12594_46348# a_2324_44458# 0.001717f
C41922 a_1208_46090# a_1337_46116# 0.062574f
C41923 a_1176_45822# a_835_46155# 3.09e-19
C41924 a_11735_46660# a_2711_45572# 1.14e-19
C41925 a_4791_45118# a_1307_43914# 0.027544f
C41926 a_1184_42692# a_2123_42473# 0.107417f
C41927 a_961_42354# a_1755_42282# 3.85e-19
C41928 a_22165_42308# a_22397_42558# 8.87e-19
C41929 a_13291_42460# a_14456_42282# 0.015899f
C41930 a_14635_42282# a_13575_42558# 5.53e-19
C41931 a_4190_30871# a_7754_38470# 8.52e-20
C41932 a_n784_42308# a_3318_42354# 1.96e-20
C41933 a_6197_43396# VDD 0.408793f
C41934 a_n2293_45010# a_n2157_42858# 3.31e-20
C41935 a_n2661_45010# a_n1991_42858# 6.37e-20
C41936 a_n863_45724# a_1606_42308# 0.20593f
C41937 a_9313_44734# a_19862_44208# 0.024263f
C41938 a_n357_42282# a_1576_42282# 1.92e-19
C41939 a_8145_46902# VDD 0.199702f
C41940 en_comp a_13887_32519# 8.37e-20
C41941 a_n755_45592# a_1067_42314# 0.047422f
C41942 a_n2661_43922# a_12429_44172# 0.004259f
C41943 a_n2661_45546# a_997_45618# 0.008847f
C41944 a_n2472_45546# a_n755_45592# 6.82e-21
C41945 a_n743_46660# a_742_44458# 3.66e-22
C41946 a_2107_46812# a_n2661_44458# 0.02628f
C41947 a_10903_43370# a_8696_44636# 0.031601f
C41948 a_n2497_47436# a_1467_44172# 0.046456f
C41949 a_n746_45260# a_n2065_43946# 2.94e-21
C41950 a_n971_45724# a_n1761_44111# 0.084835f
C41951 a_n1613_43370# a_n998_44484# 0.002879f
C41952 a_12549_44172# a_18989_43940# 0.016062f
C41953 a_20411_46873# a_413_45260# 1.63e-20
C41954 a_20202_43084# a_21542_45572# 7.05e-19
C41955 a_n1079_45724# a_n1099_45572# 0.15766f
C41956 a_n2293_45546# a_310_45028# 0.113595f
C41957 a_n2293_46634# a_4743_44484# 2.4e-20
C41958 a_5807_45002# a_13720_44458# 0.001051f
C41959 a_2324_44458# a_15037_45618# 1.52e-19
C41960 a_15227_44166# a_15415_45028# 0.222342f
C41961 a_n863_45724# a_380_45546# 4.95e-19
C41962 a_11415_45002# a_21297_45572# 2.47e-19
C41963 a_12741_44636# a_19963_31679# 2.28e-21
C41964 a_n4315_30879# a_n4064_40160# 0.363059f
C41965 a_5932_42308# VDAC_Ni 5.53e-19
C41966 a_10752_42852# VDD 4.6e-19
C41967 a_n2497_47436# a_n1151_42308# 0.156942f
C41968 a_n23_47502# a_n785_47204# 0.031198f
C41969 a_n237_47217# a_327_47204# 0.027301f
C41970 a_n971_45724# a_1239_47204# 0.022077f
C41971 a_n1741_47186# a_2553_47502# 0.010566f
C41972 a_n2109_47186# a_2905_45572# 0.124881f
C41973 a_n746_45260# a_1209_47178# 1.64e-19
C41974 a_3065_45002# a_4921_42308# 4.26e-19
C41975 a_11967_42832# a_16977_43638# 0.001333f
C41976 a_n2293_43922# a_4361_42308# 0.035634f
C41977 a_n356_44636# a_1847_42826# 3.12e-20
C41978 a_11173_44260# a_11173_43940# 8.81e-19
C41979 a_11341_43940# a_18533_43940# 0.005886f
C41980 a_20365_43914# a_21381_43940# 3.94e-20
C41981 a_5111_44636# a_5267_42460# 0.047489f
C41982 a_n1059_45260# a_8685_42308# 5.76e-19
C41983 a_n913_45002# a_8325_42308# 0.233489f
C41984 a_n2017_45002# a_8791_42308# 0.004421f
C41985 a_5066_45546# VDD 1.34058f
C41986 a_3499_42826# a_3080_42308# 4.95e-19
C41987 a_5663_43940# a_6293_42852# 7.17e-19
C41988 a_6453_43914# a_6031_43396# 0.001451f
C41989 a_1414_42308# a_3457_43396# 0.094207f
C41990 a_10057_43914# a_10341_42308# 2.07e-20
C41991 a_3537_45260# a_3905_42558# 1.27e-20
C41992 a_19862_44208# a_20974_43370# 0.026213f
C41993 a_20692_30879# a_22521_39511# 5.01e-20
C41994 a_8199_44636# a_6298_44484# 0.002319f
C41995 a_10809_44734# a_11827_44484# 0.029958f
C41996 a_2711_45572# en_comp 4.72e-20
C41997 a_15599_45572# a_15765_45572# 0.576512f
C41998 a_19692_46634# a_20679_44626# 0.010957f
C41999 a_8049_45260# a_8560_45348# 8.56e-19
C42000 a_5937_45572# a_5518_44484# 4.36e-19
C42001 a_8953_45546# a_5343_44458# 0.002817f
C42002 a_2277_45546# a_2274_45254# 0.011988f
C42003 a_1609_45822# a_2382_45260# 0.001939f
C42004 a_15227_44166# a_19279_43940# 1.77e-21
C42005 a_13661_43548# a_15301_44260# 4.13e-19
C42006 a_19900_46494# a_20193_45348# 8.77e-21
C42007 a_3483_46348# a_15004_44636# 1.48e-20
C42008 a_3877_44458# a_3820_44260# 4.75e-19
C42009 a_13059_46348# a_14581_44484# 7.41e-20
C42010 a_n357_42282# a_7229_43940# 1.8e-20
C42011 a_n2216_38778# VDD 0.004173f
C42012 a_n1741_47186# a_12251_46660# 0.011505f
C42013 a_2063_45854# a_8035_47026# 0.004006f
C42014 a_n237_47217# a_8846_46660# 7.11e-19
C42015 a_2747_46873# a_n2438_43548# 8.92e-19
C42016 a_6886_37412# a_8912_37509# 0.339465f
C42017 a_4915_47217# a_10150_46912# 9.74e-20
C42018 a_6151_47436# a_8667_46634# 0.357581f
C42019 a_7227_47204# a_7715_46873# 3.86e-19
C42020 a_6575_47204# a_5257_43370# 1.06e-19
C42021 a_7903_47542# a_7411_46660# 0.001091f
C42022 a_12891_46348# a_13661_43548# 0.001729f
C42023 a_12549_44172# a_5807_45002# 0.675558f
C42024 a_5088_37509# a_11206_38545# 0.005271f
C42025 a_4338_37500# CAL_N 0.052373f
C42026 a_5700_37509# VDAC_P 0.081094f
C42027 a_19479_31679# C1_N_btm 0.043983f
C42028 a_19478_44306# a_19339_43156# 1.67e-19
C42029 a_n2661_42834# a_6123_31319# 3.51e-21
C42030 a_n2293_43922# a_6761_42308# 4.97e-20
C42031 a_5891_43370# a_10723_42308# 2.6e-20
C42032 a_15493_43940# a_16414_43172# 3.51e-21
C42033 a_11341_43940# a_17595_43084# 3.11e-20
C42034 a_9145_43396# a_9803_43646# 0.055143f
C42035 a_8685_43396# a_15095_43370# 0.064911f
C42036 a_n356_44636# a_15486_42560# 1.56e-19
C42037 a_n4318_40392# a_n4064_40160# 0.077948f
C42038 a_15493_43396# a_19164_43230# 8.79e-19
C42039 a_14539_43914# a_17124_42282# 3.94e-20
C42040 a_3626_43646# a_18783_43370# 6.43e-21
C42041 a_2982_43646# a_19268_43646# 3.9e-21
C42042 a_n97_42460# a_4361_42308# 0.15989f
C42043 a_21188_45572# VDD 0.288663f
C42044 a_n2312_38680# a_n3674_39304# 0.023501f
C42045 a_18691_45572# a_18911_45144# 0.006432f
C42046 a_18479_45785# a_18494_42460# 3.74e-20
C42047 a_768_44030# a_10083_42826# 3.74e-20
C42048 a_1823_45246# a_3992_43940# 1.48e-19
C42049 a_6171_45002# a_9482_43914# 0.016128f
C42050 a_9290_44172# a_11341_43940# 0.040892f
C42051 a_n2438_43548# a_n1641_43230# 4.44e-20
C42052 a_4883_46098# a_17583_46090# 0.012469f
C42053 a_18479_47436# a_20708_46348# 0.04299f
C42054 a_n2661_46634# a_n2840_46090# 3.35e-19
C42055 a_6491_46660# a_5066_45546# 2.85e-21
C42056 a_11453_44696# a_14493_46090# 1.13e-21
C42057 a_13507_46334# a_18189_46348# 0.001569f
C42058 a_19787_47423# a_19553_46090# 9.41e-20
C42059 a_16588_47582# a_10809_44734# 9.65e-20
C42060 a_10227_46804# a_6945_45028# 0.220094f
C42061 a_n1151_42308# a_9823_46482# 1.61e-19
C42062 a_2063_45854# a_11387_46482# 2.86e-19
C42063 a_8270_45546# a_8846_46660# 7.05e-19
C42064 a_n881_46662# a_7920_46348# 0.025724f
C42065 a_n743_46660# a_11415_45002# 0.038831f
C42066 a_768_44030# a_3483_46348# 0.281593f
C42067 a_3067_47026# a_765_45546# 0.002408f
C42068 a_6755_46942# a_3090_45724# 0.050558f
C42069 a_4791_45118# a_8034_45724# 2.34e-20
C42070 a_19386_47436# a_19335_46494# 3.45e-20
C42071 a_18597_46090# a_20075_46420# 0.073857f
C42072 a_12465_44636# a_2324_44458# 0.070016f
C42073 a_8037_42858# a_8605_42826# 0.178024f
C42074 a_7871_42858# a_9127_43156# 0.043633f
C42075 a_7765_42852# a_8387_43230# 4.21e-19
C42076 a_15095_43370# a_15953_42852# 2.26e-19
C42077 a_2982_43646# a_1755_42282# 0.051666f
C42078 a_22223_43396# a_22223_42860# 0.026152f
C42079 a_13887_32519# a_22165_42308# 0.002652f
C42080 a_11341_43940# a_21887_42336# 1.43e-20
C42081 a_3080_42308# a_3318_42354# 0.036372f
C42082 a_n1821_44484# VDD 4.61e-20
C42083 a_n97_42460# a_6761_42308# 0.012266f
C42084 a_n2661_45010# a_n1331_43914# 4.98e-21
C42085 a_n2109_45247# a_n2065_43946# 7.64e-21
C42086 a_n2293_45010# a_n1761_44111# 0.148418f
C42087 a_n2312_38680# a_5742_30871# 4.94e-21
C42088 a_n863_45724# a_3539_42460# 8.25e-22
C42089 a_9482_43914# a_14673_44172# 0.42967f
C42090 a_13556_45296# a_14581_44484# 2.18e-19
C42091 a_n2840_44458# a_n2129_44697# 6.34e-19
C42092 a_n4318_40392# a_n2433_44484# 0.001155f
C42093 a_413_45260# a_3422_30871# 3.37e-19
C42094 a_2437_43646# a_2479_44172# 0.00389f
C42095 a_3357_43084# a_1414_42308# 6.88e-19
C42096 a_4185_45028# a_4520_42826# 0.012305f
C42097 a_16680_45572# a_15682_43940# 1.27e-20
C42098 a_n443_42852# a_n229_43646# 0.001316f
C42099 a_17023_45118# a_14539_43914# 7.91e-19
C42100 a_16922_45042# a_16979_44734# 7.83e-19
C42101 a_n2293_42834# a_7640_43914# 0.040893f
C42102 a_4883_46098# a_8696_44636# 0.023202f
C42103 a_16327_47482# a_16147_45260# 0.017922f
C42104 a_3877_44458# a_3503_45724# 0.001651f
C42105 a_12549_44172# a_15143_45578# 2.08e-21
C42106 a_5257_43370# a_n2661_45546# 0.003554f
C42107 a_3090_45724# a_8049_45260# 1.23904f
C42108 a_1823_45246# a_2804_46116# 1.33e-21
C42109 a_13507_46334# a_17478_45572# 1.05e-20
C42110 a_10227_46804# a_14127_45572# 2.84e-19
C42111 a_19551_46910# a_19335_46494# 6.39e-20
C42112 a_20411_46873# a_18985_46122# 1.23e-19
C42113 a_6755_46942# a_15002_46116# 3.59e-20
C42114 a_4007_47204# a_2437_43646# 0.007098f
C42115 a_12861_44030# a_18799_45938# 6.19e-20
C42116 a_11415_45002# a_11189_46129# 0.001065f
C42117 a_167_45260# a_2521_46116# 0.328009f
C42118 a_n2497_47436# a_327_44734# 1.11e-19
C42119 a_17339_46660# a_6945_45028# 6.42e-20
C42120 a_2107_46812# a_5907_45546# 1.16e-20
C42121 a_11599_46634# a_18691_45572# 0.034093f
C42122 a_11453_44696# a_15903_45785# 0.003342f
C42123 a_5534_30871# a_13070_42354# 0.025818f
C42124 a_17517_44484# a_19006_44850# 0.016181f
C42125 a_17061_44734# a_11967_42832# 2.07e-20
C42126 a_5343_44458# a_9028_43914# 1.94e-20
C42127 a_5111_44636# a_6547_43396# 0.035842f
C42128 a_n1059_45260# a_9803_43646# 1.87e-20
C42129 a_n913_45002# a_9145_43396# 0.004598f
C42130 a_19321_45002# VDD 1.01574f
C42131 a_13747_46662# START 0.062289f
C42132 a_6171_45002# a_6031_43396# 6.47e-22
C42133 a_3232_43370# a_6293_42852# 0.004069f
C42134 a_3537_45260# a_8791_43396# 0.071369f
C42135 a_16119_47582# CLK 2.67e-19
C42136 a_8746_45002# a_10991_42826# 2.47e-21
C42137 a_10193_42453# a_10922_42852# 3.71e-21
C42138 a_n357_42282# a_4649_42852# 0.00298f
C42139 a_n1925_42282# a_961_42354# 8.52e-20
C42140 a_18494_42460# a_14021_43940# 0.026241f
C42141 a_20202_43084# a_22775_42308# 1.98e-19
C42142 a_1307_43914# a_1209_43370# 0.001241f
C42143 a_9290_44172# a_10723_42308# 8.75e-19
C42144 a_5257_43370# a_5205_44484# 0.021038f
C42145 a_13661_43548# a_15060_45348# 6.77e-19
C42146 SMPL_ON_P a_n2661_42834# 0.002304f
C42147 a_n1741_47186# a_n2661_43922# 1.28e-19
C42148 a_19466_46812# a_20731_45938# 1.24e-20
C42149 a_11453_44696# a_n2661_44458# 0.174607f
C42150 a_2324_44458# a_2711_45572# 0.804101f
C42151 a_526_44458# a_n863_45724# 0.801581f
C42152 a_14180_46482# a_14371_46494# 4.61e-19
C42153 a_7577_46660# a_3232_43370# 6.76e-22
C42154 a_7715_46873# a_6171_45002# 3.86e-20
C42155 a_n881_46662# a_11827_44484# 2.46e-20
C42156 a_16388_46812# a_18479_45785# 3.13e-19
C42157 a_15368_46634# a_2437_43646# 1.64e-19
C42158 a_15009_46634# a_3357_43084# 1.23e-20
C42159 a_7920_46348# a_8162_45546# 2.96e-19
C42160 a_3483_46348# a_11652_45724# 0.035818f
C42161 a_8049_45260# a_15002_46116# 1.39e-19
C42162 a_5342_30871# C0_N_btm 8.41e-20
C42163 a_n4318_38216# a_n2946_37984# 4.19e-20
C42164 a_5534_30871# C2_N_btm 7.46e-20
C42165 a_15890_42674# a_4958_30871# 0.017137f
C42166 a_15803_42450# a_17531_42308# 6.07e-21
C42167 a_15959_42545# a_17303_42282# 6.6e-20
C42168 a_n4318_37592# a_n4334_38304# 7.52e-20
C42169 a_n3674_38216# a_n3690_38304# 0.071735f
C42170 a_5742_30871# a_7174_31319# 0.34728f
C42171 a_10922_42852# VDD 0.216186f
C42172 a_6123_31319# a_n3565_39590# 5.77e-21
C42173 a_5934_30871# a_n4209_39590# 1.08e-21
C42174 a_18248_44752# a_18429_43548# 5.65e-19
C42175 a_11823_42460# a_16522_42674# 1.68e-21
C42176 a_10193_42453# a_17531_42308# 7.42e-19
C42177 a_n2810_45572# a_n4064_38528# 2.53e-19
C42178 a_n2017_45002# a_18707_42852# 0.026353f
C42179 a_n2840_43914# a_n2840_43370# 0.025171f
C42180 a_16979_44734# a_15743_43084# 1.34e-20
C42181 a_1307_43914# a_3059_42968# 1.72e-19
C42182 a_5891_43370# a_10341_43396# 0.087957f
C42183 a_9313_44734# a_14579_43548# 0.038528f
C42184 a_17973_43940# a_19478_44306# 0.001007f
C42185 a_18079_43940# a_15493_43396# 1.94e-19
C42186 a_10807_43548# a_11341_43940# 0.049779f
C42187 a_5068_46348# VDD 0.085085f
C42188 a_6453_43914# a_6671_43940# 0.08213f
C42189 a_5066_45546# a_5691_45260# 1.08e-20
C42190 a_6419_46155# a_n2661_43370# 1.94e-20
C42191 a_n2293_46634# a_1414_42308# 0.260739f
C42192 a_11823_42460# a_13527_45546# 0.027805f
C42193 a_12791_45546# a_13163_45724# 1.53e-19
C42194 a_2711_45572# a_16855_45546# 2.31e-22
C42195 a_9049_44484# a_9241_45822# 3.68e-20
C42196 a_n2438_43548# a_n809_44244# 3.12e-21
C42197 a_10227_46804# a_11173_44260# 3.86e-20
C42198 a_12741_44636# a_16981_45144# 5.15e-19
C42199 a_6755_46942# a_14815_43914# 1.72e-19
C42200 a_n971_45724# a_n2267_43396# 3.28e-19
C42201 a_n2497_47436# a_n1809_43762# 0.005726f
C42202 a_n746_45260# a_n2129_43609# 1.13e-21
C42203 a_6945_45028# a_1307_43914# 3.38e-20
C42204 a_n2109_47186# a_2443_46660# 2.98e-19
C42205 a_n1151_42308# a_n2104_46634# 3.6e-20
C42206 a_4007_47204# a_n2661_46634# 1.08e-19
C42207 a_n1435_47204# a_13569_47204# 0.011393f
C42208 a_13381_47204# a_13675_47204# 1.29e-20
C42209 a_6575_47204# a_5807_45002# 1.65e-19
C42210 a_13487_47204# a_768_44030# 0.371206f
C42211 a_n4315_30879# C10_P_btm 1.5848f
C42212 a_7174_31319# C0_dummy_P_btm 0.029132f
C42213 a_11599_46634# a_11309_47204# 0.008095f
C42214 a_n3420_39616# a_n1532_35090# 1.07e-19
C42215 a_n1741_47186# a_1799_45572# 2.42e-19
C42216 a_n1920_47178# a_n2661_46098# 3.04e-20
C42217 a_n746_45260# a_288_46660# 0.010226f
C42218 SMPL_ON_N a_22959_47212# 0.007483f
C42219 a_584_46384# a_n133_46660# 2.89e-19
C42220 a_2063_45854# a_n2438_43548# 0.033724f
C42221 a_7754_39964# a_7754_39300# 3.86e-20
C42222 a_17531_42308# VDD 0.262303f
C42223 a_13258_32519# C1_N_btm 0.001902f
C42224 a_14311_47204# a_12549_44172# 7.38e-20
C42225 a_n4334_38304# a_n4334_37440# 0.050585f
C42226 a_n3565_38216# a_n4209_37414# 5.88577f
C42227 a_n4209_38216# a_n3565_37414# 0.031622f
C42228 a_2905_45572# a_n1925_46634# 0.029452f
C42229 a_n237_47217# a_1983_46706# 8.91e-19
C42230 a_17303_42282# RST_Z 0.002907f
C42231 a_3499_42826# a_2075_43172# 1.63e-19
C42232 a_4223_44672# a_5932_42308# 1.08e-20
C42233 a_n1557_42282# a_1512_43396# 1.26e-20
C42234 a_15493_43940# a_21487_43396# 1.34e-19
C42235 a_11341_43940# a_13467_32519# 0.001199f
C42236 a_3080_42308# a_6197_43396# 3.94e-21
C42237 a_n97_42460# a_7274_43762# 4.27e-20
C42238 SMPL_ON_P a_n2293_42282# 1.31e-19
C42239 a_2107_46812# a_9145_43396# 1.58e-19
C42240 a_n357_42282# a_15004_44636# 2.78e-22
C42241 a_3090_45724# a_15037_43940# 0.007895f
C42242 a_5907_45546# a_n2661_44458# 6.68e-20
C42243 a_12549_44172# a_16867_43762# 7.49e-20
C42244 a_n2293_45010# a_n2956_37592# 0.005894f
C42245 a_n2472_45002# en_comp 0.117861f
C42246 a_19963_31679# a_413_45260# 0.0432f
C42247 a_n2661_45010# a_n967_45348# 0.019427f
C42248 a_13661_43548# a_16409_43396# 0.001637f
C42249 a_11415_45002# a_11750_44172# 6.76e-21
C42250 a_n1059_45260# a_n913_45002# 1.19505f
C42251 a_n2017_45002# a_n745_45366# 7.49e-21
C42252 a_n2109_45247# a_n2810_45028# 4.84e-19
C42253 a_10193_42453# a_18184_42460# 0.216199f
C42254 a_16147_45260# a_14537_43396# 5.04e-19
C42255 a_10586_45546# a_n2661_43922# 6.49e-20
C42256 a_10907_45822# a_n2661_43370# 0.057449f
C42257 a_13059_46348# a_14485_44260# 1.96e-19
C42258 a_n2293_46634# a_12281_43396# 0.007661f
C42259 a_4646_46812# a_6197_43396# 0.601282f
C42260 a_20916_46384# a_15227_44166# 0.681561f
C42261 a_5807_45002# a_10861_46660# 0.00101f
C42262 a_768_44030# a_14513_46634# 8.17e-21
C42263 a_12549_44172# a_14226_46987# 3.77e-19
C42264 a_9067_47204# a_3483_46348# 9.45e-22
C42265 a_5732_46660# a_5894_47026# 0.006453f
C42266 a_5167_46660# a_5429_46660# 0.001705f
C42267 a_4817_46660# a_7411_46660# 1.88e-20
C42268 a_5385_46902# a_5257_43370# 5.44e-20
C42269 a_2063_45854# a_11133_46155# 0.026232f
C42270 a_n1435_47204# a_2202_46116# 1.01e-21
C42271 a_3094_47243# a_765_45546# 4.26e-19
C42272 a_11453_44696# a_17639_46660# 2.16e-19
C42273 a_13507_46334# a_20202_43084# 0.205796f
C42274 a_6151_47436# a_5204_45822# 1.22e-19
C42275 a_4791_45118# a_8016_46348# 0.001293f
C42276 a_n1151_42308# a_9569_46155# 0.05766f
C42277 a_19594_46812# a_19692_46634# 0.134424f
C42278 a_n743_46660# a_12251_46660# 3.96e-20
C42279 a_3877_44458# a_7927_46660# 3.05e-20
C42280 a_4646_46812# a_8145_46902# 1.81e-20
C42281 a_21381_43940# a_22400_42852# 1.44e-20
C42282 a_18184_42460# VDD 2.05053f
C42283 a_10729_43914# a_5742_30871# 1.45e-20
C42284 a_3422_30871# a_n4064_39616# 0.003743f
C42285 a_10807_43548# a_10723_42308# 8.52e-19
C42286 a_10341_43396# a_17595_43084# 3.94e-20
C42287 a_20202_43084# a_21855_43396# 3.14e-20
C42288 a_3090_45724# a_15279_43071# 4.84e-21
C42289 a_n2956_39768# a_n3674_38216# 0.023755f
C42290 a_9290_44172# a_10341_43396# 0.157042f
C42291 a_8199_44636# a_9885_43396# 0.002068f
C42292 a_2711_45572# a_19862_44208# 0.002631f
C42293 a_5111_44636# a_n356_44636# 1.45e-19
C42294 a_10227_46804# a_14456_42282# 6.75e-20
C42295 a_13159_45002# a_13076_44458# 3.32e-19
C42296 a_9482_43914# a_12607_44458# 0.151452f
C42297 a_13017_45260# a_13720_44458# 2.63e-20
C42298 a_n1925_42282# a_2982_43646# 0.036209f
C42299 a_19431_45546# a_11967_42832# 1.18e-20
C42300 a_20107_45572# a_17517_44484# 2.01e-21
C42301 a_1423_45028# a_4223_44672# 0.013079f
C42302 SMPL_ON_P a_n3565_39590# 0.001613f
C42303 a_n2442_46660# a_n2472_42282# 4.03e-20
C42304 a_21588_30879# COMP_P 0.001821f
C42305 a_20916_46384# a_21071_46482# 0.006088f
C42306 a_11735_46660# a_12005_46116# 2.1e-19
C42307 a_11813_46116# a_10903_43370# 0.006138f
C42308 a_12861_44030# a_11962_45724# 0.184706f
C42309 a_3090_45724# a_8953_45546# 0.032771f
C42310 a_11599_46634# a_10490_45724# 1.42e-20
C42311 a_4646_46812# a_5066_45546# 0.020397f
C42312 a_768_44030# a_n357_42282# 0.175577f
C42313 a_6151_47436# a_8697_45822# 1.19e-20
C42314 a_4915_47217# a_10907_45822# 2e-21
C42315 a_20107_46660# a_12741_44636# 0.527863f
C42316 a_4883_46098# a_7227_45028# 1.07e-19
C42317 a_20623_46660# a_20202_43084# 1.78e-20
C42318 a_20273_46660# a_22591_46660# 6.79e-20
C42319 a_10467_46802# a_6945_45028# 1.12e-19
C42320 a_n743_46660# a_13259_45724# 0.025444f
C42321 a_4955_46873# a_5210_46482# 9.61e-19
C42322 a_2905_42968# a_2903_42308# 1.75e-19
C42323 a_16547_43609# a_4958_30871# 6.55e-19
C42324 a_16243_43396# a_17303_42282# 2.6e-19
C42325 a_16137_43396# a_17531_42308# 0.001298f
C42326 a_4361_42308# a_10533_42308# 0.017218f
C42327 a_743_42282# a_11633_42558# 0.005183f
C42328 a_1847_42826# a_3823_42558# 1.7e-20
C42329 a_10922_42852# a_n784_42308# 4.32e-21
C42330 a_10341_43396# a_21887_42336# 2.25e-20
C42331 a_n357_42282# a_5755_42852# 0.179701f
C42332 a_n755_45592# a_5111_42852# 2.12e-20
C42333 a_1307_43914# a_11173_44260# 1.43e-19
C42334 a_5891_43370# a_n2293_43922# 1.56e-19
C42335 a_14539_43914# a_17061_44484# 0.003953f
C42336 a_8238_44734# a_n2661_43922# 7.85e-20
C42337 a_11459_47204# DATA[5] 0.370451f
C42338 a_13259_45724# a_17701_42308# 0.137488f
C42339 a_15811_47375# VDD 0.979053f
C42340 a_526_44458# a_7309_42852# 8.78e-19
C42341 a_1823_45246# a_1755_42282# 9.08e-19
C42342 a_5111_44636# a_9165_43940# 1.1e-19
C42343 en_comp a_14401_32519# 7.39e-20
C42344 a_484_44484# a_556_44484# 0.003395f
C42345 a_n1435_47204# DATA[3] 0.02843f
C42346 a_n4318_40392# a_n2840_43914# 4.88e-19
C42347 a_11823_42460# a_15743_43084# 1.48e-19
C42348 a_n2661_43370# a_n2661_42282# 1.08e-20
C42349 a_n2661_45010# a_n1917_43396# 3.02e-20
C42350 a_n2017_45002# a_n2433_43396# 0.035979f
C42351 a_15507_47210# RST_Z 2.28e-19
C42352 a_18374_44850# a_17517_44484# 0.019155f
C42353 a_8696_44636# a_8685_43396# 2.24e-19
C42354 a_11599_46634# START 2.57e-19
C42355 a_11031_47542# CLK 4.33e-19
C42356 a_6945_45028# a_8034_45724# 4.34e-21
C42357 a_20075_46420# a_8049_45260# 0.005224f
C42358 a_1208_46090# a_n755_45592# 0.004994f
C42359 a_2521_46116# a_n863_45724# 9.29e-20
C42360 a_1176_45822# a_n357_42282# 0.001329f
C42361 a_13747_46662# a_6171_45002# 1.31e-19
C42362 a_n2293_46634# a_1667_45002# 0.009008f
C42363 a_13059_46348# a_10193_42453# 6.88e-21
C42364 a_13925_46122# a_14371_46494# 2.28e-19
C42365 a_n746_45260# a_n2129_44697# 0.17701f
C42366 a_n971_45724# a_n2267_44484# 4.09e-19
C42367 a_5807_45002# a_5205_44484# 3.77e-19
C42368 a_n743_46660# a_n467_45028# 0.001437f
C42369 a_3699_46348# a_n2661_45546# 1.29e-20
C42370 a_n881_46662# a_15595_45028# 7.5e-20
C42371 a_12861_44030# a_13807_45067# 7.89e-20
C42372 a_11813_46116# a_12016_45572# 7.88e-20
C42373 a_n1925_46634# a_n37_45144# 1.2e-20
C42374 a_n1853_46287# a_n310_45899# 9.42e-19
C42375 a_n2497_47436# a_4223_44672# 0.047068f
C42376 a_768_44030# a_11963_45334# 2.59e-20
C42377 a_12891_46348# a_13159_45002# 0.031652f
C42378 a_12549_44172# a_13017_45260# 8.3e-19
C42379 a_12594_46348# a_12839_46116# 0.002912f
C42380 a_5934_30871# a_9293_42558# 0.001273f
C42381 a_4190_30871# C2_N_btm 9.13e-20
C42382 a_5932_42308# a_5742_30871# 1.14154f
C42383 a_8337_42558# a_8685_42308# 4.27e-19
C42384 a_11823_42460# a_1606_42308# 4.73e-20
C42385 a_n443_42852# a_13070_42354# 7.16e-20
C42386 a_n913_45002# a_19987_42826# 4.56e-20
C42387 a_n2017_45002# a_21356_42826# 1.31e-20
C42388 a_8701_44490# a_8791_43396# 1.69e-20
C42389 a_5883_43914# a_8147_43396# 3.36e-20
C42390 a_n2661_44458# a_9145_43396# 2.4e-20
C42391 a_13259_45724# a_21613_42308# 0.077442f
C42392 a_20512_43084# a_20269_44172# 2.47e-20
C42393 a_n356_44636# a_4235_43370# 5.73e-21
C42394 a_13059_46348# VDD 0.955445f
C42395 a_17613_45144# a_17499_43370# 5.51e-21
C42396 a_18184_42460# a_16137_43396# 0.029846f
C42397 a_5891_43370# a_n97_42460# 0.957548f
C42398 a_3422_30871# a_22223_43948# 0.011616f
C42399 a_20640_44752# a_14021_43940# 8.61e-21
C42400 en_comp a_18817_42826# 4.89e-21
C42401 a_5263_45724# a_6194_45824# 1.4e-19
C42402 a_2711_45572# a_6667_45809# 0.010894f
C42403 a_13661_43548# a_16241_44734# 0.047309f
C42404 a_13747_46662# a_14673_44172# 4.77e-21
C42405 a_5204_45822# a_5111_44636# 8.78e-19
C42406 a_5164_46348# a_4927_45028# 0.09665f
C42407 a_5497_46414# a_5147_45002# 4.57e-19
C42408 a_9823_46155# a_413_45260# 2.74e-21
C42409 a_3483_46348# a_7276_45260# 0.003843f
C42410 a_12549_44172# a_19006_44850# 5.76e-20
C42411 a_12891_46348# a_11967_42832# 3.62e-21
C42412 a_19335_46494# a_3357_43084# 2.49e-21
C42413 a_3090_45724# a_20193_45348# 1.53e-20
C42414 a_14976_45028# a_11691_44458# 6.38e-19
C42415 a_19692_46634# a_18494_42460# 6.49e-19
C42416 a_7920_46348# a_3537_45260# 5.32e-20
C42417 a_n2438_43548# a_n2661_42834# 0.057776f
C42418 a_n743_46660# a_n2661_43922# 1.41e-20
C42419 a_n4209_39304# a_n4209_38216# 0.029694f
C42420 a_5932_42308# C0_dummy_P_btm 1.2e-19
C42421 a_2063_45854# a_13507_46334# 7.95e-20
C42422 a_9313_45822# a_n1435_47204# 5.93e-19
C42423 a_11459_47204# a_13381_47204# 3.65e-21
C42424 a_n2302_39072# a_n2302_38778# 0.050477f
C42425 a_n971_45724# a_n2312_39304# 8.21e-21
C42426 a_n452_47436# a_n310_47570# 0.007833f
C42427 a_5934_30871# C6_P_btm 0.004563f
C42428 a_6151_47436# a_16241_47178# 5.05e-20
C42429 a_6123_31319# C4_P_btm 0.132906f
C42430 a_n815_47178# a_n89_47570# 3.25e-20
C42431 a_2903_42308# VDD 0.22017f
C42432 a_n1741_47186# a_2747_46873# 0.00508f
C42433 a_19237_31679# a_17364_32525# 0.054573f
C42434 a_10057_43914# a_10752_42852# 1.23e-20
C42435 a_n2293_42834# a_5932_42308# 2.23e-19
C42436 a_3218_45724# VDD 0.133843f
C42437 a_10807_43548# a_10341_43396# 0.042318f
C42438 a_1414_42308# a_743_42282# 0.004767f
C42439 a_14955_43940# a_14205_43396# 4.77e-19
C42440 a_n2840_43370# a_n4318_39304# 0.158695f
C42441 a_14537_43396# a_15051_42282# 7.92e-20
C42442 a_9313_44734# a_21671_42860# 0.012466f
C42443 a_11322_45546# a_13159_45002# 4.52e-20
C42444 a_13259_45724# a_17969_45144# 8.9e-19
C42445 a_n1613_43370# a_8791_43396# 4.34e-20
C42446 SMPL_ON_P a_n1423_42826# 8.78e-21
C42447 a_n2497_47436# a_n3674_39304# 4.4e-20
C42448 a_11823_42460# a_10775_45002# 2.94e-20
C42449 a_6469_45572# a_6171_45002# 4.62e-19
C42450 a_3483_46348# a_17517_44484# 0.004031f
C42451 a_11415_45002# a_20397_44484# 2.5e-20
C42452 a_11453_44696# a_9145_43396# 2.08e-20
C42453 a_12465_44636# a_14579_43548# 1.92e-21
C42454 a_18175_45572# a_20528_45572# 2.64e-21
C42455 a_19256_45572# a_20107_45572# 4.08e-19
C42456 a_3090_45724# a_9028_43914# 0.00399f
C42457 a_9290_44172# a_n2293_43922# 0.369185f
C42458 a_8746_45002# a_9482_43914# 0.002141f
C42459 a_11652_45724# a_11963_45334# 8.93e-19
C42460 a_11962_45724# a_11787_45002# 4.92e-19
C42461 a_n1925_46634# a_2443_46660# 0.054751f
C42462 a_n743_46660# a_1799_45572# 0.034264f
C42463 a_n133_46660# a_479_46660# 3.82e-19
C42464 a_22459_39145# VDD 0.682253f
C42465 a_4883_46098# a_11813_46116# 0.019696f
C42466 a_10227_46804# a_15559_46634# 7.04e-19
C42467 a_601_46902# a_491_47026# 0.097745f
C42468 a_383_46660# a_288_46660# 0.049827f
C42469 a_n1021_46688# a_n2661_46098# 3.91e-20
C42470 a_n2661_46634# a_2864_46660# 0.002851f
C42471 a_n2293_46634# a_2959_46660# 1.76e-20
C42472 a_8128_46384# a_7927_46660# 0.007223f
C42473 a_12861_44030# a_12978_47026# 6.43e-21
C42474 a_11599_46634# a_12156_46660# 2.63e-20
C42475 a_1123_46634# a_1983_46706# 9.93e-19
C42476 a_948_46660# a_2107_46812# 1.97e-20
C42477 a_5807_45002# a_5385_46902# 2.87e-19
C42478 EN_VIN_BSTR_P C4_P_btm 0.116925f
C42479 a_4915_47217# a_14226_46660# 1.65e-19
C42480 a_4007_47204# a_765_45546# 0.00663f
C42481 a_n97_42460# a_17595_43084# 0.0027f
C42482 a_20974_43370# a_21671_42860# 8.3e-20
C42483 a_3905_42865# a_5267_42460# 9.02e-20
C42484 a_n2661_42282# COMP_P 0.02767f
C42485 a_16977_43638# a_16867_43762# 0.097745f
C42486 a_16759_43396# a_16664_43396# 0.049827f
C42487 a_16137_43396# a_15868_43402# 5.04e-20
C42488 a_13556_45296# VDD 0.569056f
C42489 a_18525_43370# a_18783_43370# 0.22264f
C42490 a_18429_43548# a_15743_43084# 0.053516f
C42491 a_14205_43396# a_5649_42852# 4.06e-21
C42492 a_10341_43396# a_13467_32519# 0.007243f
C42493 a_3626_43646# a_8037_42858# 5.94e-20
C42494 a_2982_43646# a_8387_43230# 3.53e-20
C42495 a_12281_43396# a_743_42282# 0.036414f
C42496 a_n2017_45002# a_n2433_44484# 0.039498f
C42497 a_n1059_45260# a_n2661_44458# 0.028647f
C42498 a_3357_43084# a_n699_43396# 0.004379f
C42499 a_8049_45260# a_9248_44260# 1.1e-21
C42500 a_9290_44172# a_n97_42460# 0.351467f
C42501 a_n2293_45010# a_n2267_44484# 0.0118f
C42502 a_n2109_45247# a_n2129_44697# 0.003166f
C42503 a_n2661_45010# a_n1917_44484# 0.015623f
C42504 a_n2438_43548# a_n2293_42282# 1.27e-19
C42505 a_4791_45118# a_3905_42558# 8.4e-21
C42506 a_18596_45572# a_18443_44721# 1.58e-20
C42507 a_18799_45938# a_18287_44626# 2.22e-20
C42508 a_8696_44636# a_8783_44734# 7.48e-19
C42509 a_n443_42852# a_2127_44172# 5.26e-20
C42510 a_1423_45028# a_n2293_42834# 0.033636f
C42511 a_n237_47217# a_6194_45824# 2.56e-20
C42512 a_n971_45724# a_6511_45714# 0.001043f
C42513 a_3877_44458# a_5164_46348# 7.65e-19
C42514 a_4646_46812# a_5068_46348# 5.4e-20
C42515 a_9804_47204# a_5066_45546# 1.22e-21
C42516 a_4883_46098# a_14949_46494# 2.19e-19
C42517 a_21588_30879# a_10809_44734# 0.110956f
C42518 a_20916_46384# a_22959_46124# 7.06e-20
C42519 a_4651_46660# a_4704_46090# 0.013135f
C42520 a_18597_46090# a_19431_46494# 0.004523f
C42521 a_n743_46660# a_18189_46348# 1.08e-19
C42522 a_5167_46660# a_3483_46348# 1.48e-21
C42523 a_4955_46873# a_4419_46090# 7.36e-20
C42524 a_16327_47482# a_20062_46116# 1.2e-19
C42525 a_12465_44636# a_12839_46116# 4.88e-21
C42526 a_3090_45724# a_18285_46348# 1.81e-20
C42527 a_15559_46634# a_17339_46660# 1.11e-20
C42528 a_15368_46634# a_765_45546# 5.6e-19
C42529 a_n881_46662# a_8062_46482# 0.001601f
C42530 a_3422_30871# C0_P_btm 6.53e-20
C42531 a_19987_42826# a_20922_43172# 0.001853f
C42532 a_3626_43646# a_13921_42308# 5.3e-19
C42533 a_20362_44736# VDD 0.275577f
C42534 a_13467_32519# a_20356_42852# 1.53e-20
C42535 a_13678_32519# a_14097_32519# 0.04945f
C42536 a_5649_42852# a_22400_42852# 6.16e-20
C42537 a_16979_44734# a_17970_44736# 5.21e-19
C42538 a_14539_43914# a_18248_44752# 5.77e-20
C42539 a_4223_44672# a_6109_44484# 0.003455f
C42540 a_n2129_44697# a_n310_44484# 2.88e-19
C42541 a_11827_44484# a_11541_44484# 0.0442f
C42542 a_1423_45028# a_1115_44172# 3.06e-20
C42543 a_5147_45002# a_5841_44260# 1.74e-19
C42544 a_n357_42282# a_16759_43396# 0.007988f
C42545 a_13259_45724# a_4361_42308# 0.054653f
C42546 a_n443_42852# a_8945_43396# 3.77e-20
C42547 a_n2442_46660# a_n2216_39866# 0.003462f
C42548 a_17719_45144# a_17517_44484# 1.47e-19
C42549 a_1307_43914# a_895_43940# 0.754684f
C42550 a_626_44172# a_1414_42308# 0.002821f
C42551 a_7499_43078# a_7287_43370# 0.057949f
C42552 a_8270_45546# a_8685_42308# 2.23e-21
C42553 a_526_44458# a_7765_42852# 0.023934f
C42554 a_n1059_45260# a_18451_43940# 2.97e-21
C42555 a_11691_44458# a_15433_44458# 0.110923f
C42556 a_12005_46116# a_2324_44458# 9.1e-21
C42557 a_8016_46348# a_6945_45028# 4.6e-20
C42558 a_11453_44696# a_n1059_45260# 1.65e-20
C42559 a_19787_47423# a_413_45260# 8.86e-20
C42560 a_13759_46122# a_14275_46494# 0.105995f
C42561 a_13925_46122# a_14493_46090# 0.17072f
C42562 a_167_45260# a_2981_46116# 4.98e-19
C42563 a_21076_30879# a_8049_45260# 6.53e-20
C42564 a_3090_45724# a_1609_45822# 3.9e-19
C42565 a_19321_45002# a_18479_45785# 0.114441f
C42566 a_13661_43548# a_18691_45572# 0.020905f
C42567 a_5807_45002# a_19431_45546# 0.01527f
C42568 a_13747_46662# a_18909_45814# 0.025022f
C42569 a_12549_44172# a_20107_45572# 2.47e-19
C42570 a_5063_47570# a_2437_43646# 8.52e-19
C42571 a_11599_46634# a_6171_45002# 3.62e-19
C42572 a_n2497_47436# a_n2293_42834# 0.010004f
C42573 a_1823_45246# a_n1925_42282# 0.099018f
C42574 a_2202_46116# a_526_44458# 2.44e-20
C42575 a_8492_46660# a_7499_43078# 1.8e-19
C42576 a_n743_46660# a_17478_45572# 9.46e-19
C42577 a_1576_42282# a_2123_42473# 4.32e-19
C42578 a_1184_42692# a_1755_42282# 0.016329f
C42579 a_13291_42460# a_13575_42558# 0.074792f
C42580 a_14635_42282# a_13070_42354# 2.81e-20
C42581 a_14097_32519# a_6123_31319# 0.003315f
C42582 a_6293_42852# VDD 0.401011f
C42583 a_n784_42308# a_2903_42308# 3.86e-20
C42584 a_n4318_40392# a_n4318_39304# 0.024428f
C42585 a_n2661_45010# a_n1853_43023# 1.08e-20
C42586 a_n863_45724# a_1221_42558# 0.003967f
C42587 a_16922_45042# a_2982_43646# 0.010868f
C42588 a_9313_44734# a_19478_44306# 5.64e-21
C42589 a_9838_44484# a_9801_43940# 2.53e-21
C42590 a_n755_45592# a_n1630_35242# 0.044103f
C42591 a_n357_42282# a_1067_42314# 5.85e-20
C42592 a_n2293_43922# a_10807_43548# 1.85e-21
C42593 a_n2661_42834# a_12429_44172# 0.002835f
C42594 a_n2661_43922# a_11750_44172# 3.46e-20
C42595 a_7577_46660# VDD 0.249866f
C42596 a_n2661_45546# a_n755_45592# 0.14317f
C42597 a_n743_46660# a_n452_44636# 3.36e-20
C42598 a_n2293_46634# a_n699_43396# 0.016884f
C42599 a_n971_45724# a_n2065_43946# 0.016306f
C42600 a_n2497_47436# a_1115_44172# 0.069778f
C42601 a_n1613_43370# a_n1243_44484# 6.03e-19
C42602 a_n863_45724# a_n452_45724# 0.046903f
C42603 a_12549_44172# a_18374_44850# 2.67e-20
C42604 a_20107_46660# a_413_45260# 1.46e-20
C42605 a_10227_46804# a_15463_44811# 1.33e-19
C42606 a_n2293_45546# a_n1099_45572# 0.004814f
C42607 a_10809_44734# a_10907_45822# 0.003912f
C42608 a_14840_46494# a_15037_45618# 1.08e-19
C42609 a_15227_44166# a_14797_45144# 0.011685f
C42610 a_11599_46634# a_14673_44172# 3.2e-21
C42611 a_20202_43084# a_21297_45572# 2.32e-19
C42612 a_11415_45002# a_20447_31679# 2.6e-19
C42613 a_21076_30879# a_19479_31679# 0.054875f
C42614 a_20820_30879# a_19963_31679# 0.057032f
C42615 a_11554_42852# VDD 0.078978f
C42616 COMP_P a_22469_39537# 0.0359f
C42617 a_n4315_30879# a_n4334_40480# 0.253307f
C42618 a_n237_47217# a_n785_47204# 0.018044f
C42619 a_n971_45724# a_1209_47178# 0.034982f
C42620 a_n1741_47186# a_2063_45854# 0.037801f
C42621 a_n2109_47186# a_2952_47436# 0.050821f
C42622 a_n746_45260# a_327_47204# 0.022743f
C42623 a_n452_47436# a_1239_47204# 7.81e-21
C42624 a_n2833_47464# a_n1151_42308# 2.4e-19
C42625 a_22315_44484# a_10341_43396# 7.96e-19
C42626 a_11967_42832# a_16409_43396# 0.004815f
C42627 a_n356_44636# a_791_42968# 0.003419f
C42628 a_20365_43914# a_19741_43940# 8.59e-20
C42629 a_11341_43940# a_19319_43548# 0.042701f
C42630 a_20269_44172# a_21381_43940# 1.62e-20
C42631 en_comp a_5934_30871# 0.028694f
C42632 a_n1059_45260# a_8325_42308# 6.3e-20
C42633 a_n2017_45002# a_8685_42308# 0.016058f
C42634 a_n913_45002# a_8337_42558# 5.84e-19
C42635 a_3499_42826# a_4699_43561# 4.46e-21
C42636 a_n2661_42282# a_1568_43370# 1.94e-21
C42637 a_10807_43548# a_n97_42460# 5.41e-19
C42638 a_5663_43940# a_6031_43396# 1.67e-19
C42639 a_1414_42308# a_2813_43396# 0.00815f
C42640 a_19862_44208# a_14401_32519# 2.61e-20
C42641 a_20205_31679# a_22521_39511# 3.28e-20
C42642 a_n1925_42282# DATA[2] 9.03e-20
C42643 a_8016_46348# a_8103_44636# 8.07e-22
C42644 a_22223_46124# a_11827_44484# 4.45e-19
C42645 a_15599_45572# a_15903_45785# 0.161702f
C42646 a_15297_45822# a_15765_45572# 3.14e-20
C42647 a_19692_46634# a_20640_44752# 0.001236f
C42648 a_8049_45260# a_8488_45348# 7.56e-19
C42649 a_5937_45572# a_5343_44458# 0.024374f
C42650 a_1609_45822# a_2274_45254# 0.11737f
C42651 a_n443_42852# a_2382_45260# 0.020006f
C42652 a_15227_44166# a_20766_44850# 3.54e-21
C42653 a_4791_45118# a_8791_43396# 1.84e-20
C42654 a_19321_45002# a_14021_43940# 1.97e-19
C42655 a_13661_43548# a_15037_44260# 0.003411f
C42656 a_20075_46420# a_20193_45348# 4.06e-21
C42657 a_3483_46348# a_13720_44458# 0.010665f
C42658 a_n2860_38778# VDD 0.004252f
C42659 a_n1741_47186# a_12469_46902# 4.21e-19
C42660 a_2063_45854# a_7832_46660# 0.011867f
C42661 a_n237_47217# a_8601_46660# 1.58e-19
C42662 a_2747_46873# a_n743_46660# 1.24e-19
C42663 a_n1151_42308# a_6969_46634# 2.33e-19
C42664 a_4915_47217# a_9863_46634# 8.01e-20
C42665 a_6151_47436# a_7927_46660# 0.182356f
C42666 a_6491_46660# a_7577_46660# 4.53e-20
C42667 a_12891_46348# a_5807_45002# 0.044188f
C42668 a_n1435_47204# a_6540_46812# 2.44e-21
C42669 a_7227_47204# a_7411_46660# 0.011806f
C42670 a_4338_37500# a_11206_38545# 0.072616f
C42671 a_5700_37509# a_8912_37509# 15.051701f
C42672 a_8530_39574# CAL_P 0.037066f
C42673 a_3726_37500# CAL_N 0.036205f
C42674 a_5088_37509# VDAC_P 1.15441f
C42675 a_6886_37412# VDAC_N 0.067053f
C42676 a_15493_43396# a_19339_43156# 3.83e-19
C42677 a_19328_44172# a_19164_43230# 2.78e-20
C42678 a_n4318_40392# a_n4334_40480# 0.089305f
C42679 a_3422_30871# a_20753_42852# 0.048434f
C42680 a_5891_43370# a_10533_42308# 5.45e-19
C42681 a_20512_43084# a_20836_43172# 8.79e-20
C42682 a_8685_43396# a_14205_43396# 0.011249f
C42683 a_n356_44636# a_15051_42282# 8.17e-19
C42684 a_2982_43646# a_15743_43084# 0.023587f
C42685 a_15493_43940# a_15567_42826# 6.99e-20
C42686 a_21363_45546# VDD 0.36538f
C42687 a_6171_45002# a_13348_45260# 0.009869f
C42688 a_3232_43370# a_9482_43914# 0.129525f
C42689 a_3065_45002# a_1307_43914# 0.033168f
C42690 a_413_45260# a_1423_45028# 0.194002f
C42691 a_8191_45002# a_8953_45002# 1.72e-19
C42692 a_8199_44636# a_9895_44260# 0.002714f
C42693 a_8953_45546# a_9248_44260# 4.19e-20
C42694 a_n443_42852# a_15433_44458# 1.08e-21
C42695 a_1667_45002# a_626_44172# 1.79e-19
C42696 a_18909_45814# a_18911_45144# 0.0027f
C42697 a_18479_45785# a_18184_42460# 3.17e-20
C42698 a_768_44030# a_8952_43230# 2.43e-19
C42699 a_8270_45546# a_9803_43646# 0.066865f
C42700 a_2324_44458# a_15682_43940# 0.321744f
C42701 a_n2293_45010# a_117_45144# 2.83e-21
C42702 a_1823_45246# a_3737_43940# 8.92e-19
C42703 a_n2438_43548# a_n1423_42826# 9.01e-21
C42704 a_4883_46098# a_15682_46116# 0.06363f
C42705 a_18479_47436# a_19900_46494# 0.001423f
C42706 a_16763_47508# a_10809_44734# 2.22e-19
C42707 a_n2956_39768# a_n2840_46090# 6.87e-19
C42708 a_6545_47178# a_5066_45546# 0.021464f
C42709 a_11453_44696# a_13925_46122# 3.96e-21
C42710 a_13507_46334# a_17715_44484# 0.003011f
C42711 a_19787_47423# a_18985_46122# 5.06e-20
C42712 a_10227_46804# a_21137_46414# 1.29e-19
C42713 a_17591_47464# a_6945_45028# 0.025004f
C42714 a_2063_45854# a_10586_45546# 0.056181f
C42715 a_8270_45546# a_8601_46660# 8.69e-20
C42716 a_n881_46662# a_6419_46155# 0.019005f
C42717 a_n1151_42308# a_9241_46436# 5.09e-19
C42718 a_12549_44172# a_3483_46348# 0.185475f
C42719 a_2864_46660# a_765_45546# 8.25e-19
C42720 a_6755_46942# a_15009_46634# 0.012747f
C42721 a_19386_47436# a_19553_46090# 2.56e-20
C42722 a_18597_46090# a_19335_46494# 0.036056f
C42723 a_12465_44636# a_14840_46494# 2.12e-20
C42724 a_648_43396# a_564_42282# 1.99e-20
C42725 a_7871_42858# a_8387_43230# 0.106107f
C42726 a_7765_42852# a_8605_42826# 6.55e-19
C42727 a_15095_43370# a_15597_42852# 0.071983f
C42728 a_14579_43548# a_16877_42852# 2.78e-22
C42729 a_2982_43646# a_1606_42308# 0.021878f
C42730 a_13887_32519# a_21671_42860# 5.19e-19
C42731 a_22223_43396# a_22165_42308# 0.00197f
C42732 a_4235_43370# a_3823_42558# 3.1e-19
C42733 a_3080_42308# a_2903_42308# 0.154008f
C42734 a_n1190_44850# VDD 5.02e-19
C42735 a_14021_43940# a_17531_42308# 1.76e-21
C42736 a_n97_42460# a_6773_42558# 6.7e-19
C42737 a_13678_32519# a_22959_42860# 4.44e-20
C42738 a_5649_42852# a_22223_42860# 5.33e-19
C42739 a_16922_45042# a_14539_43914# 0.001347f
C42740 a_7639_45394# a_7640_43914# 2.67e-20
C42741 a_n2840_44458# a_n2433_44484# 0.039807f
C42742 a_n2293_45010# a_n2065_43946# 0.023134f
C42743 a_n2661_45010# a_n1899_43946# 2.77e-19
C42744 a_n863_45724# a_3626_43646# 1.16e-20
C42745 a_13556_45296# a_13940_44484# 8.88e-19
C42746 a_n4318_40392# a_n2661_44458# 0.026979f
C42747 a_2437_43646# a_2127_44172# 0.017247f
C42748 a_12741_44636# a_15567_42826# 1.49e-21
C42749 a_n2661_43370# a_n310_44811# 3.23e-19
C42750 en_comp a_20512_43084# 4.89e-21
C42751 a_8696_44636# a_13483_43940# 9.44e-22
C42752 a_16855_45546# a_15682_43940# 4.92e-20
C42753 a_16327_47482# a_17786_45822# 1.4e-20
C42754 a_3877_44458# a_3316_45546# 9.66e-20
C42755 a_15009_46634# a_8049_45260# 2.77e-21
C42756 a_1823_45246# a_2698_46116# 2.13e-21
C42757 a_n1151_42308# a_3357_43084# 0.028306f
C42758 a_10227_46804# a_14033_45572# 2.4e-19
C42759 a_12549_44172# a_14495_45572# 4.78e-19
C42760 a_768_44030# a_13249_42308# 0.012496f
C42761 a_20411_46873# a_18819_46122# 2.15e-20
C42762 a_19551_46910# a_19553_46090# 2.94e-19
C42763 a_11813_46116# a_11608_46482# 9.21e-19
C42764 a_19123_46287# a_19335_46494# 3.12e-19
C42765 a_3815_47204# a_2437_43646# 0.012198f
C42766 a_12861_44030# a_18596_45572# 0.007922f
C42767 a_11415_45002# a_9290_44172# 0.031886f
C42768 a_n2497_47436# a_413_45260# 0.028795f
C42769 a_n746_45260# a_n745_45366# 0.119822f
C42770 a_2107_46812# a_5263_45724# 7.2e-22
C42771 a_11599_46634# a_18909_45814# 0.042943f
C42772 a_11453_44696# a_15599_45572# 4.53e-20
C42773 a_7499_43940# VDD 0.193884f
C42774 a_5534_30871# a_12563_42308# 0.179331f
C42775 a_13460_43230# a_13575_42558# 1.38e-19
C42776 a_5343_44458# a_8333_44056# 0.092296f
C42777 a_n356_44636# a_3905_42865# 3.95e-20
C42778 a_17517_44484# a_18588_44850# 0.026595f
C42779 a_5111_44636# a_6765_43638# 0.022146f
C42780 a_5147_45002# a_6547_43396# 2e-19
C42781 a_4185_45028# a_15890_42674# 6.54e-20
C42782 a_21076_30879# a_13258_32519# 0.059077f
C42783 a_n1059_45260# a_9145_43396# 0.016142f
C42784 a_n913_45002# a_8423_43396# 7.65e-20
C42785 a_13661_43548# START 0.012406f
C42786 a_3232_43370# a_6031_43396# 4.81e-20
C42787 a_5883_43914# a_n2661_42282# 0.107496f
C42788 a_3537_45260# a_8147_43396# 0.088185f
C42789 a_13747_46662# RST_Z 0.001276f
C42790 a_10193_42453# a_10991_42826# 5.97e-20
C42791 a_n357_42282# a_4149_42891# 2.65e-19
C42792 a_n1925_42282# a_1184_42692# 5.67e-20
C42793 a_526_44458# a_961_42354# 2.74e-21
C42794 a_13259_45724# a_13622_42852# 1.68e-19
C42795 a_18184_42460# a_14021_43940# 0.029776f
C42796 a_20202_43084# a_21613_42308# 0.07574f
C42797 a_1307_43914# a_458_43396# 3.65e-20
C42798 a_9290_44172# a_10533_42308# 0.001105f
C42799 a_7499_43078# a_12089_42308# 9.57e-21
C42800 a_n443_42852# a_1709_42852# 5.75e-21
C42801 a_14976_45028# a_2437_43646# 1.11e-19
C42802 a_11599_46634# a_12607_44458# 1.01e-22
C42803 a_13661_43548# a_14976_45348# 9.13e-21
C42804 a_3483_46348# a_11525_45546# 2.41e-19
C42805 a_8270_45546# a_n913_45002# 1.44e-20
C42806 a_19692_46634# a_21188_45572# 7.15e-19
C42807 a_19466_46812# a_20528_45572# 0.157758f
C42808 a_7715_46873# a_3232_43370# 1.19e-20
C42809 a_16388_46812# a_18175_45572# 1.3e-20
C42810 a_5937_45572# a_4880_45572# 1.79e-19
C42811 a_12549_44172# a_17719_45144# 2.85e-20
C42812 a_7411_46660# a_6171_45002# 4.46e-21
C42813 a_5342_30871# C0_dummy_N_btm 1.91e-20
C42814 a_n4318_38216# a_n3420_37984# 0.001387f
C42815 a_n3674_37592# a_n4064_38528# 0.019942f
C42816 a_5534_30871# C1_N_btm 1.06e-19
C42817 a_15959_42545# a_4958_30871# 0.043235f
C42818 a_15803_42450# a_17303_42282# 0.00508f
C42819 a_n4318_37592# a_n4209_38216# 1.11e-19
C42820 a_15890_42674# a_16269_42308# 3.16e-19
C42821 a_n3674_38216# a_n3565_38216# 0.128699f
C42822 a_11323_42473# a_7174_31319# 4.88e-21
C42823 a_10991_42826# VDD 0.201891f
C42824 a_n699_43396# a_743_42282# 3.69e-20
C42825 a_10193_42453# a_17303_42282# 0.028322f
C42826 a_4704_46090# VDD 0.225404f
C42827 a_17973_43940# a_15493_43396# 8.43e-20
C42828 a_14539_43914# a_15743_43084# 0.024623f
C42829 a_1307_43914# a_2987_42968# 3.55e-20
C42830 a_9313_44734# a_13667_43396# 2.37e-20
C42831 a_5891_43370# a_9885_43646# 0.004104f
C42832 a_n2956_38216# a_n3565_38502# 0.072968f
C42833 a_9028_43914# a_9248_44260# 0.009965f
C42834 a_10949_43914# a_11341_43940# 0.0383f
C42835 a_18326_43940# a_18451_43940# 0.145292f
C42836 a_11453_44696# a_18326_43940# 3.74e-20
C42837 a_5937_45572# a_8560_45348# 0.045711f
C42838 a_6165_46155# a_n2661_43370# 9.24e-21
C42839 a_n2293_46634# a_1467_44172# 3.1e-20
C42840 a_n1613_43370# a_6756_44260# 0.00105f
C42841 a_11823_42460# a_13163_45724# 0.038493f
C42842 a_2711_45572# a_16115_45572# 0.00431f
C42843 a_9049_44484# a_8697_45822# 7.16e-20
C42844 a_n2438_43548# a_n1549_44318# 3.51e-20
C42845 a_12741_44636# a_16886_45144# 4.07e-19
C42846 a_5066_45546# a_4927_45028# 0.001602f
C42847 a_n2497_47436# a_n2012_43396# 1.4e-19
C42848 a_n971_45724# a_n2129_43609# 0.173854f
C42849 a_10227_46804# a_10555_44260# 1.96e-19
C42850 a_n1151_42308# a_n2293_46634# 0.02925f
C42851 a_3815_47204# a_n2661_46634# 9.75e-20
C42852 a_7903_47542# a_5807_45002# 1.29e-20
C42853 a_13381_47204# a_13569_47204# 3.03e-20
C42854 a_12861_44030# a_768_44030# 0.260776f
C42855 a_13487_47204# a_12549_44172# 0.036506f
C42856 a_7174_31319# C0_P_btm 0.050478f
C42857 a_n2109_47186# a_n2661_46098# 3.71e-19
C42858 a_n971_45724# a_288_46660# 9.88e-20
C42859 SMPL_ON_N a_11453_44696# 0.147722f
C42860 a_22731_47423# a_22959_47212# 0.08444f
C42861 a_584_46384# a_n2438_43548# 0.099362f
C42862 a_2063_45854# a_n743_46660# 1.58762f
C42863 a_17303_42282# VDD 0.379254f
C42864 a_13258_32519# C0_N_btm 0.033333f
C42865 a_n4209_38216# a_n4334_37440# 5.82e-19
C42866 a_n4334_38304# a_n4209_37414# 6.38e-20
C42867 a_327_47204# a_383_46660# 0.001388f
C42868 a_n237_47217# a_2107_46812# 0.086093f
C42869 a_4958_30871# RST_Z 0.087554f
C42870 a_3499_42826# a_1847_42826# 0.006199f
C42871 en_comp a_7754_40130# 0.011333f
C42872 a_2982_43646# a_3539_42460# 0.01563f
C42873 a_3540_43646# a_3626_43646# 0.100706f
C42874 a_n1557_42282# a_648_43396# 0.048175f
C42875 a_4699_43561# a_6197_43396# 9.72e-21
C42876 a_19319_43548# a_10341_43396# 0.027205f
C42877 a_n97_42460# a_5837_43396# 6.05e-19
C42878 a_9313_44734# a_20256_43172# 0.0039f
C42879 a_n2017_45002# a_n913_45002# 0.275686f
C42880 a_n2293_45010# a_n2810_45028# 7.12e-19
C42881 a_22591_45572# a_413_45260# 0.003236f
C42882 a_12549_44172# a_16664_43396# 9.47e-20
C42883 a_n443_42852# a_5343_44458# 0.057128f
C42884 a_4646_46812# a_6293_42852# 0.030189f
C42885 a_n2472_45002# a_n2956_37592# 0.152938f
C42886 a_n2661_45010# en_comp 0.10363f
C42887 a_13661_43548# a_16547_43609# 1.23e-19
C42888 a_2437_43646# a_2382_45260# 0.005858f
C42889 a_10193_42453# a_19778_44110# 8.12e-21
C42890 a_16147_45260# a_14180_45002# 4.1e-21
C42891 a_10907_45822# a_11361_45348# 1.86e-19
C42892 a_10586_45546# a_n2661_42834# 3.13e-20
C42893 SMPL_ON_N a_17364_32525# 0.029237f
C42894 a_13059_46348# a_14021_43940# 0.082427f
C42895 a_n2293_46634# a_12293_43646# 0.001258f
C42896 a_2107_46812# a_8270_45546# 0.047835f
C42897 a_12549_44172# a_14513_46634# 0.008065f
C42898 a_768_44030# a_14180_46812# 0.009222f
C42899 a_4817_46660# a_5257_43370# 4.13e-19
C42900 a_5167_46660# a_5263_46660# 0.013793f
C42901 a_5385_46902# a_5429_46660# 3.69e-19
C42902 a_2063_45854# a_11189_46129# 0.294233f
C42903 a_n1435_47204# a_1823_45246# 1.9e-20
C42904 a_6151_47436# a_5164_46348# 5.71e-20
C42905 a_4915_47217# a_6165_46155# 3.17e-20
C42906 a_4791_45118# a_7920_46348# 1.09e-19
C42907 a_n1151_42308# a_9625_46129# 0.046431f
C42908 a_19594_46812# a_19466_46812# 0.100902f
C42909 a_19321_45002# a_19692_46634# 0.040279f
C42910 a_3877_44458# a_8145_46902# 1.22e-20
C42911 a_4646_46812# a_7577_46660# 0.002516f
C42912 a_13507_46334# a_22365_46825# 0.033904f
C42913 a_n97_42460# a_18695_43230# 0.001854f
C42914 a_19778_44110# VDD 0.469922f
C42915 a_22959_43396# a_17364_32525# 0.156288f
C42916 a_10807_43548# a_10533_42308# 4.25e-19
C42917 a_10341_43396# a_16795_42852# 1.46e-20
C42918 a_3090_45724# a_5534_30871# 0.001578f
C42919 a_9290_44172# a_9885_43646# 0.008596f
C42920 a_n357_42282# a_726_44056# 4.98e-19
C42921 a_8016_46348# a_10149_43396# 1.24e-19
C42922 a_626_44172# a_n699_43396# 0.042617f
C42923 a_10227_46804# a_13575_42558# 0.001718f
C42924 a_20202_43084# a_4361_42308# 0.472299f
C42925 a_n2956_39768# a_n2104_42282# 3.63e-20
C42926 a_2711_45572# a_19478_44306# 0.006321f
C42927 a_13348_45260# a_12607_44458# 5.28e-21
C42928 a_13017_45260# a_13076_44458# 0.011055f
C42929 a_526_44458# a_2982_43646# 0.048644f
C42930 a_1423_45028# a_2779_44458# 0.246285f
C42931 a_2382_45260# a_4181_44734# 7.54e-21
C42932 a_18479_45785# a_20362_44736# 2.03e-36
C42933 a_9482_43914# a_8975_43940# 0.186623f
C42934 a_1307_43914# a_6298_44484# 4.3e-19
C42935 a_n2442_46660# a_n3674_38680# 0.023617f
C42936 a_3483_46348# a_16977_43638# 4.05e-19
C42937 a_4883_46098# a_6598_45938# 6.94e-20
C42938 a_20916_46384# a_20850_46482# 4.71e-19
C42939 a_11813_46116# a_11387_46155# 0.080527f
C42940 a_11735_46660# a_10903_43370# 0.002577f
C42941 a_3090_45724# a_5937_45572# 0.002157f
C42942 a_3877_44458# a_5066_45546# 6.79e-20
C42943 a_12549_44172# a_n357_42282# 1.1e-19
C42944 a_2063_45854# a_11136_45572# 0.054713f
C42945 a_6545_47178# a_6977_45572# 9.76e-20
C42946 a_20107_46660# a_20820_30879# 2.92e-20
C42947 a_19551_46910# a_12741_44636# 2.24e-19
C42948 a_20841_46902# a_20202_43084# 3.14e-20
C42949 a_20273_46660# a_11415_45002# 2.53e-20
C42950 a_n881_46662# a_n310_45899# 5.94e-19
C42951 a_n743_46660# a_14383_46116# 0.00314f
C42952 a_10428_46928# a_6945_45028# 8.06e-21
C42953 a_4955_46873# a_4365_46436# 7.84e-21
C42954 a_2905_42968# a_2713_42308# 1.96e-19
C42955 a_16243_43396# a_4958_30871# 2.01e-19
C42956 a_16137_43396# a_17303_42282# 8.65e-19
C42957 a_1847_42826# a_3318_42354# 9.4e-21
C42958 a_743_42282# a_11551_42558# 0.014689f
C42959 a_10991_42826# a_n784_42308# 4.32e-21
C42960 a_n755_45592# a_4520_42826# 2.49e-20
C42961 a_n357_42282# a_5111_42852# 0.011577f
C42962 a_1307_43914# a_10555_44260# 5.81e-19
C42963 a_5891_43370# a_n2661_43922# 0.042536f
C42964 a_14539_43914# a_16789_44484# 3.44e-19
C42965 a_n2840_44458# a_n2840_43914# 0.026152f
C42966 SMPL_ON_N a_21589_35634# 0.399184f
C42967 a_9313_45822# DATA[5] 0.055804f
C42968 a_13259_45724# a_17595_43084# 0.118887f
C42969 a_526_44458# a_5837_42852# 0.057897f
C42970 a_1823_45246# a_1606_42308# 6.6e-20
C42971 a_13556_45296# a_14021_43940# 1.12e-19
C42972 a_5111_44636# a_8487_44056# 0.004423f
C42973 en_comp a_21381_43940# 3.87e-21
C42974 a_n1435_47204# DATA[2] 0.028258f
C42975 a_n2293_45010# a_n2129_43609# 8.68e-20
C42976 a_n2661_45010# a_n1699_43638# 6.02e-20
C42977 a_n2017_45002# a_n4318_39304# 9.41e-20
C42978 a_11599_46634# RST_Z 2.3e-19
C42979 a_18443_44721# a_17517_44484# 0.029904f
C42980 a_9863_47436# CLK 0.00103f
C42981 a_15507_47210# VDD 0.441662f
C42982 a_19335_46494# a_8049_45260# 0.001373f
C42983 a_12005_46116# a_12839_46116# 6e-19
C42984 a_472_46348# a_997_45618# 6.4e-19
C42985 a_167_45260# a_n863_45724# 0.424358f
C42986 a_n2293_46098# a_7_45899# 3.19e-19
C42987 a_n237_47217# a_n2661_44458# 1.04e-19
C42988 a_n746_45260# a_n2433_44484# 2.7e-20
C42989 a_5807_45002# a_6431_45366# 0.018543f
C42990 a_13661_43548# a_6171_45002# 0.032575f
C42991 a_n2293_46634# a_327_44734# 0.024588f
C42992 a_13925_46122# a_14180_46482# 0.056391f
C42993 a_13759_46122# a_14371_46494# 3.82e-19
C42994 a_n971_45724# a_n2129_44697# 0.017407f
C42995 a_n2497_47436# a_2779_44458# 0.034441f
C42996 a_1138_42852# a_n1099_45572# 3.41e-20
C42997 a_3483_46348# a_n2661_45546# 0.163728f
C42998 a_n2661_46634# a_2382_45260# 2.63e-21
C42999 a_n881_46662# a_15415_45028# 3.95e-20
C43000 a_3524_46660# a_2437_43646# 1.78e-20
C43001 a_n1925_46634# a_n143_45144# 1.28e-21
C43002 a_n1853_46287# a_n23_45546# 7.5e-20
C43003 a_9290_44172# a_13259_45724# 0.272297f
C43004 a_12891_46348# a_13017_45260# 0.210934f
C43005 a_768_44030# a_11787_45002# 3.39e-21
C43006 a_5934_30871# a_9803_42558# 0.001422f
C43007 a_4190_30871# C1_N_btm 7.67e-20
C43008 a_14097_32519# a_22775_42308# 0.001341f
C43009 a_6171_42473# a_5742_30871# 1.16e-20
C43010 a_8337_42558# a_8325_42308# 0.01416f
C43011 a_n913_45002# a_19164_43230# 8.4e-21
C43012 a_n2017_45002# a_20922_43172# 1.61e-20
C43013 a_5883_43914# a_7112_43396# 2.7e-20
C43014 a_n699_43396# a_2813_43396# 0.001609f
C43015 a_21076_30879# a_22609_37990# 1.29e-20
C43016 a_13259_45724# a_21887_42336# 6.84e-19
C43017 a_n356_44636# a_4093_43548# 1.07e-21
C43018 a_15227_46910# VDD 0.229766f
C43019 a_20512_43084# a_19862_44208# 0.023947f
C43020 a_3422_30871# a_11341_43940# 0.030182f
C43021 en_comp a_18249_42858# 8.38e-21
C43022 a_3232_43370# a_10796_42968# 1.9e-20
C43023 a_5263_45724# a_5907_45546# 0.001537f
C43024 a_4185_45028# a_6171_45002# 2.76e-20
C43025 a_2324_44458# a_n2661_45010# 0.001752f
C43026 a_4419_46090# a_3232_43370# 4.56e-21
C43027 a_2711_45572# a_6511_45714# 0.04109f
C43028 a_13661_43548# a_14673_44172# 0.36897f
C43029 a_5164_46348# a_5111_44636# 0.024532f
C43030 a_5204_45822# a_5147_45002# 3.69e-19
C43031 a_3483_46348# a_5205_44484# 0.065176f
C43032 a_8270_45546# a_n2661_44458# 0.019483f
C43033 a_10903_43370# en_comp 4.34e-21
C43034 a_12549_44172# a_18588_44850# 1.05e-20
C43035 a_19553_46090# a_3357_43084# 4.81e-21
C43036 a_13059_46348# a_13711_45394# 6.86e-19
C43037 a_n443_46116# a_n2661_42282# 2.25e-20
C43038 SMPL_ON_N a_19237_31679# 0.029331f
C43039 a_19466_46812# a_18494_42460# 1.2e-19
C43040 a_19692_46634# a_18184_42460# 1.68e-19
C43041 a_3090_45724# a_11691_44458# 0.245063f
C43042 a_9569_46155# a_413_45260# 1.76e-20
C43043 a_15227_44166# a_21005_45260# 3.8e-19
C43044 a_5932_42308# C0_P_btm 0.015561f
C43045 a_6151_47436# a_15673_47210# 0.002744f
C43046 a_11031_47542# a_n1435_47204# 2.39e-19
C43047 a_n4064_39072# a_n2302_38778# 2.59e-20
C43048 a_n2302_39072# a_n4064_38528# 2.59e-20
C43049 a_n815_47178# a_n310_47570# 9.52e-19
C43050 a_5934_30871# C7_P_btm 0.007575f
C43051 a_6123_31319# C5_P_btm 0.022099f
C43052 a_2713_42308# VDD 0.208275f
C43053 a_n1741_47186# a_2487_47570# 2.13e-19
C43054 a_n1630_35242# VIN_N 0.040646f
C43055 a_n2293_42834# a_6171_42473# 2.63e-20
C43056 a_2957_45546# VDD 0.192471f
C43057 a_10949_43914# a_10341_43396# 4.22e-20
C43058 a_10807_43548# a_9885_43646# 1.34e-20
C43059 a_1467_44172# a_743_42282# 3.61e-22
C43060 a_310_45028# DATA[0] 1.08e-20
C43061 a_19319_43548# a_n97_42460# 0.029676f
C43062 a_9313_44734# a_21195_42852# 0.02195f
C43063 a_12861_44030# a_16759_43396# 2.75e-20
C43064 a_4646_46812# a_7499_43940# 0.002542f
C43065 a_11525_45546# a_11963_45334# 2.67e-19
C43066 a_11322_45546# a_13017_45260# 0.003434f
C43067 a_13259_45724# a_17896_45144# 9.29e-19
C43068 a_n1613_43370# a_8147_43396# 3.58e-19
C43069 a_16327_47482# a_15781_43660# 7.49e-21
C43070 a_n2497_47436# a_n13_43084# 1.74e-20
C43071 a_n1151_42308# a_743_42282# 1.08e-19
C43072 a_n23_45546# a_n2661_43370# 3.29e-20
C43073 a_11823_42460# a_8953_45002# 1.65e-20
C43074 a_3483_46348# a_17061_44734# 0.009179f
C43075 a_12465_44636# a_13667_43396# 2.31e-21
C43076 a_2063_45854# a_4361_42308# 1.32e-20
C43077 a_18596_45572# a_18787_45572# 4.61e-19
C43078 a_19431_45546# a_20107_45572# 0.001119f
C43079 a_3090_45724# a_8333_44056# 0.001679f
C43080 a_11415_45002# a_22315_44484# 0.001541f
C43081 a_9290_44172# a_n2661_43922# 0.029391f
C43082 a_10193_42453# a_9482_43914# 0.029531f
C43083 a_11652_45724# a_11787_45002# 0.077604f
C43084 a_n743_46660# a_645_46660# 0.002128f
C43085 a_22521_40055# VDD 1.04757f
C43086 a_19864_35138# a_21589_35634# 0.150796f
C43087 a_4883_46098# a_11735_46660# 2.67e-19
C43088 a_10227_46804# a_15368_46634# 0.003141f
C43089 a_18479_47436# a_3090_45724# 1.24e-20
C43090 a_33_46660# a_491_47026# 0.027606f
C43091 a_n1925_46634# a_n2661_46098# 0.059432f
C43092 a_n2661_46634# a_3524_46660# 0.0105f
C43093 a_n2293_46634# a_3177_46902# 1.62e-20
C43094 a_8128_46384# a_8145_46902# 0.012246f
C43095 a_n881_46662# a_9863_46634# 0.001329f
C43096 a_1123_46634# a_2107_46812# 0.002783f
C43097 a_5807_45002# a_4817_46660# 2.58e-19
C43098 a_16327_47482# a_15227_44166# 0.239667f
C43099 EN_VIN_BSTR_P C5_P_btm 0.115337f
C43100 a_3815_47204# a_765_45546# 0.003873f
C43101 a_n97_42460# a_16795_42852# 0.126591f
C43102 a_20974_43370# a_21195_42852# 1.06e-20
C43103 a_21381_43940# a_22165_42308# 1.75e-19
C43104 a_3905_42865# a_3823_42558# 1.35e-19
C43105 a_n2661_42282# a_n4318_37592# 0.03806f
C43106 a_16409_43396# a_16867_43762# 0.027606f
C43107 a_9482_43914# VDD 1.75061f
C43108 a_17324_43396# a_15743_43084# 0.050725f
C43109 a_18429_43548# a_18783_43370# 0.001885f
C43110 a_10341_43396# a_19095_43396# 0.004123f
C43111 a_3626_43646# a_7765_42852# 3.92e-20
C43112 a_2982_43646# a_8605_42826# 2.81e-20
C43113 a_14955_43396# a_4361_42308# 3.74e-21
C43114 a_11967_42832# a_15890_42674# 0.001386f
C43115 a_3090_45724# a_4190_30871# 1.55e-21
C43116 a_526_44458# a_2253_43940# 9.54e-20
C43117 a_13556_45296# a_13711_45394# 0.005081f
C43118 a_13017_45260# a_15060_45348# 7e-21
C43119 a_n2017_45002# a_n2661_44458# 0.034362f
C43120 a_n2109_45247# a_n2433_44484# 1.13e-19
C43121 a_3357_43084# a_4223_44672# 0.029613f
C43122 a_8049_45260# a_22959_43948# 1.04e-19
C43123 a_1823_45246# a_3539_42460# 0.678673f
C43124 a_n2293_45010# a_n2129_44697# 0.021404f
C43125 a_n2661_45010# a_n1699_44726# 0.04137f
C43126 a_13507_46334# a_14097_32519# 0.001207f
C43127 a_18691_45572# a_18989_43940# 1.88e-19
C43128 a_18799_45938# a_18248_44752# 5.06e-22
C43129 a_n357_42282# a_7542_44172# 2.72e-19
C43130 a_n443_42852# a_453_43940# 0.005083f
C43131 a_n237_47217# a_5907_45546# 1.7e-19
C43132 a_n971_45724# a_6472_45840# 5.6e-19
C43133 a_3877_44458# a_5068_46348# 1.58e-19
C43134 a_n1151_42308# a_2277_45546# 1.18e-22
C43135 a_3633_46660# a_1823_45246# 6.58e-20
C43136 a_8128_46384# a_5066_45546# 0.032968f
C43137 a_n1435_47204# a_n2293_45546# 1.57e-19
C43138 a_14976_45028# a_765_45546# 3.1e-19
C43139 a_4883_46098# a_14537_46482# 1.2e-19
C43140 a_21588_30879# a_22223_46124# 1.77e-19
C43141 a_20916_46384# a_10809_44734# 0.038071f
C43142 a_2905_45572# a_2307_45899# 9.36e-20
C43143 a_584_46384# a_603_45572# 3.31e-19
C43144 a_4646_46812# a_4704_46090# 0.01107f
C43145 a_13507_46334# a_15194_46482# 2.67e-19
C43146 a_18597_46090# a_19240_46482# 0.025784f
C43147 a_n743_46660# a_17715_44484# 0.01357f
C43148 a_3090_45724# a_17829_46910# 1.43e-19
C43149 a_3422_30871# C1_P_btm 7.67e-20
C43150 a_19164_43230# a_20922_43172# 8.1e-20
C43151 a_3626_43646# a_13657_42308# 0.00116f
C43152 a_20159_44458# VDD 0.345429f
C43153 a_7871_42858# a_9061_43230# 2.56e-19
C43154 a_13467_32519# a_20256_42852# 2.92e-20
C43155 a_13678_32519# a_22400_42852# 0.035124f
C43156 a_16979_44734# a_17767_44458# 0.011457f
C43157 a_14539_43914# a_17970_44736# 2.85e-19
C43158 a_11823_42460# a_3626_43646# 0.011402f
C43159 a_375_42282# a_453_43940# 0.021162f
C43160 a_11827_44484# a_10809_44484# 2.9e-20
C43161 a_n357_42282# a_16977_43638# 6.48e-19
C43162 a_13259_45724# a_13467_32519# 0.030863f
C43163 a_17715_44484# a_17701_42308# 0.002546f
C43164 a_n2312_38680# a_n2946_39866# 3.47e-20
C43165 a_n2442_46660# a_n2860_39866# 6.14e-19
C43166 a_17613_45144# a_17517_44484# 1.32e-20
C43167 a_1307_43914# a_2479_44172# 0.300587f
C43168 a_626_44172# a_1467_44172# 4.19e-19
C43169 a_7499_43078# a_6547_43396# 1.37e-19
C43170 a_3537_45260# a_n2661_42282# 0.105917f
C43171 a_n443_42852# a_8873_43396# 8.24e-20
C43172 a_526_44458# a_7871_42858# 0.031818f
C43173 a_n1059_45260# a_18326_43940# 7.46e-21
C43174 a_n2017_45002# a_18451_43940# 4.02e-22
C43175 a_11691_44458# a_14815_43914# 0.018499f
C43176 w_11334_34010# C0_dummy_N_btm 3.87e-21
C43177 a_10903_43370# a_2324_44458# 0.038342f
C43178 a_1138_42852# a_n1925_42282# 1.19e-20
C43179 a_22959_46660# a_8049_45260# 2.87e-20
C43180 a_13759_46122# a_14493_46090# 0.053479f
C43181 a_n1151_42308# a_626_44172# 3.18e-21
C43182 a_3090_45724# a_n443_42852# 0.269331f
C43183 a_19321_45002# a_18175_45572# 0.01259f
C43184 a_19123_46287# a_19240_46482# 0.157972f
C43185 a_13661_43548# a_18909_45814# 0.006912f
C43186 a_5807_45002# a_18691_45572# 0.001465f
C43187 a_13747_46662# a_18341_45572# 0.554429f
C43188 a_4842_47570# a_2437_43646# 8.98e-19
C43189 a_19386_47436# a_413_45260# 1.03e-19
C43190 a_1823_45246# a_526_44458# 1.93329f
C43191 a_472_46348# a_1337_46116# 2.04e-19
C43192 a_8667_46634# a_7499_43078# 1.51e-19
C43193 a_8492_46660# a_8568_45546# 2.74e-20
C43194 a_n743_46660# a_15861_45028# 0.005332f
C43195 a_9313_45822# a_8953_45002# 0.001732f
C43196 a_765_45546# a_18051_46116# 0.006713f
C43197 a_22959_42860# a_22775_42308# 0.019713f
C43198 a_1576_42282# a_1755_42282# 0.168925f
C43199 a_1184_42692# a_1606_42308# 0.125247f
C43200 a_n3674_37592# a_n39_42308# 0.003612f
C43201 a_13291_42460# a_13070_42354# 0.155164f
C43202 a_6031_43396# VDD 0.47547f
C43203 a_n784_42308# a_2713_42308# 2.26e-20
C43204 a_n357_42282# a_n1630_35242# 0.086672f
C43205 a_22959_44484# a_19237_31679# 0.155744f
C43206 en_comp a_5649_42852# 2.63e-19
C43207 a_n2661_45010# a_n2157_42858# 4.56e-21
C43208 a_n755_45592# a_564_42282# 0.036154f
C43209 a_n863_45724# a_1149_42558# 0.002168f
C43210 a_9313_44734# a_15493_43396# 0.001749f
C43211 a_n2293_43922# a_10949_43914# 0.008394f
C43212 a_n2661_42834# a_11750_44172# 0.006203f
C43213 a_n2661_43922# a_10807_43548# 2.2e-19
C43214 a_n2661_43370# a_7287_43370# 3.73e-21
C43215 a_7715_46873# VDD 0.414019f
C43216 a_n2661_45546# a_n357_42282# 0.044767f
C43217 a_n1079_45724# a_n452_45724# 6.61e-19
C43218 a_n2293_46634# a_4223_44672# 3.24e-21
C43219 a_8492_46660# a_n2661_43370# 1.86e-21
C43220 a_14976_45028# a_16751_45260# 1.25e-20
C43221 a_n2497_47436# a_644_44056# 0.016428f
C43222 a_11415_45002# a_22959_45572# 0.001334f
C43223 a_22591_46660# a_19963_31679# 1.81e-20
C43224 a_12549_44172# a_18443_44721# 1.36e-19
C43225 a_12741_44636# a_3357_43084# 0.036536f
C43226 a_20820_30879# a_22591_45572# 9.76e-21
C43227 a_10227_46804# a_15146_44811# 6.31e-20
C43228 a_n2293_45546# a_380_45546# 4.68e-20
C43229 a_n2956_38216# a_n1099_45572# 3.28e-19
C43230 a_13661_43548# a_12607_44458# 0.00102f
C43231 a_15015_46420# a_15037_45618# 0.001025f
C43232 a_2324_44458# a_12016_45572# 2.57e-19
C43233 a_15227_44166# a_14537_43396# 0.105881f
C43234 a_20202_43084# a_20447_31679# 8.03e-21
C43235 a_12861_44030# a_17517_44484# 0.069119f
C43236 a_n1630_35242# CAL_N 1.66e-19
C43237 COMP_P a_22821_38993# 2.95e-19
C43238 a_n237_47217# a_n23_47502# 0.056864f
C43239 a_n746_45260# a_n785_47204# 0.198992f
C43240 a_n971_45724# a_327_47204# 0.075444f
C43241 a_n1741_47186# a_584_46384# 0.021978f
C43242 a_n2109_47186# a_2553_47502# 0.04572f
C43243 a_3065_45002# a_3905_42558# 0.044632f
C43244 a_3422_30871# a_10341_43396# 0.029183f
C43245 a_11967_42832# a_16547_43609# 0.176385f
C43246 a_n356_44636# a_685_42968# 3.75e-19
C43247 a_n2017_45002# a_8325_42308# 0.009217f
C43248 a_3499_42826# a_4235_43370# 4.6e-20
C43249 a_19862_44208# a_21381_43940# 0.113704f
C43250 a_20692_30879# a_22459_39145# 3e-20
C43251 a_15493_43396# a_20974_43370# 1.15e-20
C43252 a_18479_45785# a_17303_42282# 1.31e-20
C43253 a_n357_42282# a_5205_44484# 3.84e-20
C43254 a_6945_45028# a_11827_44484# 8.14e-20
C43255 a_1609_45822# a_1667_45002# 0.001741f
C43256 a_15225_45822# a_15765_45572# 2.89e-20
C43257 a_19692_46634# a_20362_44736# 3.19e-21
C43258 a_8199_44636# a_5343_44458# 7.94e-19
C43259 a_n443_42852# a_2274_45254# 1.98e-21
C43260 a_15227_44166# a_20835_44721# 4.95e-20
C43261 a_n2293_46634# a_15493_43940# 0.003183f
C43262 a_13661_43548# a_14761_44260# 5.06e-19
C43263 a_768_44030# a_3992_43940# 0.006422f
C43264 a_8049_45260# a_8137_45348# 2.64e-19
C43265 a_3483_46348# a_13076_44458# 4.08e-21
C43266 a_n2302_38778# VDD 0.35162f
C43267 a_5700_37509# VDAC_N 1.09421f
C43268 a_n1741_47186# a_11901_46660# 0.034005f
C43269 a_n971_45724# a_8846_46660# 5.95e-19
C43270 a_n4064_39072# VCM 0.035838f
C43271 a_6491_46660# a_7715_46873# 1.43e-20
C43272 a_n1151_42308# a_6755_46942# 0.142929f
C43273 a_6151_47436# a_8145_46902# 0.178565f
C43274 a_6545_47178# a_7577_46660# 3.97e-20
C43275 a_4338_37500# VDAC_P 0.037246f
C43276 a_5088_37509# a_8912_37509# 16.1906f
C43277 a_3726_37500# a_11206_38545# 0.11542f
C43278 a_7754_38470# CAL_P 1.73e-19
C43279 a_11309_47204# a_5807_45002# 0.032739f
C43280 a_n1435_47204# a_5732_46660# 1.28e-20
C43281 a_19328_44172# a_19339_43156# 1.37e-19
C43282 a_15493_43396# a_18599_43230# 5.54e-20
C43283 a_n4318_40392# a_n4315_30879# 0.151169f
C43284 a_3422_30871# a_20356_42852# 3.72e-19
C43285 a_5891_43370# a_10545_42558# 1.64e-20
C43286 a_20512_43084# a_20573_43172# 0.00112f
C43287 a_11341_43940# a_16414_43172# 3.69e-21
C43288 a_8685_43396# a_14358_43442# 0.002184f
C43289 a_n356_44636# a_14113_42308# 0.019853f
C43290 a_2982_43646# a_18783_43370# 4.48e-21
C43291 a_n97_42460# a_19095_43396# 0.003217f
C43292 a_20623_45572# VDD 0.200978f
C43293 a_9396_43370# a_9885_43396# 4.89e-20
C43294 a_1823_45246# a_3353_43940# 4.96e-20
C43295 a_6171_45002# a_13159_45002# 0.012283f
C43296 a_8192_45572# a_5343_44458# 6.07e-21
C43297 a_2680_45002# a_1307_43914# 9.4e-20
C43298 a_7705_45326# a_8953_45002# 1.82e-20
C43299 a_3357_43084# a_n2293_42834# 0.045124f
C43300 a_8016_46348# a_10555_44260# 0.007104f
C43301 a_8199_44636# a_9801_44260# 6.23e-19
C43302 a_13249_42308# a_13720_44458# 1.19e-19
C43303 a_n443_42852# a_14815_43914# 8.61e-20
C43304 a_11415_45002# a_19319_43548# 2.49e-20
C43305 a_327_44734# a_626_44172# 0.120093f
C43306 a_18341_45572# a_18911_45144# 0.006584f
C43307 a_18479_45785# a_19778_44110# 0.009f
C43308 a_13507_46334# a_22959_42860# 0.004407f
C43309 a_n2442_46660# a_n4318_38680# 0.023781f
C43310 a_768_44030# a_9127_43156# 1.24e-19
C43311 a_8270_45546# a_9145_43396# 0.02247f
C43312 a_3483_46348# a_15301_44260# 6.81e-19
C43313 a_7499_43078# a_n356_44636# 4.62e-19
C43314 a_n2438_43548# a_n1991_42858# 9.37e-19
C43315 a_3090_45724# a_6655_43762# 0.002552f
C43316 a_n2293_45010# a_45_45144# 3.59e-21
C43317 a_2324_44458# a_14955_43940# 0.029449f
C43318 a_4883_46098# a_2324_44458# 0.074521f
C43319 a_18479_47436# a_20075_46420# 0.061108f
C43320 a_16023_47582# a_10809_44734# 5.41e-20
C43321 a_n2840_46634# a_n2840_46090# 0.026152f
C43322 a_6151_47436# a_5066_45546# 0.019067f
C43323 a_n2293_46634# a_12741_44636# 3.52e-21
C43324 a_11453_44696# a_13759_46122# 9.57e-21
C43325 a_13507_46334# a_17583_46090# 0.004113f
C43326 a_19787_47423# a_18819_46122# 1.83e-20
C43327 a_10227_46804# a_20708_46348# 0.001063f
C43328 a_16588_47582# a_6945_45028# 0.011591f
C43329 a_n881_46662# a_6165_46155# 2.6e-19
C43330 a_n1613_43370# a_6419_46155# 0.013016f
C43331 a_n1151_42308# a_8049_45260# 0.075767f
C43332 a_12891_46348# a_3483_46348# 0.053153f
C43333 a_768_44030# a_2804_46116# 0.001471f
C43334 a_3524_46660# a_765_45546# 0.002975f
C43335 a_6755_46942# a_14084_46812# 0.052304f
C43336 a_19386_47436# a_18985_46122# 6.11e-19
C43337 a_18597_46090# a_19553_46090# 0.021441f
C43338 a_12465_44636# a_15015_46420# 8.41e-21
C43339 a_7765_42852# a_8037_42858# 0.309282f
C43340 a_7871_42858# a_8605_42826# 0.06628f
C43341 a_4361_42308# a_n2293_42282# 2.71e-21
C43342 a_15095_43370# a_14853_42852# 6.13e-21
C43343 a_14579_43548# a_16245_42852# 6.32e-20
C43344 a_15493_43940# a_20107_42308# 7.88e-22
C43345 a_13887_32519# a_21195_42852# 9.75e-21
C43346 a_4093_43548# a_3823_42558# 1.14e-20
C43347 a_3080_42308# a_2713_42308# 0.004874f
C43348 a_14021_43940# a_17303_42282# 3.16e-21
C43349 a_13678_32519# a_22223_42860# 0.002285f
C43350 a_5649_42852# a_22165_42308# 0.077779f
C43351 a_n1809_44850# VDD 0.132538f
C43352 a_n2661_43370# a_n23_44458# 9.21e-19
C43353 a_n2840_44458# a_n2661_44458# 0.179135f
C43354 a_n2293_45010# a_n2472_43914# 1.49e-19
C43355 a_n2661_45010# a_n1761_44111# 8.36e-20
C43356 a_17715_44484# a_4361_42308# 6.15e-21
C43357 a_2437_43646# a_453_43940# 1.7e-19
C43358 a_12741_44636# a_5342_30871# 1.14e-22
C43359 a_n2293_46634# a_5742_30871# 2.68e-19
C43360 a_3090_45724# a_14635_42282# 0.007468f
C43361 a_n755_45592# a_n1557_42282# 0.199254f
C43362 a_5837_45028# a_5891_43370# 6.5e-21
C43363 a_6171_45002# a_11967_42832# 5.32e-19
C43364 a_8696_44636# a_12429_44172# 2.76e-20
C43365 a_16115_45572# a_15682_43940# 2.15e-19
C43366 a_n971_45724# a_n745_45366# 1.48e-20
C43367 a_n746_45260# a_n913_45002# 0.051081f
C43368 a_16327_47482# a_16377_45572# 0.001903f
C43369 a_n2293_46634# a_3260_45572# 3.64e-19
C43370 a_1823_45246# a_2521_46116# 5.42e-19
C43371 a_2202_46116# a_167_45260# 0.159883f
C43372 a_13507_46334# a_8696_44636# 3.72e-19
C43373 a_n743_46660# a_3775_45552# 3.52e-20
C43374 a_12549_44172# a_13249_42308# 0.066967f
C43375 a_768_44030# a_13904_45546# 0.005947f
C43376 a_18285_46348# a_19335_46494# 1.12e-20
C43377 a_19123_46287# a_19553_46090# 1.56e-20
C43378 SMPL_ON_P a_n967_45348# 5.24e-20
C43379 a_3785_47178# a_2437_43646# 0.015875f
C43380 a_5807_45002# a_10490_45724# 4.75e-23
C43381 a_13747_46662# a_10193_42453# 7.93e-21
C43382 a_11813_46116# a_11387_46482# 1.25e-20
C43383 a_16751_46987# a_10809_44734# 4.31e-19
C43384 a_n2497_47436# a_n37_45144# 2.82e-20
C43385 a_2107_46812# a_4099_45572# 4.87e-20
C43386 a_11599_46634# a_18341_45572# 0.588263f
C43387 a_6671_43940# VDD 0.227011f
C43388 a_5342_30871# a_5742_30871# 0.031909f
C43389 a_13635_43156# a_13575_42558# 0.00691f
C43390 a_21588_30879# C5_N_btm 5.07e-20
C43391 a_14673_44172# a_11967_42832# 3.97e-20
C43392 a_17517_44484# a_17325_44484# 1.97e-19
C43393 a_5343_44458# a_8018_44260# 0.003899f
C43394 a_5111_44636# a_6197_43396# 0.025934f
C43395 a_4185_45028# a_15959_42545# 1.27e-19
C43396 a_n2017_45002# a_9145_43396# 2.64e-19
C43397 a_13747_46662# VDD 3.70214f
C43398 a_5807_45002# START 1.22e-19
C43399 a_5691_45260# a_6031_43396# 1.62e-21
C43400 a_5883_43914# a_6101_44260# 0.001046f
C43401 a_4223_44672# a_9672_43914# 4.35e-21
C43402 a_3537_45260# a_7112_43396# 0.046531f
C43403 a_13661_43548# RST_Z 1.9e-20
C43404 a_10193_42453# a_10796_42968# 0.015009f
C43405 a_768_44030# CLK 1.44e-19
C43406 a_n357_42282# a_3863_42891# 3.29e-19
C43407 a_n755_45592# a_8483_43230# 2.93e-19
C43408 a_526_44458# a_1184_42692# 6.23e-19
C43409 a_n1925_42282# a_1576_42282# 1.31e-19
C43410 a_19778_44110# a_14021_43940# 4.06e-19
C43411 a_20202_43084# a_21887_42336# 0.082645f
C43412 a_20193_45348# a_22959_43948# 2.96e-19
C43413 a_9290_44172# a_10545_42558# 6.22e-19
C43414 a_n443_42852# a_945_42968# 9.8e-19
C43415 a_3090_45724# a_2437_43646# 1.6e-19
C43416 a_526_44458# a_n2293_45546# 1.47e-19
C43417 a_n1925_42282# a_n2956_38216# 3.5e-20
C43418 a_n971_45724# a_3363_44484# 4.12e-21
C43419 a_n746_45260# a_556_44484# 0.045671f
C43420 a_3483_46348# a_11322_45546# 0.554731f
C43421 a_8270_45546# a_n1059_45260# 5.56e-20
C43422 a_19692_46634# a_21363_45546# 8.99e-19
C43423 a_19466_46812# a_21188_45572# 4.5e-20
C43424 a_15015_46420# a_2711_45572# 1.15e-20
C43425 a_6969_46634# a_413_45260# 2.65e-20
C43426 a_15227_44166# a_20731_45938# 3.88e-19
C43427 a_13607_46688# a_3357_43084# 1.82e-20
C43428 a_n2293_46634# a_n2293_42834# 0.027042f
C43429 a_5937_45572# a_4808_45572# 6.9e-20
C43430 a_7411_46660# a_3232_43370# 8.54e-22
C43431 a_5257_43370# a_6171_45002# 3.04e-19
C43432 a_12549_44172# a_17613_45144# 7.44e-21
C43433 a_2063_45854# a_5891_43370# 1.78e-19
C43434 a_12861_44030# a_13720_44458# 4.84e-19
C43435 a_6123_31319# a_n4209_39590# 9.76e-22
C43436 a_5342_30871# C0_dummy_P_btm 1.91e-20
C43437 a_n4318_38216# a_n3690_38304# 7.76e-19
C43438 a_5534_30871# C0_N_btm 8.49e-20
C43439 a_15803_42450# a_4958_30871# 0.093396f
C43440 a_15764_42576# a_17303_42282# 1.02e-19
C43441 a_15959_42545# a_16269_42308# 0.013793f
C43442 a_15890_42674# a_16197_42308# 3.69e-19
C43443 a_10723_42308# a_7174_31319# 9.76e-21
C43444 a_n3674_38216# a_n4334_38304# 0.059852f
C43445 a_10796_42968# VDD 0.270235f
C43446 a_5663_43940# a_5829_43940# 0.143754f
C43447 a_11823_42460# a_13921_42308# 3.14e-20
C43448 a_10193_42453# a_4958_30871# 0.108497f
C43449 a_4419_46090# VDD 0.664887f
C43450 a_3422_30871# a_n97_42460# 3.53e-20
C43451 a_17973_43940# a_19328_44172# 4.29e-20
C43452 a_17737_43940# a_15493_43396# 1.12e-19
C43453 a_4185_45028# RST_Z 0.005781f
C43454 a_9313_44734# a_10695_43548# 2.41e-19
C43455 a_n356_44636# a_15781_43660# 6.74e-21
C43456 a_10729_43914# a_11341_43940# 0.243062f
C43457 a_18079_43940# a_18451_43940# 9.65e-20
C43458 a_18597_46090# a_15493_43940# 0.024181f
C43459 a_11453_44696# a_18079_43940# 1.52e-19
C43460 a_8199_44636# a_8560_45348# 0.03862f
C43461 a_5497_46414# a_n2661_43370# 4.83e-21
C43462 a_n1613_43370# a_n2661_42282# 0.017743f
C43463 a_11962_45724# a_13527_45546# 1.48e-19
C43464 a_7499_43078# a_8697_45822# 0.038073f
C43465 a_2711_45572# a_16333_45814# 9.94e-19
C43466 a_8568_45546# a_9241_45822# 7.63e-21
C43467 a_n2438_43548# a_n1331_43914# 7.33e-21
C43468 a_15227_44166# a_n356_44636# 8.76e-20
C43469 a_3090_45724# a_4181_44734# 0.003724f
C43470 a_12741_44636# a_16237_45028# 0.00167f
C43471 a_11823_42460# a_12791_45546# 0.030093f
C43472 a_5066_45546# a_5111_44636# 7.73e-19
C43473 a_n2497_47436# a_104_43370# 0.001117f
C43474 a_n971_45724# a_n2433_43396# 8.25e-19
C43475 a_n1151_42308# a_n2442_46660# 6.91e-20
C43476 a_3785_47178# a_n2661_46634# 7.96e-20
C43477 a_7227_47204# a_5807_45002# 1.09e-19
C43478 a_12861_44030# a_12549_44172# 1.20253f
C43479 a_13717_47436# a_768_44030# 0.029731f
C43480 a_13487_47204# a_12891_46348# 1.6e-19
C43481 a_7174_31319# C1_P_btm 5.34e-20
C43482 a_n2109_47186# a_1799_45572# 1.89e-19
C43483 a_n2288_47178# a_n2661_46098# 2.56e-20
C43484 a_22731_47423# a_11453_44696# 0.048111f
C43485 a_584_46384# a_n743_46660# 0.42078f
C43486 a_2124_47436# a_n2438_43548# 3.55e-19
C43487 a_4958_30871# VDD 1.06745f
C43488 VDAC_Pi a_3754_39466# 0.308867f
C43489 a_n4209_38216# a_n4209_37414# 0.041723f
C43490 a_2553_47502# a_n1925_46634# 4.04e-20
C43491 a_n971_45724# a_1983_46706# 0.004287f
C43492 a_327_47204# a_601_46902# 0.003002f
C43493 a_n785_47204# a_383_46660# 0.001568f
C43494 a_n237_47217# a_948_46660# 6.91e-20
C43495 a_16023_47582# a_n881_46662# 1.58e-20
C43496 a_20512_43084# a_21671_42860# 2.28e-19
C43497 a_4223_44672# a_5755_42308# 7.11e-21
C43498 a_3080_42308# a_6031_43396# 9.6e-22
C43499 a_4699_43561# a_6293_42852# 5.22e-21
C43500 a_2982_43646# a_3626_43646# 6.553431f
C43501 a_766_43646# a_648_43396# 1.98e-20
C43502 a_n1557_42282# a_548_43396# 0.005988f
C43503 a_20623_43914# a_4361_42308# 3.31e-21
C43504 a_11341_43940# a_21487_43396# 0.005254f
C43505 a_19862_44208# a_5649_42852# 1.34e-20
C43506 a_14815_43914# a_14635_42282# 1.04e-19
C43507 a_15493_43940# a_743_42282# 5.64e-20
C43508 a_11415_45002# a_10949_43914# 1.43e-20
C43509 a_2437_43646# a_2274_45254# 0.01398f
C43510 a_n2293_45010# a_n745_45366# 5.55e-20
C43511 a_n2017_45002# a_n1059_45260# 6.27837f
C43512 a_n2472_45002# a_n2810_45028# 0.002586f
C43513 a_3090_45724# a_11257_43940# 6.36e-20
C43514 a_4099_45572# a_n2661_44458# 2.29e-20
C43515 a_3357_43084# a_413_45260# 7.24598f
C43516 a_12549_44172# a_19700_43370# 7.13e-19
C43517 a_n443_42852# a_4743_44484# 1.62e-20
C43518 a_4646_46812# a_6031_43396# 0.849684f
C43519 a_n2293_46098# a_n2661_42282# 0.182071f
C43520 a_n2661_45010# a_n2956_37592# 0.163638f
C43521 a_n2840_45002# en_comp 8.04e-20
C43522 a_13059_46348# a_13829_44260# 0.002505f
C43523 a_n2293_46634# a_10849_43646# 0.001727f
C43524 a_13661_43548# a_16243_43396# 0.001958f
C43525 VDD VCM 1.51164f
C43526 a_4651_46660# a_7411_46660# 1.59e-21
C43527 a_19594_46812# a_19333_46634# 0.060858f
C43528 a_5807_45002# a_12156_46660# 0.002125f
C43529 a_768_44030# a_14035_46660# 0.270355f
C43530 a_12549_44172# a_14180_46812# 0.023435f
C43531 a_10227_46804# a_21542_46660# 0.002879f
C43532 a_5385_46902# a_5263_46660# 3.16e-19
C43533 a_4955_46873# a_5257_43370# 2.43e-21
C43534 a_2063_45854# a_9290_44172# 0.655982f
C43535 a_n2661_46634# a_3090_45724# 6.05e-20
C43536 DATA[3] DATA[4] 0.001426f
C43537 a_n1435_47204# a_1138_42852# 1.06e-20
C43538 a_4791_45118# a_6419_46155# 0.371259f
C43539 a_5129_47502# a_5204_45822# 2.88e-19
C43540 a_n1151_42308# a_8953_45546# 0.120628f
C43541 a_19321_45002# a_19466_46812# 0.130025f
C43542 a_n743_46660# a_11901_46660# 9.04e-20
C43543 a_3877_44458# a_7577_46660# 2.44e-19
C43544 a_4646_46812# a_7715_46873# 0.058457f
C43545 a_13507_46334# a_20885_46660# 4.28e-19
C43546 a_18597_46090# a_12741_44636# 0.267775f
C43547 a_6293_42852# a_6101_43172# 9.07e-19
C43548 a_n97_42460# a_18504_43218# 0.002932f
C43549 a_18911_45144# VDD 0.218047f
C43550 a_12281_43396# a_5534_30871# 0.012136f
C43551 a_14209_32519# a_17364_32525# 0.056697f
C43552 a_3422_30871# a_n3420_39616# 0.005543f
C43553 a_10341_43396# a_16414_43172# 8.63e-20
C43554 a_3090_45724# a_14543_43071# 0.003291f
C43555 a_768_44030# a_1755_42282# 2.83e-20
C43556 SMPL_ON_P a_n4209_39590# 0.007959f
C43557 a_1307_43914# a_5518_44484# 0.01058f
C43558 a_2711_45572# a_15493_43396# 0.054674f
C43559 a_n2312_39304# a_5934_30871# 5.64e-21
C43560 a_10227_46804# a_13070_42354# 7.16e-20
C43561 a_20202_43084# a_13467_32519# 0.333168f
C43562 a_n2956_39768# a_n4318_38216# 0.023554f
C43563 a_13017_45260# a_12883_44458# 7.59e-19
C43564 a_13159_45002# a_12607_44458# 4.65e-20
C43565 a_1423_45028# a_949_44458# 0.06121f
C43566 a_18909_45814# a_11967_42832# 4.13e-21
C43567 a_9482_43914# a_10057_43914# 0.401746f
C43568 a_n2442_46660# a_n2840_42282# 4.03e-20
C43569 a_4185_45028# a_16243_43396# 8.86e-21
C43570 a_3483_46348# a_16409_43396# 3.88e-19
C43571 a_4883_46098# a_6667_45809# 6.08e-20
C43572 a_11735_46660# a_11387_46155# 1.2e-19
C43573 a_3090_45724# a_8199_44636# 0.030057f
C43574 a_11599_46634# a_10193_42453# 0.100544f
C43575 a_6151_47436# a_6977_45572# 9.54e-19
C43576 a_2063_45854# a_11064_45572# 0.001139f
C43577 a_6545_47178# a_6905_45572# 1.54e-20
C43578 a_19123_46287# a_12741_44636# 3.1e-21
C43579 a_21188_46660# a_21350_47026# 0.006453f
C43580 a_20623_46660# a_20885_46660# 0.001705f
C43581 a_20411_46873# a_11415_45002# 4.84e-20
C43582 a_20273_46660# a_20202_43084# 8.55e-20
C43583 a_20107_46660# a_22591_46660# 3.89e-21
C43584 a_n881_46662# a_n23_45546# 3.9e-19
C43585 a_10150_46912# a_6945_45028# 5.48e-20
C43586 a_5649_42852# a_9803_42558# 6.94e-20
C43587 a_16759_43396# a_17124_42282# 7.27e-19
C43588 a_16137_43396# a_4958_30871# 0.008832f
C43589 a_10341_43396# a_7174_31319# 4.2e-20
C43590 a_1847_42826# a_2903_42308# 4.53e-19
C43591 a_19164_43230# a_19273_43230# 0.007416f
C43592 a_19339_43156# a_19518_43218# 0.007399f
C43593 a_18599_43230# a_18707_42852# 0.057222f
C43594 a_10796_42968# a_n784_42308# 8.64e-21
C43595 a_5755_42852# a_1755_42282# 7.33e-21
C43596 a_743_42282# a_5742_30871# 0.02341f
C43597 a_n755_45592# a_3935_42891# 3.21e-22
C43598 a_n357_42282# a_4520_42826# 0.005592f
C43599 a_19692_46634# a_17303_42282# 6.55e-21
C43600 a_8375_44464# a_n2661_43922# 0.007585f
C43601 a_5891_43370# a_n2661_42834# 0.091553f
C43602 a_11031_47542# DATA[5] 0.006702f
C43603 SMPL_ON_N a_19864_35138# 0.01194f
C43604 a_n443_42852# a_n1736_43218# 5.95e-22
C43605 a_13259_45724# a_16795_42852# 2.94e-19
C43606 a_526_44458# a_5193_42852# 0.058324f
C43607 a_9313_45822# DATA[4] 0.0373f
C43608 a_9482_43914# a_14021_43940# 3.32e-19
C43609 a_5111_44636# a_8415_44056# 0.003443f
C43610 a_14955_47212# RST_Z 1.35e-19
C43611 a_n2661_45010# a_n2267_43396# 2.61e-20
C43612 a_18248_44752# a_18204_44850# 1.46e-19
C43613 a_18287_44626# a_17517_44484# 0.031756f
C43614 a_n1435_47204# DATA[1] 0.037154f
C43615 a_3232_43370# a_5829_43940# 5.72e-19
C43616 a_9067_47204# CLK 1.63e-19
C43617 a_11599_46634# VDD 5.64965f
C43618 a_19553_46090# a_8049_45260# 0.002856f
C43619 a_10903_43370# a_12839_46116# 0.115226f
C43620 a_472_46348# a_n755_45592# 3.56e-20
C43621 a_805_46414# a_n357_42282# 6.63e-19
C43622 a_n2293_46098# a_n310_45899# 7.73e-19
C43623 a_n746_45260# a_n2661_44458# 0.079054f
C43624 a_n971_45724# a_n2433_44484# 4.54e-20
C43625 a_5807_45002# a_6171_45002# 0.193427f
C43626 a_n2438_43548# a_n967_45348# 4.25e-21
C43627 a_n2293_46634# a_413_45260# 0.497204f
C43628 a_13759_46122# a_14180_46482# 0.086708f
C43629 a_n2497_47436# a_949_44458# 0.127971f
C43630 a_1176_45822# a_n1099_45572# 5.28e-20
C43631 a_3147_46376# a_n2661_45546# 6.59e-20
C43632 a_n881_46662# a_14797_45144# 1.1e-19
C43633 a_12861_44030# a_15685_45394# 5.1e-20
C43634 a_3699_46634# a_2437_43646# 5.21e-20
C43635 a_n1853_46287# a_n356_45724# 0.011459f
C43636 a_768_44030# a_10951_45334# 7.27e-21
C43637 a_8515_42308# a_8791_42308# 0.001038f
C43638 a_5934_30871# a_9223_42460# 0.051891f
C43639 a_20753_42852# a_20712_42282# 5.65e-19
C43640 a_4190_30871# C0_N_btm 6.53e-20
C43641 a_n784_42308# a_4958_30871# 0.020733f
C43642 a_22400_42852# a_22775_42308# 0.003696f
C43643 a_5755_42308# a_5742_30871# 2.87e-20
C43644 a_16922_45042# a_17499_43370# 4.92e-21
C43645 a_n2293_42834# a_743_42282# 2.24e-19
C43646 a_n913_45002# a_19339_43156# 3.67e-21
C43647 a_n2017_45002# a_19987_42826# 0.142839f
C43648 a_n1059_45260# a_19164_43230# 8.48e-22
C43649 a_5883_43914# a_7287_43370# 2.97e-19
C43650 a_n1644_44306# a_n1453_44318# 4.61e-19
C43651 a_3600_43914# a_3820_44260# 0.009965f
C43652 a_3905_42865# a_3499_42826# 6.78e-19
C43653 a_3422_30871# a_21115_43940# 1.12e-21
C43654 a_20159_44458# a_14021_43940# 7.12e-20
C43655 a_13259_45724# a_21335_42336# 5.02e-20
C43656 a_n2956_38680# a_n2216_38778# 0.001511f
C43657 en_comp a_17333_42852# 1.3e-21
C43658 a_10933_46660# CLK 0.002047f
C43659 a_3232_43370# a_10835_43094# 2.81e-20
C43660 a_n2312_38680# a_n2293_43922# 3.87e-20
C43661 a_3483_46348# a_6431_45366# 0.002186f
C43662 a_4185_45028# a_3232_43370# 0.018743f
C43663 a_2711_45572# a_6472_45840# 0.049759f
C43664 a_5807_45002# a_14673_44172# 0.001217f
C43665 a_5164_46348# a_5147_45002# 0.060833f
C43666 a_5068_46348# a_5111_44636# 2.11e-19
C43667 a_18985_46122# a_3357_43084# 2.92e-20
C43668 a_13059_46348# a_13490_45394# 4.86e-19
C43669 a_2063_45854# a_10807_43548# 0.094631f
C43670 a_4791_45118# a_n2661_42282# 9.1e-19
C43671 a_3090_45724# a_19113_45348# 0.128103f
C43672 a_15227_44166# a_20567_45036# 2.08e-20
C43673 a_19466_46812# a_18184_42460# 0.006722f
C43674 a_9625_46129# a_413_45260# 4.85e-21
C43675 a_20075_46420# a_2437_43646# 1.37e-20
C43676 a_19692_46634# a_19778_44110# 1.92e-20
C43677 a_10586_45546# a_8696_44636# 1.39e-19
C43678 a_5932_42308# C1_P_btm 0.011049f
C43679 a_6151_47436# a_15811_47375# 1.9e-19
C43680 a_9863_47436# a_n1435_47204# 2.39e-19
C43681 a_9313_45822# a_11459_47204# 0.210847f
C43682 a_n4064_39072# a_n4064_38528# 0.05966f
C43683 a_n815_47178# a_n2312_39304# 8.4e-20
C43684 a_5934_30871# C8_P_btm 1.41e-19
C43685 a_n1630_35242# VIN_P 0.049047f
C43686 a_n784_42308# VCM 0.195503f
C43687 a_6123_31319# C6_P_btm 6.31e-19
C43688 a_2725_42558# VDD 0.005543f
C43689 a_n1741_47186# a_2266_47570# 2.25e-19
C43690 a_n2109_47186# a_2747_46873# 0.087441f
C43691 a_n2293_42834# a_5755_42308# 7.41e-20
C43692 a_1848_45724# VDD 0.100884f
C43693 a_10729_43914# a_10341_43396# 2.83e-20
C43694 a_n913_45002# a_22465_38105# 2.35e-19
C43695 a_17730_32519# a_17364_32525# 0.054843f
C43696 a_19237_31679# a_14209_32519# 0.052426f
C43697 a_n1099_45572# DATA[0] 1.56e-20
C43698 a_9313_44734# a_21356_42826# 0.009873f
C43699 a_584_46384# a_4361_42308# 6.47e-21
C43700 a_12861_44030# a_16977_43638# 5.41e-21
C43701 a_6755_46942# a_15493_43940# 0.001348f
C43702 a_11322_45546# a_11963_45334# 0.028732f
C43703 a_11525_45546# a_11787_45002# 5.53e-19
C43704 a_n2293_46634# a_n2012_43396# 1.17e-21
C43705 a_13259_45724# a_17801_45144# 3.04e-19
C43706 a_n1613_43370# a_7112_43396# 0.245085f
C43707 a_n2497_47436# a_n1076_43230# 2.48e-20
C43708 SMPL_ON_P a_n1853_43023# 8.05e-21
C43709 a_n2438_43548# a_n1917_43396# 2.8e-19
C43710 a_n356_45724# a_n2661_43370# 7.45e-20
C43711 a_16375_45002# a_16237_45028# 0.035582f
C43712 a_11415_45002# a_3422_30871# 0.002932f
C43713 a_9290_44172# a_n2661_42834# 0.046011f
C43714 a_10180_45724# a_9482_43914# 0.001194f
C43715 a_8049_45260# a_4223_44672# 1.63e-20
C43716 a_11652_45724# a_10951_45334# 1.16e-21
C43717 a_16327_47482# a_18834_46812# 3.5e-20
C43718 a_n743_46660# a_479_46660# 0.004337f
C43719 a_n2438_43548# a_1110_47026# 2.49e-19
C43720 a_22780_40945# VDD 1.38e-19
C43721 a_22469_40625# RST_Z 8.08e-20
C43722 a_33_46660# a_288_46660# 0.056391f
C43723 a_n2312_38680# a_n2661_46098# 0.003978f
C43724 a_n1925_46634# a_1799_45572# 0.035794f
C43725 a_n2661_46634# a_3699_46634# 0.009256f
C43726 a_n2293_46634# a_2609_46660# 1.11e-20
C43727 a_8128_46384# a_7577_46660# 0.023306f
C43728 a_6151_47436# a_13059_46348# 1.9e-19
C43729 a_13507_46334# a_11813_46116# 1.34e-19
C43730 a_10227_46804# a_14976_45028# 0.536884f
C43731 a_1123_46634# a_948_46660# 0.234322f
C43732 EN_VIN_BSTR_P C6_P_btm 0.118916f
C43733 a_3785_47178# a_765_45546# 0.004672f
C43734 a_5807_45002# a_4955_46873# 4.29e-20
C43735 a_n97_42460# a_16414_43172# 0.044625f
C43736 a_20974_43370# a_21356_42826# 8.97e-20
C43737 a_21381_43940# a_21671_42860# 0.001657f
C43738 a_16409_43396# a_16664_43396# 0.056391f
C43739 a_13348_45260# VDD 0.083657f
C43740 a_n2661_42282# a_n1736_42282# 3.68e-19
C43741 a_18429_43548# a_18525_43370# 0.419086f
C43742 a_17499_43370# a_15743_43084# 0.049383f
C43743 a_14579_43548# a_5649_42852# 3.24e-21
C43744 a_10341_43396# a_21487_43396# 0.010314f
C43745 a_15095_43370# a_4361_42308# 1.65e-19
C43746 a_11967_42832# a_15959_42545# 6.6e-19
C43747 a_2982_43646# a_8037_42858# 5.75e-20
C43748 a_3626_43646# a_7871_42858# 3.84e-20
C43749 a_526_44458# a_1443_43940# 0.001014f
C43750 a_626_44172# a_n2293_42834# 2.37e-20
C43751 a_13017_45260# a_14976_45348# 5.79e-21
C43752 a_4185_45028# a_4905_42826# 0.039846f
C43753 a_n443_42852# a_1414_42308# 0.193113f
C43754 a_6171_45002# a_18315_45260# 5.25e-20
C43755 a_n2293_45010# a_n2433_44484# 0.016908f
C43756 a_n2109_45247# a_n2661_44458# 0.001495f
C43757 a_n2017_45002# a_n4318_40392# 2.16e-20
C43758 w_11334_34010# a_5742_30871# 1.73e-19
C43759 a_8049_45260# a_15493_43940# 4.49e-20
C43760 a_1823_45246# a_3626_43646# 0.033967f
C43761 a_n2661_45010# a_n2267_44484# 0.260289f
C43762 a_13507_46334# a_22400_42852# 0.235269f
C43763 a_15227_44166# a_17486_43762# 1.43e-19
C43764 a_18909_45814# a_18989_43940# 4.16e-19
C43765 a_18691_45572# a_18374_44850# 2.44e-20
C43766 a_n237_47217# a_5263_45724# 1.16e-19
C43767 a_n443_46116# a_n23_45546# 0.118272f
C43768 a_3090_45724# a_765_45546# 0.001007f
C43769 a_4883_46098# a_12839_46116# 1.63e-19
C43770 a_20916_46384# a_22223_46124# 5.13e-19
C43771 a_21588_30879# a_6945_45028# 1.26e-19
C43772 a_768_44030# a_n1925_42282# 0.145535f
C43773 a_2905_45572# a_1990_45899# 1.24e-19
C43774 a_584_46384# a_509_45572# 3.56e-19
C43775 a_3877_44458# a_4704_46090# 3.8e-19
C43776 a_4646_46812# a_4419_46090# 1.97e-19
C43777 a_13507_46334# a_14949_46494# 2.9e-19
C43778 a_18597_46090# a_16375_45002# 0.105669f
C43779 a_11599_46634# a_20850_46155# 7e-21
C43780 a_n743_46660# a_17583_46090# 4.13e-19
C43781 a_16327_47482# a_20850_46482# 2.1e-19
C43782 a_15368_46634# a_15312_46660# 1.11e-19
C43783 a_n881_46662# a_5210_46155# 1.33e-19
C43784 a_6755_46942# a_12741_44636# 0.131965f
C43785 a_4955_46873# a_3699_46348# 1.24e-20
C43786 a_11967_42832# RST_Z 4.49e-20
C43787 a_3422_30871# C2_P_btm 9.13e-20
C43788 a_19164_43230# a_19987_42826# 3.85e-19
C43789 a_n97_42460# a_7174_31319# 6.58e-20
C43790 a_3626_43646# a_11897_42308# 3.42e-19
C43791 a_3080_42308# a_4958_30871# 0.01856f
C43792 a_7765_42852# a_7309_42852# 0.00456f
C43793 a_19615_44636# VDD 0.203841f
C43794 a_3483_46348# a_8483_43230# 1.15e-21
C43795 a_3090_45724# a_4921_42308# 0.001886f
C43796 a_16112_44458# a_17970_44736# 6.26e-20
C43797 a_14539_43914# a_17767_44458# 3.19e-19
C43798 a_4223_44672# a_5289_44734# 0.009506f
C43799 a_n357_42282# a_16409_43396# 1.19e-20
C43800 a_17715_44484# a_17595_43084# 7.53e-21
C43801 a_n2312_38680# a_n3420_39616# 1.39e-19
C43802 a_626_44172# a_1115_44172# 0.00354f
C43803 a_1307_43914# a_2127_44172# 0.127867f
C43804 a_375_42282# a_1414_42308# 6.78e-21
C43805 a_7499_43078# a_6765_43638# 3.15e-19
C43806 a_n443_42852# a_12281_43396# 0.030395f
C43807 a_526_44458# a_7227_42852# 0.062474f
C43808 a_n1059_45260# a_18079_43940# 5.09e-19
C43809 a_11691_44458# a_14112_44734# 0.005155f
C43810 a_n2442_46660# a_n2302_39866# 0.161638f
C43811 a_10903_43370# a_14840_46494# 8.02e-21
C43812 a_6419_46155# a_6945_45028# 1.24e-19
C43813 a_1138_42852# a_526_44458# 0.039045f
C43814 a_12741_44636# a_8049_45260# 0.037594f
C43815 a_13759_46122# a_13925_46122# 0.576786f
C43816 a_19321_45002# a_16147_45260# 1.91e-21
C43817 a_19123_46287# a_16375_45002# 1.65e-19
C43818 a_18285_46348# a_19240_46482# 2.07e-21
C43819 a_13661_43548# a_18341_45572# 0.037017f
C43820 a_5807_45002# a_18909_45814# 0.001758f
C43821 a_13747_46662# a_18479_45785# 0.020713f
C43822 a_n2312_39304# a_n2661_45010# 1.13e-20
C43823 a_18597_46090# a_413_45260# 1.48e-19
C43824 a_17339_46660# a_18051_46116# 0.040259f
C43825 a_4915_47217# a_14537_43396# 5.76e-19
C43826 a_n743_46660# a_8696_44636# 0.032893f
C43827 a_472_46348# a_835_46155# 0.005265f
C43828 a_2063_45854# a_2304_45348# 0.001671f
C43829 a_n2109_47186# a_5837_45028# 0.001685f
C43830 a_1576_42282# a_1606_42308# 0.176925f
C43831 a_961_42354# a_1149_42558# 7.47e-21
C43832 a_n3674_37592# a_n327_42308# 0.002227f
C43833 a_1184_42692# a_1221_42558# 3.52e-19
C43834 a_1067_42314# a_1755_42282# 8.86e-19
C43835 a_3080_42308# VCM 0.148824f
C43836 a_14537_43396# a_15681_43442# 2.41e-19
C43837 a_7411_46660# VDD 0.41059f
C43838 a_17730_32519# a_19237_31679# 0.058836f
C43839 en_comp a_13678_32519# 1.37e-19
C43840 a_n755_45592# a_n3674_37592# 0.063692f
C43841 a_n863_45724# a_961_42354# 0.038222f
C43842 a_n357_42282# a_564_42282# 0.026735f
C43843 a_2711_45572# a_18707_42852# 2.52e-19
C43844 a_n2293_43922# a_10729_43914# 1.27e-20
C43845 a_n2661_42834# a_10807_43548# 0.003836f
C43846 a_n2661_43922# a_10949_43914# 9.62e-19
C43847 a_5883_43914# a_9420_43940# 0.001123f
C43848 a_n2293_45546# a_n452_45724# 2.19e-20
C43849 a_n1079_45724# a_n863_45724# 0.091159f
C43850 a_n2438_43548# a_n1917_44484# 2.8e-19
C43851 a_14976_45028# a_1307_43914# 4.47e-20
C43852 a_n2497_47436# a_175_44278# 0.05097f
C43853 a_11415_45002# a_19963_31679# 0.033926f
C43854 a_21076_30879# a_2437_43646# 3e-20
C43855 a_5066_45546# a_9049_44484# 3.93e-19
C43856 a_n2661_45546# a_310_45028# 0.035423f
C43857 a_n2472_45546# a_n1099_45572# 9.27e-20
C43858 a_12549_44172# a_18287_44626# 0.006594f
C43859 a_19123_46287# a_413_45260# 4.85e-21
C43860 a_10227_46804# a_15433_44458# 0.001023f
C43861 a_5807_45002# a_12607_44458# 5.72e-21
C43862 a_12861_44030# a_17061_44734# 1.88e-19
C43863 a_15227_44166# a_14180_45002# 2.28e-19
C43864 a_n2293_46634# a_2779_44458# 0.004655f
C43865 a_2324_44458# a_11778_45572# 8.28e-19
C43866 a_n971_45724# a_n785_47204# 0.385455f
C43867 a_n746_45260# a_n23_47502# 0.148631f
C43868 a_n1741_47186# a_2124_47436# 0.009997f
C43869 a_n2109_47186# a_2063_45854# 0.045645f
C43870 a_5742_30871# a_n4064_37984# 0.004679f
C43871 COMP_P a_22545_38993# 4.2e-21
C43872 a_3905_42865# a_6197_43396# 1.51e-20
C43873 a_3065_45002# a_3581_42558# 0.003532f
C43874 a_11967_42832# a_16243_43396# 0.269605f
C43875 a_17517_44484# a_19268_43646# 3.12e-21
C43876 a_10555_44260# a_10651_43940# 0.001863f
C43877 a_15493_43940# a_15037_43940# 0.004121f
C43878 a_n2017_45002# a_8337_42558# 4.83e-19
C43879 a_n2661_42282# a_1209_43370# 2.03e-21
C43880 a_10729_43914# a_n97_42460# 2.13e-20
C43881 a_10057_43914# a_10796_42968# 1.53e-19
C43882 a_3537_45260# a_5379_42460# 6.86e-20
C43883 a_20205_31679# a_22459_39145# 2.38e-20
C43884 a_20692_30879# a_22521_40055# 1.07e-20
C43885 en_comp a_6123_31319# 0.028738f
C43886 a_19862_44208# a_19741_43940# 0.038152f
C43887 a_7920_46348# a_6298_44484# 1.48e-19
C43888 a_6945_45028# a_21359_45002# 1.23e-21
C43889 a_17715_44484# a_17896_45144# 3.62e-20
C43890 a_2277_45546# a_413_45260# 1.14e-20
C43891 a_n443_42852# a_1667_45002# 3.6e-19
C43892 a_5257_43370# a_5663_43940# 0.014098f
C43893 a_15037_45618# a_15765_45572# 3.63e-20
C43894 a_19466_46812# a_20362_44736# 3.02e-19
C43895 a_19692_46634# a_20159_44458# 0.001725f
C43896 a_n971_45724# a_9803_43646# 5.86e-21
C43897 a_15227_44166# a_20679_44626# 1.44e-21
C43898 a_4791_45118# a_7112_43396# 1.4e-19
C43899 a_13747_46662# a_14021_43940# 1.12e-19
C43900 a_13661_43548# a_14485_44260# 4.85e-19
C43901 a_768_44030# a_3737_43940# 0.038628f
C43902 a_8049_45260# a_n2293_42834# 0.224469f
C43903 a_8953_45546# a_4223_44672# 5.72e-21
C43904 a_n4064_38528# VDD 1.69517f
C43905 a_5700_37509# a_6886_37412# 0.13762f
C43906 a_5088_37509# VDAC_N 0.420254f
C43907 a_n4064_39072# VREF_GND 0.048253f
C43908 a_3726_37500# VDAC_P 0.059581f
C43909 a_4338_37500# a_8912_37509# 0.331796f
C43910 a_6491_46660# a_7411_46660# 2.68e-21
C43911 a_n1435_47204# a_5907_46634# 3.08e-20
C43912 a_n1741_47186# a_11813_46116# 0.004098f
C43913 a_n237_47217# a_8270_45546# 0.552109f
C43914 a_n971_45724# a_8601_46660# 5.7e-19
C43915 a_n1151_42308# a_10249_46116# 0.060327f
C43916 a_6151_47436# a_7577_46660# 0.578207f
C43917 a_4915_47217# a_8667_46634# 4.1e-20
C43918 a_6545_47178# a_7715_46873# 0.003195f
C43919 a_2747_46873# a_n1925_46634# 0.007371f
C43920 a_3422_30871# a_20256_42852# 1.38e-20
C43921 a_5891_43370# a_9885_42558# 0.001022f
C43922 a_20512_43084# a_20256_43172# 0.047194f
C43923 a_17538_32519# a_17364_32525# 9.64512f
C43924 a_8685_43396# a_14579_43548# 0.03481f
C43925 a_n2293_43922# a_5932_42308# 0.178011f
C43926 a_3626_43646# a_17324_43396# 4.75e-21
C43927 a_11341_43940# a_15567_42826# 3.04e-20
C43928 a_20841_45814# VDD 0.209907f
C43929 a_20974_43370# a_20749_43396# 0.0837f
C43930 a_1823_45246# a_3052_44056# 2.45e-20
C43931 a_6171_45002# a_13017_45260# 0.045098f
C43932 a_2382_45260# a_1307_43914# 0.53878f
C43933 a_7705_45326# a_8191_45002# 5.55e-19
C43934 a_13904_45546# a_13720_44458# 2.89e-21
C43935 a_13249_42308# a_13076_44458# 1.5e-19
C43936 a_n443_42852# a_14112_44734# 2.65e-20
C43937 a_20202_43084# a_19319_43548# 2.44e-19
C43938 a_1667_45002# a_375_42282# 2.16e-20
C43939 a_413_45260# a_626_44172# 0.032584f
C43940 a_18341_45572# a_18587_45118# 8.86e-19
C43941 a_18479_45785# a_18911_45144# 0.00112f
C43942 a_13507_46334# a_22223_42860# 0.049534f
C43943 a_n2442_46660# a_n3674_39304# 0.024039f
C43944 a_768_44030# a_8387_43230# 1.54e-20
C43945 a_3483_46348# a_15037_44260# 6.29e-19
C43946 a_n2438_43548# a_n1853_43023# 0.001525f
C43947 a_3090_45724# a_6452_43396# 0.001752f
C43948 a_13259_45724# a_3422_30871# 0.587088f
C43949 a_2324_44458# a_13483_43940# 3.39e-21
C43950 a_5066_45546# a_3905_42865# 0.001745f
C43951 a_768_44030# a_2698_46116# 0.001262f
C43952 a_3699_46634# a_765_45546# 0.002795f
C43953 a_6755_46942# a_13607_46688# 0.129798f
C43954 a_11309_47204# a_3483_46348# 1.47e-20
C43955 a_4883_46098# a_14840_46494# 0.004918f
C43956 a_18479_47436# a_19335_46494# 1.52e-20
C43957 a_16327_47482# a_10809_44734# 0.036039f
C43958 a_16763_47508# a_6945_45028# 0.01658f
C43959 a_13507_46334# a_15682_46116# 0.022078f
C43960 a_n881_46662# a_5497_46414# 0.001017f
C43961 a_n1613_43370# a_6165_46155# 3.04e-19
C43962 a_4791_45118# a_5527_46155# 2.63e-19
C43963 a_18597_46090# a_18985_46122# 0.027318f
C43964 a_19386_47436# a_18819_46122# 1.81e-21
C43965 a_12465_44636# a_14275_46494# 0.00587f
C43966 a_11453_44696# a_13351_46090# 8.02e-21
C43967 a_14021_43940# a_4958_30871# 2.74e-20
C43968 a_7871_42858# a_8037_42858# 0.772842f
C43969 a_14579_43548# a_15953_42852# 1.82e-19
C43970 a_n97_42460# a_5932_42308# 2.52e-19
C43971 a_1987_43646# a_1606_42308# 3.6e-36
C43972 a_13678_32519# a_22165_42308# 0.018986f
C43973 a_5649_42852# a_21671_42860# 0.003655f
C43974 a_n2012_44484# VDD 0.077632f
C43975 a_1307_43914# a_15433_44458# 2.11e-20
C43976 a_n2661_43370# a_n356_44636# 0.002184f
C43977 a_n2840_44458# a_n4318_40392# 0.161548f
C43978 a_n2472_45002# a_n2472_43914# 0.001034f
C43979 a_n2661_45010# a_n2065_43946# 0.001138f
C43980 a_13661_43548# a_15803_42450# 3.06e-22
C43981 a_n863_45724# a_2982_43646# 2.39e-20
C43982 a_n2293_45010# a_n2840_43914# 4.9e-20
C43983 a_n2442_46660# a_5742_30871# 8.02e-21
C43984 a_3090_45724# a_13291_42460# 0.002769f
C43985 a_n357_42282# a_n1557_42282# 0.384406f
C43986 a_n755_45592# a_766_43646# 3.04e-19
C43987 a_10907_45822# a_11173_44260# 7.74e-20
C43988 a_2437_43646# a_1414_42308# 0.023872f
C43989 a_8696_44636# a_11750_44172# 3.79e-20
C43990 a_16333_45814# a_15682_43940# 2.17e-19
C43991 a_n2497_47436# a_n143_45144# 1.83e-21
C43992 a_n971_45724# a_n913_45002# 0.101346f
C43993 a_n746_45260# a_n1059_45260# 0.138039f
C43994 a_12465_44636# a_15765_45572# 2.53e-21
C43995 a_16327_47482# a_16211_45572# 1.79e-19
C43996 a_n2293_46634# a_2211_45572# 3.32e-19
C43997 a_1823_45246# a_167_45260# 0.155648f
C43998 a_n743_46660# a_7227_45028# 0.001306f
C43999 a_768_44030# a_13527_45546# 1.49e-20
C44000 a_12549_44172# a_13904_45546# 5.84e-19
C44001 a_12891_46348# a_13249_42308# 0.166217f
C44002 a_19123_46287# a_18985_46122# 0.215692f
C44003 a_6755_46942# a_16375_45002# 8.39e-21
C44004 a_18285_46348# a_19553_46090# 7.38e-22
C44005 SMPL_ON_P en_comp 0.034192f
C44006 a_3381_47502# a_2437_43646# 0.004114f
C44007 a_12861_44030# a_19431_45546# 1.85e-20
C44008 a_5807_45002# a_8746_45002# 7.32e-20
C44009 a_13661_43548# a_10193_42453# 0.211481f
C44010 a_11813_46116# a_10586_45546# 7.37e-19
C44011 a_16434_46987# a_10809_44734# 9.15e-19
C44012 a_11599_46634# a_18479_45785# 0.028968f
C44013 a_5829_43940# VDD 0.156797f
C44014 a_5534_30871# a_11551_42558# 5.08e-19
C44015 a_12089_42308# a_13333_42558# 2.22e-19
C44016 a_17364_32525# a_22465_38105# 2.07e-19
C44017 a_20202_43084# a_21335_42336# 0.227943f
C44018 a_5111_44636# a_6293_42852# 0.072755f
C44019 a_5343_44458# a_7911_44260# 0.005844f
C44020 a_5147_45002# a_6197_43396# 9.61e-19
C44021 a_8953_45546# a_5742_30871# 1.11e-19
C44022 a_4185_45028# a_15803_42450# 2.86e-19
C44023 a_13661_43548# VDD 3.93017f
C44024 a_5883_43914# a_5841_44260# 2.9e-21
C44025 a_4223_44672# a_9028_43914# 5.03e-20
C44026 a_3537_45260# a_7287_43370# 0.400907f
C44027 a_413_45260# a_2813_43396# 6.05e-21
C44028 a_5807_45002# RST_Z 1.85e-19
C44029 a_10193_42453# a_10835_43094# 0.041273f
C44030 a_12549_44172# CLK 3.33e-19
C44031 a_n357_42282# a_8483_43230# 7.88e-19
C44032 a_n755_45592# a_8292_43218# 0.010247f
C44033 a_526_44458# a_1576_42282# 2.98e-20
C44034 a_13259_45724# a_18504_43218# 9.31e-20
C44035 a_18911_45144# a_14021_43940# 1.04e-20
C44036 a_n1925_42282# a_1067_42314# 5.5e-20
C44037 a_9290_44172# a_9885_42558# 0.021204f
C44038 a_20193_45348# a_15493_43940# 0.10893f
C44039 a_n443_42852# a_873_42968# 5.2e-19
C44040 a_7499_43078# a_10341_42308# 0.42152f
C44041 a_12861_44030# a_13076_44458# 0.01178f
C44042 a_15009_46634# a_2437_43646# 7.72e-21
C44043 a_5807_45002# a_14403_45348# 0.002634f
C44044 a_n2497_47436# a_n2293_43922# 9.38e-20
C44045 a_12549_44172# a_17023_45118# 5.36e-21
C44046 a_8270_45546# a_n2017_45002# 4.47e-21
C44047 a_19692_46634# a_20623_45572# 5.14e-19
C44048 a_19466_46812# a_21363_45546# 9.08e-21
C44049 a_14275_46494# a_2711_45572# 1.13e-20
C44050 a_6755_46942# a_413_45260# 6.02e-20
C44051 a_13059_46348# a_16147_45260# 1.3e-19
C44052 a_12816_46660# a_3357_43084# 5.53e-21
C44053 a_8049_45260# a_16375_45002# 0.026933f
C44054 a_6419_46155# a_6812_45938# 7.41e-19
C44055 a_5257_43370# a_3232_43370# 0.022872f
C44056 a_3483_46348# a_10490_45724# 0.207668f
C44057 a_4185_45028# a_10193_42453# 3.16135f
C44058 a_n1630_35242# a_n3565_38502# 1.85e-19
C44059 a_5742_30871# a_13258_32519# 0.004591f
C44060 a_n4318_38216# a_n3565_38216# 3.9e-19
C44061 a_5342_30871# C0_P_btm 8.41e-20
C44062 a_n3674_37592# a_n3420_38528# 0.020112f
C44063 a_5534_30871# C0_dummy_N_btm 2.22e-20
C44064 a_15764_42576# a_4958_30871# 0.413236f
C44065 a_15486_42560# a_17303_42282# 3.91e-21
C44066 a_15890_42674# a_15761_42308# 4.2e-19
C44067 a_15959_42545# a_16197_42308# 0.001705f
C44068 a_15803_42450# a_16269_42308# 3.82e-19
C44069 a_n3674_38680# a_n3420_37984# 2.36e-20
C44070 a_1606_42308# a_1736_39043# 7.77e-20
C44071 a_10835_43094# VDD 0.43308f
C44072 a_10533_42308# a_7174_31319# 4.88e-21
C44073 a_14113_42308# a_18057_42282# 2.13e-20
C44074 a_n784_42308# a_n4064_38528# 0.004411f
C44075 a_n3674_38216# a_n4209_38216# 0.059407f
C44076 a_10405_44172# a_11341_43940# 0.001372f
C44077 a_5495_43940# a_5829_43940# 0.001349f
C44078 a_5663_43940# a_5745_43940# 0.096132f
C44079 a_17970_44736# a_17499_43370# 9.31e-19
C44080 a_11823_42460# a_13657_42308# 4.58e-19
C44081 a_n1059_45260# a_17749_42852# 8.24e-19
C44082 a_4185_45028# VDD 1.65665f
C44083 a_19237_31679# a_17538_32519# 0.060188f
C44084 a_15682_43940# a_15493_43396# 9.79e-19
C44085 a_17973_43940# a_18451_43940# 0.0015f
C44086 a_19721_31679# a_17364_32525# 0.053872f
C44087 a_n2956_38216# a_n4209_38502# 0.023653f
C44088 a_20447_31679# a_14097_32519# 0.05131f
C44089 a_9313_44734# a_9803_43646# 2.3e-19
C44090 a_18079_43940# a_18326_43940# 0.152347f
C44091 a_5204_45822# a_n2661_43370# 4.54e-21
C44092 a_8199_44636# a_8488_45348# 0.001482f
C44093 a_5807_45002# a_5663_43940# 2.36e-20
C44094 a_11962_45724# a_13163_45724# 0.113317f
C44095 a_8568_45546# a_8697_45822# 0.062574f
C44096 a_8953_45546# a_n2293_42834# 4.91e-20
C44097 a_n2438_43548# a_n1899_43946# 8.61e-19
C44098 a_12741_44636# a_20193_45348# 0.012699f
C44099 a_n2497_47436# a_n97_42460# 0.026966f
C44100 a_12427_45724# a_12791_45546# 0.124682f
C44101 a_2711_45572# a_15765_45572# 0.005291f
C44102 a_5066_45546# a_5147_45002# 5.3e-19
C44103 a_5431_46482# a_5111_44636# 6.74e-20
C44104 a_14035_46660# a_13720_44458# 7.64e-21
C44105 a_8049_45260# a_413_45260# 0.140877f
C44106 a_11453_44696# a_17973_43940# 1.73e-21
C44107 a_n1151_42308# a_n2472_46634# 1.07e-20
C44108 a_3381_47502# a_n2661_46634# 2.12e-20
C44109 a_2905_45572# a_n2293_46634# 8.29e-19
C44110 a_6851_47204# a_5807_45002# 7.21e-20
C44111 a_12861_44030# a_12891_46348# 0.053595f
C44112 a_13717_47436# a_12549_44172# 0.002227f
C44113 a_n1435_47204# a_768_44030# 6.95e-20
C44114 a_7174_31319# C2_P_btm 1.86e-20
C44115 a_n2497_47436# a_n2661_46098# 0.026032f
C44116 a_22731_47423# SMPL_ON_N 0.194951f
C44117 a_1431_47204# a_n2438_43548# 5.68e-21
C44118 a_2063_45854# a_n1925_46634# 0.064288f
C44119 a_12465_44636# a_22959_47212# 3.19e-20
C44120 a_22223_47212# a_11453_44696# 0.057984f
C44121 a_n746_45260# a_948_46660# 0.001665f
C44122 a_n971_45724# a_2107_46812# 0.06261f
C44123 a_327_47204# a_33_46660# 0.001418f
C44124 a_n237_47217# a_1123_46634# 0.003027f
C44125 a_n3565_39590# a_n1386_35608# 1.44e-19
C44126 a_16327_47482# a_n881_46662# 0.195459f
C44127 a_20512_43084# a_21195_42852# 2.47e-19
C44128 a_9313_44734# a_19518_43218# 1.42e-19
C44129 a_11341_43940# a_20556_43646# 0.004978f
C44130 a_11415_45002# a_10729_43914# 1.25e-20
C44131 a_n2661_45010# a_n2810_45028# 0.009249f
C44132 a_n2293_45010# a_n913_45002# 0.015951f
C44133 a_n2109_45247# a_n1059_45260# 1.05e-19
C44134 SMPL_ON_N a_14209_32519# 0.02932f
C44135 a_3090_45724# a_11173_43940# 1.22e-19
C44136 a_19479_31679# a_413_45260# 0.055869f
C44137 a_6945_45028# a_19279_43940# 1.94e-21
C44138 a_n2293_46098# a_6101_44260# 1.56e-19
C44139 a_n2840_45002# a_n2956_37592# 0.035532f
C44140 a_2437_43646# a_1667_45002# 0.005688f
C44141 a_n443_42852# a_n699_43396# 0.333516f
C44142 a_5257_43370# a_4905_42826# 0.254437f
C44143 a_10193_42453# a_18587_45118# 7.6e-21
C44144 a_13059_46348# a_13565_44260# 8.69e-19
C44145 a_n2293_46634# a_10765_43646# 0.001573f
C44146 a_12549_44172# a_19268_43646# 3.27e-20
C44147 a_13661_43548# a_16137_43396# 2.21e-19
C44148 VDD VREF_GND 0.482759f
C44149 a_4646_46812# a_7411_46660# 0.266058f
C44150 a_4651_46660# a_5257_43370# 2.06e-19
C44151 a_19594_46812# a_15227_44166# 0.073663f
C44152 a_19321_45002# a_19333_46634# 0.001085f
C44153 a_5807_45002# a_10425_46660# 2.9e-19
C44154 a_12549_44172# a_14035_46660# 0.026143f
C44155 a_768_44030# a_13885_46660# 0.029614f
C44156 a_5385_46902# a_5894_47026# 2.6e-19
C44157 a_4817_46660# a_5263_46660# 2.28e-19
C44158 a_2063_45854# a_10355_46116# 9.15e-21
C44159 a_2583_47243# a_765_45546# 2e-19
C44160 a_n1435_47204# a_1176_45822# 2.97e-20
C44161 a_19452_47524# a_19466_46812# 4e-19
C44162 a_13747_46662# a_19692_46634# 0.001071f
C44163 a_4915_47217# a_5204_45822# 4.09e-20
C44164 a_4791_45118# a_6165_46155# 0.291653f
C44165 a_n1151_42308# a_5937_45572# 0.11638f
C44166 a_n743_46660# a_11813_46116# 0.003585f
C44167 a_3877_44458# a_7715_46873# 2.82e-20
C44168 a_13507_46334# a_20719_46660# 7.51e-19
C44169 a_10227_46804# a_21297_46660# 6.03e-19
C44170 a_11453_44696# a_20731_47026# 0.026307f
C44171 a_14209_32519# a_22959_43396# 0.015679f
C44172 a_22591_43396# a_17364_32525# 7.75e-19
C44173 a_19721_31679# a_21589_35634# 1.38e-20
C44174 a_10341_43396# a_15567_42826# 0.004039f
C44175 a_21381_43940# a_20256_43172# 6.27e-20
C44176 a_3539_42460# a_4649_42852# 0.006668f
C44177 a_n97_42460# a_17141_43172# 3.1e-19
C44178 a_18587_45118# VDD 0.085535f
C44179 a_19237_31679# a_22465_38105# 2.6e-19
C44180 a_10729_43914# a_10533_42308# 2.31e-20
C44181 a_18341_45572# a_11967_42832# 6.68e-21
C44182 a_18479_45785# a_19615_44636# 0.006445f
C44183 a_3090_45724# a_13460_43230# 0.004635f
C44184 a_768_44030# a_1606_42308# 0.00182f
C44185 a_1307_43914# a_5343_44458# 0.02568f
C44186 a_375_42282# a_n699_43396# 0.127058f
C44187 a_2711_45572# a_19328_44172# 0.010017f
C44188 a_n2312_40392# a_5934_30871# 8.24e-21
C44189 a_4883_46098# a_9223_42460# 2.45e-19
C44190 a_11415_45002# a_21487_43396# 1.71e-21
C44191 a_526_44458# a_1987_43646# 3.41e-20
C44192 a_1423_45028# a_742_44458# 0.019572f
C44193 a_n913_45002# a_9313_44734# 0.055701f
C44194 a_9482_43914# a_10440_44484# 0.001083f
C44195 a_n2956_39768# a_n2472_42282# 3.63e-20
C44196 a_10903_43370# a_13667_43396# 7.81e-20
C44197 a_3483_46348# a_16547_43609# 5.46e-20
C44198 a_4185_45028# a_16137_43396# 1.37e-19
C44199 w_1575_34946# VDAC_Pi 5.84e-19
C44200 a_4883_46098# a_6511_45714# 6.24e-20
C44201 a_10768_47026# a_10903_43370# 7.21e-21
C44202 a_5807_45002# a_21167_46155# 1.15e-20
C44203 a_6151_47436# a_6905_45572# 0.003156f
C44204 a_12861_44030# a_11322_45546# 7.65e-19
C44205 a_18285_46348# a_12741_44636# 8.73e-21
C44206 a_20107_46660# a_11415_45002# 2.81e-22
C44207 a_20411_46873# a_20202_43084# 1.99e-21
C44208 a_20623_46660# a_20719_46660# 0.013793f
C44209 a_20841_46902# a_20885_46660# 3.69e-19
C44210 a_20273_46660# a_22365_46825# 7.72e-20
C44211 a_n881_46662# a_n356_45724# 0.002904f
C44212 a_11813_46116# a_11189_46129# 0.009001f
C44213 a_9863_46634# a_6945_45028# 1.05e-19
C44214 a_5649_42852# a_9223_42460# 6.66e-20
C44215 a_16977_43638# a_17124_42282# 4.32e-20
C44216 a_10341_43396# a_20712_42282# 2.59e-20
C44217 a_4361_42308# a_9377_42558# 8.36e-20
C44218 a_1847_42826# a_2713_42308# 0.015903f
C44219 a_18817_42826# a_18707_42852# 0.097745f
C44220 a_3080_42308# a_n4064_38528# 0.001913f
C44221 a_10835_43094# a_n784_42308# 1.43e-21
C44222 a_5111_42852# a_1755_42282# 2.49e-20
C44223 a_743_42282# a_11323_42473# 0.008466f
C44224 a_n755_45592# a_3681_42891# 1.63e-20
C44225 a_n357_42282# a_3935_42891# 0.007216f
C44226 a_4185_45028# a_n784_42308# 7.16e-20
C44227 a_8375_44464# a_n2661_42834# 3.77e-20
C44228 a_16112_44458# a_16335_44484# 0.011458f
C44229 a_14311_47204# RST_Z 0.184572f
C44230 a_19721_31679# a_19237_31679# 0.071506f
C44231 a_13259_45724# a_16414_43172# 3.58e-20
C44232 a_526_44458# a_4649_42852# 0.028795f
C44233 a_2324_44458# a_15597_42852# 3.41e-19
C44234 a_8975_43940# a_11967_42832# 1.12e-20
C44235 a_7640_43914# a_n2661_43922# 0.019048f
C44236 a_n1435_47204# DATA[0] 0.053257f
C44237 a_18248_44752# a_17517_44484# 0.561898f
C44238 a_17970_44736# a_18204_44850# 0.006453f
C44239 a_n913_45002# a_20974_43370# 2.82e-20
C44240 a_n2661_45010# a_n2129_43609# 1.46e-20
C44241 a_3232_43370# a_5745_43940# 1.59e-19
C44242 a_1138_42852# a_1221_42558# 6.61e-20
C44243 a_14955_47212# VDD 0.301751f
C44244 a_18985_46122# a_8049_45260# 0.006692f
C44245 a_10903_43370# a_11601_46155# 2.78e-19
C44246 a_n2293_46098# a_n23_45546# 0.00525f
C44247 a_472_46348# a_n357_42282# 0.001836f
C44248 a_376_46348# a_n755_45592# 1.77e-21
C44249 a_n971_45724# a_n2661_44458# 0.051008f
C44250 a_5807_45002# a_3232_43370# 0.091049f
C44251 a_n2438_43548# en_comp 0.915368f
C44252 a_n2293_46634# a_n37_45144# 0.006632f
C44253 a_13759_46122# a_12638_46436# 1.15e-20
C44254 a_768_44030# a_10775_45002# 1.05e-21
C44255 a_n2497_47436# a_742_44458# 0.153038f
C44256 a_1823_45246# a_n863_45724# 0.207189f
C44257 a_1176_45822# a_380_45546# 2.97e-19
C44258 a_2804_46116# a_n2661_45546# 1.07e-20
C44259 a_n881_46662# a_14537_43396# 1.17e-21
C44260 a_167_45260# a_n2293_45546# 0.681309f
C44261 a_8515_42308# a_8685_42308# 0.108744f
C44262 a_5934_30871# a_8791_42308# 0.223675f
C44263 a_4190_30871# C0_dummy_N_btm 1.45e-20
C44264 a_22400_42852# a_21613_42308# 0.024416f
C44265 a_17364_32525# a_18194_35068# 9.45e-20
C44266 a_n913_45002# a_18599_43230# 1.4e-20
C44267 a_n2017_45002# a_19164_43230# 0.048221f
C44268 a_3357_43084# a_4156_43218# 2.37e-19
C44269 a_19615_44636# a_14021_43940# 4.32e-21
C44270 a_5883_43914# a_6547_43396# 2.84e-19
C44271 a_3600_43914# a_3499_42826# 0.125876f
C44272 a_2998_44172# a_3820_44260# 1.27e-20
C44273 a_21076_30879# a_22609_38406# 5.77e-21
C44274 a_n356_44636# a_1568_43370# 7.66e-20
C44275 a_14543_46987# VDD 8.63e-19
C44276 a_2779_44458# a_2813_43396# 3.22e-21
C44277 a_13259_45724# a_7174_31319# 0.033027f
C44278 a_n2956_38680# a_n2860_38778# 0.001355f
C44279 a_n357_42282# a_15890_42674# 1.81e-20
C44280 en_comp a_18083_42858# 1.15e-20
C44281 a_10861_46660# CLK 9.26e-19
C44282 SMPL_ON_N a_17730_32519# 0.029186f
C44283 a_n2312_38680# a_n2661_43922# 1.97e-21
C44284 a_3483_46348# a_6171_45002# 0.153232f
C44285 a_3699_46348# a_3232_43370# 6.75e-20
C44286 a_4185_45028# a_5691_45260# 1.6e-19
C44287 a_15227_44166# a_18494_42460# 3.03e-20
C44288 a_2711_45572# a_6194_45824# 0.013872f
C44289 a_2107_46812# a_9313_44734# 0.023852f
C44290 a_13661_43548# a_13940_44484# 0.002141f
C44291 a_5068_46348# a_5147_45002# 5.26e-21
C44292 a_5164_46348# a_4558_45348# 0.002407f
C44293 a_18819_46122# a_3357_43084# 3.26e-20
C44294 a_2063_45854# a_10949_43914# 0.129837f
C44295 a_8953_45546# a_413_45260# 4.56e-21
C44296 a_19466_46812# a_19778_44110# 0.116901f
C44297 a_19335_46494# a_2437_43646# 5.23e-21
C44298 a_15890_42674# CAL_N 6.88e-19
C44299 a_5932_42308# C2_P_btm 0.011289f
C44300 a_9067_47204# a_n1435_47204# 0.001005f
C44301 a_11031_47542# a_11459_47204# 0.001175f
C44302 a_n2946_39072# a_n4064_38528# 3.78e-20
C44303 a_n4064_39072# a_n2946_38778# 3.78e-20
C44304 a_n3565_39304# a_n2216_38778# 1e-19
C44305 a_n4064_39616# a_n4064_37984# 0.048968f
C44306 a_4958_30871# a_n4064_37440# 0.031235f
C44307 a_n1605_47204# a_n2312_39304# 0.001342f
C44308 a_5934_30871# C9_P_btm 1.37e-19
C44309 a_6151_47436# a_15507_47210# 0.003878f
C44310 a_6123_31319# C7_P_btm 0.005631f
C44311 a_n784_42308# VREF_GND 0.068593f
C44312 a_n1741_47186# a_n89_47570# 3.69e-19
C44313 a_n39_42308# VDD 0.00143f
C44314 a_10405_44172# a_10341_43396# 6.35e-20
C44315 a_n913_45002# a_22397_42558# 1.07e-20
C44316 a_644_44056# a_743_42282# 5.65e-22
C44317 a_20692_30879# VCM 0.035438f
C44318 a_997_45618# VDD 0.12359f
C44319 en_comp a_22775_42308# 9.56e-20
C44320 a_9313_44734# a_20922_43172# 0.011702f
C44321 a_17730_32519# a_22959_43396# 0.001049f
C44322 a_12861_44030# a_16409_43396# 9.01e-20
C44323 a_4646_46812# a_5829_43940# 2.16e-19
C44324 a_11322_45546# a_11787_45002# 0.035999f
C44325 a_2711_45572# a_6517_45366# 3.03e-19
C44326 a_n881_46662# a_6547_43396# 1.22e-20
C44327 a_n1613_43370# a_7287_43370# 0.337957f
C44328 a_n2497_47436# a_n901_43156# 0.006149f
C44329 SMPL_ON_P a_n2157_42858# 6.32e-21
C44330 a_n2438_43548# a_n1699_43638# 4.93e-19
C44331 a_8034_45724# a_5343_44458# 2.52e-21
C44332 a_3503_45724# a_n2661_43370# 3.04e-20
C44333 a_3483_46348# a_14673_44172# 0.026455f
C44334 a_19256_45572# a_19418_45938# 0.006453f
C44335 a_18691_45572# a_18953_45572# 0.001705f
C44336 a_11415_45002# a_21398_44850# 9.56e-19
C44337 a_20202_43084# a_3422_30871# 0.527141f
C44338 a_14495_45572# a_6171_45002# 0.002012f
C44339 a_4880_45572# a_1307_43914# 2.88e-21
C44340 a_10490_45724# a_11963_45334# 2.16e-19
C44341 a_18194_35068# a_21589_35634# 4.88e-19
C44342 a_22469_40625# VDD 0.564837f
C44343 a_19120_35138# a_19864_35138# 0.081924f
C44344 a_22521_40599# RST_Z 2.23e-19
C44345 a_n4064_37440# VCM 0.020152f
C44346 EN_VIN_BSTR_P C7_P_btm 0.115875f
C44347 a_16327_47482# a_17609_46634# 0.001241f
C44348 a_16023_47582# a_16292_46812# 7.28e-19
C44349 a_n133_46660# a_491_47026# 9.73e-19
C44350 a_n2438_43548# a_n935_46688# 6.37e-19
C44351 a_11599_46634# a_19692_46634# 0.069066f
C44352 a_171_46873# a_288_46660# 0.159893f
C44353 a_n1925_46634# a_645_46660# 4.33e-19
C44354 a_n2661_46634# a_2959_46660# 0.006729f
C44355 a_n2293_46634# a_2443_46660# 1.47e-20
C44356 a_5807_45002# a_4651_46660# 8.13e-19
C44357 a_8128_46384# a_7715_46873# 0.006283f
C44358 a_n881_46662# a_8667_46634# 5.47e-20
C44359 a_10227_46804# a_3090_45724# 0.320681f
C44360 a_3381_47502# a_765_45546# 0.002383f
C44361 a_n2104_46634# a_n2661_46098# 1.32e-19
C44362 a_383_46660# a_948_46660# 7.99e-20
C44363 a_15781_43660# a_15940_43402# 0.002605f
C44364 a_10341_43396# a_20556_43646# 0.008164f
C44365 a_20974_43370# a_20922_43172# 0.002377f
C44366 a_21381_43940# a_21195_42852# 0.238789f
C44367 a_16547_43609# a_16664_43396# 0.161376f
C44368 a_16243_43396# a_16867_43762# 9.73e-19
C44369 a_13159_45002# VDD 0.321035f
C44370 a_n97_42460# a_15567_42826# 0.040819f
C44371 a_2998_44172# a_3823_42558# 8.6e-22
C44372 a_n2661_42282# a_n3674_38216# 0.051505f
C44373 a_16759_43396# a_15743_43084# 0.033478f
C44374 a_17324_43396# a_18525_43370# 0.003432f
C44375 a_11967_42832# a_15803_42450# 0.258862f
C44376 a_2982_43646# a_7765_42852# 3.2e-20
C44377 a_13017_45260# a_14403_45348# 0.001556f
C44378 a_14495_45572# a_14673_44172# 5.52e-19
C44379 a_4185_45028# a_3080_42308# 0.030391f
C44380 a_8696_44636# a_5891_43370# 0.084594f
C44381 a_n443_42852# a_1467_44172# 0.008372f
C44382 a_n2293_45546# a_n1453_44318# 1.08e-19
C44383 a_6171_45002# a_17719_45144# 8.44e-20
C44384 a_n2472_45002# a_n2433_44484# 7.88e-19
C44385 a_n2293_45010# a_n2661_44458# 0.031066f
C44386 a_18597_46090# a_20753_42852# 3.09e-19
C44387 a_n971_45724# a_8325_42308# 4.93e-20
C44388 a_2903_45348# a_2809_45028# 1.26e-19
C44389 a_1823_45246# a_3540_43646# 8.6e-19
C44390 a_10193_42453# a_11967_42832# 0.752992f
C44391 a_n2661_45010# a_n2129_44697# 0.18531f
C44392 a_2437_43646# a_n699_43396# 0.037149f
C44393 a_15227_44166# a_15940_43402# 6.38e-19
C44394 a_18341_45572# a_18989_43940# 7.86e-20
C44395 a_19431_45546# a_18287_44626# 6.77e-21
C44396 a_3503_45724# a_2998_44172# 3.02e-21
C44397 a_4791_45118# a_5379_42460# 0.197725f
C44398 a_16327_47482# a_19443_46116# 0.012553f
C44399 a_n1741_47186# a_6598_45938# 1.67e-22
C44400 a_n237_47217# a_4099_45572# 1.6e-19
C44401 a_n443_46116# a_n356_45724# 0.113738f
C44402 a_n1151_42308# a_n443_42852# 0.001061f
C44403 a_2905_45572# a_2277_45546# 5.92e-19
C44404 a_3090_45724# a_17339_46660# 0.019979f
C44405 a_15009_46634# a_765_45546# 6.36e-21
C44406 a_14976_45028# a_15312_46660# 0.01024f
C44407 a_10227_46804# a_15002_46116# 4.37e-19
C44408 a_20916_46384# a_6945_45028# 0.036695f
C44409 a_20843_47204# a_10809_44734# 9.21e-19
C44410 a_768_44030# a_526_44458# 0.341438f
C44411 a_3877_44458# a_4419_46090# 6.31e-19
C44412 a_4646_46812# a_4185_45028# 1.6e-20
C44413 a_15227_44166# a_16388_46812# 0.02839f
C44414 a_13507_46334# a_14537_46482# 7.17e-19
C44415 a_18597_46090# a_18243_46436# 6.59e-20
C44416 a_16292_46812# a_16751_46987# 6.64e-19
C44417 a_n881_46662# a_6640_46482# 6.85e-19
C44418 a_4955_46873# a_3483_46348# 1.84e-20
C44419 a_n2438_43548# a_2324_44458# 0.00362f
C44420 a_n743_46660# a_15682_46116# 0.051046f
C44421 a_8685_43396# a_9223_42460# 2.83e-20
C44422 a_3422_30871# C3_P_btm 1.1e-19
C44423 a_19339_43156# a_19987_42826# 0.016188f
C44424 a_13467_32519# a_14097_32519# 0.048755f
C44425 a_4361_42308# a_22400_42852# 4.45e-21
C44426 a_19237_31679# a_18194_35068# 7.27e-20
C44427 a_3626_43646# a_11633_42308# 9.09e-19
C44428 a_11967_42832# VDD 2.67441f
C44429 a_526_44458# a_5755_42852# 0.054788f
C44430 a_3090_45724# a_4933_42558# 1.87e-19
C44431 a_11823_42460# a_2982_43646# 9.47e-19
C44432 a_4223_44672# a_5205_44734# 7.73e-19
C44433 a_n357_42282# a_16547_43609# 0.004365f
C44434 a_n2956_39768# a_n2216_39866# 0.001489f
C44435 a_14539_43914# a_16979_44734# 0.132799f
C44436 a_626_44172# a_644_44056# 0.126386f
C44437 a_1307_43914# a_453_43940# 0.05952f
C44438 a_n1059_45260# a_17973_43940# 0.004269f
C44439 a_7499_43078# a_6197_43396# 1.44e-19
C44440 a_n2017_45002# a_18079_43940# 1.02e-20
C44441 a_3065_45002# a_n2661_42282# 1.81e-19
C44442 a_16922_45042# a_17517_44484# 0.020096f
C44443 a_17023_45118# a_17061_44734# 1.21e-19
C44444 a_11691_44458# a_13857_44734# 0.049356f
C44445 a_n2661_44458# a_9313_44734# 0.00487f
C44446 a_n2442_46660# a_n4064_39616# 0.224005f
C44447 a_n443_42852# a_12293_43646# 7.27e-19
C44448 a_18780_47178# a_413_45260# 2.11e-19
C44449 a_20820_30879# a_8049_45260# 1.76e-19
C44450 a_n1151_42308# a_375_42282# 1.19e-19
C44451 a_18285_46348# a_16375_45002# 0.003864f
C44452 a_13661_43548# a_18479_45785# 0.087389f
C44453 a_13747_46662# a_18175_45572# 0.03273f
C44454 a_5807_45002# a_18341_45572# 0.0023f
C44455 a_2266_47243# a_2437_43646# 4.08e-19
C44456 a_n2312_40392# a_n2661_45010# 1.45e-20
C44457 a_13507_46334# en_comp 1.11e-19
C44458 a_4915_47217# a_14180_45002# 0.007501f
C44459 a_n743_46660# a_16680_45572# 0.011176f
C44460 a_376_46348# a_835_46155# 6.64e-19
C44461 a_472_46348# a_518_46155# 0.006879f
C44462 a_22223_42860# a_21613_42308# 2.06e-21
C44463 a_1184_42692# a_1149_42558# 1.16e-20
C44464 a_22165_42308# a_22775_42308# 5.13e-19
C44465 a_648_43396# VDD 9.68e-19
C44466 a_n1630_35242# a_1755_42282# 6.88e-21
C44467 a_n784_42308# a_n39_42308# 4.51e-19
C44468 a_1067_42314# a_1606_42308# 0.001471f
C44469 a_3080_42308# VREF_GND 0.001083f
C44470 a_14537_43396# a_14621_43646# 0.004541f
C44471 a_5257_43370# VDD 0.922495f
C44472 a_6540_46812# DATA[3] 1.02e-20
C44473 a_22591_44484# a_19237_31679# 6.8e-19
C44474 a_n913_45002# a_13887_32519# 1.87e-19
C44475 a_n357_42282# a_n3674_37592# 0.327427f
C44476 a_n863_45724# a_1184_42692# 0.563857f
C44477 a_7499_43078# a_10752_42852# 1.98e-19
C44478 a_9313_44734# a_18451_43940# 4.06e-21
C44479 a_17730_32519# a_22959_44484# 0.015145f
C44480 a_6171_45002# a_16664_43396# 9.32e-20
C44481 a_n755_45592# a_n327_42558# 0.003126f
C44482 a_n2661_42834# a_10949_43914# 0.037251f
C44483 a_n2661_43922# a_10729_43914# 1.53e-19
C44484 a_5883_43914# a_9165_43940# 0.019684f
C44485 a_2711_45572# a_19518_43218# 1.67e-19
C44486 a_526_44458# a_10149_42308# 1.05e-19
C44487 a_1423_45028# a_9885_43646# 1.07e-21
C44488 a_n2293_45546# a_n863_45724# 0.17075f
C44489 a_n2438_43548# a_n1699_44726# 3.52e-19
C44490 a_3090_45724# a_1307_43914# 2.66267f
C44491 a_15227_44166# a_13777_45326# 4.73e-20
C44492 a_14976_45028# a_16019_45002# 2.19e-19
C44493 a_n2497_47436# a_n984_44318# 8.35e-19
C44494 a_20202_43084# a_19963_31679# 5.55e-20
C44495 a_5066_45546# a_7499_43078# 0.002848f
C44496 a_n2661_45546# a_n1099_45572# 0.068604f
C44497 a_12549_44172# a_18248_44752# 2.68e-19
C44498 a_14513_46634# a_6171_45002# 1.88e-21
C44499 a_4185_45028# a_18479_45785# 9.87e-21
C44500 a_18285_46348# a_413_45260# 1.46e-20
C44501 a_20820_30879# a_19479_31679# 0.052973f
C44502 a_n1613_43370# a_n23_44458# 2.25e-20
C44503 a_10227_46804# a_14815_43914# 0.004604f
C44504 a_22959_46660# a_2437_43646# 8.36e-21
C44505 a_22591_46660# a_3357_43084# 3.95e-20
C44506 a_11415_45002# a_22591_45572# 0.02488f
C44507 a_15559_46634# a_15415_45028# 3.5e-19
C44508 a_9290_44172# a_8696_44636# 0.032264f
C44509 a_n2293_46634# a_949_44458# 4.57e-19
C44510 a_2324_44458# a_11688_45572# 7.44e-19
C44511 a_n746_45260# a_n237_47217# 0.285294f
C44512 a_n971_45724# a_n23_47502# 0.225828f
C44513 a_n452_47436# a_n785_47204# 0.03755f
C44514 a_n1741_47186# a_1431_47204# 0.014137f
C44515 a_n2109_47186# a_584_46384# 0.352889f
C44516 a_n815_47178# a_327_47204# 1.12e-19
C44517 a_4958_30871# a_n3420_39072# 0.079459f
C44518 a_n1630_35242# VDAC_P 0.00281f
C44519 a_9114_42852# VDD 4.6e-19
C44520 COMP_P a_22521_39511# 1.79e-19
C44521 a_19478_44306# a_19741_43940# 0.005795f
C44522 a_2382_45260# a_3905_42558# 0.002037f
C44523 a_3065_45002# a_3497_42558# 0.002517f
C44524 a_11967_42832# a_16137_43396# 0.300696f
C44525 a_17517_44484# a_15743_43084# 7.31e-22
C44526 a_2253_43940# a_2455_43940# 0.092725f
C44527 a_10555_44260# a_10555_43940# 0.001656f
C44528 a_1337_46116# VDD 0.20087f
C44529 a_n2661_42282# a_458_43396# 7.55e-21
C44530 a_10057_43914# a_10835_43094# 9.83e-19
C44531 a_20205_31679# a_22521_40055# 9e-21
C44532 a_3905_42865# a_6293_42852# 2.22e-20
C44533 a_n913_45002# a_8515_42308# 0.01424f
C44534 a_3537_45260# a_5267_42460# 3.61e-20
C44535 a_6419_46155# a_6298_44484# 4.03e-19
C44536 a_10809_44734# a_20567_45036# 5.98e-22
C44537 a_21137_46414# a_21359_45002# 8.41e-21
C44538 a_17715_44484# a_17801_45144# 2.78e-19
C44539 a_n443_42852# a_327_44734# 0.005815f
C44540 a_1609_45822# a_413_45260# 0.001816f
C44541 a_15037_45618# a_15903_45785# 2.5e-20
C44542 a_5257_43370# a_5495_43940# 0.009999f
C44543 a_19466_46812# a_20159_44458# 1.25e-19
C44544 SMPL_ON_N a_17538_32519# 0.029166f
C44545 a_n971_45724# a_9145_43396# 2.62e-19
C44546 a_2711_45572# a_n913_45002# 3.09e-19
C44547 a_15227_44166# a_20640_44752# 3.05e-21
C44548 a_4791_45118# a_7287_43370# 3.82e-21
C44549 a_n2293_46634# a_11341_43940# 0.487839f
C44550 a_13661_43548# a_14021_43940# 0.103152f
C44551 a_5807_45002# a_14485_44260# 1.16e-20
C44552 a_768_44030# a_3353_43940# 4.43e-19
C44553 a_3090_45724# a_18579_44172# 0.16932f
C44554 a_5937_45572# a_4223_44672# 0.016442f
C44555 a_3483_46348# a_12607_44458# 0.001786f
C44556 a_n755_45592# a_3232_43370# 4.34e-19
C44557 a_8049_45260# a_7639_45394# 2.57e-19
C44558 a_768_44030# a_13759_47204# 5.98e-19
C44559 a_6491_46660# a_5257_43370# 0.1719f
C44560 a_n1435_47204# a_5167_46660# 2.1e-20
C44561 a_n2946_38778# VDD 0.383009f
C44562 a_5088_37509# a_6886_37412# 0.136505f
C44563 a_4338_37500# VDAC_N 0.046178f
C44564 a_n1741_47186# a_11735_46660# 0.029236f
C44565 a_2063_45854# a_6999_46987# 4.27e-21
C44566 a_n3420_39072# VCM 0.007907f
C44567 a_n1151_42308# a_10554_47026# 2.53e-20
C44568 a_6151_47436# a_7715_46873# 0.025823f
C44569 a_3726_37500# a_8912_37509# 0.267651f
C44570 a_18451_43940# a_18599_43230# 2.19e-19
C44571 a_15493_43396# a_18249_42858# 3.35e-20
C44572 a_5891_43370# a_9377_42558# 0.003627f
C44573 a_20974_43370# a_17364_32525# 0.002207f
C44574 a_8685_43396# a_13667_43396# 0.005337f
C44575 a_11341_43940# a_5342_30871# 8.14e-20
C44576 a_17538_32519# a_22959_43396# 4.74e-19
C44577 a_3626_43646# a_17499_43370# 4.06e-20
C44578 a_20273_45572# VDD 0.571099f
C44579 a_8791_43396# a_8945_43396# 0.004009f
C44580 a_11967_42832# a_n784_42308# 4.29e-21
C44581 a_n2293_43922# a_6171_42473# 3.54e-20
C44582 a_6171_45002# a_11963_45334# 0.005724f
C44583 a_n357_42282# a_14673_44172# 4.84e-20
C44584 a_2274_45254# a_1307_43914# 1.47e-19
C44585 a_7229_43940# a_8953_45002# 7.01e-19
C44586 a_6709_45028# a_8191_45002# 9.89e-20
C44587 a_15861_45028# a_17801_45144# 4.92e-20
C44588 a_13527_45546# a_13720_44458# 3.69e-21
C44589 a_10193_42453# a_18989_43940# 0.003937f
C44590 a_327_44734# a_375_42282# 0.067169f
C44591 a_413_45260# a_501_45348# 1.71e-19
C44592 a_18479_45785# a_18587_45118# 0.003753f
C44593 a_18341_45572# a_18315_45260# 3.86e-19
C44594 a_18175_45572# a_18911_45144# 7.25e-20
C44595 a_13507_46334# a_22165_42308# 0.126777f
C44596 a_4185_45028# a_14021_43940# 0.038946f
C44597 a_n2438_43548# a_n2157_42858# 0.266513f
C44598 a_3090_45724# a_9396_43370# 0.003506f
C44599 a_2324_44458# a_12429_44172# 1.55e-21
C44600 a_5111_44636# a_9482_43914# 2.65e-19
C44601 a_11823_42460# a_14539_43914# 1.51e-19
C44602 a_4791_45118# a_5210_46155# 6.75e-22
C44603 a_768_44030# a_2521_46116# 0.008186f
C44604 a_2959_46660# a_765_45546# 0.002438f
C44605 a_6755_46942# a_12816_46660# 0.061031f
C44606 a_4883_46098# a_15015_46420# 0.010147f
C44607 a_18479_47436# a_19553_46090# 1.71e-19
C44608 a_16241_47178# a_10809_44734# 7.12e-21
C44609 a_16023_47582# a_6945_45028# 0.00884f
C44610 a_13507_46334# a_2324_44458# 0.033576f
C44611 a_10227_46804# a_20075_46420# 1.19e-20
C44612 a_n881_46662# a_5204_45822# 0.089827f
C44613 a_18597_46090# a_18819_46122# 0.230891f
C44614 a_12465_44636# a_14493_46090# 0.008365f
C44615 a_11453_44696# a_12594_46348# 2.02e-20
C44616 a_n1613_43370# a_5497_46414# 0.003931f
C44617 a_7871_42858# a_7765_42852# 0.379881f
C44618 a_13467_32519# a_22959_42860# 2.89e-21
C44619 a_14579_43548# a_15597_42852# 9.38e-19
C44620 a_15493_43940# a_19647_42308# 1.44e-21
C44621 a_11341_43940# a_20107_42308# 2.35e-21
C44622 a_n97_42460# a_6171_42473# 1.26e-20
C44623 a_1891_43646# a_1606_42308# 1.3e-20
C44624 a_12281_43396# a_13291_42460# 6.57e-21
C44625 a_5649_42852# a_21195_42852# 5.03e-19
C44626 a_13678_32519# a_21671_42860# 0.014189f
C44627 a_18989_43940# VDD 0.342796f
C44628 a_1307_43914# a_14815_43914# 0.008091f
C44629 a_15765_45572# a_15682_43940# 8.25e-19
C44630 a_n2661_45010# a_n2472_43914# 1.79e-21
C44631 a_n863_45724# a_2896_43646# 1.77e-20
C44632 a_1423_45028# a_n2661_43922# 0.099477f
C44633 SMPL_ON_N a_22465_38105# 0.001357f
C44634 a_n755_45592# a_4905_42826# 7.37e-20
C44635 a_n357_42282# a_766_43646# 0.004396f
C44636 a_8696_44636# a_10807_43548# 1.09e-19
C44637 a_5807_45002# a_10193_42453# 5.69e-19
C44638 a_11735_46660# a_10586_45546# 0.001215f
C44639 a_n2497_47436# a_n467_45028# 2.36e-19
C44640 a_n971_45724# a_n1059_45260# 0.322275f
C44641 a_n746_45260# a_n2017_45002# 2.03e-19
C44642 a_2107_46812# a_2711_45572# 0.034922f
C44643 a_n2293_46634# a_1990_45572# 1.08e-19
C44644 a_13507_46334# a_16855_45546# 2.29e-21
C44645 a_n743_46660# a_6598_45938# 0.001817f
C44646 a_12549_44172# a_13527_45546# 0.09647f
C44647 a_768_44030# a_13163_45724# 3.17e-20
C44648 a_19123_46287# a_18819_46122# 0.172712f
C44649 a_18285_46348# a_18985_46122# 5.57e-21
C44650 a_16721_46634# a_10809_44734# 0.004449f
C44651 a_1138_42852# a_167_45260# 0.250282f
C44652 a_1823_45246# a_2202_46116# 0.25354f
C44653 SMPL_ON_P a_n2956_37592# 0.03953f
C44654 a_1799_45572# a_2307_45899# 1.33e-19
C44655 a_n1925_46634# a_3775_45552# 4.34e-21
C44656 a_11599_46634# a_18175_45572# 0.844188f
C44657 a_11453_44696# a_15037_45618# 1.16e-20
C44658 a_12861_44030# a_18691_45572# 0.007387f
C44659 a_n1151_42308# a_2437_43646# 0.036608f
C44660 a_5745_43940# VDD 0.144352f
C44661 a_5534_30871# a_5742_30871# 0.069311f
C44662 a_12089_42308# a_13249_42558# 2.78e-19
C44663 a_12895_43230# a_13070_42354# 0.006332f
C44664 a_20193_45348# a_22223_43948# 0.041425f
C44665 a_11691_44458# a_15493_43940# 4.95e-19
C44666 a_20202_43084# a_7174_31319# 5.3e-20
C44667 a_20820_30879# a_13258_32519# 0.056725f
C44668 a_5147_45002# a_6293_42852# 8.04e-19
C44669 a_5111_44636# a_6031_43396# 0.207345f
C44670 a_4185_45028# a_15764_42576# 1.97e-19
C44671 a_5807_45002# VDD 1.75047f
C44672 a_4223_44672# a_8333_44056# 0.122173f
C44673 a_3537_45260# a_6547_43396# 0.03331f
C44674 a_12891_46348# CLK 8.04e-20
C44675 a_n357_42282# a_8292_43218# 0.002687f
C44676 a_18587_45118# a_14021_43940# 6.84e-23
C44677 a_n1925_42282# a_n1630_35242# 0.049072f
C44678 a_n443_42852# a_133_42852# 0.004247f
C44679 a_7499_43078# a_10922_42852# 0.008102f
C44680 a_5257_43370# a_5691_45260# 0.009554f
C44681 a_3483_46348# a_8746_45002# 0.605995f
C44682 a_12861_44030# a_12883_44458# 0.041056f
C44683 SMPL_ON_N a_19721_31679# 0.029197f
C44684 a_5807_45002# a_14309_45348# 7.13e-19
C44685 a_13661_43548# a_13711_45394# 4.59e-20
C44686 a_n2497_47436# a_n2661_43922# 0.095407f
C44687 a_12549_44172# a_16922_45042# 0.803336f
C44688 a_2063_45854# a_7640_43914# 1.19e-20
C44689 a_19692_46634# a_20841_45814# 0.003435f
C44690 a_19466_46812# a_20623_45572# 2.08e-19
C44691 a_14493_46090# a_2711_45572# 7.68e-21
C44692 a_1799_45572# a_1423_45028# 2.07e-20
C44693 a_12379_46436# a_12638_46436# 0.093752f
C44694 a_n443_46116# a_n356_44636# 0.004124f
C44695 a_10249_46116# a_413_45260# 4.88e-20
C44696 a_n1925_42282# a_n2661_45546# 0.181908f
C44697 a_12465_44636# a_n2661_44458# 3.22e-19
C44698 a_12991_46634# a_3357_43084# 5.11e-20
C44699 a_n4318_38216# a_n4334_38304# 0.081663f
C44700 a_5342_30871# C1_P_btm 9.04e-20
C44701 a_5534_30871# C0_dummy_P_btm 2.22e-20
C44702 a_15486_42560# a_4958_30871# 0.004787f
C44703 a_14113_42308# a_17531_42308# 8.59e-20
C44704 COMP_P a_1177_38525# 2.71e-19
C44705 a_15764_42576# a_16269_42308# 2.28e-19
C44706 a_n3674_38680# a_n3690_38304# 3.4e-19
C44707 a_10518_42984# VDD 0.273357f
C44708 a_5495_43940# a_5745_43940# 0.014406f
C44709 a_17767_44458# a_17499_43370# 6.82e-20
C44710 a_375_42282# a_133_42852# 0.005083f
C44711 a_11823_42460# a_11897_42308# 0.00139f
C44712 a_n2810_45572# a_n3565_38502# 0.409424f
C44713 a_n2017_45002# a_17749_42852# 0.00371f
C44714 a_n1059_45260# a_17665_42852# 8.77e-19
C44715 a_3699_46348# VDD 0.208984f
C44716 a_14955_43940# a_15493_43396# 2.56e-19
C44717 a_17973_43940# a_18326_43940# 0.009992f
C44718 a_16979_44734# a_17324_43396# 1.03e-19
C44719 a_18114_32519# a_17364_32525# 0.052488f
C44720 a_167_45260# DATA[1] 1.13e-20
C44721 a_20447_31679# a_22400_42852# 5.3e-20
C44722 a_22959_44484# a_17538_32519# 9.27e-19
C44723 a_9313_44734# a_9145_43396# 0.021257f
C44724 a_18597_46090# a_11341_43940# 0.033543f
C44725 a_13507_46334# a_19862_44208# 5.48e-20
C44726 a_5164_46348# a_n2661_43370# 0.010428f
C44727 a_3483_46348# a_14403_45348# 2.17e-20
C44728 a_5807_45002# a_5495_43940# 3.78e-19
C44729 a_18479_47436# a_15493_43940# 0.05409f
C44730 a_5937_45572# a_n2293_42834# 0.097247f
C44731 a_8199_44636# a_8137_45348# 1.55e-21
C44732 a_n2438_43548# a_n1761_44111# 0.001148f
C44733 a_12741_44636# a_11691_44458# 0.81445f
C44734 a_n2497_47436# a_n447_43370# 0.192476f
C44735 SMPL_ON_P a_n2267_43396# 0.001234f
C44736 a_n971_45724# a_n2840_43370# 3.49e-20
C44737 a_11962_45724# a_12791_45546# 0.124167f
C44738 a_12427_45724# a_11823_42460# 0.17307f
C44739 a_2711_45572# a_15903_45785# 0.028735f
C44740 a_5066_45546# a_4558_45348# 0.009388f
C44741 a_11453_44696# a_17737_43940# 2.12e-20
C44742 a_n4064_38528# a_n4064_37440# 0.045121f
C44743 a_n4209_39590# a_n1532_35090# 1.12e-19
C44744 a_n1151_42308# a_n2661_46634# 0.832521f
C44745 a_6151_47436# a_13747_46662# 1.38e-19
C44746 a_6491_46660# a_5807_45002# 0.01567f
C44747 a_n1435_47204# a_12549_44172# 0.072753f
C44748 a_13717_47436# a_12891_46348# 3.83e-20
C44749 a_13381_47204# a_768_44030# 5.3e-20
C44750 a_4958_30871# C10_N_btm 6.95e-19
C44751 a_7174_31319# C3_P_btm 3.5e-20
C44752 a_n2833_47464# a_n2661_46098# 1.96e-20
C44753 a_n2497_47436# a_1799_45572# 1.83e-20
C44754 a_1239_47204# a_n2438_43548# 1.77e-19
C44755 a_1431_47204# a_n743_46660# 0.00119f
C44756 a_7754_39964# a_7754_39632# 0.296522f
C44757 a_584_46384# a_n1925_46634# 0.047378f
C44758 a_22223_47212# SMPL_ON_N 0.00103f
C44759 a_12465_44636# a_11453_44696# 0.084038f
C44760 a_n746_45260# a_1123_46634# 4.1e-19
C44761 a_n785_47204# a_33_46660# 0.008206f
C44762 a_n237_47217# a_383_46660# 3.31e-20
C44763 a_n971_45724# a_948_46660# 6.67e-20
C44764 a_n3565_39590# a_n1838_35608# 2.37e-19
C44765 a_16241_47178# a_n881_46662# 1.39e-21
C44766 a_15761_42308# RST_Z 2.8e-20
C44767 a_15493_43940# a_4190_30871# 8.96e-20
C44768 a_11652_45724# DATA[5] 1.16e-19
C44769 a_20512_43084# a_21356_42826# 4.04e-19
C44770 a_18184_42460# a_14113_42308# 1.64e-20
C44771 a_n97_42460# a_3457_43396# 1.01e-19
C44772 a_15143_45578# VDD 0.12071f
C44773 a_9313_44734# a_19273_43230# 2.85e-21
C44774 a_11322_45546# CLK 0.003637f
C44775 a_11341_43940# a_743_42282# 3.35e-20
C44776 a_n2109_45247# a_n2017_45002# 0.193269f
C44777 a_n2840_45002# a_n2810_45028# 0.161831f
C44778 a_n2293_45010# a_n1059_45260# 0.020223f
C44779 a_n2661_45010# a_n745_45366# 1.07e-20
C44780 a_3090_45724# a_10867_43940# 0.00115f
C44781 a_3483_46348# a_5663_43940# 0.00218f
C44782 a_4185_45028# a_5013_44260# 3.66e-19
C44783 a_2277_45546# a_949_44458# 6.13e-20
C44784 a_2711_45572# a_n2661_44458# 3.52e-21
C44785 a_n2293_46098# a_5841_44260# 8.09e-20
C44786 a_13059_46348# a_12710_44260# 1.05e-20
C44787 a_n443_42852# a_4223_44672# 0.001694f
C44788 a_5257_43370# a_3080_42308# 0.00466f
C44789 a_10586_45546# a_10617_44484# 9.55e-19
C44790 a_n2293_46634# a_10341_43396# 2.04894f
C44791 a_12549_44172# a_15743_43084# 0.021095f
C44792 VDD VREF 4.8299f
C44793 C10_N_btm VCM 10.3108f
C44794 a_18479_47436# a_12741_44636# 0.020666f
C44795 a_4646_46812# a_5257_43370# 0.024804f
C44796 a_3877_44458# a_7411_46660# 4.74e-19
C44797 a_19321_45002# a_15227_44166# 0.145462f
C44798 a_12891_46348# a_14035_46660# 1.12e-20
C44799 a_12549_44172# a_13885_46660# 0.036345f
C44800 a_6151_47436# a_4419_46090# 4.28e-20
C44801 a_4817_46660# a_5894_47026# 1.46e-19
C44802 a_2063_45854# a_9823_46155# 3.28e-19
C44803 a_2266_47243# a_765_45546# 3.3e-19
C44804 a_13661_43548# a_19692_46634# 0.093373f
C44805 a_13747_46662# a_19466_46812# 0.869986f
C44806 a_5807_45002# a_10185_46660# 6.99e-19
C44807 a_4915_47217# a_5164_46348# 2.37e-20
C44808 a_n443_46116# a_5204_45822# 0.020803f
C44809 a_4791_45118# a_5497_46414# 0.056648f
C44810 a_n1151_42308# a_8199_44636# 0.161616f
C44811 a_n743_46660# a_11735_46660# 1.24e-19
C44812 a_13507_46334# a_21350_47026# 3.44e-19
C44813 a_11453_44696# a_20528_46660# 0.016145f
C44814 a_10405_44172# a_10533_42308# 2.11e-21
C44815 a_13887_32519# a_17364_32525# 0.050078f
C44816 a_19721_31679# a_19864_35138# 1.22e-21
C44817 a_10341_43396# a_5342_30871# 0.001109f
C44818 a_n97_42460# a_16877_43172# 0.002787f
C44819 a_22591_43396# a_22959_43396# 7.52e-19
C44820 a_18315_45260# VDD 0.12623f
C44821 a_18479_45785# a_11967_42832# 0.038105f
C44822 a_3090_45724# a_13635_43156# 0.00703f
C44823 a_1307_43914# a_4743_44484# 0.011512f
C44824 a_2711_45572# a_18451_43940# 0.010207f
C44825 a_n2661_45010# a_3363_44484# 2.68e-20
C44826 a_20202_43084# a_21487_43396# 0.019942f
C44827 a_n443_42852# a_15493_43940# 0.301211f
C44828 a_9290_44172# a_14205_43396# 0.010382f
C44829 a_526_44458# a_1891_43646# 4.7e-19
C44830 a_3537_45260# a_n356_44636# 4.16e-19
C44831 a_n2312_39304# a_6123_31319# 5.16e-21
C44832 a_n1059_45260# a_9313_44734# 0.089245f
C44833 a_3357_43084# a_n2293_43922# 9.05e-21
C44834 a_9482_43914# a_10334_44484# 0.015932f
C44835 a_626_44172# a_949_44458# 0.006992f
C44836 a_n863_45724# a_1443_43940# 0.005869f
C44837 a_n2956_39768# a_n3674_38680# 0.023454f
C44838 a_10903_43370# a_10695_43548# 0.041719f
C44839 a_3483_46348# a_16243_43396# 0.001863f
C44840 a_4883_46098# a_6472_45840# 4.6e-20
C44841 a_5807_45002# a_20850_46155# 6.12e-21
C44842 a_3090_45724# a_8016_46348# 0.0122f
C44843 a_12861_44030# a_10490_45724# 2.29e-20
C44844 a_3877_44458# a_4365_46436# 9.48e-20
C44845 a_n1151_42308# a_8192_45572# 9.32e-20
C44846 a_6151_47436# a_6469_45572# 6.03e-19
C44847 a_11453_44696# a_2711_45572# 0.033654f
C44848 a_n881_46662# a_3503_45724# 0.001143f
C44849 a_19692_46634# a_4185_45028# 4.25e-20
C44850 a_n1613_43370# a_n356_45724# 4.43e-20
C44851 a_20107_46660# a_20202_43084# 4.38e-20
C44852 a_20841_46902# a_20719_46660# 3.16e-19
C44853 a_11813_46116# a_9290_44172# 4.46e-19
C44854 a_11186_47026# a_11133_46155# 1.37e-19
C44855 a_5649_42852# a_8791_42308# 1.31e-19
C44856 a_16409_43396# a_17124_42282# 1.26e-20
C44857 a_4190_30871# a_5742_30871# 0.029789f
C44858 a_4361_42308# a_9293_42558# 5.9e-20
C44859 a_1847_42826# a_2725_42558# 7.35e-19
C44860 a_18249_42858# a_18707_42852# 0.027606f
C44861 a_10341_43396# a_20107_42308# 2.81e-20
C44862 a_n822_43940# VDD 5.19e-19
C44863 a_10518_42984# a_n784_42308# 2.16e-21
C44864 a_4520_42826# a_1755_42282# 2.93e-20
C44865 a_743_42282# a_10723_42308# 0.008155f
C44866 a_n755_45592# a_2905_42968# 4.85e-20
C44867 a_n357_42282# a_3681_42891# 0.005491f
C44868 a_14311_47204# VDD 0.241476f
C44869 SMPL_ON_N a_18194_35068# 3.71e-19
C44870 a_5891_43370# a_9159_44484# 6.38e-20
C44871 a_16112_44458# a_16241_44484# 0.010132f
C44872 a_3357_43084# a_n97_42460# 0.113127f
C44873 a_18114_32519# a_19237_31679# 8.86333f
C44874 a_526_44458# a_4149_42891# 2.3e-20
C44875 a_9863_47436# DATA[4] 7.9e-19
C44876 a_9482_43914# a_13565_44260# 0.003452f
C44877 a_6109_44484# a_n2661_43922# 0.021636f
C44878 a_7640_43914# a_n2661_42834# 0.030156f
C44879 a_19721_31679# a_22959_44484# 4.31e-19
C44880 a_12861_44030# START 0.006864f
C44881 a_n1435_47204# CLK_DATA 8.83e-21
C44882 a_17970_44736# a_17517_44484# 0.075165f
C44883 a_n2661_45010# a_n2433_43396# 1.83e-20
C44884 a_5691_45260# a_5745_43940# 3.63e-21
C44885 a_13717_47436# SINGLE_ENDED 0.032092f
C44886 a_13487_47204# RST_Z 0.07884f
C44887 a_18819_46122# a_8049_45260# 0.003213f
C44888 a_11387_46155# a_11601_46155# 0.005572f
C44889 a_n2293_46098# a_n356_45724# 0.022803f
C44890 a_376_46348# a_n357_42282# 2.8e-19
C44891 a_n1076_46494# a_n755_45592# 6.77e-20
C44892 a_5807_45002# a_5691_45260# 0.19412f
C44893 a_12741_44636# a_n443_42852# 7.1e-20
C44894 a_n2438_43548# a_n2956_37592# 0.004958f
C44895 a_n2661_46634# a_327_44734# 5.27e-21
C44896 a_n2293_46634# a_n143_45144# 0.00576f
C44897 a_4185_45028# a_20692_30879# 1.35e-19
C44898 a_n2497_47436# a_n452_44636# 0.001121f
C44899 SMPL_ON_P a_n2267_44484# 5.37e-21
C44900 a_472_46348# a_310_45028# 3.57e-19
C44901 a_2698_46116# a_n2661_45546# 9.6e-20
C44902 a_768_44030# a_8953_45002# 3.3e-19
C44903 a_n1021_46688# a_n967_45348# 5.18e-21
C44904 a_6755_46942# a_16223_45938# 0.002064f
C44905 a_1138_42852# a_n863_45724# 0.135594f
C44906 a_13351_46090# a_12638_46436# 0.001216f
C44907 a_2324_44458# a_10586_45546# 0.436403f
C44908 a_8515_42308# a_8325_42308# 0.134955f
C44909 a_5934_30871# a_8685_42308# 0.186981f
C44910 a_4190_30871# C0_dummy_P_btm 1.45e-20
C44911 a_17364_32525# EN_VIN_BSTR_N 0.959329f
C44912 a_16867_43762# VDD 0.132317f
C44913 a_n3674_39768# a_n1644_44306# 1.74e-19
C44914 a_20820_30879# a_22609_37990# 1.17e-20
C44915 a_n2017_45002# a_19339_43156# 0.028127f
C44916 a_n913_45002# a_18817_42826# 2.27e-20
C44917 a_n1059_45260# a_18599_43230# 2.93e-19
C44918 a_3357_43084# a_3935_43218# 2.32e-19
C44919 a_11967_42832# a_14021_43940# 0.030676f
C44920 a_5883_43914# a_6765_43638# 1.3e-19
C44921 a_2479_44172# a_n2661_42282# 3.48e-21
C44922 a_2998_44172# a_3499_42826# 0.027036f
C44923 a_n443_42852# a_5742_30871# 2.05e-19
C44924 a_n356_44636# a_1049_43396# 0.042597f
C44925 a_14226_46987# VDD 6.34e-20
C44926 a_6298_44484# a_7112_43396# 7.71e-19
C44927 a_13259_45724# a_20712_42282# 1.03e-19
C44928 a_n2956_39304# a_n2860_38778# 8.73e-19
C44929 a_n2956_38680# a_n2302_38778# 0.038021f
C44930 a_n357_42282# a_15959_42545# 9.81e-20
C44931 en_comp a_17701_42308# 1.94e-20
C44932 a_14513_46634# RST_Z 1.53e-20
C44933 a_1609_45822# a_2211_45572# 8.16e-20
C44934 a_n2312_38680# a_n2661_42834# 1.97e-21
C44935 a_8049_45260# a_16223_45938# 0.004651f
C44936 a_3483_46348# a_3232_43370# 0.220803f
C44937 a_15227_44166# a_18184_42460# 3.08e-21
C44938 a_14976_45028# a_11827_44484# 7.51e-20
C44939 a_2711_45572# a_5907_45546# 0.01826f
C44940 a_2107_46812# a_9241_44734# 1.31e-19
C44941 a_n2293_46634# a_n2293_43922# 0.02819f
C44942 a_2063_45854# a_10729_43914# 0.004795f
C44943 a_5937_45572# a_413_45260# 4.56e-21
C44944 a_19466_46812# a_18911_45144# 1.84e-19
C44945 a_4185_45028# a_4927_45028# 0.004584f
C44946 a_5164_46348# a_4574_45260# 1.44e-19
C44947 a_5204_45822# a_3537_45260# 2.3e-20
C44948 a_15959_42545# CAL_N 3.77e-19
C44949 a_5934_30871# C10_P_btm 1.89e-19
C44950 a_1343_38525# a_2684_37794# 0.224374f
C44951 a_5932_42308# C3_P_btm 0.121156f
C44952 a_6575_47204# a_n1435_47204# 5.93e-19
C44953 a_11031_47542# a_9313_45822# 0.063846f
C44954 a_n3420_39072# a_n4064_38528# 7.47287f
C44955 a_n2946_39072# a_n2946_38778# 0.050477f
C44956 a_1736_39043# a_2112_39137# 0.554188f
C44957 a_n4064_39072# a_n3420_38528# 0.048218f
C44958 SMPL_ON_P a_n2312_39304# 0.040801f
C44959 a_n1605_47204# a_n2312_40392# 2.12e-19
C44960 a_n1741_47186# a_n310_47570# 5.79e-19
C44961 a_6151_47436# a_11599_46634# 0.008629f
C44962 a_6123_31319# C8_P_btm 6.73e-20
C44963 a_n327_42308# VDD 1.42e-19
C44964 a_n357_42282# RST_Z 2.38e-20
C44965 a_20193_45348# a_20753_42852# 0.04748f
C44966 a_n913_45002# a_21421_42336# 0.001645f
C44967 a_13483_43940# a_13667_43396# 9.11e-19
C44968 a_15493_43396# a_8685_43396# 0.011009f
C44969 a_20205_31679# VCM 0.035399f
C44970 a_20692_30879# VREF_GND 0.010456f
C44971 a_20512_43084# a_20749_43396# 0.008222f
C44972 a_n755_45592# VDD 2.41485f
C44973 en_comp a_21613_42308# 2.05e-20
C44974 a_375_42282# a_5742_30871# 1.69e-20
C44975 a_n2293_43922# a_5342_30871# 1.2e-20
C44976 a_9313_44734# a_19987_42826# 0.009103f
C44977 a_22485_44484# a_17364_32525# 1e-18
C44978 a_19237_31679# a_13887_32519# 0.052352f
C44979 a_17730_32519# a_14209_32519# 0.054558f
C44980 a_10227_46804# a_12281_43396# 6.09e-20
C44981 a_12861_44030# a_16547_43609# 3.22e-19
C44982 a_6755_46942# a_11341_43940# 3.7e-19
C44983 a_11322_45546# a_10951_45334# 4.5e-19
C44984 a_2711_45572# a_6125_45348# 7.07e-19
C44985 a_n2293_46634# a_n97_42460# 0.108602f
C44986 a_9049_44484# a_9482_43914# 3.58e-19
C44987 a_768_44030# a_3626_43646# 0.002415f
C44988 a_n1613_43370# a_6547_43396# 0.154311f
C44989 a_18597_46090# a_10341_43396# 0.027979f
C44990 a_n2497_47436# a_n1641_43230# 0.001225f
C44991 SMPL_ON_P a_n2472_42826# 3.03e-19
C44992 a_n2438_43548# a_n2267_43396# 0.120634f
C44993 a_3316_45546# a_n2661_43370# 0.022024f
C44994 a_16375_45002# a_11691_44458# 1.43e-19
C44995 a_20202_43084# a_21398_44850# 4.42e-20
C44996 a_11415_45002# a_20980_44850# 0.00141f
C44997 a_18691_45572# a_18787_45572# 0.013793f
C44998 a_18909_45814# a_18953_45572# 3.69e-19
C44999 a_18479_45785# a_20273_45572# 1.17e-20
C45000 a_12465_44636# a_9145_43396# 9.6e-20
C45001 a_4883_46098# a_10695_43548# 3.82e-20
C45002 a_13249_42308# a_6171_45002# 0.026329f
C45003 a_9290_44172# a_9159_44484# 7.16e-20
C45004 a_10193_42453# a_13017_45260# 5.13e-21
C45005 a_n443_42852# a_n2293_42834# 1.60683f
C45006 a_10490_45724# a_11787_45002# 1.44e-19
C45007 a_n4064_37440# VREF_GND 0.048151f
C45008 a_16327_47482# a_16292_46812# 0.027563f
C45009 a_n133_46660# a_288_46660# 0.086708f
C45010 a_n743_46660# a_n935_46688# 0.001334f
C45011 a_n2438_43548# a_491_47026# 8.49e-19
C45012 EN_VIN_BSTR_N a_21589_35634# 2.66e-19
C45013 a_22521_40599# VDD 0.804442f
C45014 a_18194_35068# a_19864_35138# 0.045378f
C45015 CAL_N RST_Z 0.058301f
C45016 a_11599_46634# a_19466_46812# 0.453656f
C45017 a_n1925_46634# a_479_46660# 8.56e-19
C45018 a_n2661_46634# a_3177_46902# 0.00699f
C45019 a_5807_45002# a_4646_46812# 0.032485f
C45020 a_n881_46662# a_7927_46660# 0.017621f
C45021 a_10227_46804# a_15009_46634# 0.02057f
C45022 a_17591_47464# a_3090_45724# 5.31e-19
C45023 EN_VIN_BSTR_P C8_P_btm 0.090252f
C45024 a_n1151_42308# a_765_45546# 1.7705f
C45025 a_8128_46384# a_7411_46660# 0.019875f
C45026 a_n2293_46634# a_n2661_46098# 0.022053f
C45027 a_601_46902# a_948_46660# 0.051162f
C45028 a_14358_43442# a_4361_42308# 1.13e-20
C45029 a_15781_43660# a_15868_43402# 0.004898f
C45030 a_10341_43396# a_743_42282# 0.017833f
C45031 a_21381_43940# a_21356_42826# 0.196864f
C45032 a_16243_43396# a_16664_43396# 0.090164f
C45033 a_13017_45260# VDD 0.263701f
C45034 a_n97_42460# a_5342_30871# 0.068562f
C45035 a_16977_43638# a_15743_43084# 0.042866f
C45036 a_17324_43396# a_18429_43548# 1.43e-19
C45037 a_17499_43370# a_18525_43370# 1.4e-19
C45038 a_n2661_42282# a_n2104_42282# 4.14e-19
C45039 a_11967_42832# a_15764_42576# 0.012941f
C45040 a_2982_43646# a_7871_42858# 4.24e-20
C45041 a_3626_43646# a_5755_42852# 1.23e-20
C45042 a_n2312_38680# a_n2293_42282# 3.75e-20
C45043 a_375_42282# a_n2293_42834# 0.027465f
C45044 a_13348_45260# a_13490_45394# 0.007833f
C45045 a_13017_45260# a_14309_45348# 0.002224f
C45046 a_13249_42308# a_14673_44172# 0.026424f
C45047 a_4185_45028# a_4699_43561# 0.010947f
C45048 a_8696_44636# a_8375_44464# 0.006586f
C45049 a_n443_42852# a_1115_44172# 4.54e-19
C45050 a_6171_45002# a_17613_45144# 3.24e-19
C45051 a_n2472_45002# a_n2661_44458# 0.002026f
C45052 a_n2661_45010# a_n2433_44484# 0.217176f
C45053 a_2809_45348# a_2809_45028# 6.96e-20
C45054 a_1823_45246# a_2982_43646# 0.022597f
C45055 a_15227_44166# a_15868_43402# 3.62e-19
C45056 a_3357_43084# a_742_44458# 7.16e-19
C45057 a_18479_45785# a_18989_43940# 3.49e-19
C45058 a_18691_45572# a_18287_44626# 1.75e-20
C45059 a_18341_45572# a_18374_44850# 7.8e-19
C45060 a_18909_45814# a_18443_44721# 5.48e-20
C45061 a_n357_42282# a_5663_43940# 1.55e-19
C45062 a_3316_45546# a_2998_44172# 4.99e-19
C45063 a_4791_45118# a_5267_42460# 0.138738f
C45064 a_18479_47436# a_16375_45002# 2.07e-21
C45065 a_18597_46090# a_18147_46436# 5.21e-20
C45066 a_16327_47482# a_20254_46482# 0.001965f
C45067 a_n971_45724# a_5263_45724# 1.03e-20
C45068 a_n443_46116# a_3503_45724# 1.86e-19
C45069 a_n881_46662# a_6419_46482# 3.32e-21
C45070 a_14084_46812# a_765_45546# 7.01e-21
C45071 a_3090_45724# a_15312_46660# 9.66e-19
C45072 a_20916_46384# a_21137_46414# 0.118131f
C45073 a_19594_46812# a_10809_44734# 0.042242f
C45074 a_16750_47204# a_6945_45028# 7.64e-20
C45075 a_2063_45854# a_2307_45899# 4.37e-19
C45076 a_3877_44458# a_4185_45028# 0.338483f
C45077 a_15227_44166# a_13059_46348# 5.76e-19
C45078 a_n1613_43370# a_6640_46482# 7.81e-19
C45079 a_16292_46812# a_16434_46987# 0.005572f
C45080 a_n743_46660# a_2324_44458# 0.036195f
C45081 a_743_42282# a_20356_42852# 0.001934f
C45082 a_3422_30871# C4_P_btm 1.36e-19
C45083 a_19339_43156# a_19164_43230# 0.233657f
C45084 a_13467_32519# a_22400_42852# 0.029855f
C45085 a_19237_31679# EN_VIN_BSTR_N 0.069167f
C45086 a_3626_43646# a_10149_42308# 5.71e-19
C45087 a_7227_42852# a_7309_42852# 0.171361f
C45088 a_19006_44850# VDD 0.077608f
C45089 a_526_44458# a_5111_42852# 0.265994f
C45090 a_n1925_42282# a_4520_42826# 6.4e-19
C45091 a_2437_43646# a_15493_43940# 1.05e-21
C45092 a_21297_45572# a_19862_44208# 3.66e-20
C45093 a_11827_44484# a_15433_44458# 0.002592f
C45094 a_n357_42282# a_16243_43396# 1.3e-19
C45095 a_n2956_39768# a_n2860_39866# 0.001355f
C45096 a_7499_43078# a_6293_42852# 1.55e-20
C45097 a_626_44172# a_175_44278# 0.017096f
C45098 a_3537_45260# a_3820_44260# 0.001488f
C45099 a_n1059_45260# a_17737_43940# 6.9e-19
C45100 a_1307_43914# a_1414_42308# 0.147738f
C45101 a_n2661_44458# a_9241_44734# 2.59e-19
C45102 a_11691_44458# a_13468_44734# 0.004179f
C45103 a_n2442_46660# a_n2946_39866# 0.024649f
C45104 a_n2312_38680# a_n3565_39590# 0.031736f
C45105 a_18479_47436# a_413_45260# 2.86e-19
C45106 a_10903_43370# a_14275_46494# 3.08e-20
C45107 a_2063_45854# a_1423_45028# 4.66e-20
C45108 a_1138_42852# a_1431_46436# 6.23e-19
C45109 a_4915_47217# a_13777_45326# 8.78e-22
C45110 a_18285_46348# a_18243_46436# 0.002179f
C45111 a_17829_46910# a_16375_45002# 1.99e-19
C45112 a_13661_43548# a_18175_45572# 0.029369f
C45113 a_5807_45002# a_18479_45785# 0.174313f
C45114 a_13747_46662# a_16147_45260# 0.027471f
C45115 a_12549_44172# a_17668_45572# 5.63e-20
C45116 a_12861_44030# a_6171_45002# 0.05507f
C45117 a_3315_47570# a_2437_43646# 8.57e-19
C45118 a_n743_46660# a_16855_45546# 0.005475f
C45119 a_376_46348# a_518_46155# 0.005572f
C45120 a_11189_46129# a_2324_44458# 2.84e-19
C45121 a_13351_46090# a_13759_46122# 0.043782f
C45122 a_564_42282# a_1755_42282# 2.36e-20
C45123 a_22165_42308# a_21613_42308# 0.027246f
C45124 a_1184_42692# a_961_42354# 0.100246f
C45125 a_548_43396# VDD 4.01e-19
C45126 a_n784_42308# a_n327_42308# 1.52e-19
C45127 a_n1630_35242# a_1606_42308# 0.032246f
C45128 a_1067_42314# a_1221_42558# 0.008535f
C45129 a_n2661_43370# a_6197_43396# 5.24e-22
C45130 a_14537_43396# a_14537_43646# 0.003096f
C45131 a_18989_43940# a_14021_43940# 5.23e-19
C45132 a_n913_45002# a_22223_43396# 2.71e-20
C45133 a_n863_45724# a_1576_42282# 0.05148f
C45134 a_1307_43914# a_12281_43396# 1.31e-19
C45135 a_9313_44734# a_18326_43940# 1.97e-20
C45136 a_22591_44484# a_22959_44484# 7.52e-19
C45137 a_22485_44484# a_19237_31679# 3.62e-20
C45138 en_comp a_4361_42308# 2.27e-19
C45139 a_n2661_42834# a_10729_43914# 0.01161f
C45140 a_n2661_43922# a_10405_44172# 2.51e-20
C45141 a_5883_43914# a_8487_44056# 6.48e-19
C45142 a_n755_45592# a_n784_42308# 0.711298f
C45143 a_n357_42282# a_n327_42558# 0.006254f
C45144 a_n2438_43548# a_n2267_44484# 0.120608f
C45145 a_n2956_38216# a_n863_45724# 0.001226f
C45146 a_3090_45724# a_16019_45002# 3.78e-20
C45147 a_15227_44166# a_13556_45296# 0.047404f
C45148 a_14976_45028# a_15595_45028# 3.96e-19
C45149 a_n2497_47436# a_n809_44244# 0.029871f
C45150 a_5066_45546# a_8568_45546# 0.04527f
C45151 a_n2661_45546# a_380_45546# 0.012814f
C45152 a_n2810_45572# a_n1099_45572# 0.001228f
C45153 a_12549_44172# a_17970_44736# 3.76e-20
C45154 a_n1613_43370# a_n356_44636# 5.31e-19
C45155 a_10227_46804# a_14112_44734# 1.24e-19
C45156 SMPL_ON_N a_9313_44734# 2.16e-20
C45157 a_12741_44636# a_2437_43646# 0.023858f
C45158 a_11415_45002# a_3357_43084# 0.053912f
C45159 a_765_45546# a_327_44734# 5.49e-20
C45160 a_12861_44030# a_14673_44172# 0.015418f
C45161 a_15368_46634# a_15415_45028# 2.5e-19
C45162 a_n2293_46634# a_742_44458# 2.95e-19
C45163 a_n2293_45546# a_n1079_45724# 5.25e-19
C45164 a_14180_46482# a_2711_45572# 3.42e-20
C45165 a_5742_30871# a_n3420_37984# 0.004679f
C45166 a_7174_31319# a_n3565_39590# 5.27e-21
C45167 a_n2497_47436# a_2063_45854# 4e-20
C45168 a_n815_47178# a_n785_47204# 0.123817f
C45169 a_n971_45724# a_n237_47217# 0.134971f
C45170 a_n1741_47186# a_1239_47204# 0.022889f
C45171 a_n2109_47186# a_2124_47436# 0.037038f
C45172 a_2382_45260# a_3581_42558# 0.001326f
C45173 a_17517_44484# a_18783_43370# 9.36e-21
C45174 a_20365_43914# a_19319_43548# 0.007317f
C45175 a_11341_43940# a_15037_43940# 0.00577f
C45176 a_835_46155# VDD 7.28e-19
C45177 a_3499_42826# a_1568_43370# 3.66e-21
C45178 a_9313_44734# a_22959_43396# 0.002204f
C45179 a_n2293_43922# a_743_42282# 0.034167f
C45180 a_10057_43914# a_10518_42984# 4.8e-19
C45181 a_8975_43940# a_10083_42826# 5.33e-21
C45182 a_20692_30879# a_22469_40625# 2.12e-20
C45183 a_3905_42865# a_6031_43396# 4.79e-21
C45184 a_n1059_45260# a_8515_42308# 1.02e-20
C45185 a_n913_45002# a_5934_30871# 0.126791f
C45186 a_19862_44208# a_19478_44056# 4.77e-20
C45187 a_3537_45260# a_3823_42558# 2.53e-21
C45188 a_19900_46494# a_11827_44484# 1.49e-22
C45189 a_21137_46414# a_21101_45002# 1.79e-19
C45190 a_6165_46155# a_6298_44484# 2.52e-20
C45191 a_3503_45724# a_3537_45260# 0.00137f
C45192 a_3483_46348# a_8975_43940# 0.016137f
C45193 a_n443_42852# a_413_45260# 0.005091f
C45194 a_509_45822# a_327_44734# 5.3e-20
C45195 a_15037_45618# a_15599_45572# 6.39e-21
C45196 a_5257_43370# a_5013_44260# 0.002385f
C45197 a_n971_45724# a_8423_43396# 0.001593f
C45198 a_10809_44734# a_18494_42460# 8.81e-22
C45199 a_2711_45572# a_n1059_45260# 2.83e-19
C45200 a_19692_46634# a_11967_42832# 0.032909f
C45201 a_15227_44166# a_20362_44736# 4.57e-21
C45202 a_19466_46812# a_19615_44636# 3.92e-20
C45203 a_5807_45002# a_14021_43940# 0.001299f
C45204 a_13661_43548# a_13829_44260# 0.001195f
C45205 a_768_44030# a_3052_44056# 1.06e-19
C45206 a_n1613_43370# a_9165_43940# 2.36e-20
C45207 a_8199_44636# a_4223_44672# 4.87e-19
C45208 a_n357_42282# a_3232_43370# 4.05e-19
C45209 a_18985_46122# a_11691_44458# 2.44e-22
C45210 a_5066_45546# a_n2661_43370# 4.51e-19
C45211 a_768_44030# a_13675_47204# 5.16e-20
C45212 a_12549_44172# a_13759_47204# 3.89e-19
C45213 a_9804_47204# a_5807_45002# 0.039093f
C45214 a_6151_47436# a_7411_46660# 0.330209f
C45215 a_n1435_47204# a_5385_46902# 3.12e-20
C45216 a_6545_47178# a_5257_43370# 8.38e-19
C45217 a_n2312_39304# a_n2438_43548# 0.052323f
C45218 a_n3420_38528# VDD 0.522772f
C45219 a_4338_37500# a_6886_37412# 1.95816f
C45220 a_3726_37500# VDAC_N 0.06247f
C45221 a_n971_45724# a_8270_45546# 0.251101f
C45222 a_n237_47217# a_8023_46660# 1.98e-19
C45223 a_2063_45854# a_6682_46987# 8.35e-21
C45224 a_5088_37509# a_5700_37509# 1.48771f
C45225 a_n3420_39072# VREF_GND 0.066097f
C45226 a_n1151_42308# a_10623_46897# 1.42e-19
C45227 a_4915_47217# a_8145_46902# 5.23e-20
C45228 a_n4064_37984# C1_P_btm 8.65e-20
C45229 a_2982_43646# a_17324_43396# 2.59e-21
C45230 a_18451_43940# a_18817_42826# 4.37e-22
C45231 a_15493_43396# a_17333_42852# 1.04e-20
C45232 a_8791_43396# a_8873_43396# 0.005167f
C45233 a_n97_42460# a_743_42282# 0.107736f
C45234 a_5891_43370# a_9293_42558# 0.001253f
C45235 a_14401_32519# a_17364_32525# 7.51978f
C45236 a_8685_43396# a_10695_43548# 0.00269f
C45237 a_17538_32519# a_14209_32519# 0.051332f
C45238 a_20107_45572# VDD 0.458237f
C45239 a_3422_30871# a_14097_32519# 0.031284f
C45240 a_22315_44484# a_22400_42852# 1.35e-22
C45241 a_n2293_43922# a_5755_42308# 8.6e-20
C45242 a_6171_45002# a_11787_45002# 0.01986f
C45243 a_6709_45028# a_7705_45326# 0.099282f
C45244 a_7229_43940# a_8191_45002# 6.79e-19
C45245 a_15861_45028# a_16981_45144# 9.5e-19
C45246 a_6755_46942# a_10341_43396# 8.9e-20
C45247 a_13527_45546# a_13076_44458# 2.47e-21
C45248 a_13249_42308# a_12607_44458# 3.94e-19
C45249 a_10193_42453# a_18374_44850# 1.66e-20
C45250 a_413_45260# a_375_42282# 0.112554f
C45251 a_18479_45785# a_18315_45260# 3.67e-19
C45252 a_18175_45572# a_18587_45118# 0.003125f
C45253 a_13507_46334# a_21671_42860# 0.001831f
C45254 a_n2956_39768# a_n4318_38680# 0.023624f
C45255 a_768_44030# a_8037_42858# 4.29e-23
C45256 a_n2438_43548# a_n2472_42826# 0.026866f
C45257 a_3090_45724# a_8791_43396# 0.00173f
C45258 a_19431_45546# a_16922_45042# 2.16e-20
C45259 a_2324_44458# a_11750_44172# 4.42e-21
C45260 a_526_44458# a_7542_44172# 7.82e-21
C45261 a_4791_45118# a_6640_46482# 0.001342f
C45262 a_768_44030# a_167_45260# 0.014856f
C45263 a_3177_46902# a_765_45546# 0.001508f
C45264 a_6755_46942# a_12991_46634# 0.077634f
C45265 a_10249_46116# a_12816_46660# 4.52e-20
C45266 a_11453_44696# a_12005_46116# 4.21e-21
C45267 a_4883_46098# a_14275_46494# 0.006919f
C45268 a_18479_47436# a_18985_46122# 2.08e-19
C45269 a_18780_47178# a_18819_46122# 1.69e-19
C45270 a_16327_47482# a_6945_45028# 0.111399f
C45271 a_n1741_47186# a_12839_46116# 0.113988f
C45272 a_n2661_46634# a_12741_44636# 2.1e-19
C45273 a_13507_46334# a_14840_46494# 0.005149f
C45274 a_10227_46804# a_19335_46494# 8.56e-21
C45275 a_15673_47210# a_10809_44734# 4.01e-20
C45276 a_2063_45854# a_9823_46482# 1.18e-21
C45277 a_n1435_47204# a_n1533_46116# 3.18e-20
C45278 a_n2293_46634# a_11415_45002# 0.001066f
C45279 a_18597_46090# a_17957_46116# 0.018356f
C45280 a_12465_44636# a_13925_46122# 0.018086f
C45281 a_n1613_43370# a_5204_45822# 0.002482f
C45282 a_n881_46662# a_5164_46348# 0.03104f
C45283 a_7227_42852# a_7765_42852# 0.118623f
C45284 a_13467_32519# a_22223_42860# 3.77e-19
C45285 a_4361_42308# a_22165_42308# 1.92e-21
C45286 a_14579_43548# a_14853_42852# 0.002493f
C45287 a_15493_43940# a_19511_42282# 1.21e-21
C45288 a_n97_42460# a_5755_42308# 0.009194f
C45289 a_1427_43646# a_1606_42308# 6.56e-20
C45290 a_5649_42852# a_21356_42826# 1.42e-20
C45291 a_13678_32519# a_21195_42852# 0.001094f
C45292 a_21855_43396# a_21671_42860# 3.61e-19
C45293 a_18374_44850# VDD 0.203584f
C45294 a_7499_43078# a_7499_43940# 0.003097f
C45295 a_15903_45785# a_15682_43940# 1.25e-19
C45296 a_n913_45002# a_20512_43084# 1.33e-19
C45297 a_1423_45028# a_n2661_42834# 1e-18
C45298 a_n2293_46634# a_10533_42308# 2.12e-21
C45299 a_3090_45724# a_13814_43218# 2.67e-19
C45300 a_8696_44636# a_10949_43914# 4.65e-20
C45301 a_n2661_45546# a_3539_42460# 0.091495f
C45302 a_n755_45592# a_3080_42308# 0.237742f
C45303 a_n357_42282# a_4905_42826# 0.026713f
C45304 a_n1925_46634# a_7227_45028# 5.87e-19
C45305 a_4646_46812# a_n755_45592# 8.29e-20
C45306 a_5807_45002# a_10180_45724# 6.9e-20
C45307 a_n2293_46098# a_5204_45822# 0.008417f
C45308 a_n971_45724# a_n2017_45002# 0.048447f
C45309 a_n746_45260# a_n2109_45247# 1.91e-20
C45310 SMPL_ON_P a_n2810_45028# 0.039597f
C45311 a_12991_46634# a_8049_45260# 1.12e-20
C45312 a_n2661_46098# a_2277_45546# 5.6e-20
C45313 a_n743_46660# a_6667_45809# 0.001764f
C45314 a_12891_46348# a_13527_45546# 0.002777f
C45315 a_12549_44172# a_13163_45724# 0.172293f
C45316 a_19123_46287# a_17957_46116# 2.21e-20
C45317 a_18285_46348# a_18819_46122# 1.08e-19
C45318 a_16388_46812# a_10809_44734# 0.013923f
C45319 a_1176_45822# a_167_45260# 0.091673f
C45320 a_11599_46634# a_16147_45260# 0.065926f
C45321 a_1799_45572# a_1990_45899# 8.94e-19
C45322 a_12861_44030# a_18909_45814# 2.11e-19
C45323 a_3160_47472# a_2437_43646# 0.003877f
C45324 a_5326_44056# VDD 0.001151f
C45325 a_14209_32519# a_22465_38105# 6.41e-20
C45326 a_13113_42826# a_13070_42354# 4.26e-19
C45327 a_12545_42858# a_13575_42558# 0.001596f
C45328 a_20193_45348# a_11341_43940# 0.21261f
C45329 a_20202_43084# a_20712_42282# 0.028679f
C45330 a_5147_45002# a_6031_43396# 0.003581f
C45331 a_12549_44172# DATA[5] 3.42e-20
C45332 a_n863_45724# a_4649_42852# 8.36e-21
C45333 a_n1925_42282# a_564_42282# 2.11e-19
C45334 a_8199_44636# a_5742_30871# 5.25e-20
C45335 a_8953_45546# a_10723_42308# 2.61e-20
C45336 a_4185_45028# a_15486_42560# 6.43e-20
C45337 a_626_44172# a_n97_42460# 0.005505f
C45338 a_16131_47204# VDD 0.142103f
C45339 a_9313_44734# a_22959_44484# 1.37e-19
C45340 a_3537_45260# a_6765_43638# 0.025724f
C45341 a_10193_42453# a_10083_42826# 0.002709f
C45342 a_2711_45572# a_19987_42826# 0.003709f
C45343 a_n357_42282# a_7573_43172# 9.51e-19
C45344 a_11309_47204# CLK 0.01087f
C45345 a_7499_43078# a_10991_42826# 0.004793f
C45346 a_526_44458# a_n1630_35242# 9.42e-21
C45347 a_526_44458# a_n2661_45546# 0.071855f
C45348 a_n1925_42282# a_n2810_45572# 3.89e-20
C45349 a_3483_46348# a_10193_42453# 0.359034f
C45350 a_12861_44030# a_12607_44458# 0.020604f
C45351 a_13607_46688# a_2437_43646# 1.22e-21
C45352 SMPL_ON_N a_18114_32519# 0.02927f
C45353 a_n2497_47436# a_n2661_42834# 0.099608f
C45354 a_2063_45854# a_6109_44484# 1.19e-20
C45355 a_19692_46634# a_20273_45572# 0.004885f
C45356 a_19466_46812# a_20841_45814# 1.64e-19
C45357 a_13925_46122# a_2711_45572# 5.04e-19
C45358 a_5257_43370# a_4927_45028# 0.003815f
C45359 a_4791_45118# a_n356_44636# 0.001203f
C45360 a_10554_47026# a_413_45260# 1.94e-20
C45361 a_15227_44166# a_21363_45546# 6.55e-20
C45362 a_n784_42308# a_n3420_38528# 0.005039f
C45363 a_n3674_38216# a_n4251_38528# 5.77e-20
C45364 a_n1630_35242# a_n4209_38502# 3.02e-19
C45365 a_5932_42308# a_n3565_39590# 4.83e-21
C45366 a_n4318_38216# a_n4209_38216# 0.135236f
C45367 a_5342_30871# C2_P_btm 7.86e-20
C45368 a_n3674_37592# a_n3565_38502# 9.8e-20
C45369 a_15051_42282# a_4958_30871# 0.003379f
C45370 a_14113_42308# a_17303_42282# 1.39e-19
C45371 a_15803_42450# a_15761_42308# 2.56e-19
C45372 a_5534_30871# C0_P_btm 8.49e-20
C45373 a_10083_42826# VDD 0.461256f
C45374 a_19963_31679# a_14097_32519# 0.051059f
C45375 a_5013_44260# a_5745_43940# 0.007387f
C45376 a_5495_43940# a_5326_44056# 4.96e-19
C45377 a_n1059_45260# a_16877_42852# 0.058551f
C45378 a_n2017_45002# a_17665_42852# 0.004242f
C45379 a_3483_46348# VDD 2.29096f
C45380 a_19237_31679# a_14401_32519# 0.055111f
C45381 a_17973_43940# a_18079_43940# 0.419086f
C45382 a_17737_43940# a_18326_43940# 4.1e-19
C45383 a_16979_44734# a_17499_43370# 6.72e-19
C45384 a_14539_43914# a_17324_43396# 0.008599f
C45385 a_19721_31679# a_14209_32519# 0.051313f
C45386 a_742_44458# a_743_42282# 6.63e-20
C45387 a_17730_32519# a_17538_32519# 9.37324f
C45388 a_11962_45724# a_11823_42460# 0.177935f
C45389 a_526_44458# a_5205_44484# 2.73e-20
C45390 a_2711_45572# a_15599_45572# 0.045207f
C45391 a_8270_45546# a_9313_44734# 7.8e-20
C45392 a_11415_45002# a_16237_45028# 1.72e-19
C45393 a_18597_46090# a_21115_43940# 0.015966f
C45394 a_3483_46348# a_14309_45348# 2.79e-20
C45395 a_n2293_46634# a_n984_44318# 2.17e-21
C45396 a_18479_47436# a_22223_43948# 1.31e-20
C45397 a_8162_45546# a_8336_45822# 9.93e-20
C45398 a_8199_44636# a_n2293_42834# 0.048304f
C45399 a_5937_45572# a_7639_45394# 2.11e-19
C45400 a_n2438_43548# a_n2065_43946# 0.265458f
C45401 a_12741_44636# a_19113_45348# 0.003982f
C45402 a_16375_45002# a_2437_43646# 2.49e-20
C45403 a_n2497_47436# a_n1352_43396# 0.061218f
C45404 a_11453_44696# a_15682_43940# 1.72e-19
C45405 a_15673_47210# a_n881_46662# 7.77e-20
C45406 a_n4209_39590# a_n1386_35608# 1.02e-19
C45407 a_3160_47472# a_n2661_46634# 0.026361f
C45408 a_21811_47423# a_11453_44696# 0.005338f
C45409 a_4883_46098# a_22959_47212# 8.05e-21
C45410 a_6545_47178# a_5807_45002# 0.030195f
C45411 a_n1435_47204# a_12891_46348# 0.001028f
C45412 a_13381_47204# a_12549_44172# 0.135267f
C45413 a_4958_30871# C9_N_btm 0.209166f
C45414 a_7174_31319# C4_P_btm 2.64e-20
C45415 a_327_47204# a_n133_46660# 0.006131f
C45416 a_1209_47178# a_n2438_43548# 4.34e-19
C45417 a_1239_47204# a_n743_46660# 8.16e-20
C45418 a_22223_47212# a_22731_47423# 0.011229f
C45419 a_12465_44636# SMPL_ON_N 0.006167f
C45420 a_n746_45260# a_383_46660# 0.011439f
C45421 a_n23_47502# a_33_46660# 0.001405f
C45422 a_n785_47204# a_171_46873# 1.04e-19
C45423 a_n971_45724# a_1123_46634# 1.3e-19
C45424 a_15521_42308# RST_Z 4.66e-20
C45425 a_9313_44734# a_18861_43218# 2.63e-19
C45426 a_14495_45572# VDD 0.238674f
C45427 a_15493_43940# a_21259_43561# 8.06e-20
C45428 a_14021_43940# a_16867_43762# 0.004651f
C45429 a_11341_43940# a_20301_43646# 0.001136f
C45430 a_20512_43084# a_20922_43172# 0.001051f
C45431 a_n2956_37592# a_n2216_37984# 1.2e-19
C45432 a_2896_43646# a_2982_43646# 0.100706f
C45433 a_n97_42460# a_2813_43396# 0.001563f
C45434 a_10490_45724# CLK 0.029352f
C45435 a_19862_44208# a_4361_42308# 0.006467f
C45436 a_5257_43370# a_4699_43561# 2.14e-19
C45437 a_13249_42308# a_14403_45348# 8.12e-19
C45438 a_20447_31679# en_comp 2.2e-19
C45439 a_n2293_45010# a_n2017_45002# 0.076023f
C45440 a_n2661_45010# a_n913_45002# 0.019536f
C45441 a_n2472_45002# a_n1059_45260# 7.79e-20
C45442 a_n2497_47436# a_n2293_42282# 1.08e-20
C45443 a_3090_45724# a_10651_43940# 0.014051f
C45444 a_11823_42460# a_13807_45067# 1.27e-21
C45445 a_3483_46348# a_5495_43940# 3.25e-20
C45446 a_n357_42282# a_8975_43940# 1.39e-20
C45447 SMPL_ON_N a_13887_32519# 0.029238f
C45448 a_6755_46942# a_n97_42460# 2.11e-19
C45449 a_1609_45822# a_949_44458# 0.005374f
C45450 a_n443_42852# a_2779_44458# 1.63e-20
C45451 a_13059_46348# a_12603_44260# 3.73e-20
C45452 a_n2293_46634# a_9885_43646# 0.005638f
C45453 a_12549_44172# a_18783_43370# 2.61e-20
C45454 a_13661_43548# a_13837_43396# 1.48e-20
C45455 a_2437_43646# a_413_45260# 0.20387f
C45456 a_18597_46090# a_11415_45002# 0.061694f
C45457 a_3877_44458# a_5257_43370# 0.142219f
C45458 a_13747_46662# a_19333_46634# 0.011849f
C45459 a_12549_44172# a_13170_46660# 2.28e-19
C45460 a_5732_46660# a_6540_46812# 2.56e-19
C45461 a_5167_46660# a_5275_47026# 0.057222f
C45462 VDD VIN_N 1.46155f
C45463 a_n443_46116# a_5164_46348# 1.86e-20
C45464 a_2063_45854# a_9569_46155# 5.78e-20
C45465 a_n1151_42308# a_8349_46414# 0.095055f
C45466 a_4915_47217# a_5068_46348# 6.9e-20
C45467 a_4791_45118# a_5204_45822# 0.053732f
C45468 a_13661_43548# a_19466_46812# 0.011727f
C45469 a_5807_45002# a_19692_46634# 6.61e-19
C45470 C10_N_btm VREF_GND 10.3207f
C45471 C9_N_btm VCM 6.06251f
C45472 a_13507_46334# a_19636_46660# 4.68e-19
C45473 a_11453_44696# a_22000_46634# 0.008499f
C45474 a_17730_32519# a_22465_38105# 2.17e-19
C45475 a_22223_43396# a_17364_32525# 2.46e-19
C45476 a_n97_42460# a_16328_43172# 7.85e-19
C45477 a_22591_43396# a_14209_32519# 0.158752f
C45478 a_17719_45144# VDD 0.1297f
C45479 a_10341_43396# a_15279_43071# 0.001151f
C45480 a_18175_45572# a_11967_42832# 4.42e-21
C45481 a_18341_45572# a_18588_44850# 5.56e-21
C45482 a_3090_45724# a_12895_43230# 0.004563f
C45483 a_10903_43370# a_9803_43646# 2.58e-19
C45484 a_2711_45572# a_18326_43940# 0.009029f
C45485 a_327_44734# a_700_44734# 0.003235f
C45486 a_n2661_45010# a_556_44484# 0.038106f
C45487 a_9290_44172# a_14358_43442# 0.001132f
C45488 SMPL_ON_P a_n2302_40160# 1.79e-19
C45489 a_8953_45546# a_10341_43396# 0.001386f
C45490 a_n1925_42282# a_n1557_42282# 0.013245f
C45491 a_526_44458# a_1427_43646# 0.028942f
C45492 a_1307_43914# a_n699_43396# 0.094953f
C45493 en_comp a_5891_43370# 2.34e-21
C45494 a_n2312_40392# a_6123_31319# 7.4e-21
C45495 a_n2017_45002# a_9313_44734# 0.009039f
C45496 a_3357_43084# a_n2661_43922# 0.031253f
C45497 a_11963_45334# a_8975_43940# 4.93e-19
C45498 a_9482_43914# a_10157_44484# 0.321004f
C45499 a_626_44172# a_742_44458# 0.022141f
C45500 a_n863_45724# a_1241_43940# 6.18e-19
C45501 a_n2956_39768# a_n2840_42282# 3.63e-20
C45502 a_3483_46348# a_16137_43396# 6.08e-20
C45503 a_20107_46660# a_22365_46825# 4.87e-21
C45504 a_20841_46902# a_21350_47026# 2.6e-19
C45505 a_20273_46660# a_20719_46660# 2.28e-19
C45506 a_4883_46098# a_6194_45824# 9.26e-21
C45507 a_19594_46812# a_19443_46116# 1.96e-19
C45508 a_768_44030# a_n863_45724# 0.020071f
C45509 a_11459_47204# a_11652_45724# 7.77e-21
C45510 a_n2293_46634# a_13259_45724# 0.032341f
C45511 a_4791_45118# a_8697_45822# 1.06e-20
C45512 a_6151_47436# a_6229_45572# 0.002879f
C45513 a_n1151_42308# a_8120_45572# 5.11e-19
C45514 a_11186_47026# a_11189_46129# 3.64e-19
C45515 a_n881_46662# a_3316_45546# 6.79e-20
C45516 a_19123_46287# a_11415_45002# 5.55e-20
C45517 a_n743_46660# a_12839_46116# 0.011568f
C45518 a_8667_46634# a_6945_45028# 5.95e-20
C45519 a_4955_46873# a_3873_46454# 1.98e-20
C45520 a_5649_42852# a_8685_42308# 5.5e-20
C45521 a_4361_42308# a_9803_42558# 0.011987f
C45522 a_18083_42858# a_20256_43172# 9.94e-21
C45523 a_18599_43230# a_18861_43218# 0.001705f
C45524 a_18817_42826# a_19273_43230# 4.2e-19
C45525 a_10341_43396# a_13258_32519# 2.74e-20
C45526 a_3080_42308# a_n3420_38528# 1.75e-20
C45527 a_10083_42826# a_n784_42308# 8.21e-21
C45528 a_3935_42891# a_1755_42282# 3.67e-22
C45529 a_743_42282# a_10533_42308# 0.016446f
C45530 a_261_44278# VDD 2.43e-19
C45531 a_n913_45002# a_21381_43940# 5.97e-20
C45532 a_n357_42282# a_2905_42968# 0.011153f
C45533 SMPL_ON_N EN_VIN_BSTR_N 1.61e-19
C45534 a_n2293_42834# a_8018_44260# 0.001899f
C45535 a_n443_42852# a_n13_43084# 0.13203f
C45536 a_526_44458# a_3863_42891# 8.86e-21
C45537 a_9067_47204# DATA[4] 0.354356f
C45538 a_9482_43914# a_12710_44260# 0.001272f
C45539 a_13059_46348# a_13657_42558# 3.57e-21
C45540 a_15227_44166# a_17303_42282# 1.37e-19
C45541 a_5111_44636# a_5829_43940# 1.13e-20
C45542 a_6109_44484# a_n2661_42834# 0.026239f
C45543 a_13487_47204# VDD 0.273369f
C45544 a_18114_32519# a_22959_44484# 0.016108f
C45545 a_19721_31679# a_17730_32519# 0.051334f
C45546 a_13717_47436# START 0.034426f
C45547 a_3537_45260# a_8487_44056# 2.95e-19
C45548 a_17970_44736# a_17061_44734# 1.93e-19
C45549 a_17767_44458# a_17517_44484# 0.055175f
C45550 a_1138_42852# a_961_42354# 2.56e-20
C45551 a_13259_45724# a_5342_30871# 2.89e-19
C45552 a_12861_44030# RST_Z 0.290405f
C45553 a_17957_46116# a_8049_45260# 4.87e-20
C45554 a_11387_46155# a_11315_46155# 6.64e-19
C45555 a_n2293_46098# a_3503_45724# 0.01404f
C45556 a_n901_46420# a_n755_45592# 0.002034f
C45557 a_1823_45246# a_n2293_45546# 0.234971f
C45558 a_4185_45028# a_20205_31679# 8.52e-20
C45559 a_n2293_46634# a_n467_45028# 0.008099f
C45560 a_n2661_46634# a_413_45260# 0.029743f
C45561 a_n2497_47436# a_n1352_44484# 0.006874f
C45562 a_472_46348# a_n1099_45572# 0.005608f
C45563 a_805_46414# a_380_45546# 5.77e-19
C45564 a_376_46348# a_310_45028# 5.66e-19
C45565 a_768_44030# a_8191_45002# 1.08e-20
C45566 a_n2438_43548# a_n2810_45028# 0.009971f
C45567 a_5807_45002# a_4927_45028# 6.39e-19
C45568 a_6755_46942# a_16020_45572# 0.010518f
C45569 a_2609_46660# a_2437_43646# 9.86e-20
C45570 a_1176_45822# a_n863_45724# 2.47e-19
C45571 a_11189_46129# a_12839_46116# 8.15e-20
C45572 a_13351_46090# a_12379_46436# 2.98e-20
C45573 a_12594_46348# a_12638_46436# 0.049443f
C45574 a_5934_30871# a_8325_42308# 0.173576f
C45575 a_8515_42308# a_8337_42558# 6.01e-20
C45576 a_4921_42308# a_5742_30871# 3.53e-20
C45577 a_7963_42308# a_8685_42308# 2.62e-19
C45578 a_4190_30871# C0_P_btm 6.53e-20
C45579 a_17364_32525# a_11530_34132# 0.007158f
C45580 a_16664_43396# VDD 0.077608f
C45581 a_5343_44458# a_8147_43396# 0.014327f
C45582 a_742_44458# a_2813_43396# 1.77e-19
C45583 a_16922_45042# a_16409_43396# 4.18e-21
C45584 a_n913_45002# a_18249_42858# 4.01e-20
C45585 a_n2017_45002# a_18599_43230# 0.029677f
C45586 a_n1059_45260# a_18817_42826# 1.2e-20
C45587 a_20193_45348# a_10341_43396# 0.086741f
C45588 a_13259_45724# a_20107_42308# 1.03e-19
C45589 a_2998_44172# a_2537_44260# 3.26e-21
C45590 a_5883_43914# a_6197_43396# 0.001031f
C45591 a_3357_43084# a_3445_43172# 5.23e-19
C45592 a_n356_44636# a_1209_43370# 0.025313f
C45593 a_14513_46634# VDD 0.223375f
C45594 a_6298_44484# a_7287_43370# 0.003354f
C45595 a_20980_44850# a_20935_43940# 1.59e-19
C45596 a_n2956_38680# a_n4064_38528# 0.058755f
C45597 a_n357_42282# a_15803_42450# 1.12e-19
C45598 en_comp a_17595_43084# 2.61e-21
C45599 a_375_42282# a_n13_43084# 0.006217f
C45600 a_14180_46812# RST_Z 5.82e-19
C45601 a_1609_45822# a_1990_45572# 0.002458f
C45602 a_8049_45260# a_16020_45572# 0.002165f
C45603 a_3483_46348# a_5691_45260# 0.005653f
C45604 a_9290_44172# en_comp 1.1e-20
C45605 a_15227_44166# a_19778_44110# 6.82e-20
C45606 a_3090_45724# a_11827_44484# 0.066595f
C45607 a_2711_45572# a_5263_45724# 0.013854f
C45608 a_n357_42282# a_10193_42453# 0.634772f
C45609 a_n2293_46634# a_n2661_43922# 0.023539f
C45610 a_n2442_46660# a_n2293_43922# 7.85e-20
C45611 a_18189_46348# a_3357_43084# 4.56e-21
C45612 a_2063_45854# a_10405_44172# 0.001338f
C45613 a_n443_46116# a_3499_42826# 4.85e-21
C45614 a_4704_46090# a_4558_45348# 6.71e-22
C45615 a_18985_46122# a_2437_43646# 4.38e-21
C45616 a_19466_46812# a_18587_45118# 7.19e-20
C45617 a_10903_43370# a_n913_45002# 0.021559f
C45618 a_4185_45028# a_5111_44636# 3.83e-19
C45619 a_8199_44636# a_413_45260# 4.56e-21
C45620 a_5164_46348# a_3537_45260# 0.003403f
C45621 a_12741_44636# a_16751_45260# 0.01378f
C45622 a_15803_42450# CAL_N 0.002185f
C45623 a_1343_38525# a_1177_38525# 0.238422f
C45624 a_5932_42308# C4_P_btm 0.032349f
C45625 a_n784_42308# VIN_N 0.004358f
C45626 a_n3690_39392# a_n4064_38528# 6.81e-20
C45627 a_n3420_39072# a_n2946_38778# 2.59e-20
C45628 a_n3565_39304# a_n2302_38778# 8.25e-19
C45629 a_n4064_39072# a_n3690_38528# 6.81e-20
C45630 a_n2946_39072# a_n3420_38528# 2.59e-20
C45631 a_n4064_39616# a_n3420_37984# 0.050009f
C45632 a_n3420_39616# a_n4064_37984# 0.046151f
C45633 a_4958_30871# a_n3420_37440# 0.033151f
C45634 a_6123_31319# C9_P_btm 9.33e-20
C45635 a_2351_42308# VDD 0.188239f
C45636 a_n1151_42308# a_10227_46804# 0.458569f
C45637 a_7903_47542# a_n1435_47204# 2.39e-19
C45638 a_9863_47436# a_9313_45822# 0.049145f
C45639 a_n1741_47186# a_n2312_39304# 0.005742f
C45640 SMPL_ON_P a_n2312_40392# 4.89949f
C45641 a_n2109_47186# a_n89_47570# 2.32e-19
C45642 a_6151_47436# a_14955_47212# 0.192081f
C45643 a_20205_31679# VREF_GND 0.001993f
C45644 a_17730_32519# a_22591_43396# 7.33e-19
C45645 a_n2293_42834# a_4921_42308# 2.38e-19
C45646 en_comp a_21887_42336# 2.22e-20
C45647 a_n357_42282# VDD 1.90108f
C45648 a_9313_44734# a_19164_43230# 0.004691f
C45649 a_20692_30879# VREF 0.098117f
C45650 a_20512_43084# a_17364_32525# 1.45e-20
C45651 a_10193_42453# CAL_N 0.00219f
C45652 a_12861_44030# a_16243_43396# 9.34e-20
C45653 a_3775_45552# a_1423_45028# 4.78e-21
C45654 a_2711_45572# a_5837_45348# 3.63e-19
C45655 a_2324_44458# a_5891_43370# 7.07e-20
C45656 a_7499_43078# a_9482_43914# 0.062333f
C45657 a_768_44030# a_3540_43646# 0.002561f
C45658 a_n1613_43370# a_6765_43638# 0.164755f
C45659 a_4883_46098# a_9803_43646# 0.002651f
C45660 a_n881_46662# a_6197_43396# 6.52e-20
C45661 a_n2438_43548# a_n2129_43609# 0.068602f
C45662 a_3218_45724# a_n2661_43370# 6.79e-20
C45663 a_3483_46348# a_13940_44484# 1.24e-19
C45664 a_18175_45572# a_20273_45572# 3.92e-21
C45665 a_18479_45785# a_20107_45572# 3.61e-20
C45666 a_18909_45814# a_18787_45572# 3.16e-19
C45667 a_13904_45546# a_6171_45002# 3.3e-20
C45668 a_11322_45546# a_10775_45002# 6.82e-20
C45669 a_10193_42453# a_11963_45334# 0.007668f
C45670 a_10490_45724# a_10951_45334# 1.32e-19
C45671 SMPL_ON_P a_n2840_42826# 7.81e-19
C45672 a_n3420_37440# VCM 0.033198f
C45673 a_16241_47178# a_16292_46812# 3.13e-19
C45674 a_16327_47482# a_15559_46634# 0.001169f
C45675 a_n743_46660# a_491_47026# 6.49e-20
C45676 a_n2438_43548# a_288_46660# 0.013776f
C45677 CAL_N VDD 26.069302f
C45678 EN_VIN_BSTR_N a_19864_35138# 0.573134f
C45679 a_11206_38545# RST_Z 0.382319f
C45680 a_n133_46660# a_1983_46706# 6.11e-21
C45681 a_n1021_46688# a_n935_46688# 0.006584f
C45682 a_n2661_46634# a_2609_46660# 0.045654f
C45683 a_5807_45002# a_3877_44458# 0.034811f
C45684 a_n881_46662# a_8145_46902# 0.003327f
C45685 a_4915_47217# a_13059_46348# 0.021189f
C45686 a_18194_35068# a_19120_35138# 0.558402f
C45687 EN_VIN_BSTR_P C9_P_btm 0.226529f
C45688 a_3160_47472# a_765_45546# 0.027219f
C45689 a_n4064_37440# VREF 1.56e-19
C45690 a_n2293_46634# a_1799_45572# 0.001265f
C45691 a_n2442_46660# a_n2661_46098# 6.94e-20
C45692 a_33_46660# a_948_46660# 0.117156f
C45693 a_11599_46634# a_19333_46634# 0.001374f
C45694 a_10227_46804# a_14084_46812# 1.42e-19
C45695 a_14579_43548# a_4361_42308# 2.32e-19
C45696 a_15681_43442# a_15868_43402# 1.84e-19
C45697 a_21381_43940# a_20922_43172# 0.00196f
C45698 a_16137_43396# a_16664_43396# 0.002125f
C45699 a_11963_45334# VDD 0.229584f
C45700 a_10341_43396# a_20301_43646# 0.002799f
C45701 a_2998_44172# a_2903_42308# 4.71e-20
C45702 a_17499_43370# a_18429_43548# 0.012474f
C45703 a_16409_43396# a_15743_43084# 0.586918f
C45704 a_n2661_42282# a_n4318_38216# 0.023731f
C45705 a_11967_42832# a_15486_42560# 1.23e-19
C45706 a_6171_45002# CLK 0.032376f
C45707 a_n97_42460# a_15279_43071# 0.001255f
C45708 a_3626_43646# a_5111_42852# 3.39e-20
C45709 a_3539_42460# a_4520_42826# 0.003363f
C45710 a_13159_45002# a_13490_45394# 2.88e-19
C45711 a_13017_45260# a_13711_45394# 2.64e-19
C45712 a_13249_42308# a_14581_44484# 1.15e-19
C45713 a_3483_46348# a_3080_42308# 2.72e-21
C45714 a_n443_42852# a_644_44056# 1.15e-19
C45715 a_n2661_45010# a_n2661_44458# 0.090852f
C45716 a_1823_45246# a_2896_43646# 6.58e-19
C45717 a_8696_44636# a_7640_43914# 9.09e-20
C45718 a_6171_45002# a_17023_45118# 7.32e-19
C45719 a_18479_47436# a_20753_42852# 2.93e-20
C45720 a_18175_45572# a_18989_43940# 6.34e-20
C45721 a_18691_45572# a_18248_44752# 2.36e-21
C45722 a_18341_45572# a_18443_44721# 3.12e-21
C45723 a_18479_45785# a_18374_44850# 3.69e-20
C45724 a_18909_45814# a_18287_44626# 8.28e-19
C45725 a_n357_42282# a_5495_43940# 1.86e-21
C45726 a_3218_45724# a_2998_44172# 1.18e-19
C45727 a_8953_45546# a_n97_42460# 0.015611f
C45728 a_13059_46348# a_15681_43442# 2.56e-21
C45729 a_4791_45118# a_3823_42558# 0.005746f
C45730 a_18597_46090# a_13259_45724# 1.02e-19
C45731 a_16327_47482# a_20009_46494# 2.95e-19
C45732 a_n2497_47436# a_3775_45552# 4.13e-21
C45733 a_n1741_47186# a_6511_45714# 4.36e-21
C45734 a_n971_45724# a_4099_45572# 8.72e-19
C45735 a_n443_46116# a_3316_45546# 3.74e-19
C45736 a_n1151_42308# a_n906_45572# 0.002303f
C45737 a_6755_46942# a_11415_45002# 0.02226f
C45738 a_n881_46662# a_5066_45546# 0.801045f
C45739 a_13607_46688# a_765_45546# 2.05e-20
C45740 a_15009_46634# a_15312_46660# 0.001377f
C45741 a_4883_46098# a_14371_46494# 2.3e-19
C45742 a_20916_46384# a_20708_46348# 0.189941f
C45743 a_19321_45002# a_10809_44734# 0.035502f
C45744 a_20843_47204# a_6945_45028# 0.003967f
C45745 a_n237_47217# a_2711_45572# 0.025745f
C45746 a_3877_44458# a_3699_46348# 0.084544f
C45747 a_4646_46812# a_3483_46348# 0.048267f
C45748 a_17609_46634# a_16388_46812# 2.5e-19
C45749 a_11599_46634# a_20062_46116# 6.27e-19
C45750 a_2107_46812# a_10903_43370# 9.6e-21
C45751 a_n743_46660# a_14840_46494# 0.010488f
C45752 a_743_42282# a_20256_42852# 1.03e-20
C45753 a_8685_43396# a_8685_42308# 9.74e-19
C45754 a_9145_43396# a_5934_30871# 3.25e-19
C45755 a_17538_32519# a_22465_38105# 2e-19
C45756 a_3422_30871# C5_P_btm 1.71e-19
C45757 a_18599_43230# a_19164_43230# 7.99e-20
C45758 a_3626_43646# a_9885_42308# 0.001057f
C45759 a_8387_43230# a_8483_43230# 0.013793f
C45760 a_18588_44850# VDD 0.132317f
C45761 a_17730_32519# a_18194_35068# 1.21e-19
C45762 a_n1925_42282# a_3935_42891# 0.010366f
C45763 a_526_44458# a_4520_42826# 0.247914f
C45764 a_11827_44484# a_14815_43914# 0.029578f
C45765 a_n357_42282# a_16137_43396# 1.09442f
C45766 a_16112_44458# a_14539_43914# 0.13299f
C45767 a_7499_43078# a_6031_43396# 7.11e-20
C45768 a_626_44172# a_n984_44318# 7.42e-19
C45769 a_3537_45260# a_3499_42826# 0.001528f
C45770 a_n1059_45260# a_15682_43940# 0.001131f
C45771 a_n2017_45002# a_17737_43940# 1.87e-21
C45772 a_13259_45724# a_743_42282# 0.066992f
C45773 a_2382_45260# a_n2661_42282# 2.02e-19
C45774 a_8191_45002# a_7845_44172# 4.75e-20
C45775 a_11691_44458# a_13213_44734# 0.046347f
C45776 a_1307_43914# a_1467_44172# 0.228571f
C45777 a_n2661_44458# a_8855_44734# 3.59e-19
C45778 a_n2442_46660# a_n3420_39616# 0.00978f
C45779 a_n2956_39768# a_n2302_39866# 0.037924f
C45780 a_n443_42852# a_10765_43646# 6.06e-19
C45781 a_4883_46098# a_n913_45002# 1.34e-19
C45782 a_10903_43370# a_14493_46090# 1.62e-20
C45783 a_584_46384# a_1423_45028# 1.63e-19
C45784 a_1138_42852# a_1337_46436# 1.4e-19
C45785 a_4915_47217# a_13556_45296# 0.146395f
C45786 a_18143_47464# a_413_45260# 4.35e-19
C45787 a_11415_45002# a_8049_45260# 0.426371f
C45788 a_5807_45002# a_18175_45572# 0.004334f
C45789 a_13661_43548# a_16147_45260# 0.002524f
C45790 a_13747_46662# a_17786_45822# 0.005559f
C45791 a_12861_44030# a_3232_43370# 2.11e-21
C45792 a_3094_47570# a_2437_43646# 9.06e-19
C45793 a_18285_46348# a_18147_46436# 0.001014f
C45794 a_765_45546# a_16375_45002# 0.008153f
C45795 a_19123_46287# a_13259_45724# 6.59e-21
C45796 a_n1151_42308# a_1307_43914# 3.38e-20
C45797 a_7577_46660# a_8568_45546# 1.67e-20
C45798 a_8270_45546# a_2711_45572# 0.063301f
C45799 a_n743_46660# a_16115_45572# 0.012735f
C45800 a_9290_44172# a_2324_44458# 0.026216f
C45801 a_12594_46348# a_13759_46122# 9.6e-19
C45802 a_21671_42860# a_21613_42308# 9.03e-20
C45803 a_22165_42308# a_21887_42336# 0.110763f
C45804 a_3080_42308# VIN_N 0.025929f
C45805 a_16137_43396# CAL_N 7.09e-19
C45806 a_n144_43396# VDD 3.23e-19
C45807 a_14097_32519# a_5932_42308# 0.001859f
C45808 a_n1630_35242# a_1221_42558# 2.09e-20
C45809 a_n473_42460# a_n39_42308# 0.003935f
C45810 a_1067_42314# a_1149_42558# 0.004937f
C45811 a_n784_42308# a_2351_42308# 0.0035f
C45812 a_18374_44850# a_14021_43940# 6.68e-21
C45813 a_9313_44734# a_18079_43940# 1.98e-20
C45814 a_22591_44484# a_17730_32519# 0.156987f
C45815 a_20512_43084# a_19237_31679# 1.14e-20
C45816 a_n2661_42834# a_10405_44172# 0.005797f
C45817 a_n2661_43922# a_9672_43914# 8.49e-20
C45818 a_19721_31679# a_17538_32519# 0.051191f
C45819 a_5883_43914# a_8415_44056# 6.67e-19
C45820 a_n863_45724# a_1067_42314# 0.289393f
C45821 a_n755_45592# a_196_42282# 0.090568f
C45822 a_n357_42282# a_n784_42308# 0.008228f
C45823 a_n913_45002# a_5649_42852# 0.0586f
C45824 en_comp a_13467_32519# 1.89e-19
C45825 a_n2438_43548# a_n2129_44697# 0.060059f
C45826 a_7577_46660# a_n2661_43370# 3.63e-21
C45827 a_3090_45724# a_15595_45028# 0.00235f
C45828 a_15227_44166# a_9482_43914# 0.020073f
C45829 a_14976_45028# a_15415_45028# 0.027906f
C45830 a_n2497_47436# a_n1549_44318# 0.018493f
C45831 SMPL_ON_P a_n2472_43914# 3.53e-19
C45832 a_5066_45546# a_8162_45546# 0.025437f
C45833 a_n2840_45546# a_n1099_45572# 3.93e-20
C45834 a_12549_44172# a_17767_44458# 1.63e-20
C45835 a_14035_46660# a_6171_45002# 3.2e-20
C45836 a_n1613_43370# a_n1655_44484# 0.003155f
C45837 a_10227_46804# a_13857_44734# 4.26e-19
C45838 a_20820_30879# a_2437_43646# 0.006482f
C45839 a_12741_44636# a_21513_45002# 1.26e-19
C45840 a_20202_43084# a_3357_43084# 0.029548f
C45841 a_11415_45002# a_19479_31679# 0.224531f
C45842 a_765_45546# a_413_45260# 0.031429f
C45843 a_n2293_46634# a_n452_44636# 3.66e-20
C45844 a_n2472_45546# a_n863_45724# 1.45e-19
C45845 a_n2956_38216# a_n1079_45724# 5.55e-20
C45846 a_13925_46122# a_14033_45822# 0.001241f
C45847 a_n2661_45546# a_n452_45724# 0.007419f
C45848 a_n971_45724# a_n746_45260# 0.393354f
C45849 a_n1605_47204# a_n785_47204# 2e-19
C45850 a_n452_47436# a_n237_47217# 0.061523f
C45851 a_n1741_47186# a_1209_47178# 0.046323f
C45852 a_n2109_47186# a_1431_47204# 0.050586f
C45853 a_n2497_47436# a_584_46384# 0.06459f
C45854 a_n815_47178# a_n23_47502# 9.5e-20
C45855 a_n1630_35242# VDAC_N 0.003372f
C45856 COMP_P a_22459_39145# 0.032214f
C45857 a_n784_42308# CAL_N 0.00432f
C45858 a_20205_31679# a_22469_40625# 1.74e-20
C45859 a_20692_30879# a_22521_40599# 2.53e-20
C45860 a_19478_44306# a_19478_44056# 0.001278f
C45861 a_2382_45260# a_3497_42558# 0.001486f
C45862 a_n913_45002# a_7963_42308# 0.044607f
C45863 a_20269_44172# a_19319_43548# 0.12985f
C45864 a_9895_44260# a_9801_43940# 1.26e-19
C45865 a_11341_43940# a_13565_43940# 0.00518f
C45866 a_518_46155# VDD 0.00166f
C45867 a_9313_44734# a_14209_32519# 0.068114f
C45868 a_10440_44484# a_10518_42984# 1.11e-21
C45869 a_8975_43940# a_8952_43230# 2.23e-20
C45870 a_10057_43914# a_10083_42826# 0.001039f
C45871 a_19328_44172# a_19741_43940# 0.04732f
C45872 a_n2017_45002# a_8515_42308# 0.002597f
C45873 a_n1059_45260# a_5934_30871# 0.010576f
C45874 a_21137_46414# a_21005_45260# 1.84e-20
C45875 a_10903_43370# a_n2661_44458# 4.92e-19
C45876 a_3316_45546# a_3537_45260# 0.078381f
C45877 a_3483_46348# a_10057_43914# 0.00873f
C45878 a_n443_42852# a_n37_45144# 0.137227f
C45879 a_509_45822# a_413_45260# 1.95e-19
C45880 SMPL_ON_N a_14401_32519# 0.029323f
C45881 a_3503_45724# a_3429_45260# 2.71e-19
C45882 a_5257_43370# a_5244_44056# 6.32e-19
C45883 a_2711_45572# a_n2017_45002# 0.02728f
C45884 a_19466_46812# a_11967_42832# 8.14e-20
C45885 a_2211_45572# a_2437_43646# 5.1e-19
C45886 a_n1613_43370# a_8487_44056# 3.38e-21
C45887 a_16375_45002# a_16751_45260# 0.047561f
C45888 a_18819_46122# a_11691_44458# 2.75e-19
C45889 a_18985_46122# a_19113_45348# 6.36e-21
C45890 a_768_44030# a_2455_43940# 0.005192f
C45891 a_13661_43548# a_13565_44260# 3.81e-19
C45892 a_n4064_39072# VIN_P 0.039352f
C45893 a_15928_47570# a_16119_47582# 4.61e-19
C45894 a_12891_46348# a_13759_47204# 1.25e-20
C45895 a_768_44030# a_13569_47204# 8.63e-20
C45896 a_12549_44172# a_13675_47204# 5.51e-19
C45897 a_n1435_47204# a_4817_46660# 1.96e-20
C45898 a_6151_47436# a_5257_43370# 0.009542f
C45899 a_8128_46384# a_5807_45002# 0.023925f
C45900 a_n2312_40392# a_n2438_43548# 6.39e-22
C45901 a_n3690_38528# VDD 0.363159f
C45902 a_3726_37500# a_6886_37412# 0.702909f
C45903 a_4338_37500# a_5700_37509# 2.69237f
C45904 a_n3565_39304# VCM 0.035438f
C45905 a_4883_46098# a_2107_46812# 2.95673f
C45906 a_4915_47217# a_7577_46660# 1.88e-19
C45907 a_2063_45854# a_6969_46634# 0.00119f
C45908 a_n1151_42308# a_10467_46802# 0.031981f
C45909 a_3626_43646# a_16977_43638# 2.8e-21
C45910 a_2982_43646# a_17499_43370# 4.15e-20
C45911 a_8685_43396# a_9803_43646# 0.008605f
C45912 a_18451_43940# a_18249_42858# 2.07e-20
C45913 a_15493_43396# a_18083_42858# 6.8e-21
C45914 a_19721_31679# a_22465_38105# 3.17e-19
C45915 a_11341_43940# a_5534_30871# 6.54e-20
C45916 a_5891_43370# a_9803_42558# 0.002774f
C45917 a_14401_32519# a_22959_43396# 0.016242f
C45918 a_20974_43370# a_14209_32519# 0.049701f
C45919 a_3422_30871# a_22400_42852# 0.023064f
C45920 a_n356_44636# a_14456_42282# 2.77e-19
C45921 a_n2661_42834# a_6171_42473# 9.02e-22
C45922 a_6171_45002# a_10951_45334# 0.00438f
C45923 a_3232_43370# a_11787_45002# 0.001844f
C45924 a_7229_43940# a_7705_45326# 0.203098f
C45925 a_7276_45260# a_8191_45002# 3.64e-20
C45926 a_8696_44636# a_16981_45144# 0.003008f
C45927 a_15861_45028# a_16886_45144# 8.28e-19
C45928 a_3357_43084# a_5837_45028# 0.006851f
C45929 a_n2438_43548# a_n2840_42826# 2.22e-21
C45930 a_10193_42453# a_18443_44721# 8.46e-19
C45931 a_n37_45144# a_375_42282# 7.33e-19
C45932 a_18175_45572# a_18315_45260# 0.008723f
C45933 a_13507_46334# a_21195_42852# 0.005401f
C45934 a_n2956_39768# a_n3674_39304# 0.023853f
C45935 a_768_44030# a_7765_42852# 1.22e-20
C45936 a_3090_45724# a_8147_43396# 0.002892f
C45937 a_2324_44458# a_10807_43548# 1.65e-20
C45938 a_11823_42460# a_15004_44636# 2.75e-20
C45939 a_3483_46348# a_14021_43940# 0.066924f
C45940 w_1575_34946# a_5934_30871# 0.002787f
C45941 a_n1151_42308# a_8034_45724# 0.040415f
C45942 a_2609_46660# a_765_45546# 0.009946f
C45943 a_6755_46942# a_12251_46660# 0.033714f
C45944 a_9804_47204# a_3483_46348# 6.33e-21
C45945 a_11453_44696# a_10903_43370# 0.040346f
C45946 a_4883_46098# a_14493_46090# 0.00233f
C45947 a_18479_47436# a_18819_46122# 6.05e-20
C45948 a_16327_47482# a_21137_46414# 1.42e-20
C45949 a_16241_47178# a_6945_45028# 0.011279f
C45950 a_n443_46116# a_5066_45546# 0.130975f
C45951 a_4791_45118# a_6419_46482# 9.06e-19
C45952 a_13507_46334# a_15015_46420# 0.005128f
C45953 a_10227_46804# a_19553_46090# 4.1e-21
C45954 a_15811_47375# a_10809_44734# 0.049971f
C45955 a_22612_30879# a_21076_30879# 0.056101f
C45956 a_18597_46090# a_18189_46348# 4.44e-19
C45957 a_12465_44636# a_13759_46122# 0.018063f
C45958 a_n1613_43370# a_5164_46348# 3.39e-19
C45959 a_n881_46662# a_5068_46348# 0.078135f
C45960 a_10341_43396# a_15785_43172# 5.75e-19
C45961 a_20623_43914# a_20712_42282# 1.64e-19
C45962 a_7227_42852# a_7871_42858# 2.32e-20
C45963 a_4361_42308# a_21671_42860# 0.012186f
C45964 a_13467_32519# a_22165_42308# 0.009474f
C45965 a_21115_43940# a_13258_32519# 1.2e-21
C45966 a_5649_42852# a_20922_43172# 8.67e-21
C45967 a_18443_44721# VDD 0.193515f
C45968 a_3080_42308# a_2351_42308# 1.79e-19
C45969 a_n443_42852# a_104_43370# 0.003607f
C45970 a_15415_45028# a_15433_44458# 9.2e-19
C45971 a_n2661_43370# a_n1190_44850# 1.23e-19
C45972 a_15599_45572# a_15682_43940# 4.45e-19
C45973 a_13661_43548# a_15051_42282# 1.21e-20
C45974 a_13249_42308# a_14485_44260# 6.05e-19
C45975 a_n2956_39768# a_5742_30871# 7.02e-21
C45976 a_3090_45724# a_13569_43230# 1.94e-19
C45977 a_8696_44636# a_10729_43914# 7.58e-20
C45978 a_n2661_45546# a_3626_43646# 0.009175f
C45979 a_626_44172# a_n2661_43922# 0.03074f
C45980 a_n357_42282# a_3080_42308# 0.023702f
C45981 a_n755_45592# a_4699_43561# 2.57e-21
C45982 a_n1925_46634# a_6598_45938# 8.63e-21
C45983 a_3877_44458# a_n755_45592# 0.001347f
C45984 a_4646_46812# a_n357_42282# 0.030404f
C45985 a_768_44030# a_11823_42460# 0.066425f
C45986 a_12549_44172# a_12791_45546# 0.083854f
C45987 a_5807_45002# a_10053_45546# 3.59e-20
C45988 a_6755_46942# a_13259_45724# 0.021651f
C45989 a_n2293_46098# a_5164_46348# 2.77e-19
C45990 a_1138_42852# a_1823_45246# 7.31e-20
C45991 a_n746_45260# a_n2293_45010# 0.023201f
C45992 a_2063_45854# a_3357_43084# 0.023045f
C45993 a_4883_46098# a_15903_45785# 1.41e-19
C45994 a_n743_46660# a_6511_45714# 0.003331f
C45995 a_1799_45572# a_2277_45546# 2.46e-19
C45996 a_12891_46348# a_13163_45724# 0.009037f
C45997 a_19123_46287# a_18189_46348# 1.43e-20
C45998 a_18285_46348# a_17957_46116# 0.12677f
C45999 a_8270_45546# a_10037_46155# 4.27e-20
C46000 a_13059_46348# a_10809_44734# 0.003202f
C46001 a_16721_46634# a_6945_45028# 6e-20
C46002 a_11599_46634# a_17786_45822# 2.55e-20
C46003 a_2905_45572# a_2437_43646# 0.003457f
C46004 a_12861_44030# a_18341_45572# 0.026945f
C46005 a_1208_46090# a_167_45260# 0.001892f
C46006 a_5025_43940# VDD 0.004306f
C46007 a_17538_32519# a_18194_35068# 1.07e-19
C46008 a_12545_42858# a_13070_42354# 5.71e-19
C46009 a_9290_44172# a_9803_42558# 0.094028f
C46010 a_11691_44458# a_11341_43940# 4.94e-19
C46011 a_20193_45348# a_21115_43940# 0.01963f
C46012 a_12891_46348# DATA[5] 0.001817f
C46013 a_526_44458# a_564_42282# 1.5e-19
C46014 a_n1925_42282# a_n3674_37592# 0.072052f
C46015 a_8953_45546# a_10533_42308# 7.15e-20
C46016 a_4185_45028# a_15051_42282# 4.66e-19
C46017 a_20202_43084# a_20107_42308# 0.002968f
C46018 a_375_42282# a_104_43370# 0.001385f
C46019 a_n356_44636# a_895_43940# 0.026898f
C46020 a_9313_44734# a_17730_32519# 3.13e-20
C46021 a_2711_45572# a_19164_43230# 0.006484f
C46022 a_3537_45260# a_6197_43396# 0.337459f
C46023 a_7499_43078# a_10796_42968# 0.030705f
C46024 a_n913_45002# a_8685_43396# 0.03156f
C46025 a_3483_46348# a_10180_45724# 0.047643f
C46026 a_12816_46660# a_2437_43646# 1.78e-20
C46027 a_4883_46098# a_n2661_44458# 0.019556f
C46028 a_8049_45260# a_13259_45724# 0.895805f
C46029 a_n1151_42308# a_n998_44484# 7.11e-19
C46030 a_19692_46634# a_20107_45572# 0.001896f
C46031 a_19466_46812# a_20273_45572# 0.328586f
C46032 a_13759_46122# a_2711_45572# 2.27e-19
C46033 a_5257_43370# a_5111_44636# 0.22597f
C46034 a_15227_44166# a_20623_45572# 0.002557f
C46035 a_8952_43230# VDD 0.273404f
C46036 a_5342_30871# C3_P_btm 8.34e-20
C46037 a_n3674_37592# a_n4334_38528# 6.44e-20
C46038 a_5934_30871# a_n4315_30879# 8.24e-21
C46039 a_14113_42308# a_4958_30871# 0.058048f
C46040 a_15764_42576# a_15761_42308# 2.36e-20
C46041 a_5534_30871# C1_P_btm 1.06e-19
C46042 a_19963_31679# a_22400_42852# 3.97e-20
C46043 a_5013_44260# a_5326_44056# 7.61e-19
C46044 a_n2810_45572# a_n4209_38502# 0.066112f
C46045 a_n1059_45260# a_16245_42852# 0.130348f
C46046 a_n913_45002# a_15953_42852# 1.61e-20
C46047 a_n2017_45002# a_16877_42852# 5.23e-19
C46048 a_3147_46376# VDD 0.341038f
C46049 a_17737_43940# a_18079_43940# 0.001885f
C46050 a_14539_43914# a_17499_43370# 0.005043f
C46051 a_18114_32519# a_14209_32519# 0.054602f
C46052 a_17730_32519# a_20974_43370# 0.016457f
C46053 a_2324_44458# a_2304_45348# 1.74e-19
C46054 a_n2497_47436# a_n1177_43370# 0.062743f
C46055 SMPL_ON_P a_n2433_43396# 2.87e-19
C46056 a_11652_45724# a_11823_42460# 0.035142f
C46057 a_11962_45724# a_12427_45724# 0.064229f
C46058 a_2711_45572# a_15297_45822# 1.6e-19
C46059 a_n357_42282# a_18479_45785# 2.83e-19
C46060 a_11415_45002# a_20193_45348# 0.007211f
C46061 a_18597_46090# a_20935_43940# 0.008467f
C46062 a_13507_46334# a_15493_43396# 2.29e-20
C46063 a_5066_45546# a_3537_45260# 1.14e-19
C46064 a_3483_46348# a_13711_45394# 0.002278f
C46065 a_n2293_46634# a_n809_44244# 5.01e-20
C46066 a_18479_47436# a_11341_43940# 0.009284f
C46067 a_10193_42453# a_13249_42308# 0.001874f
C46068 a_8162_45546# a_6977_45572# 1.1e-19
C46069 a_5937_45572# a_7418_45394# 2.23e-19
C46070 a_n2438_43548# a_n2472_43914# 0.032003f
C46071 a_10227_46804# a_15493_43940# 0.00594f
C46072 a_n4064_38528# a_n3420_37440# 0.050813f
C46073 a_n3420_38528# a_n4064_37440# 0.045626f
C46074 a_n4209_39590# a_n1838_35608# 2.05e-19
C46075 a_4958_30871# C8_N_btm 0.001147f
C46076 a_7174_31319# C5_P_btm 3.27e-20
C46077 a_n4064_40160# EN_VIN_BSTR_P 0.187697f
C46078 a_17124_42282# RST_Z 4.07e-20
C46079 a_7754_39964# VDAC_Pi 0.001576f
C46080 a_15811_47375# a_n881_46662# 1.05e-19
C46081 a_2063_45854# a_n2293_46634# 0.004931f
C46082 a_2905_45572# a_n2661_46634# 0.029475f
C46083 a_4883_46098# a_11453_44696# 0.071224f
C46084 a_6151_47436# a_5807_45002# 0.099462f
C46085 a_13381_47204# a_12891_46348# 0.002658f
C46086 a_11459_47204# a_12549_44172# 1.19e-20
C46087 a_9313_45822# a_768_44030# 2.99e-20
C46088 a_n1435_47204# a_11309_47204# 1.78e-20
C46089 a_n785_47204# a_n133_46660# 0.001087f
C46090 a_327_47204# a_n2438_43548# 2.1e-19
C46091 a_1209_47178# a_n743_46660# 9.52e-20
C46092 a_n971_45724# a_383_46660# 1.21e-19
C46093 a_n237_47217# a_33_46660# 7.19e-21
C46094 a_n23_47502# a_171_46873# 0.001553f
C46095 a_n746_45260# a_601_46902# 0.004287f
C46096 a_12465_44636# a_22731_47423# 0.002949f
C46097 a_1431_47204# a_n1925_46634# 1.02e-20
C46098 a_9313_44734# a_17749_42852# 6.88e-20
C46099 a_13249_42308# VDD 0.653917f
C46100 a_11341_43940# a_4190_30871# 0.00376f
C46101 a_14021_43940# a_16664_43396# 0.003073f
C46102 a_20512_43084# a_19987_42826# 0.11919f
C46103 a_n97_42460# a_2437_43396# 1.3e-19
C46104 a_8746_45002# CLK 0.018523f
C46105 a_3422_30871# a_22223_42860# 0.002205f
C46106 a_7845_44172# a_7765_42852# 1.24e-19
C46107 a_19862_44208# a_13467_32519# 2.46e-19
C46108 a_20623_43914# a_20556_43646# 3.65e-19
C46109 a_n2810_45028# a_n2216_37984# 3.1e-19
C46110 a_n2956_37592# a_n2860_37984# 9.05e-19
C46111 a_10193_42453# a_17613_45144# 2.06e-20
C46112 a_n2293_45010# a_n2109_45247# 0.068458f
C46113 a_n2661_45010# a_n1059_45260# 0.021417f
C46114 a_n2472_45002# a_n2017_45002# 4.25e-20
C46115 a_n2293_46634# a_14955_43396# 0.002132f
C46116 a_17339_46660# a_15493_43940# 0.020994f
C46117 a_3090_45724# a_10555_43940# 0.005028f
C46118 a_8049_45260# a_n2661_43922# 2.89e-19
C46119 a_8696_44636# a_1423_45028# 0.095059f
C46120 a_11823_42460# a_13490_45067# 6.19e-21
C46121 a_3483_46348# a_5013_44260# 0.002821f
C46122 a_13661_43548# a_13749_43396# 1.53e-20
C46123 a_n357_42282# a_10057_43914# 9.91e-20
C46124 a_n443_42852# a_949_44458# 0.0015f
C46125 a_1609_45822# a_742_44458# 2.73e-20
C46126 a_13059_46348# a_12495_44260# 2e-20
C46127 a_12549_44172# a_18525_43370# 3.14e-20
C46128 a_21513_45002# a_413_45260# 2.28e-21
C46129 a_4185_45028# a_3905_42865# 0.09316f
C46130 RST_Z CLK 0.064624f
C46131 a_18597_46090# a_20202_43084# 0.04177f
C46132 a_n2109_47186# a_2324_44458# 0.004259f
C46133 a_3877_44458# a_5429_46660# 0.00211f
C46134 a_13661_43548# a_19333_46634# 0.011985f
C46135 a_13747_46662# a_15227_44166# 0.05203f
C46136 a_12891_46348# a_13170_46660# 2.99e-19
C46137 a_12549_44172# a_12925_46660# 3.4e-20
C46138 a_4915_47217# a_4704_46090# 5.74e-20
C46139 a_6545_47178# a_3483_46348# 2.08e-20
C46140 a_n881_46662# a_13059_46348# 0.642888f
C46141 a_10227_46804# a_12741_44636# 0.188309f
C46142 a_5385_46902# a_5275_47026# 0.097745f
C46143 a_5907_46634# a_6540_46812# 0.017547f
C46144 a_5167_46660# a_5072_46660# 0.049827f
C46145 VDD VIN_P 1.47957f
C46146 a_n2661_46634# a_12816_46660# 5.55e-19
C46147 C10_N_btm VREF 14.773f
C46148 a_n1151_42308# a_8016_46348# 0.580516f
C46149 a_4791_45118# a_5164_46348# 0.42219f
C46150 a_n443_46116# a_5068_46348# 9.9e-19
C46151 a_2063_45854# a_9625_46129# 0.001267f
C46152 a_5807_45002# a_19466_46812# 0.178376f
C46153 C9_N_btm VREF_GND 5.18245f
C46154 C8_N_btm VCM 2.61094f
C46155 a_13507_46334# a_18900_46660# 9.83e-19
C46156 a_11453_44696# a_21188_46660# 0.047802f
C46157 a_3626_43646# a_3863_42891# 5.26e-19
C46158 a_n97_42460# a_15785_43172# 3.4e-19
C46159 a_13887_32519# a_14209_32519# 0.086073f
C46160 a_5649_42852# a_17364_32525# 6.86e-20
C46161 a_17613_45144# VDD 0.094022f
C46162 a_14955_43396# a_5342_30871# 0.002466f
C46163 a_10341_43396# a_5534_30871# 2.97e-19
C46164 a_15095_43370# a_15567_42826# 0.167909f
C46165 a_3457_43396# a_n2293_42282# 3.86e-19
C46166 a_19721_31679# a_18194_35068# 1e-19
C46167 a_3065_45002# a_n356_44636# 2.39e-19
C46168 a_16147_45260# a_11967_42832# 6.48e-20
C46169 a_3090_45724# a_13113_42826# 0.003304f
C46170 a_768_44030# a_961_42354# 1.48e-21
C46171 a_10903_43370# a_9145_43396# 0.041756f
C46172 a_n357_42282# a_14021_43940# 3.16e-19
C46173 a_2711_45572# a_18079_43940# 0.006173f
C46174 a_413_45260# a_700_44734# 3.75e-19
C46175 a_n2661_45010# a_484_44484# 0.002755f
C46176 a_n443_42852# a_11341_43940# 0.51832f
C46177 a_9290_44172# a_14579_43548# 0.007608f
C46178 SMPL_ON_P a_n4064_40160# 2.22e-19
C46179 a_8953_45546# a_9885_43646# 0.011162f
C46180 a_12861_44030# a_15803_42450# 5.43e-20
C46181 a_526_44458# a_n1557_42282# 0.31675f
C46182 a_1307_43914# a_4223_44672# 0.747516f
C46183 a_6945_45028# a_6765_43638# 4.3e-20
C46184 a_11787_45002# a_8975_43940# 4.91e-20
C46185 a_9482_43914# a_9838_44484# 0.175591f
C46186 a_5257_43370# a_5837_43172# 3.27e-20
C46187 a_20202_43084# a_743_42282# 0.135735f
C46188 a_10227_46804# a_5742_30871# 6.15e-19
C46189 a_3357_43084# a_n2661_42834# 0.081135f
C46190 a_17339_46660# a_12741_44636# 0.032832f
C46191 a_18285_46348# a_11415_45002# 1.48e-20
C46192 a_20273_46660# a_21350_47026# 1.46e-19
C46193 a_20411_46873# a_20719_46660# 2.12e-19
C46194 a_4883_46098# a_5907_45546# 2.75e-20
C46195 a_4817_46660# a_526_44458# 4.05e-20
C46196 a_4955_46873# a_n1925_42282# 6.24e-20
C46197 a_19321_45002# a_19443_46116# 0.003684f
C46198 a_12861_44030# a_10193_42453# 1.83e-19
C46199 a_11459_47204# a_11525_45546# 1.91e-21
C46200 a_n743_46660# a_11601_46155# 6.77e-19
C46201 a_5649_42852# a_8325_42308# 7.52e-20
C46202 a_16547_43609# a_16522_42674# 4.2e-20
C46203 a_16243_43396# a_17124_42282# 1.48e-20
C46204 a_15743_43084# a_15890_42674# 0.001174f
C46205 a_4361_42308# a_9223_42460# 0.009506f
C46206 a_18083_42858# a_18707_42852# 9.73e-19
C46207 a_18817_42826# a_18861_43218# 3.69e-19
C46208 a_18249_42858# a_19273_43230# 2.36e-20
C46209 a_10341_43396# a_19647_42308# 2.22e-20
C46210 a_8952_43230# a_n784_42308# 1.44e-22
C46211 a_3681_42891# a_1755_42282# 1.9e-20
C46212 a_743_42282# a_10545_42558# 7.22e-19
C46213 a_n1441_43940# VDD 0.142719f
C46214 a_17970_44736# a_16241_44734# 1.65e-20
C46215 a_1307_43914# a_15493_43940# 0.057588f
C46216 SMPL_ON_N a_11530_34132# 2.32e-19
C46217 a_16979_44734# a_17517_44484# 0.109784f
C46218 a_5891_43370# a_5708_44484# 4.97e-20
C46219 a_n2293_42834# a_7911_44260# 0.00163f
C46220 a_10193_42453# a_19700_43370# 7.43e-21
C46221 a_n443_42852# a_n1076_43230# 0.003517f
C46222 a_n755_45592# a_1847_42826# 0.053279f
C46223 a_526_44458# a_8483_43230# 0.004236f
C46224 a_6575_47204# DATA[4] 0.15718f
C46225 a_9482_43914# a_12603_44260# 0.002516f
C46226 a_15227_44166# a_4958_30871# 1.39e-20
C46227 a_5111_44636# a_5745_43940# 5.27e-19
C46228 a_5147_45002# a_5829_43940# 6.15e-19
C46229 a_7640_43914# a_9159_44484# 8.4e-20
C46230 a_5289_44734# a_n2661_43922# 1.98e-35
C46231 a_12861_44030# VDD 3.56689f
C46232 a_18114_32519# a_17730_32519# 9.1497f
C46233 a_3537_45260# a_8415_44056# 3.72e-19
C46234 a_1138_42852# a_1184_42692# 0.00134f
C46235 a_13717_47436# RST_Z 4.51263f
C46236 a_18189_46348# a_8049_45260# 0.030061f
C46237 a_10903_43370# a_14180_46482# 0.001228f
C46238 a_n2293_46098# a_3316_45546# 0.008121f
C46239 SMPL_ON_P a_n2433_44484# 2.73e-19
C46240 a_n2661_46634# a_n37_45144# 2.93e-21
C46241 a_n2293_46634# a_n955_45028# 4.55e-21
C46242 a_n2497_47436# a_n1177_44458# 1.74e-19
C46243 a_472_46348# a_380_45546# 3.1e-21
C46244 a_376_46348# a_n1099_45572# 6.04e-21
C46245 a_167_45260# a_n2661_45546# 0.084316f
C46246 a_1138_42852# a_n2293_45546# 0.021487f
C46247 a_5807_45002# a_5111_44636# 0.204193f
C46248 a_2443_46660# a_2437_43646# 3.88e-20
C46249 a_n881_46662# a_13556_45296# 4.04e-20
C46250 a_11189_46129# a_11601_46155# 0.007009f
C46251 a_12594_46348# a_12379_46436# 0.04209f
C46252 a_14209_32519# EN_VIN_BSTR_N 0.032853f
C46253 a_7963_42308# a_8325_42308# 0.002341f
C46254 a_6123_31319# a_8685_42308# 1.64e-19
C46255 a_4190_30871# C1_P_btm 7.67e-20
C46256 a_19700_43370# VDD 0.28578f
C46257 a_5343_44458# a_7112_43396# 1.78e-21
C46258 a_n4318_39768# a_n3674_39768# 3.06574f
C46259 a_20820_30879# a_22609_38406# 5.26e-21
C46260 a_n1059_45260# a_18249_42858# 0.002769f
C46261 a_n913_45002# a_17333_42852# 2.15e-20
C46262 a_n2017_45002# a_18817_42826# 0.018518f
C46263 a_11691_44458# a_10341_43396# 1.54e-19
C46264 a_13259_45724# a_13258_32519# 0.037974f
C46265 a_5883_43914# a_6293_42852# 4.78e-19
C46266 a_2675_43914# a_3499_42826# 0.010775f
C46267 a_2998_44172# a_2253_44260# 2.04e-20
C46268 a_3357_43084# a_n2293_42282# 0.146926f
C46269 a_n23_44458# a_n229_43646# 8.22e-20
C46270 a_n356_44636# a_458_43396# 0.001988f
C46271 a_14180_46812# VDD 0.755623f
C46272 a_6298_44484# a_6547_43396# 0.002809f
C46273 a_18579_44172# a_15493_43940# 0.377126f
C46274 a_n2661_44458# a_8685_43396# 3.35e-20
C46275 a_n2956_38680# a_n2946_38778# 0.14863f
C46276 a_n2956_39304# a_n4064_38528# 0.001421f
C46277 a_13249_42308# a_n784_42308# 1.26e-20
C46278 a_n357_42282# a_15764_42576# 8.52e-20
C46279 a_10425_46660# CLK 1.87e-19
C46280 a_3232_43370# a_9127_43156# 4.38e-21
C46281 a_375_42282# a_n1076_43230# 1.84e-20
C46282 a_14035_46660# RST_Z 1.33e-19
C46283 a_8049_45260# a_17478_45572# 0.010438f
C46284 a_4704_46090# a_4574_45260# 1.1e-20
C46285 a_15227_44166# a_18911_45144# 3.32e-20
C46286 a_2711_45572# a_4099_45572# 0.176427f
C46287 a_n2442_46660# a_n2661_43922# 1.33e-20
C46288 a_n2293_46634# a_n2661_42834# 0.025484f
C46289 a_17715_44484# a_3357_43084# 9.87e-21
C46290 a_n443_46116# a_2537_44260# 5.68e-19
C46291 a_n1151_42308# a_7584_44260# 9.64e-20
C46292 a_12741_44636# a_1307_43914# 0.05146f
C46293 a_5068_46348# a_3537_45260# 1.38e-20
C46294 a_4419_46090# a_4558_45348# 0.00116f
C46295 a_18819_46122# a_2437_43646# 2.62e-20
C46296 a_3483_46348# a_4927_45028# 0.032156f
C46297 a_4185_45028# a_5147_45002# 5.45e-19
C46298 a_10903_43370# a_n1059_45260# 0.028694f
C46299 a_19466_46812# a_18315_45260# 9.44e-20
C46300 a_6151_47436# a_14311_47204# 0.136645f
C46301 a_15764_42576# CAL_N 9.17e-19
C46302 a_5932_42308# C5_P_btm 5.59e-19
C46303 a_n784_42308# VIN_P 0.004358f
C46304 a_7227_47204# a_n1435_47204# 0.001005f
C46305 a_9067_47204# a_9313_45822# 0.013659f
C46306 a_n3565_39304# a_n4064_38528# 0.029566f
C46307 a_n3420_39072# a_n3420_38528# 0.127439f
C46308 a_n4064_39072# a_n3565_38502# 0.030685f
C46309 a_6123_31319# C10_P_btm 1.34e-19
C46310 a_2123_42473# VDD 0.1936f
C46311 a_n1920_47178# a_n2312_39304# 0.157528f
C46312 a_n1741_47186# a_n2312_40392# 4.79e-19
C46313 a_n2109_47186# a_n310_47570# 9.67e-19
C46314 a_n3565_39590# a_n2302_37984# 8.95e-20
C46315 a_22591_44484# a_22591_43396# 2.73e-20
C46316 a_22485_44484# a_14209_32519# 4.86e-19
C46317 a_17730_32519# a_13887_32519# 0.053953f
C46318 a_13857_44734# a_13635_43156# 2.1e-21
C46319 a_n2293_43922# a_5534_30871# 0.271171f
C46320 a_1307_43914# a_5742_30871# 2.36e-20
C46321 en_comp a_21335_42336# 2.22e-20
C46322 a_310_45028# VDD 0.360949f
C46323 a_20692_30879# VIN_N 0.039f
C46324 a_13565_43940# a_n97_42460# 1.86e-21
C46325 a_20974_43370# a_17538_32519# 0.001842f
C46326 a_14955_43940# a_9145_43396# 1.77e-19
C46327 a_9313_44734# a_19339_43156# 0.01152f
C46328 a_20205_31679# VREF 0.056031f
C46329 a_18175_45572# a_20107_45572# 4.32e-19
C46330 a_18909_45814# a_19418_45938# 2.6e-19
C46331 a_18341_45572# a_18787_45572# 2.28e-19
C46332 a_18479_45785# a_18953_45572# 0.002424f
C46333 a_11453_44696# a_8685_43396# 9.12e-22
C46334 a_12861_44030# a_16137_43396# 3.28e-19
C46335 a_7227_45028# a_1423_45028# 0.009712f
C46336 a_2711_45572# a_5365_45348# 3.34e-19
C46337 a_768_44030# a_2982_43646# 0.0012f
C46338 a_8953_45546# a_n2661_43922# 0.024071f
C46339 a_20254_46482# a_18494_42460# 2.45e-20
C46340 a_4883_46098# a_9145_43396# 0.02956f
C46341 a_n2497_47436# a_n1991_42858# 9.6e-20
C46342 a_2063_45854# a_743_42282# 1.93e-20
C46343 a_n1613_43370# a_6197_43396# 0.03252f
C46344 a_n2438_43548# a_n2433_43396# 0.415301f
C46345 a_2957_45546# a_n2661_43370# 3.26e-20
C46346 a_10490_45724# a_10775_45002# 1.62e-19
C46347 a_12741_44636# a_18579_44172# 0.002357f
C46348 a_18479_47436# a_10341_43396# 1.96e-19
C46349 a_13259_45724# a_20193_45348# 0.014145f
C46350 a_11415_45002# a_20596_44850# 8.83e-20
C46351 a_3090_45724# a_n2661_42282# 0.039366f
C46352 a_13527_45546# a_6171_45002# 3.83e-20
C46353 a_8746_45002# a_10951_45334# 7.44e-20
C46354 a_10193_42453# a_11787_45002# 0.0195f
C46355 a_n3420_37440# VREF_GND 0.033872f
C46356 a_16327_47482# a_15368_46634# 2.32e-20
C46357 a_n743_46660# a_288_46660# 0.024827f
C46358 a_11206_38545# VDD 8.87267f
C46359 a_11530_34132# a_19864_35138# 0.201937f
C46360 VDAC_P RST_Z 0.158793f
C46361 a_15673_47210# a_16292_46812# 1.35e-19
C46362 a_15811_47375# a_17609_46634# 4.73e-20
C46363 a_n133_46660# a_2107_46812# 2.94e-21
C46364 a_n2438_43548# a_1983_46706# 0.057412f
C46365 a_n1925_46634# a_n935_46688# 6.05e-19
C46366 a_n2661_46634# a_2443_46660# 0.021792f
C46367 EN_VIN_BSTR_P C10_P_btm 0.320569f
C46368 a_n881_46662# a_7577_46660# 0.028487f
C46369 EN_VIN_BSTR_N a_19120_35138# 0.652984f
C46370 a_2905_45572# a_765_45546# 0.039575f
C46371 a_n2472_46634# a_n2661_46098# 2.78e-21
C46372 a_171_46873# a_948_46660# 5.47e-21
C46373 a_33_46660# a_1123_46634# 0.041798f
C46374 a_601_46902# a_383_46660# 0.209641f
C46375 a_11599_46634# a_15227_44166# 0.101252f
C46376 a_10227_46804# a_13607_46688# 0.027032f
C46377 a_21381_43940# a_19987_42826# 1.97e-19
C46378 a_n2661_42282# a_n2472_42282# 0.028691f
C46379 a_11787_45002# VDD 0.153399f
C46380 a_14955_43396# a_743_42282# 3.11e-20
C46381 a_10341_43396# a_4190_30871# 0.090771f
C46382 a_2889_44172# a_2903_42308# 3.69e-22
C46383 a_17499_43370# a_17324_43396# 0.234322f
C46384 a_16547_43609# a_15743_43084# 0.028834f
C46385 a_11967_42832# a_15051_42282# 1.9e-19
C46386 a_9313_44734# a_22465_38105# 0.002447f
C46387 a_3232_43370# CLK 2.72e-19
C46388 a_n97_42460# a_5534_30871# 0.109695f
C46389 a_2982_43646# a_5755_42852# 1.01e-20
C46390 a_3626_43646# a_4520_42826# 4.31e-20
C46391 a_3539_42460# a_3935_42891# 2.26e-20
C46392 a_11341_43940# a_14635_42282# 4.84e-20
C46393 a_4646_46812# a_8952_43230# 3.88e-21
C46394 a_3090_45724# a_16823_43084# 7.78e-20
C46395 a_13017_45260# a_13490_45394# 2.62e-19
C46396 a_3483_46348# a_4699_43561# 2.57e-21
C46397 a_4185_45028# a_4093_43548# 4.24e-20
C46398 a_n443_42852# a_175_44278# 0.003303f
C46399 a_n2840_45002# a_n2661_44458# 0.003602f
C46400 a_n2661_45010# a_n4318_40392# 8.18e-22
C46401 a_2437_43646# a_949_44458# 0.038046f
C46402 a_n2293_46634# a_n2293_42282# 7.31e-22
C46403 a_2304_45348# a_2448_45028# 6.84e-19
C46404 a_9482_43914# a_n2661_43370# 2.58e-19
C46405 a_1307_43914# a_n2293_42834# 0.089964f
C46406 a_1823_45246# a_1987_43646# 2.6e-20
C46407 a_6171_45002# a_16922_45042# 0.00895f
C46408 a_10193_42453# a_17325_44484# 1.97e-19
C46409 a_413_45260# a_22959_45036# 0.024709f
C46410 a_13507_46334# a_18707_42852# 6.67e-19
C46411 a_18909_45814# a_18248_44752# 1.74e-19
C46412 a_18479_45785# a_18443_44721# 7.52e-19
C46413 a_18175_45572# a_18374_44850# 3.73e-19
C46414 a_18341_45572# a_18287_44626# 3.7e-20
C46415 a_n2956_38216# a_n3674_39768# 0.031697f
C46416 a_n357_42282# a_5013_44260# 2.45e-20
C46417 a_3316_45546# a_2675_43914# 4.27e-20
C46418 a_5937_45572# a_n97_42460# 1.46e-20
C46419 a_13059_46348# a_14621_43646# 2.44e-20
C46420 a_4791_45118# a_3318_42354# 2.33e-20
C46421 a_n443_46116# a_2903_42308# 7.96e-21
C46422 a_16327_47482# a_19597_46482# 0.001903f
C46423 a_n1925_46634# a_2324_44458# 8.77e-20
C46424 a_n1741_47186# a_6472_45840# 9.06e-21
C46425 a_2063_45854# a_2277_45546# 0.057116f
C46426 a_n443_46116# a_3218_45724# 9.08e-19
C46427 a_n1151_42308# a_n1013_45572# 0.002324f
C46428 a_10249_46116# a_11415_45002# 1.8e-20
C46429 a_n881_46662# a_5431_46482# 9.41e-19
C46430 a_12816_46660# a_765_45546# 3.23e-20
C46431 a_n1613_43370# a_5066_45546# 0.015391f
C46432 a_4883_46098# a_14180_46482# 0.001483f
C46433 a_10227_46804# a_16375_45002# 7.63e-19
C46434 a_19594_46812# a_6945_45028# 0.014072f
C46435 a_n237_47217# a_1609_45572# 2.16e-20
C46436 a_584_46384# a_1990_45899# 4.9e-19
C46437 a_3877_44458# a_3483_46348# 0.083955f
C46438 a_16292_46812# a_16388_46812# 0.318472f
C46439 a_n743_46660# a_15015_46420# 0.007103f
C46440 a_8685_43396# a_8325_42308# 3.75e-20
C46441 a_3422_30871# C6_P_btm 2.2e-19
C46442 a_18817_42826# a_19164_43230# 0.051162f
C46443 a_5755_42852# a_5837_42852# 0.171361f
C46444 a_8387_43230# a_8292_43218# 0.049827f
C46445 a_8605_42826# a_8483_43230# 3.16e-19
C46446 a_n97_42460# a_19647_42308# 6.61e-19
C46447 a_17730_32519# EN_VIN_BSTR_N 0.072552f
C46448 a_526_44458# a_3935_42891# 0.012937f
C46449 a_n1925_42282# a_3681_42891# 9.76e-21
C46450 a_n2312_38680# a_n4209_39590# 0.020921f
C46451 a_8270_45546# a_5934_30871# 2.28e-21
C46452 a_n2442_46660# a_n3690_39616# 5.77e-19
C46453 a_1823_45246# a_4649_42852# 0.042816f
C46454 a_15004_44636# a_14539_43914# 0.001002f
C46455 a_375_42282# a_175_44278# 0.017991f
C46456 a_626_44172# a_n809_44244# 1.91e-19
C46457 a_n913_45002# a_13483_43940# 9.64e-21
C46458 a_n1059_45260# a_14955_43940# 8.05e-22
C46459 a_n2017_45002# a_15682_43940# 2.7e-20
C46460 a_11691_44458# a_n2293_43922# 0.02314f
C46461 a_1307_43914# a_1115_44172# 0.115939f
C46462 a_n2661_44458# a_8783_44734# 1.49e-19
C46463 a_n2956_39768# a_n4064_39616# 0.058734f
C46464 a_n443_42852# a_10341_43396# 0.23026f
C46465 a_4883_46098# a_n1059_45260# 0.001764f
C46466 a_10903_43370# a_13925_46122# 0.001937f
C46467 a_12594_46348# a_13351_46090# 2.97e-19
C46468 a_472_46348# a_526_44458# 3.38e-21
C46469 a_1208_46090# a_1431_46436# 0.011458f
C46470 a_1176_45822# a_1337_46436# 9.42e-19
C46471 a_4915_47217# a_9482_43914# 0.269756f
C46472 a_10227_46804# a_413_45260# 3.82e-19
C46473 a_n2293_46098# a_5066_45546# 0.140248f
C46474 a_19692_46634# a_n357_42282# 1.03e-19
C46475 a_20202_43084# a_8049_45260# 0.042894f
C46476 a_5807_45002# a_16147_45260# 3.67e-19
C46477 a_18285_46348# a_13259_45724# 3.76e-21
C46478 a_17339_46660# a_16375_45002# 0.0296f
C46479 a_7577_46660# a_8162_45546# 5.56e-21
C46480 a_n743_46660# a_16333_45814# 0.014466f
C46481 a_10355_46116# a_2324_44458# 3.32e-21
C46482 a_n4318_38680# a_n4334_38304# 3.4e-19
C46483 a_21195_42852# a_21613_42308# 7.21e-19
C46484 a_21671_42860# a_21887_42336# 1.89e-21
C46485 a_1576_42282# a_1184_42692# 0.033078f
C46486 a_3080_42308# VIN_P 0.025929f
C46487 a_n784_42308# a_2123_42473# 0.216332f
C46488 a_n998_43396# VDD 6.7e-20
C46489 a_n1630_35242# a_1149_42558# 2.88e-20
C46490 a_n473_42460# a_n327_42308# 0.013377f
C46491 a_1067_42314# a_961_42354# 0.13675f
C46492 a_6171_45002# a_15743_43084# 1.19e-20
C46493 a_5894_47026# VDD 4.6e-19
C46494 a_1307_43914# a_10849_43646# 9.39e-19
C46495 a_11691_44458# a_n97_42460# 1.21e-19
C46496 a_n2661_43922# a_9028_43914# 3.15e-20
C46497 a_n2661_42834# a_9672_43914# 0.009389f
C46498 a_22485_44484# a_17730_32519# 0.091577f
C46499 a_n2661_43370# a_6031_43396# 4.62e-21
C46500 a_18114_32519# a_17538_32519# 0.052981f
C46501 a_5883_43914# a_7499_43940# 0.04798f
C46502 a_n755_45592# a_n473_42460# 0.061354f
C46503 a_n357_42282# a_196_42282# 0.033292f
C46504 a_n863_45724# a_n1630_35242# 3.34e-20
C46505 a_n913_45002# a_13678_32519# 0.023168f
C46506 a_n1059_45260# a_5649_42852# 0.030637f
C46507 a_7715_46873# a_n2661_43370# 3.07e-20
C46508 a_14976_45028# a_14797_45144# 0.137651f
C46509 a_3090_45724# a_15415_45028# 0.009288f
C46510 a_n2497_47436# a_n1331_43914# 0.003514f
C46511 a_11415_45002# a_22223_45572# 0.021019f
C46512 a_22591_46660# a_2437_43646# 7.95e-19
C46513 SMPL_ON_P a_n2840_43914# 9.38e-19
C46514 a_n1613_43370# a_n1821_44484# 9.54e-19
C46515 a_10227_46804# a_13468_44734# 7.33e-20
C46516 a_20202_43084# a_19479_31679# 9.39e-20
C46517 a_12549_44172# a_16979_44734# 1.34e-19
C46518 a_n2293_46634# a_n1352_44484# 2.08e-20
C46519 a_2324_44458# a_10544_45572# 2.77e-19
C46520 a_n2438_43548# a_n2433_44484# 0.421822f
C46521 a_13759_46122# a_14033_45822# 1.75e-20
C46522 a_n2956_38216# a_n2293_45546# 0.005455f
C46523 a_n2661_45546# a_n863_45724# 0.045552f
C46524 a_n784_42308# a_11206_38545# 3.18e-20
C46525 a_n452_47436# a_n746_45260# 0.187792f
C46526 a_n1741_47186# a_327_47204# 0.013765f
C46527 a_n2109_47186# a_1239_47204# 0.080115f
C46528 a_n815_47178# a_n237_47217# 0.005891f
C46529 SMPL_ON_P a_n785_47204# 1.53e-19
C46530 a_n1630_35242# a_6886_37412# 2.07e-19
C46531 a_8495_42852# VDD 0.132018f
C46532 COMP_P a_22521_40055# 7.41e-20
C46533 a_7174_31319# a_n4209_39590# 8.87e-22
C46534 a_20205_31679# a_22521_40599# 2.04e-20
C46535 a_9313_44734# a_22591_43396# 0.001502f
C46536 a_19478_44306# a_18533_43940# 3.55e-20
C46537 a_3065_45002# a_3823_42558# 0.198186f
C46538 a_n913_45002# a_6123_31319# 0.21316f
C46539 a_n1059_45260# a_7963_42308# 5.71e-20
C46540 a_9801_44260# a_9801_43940# 6.96e-20
C46541 a_11341_43940# a_11257_43940# 2.31e-19
C46542 a_3232_43370# a_1755_42282# 1.63e-20
C46543 a_n2661_42834# a_743_42282# 1.34e-20
C46544 a_15493_43396# a_19478_44056# 3.41e-19
C46545 a_n2017_45002# a_5934_30871# 0.007182f
C46546 a_19862_44208# a_19319_43548# 0.049274f
C46547 a_8975_43940# a_9127_43156# 8.61e-21
C46548 a_10334_44484# a_10518_42984# 1.38e-22
C46549 a_10440_44484# a_10083_42826# 9.38e-21
C46550 a_20708_46348# a_21005_45260# 1.01e-20
C46551 a_11387_46155# a_n2661_44458# 4.75e-21
C46552 a_n443_42852# a_n143_45144# 0.104427f
C46553 a_15037_45618# a_15225_45822# 7.47e-21
C46554 a_3503_45724# a_3065_45002# 9.76e-20
C46555 a_3316_45546# a_3429_45260# 0.142842f
C46556 a_n755_45592# a_5111_44636# 0.004145f
C46557 a_5257_43370# a_3905_42865# 0.106385f
C46558 a_584_46384# a_3457_43396# 0.120485f
C46559 a_4791_45118# a_6197_43396# 1.47e-19
C46560 a_3090_45724# a_19279_43940# 0.046663f
C46561 a_n1613_43370# a_8415_44056# 4.2e-21
C46562 a_16375_45002# a_1307_43914# 0.101951f
C46563 a_18819_46122# a_19113_45348# 5.65e-21
C46564 a_8034_45724# a_n2293_42834# 0.00209f
C46565 a_768_44030# a_2253_43940# 0.004046f
C46566 a_12549_44172# a_13569_47204# 0.005506f
C46567 a_12891_46348# a_13675_47204# 2.93e-20
C46568 a_n1435_47204# a_4955_46873# 4.48e-20
C46569 a_5815_47464# a_5257_43370# 8.52e-20
C46570 a_n3565_38502# VDD 0.762011f
C46571 a_4338_37500# a_5088_37509# 0.896828f
C46572 a_3726_37500# a_5700_37509# 0.574743f
C46573 a_n3565_39304# VREF_GND 0.010456f
C46574 a_n4064_37984# C3_P_btm 0.030933f
C46575 a_n3420_37984# C1_P_btm 1.26e-19
C46576 a_2063_45854# a_6755_46942# 0.131005f
C46577 a_4915_47217# a_7715_46873# 3.51e-19
C46578 a_n1151_42308# a_10428_46928# 0.011222f
C46579 a_14401_32519# a_14209_32519# 10.7535f
C46580 a_3626_43646# a_16409_43396# 3.02e-21
C46581 a_2982_43646# a_16759_43396# 7.55e-21
C46582 a_8685_43396# a_9145_43396# 0.201058f
C46583 a_18326_43940# a_18249_42858# 8.19e-22
C46584 a_15493_43396# a_17701_42308# 4.48e-20
C46585 a_18451_43940# a_17333_42852# 4.67e-20
C46586 a_18114_32519# a_22465_38105# 2.37e-19
C46587 a_11341_43940# a_14543_43071# 8.65e-21
C46588 a_3737_43940# a_3681_42891# 2.18e-20
C46589 a_20974_43370# a_22591_43396# 0.046632f
C46590 a_17538_32519# a_13887_32519# 0.051087f
C46591 a_5891_43370# a_9223_42460# 0.13879f
C46592 a_7542_44172# a_7309_42852# 6.74e-21
C46593 a_n97_42460# a_4190_30871# 0.140814f
C46594 a_3422_30871# a_20836_43172# 2.5e-20
C46595 a_n356_44636# a_13575_42558# 1.46e-19
C46596 a_n2661_42834# a_5755_42308# 1.09e-20
C46597 a_3232_43370# a_10951_45334# 5.7e-20
C46598 a_7229_43940# a_6709_45028# 0.136786f
C46599 a_5205_44484# a_8191_45002# 2.44e-20
C46600 a_8696_44636# a_16886_45144# 0.00316f
C46601 a_1138_42852# a_1443_43940# 7.84e-21
C46602 a_13527_45546# a_12607_44458# 8.08e-22
C46603 a_10193_42453# a_18287_44626# 5.37e-19
C46604 a_n443_42852# a_n2293_43922# 0.021367f
C46605 a_1609_45822# a_n2661_43922# 7.32e-20
C46606 a_16147_45260# a_18315_45260# 4.61e-19
C46607 a_13507_46334# a_21356_42826# 1.5e-19
C46608 a_768_44030# a_7871_42858# 8.9e-21
C46609 a_3090_45724# a_7112_43396# 0.004584f
C46610 a_18909_45814# a_16922_45042# 3.62e-20
C46611 a_15861_45028# a_16237_45028# 0.062212f
C46612 a_413_45260# a_1307_43914# 0.080885f
C46613 a_6171_45002# a_10775_45002# 0.008718f
C46614 a_11823_42460# a_13720_44458# 7.98e-20
C46615 a_3483_46348# a_13829_44260# 0.002792f
C46616 a_2063_45854# a_8049_45260# 0.037406f
C46617 a_n1151_42308# a_8283_46482# 0.003687f
C46618 a_2443_46660# a_765_45546# 0.004286f
C46619 a_6755_46942# a_12469_46902# 0.042969f
C46620 a_10249_46116# a_12251_46660# 1.57e-19
C46621 a_8128_46384# a_3483_46348# 1.2e-20
C46622 a_n881_46662# a_4704_46090# 0.049125f
C46623 a_11453_44696# a_11387_46155# 3.7e-21
C46624 a_4883_46098# a_13925_46122# 0.006732f
C46625 a_16327_47482# a_20708_46348# 0.001227f
C46626 a_4791_45118# a_5066_45546# 0.238282f
C46627 a_768_44030# a_1823_45246# 0.287407f
C46628 a_22612_30879# a_22959_46660# 6.06e-19
C46629 a_13507_46334# a_14275_46494# 0.004384f
C46630 a_10227_46804# a_18985_46122# 1.14e-20
C46631 a_15673_47210# a_6945_45028# 0.056077f
C46632 a_18597_46090# a_17715_44484# 2.16e-20
C46633 a_15507_47210# a_10809_44734# 6.3e-20
C46634 a_n1613_43370# a_5068_46348# 1.7e-19
C46635 a_21588_30879# a_21076_30879# 8.21286f
C46636 a_10341_43396# a_14635_42282# 1.31e-19
C46637 a_20269_44172# a_7174_31319# 7.85e-21
C46638 a_4361_42308# a_21195_42852# 0.020952f
C46639 a_13467_32519# a_21671_42860# 0.015185f
C46640 a_11341_43940# a_19511_42282# 3.14e-21
C46641 a_19862_44208# a_21335_42336# 6.38e-20
C46642 a_4905_42826# a_1755_42282# 1.01e-19
C46643 a_3080_42308# a_2123_42473# 3.08e-20
C46644 a_743_42282# a_n2293_42282# 0.058933f
C46645 a_8975_43940# CLK 1.38e-19
C46646 a_5649_42852# a_19987_42826# 3.08e-20
C46647 a_18287_44626# VDD 0.389383f
C46648 a_12741_44636# a_13635_43156# 1.35e-21
C46649 a_n443_42852# a_n97_42460# 0.822111f
C46650 a_14537_43396# a_15146_44811# 8.25e-19
C46651 a_n2661_43370# a_n1809_44850# 0.002228f
C46652 en_comp a_3422_30871# 0.357746f
C46653 a_n2017_45002# a_20512_43084# 4.16e-19
C46654 a_11415_45002# a_5534_30871# 4.51e-21
C46655 a_13249_42308# a_14021_43940# 0.07296f
C46656 a_n863_45724# a_1427_43646# 0.006268f
C46657 a_1423_45028# a_9159_44484# 0.037664f
C46658 a_17715_44484# a_743_42282# 1.09e-20
C46659 a_8696_44636# a_10405_44172# 2.24e-20
C46660 a_18114_32519# a_19721_31679# 0.051894f
C46661 a_375_42282# a_n2293_43922# 3e-19
C46662 a_626_44172# a_n2661_42834# 0.032386f
C46663 a_n357_42282# a_4699_43561# 1.83e-20
C46664 a_n755_45592# a_4235_43370# 6.26e-21
C46665 w_1575_34946# a_n83_35174# 0.001523f
C46666 a_n1925_46634# a_6667_45809# 1.11e-20
C46667 a_3877_44458# a_n357_42282# 1.85e-23
C46668 a_12549_44172# a_11823_42460# 0.624462f
C46669 a_768_44030# a_12427_45724# 1.64e-22
C46670 a_12891_46348# a_12791_45546# 0.012918f
C46671 a_1176_45822# a_1823_45246# 1.52e-20
C46672 a_1208_46090# a_2202_46116# 0.001619f
C46673 a_n971_45724# a_n2293_45010# 0.549225f
C46674 a_n746_45260# a_n2472_45002# 9.92e-21
C46675 SMPL_ON_P a_n913_45002# 1.07e-20
C46676 a_5807_45002# a_9049_44484# 8.47e-20
C46677 a_584_46384# a_3357_43084# 0.060446f
C46678 a_n1613_43370# a_6977_45572# 0.001505f
C46679 a_n743_46660# a_6472_45840# 0.006296f
C46680 a_n2661_46098# a_n443_42852# 9.75e-20
C46681 a_1799_45572# a_1609_45822# 0.079527f
C46682 a_2952_47436# a_2437_43646# 0.007981f
C46683 a_12861_44030# a_18479_45785# 0.058482f
C46684 a_n2497_47436# a_n967_45348# 0.021003f
C46685 a_472_46348# a_2521_46116# 5.15e-21
C46686 a_15227_46910# a_10809_44734# 0.006323f
C46687 a_16388_46812# a_6945_45028# 3.6e-19
C46688 a_8270_45546# a_9751_46155# 3.2e-20
C46689 a_18285_46348# a_18189_46348# 0.118603f
C46690 a_3992_43940# VDD 0.004127f
C46691 a_4190_30871# a_n3420_39616# 1.16e-20
C46692 a_13887_32519# a_22465_38105# 0.005089f
C46693 a_17538_32519# EN_VIN_BSTR_N 0.06758f
C46694 a_12379_42858# a_13575_42558# 1.06e-19
C46695 a_12545_42858# a_12563_42308# 1.83e-19
C46696 a_12089_42308# a_13070_42354# 9.69e-20
C46697 a_9290_44172# a_9223_42460# 2.46e-19
C46698 a_20193_45348# a_20935_43940# 0.016238f
C46699 a_16241_44734# a_16335_44484# 1.26e-19
C46700 a_11309_47204# DATA[5] 0.080873f
C46701 a_8953_45546# a_10545_42558# 2.8e-20
C46702 a_3483_46348# a_15486_42560# 6.47e-22
C46703 a_4185_45028# a_14113_42308# 1.2e-19
C46704 a_20202_43084# a_13258_32519# 0.685083f
C46705 a_375_42282# a_n97_42460# 0.039466f
C46706 a_3537_45260# a_6293_42852# 0.01772f
C46707 a_n356_44636# a_2479_44172# 8.76e-21
C46708 a_2711_45572# a_19339_43156# 0.020184f
C46709 a_n357_42282# a_6101_43172# 0.001097f
C46710 a_10037_47542# CLK 2.34e-19
C46711 a_18479_45785# a_19700_43370# 0.004581f
C46712 a_7499_43078# a_10835_43094# 0.028158f
C46713 a_n1059_45260# a_8685_43396# 0.036086f
C46714 a_17613_45144# a_14021_43940# 4.87e-21
C46715 a_13351_46090# a_2711_45572# 6.51e-20
C46716 a_5204_45822# a_5437_45600# 5.76e-19
C46717 a_3483_46348# a_10053_45546# 0.002243f
C46718 a_12991_46634# a_2437_43646# 9.73e-20
C46719 a_11453_44696# a_18545_45144# 2.11e-20
C46720 a_8049_45260# a_14383_46116# 0.002486f
C46721 a_768_44030# a_14309_45028# 3.22e-19
C46722 a_n1151_42308# a_n1243_44484# 1.58e-19
C46723 a_4185_45028# a_7499_43078# 2.72e-19
C46724 a_19466_46812# a_20107_45572# 0.283769f
C46725 a_n971_45724# a_9313_44734# 2.29e-20
C46726 a_11901_46660# a_3357_43084# 5.71e-20
C46727 a_15227_44166# a_20841_45814# 3.03e-19
C46728 a_10467_46802# a_413_45260# 1.23e-20
C46729 a_5429_46660# a_5111_44636# 5.34e-20
C46730 a_5257_43370# a_5147_45002# 0.836149f
C46731 a_9127_43156# VDD 0.468721f
C46732 a_5342_30871# C4_P_btm 8.98e-20
C46733 a_n3674_37592# a_n4209_38502# 7.92e-20
C46734 a_5932_42308# a_n4209_39590# 8.09e-22
C46735 a_15890_42674# a_16104_42674# 0.097745f
C46736 a_15803_42450# a_17124_42282# 0.00132f
C46737 a_15486_42560# a_15761_42308# 0.007416f
C46738 a_15959_42545# a_16522_42674# 0.049827f
C46739 a_14113_42308# a_16269_42308# 0.004499f
C46740 a_5534_30871# C2_P_btm 7.46e-20
C46741 a_5013_44260# a_5025_43940# 0.011829f
C46742 a_22485_44484# a_17538_32519# 0.002174f
C46743 a_17737_43940# a_17973_43940# 0.22264f
C46744 a_18287_44626# a_16137_43396# 8.65e-23
C46745 a_19721_31679# a_13887_32519# 0.051264f
C46746 a_18114_32519# a_22591_43396# 6.25e-19
C46747 a_10193_42453# a_17124_42282# 3.1e-19
C46748 a_n1059_45260# a_15953_42852# 0.005616f
C46749 a_n913_45002# a_15597_42852# 6.49e-20
C46750 a_n2017_45002# a_16245_42852# 0.003157f
C46751 a_5244_44056# a_5326_44056# 0.004767f
C46752 a_2804_46116# VDD 0.159351f
C46753 a_14539_43914# a_16759_43396# 0.012597f
C46754 a_626_44172# a_n2293_42282# 7.4e-21
C46755 a_17730_32519# a_14401_32519# 0.086728f
C46756 a_22591_44484# a_20974_43370# 6.26e-19
C46757 a_12861_44030# a_14021_43940# 0.035798f
C46758 a_n2497_47436# a_n1917_43396# 0.012526f
C46759 SMPL_ON_P a_n4318_39304# 0.039268f
C46760 a_2711_45572# a_15225_45822# 7.31e-20
C46761 a_n2438_43548# a_n2840_43914# 1.6e-21
C46762 a_8270_45546# a_8855_44734# 1.44e-35
C46763 a_11415_45002# a_11691_44458# 0.047412f
C46764 a_20202_43084# a_20193_45348# 0.116706f
C46765 a_10809_44734# a_9482_43914# 0.001033f
C46766 a_11525_45546# a_11823_42460# 0.001062f
C46767 a_11322_45546# a_12791_45546# 5.08e-20
C46768 a_3483_46348# a_13490_45394# 0.001975f
C46769 a_n2293_46634# a_n1549_44318# 9.06e-21
C46770 a_765_45546# a_949_44458# 3.16e-19
C46771 a_18479_47436# a_21115_43940# 0.001943f
C46772 a_n1925_42282# a_3232_43370# 0.021554f
C46773 a_7230_45938# a_6977_45572# 4.61e-19
C46774 a_8162_45546# a_6905_45572# 4.64e-20
C46775 a_8016_46348# a_n2293_42834# 6.15e-21
C46776 a_11453_44696# a_13483_43940# 1.03e-20
C46777 a_4419_46090# a_n2661_43370# 0.002591f
C46778 a_n3565_38502# a_n2302_37690# 6.13e-19
C46779 a_12465_44636# a_22223_47212# 0.175138f
C46780 a_584_46384# a_n2293_46634# 0.374996f
C46781 a_4915_47217# a_13747_46662# 0.710704f
C46782 a_11459_47204# a_12891_46348# 1.33e-19
C46783 a_4958_30871# C7_N_btm 1.47e-19
C46784 a_7174_31319# C6_P_btm 2.51e-19
C46785 a_n4064_39072# VDAC_P 0.002814f
C46786 a_15507_47210# a_n881_46662# 2.15e-19
C46787 a_n23_47502# a_n133_46660# 0.001147f
C46788 a_n785_47204# a_n2438_43548# 3.7e-19
C46789 a_327_47204# a_n743_46660# 9.48e-19
C46790 a_21496_47436# a_11453_44696# 4.71e-20
C46791 a_n1741_47186# a_1983_46706# 1.98e-20
C46792 a_n971_45724# a_601_46902# 1.1e-19
C46793 a_n746_45260# a_33_46660# 0.035747f
C46794 a_n237_47217# a_171_46873# 9.39e-20
C46795 a_1239_47204# a_n1925_46634# 4.34e-20
C46796 a_17124_42282# VDD 0.28176f
C46797 a_7845_44172# a_7871_42858# 5.57e-21
C46798 a_9313_44734# a_17665_42852# 5.16e-20
C46799 a_13904_45546# VDD 0.135068f
C46800 a_21115_43940# a_4190_30871# 0.01145f
C46801 a_14021_43940# a_19700_43370# 0.007203f
C46802 a_11341_43940# a_21259_43561# 0.00271f
C46803 a_20512_43084# a_19164_43230# 1.84e-20
C46804 a_10193_42453# CLK 0.023289f
C46805 a_3422_30871# a_22165_42308# 0.00669f
C46806 a_15493_43396# a_4361_42308# 3.03e-20
C46807 a_20623_43914# a_743_42282# 1.51e-19
C46808 a_6469_45572# a_n2661_43370# 3.64e-21
C46809 a_n2472_45002# a_n2109_45247# 0.001038f
C46810 a_n2661_45010# a_n2017_45002# 0.087596f
C46811 a_n2840_45002# a_n1059_45260# 2.05e-21
C46812 a_n2293_46634# a_15095_43370# 3.1e-19
C46813 a_3090_45724# a_9801_43940# 0.004765f
C46814 a_8049_45260# a_n2661_42834# 5.27e-20
C46815 a_10193_42453# a_17023_45118# 0.027968f
C46816 a_19963_31679# en_comp 1.68e-19
C46817 a_n357_42282# a_10440_44484# 1.65e-21
C46818 a_n443_42852# a_742_44458# 0.168627f
C46819 a_20708_46348# a_20835_44721# 1.53e-20
C46820 a_12549_44172# a_18429_43548# 3.26e-20
C46821 a_3483_46348# a_5244_44056# 2.37e-21
C46822 VCM VSS 40.3061f
C46823 VREF_GND VSS 17.4801f
C46824 VREF VSS 8.26148f
C46825 VIN_N VSS 13.1286f
C46826 VIN_P VSS 13.1075f
C46827 CLK VSS 1.55797f
C46828 EN_OFFSET_CAL VSS 0.505642f
C46829 DATA[5] VSS 0.561058f
C46830 DATA[4] VSS 0.755679f
C46831 DATA[3] VSS 1.01838f
C46832 DATA[2] VSS 0.536983f
C46833 DATA[1] VSS 0.550109f
C46834 DATA[0] VSS 0.616231f
C46835 CLK_DATA VSS 0.488979f
C46836 SINGLE_ENDED VSS 0.60168f
C46837 START VSS 0.991673f
C46838 RST_Z VSS 11.389f
C46839 VDD VSS 0.586439p
C46840 C10_N_btm VSS 0.264623p 
C46841 C9_N_btm VSS 0.114604p 
C46842 C8_N_btm VSS 60.275196f 
C46843 C7_N_btm VSS 32.1635f 
C46844 C6_N_btm VSS 17.8701f 
C46845 C5_N_btm VSS 10.4595f 
C46846 C4_N_btm VSS 7.67475f 
C46847 C3_N_btm VSS 5.70165f 
C46848 C2_N_btm VSS 4.38917f 
C46849 C1_N_btm VSS 3.94093f 
C46850 C0_N_btm VSS 5.62287f 
C46851 C0_dummy_N_btm VSS 4.25425f 
C46852 C0_dummy_P_btm VSS 4.26067f 
C46853 C0_P_btm VSS 5.63256f 
C46854 C1_P_btm VSS 3.96779f 
C46855 C2_P_btm VSS 4.40877f 
C46856 C3_P_btm VSS 5.70398f 
C46857 C4_P_btm VSS 7.68867f 
C46858 C5_P_btm VSS 10.4672f 
C46859 C6_P_btm VSS 17.865099f 
C46860 C7_P_btm VSS 32.1589f 
C46861 C8_P_btm VSS 60.269897f 
C46862 C9_P_btm VSS 0.114595p 
C46863 C10_P_btm VSS 0.264633p 
C46864 a_21589_35634# VSS 0.729455f 
C46865 a_19864_35138# VSS 1.75392f 
C46866 a_19120_35138# VSS 1.69667f 
C46867 a_18194_35068# VSS 2.11801f 
C46868 EN_VIN_BSTR_N VSS 9.03857f 
C46869 a_11530_34132# VSS 13.9862f 
C46870 a_n83_35174# VSS 1.72857f 
C46871 EN_VIN_BSTR_P VSS 9.263339f 
C46872 a_n923_35174# VSS 14.088f 
C46873 a_n1532_35090# VSS 2.16074f 
C46874 a_n1386_35608# VSS 1.75773f 
C46875 a_n1838_35608# VSS 0.737725f 
C46876 a_22717_36887# VSS 0.092029f 
C46877 a_22717_37285# VSS 0.095943f 
C46878 a_22705_37990# VSS 0.007968f 
C46879 a_22609_37990# VSS 0.473213f 
C46880 a_22705_38406# VSS 0.010928f 
C46881 a_22609_38406# VSS 0.588255f 
C46882 CAL_P VSS 11.418599f 
C46883 a_22876_39857# VSS 0.00127f 
C46884 a_22780_39857# VSS 7.39e-19 
C46885 a_22469_39537# VSS 2.5954f 
C46886 a_22821_38993# VSS 0.55301f 
C46887 a_22545_38993# VSS 0.35571f 
C46888 a_22521_39511# VSS 1.85851f 
C46889 a_22780_40081# VSS 0.002233f 
C46890 a_22459_39145# VSS 2.29285f 
C46891 a_22521_40055# VSS 1.21928f 
C46892 a_22780_40945# VSS 0.002478f 
C46893 a_22469_40625# VSS 1.56643f 
C46894 a_22521_40599# VSS 1.85568f 
C46895 CAL_N VSS 8.69238f 
C46896 a_11206_38545# VSS 0.713084f 
C46897 VDAC_P VSS 79.0997f 
C46898 a_8912_37509# VSS 3.72815f 
C46899 VDAC_N VSS 79.6318f 
C46900 a_6886_37412# VSS 3.84457f 
C46901 a_5700_37509# VSS 2.08109f 
C46902 a_5088_37509# VSS 2.72043f 
C46903 a_4338_37500# VSS 2.61369f 
C46904 a_3726_37500# VSS 4.48332f 
C46905 a_n3607_37440# VSS 0.002657f 
C46906 a_n4251_37440# VSS 0.003621f 
C46907 a_n2860_37690# VSS 0.001049f 
C46908 a_n2302_37690# VSS 0.514508f 
C46909 a_n4064_37440# VSS 1.7233f 
C46910 a_n2946_37690# VSS 0.517242f 
C46911 a_n3420_37440# VSS 5.23286f 
C46912 a_n3690_37440# VSS 0.548488f 
C46913 a_n3565_37414# VSS 3.15906f 
C46914 a_n4334_37440# VSS 0.561497f 
C46915 a_n4209_37414# VSS 3.16282f 
C46916 a_8530_39574# VSS 2.76228f 
C46917 a_7754_38470# VSS 3.24598f 
C46918 a_3754_38470# VSS 4.77654f 
C46919 VDAC_Ni VSS 2.86404f 
C46920 a_7754_38636# VSS 0.353706f 
C46921 a_3754_38802# VSS 0.390074f 
C46922 a_7754_38968# VSS 0.330037f 
C46923 a_3754_39134# VSS 0.401983f 
C46924 a_7754_39300# VSS 0.330682f 
C46925 a_3754_39466# VSS 0.401172f 
C46926 a_7754_39632# VSS 0.340942f 
C46927 VDAC_Pi VSS 3.50355f 
C46928 a_7754_39964# VSS 2.62481f 
C46929 a_7754_40130# VSS 2.84104f 
C46930 a_3754_39964# VSS 0.671366f 
C46931 a_n2860_37984# VSS 0.001049f 
C46932 a_2113_38308# VSS 2.64372f 
C46933 a_n3607_38304# VSS 0.002772f 
C46934 a_n4251_38304# VSS 0.003689f 
C46935 a_n2302_37984# VSS 0.483504f 
C46936 a_n4064_37984# VSS 1.65074f 
C46937 a_n2946_37984# VSS 0.485942f 
C46938 a_n3420_37984# VSS 1.75918f 
C46939 a_n3690_38304# VSS 0.517812f 
C46940 a_n3565_38216# VSS 1.48743f 
C46941 a_n4334_38304# VSS 0.529531f 
C46942 a_n4209_38216# VSS 3.03366f 
C46943 a_n3607_38528# VSS 0.002662f 
C46944 a_n4251_38528# VSS 0.003622f 
C46945 a_2684_37794# VSS 0.414596f 
C46946 a_1177_38525# VSS 0.641945f 
C46947 a_n2860_38778# VSS 0.001049f 
C46948 a_n2302_38778# VSS 0.483515f 
C46949 a_n4064_38528# VSS 1.69554f 
C46950 a_n2946_38778# VSS 0.485895f 
C46951 a_n3420_38528# VSS 2.03238f 
C46952 a_n3690_38528# VSS 0.516979f 
C46953 a_n3565_38502# VSS 1.55586f 
C46954 a_n4334_38528# VSS 0.529888f 
C46955 a_n4209_38502# VSS 3.0175f 
C46956 a_2112_39137# VSS 0.414248f 
C46957 a_n2860_39072# VSS 0.001051f 
C46958 comp_n VSS 0.568772f 
C46959 a_1736_39043# VSS 0.897653f 
C46960 a_1239_39043# VSS 0.614001f 
C46961 a_n3607_39392# VSS 0.002762f 
C46962 a_n4251_39392# VSS 0.003686f 
C46963 a_n2302_39072# VSS 0.483504f 
C46964 a_n4064_39072# VSS 1.71745f 
C46965 a_n2946_39072# VSS 0.486447f 
C46966 a_n3420_39072# VSS 2.21624f 
C46967 a_n3690_39392# VSS 0.517965f 
C46968 a_n3565_39304# VSS 1.4403f 
C46969 a_n4334_39392# VSS 0.529516f 
C46970 a_n4209_39304# VSS 3.21429f 
C46971 a_1343_38525# VSS 3.5734f 
C46972 a_n3607_39616# VSS 0.002672f 
C46973 a_n4251_39616# VSS 0.003625f 
C46974 a_1736_39587# VSS 1.10676f 
C46975 a_1239_39587# VSS 0.634559f 
C46976 a_n2860_39866# VSS 0.001465f 
C46977 a_n2302_39866# VSS 0.483537f 
C46978 a_n4064_39616# VSS 2.17764f 
C46979 a_n2946_39866# VSS 0.527929f 
C46980 a_n3420_39616# VSS 2.11206f 
C46981 a_n3690_39616# VSS 0.574329f 
C46982 a_n3565_39590# VSS 2.04547f 
C46983 a_n4334_39616# VSS 0.529903f 
C46984 a_n4209_39590# VSS 3.92629f 
C46985 a_n4251_40480# VSS 0.003684f 
C46986 a_n2302_40160# VSS 0.522244f 
C46987 a_n4064_40160# VSS 3.2951f 
C46988 a_n4334_40480# VSS 0.578721f 
C46989 a_n4315_30879# VSS 4.84874f 
C46990 a_21973_42336# VSS 0.004685f 
C46991 a_22465_38105# VSS 1.91115f 
C46992 a_21421_42336# VSS 0.004685f 
C46993 a_18997_42308# VSS 0.004143f 
C46994 a_22775_42308# VSS 0.602961f 
C46995 a_21613_42308# VSS 0.725408f 
C46996 a_21887_42336# VSS 0.234022f 
C46997 a_21335_42336# VSS 0.259392f 
C46998 a_7174_31319# VSS 5.51134f 
C46999 a_20712_42282# VSS 0.349662f 
C47000 a_20107_42308# VSS 0.344464f 
C47001 a_13258_32519# VSS 6.359931f 
C47002 a_19647_42308# VSS 0.313304f 
C47003 a_19511_42282# VSS 0.751141f 
C47004 a_18548_42308# VSS 0.005248f 
C47005 a_18310_42308# VSS 0.005141f 
C47006 a_18220_42308# VSS 0.003723f 
C47007 a_18214_42558# VSS 0.006283f 
C47008 a_19332_42282# VSS 0.31505f 
C47009 a_18907_42674# VSS 0.209311f 
C47010 a_18727_42674# VSS 0.233526f 
C47011 a_18057_42282# VSS 0.370712f 
C47012 a_17531_42308# VSS 0.253358f 
C47013 a_17303_42282# VSS 1.19698f 
C47014 a_4958_30871# VSS 5.01268f 
C47015 a_16269_42308# VSS 0.006939f 
C47016 a_16197_42308# VSS 0.004992f 
C47017 a_15761_42308# VSS 4.65e-19 
C47018 a_15521_42308# VSS 0.001281f 
C47019 a_17124_42282# VSS 0.332693f 
C47020 a_16522_42674# VSS 0.073862f 
C47021 a_16104_42674# VSS 0.004694f 
C47022 a_13921_42308# VSS 0.002122f 
C47023 a_13657_42308# VSS 0.006177f 
C47024 a_11897_42308# VSS 0.002019f 
C47025 a_11633_42308# VSS 0.006177f 
C47026 a_10149_42308# VSS 0.003101f 
C47027 a_9885_42308# VSS 0.007915f 
C47028 a_15890_42674# VSS 0.180637f 
C47029 a_15959_42545# VSS 0.263128f 
C47030 a_15803_42450# VSS 0.566963f 
C47031 a_15764_42576# VSS 0.298494f 
C47032 a_15486_42560# VSS 0.263746f 
C47033 a_15051_42282# VSS 0.790649f 
C47034 a_14113_42308# VSS 1.42448f 
C47035 a_13657_42558# VSS 0.00274f 
C47036 a_13249_42558# VSS 7.16e-20 
C47037 a_14456_42282# VSS 0.33927f 
C47038 a_13575_42558# VSS 0.370369f 
C47039 a_13070_42354# VSS 0.222095f 
C47040 a_12563_42308# VSS 0.330976f 
C47041 a_11633_42558# VSS 0.002749f 
C47042 a_11551_42558# VSS 0.372919f 
C47043 a_5742_30871# VSS 8.193179f 
C47044 a_11323_42473# VSS 0.253445f 
C47045 a_10723_42308# VSS 0.342975f 
C47046 a_10533_42308# VSS 0.310658f 
C47047 a_9885_42558# VSS 0.00274f 
C47048 a_9377_42558# VSS 7.16e-20 
C47049 a_9803_42558# VSS 0.370474f 
C47050 a_9223_42460# VSS 0.236204f 
C47051 a_8791_42308# VSS 0.301f 
C47052 a_8685_42308# VSS 0.163732f 
C47053 a_8325_42308# VSS 0.316205f 
C47054 a_4169_42308# VSS 0.00288f 
C47055 a_3905_42308# VSS 0.007531f 
C47056 a_8515_42308# VSS 0.250762f 
C47057 a_5934_30871# VSS 5.17381f 
C47058 a_7963_42308# VSS 0.256292f 
C47059 a_6123_31319# VSS 5.0238f 
C47060 a_7227_42308# VSS 0.359705f 
C47061 a_6761_42308# VSS 0.447596f 
C47062 a_5932_42308# VSS 5.11915f 
C47063 a_6171_42473# VSS 0.257988f 
C47064 a_5755_42308# VSS 0.314735f 
C47065 a_5421_42558# VSS 7.16e-20 
C47066 a_4921_42308# VSS 0.511258f 
C47067 a_3905_42558# VSS 0.00274f 
C47068 a_3497_42558# VSS 7.16e-20 
C47069 a_5379_42460# VSS 0.564806f 
C47070 a_5267_42460# VSS 0.204309f 
C47071 a_3823_42558# VSS 0.381485f 
C47072 a_3318_42354# VSS 0.238394f 
C47073 a_2903_42308# VSS 0.340659f 
C47074 a_2713_42308# VSS 0.31991f 
C47075 a_n39_42308# VSS 0.006513f 
C47076 a_n327_42308# VSS 0.002036f 
C47077 a_2351_42308# VSS 0.210162f 
C47078 a_2123_42473# VSS 0.21778f 
C47079 a_1755_42282# VSS 3.17706f 
C47080 a_1606_42308# VSS 5.25438f 
C47081 a_1149_42558# VSS 5.47e-35 
C47082 a_961_42354# VSS 0.215753f 
C47083 a_1184_42692# VSS 0.222827f 
C47084 a_1576_42282# VSS 0.327109f 
C47085 a_1067_42314# VSS 0.32917f 
C47086 a_n1630_35242# VSS 10.134f 
C47087 a_564_42282# VSS 0.36802f 
C47088 a_n3674_37592# VSS 3.04613f 
C47089 a_n327_42558# VSS 0.00274f 
C47090 a_n784_42308# VSS 6.50095f 
C47091 a_196_42282# VSS 0.343186f 
C47092 a_n473_42460# VSS 0.366068f 
C47093 a_n961_42308# VSS 0.328065f 
C47094 a_n1329_42308# VSS 0.30898f 
C47095 COMP_P VSS 11.0245f 
C47096 a_n4318_37592# VSS 1.00428f 
C47097 a_n1736_42282# VSS 0.320711f 
C47098 a_n3674_38216# VSS 1.68571f 
C47099 a_n2104_42282# VSS 0.346472f 
C47100 a_n4318_38216# VSS 0.964502f 
C47101 a_n2472_42282# VSS 0.335792f 
C47102 a_n3674_38680# VSS 0.881032f 
C47103 a_n2840_42282# VSS 0.343361f 
C47104 a_20753_42852# VSS 0.004913f 
C47105 a_20256_42852# VSS 1.31e-19 
C47106 a_14097_32519# VSS 1.90783f 
C47107 a_22400_42852# VSS 2.02868f 
C47108 a_20836_43172# VSS 0.003225f 
C47109 a_20573_43172# VSS 6.53e-19 
C47110 a_20256_43172# VSS 0.192089f 
C47111 a_18707_42852# VSS 0.004694f 
C47112 a_19518_43218# VSS 0.001266f 
C47113 a_19273_43230# VSS 4.65e-19 
C47114 a_18861_43218# VSS 0.00579f 
C47115 a_17749_42852# VSS 7.16e-20 
C47116 a_16877_42852# VSS 0.00274f 
C47117 a_16245_42852# VSS 0.004647f 
C47118 a_15597_42852# VSS 0.001372f 
C47119 a_18695_43230# VSS 0.008634f 
C47120 a_18504_43218# VSS 0.078212f 
C47121 a_17141_43172# VSS 0.002263f 
C47122 a_16877_43172# VSS 0.007531f 
C47123 a_16328_43172# VSS 0.003574f 
C47124 a_15785_43172# VSS 0.004243f 
C47125 a_14635_42282# VSS 0.336817f 
C47126 a_13291_42460# VSS 0.197331f 
C47127 a_13003_42852# VSS 0.004694f 
C47128 a_13814_43218# VSS 0.001281f 
C47129 a_13569_43230# VSS 4.65e-19 
C47130 a_11136_42852# VSS 0.004694f 
C47131 a_13157_43218# VSS 0.004992f 
C47132 a_12991_43230# VSS 0.006939f 
C47133 a_12800_43218# VSS 0.073862f 
C47134 a_11554_42852# VSS 0.073028f 
C47135 a_11301_43218# VSS 0.006939f 
C47136 a_11229_43218# VSS 0.004992f 
C47137 a_10793_43218# VSS 4.65e-19 
C47138 a_10553_43218# VSS 0.001281f 
C47139 a_8495_42852# VSS 0.004694f 
C47140 a_9306_43218# VSS 0.001281f 
C47141 a_9061_43230# VSS 4.65e-19 
C47142 a_8649_43218# VSS 0.004992f 
C47143 a_7309_42852# VSS 0.003102f 
C47144 a_5837_42852# VSS 0.00274f 
C47145 a_5193_42852# VSS 0.00274f 
C47146 a_4649_42852# VSS 0.006211f 
C47147 a_3863_42891# VSS 2.7e-19 
C47148 a_8483_43230# VSS 0.006939f 
C47149 a_8292_43218# VSS 0.073862f 
C47150 a_7573_43172# VSS 0.002122f 
C47151 a_7309_43172# VSS 0.006207f 
C47152 a_6101_43172# VSS 0.00288f 
C47153 a_5837_43172# VSS 0.005926f 
C47154 a_5457_43172# VSS 0.002122f 
C47155 a_5193_43172# VSS 0.005926f 
C47156 a_4743_43172# VSS 0.005048f 
C47157 a_4649_43172# VSS 0.005607f 
C47158 a_1793_42852# VSS 1.13e-19 
C47159 a_1709_42852# VSS 9.12e-20 
C47160 a_873_42968# VSS 6.57e-20 
C47161 a_133_42852# VSS 0.003564f 
C47162 a_4156_43218# VSS 0.003279f 
C47163 a_3935_43218# VSS 0.002898f 
C47164 a_3445_43172# VSS 0.001905f 
C47165 a_n2293_42282# VSS 2.62914f 
C47166 a_22959_42860# VSS 0.34332f 
C47167 a_22223_42860# VSS 0.328988f 
C47168 a_22165_42308# VSS 0.354098f 
C47169 a_21671_42860# VSS 0.316857f 
C47170 a_21195_42852# VSS 0.277519f 
C47171 a_21356_42826# VSS 0.304166f 
C47172 a_20922_43172# VSS 0.266814f 
C47173 a_19987_42826# VSS 0.378798f 
C47174 a_19164_43230# VSS 0.264863f 
C47175 a_19339_43156# VSS 0.471496f 
C47176 a_18599_43230# VSS 0.266382f 
C47177 a_18817_42826# VSS 0.182139f 
C47178 a_18249_42858# VSS 0.302863f 
C47179 a_17333_42852# VSS 0.29982f 
C47180 a_18083_42858# VSS 0.578693f 
C47181 a_17701_42308# VSS 0.179963f 
C47182 a_17595_43084# VSS 0.205109f 
C47183 a_16795_42852# VSS 0.362281f 
C47184 a_16414_43172# VSS 0.270304f 
C47185 a_15567_42826# VSS 0.316627f 
C47186 a_5342_30871# VSS 4.18054f 
C47187 a_15279_43071# VSS 0.248252f 
C47188 a_5534_30871# VSS 4.58413f 
C47189 a_14543_43071# VSS 0.246071f 
C47190 a_13460_43230# VSS 0.259861f 
C47191 a_13635_43156# VSS 0.7696f 
C47192 a_12895_43230# VSS 0.250159f 
C47193 a_13113_42826# VSS 0.174096f 
C47194 a_12545_42858# VSS 0.287468f 
C47195 a_12089_42308# VSS 0.283874f 
C47196 a_12379_42858# VSS 0.549229f 
C47197 a_10341_42308# VSS 0.317389f 
C47198 a_10922_42852# VSS 0.176112f 
C47199 a_10991_42826# VSS 0.261283f 
C47200 a_10796_42968# VSS 0.29877f 
C47201 a_10835_43094# VSS 0.59174f 
C47202 a_10518_42984# VSS 0.260322f 
C47203 a_10083_42826# VSS 0.762957f 
C47204 a_8952_43230# VSS 0.261046f 
C47205 a_9127_43156# VSS 0.77314f 
C47206 a_8387_43230# VSS 0.255573f 
C47207 a_8605_42826# VSS 0.181157f 
C47208 a_8037_42858# VSS 0.293593f 
C47209 a_7765_42852# VSS 0.252651f 
C47210 a_7871_42858# VSS 0.503534f 
C47211 a_7227_42852# VSS 0.36607f 
C47212 a_5755_42852# VSS 0.383967f 
C47213 a_5111_42852# VSS 0.354197f 
C47214 a_4520_42826# VSS 0.334784f 
C47215 a_3935_42891# VSS 0.26911f 
C47216 a_3681_42891# VSS 0.301094f 
C47217 a_2905_42968# VSS 0.305424f 
C47218 a_2075_43172# VSS 0.537699f 
C47219 a_1847_42826# VSS 0.670072f 
C47220 a_791_42968# VSS 0.335942f 
C47221 a_685_42968# VSS 0.220885f 
C47222 a_421_43172# VSS 0.006487f 
C47223 a_133_43172# VSS 0.00288f 
C47224 a_n1533_42852# VSS 0.004694f 
C47225 a_n722_43218# VSS 0.001281f 
C47226 a_n967_43230# VSS 4.65e-19 
C47227 a_n1379_43218# VSS 0.004992f 
C47228 a_n1545_43230# VSS 0.006939f 
C47229 a_n1736_43218# VSS 0.073862f 
C47230 a_n4318_38680# VSS 1.39087f 
C47231 a_n3674_39304# VSS 1.06639f 
C47232 a_n13_43084# VSS 0.368998f 
C47233 a_n1076_43230# VSS 0.263204f 
C47234 a_n901_43156# VSS 0.76245f 
C47235 a_n1641_43230# VSS 0.256397f 
C47236 a_n1423_42826# VSS 0.1805f 
C47237 a_n1991_42858# VSS 0.295941f 
C47238 a_n1853_43023# VSS 1.30078f 
C47239 a_n2157_42858# VSS 0.556569f 
C47240 a_n2472_42826# VSS 0.301801f 
C47241 a_n2840_42826# VSS 0.327636f 
C47242 a_20749_43396# VSS 0.253248f 
C47243 a_17364_32525# VSS 1.89349f 
C47244 a_22959_43396# VSS 0.345439f 
C47245 a_14209_32519# VSS 2.01016f 
C47246 a_22591_43396# VSS 0.335697f 
C47247 a_13887_32519# VSS 1.94312f 
C47248 a_22223_43396# VSS 0.333609f 
C47249 a_5649_42852# VSS 1.95364f 
C47250 a_13678_32519# VSS 2.06126f 
C47251 a_21855_43396# VSS 0.334538f 
C47252 a_4361_42308# VSS 1.30251f 
C47253 a_13467_32519# VSS 2.22551f 
C47254 a_19095_43396# VSS 0.132304f 
C47255 a_21487_43396# VSS 0.293844f 
C47256 a_20556_43646# VSS 0.006736f 
C47257 a_743_42282# VSS 1.36822f 
C47258 a_20301_43646# VSS 0.002477f 
C47259 a_4190_30871# VSS 7.37741f 
C47260 a_21259_43561# VSS 0.217667f 
C47261 a_17678_43396# VSS 0.001281f 
C47262 a_17433_43396# VSS 4.65e-19 
C47263 a_16823_43084# VSS 1.23251f 
C47264 a_17021_43396# VSS 0.004992f 
C47265 a_16855_43396# VSS 0.006939f 
C47266 a_15940_43402# VSS 0.003101f 
C47267 a_15868_43402# VSS 6.07e-19 
C47268 a_15231_43396# VSS 0.003851f 
C47269 a_15125_43396# VSS 0.003584f 
C47270 a_15037_43396# VSS 0.001503f 
C47271 a_16867_43762# VSS 0.004694f 
C47272 a_16664_43396# VSS 0.080001f 
C47273 a_19700_43370# VSS 0.335707f 
C47274 a_19268_43646# VSS 0.242693f 
C47275 a_15743_43084# VSS 1.49489f 
C47276 a_18783_43370# VSS 0.360096f 
C47277 a_18525_43370# VSS 0.361236f 
C47278 a_18429_43548# VSS 0.222219f 
C47279 a_17324_43396# VSS 0.258017f 
C47280 a_17499_43370# VSS 0.762886f 
C47281 a_16759_43396# VSS 0.252915f 
C47282 a_16977_43638# VSS 0.178776f 
C47283 a_16409_43396# VSS 0.290743f 
C47284 a_16547_43609# VSS 0.561468f 
C47285 a_16243_43396# VSS 0.562369f 
C47286 a_16137_43396# VSS 0.635905f 
C47287 a_13943_43396# VSS 0.003344f 
C47288 a_13837_43396# VSS 0.003427f 
C47289 a_13749_43396# VSS 0.001647f 
C47290 a_15781_43660# VSS 0.234761f 
C47291 a_15681_43442# VSS 0.20154f 
C47292 a_14537_43646# VSS 7.16e-20 
C47293 a_10149_43396# VSS 0.003443f 
C47294 a_9885_43396# VSS 0.006177f 
C47295 a_8945_43396# VSS 0.002098f 
C47296 a_8873_43396# VSS 0.001365f 
C47297 a_12281_43396# VSS 0.691406f 
C47298 a_10849_43646# VSS 7.16e-20 
C47299 a_10341_43396# VSS 0.796012f 
C47300 a_9885_43646# VSS 0.00274f 
C47301 a_14955_43396# VSS 0.266041f 
C47302 a_15095_43370# VSS 0.436411f 
C47303 a_14205_43396# VSS 0.2933f 
C47304 a_14358_43442# VSS 0.198188f 
C47305 a_14579_43548# VSS 0.293668f 
C47306 a_13667_43396# VSS 0.265557f 
C47307 a_10695_43548# VSS 0.279385f 
C47308 a_9803_43646# VSS 0.371929f 
C47309 a_9145_43396# VSS 0.437647f 
C47310 a_8423_43396# VSS 0.003573f 
C47311 a_8317_43396# VSS 0.003562f 
C47312 a_8229_43396# VSS 0.002303f 
C47313 a_7466_43396# VSS 0.001281f 
C47314 a_7221_43396# VSS 4.65e-19 
C47315 a_8685_43396# VSS 1.0146f 
C47316 a_6809_43396# VSS 0.004992f 
C47317 a_6643_43396# VSS 0.006939f 
C47318 a_5837_43396# VSS 0.001678f 
C47319 a_5565_43396# VSS 0.00164f 
C47320 a_4181_43396# VSS 0.001635f 
C47321 a_3457_43396# VSS 0.379621f 
C47322 a_2813_43396# VSS 0.412407f 
C47323 a_2437_43396# VSS 0.001678f 
C47324 a_6655_43762# VSS 0.004694f 
C47325 a_6452_43396# VSS 0.073862f 
C47326 a_9396_43370# VSS 0.338475f 
C47327 a_8791_43396# VSS 0.235222f 
C47328 a_8147_43396# VSS 0.256103f 
C47329 a_7112_43396# VSS 0.256956f 
C47330 a_7287_43370# VSS 0.754599f 
C47331 a_6547_43396# VSS 0.253718f 
C47332 a_6765_43638# VSS 0.174622f 
C47333 a_6197_43396# VSS 0.290517f 
C47334 a_6293_42852# VSS 0.473619f 
C47335 a_6031_43396# VSS 0.541083f 
C47336 a_1512_43396# VSS 0.003304f 
C47337 a_648_43396# VSS 0.231254f 
C47338 a_548_43396# VSS 0.009033f 
C47339 a_n144_43396# VSS 0.003264f 
C47340 a_n998_43396# VSS 0.001266f 
C47341 a_n1243_43396# VSS 4.65e-19 
C47342 a_3539_42460# VSS 0.337918f 
C47343 a_3626_43646# VSS 1.9807f 
C47344 a_3540_43646# VSS 9.9e-19 
C47345 a_2982_43646# VSS 3.25953f 
C47346 a_2896_43646# VSS 0.00155f 
C47347 a_1987_43646# VSS 6.34e-20 
C47348 a_1891_43646# VSS 1.35e-19 
C47349 a_1427_43646# VSS 0.00568f 
C47350 a_n1557_42282# VSS 0.870257f 
C47351 a_766_43646# VSS 9.92e-19 
C47352 a_4905_42826# VSS 0.781685f 
C47353 a_3080_42308# VSS 5.07176f 
C47354 a_4699_43561# VSS 0.267684f 
C47355 a_4235_43370# VSS 0.33553f 
C47356 a_4093_43548# VSS 0.320586f 
C47357 a_1756_43548# VSS 0.322408f 
C47358 a_1568_43370# VSS 0.63594f 
C47359 a_1049_43396# VSS 0.216408f 
C47360 a_1209_43370# VSS 0.281234f 
C47361 a_458_43396# VSS 0.252302f 
C47362 a_n229_43646# VSS 0.004647f 
C47363 a_n1655_43396# VSS 0.004992f 
C47364 a_n1821_43396# VSS 0.006939f 
C47365 a_n1809_43762# VSS 0.004697f 
C47366 a_n2012_43396# VSS 0.073862f 
C47367 a_104_43370# VSS 0.297328f 
C47368 a_n97_42460# VSS 6.9914f 
C47369 a_n447_43370# VSS 0.269574f 
C47370 a_n1352_43396# VSS 0.260107f 
C47371 a_n1177_43370# VSS 0.478516f 
C47372 a_n1917_43396# VSS 0.258245f 
C47373 a_n1699_43638# VSS 0.175452f 
C47374 a_n2267_43396# VSS 0.297246f 
C47375 a_n2129_43609# VSS 1.07965f 
C47376 a_n2433_43396# VSS 0.56533f 
C47377 a_n4318_39304# VSS 0.959585f 
C47378 a_n2840_43370# VSS 0.316787f 
C47379 a_17538_32519# VSS 1.8877f 
C47380 a_20974_43370# VSS 0.458091f 
C47381 a_14401_32519# VSS 2.32323f 
C47382 a_21381_43940# VSS 0.358332f 
C47383 a_19741_43940# VSS 0.007693f 
C47384 a_21205_44306# VSS 0.004143f 
C47385 a_18533_43940# VSS 0.00274f 
C47386 a_19319_43548# VSS 0.229395f 
C47387 a_19808_44306# VSS 0.005362f 
C47388 a_18797_44260# VSS 0.002999f 
C47389 a_18533_44260# VSS 0.007531f 
C47390 a_15037_43940# VSS 0.00274f 
C47391 a_13565_43940# VSS 0.00274f 
C47392 a_9801_43940# VSS 0.006211f 
C47393 a_9165_43940# VSS 0.001166f 
C47394 a_7499_43940# VSS 0.004678f 
C47395 a_6671_43940# VSS 0.004647f 
C47396 a_5829_43940# VSS 0.001102f 
C47397 a_5745_43940# VSS 7.11e-19 
C47398 a_5326_44056# VSS 9.13e-22 
C47399 a_3737_43940# VSS 0.001166f 
C47400 a_3052_44056# VSS 9.13e-22 
C47401 a_2455_43940# VSS 7.44e-19 
C47402 a_2253_43940# VSS 0.001314f 
C47403 a_1443_43940# VSS 8.96e-19 
C47404 a_1241_43940# VSS 0.001786f 
C47405 a_726_44056# VSS 4.62e-19 
C47406 a_15301_44260# VSS 0.00288f 
C47407 a_15037_44260# VSS 0.006076f 
C47408 a_14761_44260# VSS 0.001738f 
C47409 a_14485_44260# VSS 0.001738f 
C47410 a_14021_43940# VSS 0.387813f 
C47411 a_13829_44260# VSS 0.003443f 
C47412 a_13565_44260# VSS 0.005972f 
C47413 a_12710_44260# VSS 0.003489f 
C47414 a_12603_44260# VSS 0.004224f 
C47415 a_12495_44260# VSS 0.003836f 
C47416 a_11816_44260# VSS 0.00475f 
C47417 a_11173_44260# VSS 0.219946f 
C47418 a_10555_44260# VSS 0.346315f 
C47419 a_9895_44260# VSS 0.0063f 
C47420 a_9801_44260# VSS 0.006656f 
C47421 a_9248_44260# VSS 0.003866f 
C47422 a_22959_43948# VSS 0.341565f 
C47423 a_15493_43940# VSS 0.460801f 
C47424 a_22223_43948# VSS 0.31992f 
C47425 a_11341_43940# VSS 0.365183f 
C47426 a_21115_43940# VSS 0.204633f 
C47427 a_20935_43940# VSS 0.222887f 
C47428 a_20623_43914# VSS 0.371294f 
C47429 a_20365_43914# VSS 0.359455f 
C47430 a_20269_44172# VSS 0.225063f 
C47431 a_19862_44208# VSS 0.562087f 
C47432 a_19478_44306# VSS 0.278384f 
C47433 a_15493_43396# VSS 0.277875f 
C47434 a_19328_44172# VSS 0.2031f 
C47435 a_18451_43940# VSS 0.377396f 
C47436 a_18326_43940# VSS 0.276559f 
C47437 a_18079_43940# VSS 0.21121f 
C47438 a_17973_43940# VSS 0.359917f 
C47439 a_17737_43940# VSS 0.386318f 
C47440 a_15682_43940# VSS 1.9643f 
C47441 a_14955_43940# VSS 0.365393f 
C47442 a_13483_43940# VSS 0.376442f 
C47443 a_12429_44172# VSS 0.389129f 
C47444 a_11750_44172# VSS 0.221782f 
C47445 a_10807_43548# VSS 0.451031f 
C47446 a_10949_43914# VSS 0.257331f 
C47447 a_10729_43914# VSS 0.34307f 
C47448 a_10405_44172# VSS 0.142993f 
C47449 a_9672_43914# VSS 0.323006f 
C47450 a_9028_43914# VSS 0.398016f 
C47451 a_8333_44056# VSS 0.331632f 
C47452 a_8018_44260# VSS 0.005204f 
C47453 a_7911_44260# VSS 0.006364f 
C47454 a_7584_44260# VSS 0.003279f 
C47455 a_6756_44260# VSS 0.003243f 
C47456 a_n2661_42282# VSS 1.51789f 
C47457 a_6101_44260# VSS 0.001611f 
C47458 a_5841_44260# VSS 0.001326f 
C47459 a_3820_44260# VSS 0.004263f 
C47460 a_3499_42826# VSS 0.380221f 
C47461 a_2537_44260# VSS 0.001558f 
C47462 a_2253_44260# VSS 0.002472f 
C47463 a_1525_44260# VSS 0.001638f 
C47464 a_1241_44260# VSS 0.001824f 
C47465 a_261_44278# VSS 0.003386f 
C47466 a_n1441_43940# VSS 0.004694f 
C47467 a_n630_44306# VSS 0.002229f 
C47468 a_n875_44318# VSS 9.68e-19 
C47469 a_n1287_44306# VSS 0.00579f 
C47470 a_n1453_44318# VSS 0.008634f 
C47471 a_n1644_44306# VSS 0.080042f 
C47472 a_n3674_39768# VSS 0.890487f 
C47473 a_n4318_39768# VSS 1.09976f 
C47474 a_7845_44172# VSS 0.239173f 
C47475 a_7542_44172# VSS 0.283767f 
C47476 a_7281_43914# VSS 0.271121f 
C47477 a_6453_43914# VSS 0.26639f 
C47478 a_5663_43940# VSS 0.488325f 
C47479 a_5495_43940# VSS 0.212229f 
C47480 a_5013_44260# VSS 0.279924f 
C47481 a_5244_44056# VSS 0.216368f 
C47482 a_3905_42865# VSS 0.9893f 
C47483 a_3600_43914# VSS 0.422049f 
C47484 a_2998_44172# VSS 0.503048f 
C47485 a_2889_44172# VSS 0.217034f 
C47486 a_2675_43914# VSS 0.2974f 
C47487 a_895_43940# VSS 0.237723f 
C47488 a_2479_44172# VSS 0.817462f 
C47489 a_2127_44172# VSS 0.517911f 
C47490 a_453_43940# VSS 0.285192f 
C47491 a_1414_42308# VSS 1.07452f 
C47492 a_1467_44172# VSS 0.187431f 
C47493 a_1115_44172# VSS 0.52592f 
C47494 a_644_44056# VSS 0.227493f 
C47495 a_175_44278# VSS 0.226801f 
C47496 a_n984_44318# VSS 0.27358f 
C47497 a_n809_44244# VSS 0.785904f 
C47498 a_n1549_44318# VSS 0.264547f 
C47499 a_n1331_43914# VSS 0.185087f 
C47500 a_n1899_43946# VSS 0.299008f 
C47501 a_n1761_44111# VSS 0.392075f 
C47502 a_n2065_43946# VSS 0.658803f 
C47503 a_n2472_43914# VSS 0.3103f 
C47504 a_n2840_43914# VSS 0.345355f 
C47505 a_19237_31679# VSS 1.48755f 
C47506 a_22959_44484# VSS 0.343897f 
C47507 a_17730_32519# VSS 2.45301f 
C47508 a_22591_44484# VSS 0.315361f 
C47509 a_22485_44484# VSS 0.590119f 
C47510 a_20512_43084# VSS 0.561552f 
C47511 a_21145_44484# VSS 0.006939f 
C47512 a_21073_44484# VSS 0.004992f 
C47513 a_20637_44484# VSS 4.65e-19 
C47514 a_20397_44484# VSS 0.001266f 
C47515 a_22315_44484# VSS 0.238239f 
C47516 a_3422_30871# VSS 9.01786f 
C47517 a_21398_44850# VSS 0.073862f 
C47518 a_20980_44850# VSS 0.004694f 
C47519 a_19789_44512# VSS 0.003386f 
C47520 a_18753_44484# VSS 0.006939f 
C47521 a_18681_44484# VSS 0.004992f 
C47522 a_18579_44172# VSS 0.812679f 
C47523 a_18245_44484# VSS 4.65e-19 
C47524 a_18005_44484# VSS 0.001266f 
C47525 a_19279_43940# VSS 1.69633f 
C47526 a_20766_44850# VSS 0.177656f 
C47527 a_20835_44721# VSS 0.260406f 
C47528 a_20679_44626# VSS 0.58931f 
C47529 a_20640_44752# VSS 0.296084f 
C47530 a_20362_44736# VSS 0.255907f 
C47531 a_20159_44458# VSS 0.483669f 
C47532 a_19615_44636# VSS 0.238459f 
C47533 a_11967_42832# VSS 6.11191f 
C47534 a_19006_44850# VSS 0.073862f 
C47535 a_18588_44850# VSS 0.004694f 
C47536 a_17325_44484# VSS 0.002122f 
C47537 a_17061_44484# VSS 0.006177f 
C47538 a_16789_44484# VSS 0.002002f 
C47539 a_16335_44484# VSS 0.005048f 
C47540 a_16241_44484# VSS 0.005441f 
C47541 a_15367_44484# VSS 0.002898f 
C47542 a_15146_44484# VSS 0.002399f 
C47543 a_17517_44484# VSS 0.244051f 
C47544 a_17061_44734# VSS 0.00274f 
C47545 a_16241_44734# VSS 0.006211f 
C47546 a_14673_44172# VSS 0.290001f 
C47547 a_14581_44484# VSS 0.001661f 
C47548 a_13940_44484# VSS 0.004195f 
C47549 a_13296_44484# VSS 0.005047f 
C47550 a_12829_44484# VSS 0.001944f 
C47551 a_12553_44484# VSS 0.00193f 
C47552 a_12189_44484# VSS 0.001627f 
C47553 a_11909_44484# VSS 0.001659f 
C47554 a_11541_44484# VSS 0.139071f 
C47555 a_10809_44484# VSS 0.001938f 
C47556 a_15463_44811# VSS 2.7e-19 
C47557 a_15433_44458# VSS 0.301508f 
C47558 a_14815_43914# VSS 0.445698f 
C47559 a_13857_44734# VSS 0.001166f 
C47560 a_13213_44734# VSS 0.001208f 
C47561 a_n2293_43922# VSS 3.31971f 
C47562 a_n2661_43922# VSS 1.51991f 
C47563 a_n2661_42834# VSS 1.20196f 
C47564 a_9159_44484# VSS 0.158168f 
C47565 a_10617_44484# VSS 0.119149f 
C47566 a_5708_44484# VSS 0.231649f 
C47567 a_5608_44484# VSS 0.007818f 
C47568 a_3363_44484# VSS 0.27629f 
C47569 a_556_44484# VSS 0.201935f 
C47570 a_484_44484# VSS 0.004815f 
C47571 a_n89_44484# VSS 0.002857f 
C47572 a_n310_44484# VSS 0.002596f 
C47573 a_9313_44734# VSS 1.31461f 
C47574 a_5891_43370# VSS 2.82295f 
C47575 a_8375_44464# VSS 0.211867f 
C47576 a_7640_43914# VSS 0.542377f 
C47577 a_6109_44484# VSS 0.648821f 
C47578 a_700_44734# VSS 0.001076f 
C47579 a_n998_44484# VSS 0.002215f 
C47580 a_n1243_44484# VSS 9.68e-19 
C47581 a_7_44811# VSS 2.7e-19 
C47582 a_n23_44458# VSS 0.278255f 
C47583 a_n356_44636# VSS 2.91333f 
C47584 a_n1655_44484# VSS 0.00579f 
C47585 a_n1821_44484# VSS 0.008634f 
C47586 a_n1809_44850# VSS 0.007269f 
C47587 a_n2012_44484# VSS 0.080001f 
C47588 a_18989_43940# VSS 0.423174f 
C47589 a_18374_44850# VSS 0.179731f 
C47590 a_18443_44721# VSS 0.253971f 
C47591 a_18287_44626# VSS 0.507939f 
C47592 a_18248_44752# VSS 0.294917f 
C47593 a_17970_44736# VSS 0.26161f 
C47594 a_17767_44458# VSS 0.474097f 
C47595 a_16979_44734# VSS 0.363013f 
C47596 a_14539_43914# VSS 1.18088f 
C47597 a_16112_44458# VSS 0.326339f 
C47598 a_15004_44636# VSS 0.254778f 
C47599 a_13720_44458# VSS 0.403209f 
C47600 a_13076_44458# VSS 0.38829f 
C47601 a_12883_44458# VSS 0.287544f 
C47602 a_12607_44458# VSS 0.499331f 
C47603 a_8975_43940# VSS 0.652857f 
C47604 a_10057_43914# VSS 0.654189f 
C47605 a_10440_44484# VSS 0.210149f 
C47606 a_10334_44484# VSS 0.210217f 
C47607 a_10157_44484# VSS 0.208916f 
C47608 a_9838_44484# VSS 0.276258f 
C47609 a_5883_43914# VSS 0.792825f 
C47610 a_8701_44490# VSS 0.358059f 
C47611 a_8103_44636# VSS 0.340824f 
C47612 a_6298_44484# VSS 1.93814f 
C47613 a_5518_44484# VSS 0.242995f 
C47614 a_5343_44458# VSS 1.28071f 
C47615 a_4743_44484# VSS 0.327178f 
C47616 a_n699_43396# VSS 1.82142f 
C47617 a_4223_44672# VSS 0.659279f 
C47618 a_2779_44458# VSS 0.532137f 
C47619 a_949_44458# VSS 1.97734f 
C47620 a_742_44458# VSS 1.02263f 
C47621 a_n452_44636# VSS 0.254732f 
C47622 a_n1352_44484# VSS 0.269853f 
C47623 a_n1177_44458# VSS 0.493891f 
C47624 a_n1917_44484# VSS 0.280038f 
C47625 a_n1699_44726# VSS 0.197478f 
C47626 a_n2267_44484# VSS 0.308908f 
C47627 a_n2129_44697# VSS 0.307327f 
C47628 a_n2433_44484# VSS 0.679598f 
C47629 a_n2661_44458# VSS 0.487677f 
C47630 a_n4318_40392# VSS 0.995833f 
C47631 a_n2840_44458# VSS 0.316322f 
C47632 a_19721_31679# VSS 1.61485f 
C47633 a_18114_32519# VSS 3.10957f 
C47634 a_17801_45144# VSS 8.35e-20 
C47635 a_16237_45028# VSS 0.017944f 
C47636 a_20193_45348# VSS 1.70015f 
C47637 a_11691_44458# VSS 1.78467f 
C47638 a_19113_45348# VSS 0.367248f 
C47639 a_22959_45036# VSS 0.345334f 
C47640 a_22223_45036# VSS 0.354178f 
C47641 a_11827_44484# VSS 1.28091f 
C47642 a_21359_45002# VSS 0.397791f 
C47643 a_21101_45002# VSS 0.35202f 
C47644 a_21005_45260# VSS 0.212992f 
C47645 a_20567_45036# VSS 0.31908f 
C47646 a_18494_42460# VSS 1.15626f 
C47647 a_18184_42460# VSS 0.838573f 
C47648 a_19778_44110# VSS 0.599421f 
C47649 a_18911_45144# VSS 0.307008f 
C47650 a_18587_45118# VSS 0.214925f 
C47651 a_18315_45260# VSS 0.334834f 
C47652 a_17719_45144# VSS 0.331229f 
C47653 a_17613_45144# VSS 0.244364f 
C47654 a_17023_45118# VSS 0.20885f 
C47655 a_16922_45042# VSS 0.818675f 
C47656 a_16501_45348# VSS 0.005461f 
C47657 a_16405_45348# VSS 0.003038f 
C47658 a_16321_45348# VSS 0.002956f 
C47659 a_14309_45028# VSS 0.006587f 
C47660 a_13807_45067# VSS 2.7e-19 
C47661 a_15685_45394# VSS 0.003883f 
C47662 a_15060_45348# VSS 0.006388f 
C47663 a_14976_45348# VSS 0.005191f 
C47664 a_14403_45348# VSS 0.006612f 
C47665 a_14309_45348# VSS 0.006958f 
C47666 a_13711_45394# VSS 0.002898f 
C47667 a_13490_45394# VSS 0.002596f 
C47668 a_13105_45348# VSS 0.001738f 
C47669 a_11915_45394# VSS 0.004143f 
C47670 a_n2661_43370# VSS 0.820606f 
C47671 a_11361_45348# VSS 0.001666f 
C47672 a_7735_45067# VSS 2.7e-19 
C47673 a_10903_45394# VSS 0.004143f 
C47674 a_8560_45348# VSS 0.185033f 
C47675 a_8488_45348# VSS 0.003218f 
C47676 a_8137_45348# VSS 0.001684f 
C47677 a_n2293_42834# VSS 1.1151f 
C47678 a_7639_45394# VSS 0.002898f 
C47679 a_7418_45394# VSS 0.002596f 
C47680 a_6945_45348# VSS 0.001738f 
C47681 a_5837_45028# VSS 0.00274f 
C47682 a_5093_45028# VSS 0.001102f 
C47683 a_5009_45028# VSS 7.39e-19 
C47684 a_2809_45028# VSS 0.00638f 
C47685 a_2448_45028# VSS 1.19e-20 
C47686 a_6517_45366# VSS 0.003386f 
C47687 a_6125_45348# VSS 0.007531f 
C47688 a_5837_45348# VSS 0.002999f 
C47689 a_5365_45348# VSS 0.002387f 
C47690 a_5105_45348# VSS 0.001558f 
C47691 a_4640_45348# VSS 0.006141f 
C47692 a_4185_45348# VSS 0.001865f 
C47693 a_3602_45348# VSS 0.005184f 
C47694 a_3495_45348# VSS 0.006372f 
C47695 a_2903_45348# VSS 0.005166f 
C47696 a_2809_45348# VSS 0.006958f 
C47697 a_2304_45348# VSS 0.182367f 
C47698 a_2232_45348# VSS 0.004649f 
C47699 a_1423_45028# VSS 0.980773f 
C47700 a_1145_45348# VSS 0.001816f 
C47701 a_626_44172# VSS 0.67926f 
C47702 a_501_45348# VSS 0.001778f 
C47703 a_375_42282# VSS 0.447027f 
C47704 a_16751_45260# VSS 0.316547f 
C47705 a_1307_43914# VSS 2.30311f 
C47706 a_16019_45002# VSS 0.25377f 
C47707 a_15595_45028# VSS 0.214111f 
C47708 a_15415_45028# VSS 0.221991f 
C47709 a_14797_45144# VSS 0.249222f 
C47710 a_14537_43396# VSS 1.73146f 
C47711 a_14180_45002# VSS 0.327485f 
C47712 a_13777_45326# VSS 0.272936f 
C47713 a_13556_45296# VSS 1.01916f 
C47714 a_9482_43914# VSS 3.42654f 
C47715 a_13348_45260# VSS 0.243533f 
C47716 a_13159_45002# VSS 0.265737f 
C47717 a_13017_45260# VSS 0.362048f 
C47718 a_11963_45334# VSS 0.226884f 
C47719 a_11787_45002# VSS 0.212512f 
C47720 a_10951_45334# VSS 0.228638f 
C47721 a_10775_45002# VSS 0.204487f 
C47722 a_8953_45002# VSS 1.94941f 
C47723 a_8191_45002# VSS 0.325964f 
C47724 a_7705_45326# VSS 0.273009f 
C47725 a_6709_45028# VSS 0.354418f 
C47726 a_7229_43940# VSS 0.786182f 
C47727 a_7276_45260# VSS 0.251523f 
C47728 a_5205_44484# VSS 0.546179f 
C47729 a_6431_45366# VSS 0.233718f 
C47730 a_6171_45002# VSS 0.700605f 
C47731 a_3232_43370# VSS 2.99721f 
C47732 a_5691_45260# VSS 0.370273f 
C47733 a_4927_45028# VSS 0.520892f 
C47734 a_5111_44636# VSS 3.44603f 
C47735 a_5147_45002# VSS 0.803306f 
C47736 a_4558_45348# VSS 0.446148f 
C47737 a_4574_45260# VSS 0.208274f 
C47738 a_3537_45260# VSS 2.45782f 
C47739 a_3429_45260# VSS 0.274034f 
C47740 a_3065_45002# VSS 0.864786f 
C47741 a_2680_45002# VSS 0.321351f 
C47742 a_2382_45260# VSS 1.03422f 
C47743 a_2274_45254# VSS 0.187307f 
C47744 a_1667_45002# VSS 0.345429f 
C47745 a_327_44734# VSS 0.419171f 
C47746 a_413_45260# VSS 4.87522f 
C47747 a_n37_45144# VSS 0.321746f 
C47748 a_n143_45144# VSS 0.209896f 
C47749 a_n467_45028# VSS 0.311181f 
C47750 a_n659_45366# VSS 0.004685f 
C47751 a_n967_45348# VSS 0.453992f 
C47752 en_comp VSS 7.869411f 
C47753 a_n2956_37592# VSS 2.90302f 
C47754 a_n2810_45028# VSS 1.52635f 
C47755 a_n745_45366# VSS 0.257282f 
C47756 a_n913_45002# VSS 5.04726f 
C47757 a_n1059_45260# VSS 2.30619f 
C47758 a_n2017_45002# VSS 1.09013f 
C47759 a_n2109_45247# VSS 0.252392f 
C47760 a_n2293_45010# VSS 0.614925f 
C47761 a_n2472_45002# VSS 0.298945f 
C47762 a_n2661_45010# VSS 0.839496f 
C47763 a_n2840_45002# VSS 0.340687f 
C47764 a_21542_45572# VSS 0.002215f 
C47765 a_21297_45572# VSS 9.68e-19 
C47766 a_20447_31679# VSS 1.48786f 
C47767 a_22959_45572# VSS 0.34535f 
C47768 a_19963_31679# VSS 1.43433f 
C47769 a_22591_45572# VSS 0.363695f 
C47770 a_3357_43084# VSS 2.42707f 
C47771 a_19479_31679# VSS 1.66892f 
C47772 a_22223_45572# VSS 0.334964f 
C47773 a_2437_43646# VSS 6.25635f 
C47774 a_21513_45002# VSS 0.669089f 
C47775 a_20885_45572# VSS 0.004992f 
C47776 a_20719_45572# VSS 0.006939f 
C47777 a_19610_45572# VSS 0.002215f 
C47778 a_19365_45572# VSS 4.65e-19 
C47779 a_20731_45938# VSS 0.004694f 
C47780 a_20528_45572# VSS 0.073082f 
C47781 a_21188_45572# VSS 0.284872f 
C47782 a_21363_45546# VSS 0.515994f 
C47783 a_20623_45572# VSS 0.256236f 
C47784 a_20841_45814# VSS 0.180037f 
C47785 a_20273_45572# VSS 0.288513f 
C47786 a_20107_45572# VSS 0.541125f 
C47787 a_18953_45572# VSS 0.004992f 
C47788 a_18787_45572# VSS 0.006939f 
C47789 a_17668_45572# VSS 0.217142f 
C47790 a_17568_45572# VSS 0.005817f 
C47791 a_17034_45572# VSS 0.001266f 
C47792 a_16789_45572# VSS 4.65e-19 
C47793 a_18799_45938# VSS 0.004694f 
C47794 a_18596_45572# VSS 0.073862f 
C47795 a_19256_45572# VSS 0.257674f 
C47796 a_19431_45546# VSS 0.487121f 
C47797 a_18691_45572# VSS 0.255356f 
C47798 a_18909_45814# VSS 0.178658f 
C47799 a_18341_45572# VSS 0.291608f 
C47800 a_18479_45785# VSS 1.15946f 
C47801 a_18175_45572# VSS 0.516981f 
C47802 a_16147_45260# VSS 0.506229f 
C47803 a_16377_45572# VSS 0.004992f 
C47804 a_16211_45572# VSS 0.006939f 
C47805 a_14127_45572# VSS 0.006612f 
C47806 a_14033_45572# VSS 0.006958f 
C47807 a_13485_45572# VSS 0.001696f 
C47808 a_13385_45572# VSS 0.004208f 
C47809 a_13297_45572# VSS 0.004404f 
C47810 a_12749_45572# VSS 0.00153f 
C47811 a_12649_45572# VSS 0.005051f 
C47812 a_12561_45572# VSS 0.005505f 
C47813 a_16223_45938# VSS 0.004694f 
C47814 a_16020_45572# VSS 0.073862f 
C47815 a_17478_45572# VSS 0.232341f 
C47816 a_15861_45028# VSS 0.449058f 
C47817 a_8696_44636# VSS 0.917254f 
C47818 a_16680_45572# VSS 0.258674f 
C47819 a_16855_45546# VSS 0.471485f 
C47820 a_16115_45572# VSS 0.253972f 
C47821 a_16333_45814# VSS 0.178165f 
C47822 a_15765_45572# VSS 0.291326f 
C47823 a_15903_45785# VSS 0.4164f 
C47824 a_15599_45572# VSS 0.50233f 
C47825 a_15037_45618# VSS 0.209713f 
C47826 a_14033_45822# VSS 0.006541f 
C47827 a_12016_45572# VSS 0.005248f 
C47828 a_11778_45572# VSS 0.003039f 
C47829 a_11688_45572# VSS 0.002091f 
C47830 a_11136_45572# VSS 0.17156f 
C47831 a_11064_45572# VSS 0.003188f 
C47832 a_10544_45572# VSS 0.006484f 
C47833 a_10306_45572# VSS 0.004928f 
C47834 a_10216_45572# VSS 0.003935f 
C47835 a_9159_45572# VSS 0.151638f 
C47836 a_8791_45572# VSS 0.00583f 
C47837 a_8697_45572# VSS 0.005152f 
C47838 a_8192_45572# VSS 0.17002f 
C47839 a_8120_45572# VSS 0.004768f 
C47840 a_11682_45822# VSS 0.010374f 
C47841 a_10907_45822# VSS 0.547001f 
C47842 a_10210_45822# VSS 0.012573f 
C47843 a_8697_45822# VSS 0.006221f 
C47844 a_6977_45572# VSS 0.008634f 
C47845 a_6905_45572# VSS 0.00579f 
C47846 a_6469_45572# VSS 9.68e-19 
C47847 a_6229_45572# VSS 0.002215f 
C47848 a_15143_45578# VSS 0.315994f 
C47849 a_14495_45572# VSS 0.325874f 
C47850 a_13249_42308# VSS 1.08648f 
C47851 a_13904_45546# VSS 0.327907f 
C47852 a_13527_45546# VSS 0.245514f 
C47853 a_13163_45724# VSS 0.180841f 
C47854 a_12791_45546# VSS 0.237787f 
C47855 a_11823_42460# VSS 2.45644f 
C47856 a_12427_45724# VSS 0.190531f 
C47857 a_11962_45724# VSS 0.218739f 
C47858 a_11652_45724# VSS 0.258015f 
C47859 a_11525_45546# VSS 0.346102f 
C47860 a_11322_45546# VSS 0.62914f 
C47861 a_10490_45724# VSS 0.972668f 
C47862 a_8746_45002# VSS 0.547616f 
C47863 a_10193_42453# VSS 3.59848f 
C47864 a_10180_45724# VSS 0.281135f 
C47865 a_10053_45546# VSS 0.373668f 
C47866 a_9049_44484# VSS 0.249658f 
C47867 a_7499_43078# VSS 3.22587f 
C47868 a_8568_45546# VSS 0.317032f 
C47869 a_8162_45546# VSS 0.376225f 
C47870 a_7230_45938# VSS 0.078992f 
C47871 a_6812_45938# VSS 0.004694f 
C47872 a_5437_45600# VSS 0.004685f 
C47873 a_4880_45572# VSS 0.182839f 
C47874 a_4808_45572# VSS 0.004805f 
C47875 a_5024_45822# VSS 2.99e-19 
C47876 a_3260_45572# VSS 0.003272f 
C47877 a_2211_45572# VSS 0.002983f 
C47878 a_1990_45572# VSS 0.00263f 
C47879 a_3775_45552# VSS 0.209244f 
C47880 a_7227_45028# VSS 0.439395f 
C47881 a_6598_45938# VSS 0.185967f 
C47882 a_6667_45809# VSS 0.264656f 
C47883 a_6511_45714# VSS 0.647716f 
C47884 a_6472_45840# VSS 0.310105f 
C47885 a_6194_45824# VSS 0.2717f 
C47886 a_5907_45546# VSS 0.592148f 
C47887 a_5263_45724# VSS 0.250928f 
C47888 a_4099_45572# VSS 0.33915f 
C47889 a_3175_45822# VSS 0.004647f 
C47890 a_2711_45572# VSS 1.77517f 
C47891 a_1609_45572# VSS 0.001977f 
C47892 a_1260_45572# VSS 0.006784f 
C47893 a_1176_45572# VSS 0.005484f 
C47894 a_603_45572# VSS 0.008207f 
C47895 a_509_45572# VSS 0.005519f 
C47896 a_n89_45572# VSS 0.003313f 
C47897 a_n310_45572# VSS 0.002596f 
C47898 a_2307_45899# VSS 3.38e-19 
C47899 a_1990_45899# VSS 1.9e-19 
C47900 a_2277_45546# VSS 0.303704f 
C47901 a_1609_45822# VSS 0.5528f 
C47902 a_n443_42852# VSS 4.64762f 
C47903 a_509_45822# VSS 0.010571f 
C47904 a_n906_45572# VSS 0.006201f 
C47905 a_n1013_45572# VSS 0.008252f 
C47906 a_7_45899# VSS 2.7e-19 
C47907 a_n23_45546# VSS 0.281189f 
C47908 a_n356_45724# VSS 0.32306f 
C47909 a_3503_45724# VSS 0.322319f 
C47910 a_3316_45546# VSS 0.336134f 
C47911 a_3218_45724# VSS 0.379893f 
C47912 a_2957_45546# VSS 0.276358f 
C47913 a_1848_45724# VSS 0.245258f 
C47914 a_997_45618# VSS 0.248122f 
C47915 a_n755_45592# VSS 5.8889f 
C47916 a_n357_42282# VSS 2.46134f 
C47917 a_310_45028# VSS 0.207165f 
C47918 a_n1099_45572# VSS 0.339525f 
C47919 a_380_45546# VSS 0.337145f 
C47920 a_n452_45724# VSS 0.253614f 
C47921 a_n863_45724# VSS 3.49288f 
C47922 a_n1079_45724# VSS 0.289271f 
C47923 a_n2293_45546# VSS 0.879703f 
C47924 a_n2956_38216# VSS 1.49846f 
C47925 a_n2472_45546# VSS 0.340801f 
C47926 a_n2661_45546# VSS 1.58481f 
C47927 a_n2810_45572# VSS 1.43198f 
C47928 a_n2840_45546# VSS 0.344757f 
C47929 a_21167_46155# VSS 2.7e-19 
C47930 a_20692_30879# VSS 1.59585f 
C47931 a_20205_31679# VSS 1.45349f 
C47932 a_21071_46482# VSS 0.003313f 
C47933 a_20850_46482# VSS 0.003279f 
C47934 a_19443_46116# VSS 0.004694f 
C47935 a_20254_46482# VSS 0.001266f 
C47936 a_20009_46494# VSS 4.65e-19 
C47937 a_19597_46482# VSS 0.004992f 
C47938 a_18051_46116# VSS 0.006211f 
C47939 a_19431_46494# VSS 0.006939f 
C47940 a_19240_46482# VSS 0.073862f 
C47941 a_16375_45002# VSS 1.44161f 
C47942 a_18243_46436# VSS 0.005441f 
C47943 a_18147_46436# VSS 0.005048f 
C47944 a_13259_45724# VSS 4.49011f 
C47945 a_14383_46116# VSS 0.00471f 
C47946 a_15194_46482# VSS 0.001266f 
C47947 a_14949_46494# VSS 9.68e-19 
C47948 a_14537_46482# VSS 0.004992f 
C47949 a_12839_46116# VSS 0.001465f 
C47950 a_11315_46155# VSS 2.7e-19 
C47951 a_14371_46494# VSS 0.006939f 
C47952 a_14180_46482# VSS 0.073862f 
C47953 a_12638_46436# VSS 0.162178f 
C47954 a_12379_46436# VSS 0.275423f 
C47955 a_12005_46436# VSS 0.001661f 
C47956 a_9751_46155# VSS 2.7e-19 
C47957 a_11608_46482# VSS 0.003279f 
C47958 a_11387_46482# VSS 0.002827f 
C47959 a_10586_45546# VSS 0.542658f 
C47960 a_8379_46155# VSS 2.7e-19 
C47961 a_10044_46482# VSS 0.003279f 
C47962 a_9823_46482# VSS 0.002827f 
C47963 a_9241_46436# VSS 0.001883f 
C47964 a_8049_45260# VSS 0.741927f 
C47965 a_8781_46436# VSS 0.00189f 
C47966 a_6347_46155# VSS 2.7e-19 
C47967 a_8034_45724# VSS 0.299594f 
C47968 a_8283_46482# VSS 0.002857f 
C47969 a_8062_46482# VSS 0.003279f 
C47970 a_5527_46155# VSS 2.7e-19 
C47971 a_6640_46482# VSS 0.003279f 
C47972 a_6419_46482# VSS 0.003313f 
C47973 a_5066_45546# VSS 0.436834f 
C47974 a_5431_46482# VSS 0.003543f 
C47975 a_5210_46482# VSS 0.003279f 
C47976 a_4365_46436# VSS 0.001655f 
C47977 a_1337_46116# VSS 0.007537f 
C47978 a_835_46155# VSS 0.001095f 
C47979 a_518_46155# VSS 4.91e-19 
C47980 a_3873_46454# VSS 0.00338f 
C47981 a_n1925_42282# VSS 1.34109f 
C47982 a_526_44458# VSS 6.44493f 
C47983 a_2981_46116# VSS 0.091491f 
C47984 a_1431_46436# VSS 0.005311f 
C47985 a_1337_46436# VSS 0.005657f 
C47986 a_739_46482# VSS 0.004344f 
C47987 a_518_46482# VSS 0.003651f 
C47988 a_n1533_46116# VSS 0.006086f 
C47989 a_n722_46482# VSS 0.001281f 
C47990 a_n967_46494# VSS 4.65e-19 
C47991 a_n1379_46482# VSS 0.004992f 
C47992 a_n1545_46494# VSS 0.006939f 
C47993 a_n1736_46482# VSS 0.07565f 
C47994 a_n2956_38680# VSS 1.34225f 
C47995 a_n2956_39304# VSS 1.60721f 
C47996 a_22959_46124# VSS 0.345245f 
C47997 a_10809_44734# VSS 1.05002f 
C47998 a_22223_46124# VSS 0.354467f 
C47999 a_6945_45028# VSS 0.978274f 
C48000 a_21137_46414# VSS 0.340736f 
C48001 a_20708_46348# VSS 0.268156f 
C48002 a_19900_46494# VSS 0.26164f 
C48003 a_20075_46420# VSS 0.475201f 
C48004 a_19335_46494# VSS 0.260378f 
C48005 a_19553_46090# VSS 0.179968f 
C48006 a_18985_46122# VSS 0.297132f 
C48007 a_18819_46122# VSS 0.545109f 
C48008 a_17957_46116# VSS 0.309446f 
C48009 a_18189_46348# VSS 0.296366f 
C48010 a_17715_44484# VSS 0.55862f 
C48011 a_17583_46090# VSS 0.307562f 
C48012 a_15682_46116# VSS 1.96743f 
C48013 a_2324_44458# VSS 6.12227f 
C48014 a_14840_46494# VSS 0.263367f 
C48015 a_15015_46420# VSS 0.472948f 
C48016 a_14275_46494# VSS 0.258968f 
C48017 a_14493_46090# VSS 0.176122f 
C48018 a_13925_46122# VSS 0.294602f 
C48019 a_13759_46122# VSS 0.518292f 
C48020 a_13351_46090# VSS 0.304427f 
C48021 a_12594_46348# VSS 0.284494f 
C48022 a_12005_46116# VSS 0.381711f 
C48023 a_10903_43370# VSS 2.66576f 
C48024 a_11387_46155# VSS 0.260117f 
C48025 a_11133_46155# VSS 0.299642f 
C48026 a_11189_46129# VSS 0.32558f 
C48027 a_9290_44172# VSS 4.78398f 
C48028 a_10355_46116# VSS 0.290668f 
C48029 a_9823_46155# VSS 0.261206f 
C48030 a_9569_46155# VSS 0.304755f 
C48031 a_9625_46129# VSS 0.369694f 
C48032 a_8953_45546# VSS 1.00397f 
C48033 a_5937_45572# VSS 1.8333f 
C48034 a_8199_44636# VSS 2.29742f 
C48035 a_8349_46414# VSS 0.273442f 
C48036 a_8016_46348# VSS 0.539696f 
C48037 a_7920_46348# VSS 0.269852f 
C48038 a_6419_46155# VSS 0.273686f 
C48039 a_6165_46155# VSS 0.303989f 
C48040 a_5497_46414# VSS 0.304684f 
C48041 a_5204_45822# VSS 0.338817f 
C48042 a_5164_46348# VSS 0.419282f 
C48043 a_5068_46348# VSS 0.25855f 
C48044 a_4704_46090# VSS 0.296767f 
C48045 a_4419_46090# VSS 0.357571f 
C48046 a_4185_45028# VSS 2.50501f 
C48047 a_3699_46348# VSS 0.226584f 
C48048 a_3483_46348# VSS 4.80498f 
C48049 a_3147_46376# VSS 0.52775f 
C48050 a_2804_46116# VSS 0.222855f 
C48051 a_2698_46116# VSS 0.215567f 
C48052 a_2521_46116# VSS 0.220999f 
C48053 a_167_45260# VSS 1.32487f 
C48054 a_2202_46116# VSS 0.273578f 
C48055 a_1823_45246# VSS 2.36307f 
C48056 a_1138_42852# VSS 0.456566f 
C48057 a_1176_45822# VSS 0.278365f 
C48058 a_1208_46090# VSS 0.348206f 
C48059 a_805_46414# VSS 0.27506f 
C48060 a_472_46348# VSS 0.32751f 
C48061 a_376_46348# VSS 0.285607f 
C48062 a_n1076_46494# VSS 0.262147f 
C48063 a_n901_46420# VSS 0.762523f 
C48064 a_n1641_46494# VSS 0.256945f 
C48065 a_n1423_46090# VSS 0.176189f 
C48066 a_n1991_46122# VSS 0.305274f 
C48067 a_n1853_46287# VSS 0.341802f 
C48068 a_n2157_46122# VSS 0.525314f 
C48069 a_n2293_46098# VSS 0.690447f 
C48070 a_n2472_46090# VSS 0.290925f 
C48071 a_n2840_46090# VSS 0.340313f 
C48072 a_21542_46660# VSS 0.002215f 
C48073 a_21297_46660# VSS 9.68e-19 
C48074 a_21076_30879# VSS 2.00065f 
C48075 a_22959_46660# VSS 0.338967f 
C48076 a_12741_44636# VSS 0.979225f 
C48077 a_20820_30879# VSS 1.64286f 
C48078 a_22591_46660# VSS 0.292786f 
C48079 a_11415_45002# VSS 1.63684f 
C48080 a_20202_43084# VSS 1.05073f 
C48081 a_22365_46825# VSS 0.208388f 
C48082 a_20885_46660# VSS 0.004992f 
C48083 a_20719_46660# VSS 0.006939f 
C48084 a_19636_46660# VSS 0.003657f 
C48085 a_18900_46660# VSS 0.006141f 
C48086 a_18280_46660# VSS 0.29316f 
C48087 a_17639_46660# VSS 0.308795f 
C48088 a_16655_46660# VSS 0.003226f 
C48089 a_16434_46660# VSS 0.003279f 
C48090 a_20731_47026# VSS 0.004694f 
C48091 a_20528_46660# VSS 0.07565f 
C48092 a_22000_46634# VSS 0.295895f 
C48093 a_21188_46660# VSS 0.261124f 
C48094 a_21363_46634# VSS 0.488515f 
C48095 a_20623_46660# VSS 0.258464f 
C48096 a_20841_46902# VSS 0.180869f 
C48097 a_20273_46660# VSS 0.309206f 
C48098 a_20411_46873# VSS 0.393328f 
C48099 a_20107_46660# VSS 0.575208f 
C48100 a_19551_46910# VSS 0.005326f 
C48101 a_19123_46287# VSS 0.477642f 
C48102 a_18285_46348# VSS 0.577053f 
C48103 a_17829_46910# VSS 3.25e-20 
C48104 a_765_45546# VSS 0.902406f 
C48105 a_17339_46660# VSS 0.927636f 
C48106 a_15312_46660# VSS 0.003243f 
C48107 a_14447_46660# VSS 0.002898f 
C48108 a_14226_46660# VSS 0.002596f 
C48109 a_16751_46987# VSS 2.7e-19 
C48110 a_16721_46634# VSS 0.305539f 
C48111 a_16388_46812# VSS 1.42609f 
C48112 a_13059_46348# VSS 2.36107f 
C48113 a_15227_46910# VSS 0.004775f 
C48114 a_13693_46688# VSS 0.003947f 
C48115 a_14543_46987# VSS 2.7e-19 
C48116 a_14513_46634# VSS 0.29862f 
C48117 a_14180_46812# VSS 0.368158f 
C48118 a_14035_46660# VSS 0.322858f 
C48119 a_13885_46660# VSS 0.297377f 
C48120 a_13170_46660# VSS 0.001266f 
C48121 a_12925_46660# VSS 4.65e-19 
C48122 a_12513_46660# VSS 0.004992f 
C48123 a_12347_46660# VSS 0.006939f 
C48124 a_10933_46660# VSS 0.008634f 
C48125 a_10861_46660# VSS 0.00579f 
C48126 a_12359_47026# VSS 0.007095f 
C48127 a_12156_46660# VSS 0.074642f 
C48128 a_10425_46660# VSS 9.68e-19 
C48129 a_10185_46660# VSS 0.002215f 
C48130 a_19692_46634# VSS 1.97188f 
C48131 a_19466_46812# VSS 0.675335f 
C48132 a_19333_46634# VSS 0.289568f 
C48133 a_15227_44166# VSS 2.80559f 
C48134 a_18834_46812# VSS 0.198054f 
C48135 a_17609_46634# VSS 0.205547f 
C48136 a_16292_46812# VSS 0.271203f 
C48137 a_15559_46634# VSS 0.394779f 
C48138 a_15368_46634# VSS 0.278142f 
C48139 a_14976_45028# VSS 0.479565f 
C48140 a_3090_45724# VSS 2.6372f 
C48141 a_15009_46634# VSS 0.270859f 
C48142 a_14084_46812# VSS 0.251005f 
C48143 a_13607_46688# VSS 0.218935f 
C48144 a_12816_46660# VSS 0.260317f 
C48145 a_12991_46634# VSS 0.475827f 
C48146 a_12251_46660# VSS 0.270927f 
C48147 a_12469_46902# VSS 0.193369f 
C48148 a_11901_46660# VSS 0.303844f 
C48149 a_11813_46116# VSS 0.563718f 
C48150 a_11735_46660# VSS 0.520568f 
C48151 a_11186_47026# VSS 0.078586f 
C48152 a_10768_47026# VSS 0.006047f 
C48153 a_8846_46660# VSS 0.002215f 
C48154 a_8601_46660# VSS 9.68e-19 
C48155 a_8270_45546# VSS 0.779033f 
C48156 a_8189_46660# VSS 0.004992f 
C48157 a_8023_46660# VSS 0.006939f 
C48158 a_6903_46660# VSS 0.002857f 
C48159 a_6682_46660# VSS 0.002596f 
C48160 a_8035_47026# VSS 0.004694f 
C48161 a_7832_46660# VSS 0.073862f 
C48162 a_6086_46660# VSS 0.001266f 
C48163 a_5841_46660# VSS 4.65e-19 
C48164 a_6999_46987# VSS 2.7e-19 
C48165 a_6969_46634# VSS 0.289597f 
C48166 a_6755_46942# VSS 3.33348f 
C48167 a_10249_46116# VSS 0.414443f 
C48168 a_10554_47026# VSS 0.191251f 
C48169 a_10623_46897# VSS 0.283572f 
C48170 a_10467_46802# VSS 0.523954f 
C48171 a_10428_46928# VSS 0.314538f 
C48172 a_10150_46912# VSS 0.276624f 
C48173 a_9863_46634# VSS 0.607398f 
C48174 a_8492_46660# VSS 0.283316f 
C48175 a_8667_46634# VSS 0.596387f 
C48176 a_7927_46660# VSS 0.269867f 
C48177 a_8145_46902# VSS 0.179735f 
C48178 a_7577_46660# VSS 0.314978f 
C48179 a_7715_46873# VSS 0.546182f 
C48180 a_7411_46660# VSS 0.532412f 
C48181 a_5257_43370# VSS 1.42323f 
C48182 a_5429_46660# VSS 0.004992f 
C48183 a_5263_46660# VSS 0.006939f 
C48184 a_3878_46660# VSS 0.002215f 
C48185 a_3633_46660# VSS 9.68e-19 
C48186 a_5275_47026# VSS 0.005488f 
C48187 a_5072_46660# VSS 0.073862f 
C48188 a_6540_46812# VSS 0.248814f 
C48189 a_5732_46660# VSS 0.260482f 
C48190 a_5907_46634# VSS 0.473347f 
C48191 a_5167_46660# VSS 0.263586f 
C48192 a_5385_46902# VSS 0.17737f 
C48193 a_4817_46660# VSS 0.296797f 
C48194 a_4955_46873# VSS 0.365781f 
C48195 a_4651_46660# VSS 0.548065f 
C48196 a_4646_46812# VSS 2.12519f 
C48197 a_3877_44458# VSS 2.8543f 
C48198 a_3221_46660# VSS 0.00579f 
C48199 a_3055_46660# VSS 0.008634f 
C48200 a_2162_46660# VSS 0.006278f 
C48201 a_1302_46660# VSS 0.001378f 
C48202 a_1057_46660# VSS 5.58e-19 
C48203 a_3067_47026# VSS 0.004694f 
C48204 a_2864_46660# VSS 0.080001f 
C48205 a_3524_46660# VSS 0.267612f 
C48206 a_3699_46634# VSS 0.499647f 
C48207 a_2959_46660# VSS 0.261026f 
C48208 a_3177_46902# VSS 0.184239f 
C48209 a_2609_46660# VSS 0.302878f 
C48210 a_2443_46660# VSS 0.657702f 
C48211 a_n2661_46098# VSS 2.05975f 
C48212 a_1799_45572# VSS 0.30194f 
C48213 a_645_46660# VSS 0.006691f 
C48214 a_479_46660# VSS 0.008994f 
C48215 a_1110_47026# VSS 8.17e-20 
C48216 a_n935_46688# VSS 0.004685f 
C48217 a_491_47026# VSS 0.010533f 
C48218 a_288_46660# VSS 0.075217f 
C48219 a_1983_46706# VSS 0.205951f 
C48220 a_2107_46812# VSS 1.13475f 
C48221 a_948_46660# VSS 0.263413f 
C48222 a_1123_46634# VSS 0.776627f 
C48223 a_383_46660# VSS 0.269735f 
C48224 a_601_46902# VSS 0.192316f 
C48225 a_33_46660# VSS 0.309712f 
C48226 a_171_46873# VSS 0.579977f 
C48227 a_n133_46660# VSS 0.576523f 
C48228 a_n2438_43548# VSS 2.99787f 
C48229 a_n743_46660# VSS 3.29885f 
C48230 a_n1021_46688# VSS 0.271211f 
C48231 a_n1925_46634# VSS 1.33202f 
C48232 a_n2312_38680# VSS 2.0221f 
C48233 a_n2104_46634# VSS 0.340006f 
C48234 a_n2293_46634# VSS 1.52366f 
C48235 a_n2442_46660# VSS 1.32617f 
C48236 a_n2472_46634# VSS 0.323981f 
C48237 a_n2661_46634# VSS 0.742038f 
C48238 a_n2956_39768# VSS 1.30197f 
C48239 a_n2840_46634# VSS 0.328049f 
C48240 a_22612_30879# VSS 3.18235f 
C48241 a_21588_30879# VSS 2.65298f 
C48242 a_20916_46384# VSS 0.827544f 
C48243 a_20843_47204# VSS 0.121976f 
C48244 a_19594_46812# VSS 0.277274f 
C48245 a_19321_45002# VSS 1.15234f 
C48246 a_19452_47524# VSS 0.006141f 
C48247 a_13747_46662# VSS 2.11905f 
C48248 a_13661_43548# VSS 2.82749f 
C48249 a_5807_45002# VSS 2.5828f 
C48250 a_16131_47204# VSS 0.004694f 
C48251 a_16942_47570# VSS 0.001266f 
C48252 a_16697_47582# VSS 4.65e-19 
C48253 a_16285_47570# VSS 0.004992f 
C48254 a_16119_47582# VSS 0.006939f 
C48255 a_15928_47570# VSS 0.075455f 
C48256 a_768_44030# VSS 3.03052f 
C48257 a_12549_44172# VSS 2.68201f 
C48258 a_12891_46348# VSS 1.22195f 
C48259 a_11309_47204# VSS 0.423399f 
C48260 a_11117_47542# VSS 0.003386f 
C48261 a_10037_47542# VSS 0.004685f 
C48262 a_9804_47204# VSS 0.528639f 
C48263 a_8128_46384# VSS 0.573494f 
C48264 a_5159_47243# VSS 2.7e-19 
C48265 a_7989_47542# VSS 0.004685f 
C48266 a_n881_46662# VSS 4.56296f 
C48267 a_n1613_43370# VSS 4.90074f 
C48268 a_3411_47243# VSS 4.87e-19 
C48269 a_3094_47243# VSS 3.78e-19 
C48270 a_5063_47570# VSS 0.003543f 
C48271 a_4842_47570# VSS 0.003279f 
C48272 a_2583_47243# VSS 2.7e-19 
C48273 a_2266_47243# VSS 6.13e-20 
C48274 a_3315_47570# VSS 0.003543f 
C48275 a_3094_47570# VSS 0.003279f 
C48276 a_7_47243# VSS 2.7e-19 
C48277 a_2747_46873# VSS 0.287894f 
C48278 a_2487_47570# VSS 0.003543f 
C48279 a_2266_47570# VSS 0.003328f 
C48280 a_n89_47570# VSS 0.002898f 
C48281 a_n310_47570# VSS 0.003279f 
C48282 a_n2312_39304# VSS 1.49307f 
C48283 a_n2312_40392# VSS 2.25565f 
C48284 a_22959_47212# VSS 0.322938f 
C48285 a_11453_44696# VSS 0.689179f 
C48286 SMPL_ON_N VSS 2.60102f 
C48287 a_22731_47423# VSS 0.227778f 
C48288 a_22223_47212# VSS 0.332189f 
C48289 a_12465_44636# VSS 5.61685f 
C48290 a_21811_47423# VSS 0.23358f 
C48291 a_4883_46098# VSS 1.54736f 
C48292 a_21496_47436# VSS 0.249536f 
C48293 a_13507_46334# VSS 4.83849f 
C48294 a_21177_47436# VSS 0.223524f 
C48295 a_20990_47178# VSS 0.224581f 
C48296 a_20894_47436# VSS 0.233111f 
C48297 a_19787_47423# VSS 0.258015f 
C48298 a_19386_47436# VSS 0.209882f 
C48299 a_18597_46090# VSS 2.82344f 
C48300 a_18780_47178# VSS 0.319719f 
C48301 a_18479_47436# VSS 1.19826f 
C48302 a_18143_47464# VSS 0.579061f 
C48303 a_10227_46804# VSS 8.12328f 
C48304 a_17591_47464# VSS 0.576556f 
C48305 a_16588_47582# VSS 0.263715f 
C48306 a_16763_47508# VSS 0.587861f 
C48307 a_16023_47582# VSS 0.264352f 
C48308 a_16327_47482# VSS 5.17799f 
C48309 a_16241_47178# VSS 0.18232f 
C48310 a_15673_47210# VSS 0.315684f 
C48311 a_15811_47375# VSS 0.349499f 
C48312 a_15507_47210# VSS 0.556554f 
C48313 a_11599_46634# VSS 2.84967f 
C48314 a_14955_47212# VSS 0.358339f 
C48315 a_14311_47204# VSS 0.248858f 
C48316 a_13487_47204# VSS 0.643275f 
C48317 a_12861_44030# VSS 3.64545f 
C48318 a_13717_47436# VSS 1.02478f 
C48319 a_n1435_47204# VSS 9.72476f 
C48320 a_13381_47204# VSS 0.225132f 
C48321 a_11459_47204# VSS 0.553679f 
C48322 a_9313_45822# VSS 1.04727f 
C48323 a_11031_47542# VSS 0.247302f 
C48324 a_9863_47436# VSS 0.265619f 
C48325 a_9067_47204# VSS 0.606182f 
C48326 a_6575_47204# VSS 0.798434f 
C48327 a_7903_47542# VSS 0.258657f 
C48328 a_7227_47204# VSS 0.610401f 
C48329 a_6851_47204# VSS 0.346433f 
C48330 a_6491_46660# VSS 0.343406f 
C48331 a_6545_47178# VSS 0.597936f 
C48332 a_6151_47436# VSS 2.12954f 
C48333 a_5815_47464# VSS 0.594449f 
C48334 a_5129_47502# VSS 0.361487f 
C48335 a_4915_47217# VSS 2.79467f 
C48336 a_n443_46116# VSS 4.167f 
C48337 a_4791_45118# VSS 2.65418f 
C48338 a_4700_47436# VSS 0.271201f 
C48339 a_4007_47204# VSS 0.628996f 
C48340 a_3815_47204# VSS 0.440491f 
C48341 a_3785_47178# VSS 0.541893f 
C48342 a_3381_47502# VSS 0.320926f 
C48343 a_n1151_42308# VSS 3.78206f 
C48344 a_3160_47472# VSS 0.607125f 
C48345 a_2905_45572# VSS 0.47073f 
C48346 a_2952_47436# VSS 0.275026f 
C48347 a_2553_47502# VSS 0.294118f 
C48348 a_2063_45854# VSS 1.92678f 
C48349 a_584_46384# VSS 2.10508f 
C48350 a_2124_47436# VSS 0.276508f 
C48351 a_1431_47204# VSS 0.595895f 
C48352 a_1239_47204# VSS 0.33333f 
C48353 a_1209_47178# VSS 0.474725f 
C48354 a_327_47204# VSS 0.581187f 
C48355 a_n785_47204# VSS 0.361759f 
C48356 a_n23_47502# VSS 0.278861f 
C48357 a_n237_47217# VSS 3.05697f 
C48358 a_n746_45260# VSS 0.993718f 
C48359 a_n971_45724# VSS 4.81311f 
C48360 a_n452_47436# VSS 0.28781f 
C48361 a_n815_47178# VSS 0.513835f 
C48362 a_n1605_47204# VSS 0.250546f 
C48363 SMPL_ON_P VSS 4.94844f 
C48364 a_n1741_47186# VSS 1.81488f 
C48365 a_n1920_47178# VSS 0.310881f 
C48366 a_n2109_47186# VSS 0.936844f 
C48367 a_n2288_47178# VSS 0.346995f 
C48368 a_n2497_47436# VSS 2.31207f 
C48369 a_n2833_47464# VSS 0.602779f 
C48370 w_11334_34010# VSS 51.3801f 
C48371 w_1575_34946# VSS 51.6622f 
.ends
