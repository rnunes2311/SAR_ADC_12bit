* NGSPICE file created from SAR_ADC_12bit_flat.ext - technology: sky130A

.subckt SAR_ADC_12bit VDD VCM VSS VREF VIN_P VIN_N RST_Z CLK_DATA DATA[5] DATA[4] DATA[3] DATA[2] DATA[1] DATA[0] START
+ EN_OFFSET_CAL DEBUG_MUX[3] DEBUG_MUX[2] DEBUG_MUX[1] DEBUG_MUX[0] DEBUG_OUT CLK
X0 a_n2840_46500# a_n2661_46508.t4 VSS.t2560 VSS.t2559 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1 VDAC_N.t1081 C6_N_btm.t21 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2 a_8912_37509.t27 VDAC_P.t1081 a_5088_37509.t9 VDD.t2245 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3 VSS.t2562 a_18445_42718# a_19187_42718# VSS.t2561 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VDAC_P.t2133 C10_P_btm.t44 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5 a_n1522_42718.t1 a_n1552_42692# VSS.t2570 VSS.t2569 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X6 VDAC_N.t2133 C10_N_btm.t41 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7 VDAC_N.t291 C10_N_btm.t117 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8 a_10414_43780# a_10844_44364# VSS.t2574 VSS.t2573 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.11975 ps=1.045 w=0.42 l=0.15
X9 C10_P_btm.t1072 a_n2810_44894.t4 VSS.t3272 VSS.t3271 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X10 VDD.t31 a_9521_45982.t13 a_9803_45982# VDD.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X11 VSS.t2582 a_11415_45670# a_9349_46539# VSS.t2581 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X12 VDAC_N.t2131 C10_N_btm.t83 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X13 VDAC_P.t291 C8_P_btm.t45 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X14 a_5088_37509.t12 VDAC_P.t2131 a_8912_37509.t30 VDD.t2254 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X15 VDAC_N.t1079 C9_N_btm.t41 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X16 VDAC_P.t1079 C10_P_btm.t48 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X17 VDAC_P.t2129 C9_P_btm.t70 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X18 VDAC_P.t553 C9_P_btm.t529 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X19 a_2512_45982# a_1597_45982# a_2165_46224# VSS.t2587 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X20 VDAC_P.t2127 C9_P_btm.t324 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X21 VDAC_N.t2129 C10_N_btm.t116 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X22 VSS.t2381 VSS.t2382 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X23 VDAC_P.t1077 C9_P_btm.t288 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X24 VDAC_P.t2125 C9_P_btm.t260 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X25 VDAC_P.t159 C10_P_btm.t64 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X26 VDAC_P.t2123 C8_P_btm.t93 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X27 VDAC_N.t553 C9_N_btm.t64 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X28 VDAC_P.t1075 C10_P_btm.t95 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X29 VDD.t2687 a_22521_39947# a_22469_39973# VDD.t2686 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X30 VDAC_N.t2127 C9_N_btm.t146 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X31 VDD.t2304 VSS.t3683 VDD.t2303 VDD.t2302 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X32 VSS.t2594 a_5663_45982# a_8055_45491# VSS.t2593 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X33 VDAC_N.t1077 C10_N_btm.t515 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X34 w_1375_34946.t3 a_n1123_35174.t4 w_1375_34946.t3 w_1375_34946.t2 sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X35 C10_N_btm.t33 a_22812_30659.t19 VREF.t42 VDD.t531 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X36 VSS.t2602 a_19633_43262# a_21303_42718# VSS.t2601 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X37 a_9547_46565# a_n53_44363.t13 a_9547_46892# VSS.t620 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X38 a_14194_46348# a_13524_46832.t4 VDD.t536 VDD.t535 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X39 VDAC_P.t2121 C9_P_btm.t245 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X40 a_18918_45758# a_7208_47044# a_19168_45758# VSS.t2615 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X41 a_9863_43958# a_1053_45123.t2 a_10037_43834# VSS.t579 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X42 VSS.t586 a_9096_45276.t2 a_8848_44868# VSS.t585 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X43 VDD.t2454 VSS.t3594 VDD.t2453 VDD.t2333 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X44 SMPL_ON_P.t6 a_n2038_35608# VDD.t2719 VDD.t2718 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X45 VSS.t573 a_15730_45670.t17 a_16140_44894# VSS.t572 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X46 VDD.t539 a_n1459_43236.t9 a_22959_44894# VDD.t538 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X47 a_5088_37509.t3 VSS.t3798 VDAC_Ni.t4 VDD.t2286 sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X48 a_2113_38308# VDAC_Ni.t9 a_2112_39137# VSS.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X49 a_12845_42968# a_10259_42870.t17 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X50 VDAC_N.t2125 C8_N_btm.t41 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X51 VDAC_N.t159 C8_N_btm.t94 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X52 VDD.t597 a_13273_44868.t23 a_12931_44894# VDD.t596 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X53 VDAC_N.t2123 C7_N_btm.t33 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X54 VDAC_P.t551 C7_P_btm.t65 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X55 a_20892_30659.t1 a_22959_46534# VSS.t2636 VSS.t1203 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X56 a_n1551_45412.t4 a_10259_42870.t25 VDD.t16 VDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X57 VDAC_N.t1075 C9_N_btm.t167 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X58 VDAC_P.t2119 C8_P_btm.t271 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X59 VDD.t606 a_n1735_43236.t8 a_n1741_42692# VDD.t605 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X60 VDAC_P.t1073 C8_P_btm.t46 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X61 VDAC_P.t2117 C10_P_btm.t242 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X62 VDAC_P.t289 C10_P_btm.t490 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X63 VDAC_N.t2121 C10_N_btm.t198 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X64 VCM.t41 a_3222_30651.t15 VDAC_P.t4 VSS.t666 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X65 VDAC_P.t1071 C9_P_btm.t117 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X66 VDAC_N.t551 C2_N_btm.t5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X67 a_9266_44350# a_9179_44592# a_8862_44482# VDD.t2736 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X68 VDD.t67 COMP_P.t9 a_n1237_42718# VDD.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X69 VSS.t2480 VSS.t2481 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X70 a_n2467_30659.t0 a_n2472_47044# VSS.t2648 VSS.t1669 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X71 VDAC_P.t2113 C10_P_btm.t1031 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X72 VDAC_N.t2119 C9_N_btm.t263 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X73 a_10227_47214.t5 a_11795_47044# VDD.t2753 VDD.t2752 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X74 VDAC_N.t1073 C8_N_btm.t103 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X75 VDAC_N.t2117 C10_N_btm.t361 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X76 C8_P_btm.t0 a_n2810_47070.t4 VREF.t0 VDD.t86 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X77 SMPL_ON_N.t5 a_21789_35634# VDD.t2757 VDD.t2756 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X78 a_1343_38525.t7 a_1177_38525# VDD.t2771 VDD.t2770 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X79 a_19058_43806# a_8727_47222.t4 VSS.t78 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X80 VDAC_N.t289 C9_N_btm.t267 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X81 VDAC_N.t2115 C10_N_btm.t573 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X82 VDAC_P.t549 C10_P_btm.t139 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X83 VDAC_P.t2111 C10_P_btm.t147 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X84 VDAC_P.t1069 C9_P_btm.t102 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X85 VDAC_P.t2109 C10_P_btm.t266 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X86 a_n1920_47588# a_n1741_47596.t5 VDD.t271 VDD.t270 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X87 VDAC_P.t93 C10_P_btm.t344 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X88 VDAC_N.t1071 C8_N_btm.t246 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X89 VDAC_P.t2107 C9_P_btm.t53 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X90 VSS.t2679 a_2151_45670# a_1735_46195# VSS.t2678 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X91 VDAC_N.t2113 C10_N_btm.t634 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X92 a_18958_44350# a_17881_44356# a_18796_44728# VDD.t2781 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X93 VSS.t3593 C10_N_btm.t1079 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X94 VDD.t2560 VSS.t3790 VDD.t2559 VDD.t2283 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X95 VDAC_P.t1067 C10_P_btm.t420 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X96 VSS.t2690 a_22775_42718# a_22465_38541# VSS.t2689 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X97 VDAC_N.t549 C10_N_btm.t738 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X98 VDAC_P.t2105 C9_P_btm.t46 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X99 VSS.t324 a_n1827_44868.t8 a_22223_47070# VSS.t301 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X100 VDAC_P.t547 C9_P_btm.t38 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X101 a_5142_30651.t3 a_15008_42692# VDD.t2802 VDD.t2801 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X102 VDD.t2804 a_15831_42883# a_13144_47452.t1 VDD.t2803 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X103 VSS.t3410 VDD.t3194 VSS.t3409 VSS.t3408 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X104 VDAC_N.t2111 C9_N_btm.t298 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X105 VDAC_N.t1069 C9_N_btm.t344 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X106 VDAC_N.t2109 C6_N_btm.t22 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X107 a_15589_44670# a_12769_44594.t2 VSS.t57 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X108 VDAC_P.t2103 C9_P_btm.t527 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X109 VDD.t414 a_n237_45454.t13 a_n377_45776# VDD.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X110 VSS.t3782 C6_N_btm.t66 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X111 VDD.t2097 a_8969_43582# a_9343_42718# VDD.t2096 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X112 a_22545_39429# a_22459_39581# VDD.t2132 VDD.t2131 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X113 a_10703_46526# a_10079_46532# a_10595_46904# VDD.t2218 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X114 VCM.t34 a_3222_30651.t19 VDAC_N.t6 VSS.t671 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X115 VDAC_N.t2107 C7_N_btm.t119 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X116 a_927_42692.t7 a_4527_43566# VDD.t2174 VDD.t2173 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X117 VDAC_N.t1067 C6_N_btm.t60 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X118 VDAC_P.t1065 C7_P_btm.t11 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X119 VDAC_N.t2105 C10_N_btm.t759 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X120 a_10795_43262# a_10171_43268# a_10687_43640# VDD.t2148 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X121 a_2471_45046# a_927_42692.t23 a_2617_44894# VSS.t100 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X122 a_17930_32299.t1 a_22591_44894# VSS.t2184 VSS.t2183 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X123 VDAC_P.t2101 C10_P_btm.t464 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X124 VDD.t2763 a_21789_35634# SMPL_ON_N.t7 VDD.t2762 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X125 VDAC_N.t547 C9_N_btm.t354 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X126 VDAC_P.t287 C9_P_btm.t31 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X127 VDD.t2769 a_1177_38525# a_1343_38525.t6 VDD.t2768 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X128 VDAC_P.t2099 C9_P_btm.t517 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X129 VREF.t10 a_20163_31459.t4 C3_N_btm.t1 VDD.t412 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X130 VDAC_P.t1063 C8_P_btm.t39 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X131 VDAC_P.t2097 C9_P_btm.t194 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X132 VDAC_N.t2103 C10_N_btm.t793 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X133 a_n2109_47596.t2 a_19520_46500# VDD.t2066 VDD.t2065 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X134 a_505_43640# a_n685_43268# a_396_43640# VSS.t2261 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X135 VSS.t3029 VDD.t3111 VSS.t3028 VSS.t3027 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X136 a_4833_47320# a_n53_44363.t21 VDD.t565 VDD.t564 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X137 VDAC_P.t545 C9_P_btm.t118 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X138 VSS.t2169 a_10467_47212# a_10428_47338# VSS.t2168 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X139 VDAC_N.t1065 C8_N_btm.t143 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X140 VSS.t2503 VSS.t2504 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X141 VDD.t2730 a_22959_46534# a_20892_30659.t3 VDD.t1857 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X142 VDAC_P.t2095 C10_P_btm.t1010 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X143 VSS.t2470 VSS.t2471 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X144 VDAC_N.t2101 C10_N_btm.t812 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X145 VDAC_N.t287 C10_N_btm.t903 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X146 VSS.t476 a_13248_45956.t4 a_16177_45982# VSS.t475 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.08775 ps=0.92 w=0.65 l=0.15
X147 VDAC_N.t2099 C9_N_btm.t361 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X148 VDAC_N.t1063 C9_N_btm.t379 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X149 VDAC_N.t2097 C10_N_btm.t920 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X150 VDAC_N.t545 C10_N_btm.t924 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X151 VDAC_P.t1061 C10_P_btm.t578 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X152 VDAC_P.t2093 C9_P_btm.t54 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X153 VDAC_P.t157 C9_P_btm.t521 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X154 a_5088_37509.t4 VDAC_P.t2091 a_8912_37509.t22 VDD.t2249 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X155 a_4461_43640# a_3271_43268# a_4352_43640# VSS.t2110 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X156 a_15037_46232# a_n1067_42718.t2 a_15121_46232# VDD.t266 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X157 VSS.t2197 a_n1920_42692# a_n1890_42718.t1 VSS.t2196 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X158 VDAC_P.t1059 C10_P_btm.t579 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X159 VSS.t2442 VSS.t2443 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X160 a_10949_43628# a_10905_43236# a_10783_43640# VSS.t2141 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X161 VDD.t2197 a_7195_44868# a_7182_45260# VDD.t2196 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X162 VDAC_N.t2095 C3_N_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X163 VSS.t74 a_n1551_45412.t9 a_n2293_44332# VSS.t73 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X164 VDD.t2130 a_22399_44894# a_22959_43806# VDD.t873 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X165 VDAC_P.t2089 C8_P_btm.t23 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X166 a_834_46348# a_n243_45982# a_672_45982# VDD.t854 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X167 VSS.t408 a_1334_43494.t26 a_1339_43315# VSS.t407 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X168 VDAC_N.t1061 C8_N_btm.t144 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X169 VDD.t2785 a_22775_42718# a_22465_38541# VDD.t2784 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X170 VDAC_N.t2093 C10_N_btm.t941 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X171 VDAC_P.t543 C7_P_btm.t62 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X172 VDAC_P.t2087 C10_P_btm.t664 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X173 VDAC_P.t1057 C8_P_btm.t20 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X174 VDAC_P.t2085 C8_P_btm.t256 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X175 VDAC_N.t157 C9_N_btm.t398 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X176 VDAC_P.t285 C9_P_btm.t39 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X177 a_3897_45444# a_3731_45444# VSS.t2151 VSS.t2150 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X178 VDAC_N.t2091 C10_N_btm.t975 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X179 VSS.t3574 C10_P_btm.t19 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X180 VDAC_P.t2083 C10_P_btm.t894 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X181 a_11599_42883# a_5734_30651.t4 VDD.t378 VDD.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X182 VDAC_N.t1059 C10_N_btm.t979 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X183 VDAC_N.t2089 C10_N_btm.t994 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X184 VDD.t2109 a_6635_47044# a_n690_43494.t2 VDD.t2108 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X185 VDAC_N.t543 C10_N_btm.t1055 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X186 a_n237_45454.t0 a_11971_46500# VSS.t2189 VSS.t2188 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X187 VDD.t2144 a_2216_46758# a_2167_46526# VDD.t2143 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X188 VDAC_N.t2087 C9_N_btm.t400 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X189 VDAC_N.t1057 C9_N_btm.t405 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X190 VDAC_N.t2085 C9_N_btm.t435 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X191 a_6391_46219# a_6235_46124# a_6536_46348# VDD.t2239 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X192 C8_N_btm.t4 a_17738_32299.t4 VSS.t451 VSS.t450 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X193 a_9863_43958# a_n237_45454.t15 VDD.t416 VDD.t415 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X194 VSS.t2127 a_n2840_47044# a_n2810_47070.t1 VSS.t2126 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X195 VDAC_P.t1055 C9_P_btm.t518 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X196 VSS.t2258 a_20383_42718# a_6974_31099.t1 VSS.t2257 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X197 a_n2840_45412# a_n2661_45420.t5 VDD.t307 VDD.t306 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X198 VDAC_N.t285 C10_N_btm.t54 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X199 VDAC_P.t2081 C10_P_btm.t898 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X200 VDD.t2182 a_9343_43806# a_5655_43780# VDD.t2181 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X201 VDAC_P.t541 C9_P_btm.t189 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X202 VDAC_N.t2083 C7_N_btm.t120 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X203 VDAC_P.t2079 C9_P_btm.t55 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X204 VDAC_P.t1053 C10_P_btm.t961 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X205 VDAC_N.t1055 C9_N_btm.t483 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X206 C9_P_btm.t0 a_n2442_44894.t4 VSS.t367 VSS.t366 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X207 VDAC_P.t2077 C10_P_btm.t974 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X208 VDAC_P.t2135 C7_P_btm.t10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X209 VSS.t3755 C0_dummy_N_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X210 VDAC_N.t2081 C10_N_btm.t51 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X211 VDAC_N.t541 C10_N_btm.t46 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X212 VSS.t2343 VSS.t2344 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X213 VDAC_N.t2079 C10_N_btm.t43 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X214 VDAC_N.t1053 C8_N_btm.t177 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X215 VSS.t426 a_n690_43494.t21 a_2443_43806# VSS.t425 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X216 a_14545_44569# a_14635_44324# VDD.t2160 VDD.t2159 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X217 VDAC_P.t2075 C7_P_btm.t56 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X218 VDAC_N.t2077 C9_N_btm.t254 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X219 VDAC_P.t1051 C10_P_btm.t220 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X220 VDAC_P.t2073 C10_P_btm.t1053 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X221 VDAC_P.t539 C10_P_btm.t56 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X222 VDAC_P.t2071 C9_P_btm.t509 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X223 VDAC_P.t1049 C10_P_btm.t52 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X224 VDAC_N.t2135 C8_N_btm.t186 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X225 VDAC_P.t2069 C9_P_btm.t508 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X226 a_n2661_44332# a_n1827_45412.t8 VDD.t312 VDD.t280 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X227 VDAC_P.t283 C10_P_btm.t49 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X228 VDAC_P.t2067 C10_P_btm.t45 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X229 VDAC_P.t1047 C10_P_btm.t41 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X230 VDAC_N.t2075 C10_N_btm.t39 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X231 VDAC_N.t1051 C10_N_btm.t36 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X232 VDAC_N.t2073 C10_N_btm.t1035 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X233 VDAC_N.t539 C10_N_btm.t478 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X234 a_18319_44868# a_15730_45670.t25 VDD.t504 VDD.t503 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X235 VSS.t2395 VSS.t2396 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X236 VSS.t2345 VSS.t2346 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X237 VDAC_P.t2065 C10_P_btm.t37 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X238 VSS.t2264 a_8192_44874# a_8204_45412# VSS.t2263 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X239 VDAC_N.t2071 C9_N_btm.t121 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X240 VDAC_P.t537 C10_P_btm.t34 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X241 VDAC_N.t1049 C10_N_btm.t222 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X242 VDAC_P.t2063 C8_P_btm.t111 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X243 VSS.t2351 VSS.t2352 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X244 VDAC_N.t2069 C10_N_btm.t111 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X245 VSS.t376 a_1429_47222.t4 a_1431_47070# VSS.t375 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X246 VDAC_N.t283 C10_N_btm.t95 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X247 VSS.t2193 a_14635_44324# a_15323_44894# VSS.t2192 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X248 VDAC_P.t1045 C10_P_btm.t1034 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X249 VDAC_P.t2061 C10_P_btm.t476 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X250 VSS.t3276 a_n2810_44894.t6 C10_P_btm.t1074 VSS.t3275 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X251 VDAC_N.t2067 C5_N_btm.t5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X252 VSS.t2174 a_n2472_43236# a_n2442_43262.t1 VSS.t805 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X253 VSS.t131 a_n1551_44324.t9 a_n2661_43780# VSS.t130 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X254 VDAC_N.t1047 C10_N_btm.t55 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X255 VDAC_N.t2065 VSS.t3309 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X256 a_15133_45144# a_1429_47222.t21 a_15049_45144# VDD.t329 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X257 VDAC_N.t537 C9_N_btm.t57 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X258 VDAC_N.t2063 C10_N_btm.t47 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X259 VDAC_N.t1045 C9_N_btm.t50 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X260 VDAC_N.t2061 C10_N_btm.t40 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X261 VDD.t376 a_n331_42718.t2 a_15121_46232# VDD.t375 sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X262 a_4005_46500# a_3787_46904# VDD.t2107 VDD.t2106 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X263 VDAC_N.t155 C9_N_btm.t25 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X264 VDAC_P.t155 C10_P_btm.t109 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X265 a_3754_39466# a_7754_39300# VSS.t693 sky130_fd_pr__res_high_po_0p35 l=18
X266 VDAC_P.t2059 C10_P_btm.t94 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X267 a_12121_45956# a_11788_46134# VSS.t1646 VSS.t1645 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X268 VDAC_P.t1043 C8_P_btm.t47 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X269 VDAC_P.t2057 C10_P_btm.t53 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X270 C0_dummy_P_btm.t1 a_6974_31099.t4 VCM.t22 VSS.t305 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X271 a_13157_43628# a_13113_43236# a_12991_43640# VSS.t1651 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X272 VDD.t1594 a_570_44324# a_n1459_43236.t6 VDD.t1593 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X273 VDAC_N.t2059 C10_N_btm.t1036 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X274 VDAC_P.t535 C8_P_btm.t96 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X275 VDAC_N.t1043 C10_N_btm.t223 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X276 VDAC_P.t2055 C8_P_btm.t24 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X277 a_n2840_45956# a_n2661_45956.t4 VSS.t431 VSS.t353 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X278 VSS.t3648 C10_P_btm.t16 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X279 VDAC_N.t2057 C10_N_btm.t96 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X280 VDAC_N.t535 C10_N_btm.t48 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X281 VSS.t3463 VDD.t3213 VSS.t3462 VSS.t3461 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X282 VDAC_N.t2055 C8_N_btm.t213 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X283 VDAC_P.t1041 C10_P_btm.t46 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X284 VSS.t3646 C1_P_btm.t2 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X285 VSS.t2584 a_9349_46539# a_9768_46892# VSS.t2583 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X286 VDAC_P.t2053 C9_P_btm.t507 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X287 a_15192_46500# a_15163_45670.t5 a_15415_46846# VSS.t115 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X288 VSS.t3189 VDD.t3165 VSS.t3188 VSS.t3187 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X289 VSS.t1661 a_5441_46500# a_5089_47044# VSS.t1660 sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.169 ps=1.82 w=0.65 l=0.15
X290 a_15582_45982# a_14955_45982# VDD.t1605 VDD.t1604 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X291 SMPL_ON_P.t4 a_n2038_35608# VDD.t2721 VDD.t2720 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X292 a_n2472_46500# a_n2293_46508.t4 VSS.t106 VSS.t105 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X293 VDAC_P.t281 C6_P_btm.t8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X294 a_4514_43262# a_3437_43268# a_4352_43640# VDD.t1610 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X295 a_12557_43806# a_11367_43806# a_12448_43806# VSS.t1676 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X296 VDAC_P.t2051 C10_P_btm.t38 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X297 VDAC_N.t1041 C10_N_btm.t1037 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X298 a_3787_46904# a_3271_46532# a_3692_46892# VSS.t1680 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X299 VSS.t3720 C10_P_btm.t26 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X300 VSS.t611 a_13524_46832.t23 a_14373_47070# VSS.t610 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X301 a_82_45670# a_847_45956# VSS.t1685 VSS.t1684 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X302 VDAC_N.t2053 C10_N_btm.t1028 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X303 VDAC_P.t1039 C9_P_btm.t506 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X304 VIN_N.t9 EN_VIN_BSTR_N.t7 C7_N_btm.t2 VSS.t436 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X305 VDAC_N.t281 C7_N_btm.t72 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X306 VSS.t3165 VDD.t3157 VSS.t3164 VSS.t3163 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X307 VDAC_P.t2049 C9_P_btm.t505 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X308 VDAC_P.t533 C9_P_btm.t504 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X309 VDD.t447 a_7754_40130.t9 a_11206_38545.t3 VDD.t446 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X310 VDAC_P.t2047 C10_P_btm.t1035 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X311 VDAC_N.t2051 C10_N_btm.t508 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X312 VSS.t3604 C7_N_btm.t133 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X313 VDAC_N.t1039 C10_N_btm.t1025 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X314 VSS.t491 a_13248_45956.t25 a_15079_46134# VSS.t490 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X315 VDAC_N.t2049 C10_N_btm.t1024 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X316 VDAC_N.t533 C10_N_btm.t1023 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X317 VDAC_N.t2047 C10_N_btm.t1022 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X318 VDAC_P.t1037 C10_P_btm.t221 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X319 VDAC_N.t1037 C9_N_btm.t22 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X320 VDD.t363 a_n690_43494.t15 a_2443_43806# VDD.t362 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X321 VDAC_N.t2045 C9_N_btm.t18 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X322 VDAC_P.t2045 C10_P_btm.t1026 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X323 VDD.t2298 VSS.t3713 VDD.t2297 VDD.t2296 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X324 VDAC_P.t91 C9_P_btm.t503 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X325 VDAC_P.t2043 VSS.t3380 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X326 a_n2293_43244# a_n1827_44324.t5 VDD.t261 VDD.t260 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X327 VDAC_P.t1035 C7_P_btm.t9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X328 VDAC_N.t91 VSS.t3290 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X329 a_9987_42968# a_2755_43494.t22 a_10069_42968# VDD.t432 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X330 VDAC_N.t2043 C8_N_btm.t218 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X331 a_3470_46232# a_1847_45528.t17 VDD.t2884 VDD.t2883 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X332 VREF.t45 a_22812_30659.t17 C10_N_btm.t31 VDD.t529 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X333 VDAC_N.t1035 C9_N_btm.t515 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X334 VDD.t1641 a_3823_42718# a_4000_42718.t3 VDD.t1640 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X335 a_7374_44894# a_5655_43780# VSS.t2250 VSS.t2249 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X336 a_15935_43640# a_15489_43268# a_15839_43640# VSS.t1701 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X337 VDAC_P.t2041 C3_P_btm.t5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X338 a_2755_43494.t1 a_13536_43780# VSS.t1706 VSS.t1705 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X339 VSS.t276 a_2587_44868.t33 a_4703_44894# VSS.t275 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X340 VDAC_N.t2041 C10_N_btm.t1020 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X341 a_7735_45477# a_6985_45438# a_7276_45670# VDD.t1652 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X342 VDAC_N.t531 C10_N_btm.t1019 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X343 VDD.t1656 a_6091_43780# a_6078_44172# VDD.t1655 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X344 a_927_42692.t4 a_4527_43566# VDD.t2176 VDD.t2175 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X345 VDAC_P.t531 C10_P_btm.t1025 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X346 VDAC_N.t2039 C10_N_btm.t1018 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X347 VDD.t2276 VSS.t3706 VDD.t2275 VDD.t2274 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X348 VDAC_P.t2039 VSS.t3379 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X349 VSS.t3026 VDD.t3110 VSS.t3025 VSS.t3024 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X350 VDAC_P.t1033 C10_P_btm.t1024 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X351 a_15155_47070# a_15113_47222# VSS.t1723 VSS.t1722 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X352 VDAC_P.t2037 C10_P_btm.t1023 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X353 C10_N_btm.t27 a_22812_30659.t13 VREF.t41 VDD.t525 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X354 VDD.t1668 a_4005_43236# a_3895_43262# VDD.t1667 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X355 a_8969_43582# a_1203_42692.t33 a_8981_43262# VDD.t486 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X356 a_n1551_44324.t4 a_10414_43780# VDD.t2666 VDD.t2665 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X357 VDAC_N.t1033 C10_N_btm.t1017 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X358 VSS.t3020 VDD.t3108 VSS.t3019 VSS.t3018 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X359 VSS.t1729 a_16291_44914# a_18495_44868# VSS.t1728 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X360 VDAC_N.t2037 C10_N_btm.t1016 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X361 VDD.t1684 a_7429_47044# a_7459_47397# VDD.t1683 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X362 VDAC_N.t279 C10_N_btm.t1015 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X363 VDAC_P.t279 C10_P_btm.t1022 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X364 VDD.t1686 a_21629_47833# a_14766_45596.t1 VDD.t1685 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X365 VDAC_N.t2035 C10_N_btm.t1014 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X366 VDAC_N.t1031 C8_N_btm.t223 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X367 VDAC_N.t2033 C10_N_btm.t1029 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X368 VDAC_P.t2035 C10_P_btm.t1021 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X369 VDD.t1688 a_22591_47070# a_21020_30659.t3 VDD.t1687 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X370 VDAC_P.t1031 C9_P_btm.t511 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X371 VDAC_P.t2033 C10_P_btm.t1020 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X372 VDAC_N.t529 C8_N_btm.t245 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X373 C10_N_btm.t1 a_18314_32299.t5 VSS.t248 VSS.t247 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X374 VDD.t1694 a_16475_45412# a_18759_42746# VDD.t1693 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X375 a_n519_43268# a_n685_43268# VSS.t2260 VSS.t2259 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X376 VDAC_P.t529 C9_P_btm.t510 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X377 a_n283_35174# VDD.t3120 EN_VIN_BSTR_P.t2 VSS.t3054 sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.9
X378 VDAC_N.t2031 C9_N_btm.t15 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X379 a_n2293_47044.t3 a_16576_44868# VDD.t1704 VDD.t1703 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X380 VDD.t2872 a_n2103_45412.t9 a_22959_47622# VDD.t314 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X381 a_21629_47833# DEBUG_MUX[2].t0 VDD.t2829 VDD.t2828 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X382 a_396_43640# a_n519_43268# a_49_43236# VSS.t1752 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X383 a_21755_44350# a_n2661_46508.t6 VSS.t2556 VSS.t2555 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X384 VSS.t2734 a_n1732_35090.t8 a_n283_35174# VSS.t2733 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X385 a_12562_46642# a_11455_44576.t17 VDD.t2818 VDD.t2817 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X386 a_18282_45670# a_15730_45670.t19 VSS.t575 VSS.t574 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X387 VDD.t1716 a_1239_39587# COMP_P.t4 VDD.t1715 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X388 VDAC_N.t1029 C7_N_btm.t76 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X389 VDAC_N.t2029 C10_N_btm.t1026 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X390 C10_P_btm.t4 a_3990_30651.t15 VCM.t14 VSS.t287 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X391 a_14545_44569# a_14635_44324# VSS.t2195 VSS.t2194 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X392 a_12461_44670# a_11455_44576.t25 VSS.t2722 VSS.t2721 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X393 a_n2661_46508.t3 a_10596_44324# VSS.t1777 VSS.t1776 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X394 VDAC_P.t2031 C7_P_btm.t121 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X395 VDAC_N.t153 C9_N_btm.t505 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X396 VSS.t3565 C6_P_btm.t4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X397 VDAC_N.t2027 C5_N_btm.t7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X398 VDAC_P.t1029 C9_P_btm.t501 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X399 VDD.t463 a_1736_39043.t3 a_1239_39043# VDD.t462 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X400 VDAC_P.t2029 C8_P_btm.t95 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X401 a_19274_43262# a_19003_43262# a_19191_43262# VDD.t1733 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X402 VDAC_N.t1027 C10_N_btm.t1021 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X403 VDD.t2497 VSS.t3563 VDD.t2496 VDD.t2495 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X404 VDAC_P.t153 VSS.t3374 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X405 a_4352_43640# a_3437_43268# a_4005_43236# VSS.t1671 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X406 VDAC_P.t2027 C10_P_btm.t1017 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X407 VDAC_N.t2025 C9_N_btm.t58 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X408 VDD.t1737 a_2134_44324# a_n1735_43236.t6 VDD.t1736 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X409 VDAC_N.t527 C10_N_btm.t1011 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X410 VDAC_N.t2023 C10_N_btm.t1010 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X411 VSS.t3558 C9_P_btm.t24 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X412 VDAC_N.t1025 C10_N_btm.t1009 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X413 VDAC_P.t1027 C9_P_btm.t497 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X414 a_5159_46309# a_4908_45956# a_4700_46134# VDD.t1742 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X415 VDAC_N.t2021 C10_N_btm.t1008 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X416 VDAC_P.t2025 C10_P_btm.t1016 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X417 VDAC_P.t527 C9_P_btm.t498 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X418 VDAC_P.t2023 C10_P_btm.t1015 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X419 VDAC_N.t277 C10_N_btm.t1007 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X420 VDAC_P.t1025 C9_P_btm.t496 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X421 VDAC_N.t2019 C10_N_btm.t1006 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X422 VDAC_P.t2021 C9_P_btm.t495 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X423 a_4527_46830# a_135_43540.t31 VDD.t180 VDD.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X424 VDAC_P.t277 C9_P_btm.t494 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X425 VSS.t1807 a_1387_42883# a_546_43100# VSS.t1806 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X426 VDAC_N.t1023 C10_N_btm.t1005 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X427 VDD.t2353 VSS.t3553 VDD.t2352 VDD.t2351 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X428 VSS.t45 a_13144_47452.t2 a_12896_47044# VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X429 VDAC_P.t2019 C10_P_btm.t1014 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X430 VDAC_N.t2017 C10_N_btm.t1004 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X431 VDAC_N.t525 C10_N_btm.t1003 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X432 VDAC_P.t1023 C10_P_btm.t1013 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X433 VDAC_N.t2015 C10_N_btm.t1002 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X434 VSS.t2568 a_n1552_42692# a_n1522_42718.t0 VSS.t2567 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X435 VDAC_P.t2017 C10_P_btm.t1028 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X436 a_4997_44670# a_4322_46134# a_4651_44350# VSS.t1829 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X437 VDAC_N.t1021 C10_N_btm.t1001 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X438 VDAC_N.t2013 C10_N_btm.t1000 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X439 VDAC_P.t525 C8_P_btm.t257 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X440 VDAC_N.t59 C7_N_btm.t98 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X441 a_1387_42883# a_134_42718.t4 VSS.t2705 VSS.t2704 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X442 VDAC_P.t2015 C9_P_btm.t493 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X443 VDAC_N.t2011 C8_N_btm.t97 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X444 VDAC_N.t1019 C8_N_btm.t259 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X445 VSS.t2359 VSS.t2360 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X446 a_11692_46134# a_7208_47044# a_11834_45982# VSS.t2612 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X447 a_1893_45144# a_1429_47222.t15 a_1798_45144# VDD.t324 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X448 VDAC_N.t2009 C7_N_btm.t61 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X449 VSS.t1838 a_18103_46768# a_18064_46642# VSS.t1837 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X450 VSS.t2795 a_n2810_44350.t4 C8_P_btm.t274 VSS.t2794 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X451 VDAC_P.t1021 C7_P_btm.t129 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X452 VSS.t1848 a_22400_42718# a_22780_41381# VSS.t1847 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X453 a_19168_45758# a_7208_47044# a_18918_45758# VSS.t2611 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X454 a_11265_44670# a_10259_42870.t19 VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X455 VDAC_N.t523 C8_N_btm.t9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X456 VDAC_P.t2013 C7_P_btm.t54 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X457 VSS.t1850 a_18689_45412# a_17763_44868# VSS.t1849 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X458 VSS.t1858 a_22733_47833# a_15163_45670.t0 VSS.t1857 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X459 VDAC_N.t2007 VSS.t3313 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X460 VDAC_N.t1017 C10_N_btm.t999 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X461 VSS.t1868 a_18971_44654# a_18905_44728# VSS.t1867 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X462 VDAC_P.t59 C9_P_btm.t492 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X463 a_12427_46758# a_12699_46616# VSS.t1870 VSS.t1869 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X464 a_16046_47070# a_15582_45982# a_15879_47320# VSS.t1666 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X465 VDAC_N.t2005 C10_N_btm.t998 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X466 a_2864_43806# a_2627_42718# VDD.t1343 VDD.t1342 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X467 VDAC_P.t2011 C10_P_btm.t1027 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X468 DATA[3].t3 a_4651_47614# VSS.t1420 VSS.t1419 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X469 VSS.t1831 a_4322_46134# a_4993_47044# VSS.t1830 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X470 VDD.t1367 a_14950_43958# a_15323_43268# VDD.t1366 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X471 VDAC_P.t1019 C9_P_btm.t491 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X472 VDAC_N.t275 C10_N_btm.t997 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X473 a_10227_47214.t4 a_11795_47044# VDD.t2749 VDD.t2748 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X474 VDD.t2568 VSS.t3762 VDD.t2567 VDD.t2566 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X475 VDAC_N.t2003 C9_N_btm.t26 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X476 VDAC_P.t2009 C9_P_btm.t490 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X477 VDAC_N.t1015 C10_N_btm.t996 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X478 VDAC_P.t523 C10_P_btm.t1018 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X479 VDAC_P.t2007 C10_P_btm.t1012 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X480 VDAC_P.t1017 C10_P_btm.t1008 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X481 VDAC_N.t2001 C10_N_btm.t995 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X482 VDAC_N.t521 C9_N_btm.t190 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X483 a_11143_47588# a_11299_47832# VDD.t1373 VDD.t1372 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X484 VSS.t3659 C10_N_btm.t1069 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X485 C0_N_btm.t1 EN_VIN_BSTR_N.t23 VIN_N.t11 VSS.t445 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X486 VSS.t2649 a_n2472_47044# a_n2467_30659.t1 VSS.t1667 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X487 VDAC_P.t2005 C10_P_btm.t1009 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X488 VSS.t3075 VDD.t3127 VSS.t3074 VSS.t3073 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X489 a_n2472_45412# a_n2293_45420.t5 VDD.t2867 VDD.t1422 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X490 VDAC_N.t1999 C8_N_btm.t7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X491 VSS.t1453 a_22959_43270# a_14297_32299.t1 VSS.t1452 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X492 VDAC_P.t275 C6_P_btm.t31 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X493 VDD.t2928 EN_COMP.t4 a_1177_38525# VDD.t2927 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X494 VDAC_P.t2003 C9_P_btm.t489 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X495 VDAC_P.t1015 C8_P_btm.t48 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X496 VSS.t3413 VDD.t3195 VSS.t3412 VSS.t3411 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X497 a_2655_42870# a_1847_45528.t25 a_2801_42718# VSS.t2809 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X498 a_3165_45982# a_2687_45956# VDD.t1388 VDD.t1387 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X499 VDAC_N.t1013 C7_N_btm.t127 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X500 VCM.t17 a_3990_30651.t19 C10_N_btm.t15 VSS.t292 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X501 VSS.t546 a_1203_42692.t31 a_7735_42692# VSS.t545 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X502 VDAC_N.t1997 C7_N_btm.t59 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X503 VDAC_N.t151 C10_N_btm.t990 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X504 a_713_47044# a_380_47222# VDD.t1401 VDD.t1400 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X505 VDAC_P.t2001 C5_P_btm.t18 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X506 VDAC_P.t521 C10_P_btm.t1007 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X507 VDD.t420 a_n237_45454.t19 a_5441_46500# VDD.t419 sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X508 VDAC_P.t1999 C7_P_btm.t22 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X509 VSS.t3195 VDD.t3167 VSS.t3194 VSS.t3193 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X510 VDAC_N.t1995 C9_N_btm.t19 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X511 VSS.t3732 C8_P_btm.t17 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X512 a_n2103_45412.t7 a_13273_44868.t29 VDD.t601 VDD.t600 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X513 VDAC_P.t1013 C9_P_btm.t488 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X514 VDAC_N.t1011 C9_N_btm.t189 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X515 VDAC_N.t1993 VSS.t3312 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X516 VDAC_P.t1997 C8_P_btm.t249 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X517 VDD.t1407 a_3699_43780# a_1334_43494.t4 VDD.t1406 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X518 a_15689_44048# a_15471_43806# VSS.t1487 VSS.t1486 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X519 a_7429_47044# a_885_44868.t29 VDD.t2848 VDD.t2847 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X520 VDAC_N.t519 C9_N_btm.t506 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X521 VDD.t2968 a_12651_44576.t17 a_12699_46616# VDD.t2967 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X522 a_16475_45412# a_16335_47614# VSS.t1490 VSS.t1489 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X523 C6_P_btm.t69 a_n2810_43806.t4 VSS.t2898 VSS.t2897 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X524 a_n2293_44868# a_n2103_44868.t8 VSS.t2902 VSS.t2901 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X525 VDAC_P.t151 C10_P_btm.t1006 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X526 VSS.t2521 VSS.t2522 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X527 a_8662_43806# a_5655_43780# VSS.t2240 VSS.t2239 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X528 VDAC_N.t1991 C10_N_btm.t989 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X529 VDAC_P.t1995 C10_P_btm.t1005 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X530 a_18357_46224# a_18139_45982# VSS.t1494 VSS.t1493 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X531 VDAC_P.t1011 C10_P_btm.t1004 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X532 VDAC_P.t1993 C8_P_btm.t248 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X533 VDAC_P.t519 C10_P_btm.t1003 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X534 VDAC_N.t1009 C10_N_btm.t988 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X535 VDAC_N.t1989 C10_N_btm.t987 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X536 a_5655_43780# a_9343_43806# VSS.t2215 VSS.t2214 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X537 a_18361_47320# a_14757_47614# VDD.t1429 VDD.t1428 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X538 VDAC_N.t273 C9_N_btm.t187 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X539 VDAC_P.t1991 C10_P_btm.t1002 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X540 VCM.t46 a_5840_42718.t4 C3_N_btm.t11 VSS.t2880 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X541 VDAC_N.t1987 C8_N_btm.t99 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X542 a_18235_45982# a_17789_45982# a_18139_45982# VSS.t1497 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X543 a_4080_44670# a_1847_45528.t19 VSS.t2808 VSS.t2807 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X544 VDD.t1433 a_20049_43262# a_22775_42718# VDD.t1432 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X545 VSS.t1733 a_16291_44914# a_15549_47044.t0 VSS.t1732 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X546 VDAC_P.t1009 C6_P_btm.t39 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X547 a_16177_45982# a_15328_46134# VSS.t1502 VSS.t1501 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X548 VDAC_P.t1989 C6_P_btm.t29 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X549 VDD.t2713 a_9863_43958# a_9416_43530# VDD.t2712 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X550 VDAC_N.t1007 C10_N_btm.t986 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X551 VDAC_N.t1985 C5_N_btm.t8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X552 a_6631_44582# a_7195_44868# VSS.t2228 VSS.t2227 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X553 VDAC_N.t517 C8_N_btm.t6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X554 VSS.t2495 VSS.t2496 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X555 VDD.t2076 a_2471_45046# a_171_44019# VDD.t2075 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X556 VDAC_N.t1983 C7_N_btm.t115 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X557 VDAC_N.t1005 C10_N_btm.t985 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X558 VDAC_P.t273 C7_P_btm.t47 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X559 VDAC_P.t1987 C8_P_btm.t247 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X560 VDAC_N.t1981 C9_N_btm.t27 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X561 VSS.t3490 VDD.t3223 VSS.t3489 VSS.t3488 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X562 a_n2472_45956# a_n2293_45956.t4 VSS.t2855 VSS.t2784 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X563 VDAC_P.t1007 C8_P_btm.t251 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X564 VDAC_P.t1985 C9_P_btm.t487 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X565 VDAC_P.t517 C9_P_btm.t486 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X566 VDAC_N.t89 C10_N_btm.t984 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X567 a_13937_46602# a_10259_42870.t23 VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X568 a_n2840_45956# a_n2661_45956.t6 VDD.t369 VDD.t368 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X569 a_14601_32299.t3 a_22223_44358# VDD.t1456 VDD.t1455 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X570 VDAC_N.t1979 C10_N_btm.t983 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X571 a_13457_46892# a_13427_46756# a_13207_46526# VDD.t1459 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X572 VSS.t1527 a_9343_45982# a_9521_45982.t1 VSS.t1526 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X573 VDAC_N.t1003 C9_N_btm.t498 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X574 a_3733_46348# a_n237_45454.t23 VDD.t319 VDD.t318 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X575 VDAC_P.t1983 C10_P_btm.t1001 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X576 VDAC_P.t1005 C10_P_btm.t1000 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X577 VDAC_P.t1981 C10_P_btm.t999 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X578 a_12448_43806# a_11533_43806# a_12101_44048# VSS.t1530 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X579 VDAC_P.t89 C10_P_btm.t998 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X580 VSS.t2597 a_5663_45982# a_7842_44868# VSS.t2596 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X581 VDAC_N.t1977 C10_N_btm.t982 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X582 VDAC_P.t1979 C8_P_btm.t250 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X583 VSS.t2781 a_14297_32299.t4 C4_N_btm.t1 VSS.t2082 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X584 VDAC_N.t515 C10_N_btm.t981 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X585 VDD.t2327 VSS.t3797 VDD.t2326 VDD.t2258 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X586 VSS.t2653 a_11795_47044# a_10227_47214.t0 VSS.t2652 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X587 VDAC_N.t1975 C10_N_btm.t980 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X588 VDAC_P.t1003 C10_P_btm.t997 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X589 C8_N_btm.t272 a_21276_30659.t4 VREF.t47 VDD.t2930 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X590 VSS.t1538 a_22521_40491# a_22459_39581# VSS.t1537 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X591 VDAC_N.t1001 C9_N_btm.t497 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X592 VDAC_N.t1973 C7_N_btm.t48 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X593 VSS.t3617 C10_N_btm.t1059 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X594 VSS.t1540 a_21847_43806# a_21855_42718# VSS.t1539 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X595 C7_P_btm.t137 a_n2442_44350.t4 VSS.t2826 VSS.t2825 sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X596 VDAC_P.t1977 C10_P_btm.t996 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X597 VDAC_N.t271 C9_N_btm.t496 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X598 VDAC_N.t1971 C9_N_btm.t495 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X599 VDAC_P.t515 C0_dummy_P_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X600 VDD.t33 a_9521_45982.t15 a_10171_43268# VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X601 a_13738_46032# a_13151_45956# a_13654_46032# VSS.t1546 sky130_fd_pr__nfet_01v8 ad=0.10795 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X602 VDAC_P.t1975 C9_P_btm.t485 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X603 VDAC_P.t1001 C10_P_btm.t995 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X604 a_12683_43433# a_12379_44350# VDD.t1484 VDD.t1483 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X605 VDAC_P.t1973 C10_P_btm.t994 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X606 VDAC_N.t999 C5_N_btm.t26 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X607 VDAC_N.t1969 C9_N_btm.t494 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X608 VDAC_P.t271 C10_P_btm.t753 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X609 a_10319_45982# a_9969_45982# a_10224_45982# VDD.t1488 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X610 VSS.t3663 C1_N_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X611 a_13667_32299.t3 a_21855_42718# VDD.t1478 VDD.t1477 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X612 a_7694_46309# a_7648_46134# VDD.t1494 VDD.t1493 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X613 VSS.t2541 VSS.t2542 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X614 VDAC_P.t1971 C9_P_btm.t484 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X615 VSS.t424 a_n690_43494.t19 a_3271_43268# VSS.t423 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X616 VDAC_N.t513 C8_N_btm.t244 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X617 VDAC_N.t1967 C10_N_btm.t978 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X618 VDAC_N.t997 C10_N_btm.t977 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X619 VDD.t1427 a_18357_46224# a_18247_46348# VDD.t1426 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X620 VDAC_N.t1965 C8_N_btm.t32 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X621 VDAC_N.t149 C9_N_btm.t493 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X622 a_16211_43780# a_16036_43806# a_16390_43806# VSS.t1559 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X623 VDAC_P.t999 VSS.t3349 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X624 VDAC_N.t1963 C10_N_btm.t976 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X625 VDAC_P.t1969 C7_P_btm.t46 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X626 VDAC_N.t995 C9_N_btm.t492 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X627 a_6491_44716# a_1847_45528.t23 VDD.t2894 VDD.t2893 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X628 VDAC_N.t1961 C9_N_btm.t491 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X629 VDAC_N.t511 C9_N_btm.t490 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X630 VDAC_P.t513 C10_P_btm.t992 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X631 a_13113_43236# a_12895_43640# VDD.t1504 VDD.t1503 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X632 VDAC_P.t1967 C10_P_btm.t991 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X633 VDAC_P.t997 C8_P_btm.t244 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X634 VSS.t1569 a_7705_45736# a_7639_45804# VSS.t1568 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X635 VDAC_P.t1965 C10_P_btm.t990 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X636 VDAC_P.t149 C9_P_btm.t483 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X637 VSS.t3742 C10_N_btm.t1060 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X638 a_10901_42718# a_7557_43236.t17 VSS.t224 VSS.t223 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X639 VDAC_P.t1963 C10_P_btm.t989 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X640 VSS.t250 a_18314_32299.t6 C10_N_btm.t2 VSS.t249 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X641 VSS.t1573 a_4061_45956# a_3575_46697# VSS.t1572 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X642 VDAC_N.t1959 C10_N_btm.t973 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X643 VSS.t1860 a_18971_44654# a_15730_45670.t0 VSS.t1859 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X644 VDAC_N.t993 C10_N_btm.t972 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X645 VDAC_N.t1957 C8_N_btm.t27 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X646 VDAC_N.t269 C10_N_btm.t971 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X647 VDAC_P.t995 C9_P_btm.t482 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X648 a_17786_46658# a_18064_46642# a_18020_46526# VDD.t1800 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X649 VSS.t3180 VDD.t3162 VSS.t3179 VSS.t3178 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X650 VSS.t2424 VSS.t2425 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X651 VDAC_P.t1961 C10_P_btm.t988 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X652 VDAC_N.t1955 C9_N_btm.t489 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X653 VDAC_P.t511 C10_P_btm.t987 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X654 a_426_47070# a_380_47222# VSS.t1473 VSS.t1472 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X655 VDAC_N.t991 C10_N_btm.t970 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X656 VDAC_N.t1953 C10_N_btm.t969 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X657 VCM.t19 a_3990_30651.t21 C10_P_btm.t7 VSS.t294 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X658 VDD.t1516 a_4061_47044# a_4091_47070# VDD.t1515 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X659 VDAC_P.t1959 C10_P_btm.t986 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X660 a_6793_45776# a_5663_45982# a_6707_45776# VSS.t2598 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X661 VSS.t2482 VSS.t2483 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X662 VDAC_N.t509 C8_N_btm.t11 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X663 VDAC_P.t993 C10_P_btm.t985 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X664 VDAC_P.t1957 C7_P_btm.t122 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X665 VDAC_N.t1951 C7_N_btm.t24 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X666 a_15579_44172# a_8727_47222.t19 VDD.t50 VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X667 a_n2810_43806.t1 a_n2840_43780# VSS.t1586 VSS.t945 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X668 VSS.t3084 VDD.t3130 VSS.t3083 VSS.t3082 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X669 a_8204_45412# a_5419_47258# VSS.t1587 VSS.t993 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X670 VDAC_P.t269 C6_P_btm.t5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X671 a_3470_45982# a_885_44868.t37 a_3470_46232# VDD.t2856 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X672 a_5734_30651.t1 a_9343_42718# VSS.t2268 VSS.t2267 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X673 VDAC_P.t1955 C8_P_btm.t245 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X674 a_7029_44350.t1 a_6491_44716# VDD.t1502 VDD.t1501 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X675 a_8470_44172# a_7393_43806# a_8308_43806# VDD.t1533 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X676 VDAC_P.t991 C10_P_btm.t984 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X677 a_22821_39429# a_22400_42718# VDD.t1805 VDD.t1804 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X678 a_11507_47833# RST_Z.t0 VDD.t2916 VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X679 VSS.t3465 VDD.t3214 VSS.t3464 VSS.t3145 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X680 VDAC_N.t989 C3_N_btm.t5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X681 VSS.t536 a_1203_42692.t23 a_5473_43582# VSS.t535 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X682 VDD.t2798 a_22223_47070# a_20647_31459.t3 VDD.t970 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X683 VDAC_P.t1953 C10_P_btm.t983 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X684 a_6105_44894# a_5939_44894# VDD.t1545 VDD.t1544 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X685 VDAC_N.t1949 C10_N_btm.t968 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X686 VDAC_N.t43 C9_N_btm.t488 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X687 VDAC_N.t1947 C9_N_btm.t487 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X688 VDAC_N.t987 C10_N_btm.t967 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X689 VDAC_N.t1945 C8_N_btm.t240 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X690 VDAC_P.t509 C10_P_btm.t982 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X691 VDD.t1552 a_6951_47070# a_7311_47614# VDD.t1551 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X692 VDAC_P.t1951 C8_P_btm.t243 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X693 VDAC_N.t507 C10_N_btm.t966 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X694 VDD.t1562 a_1123_43780# a_1581_43806.t7 VDD.t1561 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X695 a_10623_47307# a_10428_47338# a_10933_47070# VSS.t2119 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X696 VDAC_N.t1943 C10_N_btm.t965 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X697 w_1375_34946.t13 a_n1732_35090.t10 EN_VIN_BSTR_P.t4 w_1375_34946.t12 sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X698 VDD.t1576 a_18879_43780# a_18866_44172# VDD.t1575 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X699 a_15049_45144# a_9521_45982.t19 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X700 VDAC_N.t985 VSS.t3263 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X701 VSS.t430 a_n690_43494.t23 a_n685_46532# VSS.t429 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X702 VSS.t1644 a_9335_44324# a_9266_44350# VSS.t1643 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X703 VDAC_P.t989 VSS.t3348 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X704 a_12636_45758# a_2424_46794.t5 a_12386_45758# VSS.t2852 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X705 VDAC_P.t1949 C9_P_btm.t481 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X706 VDAC_N.t1941 VSS.t3310 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X707 VDD.t2522 VSS.t3632 VDD.t2521 VDD.t2520 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X708 VDAC_P.t43 C10_P_btm.t981 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X709 a_13273_44868.t7 a_18879_43780# VDD.t1574 VDD.t1573 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X710 VDAC_N.t267 C7_N_btm.t46 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X711 a_7552_46134# a_n53_44363.t15 a_7694_46309# VDD.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X712 VDAC_P.t1947 C6_P_btm.t54 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X713 VDAC_N.t1939 C9_N_btm.t486 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X714 VDAC_P.t987 C7_P_btm.t44 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X715 VDAC_P.t1945 C7_P_btm.t23 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X716 VSS.t3694 C10_P_btm.t18 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X717 VSS.t1202 a_22959_47070# a_21276_30659.t0 VSS.t1201 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X718 VDAC_P.t507 C9_P_btm.t480 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X719 VDAC_P.t1943 C9_P_btm.t479 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X720 VDAC_P.t985 C10_P_btm.t980 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X721 VDAC_P.t1941 C9_P_btm.t478 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X722 VDD.t279 a_n1827_44868.t10 a_n2293_43780# VDD.t278 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X723 VDAC_P.t267 C10_P_btm.t979 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X724 w_1375_34946.t4 a_n1123_35174.t6 w_1375_34946.t4 w_1375_34946.t2 sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X725 VDAC_P.t1939 VSS.t3385 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X726 VSS.t3785 C6_N_btm.t69 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X727 VDAC_N.t983 C10_N_btm.t964 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X728 a_5419_47258# a_6631_44582# VDD.t1446 VDD.t1445 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X729 VDAC_N.t1937 C10_N_btm.t963 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X730 a_1852_45982# a_1735_46195# VSS.t2681 VSS.t2680 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X731 VDD.t1147 a_8391_47044# a_135_43540.t5 VDD.t1146 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X732 VDAC_N.t505 C9_N_btm.t485 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X733 VDAC_N.t1935 C9_N_btm.t484 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X734 a_19520_46500# a_7208_47044# VSS.t2614 VSS.t2613 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X735 VDAC_P.t983 C8_P_btm.t242 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X736 VDAC_N.t981 C10_N_btm.t962 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X737 VDAC_P.t1937 C10_P_btm.t978 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X738 VDAC_P.t505 C10_P_btm.t977 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X739 VDAC_P.t1935 C9_P_btm.t477 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X740 VDAC_N.t1933 C10_N_btm.t961 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X741 VDAC_P.t981 C9_P_btm.t476 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X742 VDAC_N.t147 C10_N_btm.t960 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X743 VDAC_P.t1933 C9_P_btm.t475 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X744 VDAC_P.t147 C8_P_btm.t241 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X745 VSS.t3572 C9_N_btm.t528 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X746 VDAC_P.t1931 C10_P_btm.t976 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X747 VDAC_P.t979 VSS.t3347 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X748 a_15079_46134# a_13248_45956.t17 VSS.t485 VSS.t484 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X749 a_10612_43806# a_1053_45123.t6 a_10362_43806# VSS.t581 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X750 a_18445_42718# a_1203_42692.t29 a_18457_42968# VDD.t485 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X751 VDD.t2330 VSS.t3666 VDD.t2329 VDD.t2328 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X752 VDAC_P.t1929 C10_P_btm.t975 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X753 VDAC_N.t1931 C7_N_btm.t8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X754 a_1123_43780# a_135_43540.t23 VDD.t2862 VDD.t2861 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X755 VSS.t2081 a_5923_31099.t4 a_8423_42718# VSS.t2080 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X756 a_10069_42968# a_7557_43236.t25 a_9987_42968# VDD.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X757 VDD.t345 a_1334_43494.t24 a_1339_43315# VDD.t344 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X758 a_10703_46526# a_10227_47214.t41 VDD.t572 VDD.t571 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X759 VDAC_N.t979 C8_N_btm.t8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X760 C10_P_btm.t1071 a_n4515_30659.t19 VREF.t68 VDD.t3005 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X761 VDAC_N.t1929 C10_N_btm.t959 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X762 VDAC_N.t503 C6_N_btm.t45 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X763 a_3177_44048# a_2959_43806# VSS.t1218 VSS.t1217 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X764 VDAC_N.t1927 C8_N_btm.t239 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X765 VDAC_P.t503 C7_P_btm.t116 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X766 VDAC_P.t1927 C7_P_btm.t115 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X767 VSS.t188 a_135_43540.t43 a_369_45982# VSS.t187 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X768 a_1663_45046# a_1935_44874# a_1893_45144# VDD.t1156 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X769 VDAC_P.t977 C8_P_btm.t240 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X770 VDD.t2325 VSS.t3813 VDD.t2324 VDD.t2323 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X771 VDAC_P.t1925 C10_P_btm.t973 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X772 VDAC_P.t265 C10_P_btm.t972 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X773 a_3055_43806# a_2609_43806# a_2959_43806# VSS.t1225 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X774 VDAC_P.t1923 C9_P_btm.t474 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X775 a_2113_38308# a_1343_38525.t10 VSS.t67 VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X776 VDAC_N.t977 C10_N_btm.t958 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X777 C5_P_btm.t2 a_5734_30651.t6 VCM.t25 VSS.t457 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X778 VDAC_N.t1925 C10_N_btm.t957 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X779 C4_N_btm.t2 EN_VIN_BSTR_N.t20 VIN_N.t12 VSS.t447 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X780 a_6078_44172# a_5001_43806# a_5916_43806# VDD.t1161 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X781 VDAC_N.t265 C10_N_btm.t956 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X782 VDD.t2178 a_4527_43566# a_927_42692.t5 VDD.t2177 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X783 VDAC_N.t1923 C10_N_btm.t955 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X784 VDAC_N.t975 C10_N_btm.t954 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X785 VSS.t1236 a_7595_47614# DATA[5].t3 VSS.t1235 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X786 VDAC_P.t975 C10_P_btm.t971 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X787 VDAC_P.t1921 C10_P_btm.t970 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X788 VDAC_P.t501 C9_P_btm.t473 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X789 VDAC_P.t1919 C9_P_btm.t472 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X790 VDAC_N.t1921 C10_N_btm.t953 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X791 VSS.t141 a_20107_43806# a_2587_44868.t0 VSS.t140 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X792 a_13930_46842# a_13524_46832.t13 a_13937_46602# VDD.t547 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X793 a_21020_30659.t2 a_22591_47070# VDD.t1690 VDD.t1689 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X794 a_3726_37500# a_3754_38470.t3 VDAC_Ni.t5 VSS.t2837 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X795 a_17564_32305.t3 a_22959_43806# VDD.t2074 VDD.t1060 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X796 VDAC_P.t973 C9_P_btm.t471 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X797 VDAC_P.t1917 C10_P_btm.t969 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X798 VSS.t1240 a_n2288_47588# a_n4515_30659.t0 VSS.t1239 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X799 VDAC_N.t501 C9_N_btm.t482 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X800 VDAC_P.t87 C10_P_btm.t968 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X801 VDAC_N.t1919 C6_N_btm.t53 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X802 VSS.t1244 a_13635_43566# a_11455_44576.t1 VSS.t1243 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X803 a_4830_43958.t0 a_9395_47044# VSS.t1252 VSS.t1251 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X804 VSS.t3237 VDD.t3182 VSS.t3236 VSS.t3235 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X805 VDAC_N.t973 C4_N_btm.t16 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X806 VDAC_N.t1917 C7_N_btm.t44 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X807 COMP_P.t6 a_1239_39587# VDD.t1718 VDD.t1717 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X808 VSS.t3534 VDD.t3238 VSS.t3533 VSS.t3532 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X809 VDAC_N.t87 C10_N_btm.t952 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X810 VSS.t3090 VDD.t3132 VSS.t3089 VSS.t3088 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X811 a_15133_43582# a_11455_44576.t23 VSS.t2720 VSS.t2719 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X812 VDAC_N.t1915 C9_N_btm.t481 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X813 VDAC_P.t1915 C8_P_btm.t239 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X814 VDAC_N.t971 C9_N_btm.t480 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X815 a_5626_46846# a_1429_47222.t19 VSS.t390 VSS.t389 sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X816 a_4152_45804# a_4035_45609# VSS.t1258 VSS.t1257 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X817 VSS.t3557 C10_P_btm.t29 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X818 VDAC_P.t971 C9_P_btm.t470 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X819 VDAC_N.t1913 C10_N_btm.t951 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X820 a_2709_43262# a_1334_43494.t18 VDD.t341 VDD.t340 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X821 VSS.t1260 a_16211_44582# a_13715_43780# VSS.t1259 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X822 VDAC_P.t1913 C8_P_btm.t238 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X823 VDAC_P.t499 C9_P_btm.t469 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X824 a_2959_43806# a_2443_43806# a_2864_43806# VSS.t2098 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X825 a_2617_44894# a_2587_44868.t23 VSS.t266 VSS.t265 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X826 VDAC_N.t499 C10_N_btm.t950 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X827 VDAC_P.t1911 C10_P_btm.t964 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X828 VDAC_N.t1911 C10_N_btm.t949 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X829 VSS.t3615 C8_N_btm.t263 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X830 VDAC_N.t969 C10_N_btm.t948 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X831 VDAC_P.t969 C9_P_btm.t468 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X832 VDAC_P.t1909 C10_P_btm.t963 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X833 VDAC_P.t263 C10_P_btm.t962 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X834 VDAC_N.t1909 C10_N_btm.t947 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X835 VDAC_N.t263 C10_N_btm.t946 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X836 a_1343_38525.t1 a_1177_38525# VSS.t2669 VSS.t2668 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X837 a_n2103_44868.t1 a_16670_44324# a_16618_44670# VSS.t1267 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X838 VDD.t1205 a_16111_45412# a_15187_44868# VDD.t1204 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X839 VDAC_N.t1907 C9_N_btm.t479 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X840 VDAC_N.t967 C8_N_btm.t189 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X841 VDAC_N.t1905 C10_N_btm.t945 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X842 a_1617_45554# a_1429_47222.t23 a_1522_45554# VDD.t330 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X843 VDAC_P.t1907 C9_P_btm.t467 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X844 VDAC_P.t967 C9_P_btm.t466 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X845 VDAC_P.t1905 C9_P_btm.t465 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X846 a_12896_47044# a_4908_45956# VSS.t1790 VSS.t1789 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X847 a_7393_46532# a_7227_46532# VSS.t1276 VSS.t1275 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X848 a_10319_45982# a_9803_45982# a_10224_45982# VSS.t2577 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X849 a_7842_44868# a_8192_44874# a_8150_45144# VDD.t2230 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X850 VDAC_P.t497 C4_P_btm.t6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X851 C1_P_btm.t0 EN_VIN_BSTR_P.t23 VIN_P.t4 VSS.t559 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X852 VDD.t1664 a_6091_43780# a_1847_45528.t7 VDD.t1663 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X853 VSS.t1616 a_7311_47614# a_7595_47614# VSS.t1615 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X854 VSS.t2391 VSS.t2392 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X855 VSS.t3278 a_n2810_44894.t7 C10_P_btm.t1075 VSS.t3277 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X856 VSS.t340 a_10227_47214.t19 a_19857_43600# VSS.t339 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X857 VDAC_P.t1903 C10_P_btm.t960 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X858 VSS.t2191 a_11971_46500# a_n237_45454.t1 VSS.t2190 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X859 VDAC_P.t965 C10_P_btm.t959 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X860 a_2674_46348# a_1597_45982# a_2512_45982# VDD.t2680 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X861 a_n2472_45956# a_n2293_45956.t6 VDD.t2953 VDD.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X862 VDAC_N.t497 C3_N_btm.t4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X863 a_18971_44654# a_10227_47214.t39 VDD.t570 VDD.t569 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X864 VSS.t94 a_927_42692.t17 a_768_44670# VSS.t93 sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.08775 ps=0.92 w=0.65 l=0.15
X865 VDAC_P.t1901 C9_P_btm.t464 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X866 VDD.t1215 a_18803_47070# a_18822_46526# VDD.t1214 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X867 VDAC_N.t1903 C10_N_btm.t944 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X868 VSS.t2393 VSS.t2394 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X869 a_18044_43806# a_17515_43806# VDD.t1217 VDD.t1216 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X870 a_12802_43806# a_10227_47214.t27 VSS.t348 VSS.t347 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X871 VDAC_N.t965 C8_N_btm.t12 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X872 VDAC_N.t1901 C10_N_btm.t943 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X873 VDAC_P.t145 C10_P_btm.t958 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X874 VDAC_P.t1899 C7_P_btm.t114 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X875 a_9179_44592# a_9521_45982.t23 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X876 VDAC_P.t963 C10_P_btm.t957 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X877 VDAC_P.t1897 C8_P_btm.t237 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X878 VDAC_N.t145 C8_N_btm.t238 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X879 VDAC_P.t495 C9_P_btm.t463 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X880 a_14757_45982# a_14382_46348# VDD.t1219 VDD.t1218 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X881 a_17763_44868# a_18689_45412# VSS.t1852 VSS.t1851 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X882 VDAC_N.t1899 C10_N_btm.t942 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X883 a_8659_44324# a_8862_44482# VDD.t2739 VDD.t2738 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X884 VDAC_P.t1895 C7_P_btm.t113 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X885 a_n2288_47588# a_n2109_47596.t5 VDD.t380 VDD.t379 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X886 VDAC_P.t961 C10_P_btm.t956 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X887 VDAC_P.t1893 C9_P_btm.t462 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X888 VDAC_P.t261 C10_P_btm.t955 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X889 a_13003_43262# a_10227_47214.t37 VDD.t568 VDD.t567 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X890 VSS.t3721 C10_N_btm.t1061 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X891 VDAC_N.t963 VSS.t3262 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X892 a_20283_43262# a_1203_42692.t19 VSS.t530 VSS.t529 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X893 VDAC_N.t1897 C10_N_btm.t940 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X894 VDAC_N.t495 C9_N_btm.t478 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X895 VDD.t19 VDAC_Ni.t10 a_6886_37412# VSS.t19 sky130_fd_pr__nfet_03v3_nvt ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X896 a_7961_46500# a_7743_46904# VDD.t1229 VDD.t1228 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X897 VDAC_N.t1895 C8_N_btm.t237 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X898 CAL_P.t2 a_22465_38541# VDD.t2796 VDD.t2792 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X899 a_n2497_42870.t1 a_15549_47044.t7 VSS.t2892 VSS.t2891 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X900 VDD.t2344 VSS.t3589 VDD.t2343 VDD.t2342 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X901 VDAC_N.t961 C10_N_btm.t939 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X902 a_8192_44874# a_8423_42718# VDD.t1151 VDD.t1150 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X903 a_5945_46846# a_n237_45454.t11 a_5626_46846# VSS.t474 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X904 VDAC_P.t1891 C9_P_btm.t461 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X905 VDAC_P.t959 C10_P_btm.t954 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X906 VSS.t3528 VDD.t3236 VSS.t3527 VSS.t3526 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X907 VDAC_P.t1889 C10_P_btm.t953 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X908 VSS.t1302 a_284_47222# a_n381_46697# VSS.t1301 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X909 VDAC_P.t493 C9_P_btm.t460 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X910 VDAC_N.t1893 C9_N_btm.t477 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X911 VREF.t51 a_19679_31459.t4 C1_N_btm.t5 VDD.t2975 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X912 VDAC_P.t1887 C9_P_btm.t459 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X913 a_19320_35138# a_18394_35068.t9 VSS.t194 VSS.t193 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X914 a_13464_45758# a_4908_45956# a_13214_45758# VSS.t1793 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X915 VDAC_N.t261 C10_N_btm.t938 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X916 VDAC_P.t957 C7_P_btm.t112 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X917 VDAC_N.t1891 C8_N_btm.t236 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X918 VSS.t1314 a_12623_43780# a_12557_43806# VSS.t1313 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X919 VDAC_P.t1885 C10_P_btm.t952 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X920 a_7735_42692# a_6631_44582# VSS.t1513 VSS.t1512 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X921 VDAC_N.t959 C10_N_btm.t937 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X922 VDAC_N.t1889 C10_N_btm.t936 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X923 VCM.t45 a_134_42718.t6 C0_N_btm.t2 VSS.t2706 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X924 a_3990_30651.t2 a_19187_42718# VDD.t2655 VDD.t2654 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X925 VDD.t2399 VSS.t3598 VDD.t2398 VDD.t2397 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X926 VDAC_P.t57 C10_P_btm.t951 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X927 VDAC_P.t1883 C10_P_btm.t950 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X928 VDD.t599 a_13273_44868.t27 a_15589_44350# VDD.t598 sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X929 VDD.t220 a_7557_43236.t19 a_8651_45962# VDD.t219 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X930 VDAC_N.t493 C10_N_btm.t935 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X931 a_n2661_45956.t0 a_6126_46642# VSS.t1318 VSS.t1317 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X932 VDAC_P.t955 C9_P_btm.t458 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X933 VDAC_N.t1887 C8_N_btm.t235 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X934 VSS.t3628 C8_P_btm.t16 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X935 VDD.t2710 a_7208_47044# a_n2103_45412.t5 VDD.t2709 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X936 VDAC_P.t1881 C10_P_btm.t949 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X937 VDAC_P.t491 C9_P_btm.t457 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X938 VDAC_P.t1879 C9_P_btm.t456 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X939 VDAC_P.t953 C9_P_btm.t455 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X940 a_7743_46904# a_7227_46532# a_7648_46892# VSS.t1274 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X941 a_2332_44670# a_1334_43494.t22 VSS.t404 VSS.t403 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X942 VDAC_P.t1877 C10_P_btm.t948 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X943 a_18394_35068.t0 SMPL.t8 VDD.t3043 VDD.t3042 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X944 a_1334_43494.t5 a_3699_43780# VDD.t1409 VDD.t1408 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X945 VDAC_P.t259 C9_P_btm.t454 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X946 VDAC_N.t957 C10_N_btm.t934 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X947 VDAC_N.t1885 C10_N_btm.t933 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X948 VSS.t463 a_n2109_47596.t6 a_22455_45420# VSS.t462 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X949 VSS.t2848 a_n2103_44868.t11 a_n2293_44868# VSS.t2847 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X950 VDAC_N.t57 C10_N_btm.t932 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X951 VSS.t1324 a_2075_42870# a_2075_42718# VSS.t1323 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X952 VDAC_P.t1875 C10_P_btm.t947 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X953 a_49_46500# a_n169_46904# VDD.t1259 VDD.t1258 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X954 VDAC_P.t951 C10_P_btm.t946 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X955 a_3222_30651.t2 a_21303_42718# VDD.t2698 VDD.t2697 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X956 VSS.t1509 a_6631_44582# a_7415_44466# VSS.t1508 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X957 VDAC_P.t1873 C10_P_btm.t945 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X958 VDAC_P.t489 C9_P_btm.t453 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X959 a_8981_43262# a_6485_44582.t8 VDD.t3011 VDD.t3010 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X960 VDAC_P.t1871 C10_P_btm.t944 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X961 a_16102_47044# a_15871_47614# VDD.t1265 VDD.t1264 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X962 VREF.t35 a_22812_30659.t15 C10_N_btm.t29 VDD.t527 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X963 VSS.t2519 VSS.t2520 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X964 a_3692_43628# a_3165_43262# VDD.t1269 VDD.t1268 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X965 VDD.t2511 VSS.t3725 VDD.t2510 VDD.t2509 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X966 VDD.t1271 a_4812_45816# a_4987_45742# VDD.t1270 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X967 VDAC_N.t1883 C10_N_btm.t931 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X968 VSS.t2832 a_13667_32299.t4 C1_N_btm.t4 VSS.t2831 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X969 a_16758_43628# a_8727_47222.t21 VSS.t55 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X970 VDAC_P.t949 C10_P_btm.t943 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X971 VSS.t61 a_12769_44594.t4 a_12725_44670# VSS.t60 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X972 VDD.t1411 a_3699_43780# a_1334_43494.t6 VDD.t1410 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X973 VSS.t3745 C9_P_btm.t22 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X974 VDAC_P.t1869 C8_P_btm.t236 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X975 a_8912_37509.t11 VDAC_N.t955 a_5700_37509.t5 VDD.t2253 sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X976 VDAC_N.t1881 C5_N_btm.t31 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X977 a_7839_47222# a_n237_45454.t9 VDD.t388 VDD.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X978 VDAC_N.t491 C10_N_btm.t930 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X979 VDD.t2955 a_n2293_45956.t7 a_22087_43244# VDD.t2954 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X980 VDAC_N.t1879 C10_N_btm.t929 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X981 VDAC_N.t953 C9_N_btm.t476 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X982 VSS.t2543 VSS.t2544 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X983 a_15139_47730# a_14766_45596.t6 VSS.t2800 VSS.t2799 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X984 VDD.t1135 a_7552_46134# a_7503_45982# VDD.t1134 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X985 a_14382_46348# a_13524_46832.t21 a_13654_46032# VSS.t609 sky130_fd_pr__nfet_01v8 ad=0.151025 pd=1.285 as=0.1092 ps=1.36 w=0.42 l=0.15
X986 a_19679_31459.t3 a_22959_45446# VDD.t1287 VDD.t1286 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X987 VDAC_N.t1877 C9_N_btm.t475 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X988 VDAC_N.t259 C10_N_btm.t928 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X989 VDAC_P.t143 C10_P_btm.t942 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X990 VDAC_P.t1867 C10_P_btm.t941 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X991 VDAC_P.t947 C10_P_btm.t940 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X992 VDAC_P.t1865 C10_P_btm.t939 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X993 VDAC_N.t1875 C7_N_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X994 VDAC_P.t487 C9_P_btm.t451 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X995 a_10251_45454# a_17951_44868# VSS.t1360 VSS.t1359 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X996 VDAC_N.t951 C10_N_btm.t927 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X997 VDAC_P.t1863 C8_P_btm.t235 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X998 VDAC_N.t1873 C10_N_btm.t926 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X999 a_17153_46846# a_13248_45956.t23 a_16921_46364# VSS.t488 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1000 VDD.t226 a_7557_43236.t23 a_14103_46576# VDD.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.090125 ps=0.995 w=0.42 l=0.15
X1001 VDAC_N.t489 C10_N_btm.t925 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1002 VDAC_P.t945 C10_P_btm.t938 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1003 VDAC_N.t1871 C9_N_btm.t474 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1004 VDD.t1397 a_3165_45982# a_3733_46348# VDD.t1396 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1005 a_n2810_44894.t3 a_n2840_44868# VDD.t1304 VDD.t1303 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1006 VSS.t3758 C10_N_btm.t1062 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1007 VREF.t3 a_n2810_47070.t7 C8_P_btm.t3 VDD.t89 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1008 VDAC_P.t1861 C10_P_btm.t937 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1009 a_12610_44172# a_11533_43806# a_12448_43806# VDD.t1466 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1010 VDAC_P.t257 C1_P_btm.t4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1011 VDAC_N.t949 C9_N_btm.t473 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1012 VDAC_P.t1859 C9_P_btm.t450 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1013 VDD.t1306 a_14647_43494# a_14301_44035# VDD.t1305 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1014 VDAC_N.t1869 VSS.t3318 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1015 a_1581_43806.t1 a_1123_43780# VSS.t1624 VSS.t1623 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1016 VDD.t2442 VSS.t3763 VDD.t2441 VDD.t2440 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1017 a_15839_43640# a_15489_43268# a_15744_43628# VDD.t1645 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1018 VDAC_N.t143 C9_N_btm.t472 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1019 VDD.t2430 VSS.t3668 VDD.t2429 VDD.t2428 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1020 CLK_DATA.t4 a_n2833_47874# VDD.t1309 VDD.t1308 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1021 VDAC_P.t943 C10_P_btm.t936 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1022 VSS.t2924 a_6485_44582.t25 a_9048_45758# VSS.t2923 sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.08775 ps=0.92 w=0.65 l=0.15
X1023 VDAC_N.t1867 C10_N_btm.t923 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1024 VDAC_P.t1857 C9_P_btm.t449 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1025 VDAC_N.t947 C7_N_btm.t42 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1026 VDAC_N.t1865 C10_N_btm.t922 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1027 VDD.t1319 a_n1586_35608# a_n2038_35608# VDD.t1318 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1028 VDAC_P.t485 C10_P_btm.t935 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1029 a_n2833_47874# a_n2497_47846.t4 VSS.t2094 VSS.t2093 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X1030 VDAC_P.t1855 C10_P_btm.t934 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1031 VDAC_N.t487 VSS.t3308 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1032 VDAC_N.t1863 C10_N_btm.t921 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1033 VSS.t453 a_17738_32299.t5 C8_N_btm.t5 VSS.t452 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1034 VSS.t1634 a_18879_43780# a_13273_44868.t2 VSS.t1633 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1035 a_17515_43806# a_17242_43806# VSS.t1393 VSS.t1392 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X1036 VSS.t3623 C10_N_btm.t1063 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1037 VSS.t274 a_2587_44868.t29 a_11529_44670# VSS.t273 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X1038 a_5088_37509.t6 VDAC_P.t941 a_8912_37509.t24 VDD.t2244 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X1039 VSS.t2499 VSS.t2500 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1040 VDAC_N.t945 C10_N_btm.t919 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1041 VSS.t2224 a_1431_47070# a_1203_42692.t0 VSS.t2223 sky130_fd_pr__nfet_01v8 ad=0.20475 pd=1.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X1042 VDAC_N.t1861 C8_N_btm.t234 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1043 VDD.t2099 a_2167_46526# a_2343_47070# VDD.t2098 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1044 VDAC_N.t257 C9_N_btm.t471 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1045 VDAC_N.t1859 C9_N_btm.t470 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1046 a_18971_44654# a_18796_44728# a_19150_44716# VSS.t2684 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1047 VDAC_N.t943 C10_N_btm.t918 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1048 a_16513_43640# a_15323_43268# a_16404_43640# VSS.t1439 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1049 VDAC_P.t1853 C10_P_btm.t933 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1050 VDAC_N.t1857 VSS.t3317 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1051 VDAC_P.t85 C8_P_btm.t232 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1052 VDAC_P.t1851 VSS.t3383 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1053 VDAC_P.t939 C9_P_btm.t448 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1054 a_3692_43628# a_3165_43262# VSS.t1339 VSS.t1338 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1055 VSS.t3197 VDD.t3168 VSS.t3196 VSS.t3085 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1056 VDAC_N.t485 C8_N_btm.t233 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1057 a_15730_45670.t1 a_18971_44654# VSS.t1864 VSS.t1863 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1058 VSS.t2515 VSS.t2516 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1059 VSS.t2974 a_n1925_47044.t5 a_22591_43958# VSS.t2973 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1060 VDAC_P.t1849 C10_P_btm.t932 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1061 a_8483_46830# a_135_43540.t29 VDD.t178 VDD.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1062 VSS.t2315 VSS.t2316 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1063 VDAC_P.t483 C6_P_btm.t26 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1064 a_14757_47614# a_14587_47614# VDD.t1333 VDD.t1332 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1065 VDAC_N.t1855 C9_N_btm.t469 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1066 VDAC_P.t1847 C8_P_btm.t231 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1067 VSS.t1408 a_18766_43236# a_18541_43582# VSS.t1407 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1068 VDAC_P.t937 C8_P_btm.t230 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1069 VDAC_N.t941 C10_N_btm.t917 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1070 VDD.t334 a_1334_43494.t13 a_12931_46348# VDD.t333 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1071 a_17951_44868# a_12127_46744# VDD.t1048 VDD.t1047 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X1072 a_n1732_35090.t5 SMPL.t21 VSS.t2954 VSS.t2953 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1073 a_9898_44350# a_9140_44466# a_9335_44324# VDD.t1050 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1074 VDAC_P.t1845 C10_P_btm.t931 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1075 VDD.t1468 a_12101_44048# a_11991_44172# VDD.t1467 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1076 VDAC_N.t1853 C10_N_btm.t916 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1077 VDAC_P.t255 C8_P_btm.t229 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1078 VSS.t2331 VSS.t2332 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1079 VDAC_P.t1843 C10_P_btm.t930 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1080 VDAC_N.t85 C9_N_btm.t468 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1081 VSS.t3678 C10_P_btm.t20 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1082 VDAC_N.t1851 C10_N_btm.t915 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1083 a_12833_42718# a_10259_42870.t27 VSS.t17 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1084 a_428_42724# a_546_43100# VSS.t1809 VSS.t1808 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1085 VDAC_N.t939 C10_N_btm.t914 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1086 VDAC_P.t935 C10_P_btm.t928 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1087 VDAC_N.t1849 C10_N_btm.t913 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1088 VDAC_N.t483 C9_N_btm.t467 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1089 VDAC_P.t1841 C10_P_btm.t927 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1090 VDAC_N.t1847 C8_N_btm.t232 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1091 VDAC_N.t937 C10_N_btm.t912 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1092 a_15005_47222# a_15329_47044# a_15251_47320# VDD.t1057 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X1093 VDAC_P.t481 C9_P_btm.t447 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1094 VDAC_N.t1845 C8_N_btm.t231 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1095 a_17738_32299.t3 a_22959_44358# VDD.t1061 VDD.t1060 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1096 VDAC_P.t1839 C9_P_btm.t446 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1097 a_18190_46526# a_18064_46642# a_17786_46658# VSS.t1841 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1098 a_571_46830# a_135_43540.t41 VDD.t190 VDD.t189 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1099 VDAC_P.t933 C10_P_btm.t926 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1100 a_18866_44172# a_17789_43806# a_18704_43806# VDD.t1071 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1101 a_n519_46532# a_n685_46532# VSS.t1642 VSS.t1641 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1102 VSS.t1139 a_22223_46534# a_20163_31459.t1 VSS.t1138 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1103 VDAC_N.t255 C8_N_btm.t230 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1104 VDAC_N.t1843 C7_N_btm.t116 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1105 VDAC_N.t935 C10_N_btm.t911 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1106 VSS.t3192 VDD.t3166 VSS.t3191 VSS.t3190 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1107 VDAC_N.t1841 C10_N_btm.t910 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1108 VDAC_P.t1837 C7_P_btm.t111 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1109 VDAC_N.t481 C9_N_btm.t466 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1110 VDAC_P.t141 C7_P_btm.t110 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1111 VDAC_P.t1835 C6_P_btm.t44 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1112 VDAC_N.t1839 C4_N_btm.t17 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1113 VDAC_P.t931 C9_P_btm.t445 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1114 a_18247_46348# a_17623_45982# a_18139_45982# VDD.t1080 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1115 VDAC_P.t1833 C8_P_btm.t228 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1116 VDAC_N.t933 C10_N_btm.t909 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1117 VDAC_P.t479 VSS.t3368 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1118 a_1115_47044# a_n99_45438.t2 VDD.t2044 VDD.t2043 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X1119 VDAC_N.t1837 C9_N_btm.t465 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1120 VSS.t1149 a_3576_44364# a_3328_44324# VSS.t1148 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1121 a_13003_43262# a_12379_43268# a_12895_43640# VDD.t1095 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1122 VDAC_N.t141 C9_N_btm.t464 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1123 VDAC_P.t1831 C10_P_btm.t925 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1124 VDAC_P.t929 C9_P_btm.t444 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1125 VDAC_N.t1835 C10_N_btm.t908 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1126 VDAC_N.t931 C9_N_btm.t463 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1127 VDAC_P.t1829 C10_P_btm.t924 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1128 VDD.t1100 a_7981_45956# a_8011_46309# VDD.t1099 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1129 VDAC_P.t253 C10_P_btm.t923 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1130 a_7557_43236.t7 a_11427_43566# VDD.t1102 VDD.t1101 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1131 VDAC_N.t1833 C10_N_btm.t907 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1132 VDAC_P.t1827 C10_P_btm.t922 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1133 VDAC_N.t479 C10_N_btm.t448 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1134 a_847_45956# a_135_43540.t19 VDD.t2858 VDD.t2857 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1135 VDAC_N.t1831 C10_N_btm.t904 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1136 VDAC_P.t927 C9_P_btm.t443 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1137 VDAC_P.t1825 C10_P_btm.t921 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1138 VDD.t1112 a_18135_47588# a_13524_46832.t3 VDD.t1111 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1139 VDAC_N.t929 C8_N_btm.t229 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1140 VDAC_P.t477 C10_P_btm.t920 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1141 VSS.t3658 C10_N_btm.t1064 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1142 VSS.t3126 VDD.t3144 VSS.t3125 VSS.t3124 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1143 VDD.t449 a_7754_40130.t10 a_8912_37509.t3 VDD.t448 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X1144 a_3437_43268# a_3271_43268# VDD.t2071 VDD.t2070 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1145 VDD.t2475 VSS.t3588 VDD.t2474 VDD.t2473 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1146 a_3883_46904# a_3437_46532# a_3787_46904# VSS.t1871 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1147 VDAC_N.t1829 C9_N_btm.t462 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1148 VDAC_N.t253 C10_N_btm.t902 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1149 VDAC_P.t1823 C8_P_btm.t227 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1150 VSS.t49 a_8727_47222.t17 a_15733_43806# VSS.t48 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1151 a_13991_42883# a_5334_30651.t4 VDD.t3038 VDD.t3037 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1152 VSS.t1876 a_15468_45412# a_11788_46134# VSS.t1875 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X1153 a_1387_45670# a_1659_45528# a_1617_45554# VDD.t1834 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1154 a_16140_44894# a_16074_45046# a_14635_44324# VSS.t1881 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1155 VSS.t1885 a_13023_42718# a_5334_30651.t0 VSS.t1884 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1156 VSS.t1771 a_1239_39587# COMP_P.t2 VSS.t1770 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1157 VDD.t2319 VSS.t3571 VDD.t2318 VDD.t2317 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1158 a_10362_43806# a_10414_43780# a_n1551_44324.t2 VSS.t2576 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1159 VSS.t3422 VDD.t3198 VSS.t3421 VSS.t3420 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1160 a_13725_44350# a_10114_45276.t5 VSS.t157 VSS.t156 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X1161 a_8391_47044# a_8727_47222.t13 VDD.t85 VDD.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X1162 VDAC_N.t1827 C8_N_btm.t228 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1163 VDAC_N.t927 C10_N_btm.t901 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1164 a_3754_39134# a_7754_39300# VSS.t693 sky130_fd_pr__res_high_po_0p35 l=18
X1165 VDD.t1846 a_n268_44582# a_n381_43433# VDD.t1845 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1166 VDD.t2301 VSS.t3701 VDD.t2300 VDD.t2299 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1167 VDAC_P.t925 C10_P_btm.t919 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1168 VDAC_N.t1825 C6_N_btm.t28 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1169 VDAC_N.t477 C8_N_btm.t227 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1170 VDAC_N.t1823 C10_N_btm.t900 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1171 VDAC_P.t1821 C7_P_btm.t109 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1172 VDAC_P.t35 C10_P_btm.t918 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1173 a_5700_37509.t0 VDAC_N.t925 a_8912_37509.t6 VDD.t2254 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1174 VDAC_P.t1819 C6_P_btm.t10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1175 a_11361_43640# a_10171_43268# a_11252_43640# VSS.t2182 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1176 a_15033_46526# a_14658_46526# VDD.t1852 VDD.t1851 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1177 VREF.t24 a_21788_30659.t5 C9_N_btm.t6 VDD.t2052 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1178 a_20405_31459.t1 a_22959_45982# VSS.t1897 VSS.t1353 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1179 VDAC_N.t1821 C10_N_btm.t899 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1180 VDAC_P.t923 C9_P_btm.t442 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1181 VSS.t1905 a_5847_47614# DATA[4].t3 VSS.t1904 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1182 VDD.t1870 a_12436_44868# a_n1741_47596.t2 VDD.t1869 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X1183 VDAC_N.t35 C10_N_btm.t898 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1184 VDAC_P.t1817 C10_P_btm.t917 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1185 a_n2810_46526.t3 a_n2840_46500# VDD.t2256 VDD.t1595 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1186 a_12931_44894# a_4322_46134# VDD.t1782 VDD.t1781 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X1187 VDAC_N.t1819 C8_N_btm.t226 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1188 VDD.t1872 a_2535_45670# a_2151_45670# VDD.t1871 sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X1189 VDAC_P.t475 C9_P_btm.t441 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1190 VSS.t228 a_7557_43236.t21 a_10612_43806# VSS.t227 sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.08775 ps=0.92 w=0.65 l=0.15
X1191 VDAC_N.t923 C10_N_btm.t897 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1192 VDAC_N.t1817 C10_N_btm.t896 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1193 VDAC_N.t475 C10_N_btm.t895 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1194 VDAC_N.t1815 C10_N_btm.t894 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1195 VDAC_P.t1815 C9_P_btm.t440 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1196 VDAC_P.t921 C10_P_btm.t916 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1197 VSS.t1912 a_7754_38470# a_6886_37412# VSS.t1911 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1198 VDD.t2263 VSS.t3691 VDD.t2262 VDD.t2261 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1199 VDAC_N.t921 C10_N_btm.t893 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1200 C10_N_btm.t25 a_22812_30659.t11 VREF.t38 VDD.t523 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1201 a_4651_44350# a_2755_43494.t20 a_4733_44350# VDD.t430 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1202 a_7556_42692# a_7735_42692# VDD.t1399 VDD.t1398 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1203 VSS.t137 a_20107_43806# a_2587_44868.t1 VSS.t136 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1204 VSS.t3555 C4_P_btm.t5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1205 VDAC_P.t1813 C9_P_btm.t439 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1206 VDAC_P.t251 C8_P_btm.t226 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1207 VSS.t1928 a_15221_47044# a_15155_47070# VSS.t1927 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X1208 VDAC_P.t1811 C10_P_btm.t915 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1209 VDAC_P.t919 C10_P_btm.t914 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1210 VDAC_N.t1813 C7_N_btm.t41 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1211 VDAC_N.t251 C2_N_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1212 VDAC_N.t1811 C7_N_btm.t9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1213 VDAC_N.t919 C10_N_btm.t891 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1214 a_2801_42718# a_2587_44868.t27 VSS.t270 VSS.t269 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X1215 VDAC_N.t1809 C10_N_btm.t890 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1216 VDAC_P.t1809 C6_P_btm.t41 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1217 VSS.t356 a_n2661_45420.t6 a_21847_43806# VSS.t355 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1218 a_16145_43806# a_14955_43806# a_16036_43806# VSS.t1931 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1219 VDAC_N.t473 C8_N_btm.t225 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1220 VDD.t2307 VSS.t3673 VDD.t2306 VDD.t2305 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1221 VDAC_P.t473 C10_P_btm.t913 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1222 VDAC_P.t1807 C7_P_btm.t108 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1223 VDAC_N.t1807 C9_N_btm.t461 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1224 SMPL_ON_N.t4 a_21789_35634# VDD.t2761 VDD.t2760 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1225 VDD.t2341 VSS.t3612 VDD.t2340 VDD.t2339 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1226 VSS.t3174 VDD.t3160 VSS.t3173 VSS.t3172 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1227 VDD.t1882 a_22123_44894# a_22591_44894# VDD.t1881 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1228 VDAC_P.t917 C8_P_btm.t225 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1229 VDAC_N.t917 VSS.t3260 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1230 VDAC_P.t1805 C9_P_btm.t438 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1231 VSS.t1779 a_1239_39043# COMP_N.t3 VSS.t1772 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1232 VDAC_N.t1805 C10_N_btm.t889 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1233 a_18139_43806# a_17623_43806# a_18044_43806# VSS.t1938 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1234 VDAC_N.t139 C9_N_btm.t460 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1235 a_n283_35174# a_n1732_35090.t12 VSS.t2736 VSS.t2735 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1236 a_5700_37509.t19 VSS.t3692 VDAC_Pi.t7 VDD.t2452 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1237 VDD.t2084 a_15323_44894# a_1429_47222.t3 VDD.t2083 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1238 a_2113_38308# a_2113_38308# a_2113_38308# VSS.t2633 sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=3.02 ps=24.88 w=1 l=0.15
X1239 VSS.t1944 a_21540_43236# a_13458_32299.t1 VSS.t1943 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1240 VDAC_N.t1803 C10_N_btm.t888 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1241 VSS.t1416 a_4651_47614# DATA[3].t1 VSS.t1415 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1242 VDAC_P.t139 C9_P_btm.t437 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1243 VDAC_P.t1803 C10_P_btm.t912 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1244 VDAC_N.t915 C10_N_btm.t887 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1245 VDAC_N.t1801 VSS.t3315 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1246 VDAC_N.t471 C9_N_btm.t459 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1247 VDAC_P.t915 C10_P_btm.t911 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1248 VSS.t1948 a_17927_46195# a_18530_47070# VSS.t1947 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X1249 a_15393_45982# a_15328_46134# a_14955_45982# VSS.t1503 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1250 VDAC_P.t1801 C10_P_btm.t910 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1251 a_11160_46904# a_10079_46532# a_10813_46500# VDD.t2219 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1252 VDAC_N.t1799 C8_N_btm.t224 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1253 VSS.t3748 C8_N_btm.t264 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1254 VDD.t1778 a_4322_46134# a_4279_46232# VDD.t1777 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1255 VDAC_P.t471 C6_P_btm.t7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1256 a_18493_44716# a_18449_44324# a_18327_44728# VSS.t1953 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1257 VDAC_P.t1799 C7_P_btm.t107 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1258 VSS.t2673 a_1177_38525# a_1343_38525.t2 VSS.t2672 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1259 a_11455_44576.t6 a_13635_43566# VDD.t1182 VDD.t1181 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1260 VDAC_P.t913 C6_P_btm.t23 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1261 a_12651_44576.t4 a_16579_43566# VDD.t1911 VDD.t1910 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1262 a_1412_46794.t1 a_8483_46830# VDD.t1331 VDD.t1330 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1263 a_4247_45816# a_3731_45444# a_4152_45804# VSS.t2152 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1264 VDAC_P.t1797 C10_P_btm.t909 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1265 VDAC_N.t913 C10_N_btm.t886 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1266 VDD.t138 a_20107_43806# a_2587_44868.t7 VDD.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1267 VSS.t422 a_n690_43494.t17 a_7227_46532# VSS.t421 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1268 VDAC_N.t1797 C5_N_btm.t4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1269 VDD.t1917 a_16057_43236# a_15947_43262# VDD.t1916 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1270 VDAC_N.t249 C10_N_btm.t885 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1271 a_1847_45528.t6 a_6091_43780# VDD.t1658 VDD.t1657 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1272 VSS.t2357 VSS.t2358 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1273 VSS.t1926 a_7556_42692# a_5923_31099.t1 VSS.t1925 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1274 a_19857_43600# a_16475_45412# a_19771_43600# VSS.t1747 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1275 VSS.t3404 VDD.t3192 VSS.t3403 VSS.t3402 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1276 VDAC_N.t1795 C7_N_btm.t110 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1277 VDD.t2433 VSS.t3578 VDD.t2432 VDD.t2431 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1278 VDAC_N.t911 C10_N_btm.t884 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1279 VDAC_P.t249 C7_P_btm.t106 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1280 a_17613_44894# a_14204_44350# a_17531_44894# VSS.t1969 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1281 a_4927_47070# a_n2497_47846.t5 a_4833_47070# VSS.t2095 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1282 VDAC_P.t1795 C8_P_btm.t224 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1283 VDAC_N.t1793 C9_N_btm.t458 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1284 VDAC_P.t911 C10_P_btm.t908 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1285 VDAC_P.t1793 C8_P_btm.t223 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1286 VDAC_P.t469 C9_P_btm.t436 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1287 VDAC_N.t469 C10_N_btm.t883 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1288 VSS.t1973 a_10415_47846# a_9517_46539# VSS.t1972 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1289 VDD.t390 a_n237_45454.t10 a_83_45776# VDD.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1290 a_5700_37509.t7 VDAC_N.t1791 a_8912_37509.t13 VDD.t2249 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1291 VSS.t3168 VDD.t3158 VSS.t3167 VSS.t3166 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1292 a_2655_42870# a_1334_43494.t14 a_2801_42968# VDD.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1293 VDAC_N.t909 C9_N_btm.t457 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1294 VDAC_P.t1791 C10_P_btm.t907 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1295 VDAC_N.t1789 C10_N_btm.t882 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1296 VDAC_P.t909 C10_P_btm.t906 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1297 VDD.t2735 a_9179_44592# a_9140_44466# VDD.t2734 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1298 VDAC_P.t1789 C10_P_btm.t905 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1299 VDAC_P.t83 C8_P_btm.t222 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1300 VDAC_N.t83 C10_N_btm.t881 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1301 VDAC_N.t1787 C8_N_btm.t222 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1302 a_1334_43494.t1 a_3699_43780# VSS.t1479 VSS.t1478 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1303 C3_P_btm.t2 a_n2442_43262.t4 VSS.t127 VSS.t126 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1304 a_8727_47222.t0 a_11143_47588# VSS.t1445 VSS.t1444 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1305 a_22087_43244# a_n2293_45956.t8 VSS.t2857 VSS.t2856 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1306 VDAC_N.t907 C7_N_btm.t109 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1307 a_22465_38541# a_22775_42718# VSS.t2692 VSS.t2691 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X1308 VDD.t1056 a_428_42724# a_n2293_45420.t2 VDD.t1055 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X1309 VDAC_P.t1787 C6_P_btm.t55 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1310 VDAC_P.t907 C10_P_btm.t904 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1311 a_4322_46134# a_4527_46830# VSS.t1805 VSS.t1804 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1312 VDAC_N.t1785 C9_N_btm.t456 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1313 a_16404_43640# a_15489_43268# a_16057_43236# VSS.t1702 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1314 VSS.t3764 C8_P_btm.t15 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1315 a_n2497_42870.t7 a_13273_44868.t25 VSS.t648 VSS.t647 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1316 VDAC_P.t1785 C10_P_btm.t903 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1317 a_1522_44466# a_927_42692.t15 VDD.t98 VDD.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X1318 VDAC_P.t467 C10_P_btm.t902 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1319 VDAC_P.t1783 C9_P_btm.t435 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1320 VDAC_N.t467 C5_N_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1321 VDAC_N.t1783 C9_N_btm.t455 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1322 VDD.t1795 a_11692_46134# a_11248_47319# VDD.t1794 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1323 VDAC_P.t905 C9_P_btm.t434 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1324 a_7648_43806# a_7319_43262# VDD.t1931 VDD.t1930 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1325 VSS.t2434 VSS.t2435 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1326 VDAC_N.t905 C7_N_btm.t108 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1327 VDAC_N.t1781 C8_N_btm.t221 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1328 VDAC_P.t1781 C10_P_btm.t901 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1329 VDAC_N.t247 C10_N_btm.t880 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1330 a_7347_43494# a_6485_44582.t19 a_7493_43262# VDD.t3019 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1331 a_11322_46526# a_10245_46532# a_11160_46904# VDD.t789 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1332 VDAC_P.t247 C9_P_btm.t433 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1333 VDAC_N.t1779 C10_N_btm.t879 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1334 VDD.t1936 a_560_45670# a_n105_46195# VDD.t1935 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1335 VDAC_P.t1779 VSS.t3388 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1336 VDAC_N.t903 C10_N_btm.t878 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1337 a_11414_43262# a_10337_43268# a_11252_43640# VDD.t1940 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1338 VDAC_N.t1777 C9_N_btm.t454 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1339 VDAC_P.t903 C10_P_btm.t900 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1340 VDAC_P.t1777 C9_P_btm.t432 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1341 VDAC_N.t465 C9_N_btm.t453 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1342 VDAC_P.t465 C10_P_btm.t899 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1343 VDAC_P.t1775 C9_P_btm.t431 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1344 VDAC_P.t901 C9_P_btm.t430 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1345 VDD.t1327 a_22591_43958# a_22591_43806# VDD.t1326 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1346 VSS.t418 a_n690_43494.t11 a_3271_46532# VSS.t417 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1347 VDD.t1600 a_15192_46500# a_15113_47222# VDD.t1599 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1348 VDAC_P.t1773 C9_P_btm.t429 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1349 VDAC_P.t137 C9_P_btm.t428 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1350 VDAC_N.t1775 C10_N_btm.t877 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1351 VREF.t62 a_n4515_30659.t13 C10_P_btm.t1065 VDD.t2999 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1352 VDD.t2555 VSS.t3552 VDD.t2554 VDD.t2553 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1353 a_9266_44350# a_9140_44466# a_8862_44482# VSS.t1111 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1354 VDAC_P.t1771 C10_P_btm.t897 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1355 VDAC_P.t899 C10_P_btm.t896 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1356 VDAC_N.t901 C9_N_btm.t452 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1357 VDD.t1654 a_7276_45670# a_7016_46231# VDD.t1653 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1358 VDAC_N.t1773 C10_N_btm.t876 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1359 VDAC_N.t137 C10_N_btm.t875 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1360 a_1736_39587.t1 a_1736_39043.t4 a_2112_39137# VSS.t515 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1361 VDAC_N.t1771 C10_N_btm.t874 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1362 a_18282_45670# a_15730_45670.t21 VDD.t498 VDD.t497 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1363 VDAC_P.t1769 C10_P_btm.t895 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1364 DATA[0].t3 a_n1085_47874# VSS.t2000 VSS.t1999 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X1365 a_7142_47070# a_885_44868.t39 VSS.t2770 VSS.t2769 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1366 VDAC_N.t899 C10_N_btm.t873 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1367 VDAC_P.t463 C9_P_btm.t427 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1368 a_999_47846# a_1209_47588# VSS.t2008 VSS.t2007 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1369 VDAC_N.t1769 C6_N_btm.t29 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1370 VDAC_N.t463 C8_N_btm.t220 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1371 a_22455_45420# a_n2109_47596.t7 VSS.t465 VSS.t464 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1372 VDAC_N.t1767 C8_N_btm.t219 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1373 VDAC_P.t1767 C7_P_btm.t105 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1374 a_n331_42718.t0 a_n501_42718# VSS.t2012 VSS.t2011 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1375 VDAC_N.t897 C7_N_btm.t107 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1376 VDAC_P.t897 C6_P_btm.t11 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1377 a_13878_32299.t1 a_21908_43236# VSS.t2016 VSS.t2015 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1378 VSS.t2869 a_12651_44576.t19 a_15877_44670# VSS.t2868 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1379 a_22521_40491# EN_COMP.t5 VDD.t2929 VDD.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1380 VDAC_P.t1765 C8_P_btm.t220 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1381 VSS.t2018 a_9947_47044# a_7208_47044# VSS.t2017 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X1382 a_17786_46658# a_18103_46768# a_18061_46892# VSS.t1839 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1383 VSS.t2938 COMP_N.t8 a_n501_42718# VSS.t2937 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1384 C6_N_btm.t72 a_5542_30651.t5 VCM.t51 VSS.t2833 sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1385 C10_P_btm.t1067 a_n4515_30659.t15 VREF.t64 VDD.t3001 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1386 VDAC_P.t245 C10_P_btm.t893 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1387 VDD.t1972 a_6519_43494# a_6243_45107# VDD.t1971 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X1388 a_10173_45144# a_10114_45276.t6 a_10078_45144# VDD.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X1389 VDAC_N.t1765 C4_N_btm.t9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1390 VDD.t295 a_10227_47214.t21 a_9947_47044# VDD.t294 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1391 a_22465_38541# a_22775_42718# VDD.t2787 VDD.t2786 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1392 VSS.t2491 VSS.t2492 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1393 VDAC_P.t1763 C10_P_btm.t892 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1394 a_n2103_45412.t1 a_18970_45412# VDD.t1978 VDD.t1977 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1395 VDAC_N.t245 C9_N_btm.t451 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1396 VDAC_N.t1763 C9_N_btm.t450 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1397 VDAC_N.t895 C10_N_btm.t872 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1398 a_4987_45742# a_135_43540.t39 VDD.t188 VDD.t187 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1399 VDD.t2586 VSS.t3595 VDD.t2585 VDD.t2584 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1400 VDAC_P.t895 C10_P_btm.t891 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1401 VDAC_P.t1761 C10_P_btm.t890 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1402 a_1387_44582# a_927_42692.t13 VSS.t92 VSS.t91 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1403 a_9395_47044# a_9551_47203# VDD.t1982 VDD.t1981 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X1404 VDAC_P.t461 C10_P_btm.t889 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1405 VDAC_P.t1759 C9_P_btm.t426 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1406 VSS.t3549 VDD.t3243 VSS.t3548 VSS.t3547 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1407 DATA[0].t6 a_n1085_47874# VDD.t1954 VDD.t1953 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1408 VDAC_N.t1761 C10_N_btm.t871 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1409 VDAC_N.t461 C9_N_btm.t449 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1410 a_7557_43236.t4 a_11427_43566# VDD.t1104 VDD.t1103 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1411 VDAC_N.t1759 C10_N_btm.t870 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1412 VDD.t1741 a_4908_45956# a_n1827_45412.t5 VDD.t1740 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1413 VDAC_P.t893 VSS.t3353 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1414 a_4791_42883# a_4000_42718.t5 VSS.t296 VSS.t295 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1415 VDD.t1986 a_17671_42883# a_16824_45276# VDD.t1985 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1416 VDD.t2633 VSS.t3562 VDD.t2632 VDD.t2631 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1417 VSS.t2089 a_1651_47044.t2 a_1431_47070# VSS.t2088 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.08775 ps=0.92 w=0.65 l=0.15
X1418 VDAC_P.t1757 C10_P_btm.t888 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1419 a_n2103_43780.t5 a_3882_44324# a_3830_44670# VSS.t2040 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1420 VDAC_N.t893 C5_N_btm.t29 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1421 VDAC_P.t55 C8_P_btm.t219 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1422 VDD.t1995 a_3541_42718# a_3823_42718# VDD.t1994 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1423 VSS.t1346 a_7839_47222# a_7760_45956# VSS.t1345 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1424 a_16287_45744# a_16475_45412# VDD.t1692 VDD.t1691 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X1425 C8_N_btm.t275 a_21276_30659.t7 VREF.t50 VDD.t2933 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1426 VDAC_N.t1757 C8_N_btm.t217 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1427 VDAC_P.t1755 C6_P_btm.t56 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1428 VDD.t2002 a_2351_47614# DATA[2].t4 VDD.t2001 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1429 VDAC_P.t891 C7_P_btm.t104 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1430 VDAC_N.t55 C9_N_btm.t448 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1431 VDAC_P.t1753 C10_P_btm.t887 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1432 VDD.t2972 a_12651_44576.t23 a_16427_44894# VDD.t2971 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X1433 VDAC_P.t459 C9_P_btm.t425 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1434 VDAC_P.t1751 C9_P_btm.t424 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1435 VDAC_P.t889 C10_P_btm.t886 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1436 VDD.t1958 a_1209_47588# a_999_47846# VDD.t1957 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1437 VDAC_P.t1749 C10_P_btm.t885 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1438 a_14014_46842# a_10259_42870.t21 VSS.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1439 VDAC_N.t1755 C9_N_btm.t447 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1440 VSS.t2472 VSS.t2473 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1441 VDD.t1964 a_21908_43236# a_13878_32299.t3 VDD.t1963 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1442 VDAC_P.t243 C10_P_btm.t884 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1443 VDAC_N.t891 C10_N_btm.t869 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1444 a_11160_46904# a_10245_46532# a_10813_46500# VSS.t1984 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1445 a_1488_43236# a_1339_43315# a_1784_43378# VDD.t2142 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1446 VDAC_N.t1753 C9_N_btm.t446 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1447 a_2216_46758# a_82_45670# a_2358_46565# VDD.t1628 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1448 VDAC_N.t459 C10_N_btm.t868 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1449 VDAC_N.t1751 C10_N_btm.t867 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1450 a_5256_43806# a_5139_44019# VDD.t2013 VDD.t2012 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1451 VSS.t608 a_13524_46832.t19 a_15328_46134# VSS.t607 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1452 VDAC_N.t889 C10_N_btm.t866 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1453 a_11252_43640# a_10337_43268# a_10905_43236# VSS.t1990 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1454 VDD.t2015 a_12887_47833# a_9551_47203# VDD.t2014 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1455 VDAC_N.t1749 C9_N_btm.t445 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1456 VDAC_P.t1747 C10_P_btm.t883 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1457 VDD.t2017 a_5896_45670# a_5749_47222# VDD.t2016 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1458 VDAC_P.t887 C9_P_btm.t423 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1459 VDAC_P.t1745 C8_P_btm.t218 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1460 a_12887_47833# CLK.t0 VDD.t3060 VDD.t3059 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1461 VIN_N.t1 EN_VIN_BSTR_N.t16 C3_N_btm.t0 VSS.t445 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1462 VDAC_P.t457 C10_P_btm.t882 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1463 VSS.t2456 VSS.t2457 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1464 VDAC_P.t1743 C10_P_btm.t881 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1465 VDAC_N.t243 C7_N_btm.t106 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1466 a_6126_46642# a_5382_44582# VSS.t2073 VSS.t2072 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1467 VDAC_N.t1747 C10_N_btm.t865 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1468 VDAC_N.t887 C10_N_btm.t864 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1469 VDAC_P.t885 C7_P_btm.t103 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1470 VDAC_N.t1745 C3_N_btm.t7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1471 VDD.t2338 VSS.t3734 VDD.t2337 VDD.t2336 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1472 VDAC_N.t457 C8_N_btm.t216 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1473 VDAC_P.t1741 C8_P_btm.t217 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1474 VSS.t172 a_135_43540.t27 a_2209_45982# VSS.t171 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1475 VDAC_N.t1743 C10_N_btm.t863 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1476 a_n2497_42870.t3 a_15730_45670.t15 a_18541_43582# VSS.t571 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1477 a_22591_43958# a_n1925_47044.t6 VSS.t2976 VSS.t2975 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1478 a_15309_45438# a_14953_45554# VDD.t2029 VDD.t2028 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1479 VDAC_N.t885 C8_N_btm.t215 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1480 VDAC_Ni.t2 VSS.t3649 a_5088_37509.t1 VDD.t2646 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1481 VDAC_P.t135 C7_P_btm.t102 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1482 VDAC_P.t1739 C10_P_btm.t880 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1483 VDD.t1588 a_12121_45956# a_12151_46309# VDD.t1587 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1484 VDAC_P.t883 C8_P_btm.t216 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1485 VDAC_N.t1741 C9_N_btm.t444 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1486 VDAC_P.t1737 C9_P_btm.t422 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1487 VDAC_N.t135 C9_N_btm.t443 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1488 VDAC_P.t455 C9_P_btm.t421 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1489 a_284_47222# a_85_47070# a_426_47070# VSS.t2079 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1490 VSS.t2591 a_22521_39947# a_22469_39973# VSS.t1537 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1491 VSS.t2071 a_5382_44582# a_5387_44403# VSS.t2070 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1492 VDAC_P.t1735 C10_P_btm.t879 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1493 VDAC_N.t1739 C10_N_btm.t862 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1494 VDAC_N.t883 C10_N_btm.t861 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1495 VSS.t3611 C10_P_btm.t13 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1496 a_5063_45982# a_3165_45982# a_4700_46134# VSS.t1464 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1497 a_n2293_46508.t1 a_7842_44868# VSS.t1536 VSS.t1535 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.18525 ps=1.87 w=0.65 l=0.15
X1498 VDAC_P.t881 C10_P_btm.t878 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1499 VDAC_N.t1737 C10_N_btm.t860 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1500 VDAC_N.t455 C10_N_btm.t859 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1501 VDAC_N.t1735 C10_N_btm.t858 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1502 a_16036_43806# a_15121_43806# a_15689_44048# VSS.t918 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1503 a_15961_47980# a_15691_47614# a_15871_47614# VSS.t919 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X1504 a_18759_42746# a_1581_43806.t18 VDD.t2910 VDD.t2909 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1505 VDAC_P.t1733 C9_P_btm.t420 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1506 VDAC_P.t241 C10_P_btm.t877 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1507 VDAC_N.t881 C9_N_btm.t442 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1508 VDAC_P.t1731 C8_P_btm.t215 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1509 VDAC_N.t1733 C10_N_btm.t857 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1510 a_11335_46830# a_11160_46904# a_11514_46892# VSS.t1952 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1511 VSS.t925 a_22223_42718# a_22400_42718# VSS.t924 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1512 a_6455_44894# a_5939_44894# a_6360_44894# VSS.t1607 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1513 EN_VIN_BSTR_N.t6 VDD.t3188 a_19320_35138# VSS.t3251 sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.9
X1514 VDAC_P.t879 C9_P_btm.t419 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1515 VDAC_N.t241 C10_N_btm.t856 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1516 VSS.t1429 a_14950_43958# a_17623_43806# VSS.t1428 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1517 VDAC_P.t1729 C10_P_btm.t876 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1518 VSS.t1435 a_14950_43958# a_15323_43268# VSS.t1434 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1519 VDAC_N.t1731 C9_N_btm.t441 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1520 VSS.t2963 a_n2661_47044.t4 a_22031_45438# VSS.t2962 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1521 VDAC_N.t879 C6_N_btm.t61 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1522 VDAC_P.t453 C10_P_btm.t875 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1523 VDAC_N.t1729 C5_N_btm.t15 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1524 a_11186_47436# a_10467_47212# a_10623_47307# VSS.t2170 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1525 VDAC_P.t1727 C10_P_btm.t874 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1526 VDAC_N.t453 C10_N_btm.t855 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1527 a_1852_45982# a_1735_46195# VDD.t2779 VDD.t2778 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1528 VSS.t3581 C4_N_btm.t20 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1529 VDAC_N.t1727 C10_N_btm.t854 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1530 VDAC_N.t877 C10_N_btm.t853 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1531 VSS.t402 a_1334_43494.t21 a_12931_45982# VSS.t401 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1532 VDAC_N.t1725 C9_N_btm.t440 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1533 VDAC_P.t877 C8_P_btm.t214 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1534 VDAC_N.t81 C9_N_btm.t439 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1535 VDAC_P.t1725 C10_P_btm.t873 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1536 VDD.t876 a_104_42692# a_134_42718.t2 VDD.t875 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1537 VDAC_P.t81 C10_P_btm.t872 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1538 VDAC_P.t1723 C9_P_btm.t418 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1539 VDAC_P.t875 C10_P_btm.t871 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1540 VDAC_N.t1723 C9_N_btm.t438 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1541 VDAC_P.t1721 C8_P_btm.t213 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1542 a_n2840_44324# a_n2661_44332# VSS.t2172 VSS.t905 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1543 VDAC_P.t451 C10_P_btm.t870 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1544 a_479_43806# a_33_43806# a_383_43806# VSS.t939 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1545 VDAC_P.t1719 C10_P_btm.t869 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1546 VDAC_N.t875 C10_N_btm.t852 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1547 VDAC_P.t873 C10_P_btm.t429 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1548 VDAC_N.t1721 C10_N_btm.t851 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1549 VDAC_N.t451 C10_N_btm.t850 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1550 VDAC_P.t1717 C9_P_btm.t417 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1551 a_n2442_45982.t3 a_n2472_45956# VDD.t1454 VDD.t1453 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1552 a_n2810_43262.t1 a_n2840_43236# VSS.t946 VSS.t945 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1553 VDAC_N.t1719 C10_N_btm.t849 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1554 VDAC_N.t873 C8_N_btm.t214 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1555 VDAC_N.t1717 C9_N_btm.t437 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1556 VDAC_N.t239 C10_N_btm.t848 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1557 VDAC_P.t239 C10_P_btm.t866 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1558 a_n749_47846# a_n447_47044# VSS.t948 VSS.t947 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1559 VSS.t596 a_n1459_43236.t11 a_n1429_43262# VSS.t595 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1560 a_17789_45982# a_17623_45982# VSS.t1141 VSS.t1140 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1561 VSS.t2387 VSS.t2388 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1562 VDAC_P.t1715 C5_P_btm.t6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1563 a_5839_47070# a_5749_47222# VDD.t2021 VDD.t2020 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1564 VDD.t1942 a_22591_43806# a_14409_32299.t3 VDD.t1941 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1565 VDAC_N.t1715 C10_N_btm.t847 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1566 C2_P_btm.t0 a_n2442_45982.t4 VREF.t70 VDD.t3058 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1567 a_9208_43494# a_9416_43530# a_9350_43628# VSS.t1504 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1568 VSS.t627 a_10227_47214.t35 a_18493_44716# VSS.t626 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1569 VDAC_P.t871 C10_P_btm.t865 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1570 VSS.t268 a_2587_44868.t25 a_19358_43582# VSS.t267 sky130_fd_pr__nfet_01v8 ad=0.258375 pd=1.445 as=0.091 ps=0.93 w=0.65 l=0.15
X1571 VDAC_N.t871 C7_N_btm.t105 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1572 VDD.t908 a_8483_43780# a_6485_44582.t7 VDD.t907 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1573 a_4322_46134# a_4527_46830# VSS.t1803 VSS.t1802 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1574 VDAC_P.t1713 C10_P_btm.t864 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1575 VDD.t874 a_22031_45438# a_22959_44358# VDD.t873 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1576 VDAC_P.t449 C10_P_btm.t863 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1577 a_13266_45412# a_13144_47452.t3 VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.17575 ps=1.395 w=0.42 l=0.15
X1578 VDAC_N.t1713 C7_N_btm.t104 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1579 VDAC_N.t449 C10_N_btm.t846 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1580 VDAC_N.t1711 C10_N_btm.t845 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1581 VDAC_P.t1711 C10_P_btm.t862 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1582 VDD.t917 a_6631_42883# a_5784_44364# VDD.t246 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1583 VSS.t159 a_10114_45276.t7 a_12427_46758# VSS.t158 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1584 VDAC_N.t869 C10_N_btm.t844 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1585 C9_P_btm.t8 a_n2467_30659.t7 VREF.t14 VDD.t580 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1586 VIN_P.t14 EN_VIN_BSTR_P.t19 a_n1123_35174.t1 VSS.t560 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1587 VDAC_N.t1709 C9_N_btm.t436 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1588 VDAC_P.t869 C10_P_btm.t861 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1589 VSS.t1903 a_5847_47614# DATA[4].t0 VSS.t1902 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1590 VDAC_P.t1709 C10_P_btm.t860 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1591 a_9969_45982# a_9803_45982# VDD.t2671 VDD.t2670 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1592 VDAC_P.t133 C8_P_btm.t212 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1593 VSS.t2824 a_7029_44350.t2 a_14011_44670# VSS.t2823 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X1594 a_5382_44582# a_4987_45742# VDD.t1275 VDD.t1274 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1595 VDAC_P.t1707 C7_P_btm.t101 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1596 a_n1741_47596.t3 a_12436_44868# VDD.t1868 VDD.t1867 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X1597 a_3754_39134# a_7754_38968# VSS.t693 sky130_fd_pr__res_high_po_0p35 l=18
X1598 VSS.t2377 VSS.t2378 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1599 a_1026_45982# a_135_43540.t37 VSS.t180 VSS.t179 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1600 VDAC_N.t133 VSS.t3293 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1601 a_18449_44324# a_18231_44728# VDD.t921 VDD.t920 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1602 VDAC_N.t1707 C10_N_btm.t843 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1603 VDD.t1933 a_7347_43494# a_7319_43262# VDD.t1932 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X1604 VSS.t980 a_3320_46134# a_2535_45670# VSS.t979 sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
X1605 VSS.t3776 C2_P_btm.t4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1606 VDD.t2129 a_8204_45412# a_n2103_44324.t3 VDD.t2128 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X1607 a_7363_47070# a_5663_45982# a_7000_47222# VSS.t2595 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1608 VDD.t3051 SMPL.t17 a_18394_35068.t5 VDD.t3050 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1609 a_8862_44482# a_9179_44592# a_9137_44716# VSS.t2643 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1610 VSS.t209 a_4830_43958.t13 sky130_fd_pr__diode_pw2nd_05v5 perim=2.64e+06 area=4.347e+11
X1611 VDAC_N.t867 C10_N_btm.t842 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1612 VDD.t35 a_9521_45982.t17 a_12379_43268# VDD.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1613 VSS.t3679 C10_P_btm.t12 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1614 SMPL.t4 a_n2833_42692# VDD.t926 VDD.t925 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1615 VDAC_N.t1705 C10_N_btm.t841 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1616 VDAC_P.t867 C9_P_btm.t416 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1617 VDD.t1365 a_14950_43958# a_17623_43806# VDD.t1364 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1618 VDAC_P.t1705 C10_P_btm.t858 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1619 a_n1741_42692# a_n1735_43236.t11 VDD.t608 VDD.t607 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1620 VDAC_P.t447 C10_P_btm.t857 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1621 VSS.t982 a_7000_47222# a_6951_47070# VSS.t981 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1622 a_885_44868.t4 a_4322_46134# a_4703_44894# VSS.t1817 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1623 VDAC_P.t1703 C9_P_btm.t415 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1624 VDAC_P.t865 C9_P_btm.t414 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1625 VDAC_P.t1701 C10_P_btm.t856 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1626 VSS.t3047 VDD.t3117 VSS.t3046 VSS.t3045 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1627 VSS.t108 a_n2293_46508.t7 a_22031_44350# VSS.t107 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1628 VSS.t3627 C8_N_btm.t266 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1629 VDAC_N.t447 C10_N_btm.t840 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1630 a_3754_38802# a_7754_38968# VSS.t693 sky130_fd_pr__res_high_po_0p35 l=18
X1631 VDAC_N.t1703 C10_N_btm.t839 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1632 VDAC_N.t865 C10_N_btm.t838 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1633 a_3177_44048# a_2959_43806# VDD.t1153 VDD.t1152 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1634 a_15688_45758# a_13273_44868.t31 VSS.t655 VSS.t654 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X1635 VDAC_P.t237 C10_P_btm.t855 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1636 VDAC_N.t1701 C10_N_btm.t837 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1637 a_21847_43806# a_n2661_45420.t7 VSS.t358 VSS.t357 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1638 a_8379_46134# a_8651_45962# a_8609_46232# VDD.t1246 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1639 VDAC_N.t237 C8_N_btm.t212 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1640 VDAC_P.t1699 C9_P_btm.t413 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1641 VDAC_P.t863 C8_P_btm.t211 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1642 VDD.t2759 a_21789_35634# SMPL_ON_N.t6 VDD.t2758 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1643 VDAC_P.t1697 C9_P_btm.t412 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1644 VDAC_N.t1699 C10_N_btm.t836 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1645 VDAC_P.t445 C9_P_btm.t411 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1646 COMP_N.t2 a_1239_39043# VSS.t1778 VSS.t1766 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1647 VSS.t31 a_9521_45982.t11 a_10171_43268# VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1648 VDAC_P.t1695 C10_P_btm.t854 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1649 a_5715_45956# a_5918_46234# VDD.t938 VDD.t937 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1650 VDD.t163 a_1412_46794.t6 a_7839_47222# VDD.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1651 VSS.t1683 a_847_45956# a_781_45982# VSS.t1682 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1652 a_22123_44894# a_n2293_47044.t5 VDD.t468 VDD.t467 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1653 VSS.t598 a_n1459_43236.t12 a_22959_44894# VSS.t597 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1654 VDAC_N.t863 C8_N_btm.t211 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1655 VSS.t2531 VSS.t2532 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1656 VDAC_P.t861 C7_P_btm.t100 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1657 VDAC_N.t1697 C6_N_btm.t11 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1658 VSS.t1358 a_17951_44868# a_10251_45454# VSS.t1357 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X1659 a_11788_43806# a_11671_44019# VDD.t944 VDD.t943 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1660 VDAC_P.t1693 C10_P_btm.t853 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1661 a_5001_43806# a_4835_43806# VSS.t1004 VSS.t1003 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1662 VDAC_N.t445 C10_N_btm.t835 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1663 a_4080_44670# a_3165_45982# a_3830_44670# VSS.t1467 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1664 VDAC_P.t41 VSS.t3376 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1665 VDD.t136 a_20107_43806# a_2587_44868.t4 VDD.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1666 VDD.t1598 a_n2840_45956# a_n2810_45982.t3 VDD.t1597 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1667 a_15037_46232# a_14573_47070# a_14955_45982# VDD.t949 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1668 VDAC_N.t1695 C10_N_btm.t834 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1669 VDAC_N.t861 C10_N_btm.t412 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1670 VDAC_N.t1693 C10_N_btm.t833 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1671 VDAC_P.t1691 C10_P_btm.t852 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1672 VDD.t934 a_22031_44350# a_22959_43270# VDD.t933 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1673 VDAC_P.t859 C10_P_btm.t851 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1674 VDAC_N.t41 C10_N_btm.t832 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1675 a_7743_43806# a_7227_43806# a_7648_43806# VSS.t1011 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1676 VDAC_P.t1689 C9_P_btm.t410 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1677 VDAC_P.t443 C8_P_btm.t210 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1678 VDAC_N.t1691 C10_N_btm.t831 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1679 VDD.t2064 a_19520_46500# a_n2109_47596.t3 VDD.t2063 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X1680 a_10415_45982# a_9969_45982# a_10319_45982# VSS.t1551 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1681 VSS.t3603 C9_N_btm.t526 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1682 VDAC_N.t859 C10_N_btm.t830 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1683 a_9943_45046# a_10215_44874# a_10173_45144# VDD.t956 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1684 VDAC_N.t1689 C10_N_btm.t829 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1685 VDAC_N.t443 C9_N_btm.t434 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1686 a_5923_31099.t0 a_7556_42692# VSS.t1924 VSS.t1923 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1687 a_12725_44670# a_12651_44576.t27 a_12379_44350# VSS.t2887 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1688 VDAC_N.t1687 C10_N_btm.t828 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1689 VDAC_P.t1687 C10_P_btm.t850 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1690 a_1736_39587.t0 a_1736_39043.t5 VDD.t465 VDD.t464 sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X1691 VDAC_N.t857 C10_N_btm.t827 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1692 VDAC_N.t1685 C10_N_btm.t826 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1693 VDAC_P.t857 C10_P_btm.t849 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1694 VDAC_P.t1685 C10_P_btm.t848 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1695 VDAC_N.t235 C7_N_btm.t103 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1696 VDAC_P.t235 C8_P_btm.t209 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1697 VDAC_P.t1683 C9_P_btm.t409 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1698 VDAC_N.t1683 C10_N_btm.t825 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1699 a_83_45776# a_82_45670# VDD.t1627 VDD.t1626 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1700 VDAC_N.t855 C8_N_btm.t210 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1701 VDAC_N.t1681 C7_N_btm.t102 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1702 a_12145_43806# a_12101_44048# a_11979_43806# VSS.t1532 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1703 VDAC_P.t855 C6_P_btm.t51 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1704 a_n1890_42718.t0 a_n1920_42692# VSS.t2199 VSS.t2198 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1705 a_8011_46309# a_7760_45956# a_7552_46134# VDD.t1996 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1706 VDD.t1582 a_9335_44324# a_9266_44350# VDD.t1581 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1707 a_5441_46500# a_5382_44582# VDD.t2027 VDD.t2026 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X1708 VDAC_N.t441 C9_N_btm.t433 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1709 VSS.t3716 C7_P_btm.t7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1710 VDAC_N.t1679 VSS.t3320 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1711 VSS.t221 a_7557_43236.t13 a_8651_45962# VSS.t220 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1712 VDAC_P.t1681 C9_P_btm.t408 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1713 VDAC_N.t853 C10_N_btm.t824 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1714 VDAC_N.t1677 C9_N_btm.t432 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1715 VDAC_P.t441 C10_P_btm.t847 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1716 a_n2293_45420.t3 a_428_42724# VDD.t1054 VDD.t1053 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X1717 VDAC_N.t131 C10_N_btm.t823 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1718 VSS.t3582 C9_P_btm.t19 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1719 VDAC_N.t1675 C10_N_btm.t822 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1720 VDAC_N.t851 C10_N_btm.t821 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1721 VDAC_P.t1679 C10_P_btm.t846 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1722 VDAC_P.t853 C9_P_btm.t407 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1723 VDAC_P.t1677 C10_P_btm.t845 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1724 VDAC_N.t1673 C10_N_btm.t820 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1725 VDAC_N.t439 VSS.t3307 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1726 VDAC_P.t131 C9_P_btm.t406 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1727 VDAC_P.t1675 C9_P_btm.t405 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1728 VDAC_N.t1671 C10_N_btm.t819 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1729 VSS.t3023 VDD.t3109 VSS.t3022 VSS.t3021 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1730 VDAC_P.t851 C9_P_btm.t404 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1731 VDAC_P.t1673 C10_P_btm.t844 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1732 VDAC_N.t849 C9_N_btm.t431 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1733 a_13097_46348# a_6485_44582.t27 VDD.t3026 VDD.t3025 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1734 VDAC_P.t439 C10_P_btm.t843 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1735 VDAC_N.t1669 C8_N_btm.t209 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1736 VDAC_N.t233 C10_N_btm.t818 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1737 VDD.t2603 VSS.t3642 VDD.t2602 VDD.t2601 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1738 VSS.t9 a_10259_42870.t15 a_10215_44874# VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1739 VDAC_N.t1667 C9_N_btm.t430 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1740 VDAC_N.t847 C10_N_btm.t817 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1741 a_19037_42718# a_18759_42746# VDD.t1698 VDD.t1697 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1742 VDAC_P.t1671 C8_P_btm.t208 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1743 a_11529_44670# a_11455_44576.t21 a_11183_44350# VSS.t2716 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1744 VSS.t3087 VDD.t3131 VSS.t3086 VSS.t3085 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1745 a_16211_44582# a_15730_45670.t13 VDD.t491 VDD.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X1746 VDAC_P.t849 C9_P_btm.t403 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1747 VDAC_P.t1669 VSS.t3394 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1748 VDD.t2598 VSS.t3645 VDD.t2597 VDD.t2596 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1749 VSS.t196 a_18394_35068.t12 a_19320_35138# VSS.t195 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1750 VDAC_N.t1665 C8_N_btm.t208 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1751 VDAC_P.t233 C9_P_btm.t402 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1752 VDAC_N.t437 C8_N_btm.t207 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1753 VSS.t2444 VSS.t2445 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1754 VDD.t1836 a_1387_45670# a_656_45670# VDD.t1835 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X1755 VDAC_P.t1667 C4_P_btm.t17 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1756 VDAC_P.t847 C10_P_btm.t842 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1757 a_104_42692# a_283_42692# VDD.t967 VDD.t966 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1758 a_3692_46892# a_3575_46697# VSS.t1575 VSS.t1574 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1759 VDAC_P.t1665 C7_P_btm.t99 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1760 a_n2810_47070.t0 a_n2840_47044# VSS.t2129 VSS.t2128 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1761 C4_P_btm.t22 a_n2442_46526.t4 VREF.t72 VDD.t3078 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1762 C7_P_btm.t1 a_n1890_47614.t4 VREF.t20 VDD.t2038 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1763 VDAC_N.t1663 C9_N_btm.t429 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1764 VDAC_P.t437 C8_P_btm.t207 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1765 VDD.t2592 VSS.t3729 VDD.t2591 VDD.t2590 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1766 VDAC_P.t1663 C9_P_btm.t401 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1767 VDAC_N.t845 C10_N_btm.t816 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1768 VDAC_N.t1661 C9_N_btm.t428 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1769 a_5001_43806# a_4835_43806# VDD.t947 VDD.t946 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1770 a_21788_30659.t0 a_22223_47622# VSS.t1031 VSS.t1030 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1771 VDAC_P.t845 C10_P_btm.t841 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1772 VSS.t3206 VDD.t3171 VSS.t3205 VSS.t3204 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1773 a_16390_43806# a_8727_47222.t9 VSS.t84 VSS.t83 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1774 VSS.t1862 a_18971_44654# a_15730_45670.t2 VSS.t1861 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1775 a_2609_43806# a_2443_43806# VSS.t2100 VSS.t2099 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1776 a_13181_45982# a_13151_45956# a_13097_45982# VSS.t1545 sky130_fd_pr__nfet_01v8 ad=0.085225 pd=0.925 as=0.0567 ps=0.69 w=0.42 l=0.15
X1777 VDAC_P.t1661 C8_P_btm.t206 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1778 VDAC_P.t79 C10_P_btm.t840 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1779 VSS.t2774 a_135_43540.t21 a_4049_43628# VSS.t2773 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1780 VSS.t211 a_4830_43958.t15 a_5939_44894# VSS.t210 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1781 VDAC_N.t79 C9_N_btm.t427 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1782 VDAC_N.t1659 C10_N_btm.t815 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1783 VDAC_P.t1659 C10_P_btm.t839 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1784 VDAC_P.t843 C10_P_btm.t838 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1785 VDAC_P.t1657 C10_P_btm.t837 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1786 VSS.t2131 a_18319_44868# a_12769_44594.t0 VSS.t2130 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X1787 VDAC_P.t435 C10_P_btm.t836 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1788 VDAC_N.t843 C10_N_btm.t814 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1789 VSS.t1542 a_21855_42718# a_13667_32299.t1 VSS.t1541 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1790 VDAC_N.t1657 C10_N_btm.t813 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1791 VDAC_P.t1655 C10_P_btm.t835 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1792 a_21540_43236# a_21719_43244# VDD.t973 VDD.t972 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1793 VSS.t3135 VDD.t3147 VSS.t3134 VSS.t3133 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1794 VSS.t3744 C10_N_btm.t1065 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1795 VDAC_P.t841 C10_P_btm.t834 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1796 VDAC_N.t435 C8_N_btm.t206 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1797 a_n194_47222# a_571_46830# VDD.t1069 VDD.t1068 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1798 a_8204_45412# a_8055_45491# VSS.t2600 VSS.t2599 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1799 VDD.t2579 VSS.t3747 VDD.t2578 VDD.t2517 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1800 a_n2840_43780# a_n2661_43780# VSS.t2157 VSS.t687 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1801 VDAC_P.t1653 C9_P_btm.t400 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1802 a_3787_46904# a_3437_46532# a_3692_46892# VDD.t1829 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1803 a_n243_45982# a_n409_45982# VDD.t978 VDD.t977 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1804 a_18970_45412# a_19566_45670# VDD.t982 VDD.t981 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.17575 ps=1.395 w=0.42 l=0.15
X1805 VSS.t1045 a_16703_45982# a_16757_47070# VSS.t1044 sky130_fd_pr__nfet_01v8 ad=0.2665 pd=2.12 as=0.091 ps=0.93 w=0.65 l=0.15
X1806 a_n1827_45412.t4 a_4908_45956# VDD.t1746 VDD.t1745 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1807 VDAC_N.t1655 C5_N_btm.t14 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1808 VDAC_N.t841 C8_N_btm.t205 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1809 VSS.t613 a_13524_46832.t25 a_13427_46756# VSS.t612 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1810 VDAC_N.t1653 C8_N_btm.t204 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1811 VDAC_N.t231 C10_N_btm.t811 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1812 VDAC_P.t231 C6_P_btm.t50 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1813 VDAC_P.t1651 C7_P_btm.t96 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1814 a_1431_47070# a_n1435_47614.t2 VSS.t2997 VSS.t2996 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1815 VDD.t2004 a_2351_47614# DATA[2].t6 VDD.t2003 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1816 a_17242_43806# a_12769_44594.t6 a_17073_44056# VDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X1817 VREF.t2 a_n2810_47070.t6 C8_P_btm.t2 VDD.t88 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1818 VSS.t1047 a_9637_43560# a_9571_43628# VSS.t1046 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1819 a_n2472_44324# a_n2293_44332# VSS.t2132 VSS.t1491 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1820 VSS.t3656 C9_P_btm.t23 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1821 VDAC_N.t1651 C10_N_btm.t810 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1822 VDD.t912 a_8483_43780# a_6485_44582.t6 VDD.t911 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X1823 VDAC_P.t839 C9_P_btm.t396 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1824 VDAC_P.t1649 C8_P_btm.t205 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1825 VDD.t2937 CAL_P.t3 VDD.t2937 VDD.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X1826 VDAC_N.t839 C9_N_btm.t426 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1827 VDD.t1560 a_1123_43780# a_1581_43806.t5 VDD.t1559 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X1828 VSS.t3435 VDD.t3203 VSS.t3434 VSS.t3433 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1829 VDAC_N.t1649 C9_N_btm.t425 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1830 VDAC_N.t433 C9_N_btm.t424 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1831 VDAC_P.t433 C10_P_btm.t412 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1832 a_16273_46232# a_10251_45454# a_16085_45982# VDD.t1299 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2125 ps=1.425 w=1 l=0.15
X1833 a_9060_45144# a_1412_46794.t7 VDD.t165 VDD.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X1834 VDAC_P.t1647 C10_P_btm.t833 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1835 VSS.t1561 a_16211_43780# a_16145_43806# VSS.t1560 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1836 a_6954_46348# a_6196_46250# a_6391_46219# VDD.t993 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1837 VSS.t2303 VSS.t2304 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1838 VDAC_N.t1647 C10_N_btm.t809 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1839 VDAC_P.t837 C10_P_btm.t832 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1840 VDAC_N.t837 C10_N_btm.t808 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1841 VDAC_P.t1645 C10_P_btm.t831 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1842 VSS.t3123 VDD.t3143 VSS.t3122 VSS.t3121 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1843 VDAC_P.t129 C10_P_btm.t830 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1844 VDAC_N.t1645 C10_N_btm.t807 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1845 VDAC_Pi.t3 a_3754_38470.t5 a_4338_37500.t4 VSS.t2839 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1846 VDAC_N.t129 C9_N_btm.t423 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1847 VDAC_P.t1643 C10_P_btm.t829 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1848 VDAC_P.t835 C9_P_btm.t395 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1849 VDAC_P.t1641 C9_P_btm.t394 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1850 VDAC_N.t1643 C8_N_btm.t203 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1851 VDD.t995 a_9863_47874# DEBUG_OUT.t7 VDD.t994 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1852 VDAC_N.t835 C10_N_btm.t806 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1853 CLK_DATA.t3 a_n2833_47874# VSS.t1385 VSS.t1384 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X1854 VDAC_P.t431 C10_P_btm.t828 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1855 VDAC_N.t1641 C8_N_btm.t202 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1856 VSS.t3401 VDD.t3191 VSS.t3400 VSS.t3399 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1857 a_16750_46134# a_15187_44868# a_17053_46232# VDD.t1207 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X1858 VDD.t2558 VSS.t3569 VDD.t2557 VDD.t2556 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1859 a_2252_42718.t3 a_2075_42718# VDD.t1257 VDD.t1256 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1860 VSS.t2004 a_n1085_47874# DATA[0].t2 VSS.t2003 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1861 VDD.t257 a_3990_30651.t13 a_19555_42718# VDD.t256 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1862 VDAC_N.t431 C10_N_btm.t805 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1863 VDD.t2935 a_n2103_44868.t12 a_22223_47622# VDD.t276 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1864 a_15328_46134# a_13524_46832.t11 VSS.t603 VSS.t602 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1865 VSS.t2507 VSS.t2508 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1866 VDAC_P.t1639 C10_P_btm.t827 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1867 VSS.t2572 a_10844_44364# a_10596_44324# VSS.t2571 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1868 a_6519_43494# a_6485_44582.t15 a_6665_43582# VSS.t2913 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X1869 VDAC_N.t1639 C10_N_btm.t804 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1870 a_5626_46846# a_5419_47258# VSS.t1591 VSS.t1590 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.203125 ps=1.275 w=0.65 l=0.15
X1871 VDAC_N.t833 C3_N_btm.t6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1872 VDAC_N.t1637 C8_N_btm.t201 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1873 VDAC_P.t833 C8_P_btm.t204 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1874 VSS.t2355 VSS.t2356 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1875 VDD.t2172 a_4527_43566# a_4514_43262# VDD.t2171 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1876 VDAC_N.t229 C8_N_btm.t200 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1877 VDAC_N.t1635 C8_N_btm.t199 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1878 VDAC_N.t831 C10_N_btm.t803 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1879 VSS.t2436 VSS.t2437 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1880 VDD.t1980 a_1387_44582# a_n172_44582# VDD.t1979 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X1881 VDAC_P.t1637 C7_P_btm.t95 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1882 VDD.t2549 VSS.t3622 VDD.t2548 VDD.t2547 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1883 VSS.t974 a_5784_44364# a_6126_46642# VSS.t973 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1884 VDAC_P.t229 C8_P_btm.t203 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1885 a_6985_45438# a_6707_45776# VDD.t1521 VDD.t1520 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1886 VDAC_N.t1633 C10_N_btm.t802 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1887 VDAC_P.t1635 C9_P_btm.t393 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1888 VDAC_N.t429 C9_N_btm.t422 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1889 VDAC_N.t1631 C10_N_btm.t801 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1890 VDAC_P.t831 VSS.t3352 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1891 VSS.t1874 a_13991_42883# a_12684_45276# VSS.t1873 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1892 VSS.t2655 a_11795_47044# a_10227_47214.t3 VSS.t2654 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1893 VDAC_N.t829 C10_N_btm.t800 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1894 VDAC_N.t1629 C8_N_btm.t198 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1895 a_1203_42692.t1 a_1431_47070# VSS.t2218 VSS.t2217 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.26 ps=1.45 w=0.65 l=0.15
X1896 VDAC_P.t1633 C10_P_btm.t826 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1897 VDAC_P.t429 C9_P_btm.t392 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1898 VDAC_N.t53 C10_N_btm.t799 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1899 VDAC_N.t1627 C10_N_btm.t394 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1900 a_2609_43806# a_2443_43806# VDD.t2060 VDD.t2059 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1901 VDAC_N.t827 C10_N_btm.t798 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1902 VDD.t2918 RST_Z.t1 a_8530_39574# VDD.t2917 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1903 VDAC_P.t1631 C10_P_btm.t825 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1904 VDAC_P.t829 C10_P_btm.t824 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1905 VDAC_P.t1629 C10_P_btm.t823 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1906 VDAC_P.t53 C10_P_btm.t822 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1907 VDAC_N.t1625 C9_N_btm.t421 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1908 VDAC_P.t1627 C7_P_btm.t94 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1909 VDAC_N.t427 C10_N_btm.t797 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1910 VDD.t2540 VSS.t3600 VDD.t2539 VDD.t2538 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1911 VDAC_P.t827 C10_P_btm.t821 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1912 VDAC_P.t1625 C4_P_btm.t18 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1913 a_9179_44592# a_9521_45982.t9 VSS.t27 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1914 a_11059_45956# a_10227_47214.t33 VDD.t132 VDD.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1915 VDAC_P.t427 C9_P_btm.t391 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1916 VDAC_P.t1623 C10_P_btm.t820 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1917 a_4352_46904# a_3271_46532# a_4005_46500# VDD.t1620 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1918 VDAC_N.t1623 C7_N_btm.t101 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1919 a_4703_44894# a_2587_44868.t15 VSS.t240 VSS.t239 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1920 VDAC_N.t825 C9_N_btm.t420 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1921 VSS.t1155 a_3328_44324# a_n2293_45956.t1 VSS.t1154 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X1922 VDAC_N.t1621 C5_N_btm.t2 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1923 VDAC_P.t825 C10_P_btm.t819 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1924 VSS.t3698 C2_N_btm.t6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1925 VDAC_N.t227 C10_N_btm.t796 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1926 VSS.t2297 VSS.t2298 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1927 C10_P_btm.t1063 a_n4515_30659.t11 VREF.t60 VDD.t2997 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1928 VDAC_N.t1619 C9_N_btm.t419 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1929 VDAC_N.t823 C10_N_btm.t795 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1930 VDAC_N.t1617 C8_N_btm.t197 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1931 VDAC_P.t1621 C10_P_btm.t818 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1932 VSS.t1082 a_21997_47833# a_1651_47044.t0 VSS.t1081 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1933 VDAC_P.t227 C8_P_btm.t202 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1934 VDAC_N.t425 C9_N_btm.t418 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1935 VDD.t2170 a_4527_43566# a_927_42692.t6 VDD.t2169 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X1936 VDAC_N.t1615 VSS.t3324 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1937 VSS.t1084 a_22591_45982# a_19921_31459.t1 VSS.t1083 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1938 VDAC_P.t1619 C9_P_btm.t390 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1939 VDAC_N.t821 C10_N_btm.t794 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1940 a_13023_44716# a_10259_42870.t13 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1941 VDD.t2751 a_11795_47044# a_10227_47214.t6 VDD.t2750 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X1942 VSS.t3580 C10_N_btm.t1066 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1943 VDAC_P.t823 C10_P_btm.t817 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1944 VSS.t956 a_5839_47070# a_5847_47614# VSS.t955 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X1945 VDAC_N.t1613 C10_N_btm.t792 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1946 VDAC_P.t1617 C9_P_btm.t389 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1947 a_6701_45982# a_6322_46348# a_6629_45982# VSS.t1089 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1948 VSS.t2341 VSS.t2342 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1949 VDAC_P.t425 VSS.t3369 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1950 a_19520_46500# a_19371_46579# a_19816_46642# VDD.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1951 VDAC_N.t127 C9_N_btm.t417 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1952 VDAC_P.t1615 C10_P_btm.t816 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1953 VDAC_N.t1611 VSS.t3323 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1954 VDAC_N.t819 C9_N_btm.t416 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1955 VSS.t2959 a_14409_32299.t4 C5_N_btm.t37 VSS.t456 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1956 VDD.t2528 VSS.t3705 VDD.t2527 VDD.t2526 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1957 VDAC_P.t821 C10_P_btm.t815 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1958 VDAC_N.t1609 C8_N_btm.t196 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1959 a_2709_43582# a_927_42692.t18 VSS.t96 VSS.t95 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1960 VDD.t2525 VSS.t3708 VDD.t2524 VDD.t2523 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1961 VSS.t2287 VSS.t2288 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1962 VDAC_P.t1613 C6_P_btm.t49 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1963 VSS.t2558 a_n2661_46508.t8 a_21755_44350# VSS.t2557 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1964 VDD.t1452 a_n2472_45956# a_n2442_45982.t2 VDD.t1451 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1965 VDAC_P.t127 C7_P_btm.t93 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1966 COMP_P.t7 a_1239_39587# VDD.t1714 VDD.t1713 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1967 VDAC_P.t1611 C6_P_btm.t48 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1968 a_4000_42718.t0 a_3823_42718# VSS.t1698 VSS.t1697 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1969 a_18444_47070# a_15549_47044.t8 VSS.t2894 VSS.t2893 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1970 C6_N_btm.t0 EN_VIN_BSTR_N.t13 VIN_N.t3 VSS.t442 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1971 a_18766_43236# a_21197_42718# VSS.t1095 VSS.t1094 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1972 a_20159_47588# DEBUG_MUX[1].t0 VDD.t156 VDD.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X1973 VDAC_P.t819 C9_P_btm.t388 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1974 VSS.t2553 VSS.t2554 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1975 VDAC_P.t1609 C10_P_btm.t814 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1976 a_3165_43262# a_2627_43262# VDD.t1038 VDD.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1977 VDAC_N.t423 C9_N_btm.t415 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1978 VDD.t120 a_15163_45670.t7 a_14953_45554# VDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X1979 a_768_44670# a_927_42692.t20 VSS.t98 VSS.t97 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1980 VDAC_N.t1607 C6_N_btm.t59 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1981 VDD.t2869 a_n2293_45420.t8 a_21719_43244# VDD.t2868 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1982 VDD.t3009 a_1581_43806.t13 a_19274_43262# VDD.t3008 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X1983 a_n2442_45438.t1 a_n2472_45412# VSS.t1451 VSS.t1450 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1984 VDAC_P.t423 C8_P_btm.t201 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1985 a_14409_32299.t2 a_22591_43806# VDD.t1944 VDD.t1943 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1986 VDAC_N.t817 C10_N_btm.t791 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1987 VDAC_N.t1605 C10_N_btm.t790 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1988 VDAC_N.t225 C9_N_btm.t414 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1989 VDAC_P.t1607 C8_P_btm.t200 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1990 VSS.t2675 a_n1920_47588# a_n1890_47614.t1 VSS.t2674 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1991 VSS.t1801 a_4527_46830# a_4322_46134# VSS.t1800 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1992 VDAC_N.t1603 C9_N_btm.t413 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1993 a_4338_37500.t3 a_3754_38470.t6 VDAC_Pi.t2 VSS.t2840 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1994 a_10500_46892# a_10383_46697# VDD.t1040 VDD.t1039 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1995 VDAC_P.t817 C10_P_btm.t813 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1996 VDAC_P.t1605 C8_P_btm.t199 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X1997 a_10592_43628# a_10475_43433# VDD.t1042 VDD.t1041 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1998 VDD.t235 a_2587_44868.t13 a_4733_44350# VDD.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1999 VDAC_P.t225 C8_P_btm.t198 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2000 VDAC_N.t815 C9_N_btm.t412 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2001 VDAC_N.t1601 C10_N_btm.t789 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2002 VDAC_N.t421 C10_N_btm.t788 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2003 a_13915_44670# a_13561_44350# a_13725_44350# VSS.t1106 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2004 VDAC_N.t1599 C10_N_btm.t388 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2005 a_12896_47044# a_12747_47070# VSS.t789 VSS.t788 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2006 VDAC_P.t1603 C10_P_btm.t812 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2007 a_49_43236# a_n169_43640# VSS.t791 VSS.t790 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2008 VSS.t1582 a_4091_47070# a_4651_47614# VSS.t1581 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X2009 VDAC_P.t815 C8_P_btm.t197 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2010 EN_VIN_BSTR_N.t3 a_18394_35068.t13 w_11534_34010.t5 w_11534_34010.t4 sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2011 VDD.t305 a_10227_47214.t31 a_19771_43600# VDD.t304 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2012 VDAC_P.t1601 C10_P_btm.t811 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2013 VDAC_N.t813 C7_N_btm.t100 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2014 VDAC_P.t421 C10_P_btm.t810 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2015 VDAC_N.t1597 C9_N_btm.t411 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2016 a_5700_37509.t16 VSS.t3641 VDAC_Pi.t4 VDD.t2494 sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2017 a_9667_43301# a_9416_43530# a_9208_43494# VDD.t1437 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X2018 VDAC_N.t77 C7_N_btm.t99 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2019 VDAC_P.t1599 C6_P_btm.t47 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2020 VDD.t936 a_8379_46134# a_7648_46134# VDD.t935 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X2021 a_22717_37323# a_22459_39581# a_22609_38426# VSS.t2165 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2022 VDAC_N.t1595 C9_N_btm.t410 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2023 VDAC_P.t813 C7_P_btm.t92 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2024 a_18103_46768# a_14950_43958# VSS.t1437 VSS.t1436 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2025 VDAC_P.t1597 C8_P_btm.t196 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2026 VSS.t3643 C10_P_btm.t22 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2027 a_18135_47588# DEBUG_MUX[0].t0 VSS.t143 VSS.t142 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X2028 VDD.t231 a_2587_44868.t11 a_10069_42968# VDD.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2029 a_4005_43236# a_3787_43640# VSS.t793 VSS.t792 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2030 a_11883_43806# a_11367_43806# a_11788_43806# VSS.t1673 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2031 a_4908_45956# a_11335_46830# VSS.t923 VSS.t922 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2032 VDAC_P.t77 C10_P_btm.t809 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2033 VDD.t2970 a_12651_44576.t21 a_n2103_44868.t4 VDD.t2969 sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.135 ps=1.27 w=1 l=0.15
X2034 VDAC_P.t1595 C9_P_btm.t387 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2035 VDAC_N.t811 C4_N_btm.t7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2036 VDAC_P.t811 C9_P_btm.t386 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2037 VSS.t338 a_10227_47214.t17 a_10857_46892# VSS.t337 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2038 VDAC_P.t1593 C10_P_btm.t808 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2039 VDAC_N.t1593 C9_N_btm.t409 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2040 VDAC_N.t419 C9_N_btm.t408 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2041 VSS.t3644 C7_N_btm.t135 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2042 VDAC_P.t419 C9_P_btm.t385 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2043 VDAC_N.t1591 C10_N_btm.t787 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2044 VDAC_N.t809 C10_N_btm.t786 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2045 a_743_47397# a_85_47070# a_284_47222# VDD.t2031 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X2046 a_15489_43268# a_15323_43268# VDD.t1369 VDD.t1368 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2047 VDAC_N.t1589 C9_N_btm.t407 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2048 a_n1067_42718.t1 a_n1237_42718# VDD.t2743 VDD.t2742 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2049 VDAC_P.t1591 C10_P_btm.t807 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2050 VSS.t3250 VDD.t3187 VSS.t3249 VSS.t3248 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2051 VDAC_P.t809 C9_P_btm.t384 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2052 VDAC_N.t223 C9_N_btm.t406 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2053 VDAC_P.t1589 C9_P_btm.t383 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2054 VDAC_N.t1587 C10_N_btm.t785 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2055 VDAC_P.t223 C10_P_btm.t806 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2056 VDAC_N.t807 C10_N_btm.t784 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2057 VDAC_P.t1587 C10_P_btm.t805 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2058 VDAC_P.t807 C9_P_btm.t382 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2059 C8_P_btm.t7 EN_VIN_BSTR_P.t15 VIN_P.t11 VSS.t557 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2060 VDAC_P.t1585 C9_P_btm.t381 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2061 VDAC_P.t417 C10_P_btm.t804 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2062 VSS.t3606 C9_N_btm.t527 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2063 VDAC_P.t1583 C9_P_btm.t380 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2064 VDAC_P.t805 C10_P_btm.t803 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2065 a_7459_47397# a_7208_47044# a_7000_47222# VDD.t2706 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X2066 VDD.t3007 a_1581_43806.t11 a_13827_46298# VDD.t3006 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.090125 ps=0.995 w=0.42 l=0.15
X2067 VDAC_N.t1585 C10_N_btm.t783 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2068 a_18357_44048# a_18139_43806# VSS.t1940 VSS.t1939 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2069 a_22521_41035# COMP_P.t8 VDD.t65 VDD.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2070 VDD.t1976 a_18970_45412# a_n2103_45412.t0 VDD.t1975 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2071 VDD.t730 a_16291_46758# a_16128_46134# VDD.t729 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X2072 VDAC_N.t417 C9_N_btm.t404 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2073 VDAC_N.t1583 C6_N_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2074 VDAC_P.t1581 C10_P_btm.t802 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2075 VDAC_N.t805 C6_N_btm.t57 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2076 a_18235_43806# a_17789_43806# a_18139_43806# VSS.t1131 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2077 VDAC_N.t1581 C8_N_btm.t195 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2078 VDAC_Pi.t6 VSS.t3728 a_5700_37509.t18 VDD.t2490 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2079 DATA[3].t5 a_4651_47614# VDD.t1347 VDD.t1346 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2080 VSS.t2279 VSS.t2280 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2081 VDAC_N.t125 C10_N_btm.t782 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2082 VDAC_N.t1579 C6_N_btm.t2 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2083 a_15049_44466# a_10114_45276.t9 a_14954_44466# VDD.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X2084 VDAC_P.t125 C7_P_btm.t91 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2085 VDAC_N.t803 C9_N_btm.t403 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2086 a_4993_47044# a_4322_46134# VDD.t1772 VDD.t1771 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2087 a_10592_43628# a_10475_43433# VSS.t1105 VSS.t1104 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2088 VDAC_P.t1579 C8_P_btm.t195 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2089 VDD.t2023 a_5382_44582# a_5387_44403# VDD.t2022 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2090 a_6104_45706.t1 a_16211_43780# VDD.t1500 VDD.t1499 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2091 VDAC_N.t1577 C10_N_btm.t781 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2092 VDAC_P.t803 C10_P_btm.t801 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2093 VSS.t1232 a_7595_47614# DATA[5].t0 VSS.t1231 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2094 VSS.t213 a_4830_43958.t16 a_4835_43806# VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2095 VDAC_N.t415 C8_N_btm.t194 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2096 VDAC_N.t1575 C10_N_btm.t780 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2097 a_n2442_44350.t1 a_n2472_44324# VSS.t1049 VSS.t741 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2098 VDAC_N.t801 C10_N_btm.t779 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2099 VDAC_N.t1573 C9_N_btm.t402 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2100 VDAC_N.t221 C10_N_btm.t778 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2101 a_7347_43494# a_7557_43236.t14 a_7493_43582# VSS.t222 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X2102 a_n2472_43780# a_n2293_43780# VSS.t1206 VSS.t1205 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2103 VDAC_N.t1571 C8_N_btm.t193 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2104 VDAC_N.t799 C10_N_btm.t777 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2105 VDAC_P.t1577 C9_P_btm.t379 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2106 VDAC_N.t1569 C10_N_btm.t776 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2107 a_22609_38842# a_22521_39947# CAL_N.t0 VDD.t2685 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2108 a_7497_44466# a_7309_44466# a_7415_44466# VDD.t737 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2109 VDAC_P.t415 C10_P_btm.t800 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2110 VDAC_P.t1575 C10_P_btm.t799 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2111 VSS.t2874 a_1581_43806.t9 a_2905_44894# VSS.t2873 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2112 VDAC_P.t801 C9_P_btm.t378 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2113 C10_N_btm.t23 a_22812_30659.t9 VREF.t32 VDD.t521 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2114 VDAC_N.t413 C9_N_btm.t401 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2115 VCM.t58 a_4758_30651.t7 C9_N_btm.t537 VSS.t2988 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2116 VDD.t997 a_9863_47874# DEBUG_OUT.t6 VDD.t996 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X2117 a_4343_45816# a_3897_45444# a_4247_45816# VSS.t2158 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2118 VSS.t2213 a_9343_43806# a_5655_43780# VSS.t2212 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2119 a_11730_34132.t3 EN_VIN_BSTR_N.t9 VIN_N.t15 VSS.t438 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2120 VSS.t2106 a_n2840_45412# a_n2810_45438.t1 VSS.t1654 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2121 a_3733_46348# a_3470_45982# a_3320_46134# VDD.t1532 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2122 VSS.t2730 a_1847_45528.t15 a_4080_44670# VSS.t2729 sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.08775 ps=0.92 w=0.65 l=0.15
X2123 VSS.t1147 a_1115_47044# a_n53_44363.t0 VSS.t1146 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X2124 VCM.t21 a_4000_42718.t7 C2_N_btm.t0 VSS.t298 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2125 a_4704_47044# a_4993_47044# a_4927_47070# VSS.t1423 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2126 VDAC_P.t1573 C10_P_btm.t798 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2127 a_8912_37509.t29 VDAC_P.t221 a_5088_37509.t11 VDD.t2253 sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X2128 a_4842_45982# a_885_44868.t27 VSS.t2758 VSS.t2757 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2129 VDAC_N.t1567 C5_N_btm.t25 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2130 a_4465_45412# a_4247_45816# VDD.t1915 VDD.t1914 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2131 VDAC_P.t1571 C8_P_btm.t194 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2132 a_18813_45982# a_17623_45982# a_18704_45982# VSS.t1143 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2133 VDAC_N.t797 C6_N_btm.t55 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2134 VDAC_N.t1565 C8_N_btm.t192 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2135 a_6391_46219# a_6196_46250# a_6701_45982# VSS.t1052 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X2136 VDAC_N.t31 C10_N_btm.t771 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2137 VDAC_P.t799 C6_P_btm.t46 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2138 VDAC_P.t1569 C10_P_btm.t797 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2139 VDAC_P.t413 C8_P_btm.t193 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2140 VDAC_N.t1563 C9_N_btm.t399 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2141 a_10259_42870.t5 a_12623_43780# VDD.t1241 VDD.t1240 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2142 VSS.t3765 C9_P_btm.t15 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2143 VDAC_P.t1567 C7_P_btm.t90 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2144 a_135_43540.t2 a_8391_47044# VSS.t1208 VSS.t1207 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2145 VDAC_P.t797 C9_P_btm.t376 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2146 VSS.t3770 C9_N_btm.t529 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2147 VDAC_N.t795 C10_N_btm.t770 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2148 VDD.t1458 a_22223_44358# a_14601_32299.t2 VDD.t1457 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2149 VDAC_N.t1561 C10_N_btm.t769 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2150 VDAC_N.t411 C9_N_btm.t397 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2151 a_13373_46526# a_13524_46832.t22 a_13457_46892# VDD.t554 sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2152 VSS.t3153 VDD.t3153 VSS.t3152 VSS.t3151 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2153 VDAC_P.t1565 C10_P_btm.t796 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2154 VDAC_P.t31 C10_P_btm.t795 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2155 VDAC_N.t1559 C10_N_btm.t768 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2156 VDAC_N.t793 C10_N_btm.t767 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2157 VSS.t1057 a_9863_47874# DEBUG_OUT.t1 VSS.t1056 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2158 a_2343_47070# a_2167_46526# VDD.t2101 VDD.t2100 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2159 VDAC_N.t1557 C10_N_btm.t766 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2160 VDAC_N.t219 C10_N_btm.t765 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2161 a_14853_45438# a_14766_45596.t7 VSS.t2802 VSS.t2801 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2162 C4_P_btm.t1 a_5923_31099.t7 VCM.t27 VSS.t146 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2163 VDAC_N.t1555 C9_N_btm.t396 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2164 VDAC_P.t1563 C9_P_btm.t375 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2165 a_12438_45412# a_12684_45276# VSS.t1073 VSS.t1072 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.11975 ps=1.045 w=0.42 l=0.15
X2166 VSS.t2409 VSS.t2410 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2167 a_636_42870# a_571_43566# VSS.t817 VSS.t816 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2168 VDAC_P.t795 C10_P_btm.t794 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2169 a_10337_43268# a_10171_43268# VDD.t2146 VDD.t2145 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2170 a_2301_45758# a_1847_45528.t13 VSS.t2728 VSS.t2727 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X2171 VDAC_P.t1561 C10_P_btm.t793 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2172 VREF.t15 a_n2467_30659.t8 C9_P_btm.t9 VDD.t581 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2173 VDAC_N.t791 C9_N_btm.t395 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2174 VDD.t1810 a_18689_45412# a_18993_47320# VDD.t1809 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2175 VDAC_P.t411 C7_P_btm.t89 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2176 VDAC_N.t1553 C2_N_btm.t4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2177 VDAC_N.t409 C10_N_btm.t764 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2178 a_n264_43628# a_n381_43433# VDD.t1848 VDD.t1847 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2179 VDAC_P.t1559 C9_P_btm.t374 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2180 VDAC_N.t1551 C10_N_btm.t763 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2181 VDAC_N.t789 C10_N_btm.t762 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2182 VSS.t2407 VSS.t2408 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2183 VDAC_N.t1549 C8_N_btm.t191 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2184 VDAC_P.t793 C10_P_btm.t792 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2185 a_10425_47070# a_9947_47044# VSS.t2020 VSS.t2019 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2186 VDAC_P.t1557 C7_P_btm.t88 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2187 VDD.t1419 a_15689_44048# a_15579_44172# VDD.t1418 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2188 VDAC_P.t219 C10_P_btm.t791 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2189 a_3437_43268# a_3271_43268# VSS.t2109 VSS.t2108 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2190 VDAC_N.t123 C9_N_btm.t394 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2191 VDD.t1858 a_22959_45982# a_20405_31459.t3 VDD.t1857 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2192 VIN_P.t10 EN_VIN_BSTR_P.t13 C8_P_btm.t6 VSS.t555 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2193 a_361_45438# a_83_45776# VSS.t1976 VSS.t1975 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X2194 VDAC_P.t1555 C9_P_btm.t373 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2195 VDAC_N.t1547 C8_N_btm.t93 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2196 VSS.t2038 a_16824_45276# a_16576_44868# VSS.t2037 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2197 VDAC_P.t791 C9_P_btm.t372 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2198 VSS.t3519 VDD.t3233 VSS.t3518 VSS.t3517 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2199 VDD.t2103 a_14545_44569# a_10114_45276.t1 VDD.t2102 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2200 VDAC_P.t1553 C10_P_btm.t790 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2201 VDAC_N.t787 C10_N_btm.t761 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2202 VDD.t202 a_4830_43958.t10 a_4835_43806# VDD.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2203 VDAC_N.t1545 C10_N_btm.t760 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2204 VDAC_P.t409 C10_P_btm.t789 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2205 VDAC_P.t1551 C10_P_btm.t788 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2206 VDAC_P.t789 C10_P_btm.t787 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2207 VIN_P.t5 EN_VIN_BSTR_P.t11 C6_P_btm.t0 VSS.t553 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2208 VSS.t540 a_1203_42692.t25 a_10901_42718# VSS.t539 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2209 VSS.t3789 C10_N_btm.t1067 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2210 a_15730_45670.t3 a_18971_44654# VSS.t1866 VSS.t1865 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2211 a_19150_44716# a_10227_47214.t15 VSS.t334 VSS.t333 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2212 a_13097_45982# a_6485_44582.t13 VSS.t2910 VSS.t2909 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2213 a_5377_47320# a_1429_47222.t11 a_n2497_47846.t1 VDD.t323 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2214 VDAC_N.t407 C10_N_btm.t758 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2215 VDAC_P.t1549 C10_P_btm.t786 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2216 VDAC_N.t1543 C9_N_btm.t393 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2217 a_18044_45982# a_17927_46195# VSS.t1946 VSS.t1945 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2218 VDAC_P.t123 C8_P_btm.t189 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2219 VDAC_P.t1547 C9_P_btm.t371 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2220 VCM.t52 a_5542_30651.t6 C6_N_btm.t73 VSS.t2835 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2221 a_191_44389# a_n60_44618# a_n268_44582# VDD.t764 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X2222 VSS.t495 a_n237_45454.t12 a_6793_45776# VSS.t494 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2223 VDAC_P.t787 C10_P_btm.t785 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2224 VDAC_P.t1545 C10_P_btm.t784 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2225 a_15221_47044# a_15163_45670.t9 VSS.t119 VSS.t118 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.10075 ps=0.96 w=0.65 l=0.15
X2226 a_n1732_35090.t3 SMPL.t15 VSS.t2946 VSS.t2945 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2227 a_n2104_43236# a_n2073_43806# VDD.t766 VDD.t765 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2228 a_16561_45982# a_16085_45982# VSS.t1051 VSS.t1050 sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.12675 ps=1.04 w=0.65 l=0.15
X2229 VSS.t938 a_n2840_44324# a_n2810_44350.t1 VSS.t937 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2230 VDAC_N.t785 C10_N_btm.t374 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2231 VDAC_P.t407 C9_P_btm.t370 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2232 VDAC_P.t1543 C10_P_btm.t783 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2233 VSS.t2270 a_9343_42718# a_5734_30651.t0 VSS.t2269 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2234 VDAC_P.t785 C10_P_btm.t782 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2235 a_13469_44894# a_12931_44894# VDD.t2729 VDD.t2728 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X2236 VDAC_P.t1541 C9_P_btm.t369 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2237 VSS.t3105 VDD.t3137 VSS.t3104 VSS.t3103 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2238 VDAC_N.t1541 C5_N_btm.t24 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2239 a_13273_44868.t6 a_18879_43780# VDD.t1568 VDD.t1567 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2240 VDAC_P.t217 C9_P_btm.t368 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2241 VDAC_N.t217 C10_N_btm.t756 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2242 VDD.t904 a_8483_43780# a_8470_44172# VDD.t903 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2243 VDAC_N.t1539 C10_N_btm.t755 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2244 VDAC_N.t783 C8_N_btm.t188 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2245 VSS.t336 a_10227_47214.t16 a_10185_47070# VSS.t335 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X2246 VDAC_N.t1537 C9_N_btm.t392 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2247 VDAC_N.t405 C10_N_btm.t754 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2248 VDAC_P.t1539 C10_P_btm.t781 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2249 a_3328_44324# a_3165_45982# VSS.t1463 VSS.t1462 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X2250 VDAC_N.t1535 C9_N_btm.t391 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2251 VDAC_P.t783 C10_P_btm.t780 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2252 VDD.t1223 a_8659_44324# a_1053_45123.t1 VDD.t1222 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X2253 VDAC_N.t781 C10_N_btm.t753 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2254 VSS.t3803 C8_P_btm.t10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2255 a_5088_37509.t10 VDAC_P.t1537 a_8912_37509.t28 VDD.t2252 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2256 VSS.t839 a_14133_43780# a_14077_44133# VSS.t838 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X2257 VDAC_P.t405 C10_P_btm.t779 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2258 a_6485_44582.t5 a_8483_43780# VDD.t910 VDD.t909 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2259 a_18231_44728# a_17881_44356# a_18136_44716# VDD.t2780 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2260 a_7195_44868# a_5655_43780# VDD.t2213 VDD.t2212 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2261 VDAC_P.t1535 C8_P_btm.t187 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2262 VDAC_P.t781 C10_P_btm.t778 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2263 VSS.t3407 VDD.t3193 VSS.t3406 VSS.t3405 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2264 a_1581_43806.t6 a_1123_43780# VDD.t1558 VDD.t1557 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2265 VDAC_P.t1533 C9_P_btm.t367 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2266 VDAC_N.t1533 C9_N_btm.t390 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2267 VDAC_P.t75 C10_P_btm.t777 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2268 VDAC_N.t75 C10_N_btm.t752 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2269 VDAC_N.t1531 C10_N_btm.t751 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2270 VDAC_N.t779 C10_N_btm.t750 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2271 VDAC_P.t1531 C10_P_btm.t776 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2272 VDAC_P.t779 C10_P_btm.t775 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2273 VDAC_N.t1529 C10_N_btm.t749 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2274 CLK_DATA.t2 a_n2833_47874# VSS.t1387 VSS.t1386 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2275 a_1346_46565# a_885_44868.t33 VDD.t2852 VDD.t2851 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2276 a_10427_46348# a_9803_45982# a_10319_45982# VDD.t2669 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2277 VDD.t2645 VSS.t3596 VDD.t2644 VDD.t2643 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2278 VDAC_N.t403 C10_N_btm.t748 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2279 VSS.t29 a_9521_45982.t10 a_9803_45982# VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2280 VDAC_N.t1527 VSS.t3328 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2281 a_11645_45554# a_10114_45276.t2 a_11550_45554# VDD.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X2282 VDAC_P.t1529 C10_P_btm.t774 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2283 VDAC_P.t403 C10_P_btm.t773 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2284 VDD.t1570 a_18879_43780# a_13273_44868.t4 VDD.t1569 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2285 VDAC_P.t1527 C5_P_btm.t5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2286 VDAC_N.t777 C10_N_btm.t747 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2287 a_18803_47070# a_18530_47070# VDD.t1897 VDD.t1896 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2288 a_13460_43640# a_12379_43268# a_13113_43236# VDD.t1098 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2289 a_n1551_44324.t3 a_10414_43780# a_10362_43806# VSS.t2575 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2290 a_18495_44868# a_16291_44914# VDD.t1670 VDD.t1669 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X2291 a_14573_47070# a_14219_47070# VDD.t784 VDD.t783 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2292 VSS.t2289 VSS.t2290 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2293 VDAC_N.t1525 C7_N_btm.t97 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2294 a_10596_44324# a_1053_45123.t9 VSS.t584 VSS.t583 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X2295 VDAC_P.t777 C10_P_btm.t772 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2296 VDAC_N.t215 VSS.t3297 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2297 C10_P_btm.t9 EN_VIN_BSTR_P.t9 VIN_P.t8 VSS.t551 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X2298 a_12436_44868# a_12287_44894# VSS.t846 VSS.t845 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2299 VDAC_N.t1523 C7_N_btm.t96 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2300 VDAC_N.t775 C10_N_btm.t746 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2301 VDD.t1899 a_10813_46500# a_10703_46526# VDD.t1898 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2302 VDD.t2393 VSS.t3814 VDD.t2392 VDD.t2391 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2303 VDAC_N.t1521 C10_N_btm.t745 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2304 a_n2293_43780# a_n1827_44868.t11 VDD.t281 VDD.t280 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2305 VDAC_N.t401 C8_N_btm.t187 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2306 VSS.t2476 VSS.t2477 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2307 VDAC_P.t1525 C10_P_btm.t767 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2308 a_8848_44868# a_8699_44894# a_9144_45144# VDD.t786 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2309 VDAC_N.t1519 C9_N_btm.t389 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2310 VDD.t2105 a_10905_43236# a_10795_43262# VDD.t2104 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2311 VDD.t749 a_12438_45412# a_n1551_45412.t2 VDD.t748 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2312 VDAC_P.t215 C10_P_btm.t766 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2313 a_22812_30659.t0 a_22959_47622# VSS.t1759 VSS.t1758 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2314 VDAC_P.t1523 C8_P_btm.t186 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2315 VDAC_N.t773 C10_N_btm.t744 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2316 VDD.t2384 VSS.t3719 VDD.t2383 VDD.t2382 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2317 VDAC_N.t1517 VSS.t3327 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2318 VDAC_P.t775 VSS.t3359 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2319 VDAC_P.t1521 C10_P_btm.t765 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2320 VDAC_N.t121 C9_N_btm.t388 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2321 VSS.t2430 VSS.t2431 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2322 a_10362_43806# a_1053_45123.t4 a_10612_43806# VSS.t580 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2323 a_10884_45982# a_9803_45982# a_10537_46224# VDD.t2672 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2324 a_4733_44350# a_1847_45528.t14 a_4651_44350# VDD.t2830 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2325 a_10389_45438# a_10111_45776# VSS.t852 VSS.t851 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X2326 VDAC_P.t401 C10_P_btm.t764 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2327 a_2043_43958# a_636_42870# a_2217_43834# VSS.t824 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2328 VDAC_N.t1515 C9_N_btm.t387 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2329 VDAC_P.t1519 C2_P_btm.t6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2330 VDAC_P.t773 C8_P_btm.t185 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2331 VDAC_N.t771 C10_N_btm.t743 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2332 VDD.t797 a_948_43806# a_1123_43780# VDD.t796 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2333 DATA[1].t7 a_663_47874# VDD.t805 VDD.t804 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2334 VDD.t2201 a_5655_43780# a_5715_45956# VDD.t2200 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2335 VDAC_N.t1513 C9_N_btm.t386 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2336 VDD.t987 a_9637_43560# a_9667_43301# VDD.t986 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2337 VDAC_P.t1517 C10_P_btm.t763 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2338 a_6673_45136# a_6455_44894# VSS.t929 VSS.t928 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2339 VDAC_P.t121 C9_P_btm.t366 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2340 VSS.t2642 a_9179_44592# a_9140_44466# VSS.t2641 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2341 VDAC_N.t399 C10_N_btm.t742 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2342 VDAC_P.t1515 C10_P_btm.t762 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2343 VDAC_P.t771 C10_P_btm.t761 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2344 VSS.t238 a_2587_44868.t10 a_2973_43582# VSS.t237 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2345 VDAC_N.t1511 C10_N_btm.t741 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2346 VDD.t452 a_7754_40130.t11 VDD.t451 VDD.t450 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.5
X2347 VDAC_P.t1513 C10_P_btm.t760 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2348 a_9973_46526# a_9547_46565# VDD.t2702 VDD.t2701 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X2349 VDAC_N.t769 C10_N_btm.t740 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2350 VDAC_N.t1509 C10_N_btm.t739 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2351 a_n2293_45956.t0 a_3328_44324# VSS.t1153 VSS.t1152 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2352 VDAC_P.t399 C10_P_btm.t759 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2353 VSS.t3812 C10_N_btm.t1068 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2354 a_6551_44894# a_6105_44894# a_6455_44894# VSS.t1610 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2355 VREF.t49 a_21276_30659.t6 C8_N_btm.t274 VDD.t2932 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2356 VSS.t2311 VSS.t2312 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2357 VDAC_N.t213 C8_N_btm.t185 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2358 VDAC_N.t1507 C10_N_btm.t737 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2359 a_1204_46758# a_n194_47222# a_1346_46565# VDD.t974 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2360 VDAC_N.t767 C10_N_btm.t736 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2361 VDAC_N.t1505 C8_N_btm.t184 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2362 VSS.t323 a_n1741_47596.t8 a_22399_44894# VSS.t322 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2363 VDAC_N.t397 C10_N_btm.t735 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2364 a_13622_43262# a_12545_43268# a_13460_43640# VDD.t813 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2365 VDAC_P.t1511 C9_P_btm.t365 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2366 VDAC_N.t1503 C9_N_btm.t385 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2367 VDAC_P.t769 C9_P_btm.t364 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2368 VSS.t1459 a_2687_45956# a_2621_45982# VSS.t1458 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2369 a_19921_31459.t0 a_22591_45982# VSS.t1086 VSS.t1085 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2370 VDAC_P.t1509 C8_P_btm.t184 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2371 VDAC_P.t213 C10_P_btm.t758 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2372 VDAC_N.t765 C9_N_btm.t384 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2373 VDAC_N.t1501 C8_N_btm.t183 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2374 VDAC_N.t51 C10_N_btm.t734 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2375 VSS.t2309 VSS.t2310 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2376 EN_VIN_BSTR_P.t0 VDD.t3185 a_n1586_35608# VSS.t3244 sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.9
X2377 VDAC_P.t1507 C10_P_btm.t183 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2378 VDAC_P.t767 C7_P_btm.t87 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2379 VDD.t1705 a_22959_47622# a_22812_30659.t3 VDD.t1136 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2380 a_19816_46642# a_19566_45670# a_19732_46642# VDD.t983 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2381 VDAC_P.t1505 C6_P_btm.t21 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2382 a_1343_38525.t3 a_1177_38525# VSS.t2667 VSS.t2666 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2383 VDAC_N.t1499 C6_N_btm.t24 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2384 DATA[1].t1 a_663_47874# VSS.t858 VSS.t857 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2385 VSS.t1097 a_20159_47588# a_13248_45956.t0 VSS.t1096 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X2386 VSS.t2140 a_14545_44569# a_10114_45276.t0 VSS.t2139 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2387 VDAC_P.t397 C8_P_btm.t183 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2388 VDAC_P.t1503 C10_P_btm.t374 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2389 a_11238_45982# a_10227_47214.t11 VSS.t332 VSS.t331 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2390 VDAC_N.t763 C10_N_btm.t733 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2391 VDAC_P.t765 VSS.t3357 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2392 VSS.t1254 a_9395_47044# a_4830_43958.t1 VSS.t1253 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X2393 a_8054_45144# a_5419_47258# VDD.t1525 VDD.t1524 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.14825 ps=1.34 w=0.42 l=0.15
X2394 VDAC_N.t1497 C10_N_btm.t732 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2395 VDAC_P.t1501 C10_P_btm.t756 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2396 a_4355_45438# a_135_43540.t25 VDD.t2864 VDD.t2863 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2397 VDD.t1662 a_6091_43780# a_1847_45528.t4 VDD.t1661 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2398 VSS.t2313 VSS.t2314 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2399 VDAC_N.t395 C10_N_btm.t731 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2400 a_5142_30651.t1 a_15008_42692# VSS.t2699 VSS.t2698 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2401 VDD.t817 a_22276_45412# a_18314_32299.t3 VDD.t816 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2402 VDAC_N.t1495 C10_N_btm.t730 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2403 VSS.t2319 VSS.t2320 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2404 VDAC_P.t51 C10_P_btm.t755 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2405 VDAC_P.t1499 C8_P_btm.t182 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2406 VDAC_N.t761 C10_N_btm.t729 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2407 VSS.t1795 a_4700_46134# a_4061_47044# VSS.t1794 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2408 VSS.t3807 C10_P_btm.t23 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2409 a_n2073_43806# a_n2103_43780.t10 VDD.t3030 VDD.t3029 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2410 VDAC_N.t1493 C10_N_btm.t728 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2411 a_22545_39429# a_22459_39581# VSS.t2167 VSS.t2166 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2412 a_21719_43244# a_n2293_45420.t4 VDD.t2866 VDD.t2865 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2413 a_18704_45982# a_17789_45982# a_18357_46224# VSS.t1498 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2414 VSS.t1449 a_n2472_45412# a_n2442_45438.t0 VSS.t1448 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2415 VDAC_N.t211 C10_N_btm.t727 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2416 VDAC_P.t763 C10_P_btm.t752 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2417 VDAC_N.t1491 C10_N_btm.t726 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2418 VSS.t879 a_17583_46500# a_16291_44914# VSS.t878 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X2419 a_601_44048# a_383_43806# VDD.t886 VDD.t885 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2420 VDAC_N.t759 C10_N_btm.t725 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2421 VDAC_N.t1489 C10_N_btm.t724 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2422 VDAC_P.t1497 C10_P_btm.t751 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2423 VDAC_P.t395 C8_P_btm.t181 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2424 VDAC_N.t393 C7_N_btm.t95 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2425 VDD.t827 a_20064_35138# a_21789_35634# VDD.t826 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2426 VDD.t2466 VSS.t3577 VDD.t2465 VDD.t2464 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2427 VDAC_P.t1495 C9_P_btm.t363 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2428 VSS.t2671 a_1177_38525# a_1343_38525.t0 VSS.t2670 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2429 a_16618_44670# a_16670_44324# a_n2103_44868.t0 VSS.t1266 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2430 VDAC_N.t1487 C10_N_btm.t723 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2431 a_11455_44576.t4 a_13635_43566# VDD.t1180 VDD.t1179 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2432 a_7569_44466# a_1429_47222.t9 a_7497_44466# VDD.t322 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X2433 VSS.t3484 VDD.t3221 VSS.t3483 VSS.t3482 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2434 VDAC_P.t761 C10_P_btm.t750 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2435 a_15860_45438# a_15549_47044.t10 a_15605_45438# VDD.t2987 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X2436 VDAC_N.t757 C9_N_btm.t383 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2437 VSS.t1485 a_3699_43780# a_1334_43494.t2 VSS.t1484 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2438 VDD.t1590 a_13113_43236# a_13003_43262# VDD.t1589 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2439 VDAC_N.t1485 C7_N_btm.t94 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2440 a_n1123_35174.t0 EN_VIN_BSTR_P.t7 VIN_P.t13 VSS.t549 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2441 VDAC_N.t119 C10_N_btm.t722 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2442 VDAC_P.t1493 C6_P_btm.t43 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2443 a_19771_43600# a_16475_45412# VDD.t1696 VDD.t1695 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2444 VSS.t958 a_9208_43494# a_9159_43262# VSS.t957 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2445 VDAC_N.t1483 C9_N_btm.t382 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2446 VDAC_P.t211 C10_P_btm.t749 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2447 VSS.t3212 VDD.t3173 VSS.t3211 VSS.t3210 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2448 VDAC_P.t1491 C7_P_btm.t86 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2449 VDD.t1386 a_2687_45956# a_2674_46348# VDD.t1385 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2450 VDAC_P.t759 C9_P_btm.t362 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2451 VDAC_N.t755 C10_N_btm.t721 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2452 VDAC_N.t1481 C10_N_btm.t720 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2453 VDD.t2783 a_18796_44728# a_18971_44654# VDD.t2782 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2454 a_7743_46904# a_7393_46532# a_7648_46892# VDD.t1213 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2455 VDAC_P.t1489 C10_P_btm.t748 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2456 VDAC_P.t393 C10_P_btm.t747 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2457 VDAC_N.t391 C9_N_btm.t381 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2458 a_369_45982# a_325_46224# a_203_45982# VSS.t887 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2459 VDAC_P.t1487 C9_P_btm.t361 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2460 VDAC_N.t1479 C10_N_btm.t719 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2461 VDAC_N.t753 C10_N_btm.t718 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2462 a_n2840_46500# a_n2661_46508.t9 VDD.t2647 VDD.t368 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2463 VDAC_N.t1477 C9_N_btm.t380 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2464 VDAC_P.t757 C10_P_btm.t746 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2465 VDAC_N.t209 C10_N_btm.t717 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2466 VDAC_P.t1485 C10_P_btm.t745 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2467 VDAC_N.t1475 C10_N_btm.t716 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2468 VDAC_P.t119 C9_P_btm.t360 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2469 C2_P_btm.t1 a_4000_42718.t6 VCM.t20 VSS.t297 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2470 VDAC_N.t751 C10_N_btm.t715 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2471 VDAC_P.t1483 C9_P_btm.t359 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2472 VDAC_P.t755 C10_P_btm.t744 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2473 VDAC_N.t1473 C10_N_btm.t714 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2474 VDD.t2211 a_5655_43780# a_8659_44324# VDD.t2210 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2475 VDAC_P.t1481 C9_P_btm.t358 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2476 VDAC_P.t391 C10_P_btm.t743 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2477 VSS.t3796 C9_N_btm.t535 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2478 VSS.t2617 a_9863_43958# a_9416_43530# VSS.t2616 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X2479 VSS.t176 a_135_43540.t33 a_4509_45804# VSS.t175 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2480 a_6091_43780# a_5655_43780# VDD.t2207 VDD.t2206 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2481 VDAC_N.t389 C10_N_btm.t713 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2482 VDD.t1672 a_16291_44914# a_17981_45438# VDD.t1671 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2483 VDAC_P.t1479 C8_P_btm.t180 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2484 VSS.t548 a_1203_42692.t32 a_20283_43262# VSS.t547 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2485 a_13460_43640# a_12545_43268# a_13113_43236# VSS.t871 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2486 VDD.t2322 VSS.t3677 VDD.t2321 VDD.t2320 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2487 VDD.t2078 a_6391_46219# a_6322_46348# VDD.t2077 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X2488 a_6105_44894# a_5939_44894# VSS.t1606 VSS.t1605 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2489 VDAC_P.t753 VSS.t3356 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2490 VDAC_P.t1477 C10_P_btm.t742 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2491 VDAC_N.t1471 C7_N_btm.t93 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2492 VDAC_P.t209 C9_P_btm.t357 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2493 VDAC_N.t749 C10_N_btm.t712 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2494 VSS.t2369 VSS.t2370 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2495 VDAC_N.t1469 C8_N_btm.t182 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2496 VSS.t2915 a_6485_44582.t16 a_8699_44894# VSS.t2914 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X2497 VDAC_P.t1475 C5_P_btm.t25 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2498 a_16085_45982# a_16128_46134# VDD.t732 VDD.t731 sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.345 ps=2.69 w=1 l=0.15
X2499 VDAC_N.t73 C8_N_btm.t181 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2500 VDAC_P.t751 C7_P_btm.t85 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2501 VDAC_P.t1473 C7_P_btm.t84 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2502 VSS.t889 a_161_44648# a_95_44716# VSS.t888 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2503 VDAC_N.t1467 VSS.t3326 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2504 a_510_42968# a_468_42870# a_428_42724# VDD.t834 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2505 VDAC_N.t747 C9_N_btm.t378 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2506 a_13214_45758# a_4908_45956# a_13464_45758# VSS.t1792 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2507 a_1083_45221# a_1053_45123.t11 a_1011_45221# VDD.t515 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2508 VDAC_P.t389 C10_P_btm.t741 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2509 VDAC_P.t1471 C9_P_btm.t356 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2510 VIN_P.t1 EN_VIN_BSTR_P.t14 C4_P_btm.t2 VSS.t556 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2511 C1_P_btm.t1 a_n1890_42718.t4 VSS.t365 VSS.t364 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2512 VDD.t2657 a_19187_42718# a_3990_30651.t3 VDD.t2656 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2513 VDAC_N.t1465 C10_N_btm.t711 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2514 VSS.t2087 EN_OFFSET_CAL.t0 a_16335_47614# VSS.t2086 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2515 VDAC_N.t387 C10_N_btm.t710 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2516 VDD.t63 a_1343_38525.t13 a_2684_37794# VDD.t61 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2517 VSS.t1320 a_6126_46642# a_n2661_45956.t1 VSS.t1319 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X2518 VDAC_P.t749 C10_P_btm.t740 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2519 VDAC_P.t1469 C10_P_btm.t739 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2520 a_n237_45454.t3 a_11971_46500# VDD.t2156 VDD.t2155 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2521 C3_P_btm.t1 a_n2810_45982.t4 VREF.t22 VDD.t2040 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2522 VSS.t396 a_1334_43494.t12 a_2332_44670# VSS.t395 sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.08775 ps=0.92 w=0.65 l=0.15
X2523 VDAC_N.t1463 C8_N_btm.t180 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2524 VSS.t192 a_135_43540.t47 a_4049_46892# VSS.t191 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2525 VDAC_N.t745 VSS.t3256 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2526 a_n126_44389# a_n172_44582# VDD.t1007 VDD.t1006 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2527 VSS.t1048 a_n2472_44324# a_n2442_44350.t0 VSS.t743 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2528 VDAC_P.t73 C6_P_btm.t42 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2529 VDD.t2295 VSS.t3795 VDD.t2294 VDD.t2293 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2530 VSS.t3228 VDD.t3179 VSS.t3227 VSS.t3226 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2531 VSS.t2619 a_8848_44868# a_n1925_47044.t1 VSS.t2618 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X2532 VDD.t2700 a_21303_42718# a_3222_30651.t3 VDD.t2699 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2533 VSS.t3675 C6_P_btm.t2 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2534 VDD.t2812 a_11455_44576.t13 a_12747_47070# VDD.t2811 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2535 VDAC_P.t1467 C9_P_btm.t355 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2536 VDD.t1527 a_5419_47258# a_5377_47320# VDD.t1526 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2537 VDD.t1059 a_15005_47222# a_10199_47846.t1 VDD.t1058 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X2538 VDAC_P.t747 C10_P_btm.t738 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2539 VDAC_N.t1461 C10_N_btm.t709 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2540 a_3754_38802# a_7754_38636# VSS.t693 sky130_fd_pr__res_high_po_0p35 l=18
X2541 VDD.t916 a_13266_45412# a_n1827_45412.t3 VDD.t915 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2542 VDAC_P.t1465 VSS.t3332 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2543 VDAC_N.t207 C5_N_btm.t23 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2544 VDD.t2469 VSS.t3793 VDD.t2468 VDD.t2467 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2545 VDD.t833 a_161_44648# a_191_44389# VDD.t832 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2546 VDAC_N.t1459 C10_N_btm.t708 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2547 VDD.t2689 a_5663_45982# a_8055_45491# VDD.t2688 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2548 VDAC_N.t743 C7_N_btm.t92 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2549 VDD.t2362 VSS.t3787 VDD.t2361 VDD.t2360 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2550 VDAC_P.t387 C6_P_btm.t40 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2551 VDAC_N.t1457 C10_N_btm.t707 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2552 VDAC_N.t385 C9_N_btm.t377 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2553 VDAC_P.t1463 C10_P_btm.t737 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2554 VDAC_P.t745 C8_P_btm.t179 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2555 VDAC_P.t1461 C9_P_btm.t354 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2556 VSS.t1418 a_4651_47614# DATA[3].t0 VSS.t1417 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2557 VSS.t2804 a_14766_45596.t9 a_15961_47980# VSS.t2803 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2558 VDAC_P.t207 C9_P_btm.t353 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2559 VDAC_P.t1459 C9_P_btm.t352 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2560 VSS.t3672 C9_P_btm.t13 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2561 VDAC_N.t1455 C10_N_btm.t706 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2562 VDD.t1634 a_82_45670# a_n1735_43236.t2 VDD.t1633 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2563 VDD.t2335 VSS.t3786 VDD.t2334 VDD.t2333 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2564 VDAC_N.t741 C9_N_btm.t376 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2565 VDAC_N.t1453 C9_N_btm.t375 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2566 VDAC_P.t743 C10_P_btm.t736 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2567 a_135_43540.t3 a_8391_47044# VSS.t1210 VSS.t1209 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X2568 a_8308_46904# a_7227_46532# a_7961_46500# VDD.t1210 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2569 VDD.t751 a_571_43566# a_558_43262# VDD.t750 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2570 VDD.t586 a_13273_44868.t13 a_17073_44056# VDD.t585 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2571 VDAC_N.t117 C10_N_btm.t705 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2572 VDAC_P.t1457 C8_P_btm.t178 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2573 VDD.t840 a_5663_42718# a_5840_42718.t2 VDD.t839 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2574 VDAC_P.t385 C10_P_btm.t735 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2575 VDAC_N.t1451 C9_N_btm.t374 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2576 VDAC_P.t1455 C9_P_btm.t349 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2577 VSS.t592 a_13524_46832.t7 a_17153_46846# VSS.t591 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2578 VDAC_N.t739 C8_N_btm.t179 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2579 VDAC_P.t741 C9_P_btm.t348 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2580 VDAC_P.t1453 C9_P_btm.t347 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2581 VDD.t1761 a_1387_42883# a_546_43100# VDD.t344 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2582 VDAC_N.t1449 C8_N_btm.t178 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2583 VSS.t3777 C8_N_btm.t268 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2584 a_n2103_43780.t1 a_3165_45982# VDD.t1393 VDD.t1392 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2585 VDAC_P.t117 C10_P_btm.t734 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2586 VDAC_P.t1451 C4_P_btm.t15 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2587 VDAC_P.t739 C10_P_btm.t733 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2588 a_1387_42883# a_134_42718.t7 VDD.t2808 VDD.t2807 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2589 VDAC_P.t1449 C10_P_btm.t732 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2590 VSS.t900 a_16513_42718# a_16703_42718# VSS.t899 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2591 VDD.t1243 a_12623_43780# a_12610_44172# VDD.t1242 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2592 VDD.t2486 VSS.t3616 VDD.t2485 VDD.t2290 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2593 a_n2661_44868# a_n2103_45412.t13 VDD.t2874 VDD.t2873 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2594 VDAC_P.t383 C10_P_btm.t731 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2595 VDAC_N.t383 C6_N_btm.t4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2596 VDAC_N.t1447 C9_N_btm.t373 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2597 VDAC_N.t737 C1_N_btm.t2 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2598 VSS.t1618 a_1123_43780# a_1581_43806.t2 VSS.t1617 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2599 VDAC_P.t1447 C9_P_btm.t346 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2600 VDAC_N.t1445 C8_N_btm.t176 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2601 VDAC_N.t205 C10_N_btm.t704 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2602 VSS.t2529 VSS.t2530 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2603 VDD.t2350 VSS.t3771 VDD.t2349 VDD.t2348 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2604 a_2424_46794.t0 a_11059_45956# VSS.t1077 VSS.t1076 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2605 VDAC_N.t1443 C8_N_btm.t175 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2606 VDAC_P.t737 VSS.t3355 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2607 a_6665_43582# a_2587_44868.t17 VSS.t244 VSS.t243 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X2608 VDAC_P.t1445 C7_P_btm.t83 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2609 VDAC_N.t735 C10_N_btm.t703 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2610 VDAC_P.t205 C9_P_btm.t345 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2611 VDAC_P.t1443 C9_P_btm.t344 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2612 VDAC_P.t735 C10_P_btm.t730 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2613 VSS.t3216 VDD.t3175 VSS.t3215 VSS.t3214 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2614 VDAC_P.t1441 C8_P_btm.t177 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2615 VSS.t2738 a_n1732_35090.t14 a_n1123_35174.t2 VSS.t2737 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2616 a_33_43806# a_n133_43806# VSS.t908 VSS.t907 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2617 VDAC_P.t381 C9_P_btm.t343 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2618 VDAC_N.t1441 C10_N_btm.t702 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2619 a_396_46904# a_n685_46532# a_49_46500# VDD.t1577 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2620 C6_P_btm.t71 a_n2810_46526.t4 VREF.t69 VDD.t3039 sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=0.35
X2621 VDAC_N.t381 C9_N_btm.t372 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2622 VDAC_P.t1439 VSS.t3338 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2623 a_7276_45670# a_n99_45438.t3 a_7418_45477# VDD.t2045 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2624 a_13273_44868.t0 a_18879_43780# VSS.t1630 VSS.t1629 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2625 VDAC_N.t1439 C8_N_btm.t174 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2626 VDAC_N.t733 C10_N_btm.t701 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2627 VDAC_P.t733 C10_P_btm.t729 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2628 VDAC_P.t1437 C9_P_btm.t342 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2629 VDAC_P.t39 C10_P_btm.t728 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2630 VSS.t3060 VDD.t3122 VSS.t3059 VSS.t3058 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2631 VDD.t100 a_927_42692.t16 a_2617_45144# VDD.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X2632 a_9863_47874# a_10199_47846.t2 VSS.t3005 VSS.t3004 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X2633 VDAC_N.t1437 C10_N_btm.t700 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2634 a_16576_44868# a_6104_45706.t6 VSS.t3008 VSS.t3007 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X2635 VDAC_N.t39 C10_N_btm.t699 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2636 VDAC_N.t1435 C10_N_btm.t698 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2637 VDAC_P.t1435 C10_P_btm.t727 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2638 VDAC_P.t731 C10_P_btm.t726 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2639 a_15871_47614# a_15691_47614# VDD.t864 VDD.t863 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X2640 VDD.t2463 VSS.t3664 VDD.t2462 VDD.t2461 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2641 VDAC_N.t731 C6_N_btm.t48 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2642 VDD.t778 a_14133_43780# a_14077_44133# VDD.t777 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X2643 VDAC_N.t1433 C8_N_btm.t173 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2644 VDAC_P.t1433 C7_P_btm.t82 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2645 VDAC_N.t379 C7_N_btm.t91 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2646 VDAC_P.t379 C5_P_btm.t15 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2647 VDAC_P.t1431 C10_P_btm.t725 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2648 a_16239_45804# a_1581_43806.t12 VSS.t2904 VSS.t2903 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X2649 VDD.t2880 a_14766_45596.t4 a_15871_47614# VDD.t2879 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2650 VDD.t838 a_8308_46904# a_8483_46830# VDD.t837 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2651 a_n1827_44868.t7 a_6485_44582.t20 VDD.t3021 VDD.t3020 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2652 VSS.t1735 a_16291_44914# a_18348_45758# VSS.t1734 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X2653 VSS.t1356 a_22959_45446# a_19679_31459.t1 VSS.t1355 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2654 VSS.t3590 C8_P_btm.t8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2655 a_16074_45046# a_16291_44914# VDD.t1676 VDD.t1675 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X2656 a_5569_44048# a_5351_43806# VSS.t913 VSS.t912 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2657 VDAC_P.t729 C10_P_btm.t724 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2658 a_3524_43806# a_2609_43806# a_3177_44048# VSS.t1224 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2659 a_10415_47846# a_2424_46794.t7 a_10589_47952# VSS.t2853 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2660 VDAC_P.t1429 C10_P_btm.t723 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2661 VDD.t7 a_10259_42870.t16 a_12287_44894# VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2662 VDD.t2876 a_14766_45596.t2 a_15321_46526# VDD.t2875 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2663 a_22031_45438# a_n2661_47044.t5 VSS.t2965 VSS.t2964 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2664 VDAC_N.t1431 C5_N_btm.t22 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2665 VDAC_N.t729 C9_N_btm.t371 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2666 VDAC_N.t1429 C8_N_btm.t172 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2667 VSS.t2944 SMPL.t13 a_n1732_35090.t2 VSS.t2943 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2668 VDAC_N.t203 C10_N_btm.t697 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2669 VDAC_N.t1427 C9_N_btm.t370 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2670 VDAC_P.t203 C10_P_btm.t722 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2671 VDAC_N.t727 C9_N_btm.t369 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2672 VDAC_N.t1425 C10_N_btm.t696 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2673 a_5447_43806# a_5001_43806# a_5351_43806# VSS.t1226 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2674 a_7393_43806# a_7227_43806# VSS.t1010 VSS.t1009 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2675 VDAC_P.t1427 C10_P_btm.t721 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2676 VDAC_P.t727 C10_P_btm.t720 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2677 VSS.t1700 a_3823_42718# a_4000_42718.t1 VSS.t1699 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2678 a_134_42718.t3 a_104_42692# VDD.t878 VDD.t877 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2679 VDAC_P.t1425 C9_P_btm.t341 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2680 VDAC_N.t377 C10_N_btm.t695 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2681 VDAC_P.t377 C9_P_btm.t340 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2682 VDAC_P.t1423 C9_P_btm.t339 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2683 a_5700_37509.t13 VDAC_N.t1423 a_8912_37509.t19 VDD.t2250 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2684 VDAC_P.t725 C10_P_btm.t719 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2685 VDAC_N.t725 C8_N_btm.t171 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2686 VSS.t823 a_636_42870# a_428_42724# VSS.t822 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X2687 VDAC_N.t1421 C10_N_btm.t694 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2688 VSS.t2068 a_5749_47222# a_5839_47070# VSS.t2067 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2689 VDAC_N.t115 VSS.t3292 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2690 a_16525_42968# a_12651_44576.t15 VDD.t2964 VDD.t2963 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2691 VDAC_P.t1421 VSS.t3337 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2692 a_15947_43262# a_15323_43268# a_15839_43640# VDD.t1371 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2693 VDD.t21 SMPL_ON_P.t9 a_n1605_47614# VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2694 VDD.t2653 a_18445_42718# a_19187_42718# VDD.t2652 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2695 VSS.t33 a_9521_45982.t12 a_12379_43268# VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2696 VSS.t810 a_4704_47044# a_4035_45609# VSS.t809 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X2697 VDAC_P.t115 C9_P_btm.t338 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2698 a_11514_46892# a_10227_47214.t10 VSS.t330 VSS.t329 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2699 VDAC_P.t1419 C10_P_btm.t718 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2700 VDAC_N.t1419 C8_N_btm.t170 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2701 VDAC_P.t723 C9_P_btm.t337 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2702 VDD.t855 a_396_46904# a_571_46830# VDD.t854 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2703 VDD.t1003 a_16750_46134# a_16703_45982# VDD.t1002 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.27 ps=2.54 w=1 l=0.15
X2704 VDAC_N.t723 C8_N_btm.t169 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2705 VDAC_P.t1417 C6_P_btm.t38 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2706 a_13561_44350# a_13023_44716# VDD.t1026 VDD.t1025 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X2707 VDAC_P.t375 C5_P_btm.t10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2708 VDAC_P.t1415 C7_P_btm.t81 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2709 VREF.t39 a_22812_30659.t14 C10_N_btm.t28 VDD.t526 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2710 VCM.t28 a_3222_30651.t13 VDAC_N.t5 VSS.t665 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2711 a_15579_44172# a_14955_43806# a_15471_43806# VDD.t1878 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2712 VDAC_P.t721 C9_P_btm.t336 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2713 VDAC_P.t1413 C10_P_btm.t717 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2714 a_6485_44582.t4 a_8483_43780# VDD.t906 VDD.t905 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2715 VDD.t2696 a_19633_43262# a_21303_42718# VDD.t2695 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2716 VDAC_P.t201 C10_P_btm.t716 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2717 VSS.t3513 VDD.t3231 VSS.t3512 VSS.t3178 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2718 a_n2661_43244# a_n2103_44324.t6 VDD.t3104 VDD.t3029 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2719 VDAC_N.t375 C6_N_btm.t47 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2720 VDAC_P.t1411 C8_P_btm.t84 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2721 VSS.t1773 a_1239_39587# COMP_P.t1 VSS.t1772 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2722 VDAC_P.t719 C10_P_btm.t715 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2723 VSS.t3032 VDD.t3112 VSS.t3031 VSS.t3030 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2724 VSS.t2450 VSS.t2451 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2725 a_3328_44324# a_3179_44403# VSS.t690 VSS.t689 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2726 VDAC_N.t1415 C9_N_btm.t368 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2727 a_3541_42718# a_1203_42692.t15 a_3553_42968# VDD.t477 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2728 VDAC_P.t1409 C8_P_btm.t174 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2729 a_17564_32305.t1 a_22959_43806# VSS.t2113 VSS.t1454 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2730 a_203_45982# a_n243_45982# a_107_45982# VSS.t2225 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2731 VDAC_P.t373 C10_P_btm.t714 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2732 VDAC_P.t1407 C10_P_btm.t713 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2733 VIN_N.t0 EN_VIN_BSTR_N.t15 C0_dummy_N_btm.t0 VSS.t444 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2734 VSS.t2201 a_11599_42883# a_9096_45276.t0 VSS.t2200 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2735 VDD.t1106 a_11427_43566# a_7557_43236.t5 VDD.t1105 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2736 a_33_43806# a_n133_43806# VDD.t853 VDD.t852 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2737 VDAC_N.t721 C10_N_btm.t693 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2738 VDAC_P.t717 C8_P_btm.t173 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2739 VDAC_N.t1413 C9_N_btm.t367 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2740 a_22717_37721# a_22459_39581# a_22609_38842# VSS.t2165 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2741 VDD.t2577 VSS.t3752 VDD.t2576 VDD.t2575 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2742 VDAC_N.t201 C10_N_btm.t692 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2743 a_3754_39964# a_7754_40130.t0 VSS.t693 sky130_fd_pr__res_high_po_0p35 l=18
X2744 a_20163_31459.t3 a_22223_46534# VDD.t1079 VDD.t1078 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2745 a_n1551_45412.t3 a_12438_45412# VDD.t747 VDD.t746 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2746 VSS.t3147 VDD.t3151 VSS.t3146 VSS.t3145 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2747 VDAC_P.t1405 C10_P_btm.t712 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2748 VDD.t2292 VSS.t3750 VDD.t2291 VDD.t2290 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2749 VDAC_N.t1411 C7_N_btm.t90 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2750 VDAC_P.t71 C10_P_btm.t711 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2751 VDAC_N.t719 C5_N_btm.t21 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2752 VSS.t921 a_11335_46830# a_11269_46904# VSS.t920 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2753 a_n2103_44324.t2 a_8204_45412# VDD.t2127 VDD.t2126 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X2754 VDAC_N.t1409 C8_N_btm.t168 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2755 VDAC_P.t1403 C8_P_btm.t172 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2756 VDAC_N.t373 C10_N_btm.t691 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2757 VDAC_N.t1407 C8_N_btm.t167 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2758 VSS.t3050 VDD.t3118 VSS.t3049 VSS.t3048 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2759 VDAC_P.t715 C7_P_btm.t38 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2760 DATA[1].t5 a_663_47874# VDD.t803 VDD.t802 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2761 a_21197_42718# a_21027_42718# VSS.t695 VSS.t694 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2762 VDAC_P.t1401 C7_P_btm.t79 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2763 a_n2472_46500# a_n2293_46508.t8 VDD.t114 VDD.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2764 a_2217_43834# a_n237_45454.t4 VSS.t467 VSS.t466 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X2765 a_6193_45982# a_5715_45956# VSS.t997 VSS.t996 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2766 VDAC_N.t717 C9_N_btm.t366 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2767 VDAC_P.t371 C10_P_btm.t710 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2768 VSS.t1123 a_22959_44358# a_17738_32299.t1 VSS.t1122 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2769 a_383_43806# a_33_43806# a_288_43806# VDD.t883 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2770 VDAC_P.t1399 C10_P_btm.t709 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2771 VDAC_P.t713 C10_P_btm.t708 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2772 VDAC_N.t1405 C10_N_btm.t690 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2773 VDAC_P.t1397 C10_P_btm.t707 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2774 VDAC_N.t71 C9_N_btm.t365 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2775 VDAC_N.t1403 C10_N_btm.t689 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2776 a_22031_44350# a_n2293_46508.t9 VSS.t110 VSS.t109 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2777 VSS.t2484 VSS.t2485 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2778 VDAC_P.t199 C10_P_btm.t706 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2779 VDAC_N.t715 C10_N_btm.t688 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2780 a_7393_43806# a_7227_43806# VDD.t952 VDD.t951 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2781 VDAC_P.t1395 C10_P_btm.t705 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2782 VSS.t1604 a_5473_43582# a_5663_42718# VSS.t1603 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2783 VSS.t1715 a_6091_43780# a_1847_45528.t3 VSS.t1714 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2784 a_18259_46500# a_18103_46768# a_18404_46526# VDD.t1799 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X2785 a_4338_37500.t6 VSS.t2488 VSS.t2490 VSS.t2489 sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.589 ps=4.42 w=1.9 l=0.15
X2786 a_n61_46526# a_n685_46532# a_n169_46904# VDD.t1578 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2787 VDAC_N.t1401 C10_N_btm.t687 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2788 VDAC_N.t371 C10_N_btm.t686 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2789 VDAC_P.t711 C9_P_btm.t335 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2790 a_18993_47320# a_10251_45454# a_17927_46195# VDD.t1296 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2791 VDAC_N.t1399 C10_N_btm.t685 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2792 VDAC_P.t1393 C9_P_btm.t334 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2793 VDAC_P.t369 C10_P_btm.t704 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2794 VDAC_P.t1391 C9_P_btm.t333 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2795 VDAC_P.t709 C10_P_btm.t703 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2796 VSS.t3066 VDD.t3124 VSS.t3065 VSS.t3064 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2797 a_4247_45816# a_3897_45444# a_4152_45804# VDD.t2124 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2798 VDAC_N.t713 C10_N_btm.t684 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2799 a_22399_44894# a_n1741_47596.t4 VSS.t319 VSS.t318 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2800 a_5700_37509.t12 VDAC_N.t1397 a_8912_37509.t18 VDD.t2242 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2801 VDAC_P.t1389 C10_P_btm.t702 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2802 VDD.t772 a_16561_45982# a_16671_47320# VDD.t771 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2803 VSS.t2497 VSS.t2498 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2804 VDAC_N.t199 C6_N_btm.t46 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2805 a_n126_44716# a_n172_44582# VSS.t1067 VSS.t1066 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2806 a_11795_47044# a_8727_47222.t7 VDD.t77 VDD.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2807 a_885_44868.t5 a_4322_46134# a_4703_44894# VSS.t1821 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2808 VDAC_N.t1395 C4_N_btm.t13 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2809 VDAC_N.t711 C10_N_btm.t683 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2810 DATA[1].t3 a_663_47874# VSS.t864 VSS.t863 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X2811 a_5129_45956# a_885_44868.t31 VSS.t2762 VSS.t2761 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2812 VDAC_N.t1393 C8_N_btm.t166 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2813 VDAC_P.t113 C8_P_btm.t171 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2814 VDAC_N.t369 C10_N_btm.t682 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2815 VDAC_N.t1391 C9_N_btm.t364 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2816 VDAC_P.t1387 C8_P_btm.t170 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2817 VDAC_P.t707 C10_P_btm.t701 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2818 VSS.t2830 EN_COMP.t6 a_1177_38525# VSS.t2829 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2819 VSS.t2248 a_5655_43780# a_5953_45982# VSS.t2247 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X2820 VDAC_N.t709 C10_N_btm.t681 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2821 a_13248_45956.t1 a_20159_47588# VSS.t1099 VSS.t1098 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2822 VDAC_N.t1389 C10_N_btm.t680 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2823 VDAC_P.t1385 C8_P_btm.t169 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2824 a_18905_44728# a_17715_44356# a_18796_44728# VSS.t702 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2825 a_12651_44576.t5 a_16579_43566# VDD.t1905 VDD.t1904 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2826 COMP_N.t0 a_1239_39043# VSS.t1781 VSS.t1768 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2827 VDAC_P.t367 C10_P_btm.t700 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2828 VDAC_N.t113 C10_N_btm.t679 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2829 VSS.t3609 C10_P_btm.t25 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2830 VDAC_N.t1387 C8_N_btm.t165 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2831 VDD.t443 a_7754_40130.t7 a_11206_38545.t2 VDD.t442 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X2832 a_1847_45528.t5 a_6091_43780# VDD.t1660 VDD.t1659 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2833 VDAC_N.t707 C10_N_btm.t678 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2834 VSS.t2281 VSS.t2282 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2835 a_18314_32299.t2 a_22276_45412# VDD.t815 VDD.t814 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2836 VDAC_N.t1385 C9_N_btm.t363 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2837 VDAC_N.t367 C8_N_btm.t164 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2838 VDAC_N.t1383 C10_N_btm.t677 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2839 VDAC_P.t1383 C9_P_btm.t332 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2840 a_n690_43494.t1 a_6635_47044# VSS.t2145 VSS.t2144 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2841 VDAC_P.t705 C9_P_btm.t331 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2842 VDD.t3028 a_n2103_43780.t8 a_n2073_43806# VDD.t3027 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2843 VDAC_N.t705 C10_N_btm.t676 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2844 VDAC_P.t1381 C4_P_btm.t14 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2845 a_7493_43582# a_2587_44868.t16 VSS.t242 VSS.t241 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X2846 VDD.t635 a_18879_45956# a_18866_46348# VDD.t634 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2847 a_n2840_47044# a_n2661_47044.t6 VDD.t3062 VDD.t3061 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2848 a_n2074_43262.t1 a_n2104_43236# VSS.t831 VSS.t830 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2849 VCM.t2 a_5142_30651.t6 C8_P_btm.t5 VSS.t122 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2850 a_21789_35634# a_20064_35138# VDD.t825 VDD.t824 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2851 VDAC_Pi.t1 a_3754_38470.t7 a_4338_37500.t2 VSS.t2841 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2852 VDAC_P.t197 C10_P_btm.t698 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2853 VDD.t1186 a_13635_43566# a_11455_44576.t5 VDD.t1185 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2854 VDAC_P.t1379 C10_P_btm.t697 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2855 VDAC_N.t1381 C4_N_btm.t11 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2856 VDD.t2332 VSS.t3573 VDD.t2331 VDD.t2296 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2857 VDD.t1907 a_16579_43566# a_12651_44576.t6 VDD.t1906 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2858 VDD.t2846 a_885_44868.t25 a_829_45221# VDD.t2845 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X2859 VDAC_N.t197 C7_N_btm.t89 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2860 VDAC_P.t703 C8_P_btm.t167 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2861 VSS.t1934 a_22123_44894# a_22591_44894# VSS.t1933 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2862 VDAC_N.t1379 C10_N_btm.t675 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2863 a_1334_43494.t3 a_3699_43780# VSS.t1483 VSS.t1482 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2864 VSS.t3726 C6_N_btm.t68 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2865 a_14011_44670# a_13469_44894# a_13915_44670# VSS.t835 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
X2866 VDAC_P.t1377 C10_P_btm.t696 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2867 VDAC_N.t703 C10_N_btm.t674 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2868 VDAC_P.t365 C10_P_btm.t695 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2869 VSS.t1500 a_20049_43262# a_22775_42718# VSS.t1499 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X2870 a_13458_32299.t3 a_21540_43236# VDD.t1892 VDD.t1891 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2871 VSS.t3508 VDD.t3229 VSS.t3507 VSS.t3506 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2872 VDAC_P.t1375 C8_P_btm.t166 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2873 w_11534_34010.t1 a_18394_35068.t8 EN_VIN_BSTR_N.t0 w_11534_34010.t0 sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2874 VDAC_N.t1377 C9_N_btm.t362 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2875 VDD.t2359 VSS.t3583 VDD.t2358 VDD.t2357 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2876 VDAC_P.t701 C9_P_btm.t330 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2877 VSS.t1372 a_10251_45454# a_17613_44894# VSS.t1371 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2878 VDAC_P.t1373 C7_P_btm.t78 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2879 VDAC_P.t49 C10_P_btm.t694 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2880 VDAC_N.t365 C10_N_btm.t673 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2881 a_15437_47044# a_15139_47730# VSS.t1350 VSS.t1349 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X2882 VDAC_P.t1371 C10_P_btm.t693 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2883 VSS.t3722 C9_N_btm.t531 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2884 VSS.t714 a_22469_41061# a_22717_37323# VSS.t713 sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2885 VDAC_N.t1375 C10_N_btm.t672 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2886 VDAC_N.t701 C9_N_btm.t360 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2887 VDAC_N.t1373 VSS.t3330 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2888 VDAC_N.t49 C9_N_btm.t359 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2889 a_n4515_30659.t3 a_n2288_47588# VDD.t1176 VDD.t1175 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2890 a_n1920_42692# a_n1741_42692# VSS.t2639 VSS.t2638 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2891 a_16750_46134# a_9521_45982.t16 VSS.t37 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X2892 VDD.t1732 a_1239_39043# COMP_N.t4 VDD.t1731 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2893 VSS.t1477 a_3699_43780# a_1334_43494.t0 VSS.t1476 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2894 VCM.t32 a_3222_30651.t11 VDAC_N.t3 VSS.t663 sky130_fd_pr__nfet_01v8_lvt ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X2895 a_15133_43582# a_1203_42692.t13 a_15145_43262# VDD.t474 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2896 a_18689_45412# a_18879_45956# VDD.t637 VDD.t636 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2897 VSS.t1447 a_11143_47588# a_8727_47222.t1 VSS.t1446 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X2898 VSS.t2859 a_n2293_45956.t9 a_22087_43244# VSS.t2858 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2899 VDAC_P.t699 C10_P_btm.t692 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2900 VSS.t3234 VDD.t3181 VSS.t3233 VSS.t3232 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2901 VDAC_N.t699 C10_N_btm.t671 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2902 VDAC_P.t1369 VSS.t3335 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2903 VSS.t2493 VSS.t2494 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2904 VDAC_P.t363 C10_P_btm.t691 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2905 VDAC_N.t1369 C9_N_btm.t358 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2906 a_n2103_44868.t7 a_6104_45706.t7 VDD.t3101 VDD.t3100 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2907 a_5700_37509.t11 VDAC_N.t363 a_8912_37509.t17 VDD.t2248 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2908 VDAC_N.t1367 C10_N_btm.t670 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2909 VDD.t2033 a_5923_31099.t6 a_8423_42718# VDD.t2032 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2910 VDAC_N.t697 C8_N_btm.t163 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2911 VDAC_P.t2 a_3222_30651.t9 VCM.t40 VSS.t661 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2912 VDAC_P.t697 C8_P_btm.t165 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2913 VDAC_N.t1365 C10_N_btm.t669 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2914 VDAC_N.t195 C10_N_btm.t668 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2915 VDAC_P.t1365 C9_P_btm.t329 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2916 VDAC_P.t195 C10_P_btm.t690 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2917 a_713_47044# a_380_47222# VSS.t1471 VSS.t1470 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2918 VDAC_N.t1363 C8_N_btm.t162 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2919 VDAC_P.t1363 C10_P_btm.t689 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2920 VDD.t868 a_11335_46830# a_11322_46526# VDD.t867 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2921 VDAC_N.t695 C9_N_btm.t357 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2922 VDAC_P.t695 C9_P_btm.t328 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2923 VDAC_P.t1361 C9_P_btm.t327 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2924 VREF.t19 a_20892_30659.t4 C6_N_btm.t1 VDD.t602 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=0.35
X2925 VDD.t1448 a_6631_44582# a_6491_44716# VDD.t1447 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X2926 VDD.t1110 a_11427_43566# a_11414_43262# VDD.t1109 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2927 a_7429_47044# a_885_44868.t21 VSS.t2752 VSS.t2751 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2928 a_3437_46532# a_3271_46532# VSS.t1679 VSS.t1678 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2929 VDAC_N.t1361 C10_N_btm.t667 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2930 VDAC_N.t361 C10_N_btm.t666 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2931 VSS.t992 a_22031_44350# a_22959_43270# VSS.t991 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2932 a_13667_32299.t0 a_21855_42718# VSS.t1544 VSS.t1543 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2933 a_n2293_44332# a_n1551_45412.t11 VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2934 VSS.t3430 VDD.t3201 VSS.t3429 VSS.t3058 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2935 a_10427_46348# a_10227_47214.t34 VDD.t134 VDD.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2936 VDAC_N.t1359 C7_N_btm.t88 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2937 VSS.t1740 a_21629_47833# a_14766_45596.t0 VSS.t1739 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2938 VDAC_P.t361 C8_P_btm.t164 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2939 a_n2840_47044# a_n2661_47044.t7 VSS.t2966 VSS.t2559 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2940 a_16057_43236# a_15839_43640# VSS.t1704 VSS.t1703 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2941 C9_N_btm.t8 a_21788_30659.t7 VREF.t26 VDD.t2054 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2942 VDAC_N.t2 a_3222_30651.t7 VCM.t35 VSS.t659 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2943 a_21629_47833# DEBUG_MUX[2].t1 VSS.t2726 VSS.t2725 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2944 a_18357_44048# a_18139_43806# VDD.t1888 VDD.t1887 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2945 a_n1925_47044.t0 a_8848_44868# VSS.t2621 VSS.t2620 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2946 VSS.t716 a_12427_42883# a_10844_44364# VSS.t715 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2947 VDAC_N.t1357 C10_N_btm.t665 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2948 VDAC_N.t111 C10_N_btm.t664 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2949 VDAC_P.t1359 C9_P_btm.t326 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2950 a_22705_38842# a_22521_40491# a_22609_38842# VDD.t1474 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2951 C7_N_btm.t0 a_21020_30659.t4 VREF.t8 VDD.t254 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2952 VDAC_P.t693 C10_P_btm.t688 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2953 VDAC_P.t1357 C10_P_btm.t687 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2954 VDAC_P.t111 C7_P_btm.t77 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2955 VDAC_N.t1355 C10_N_btm.t663 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2956 VDD.t1806 a_22400_42718# a_22521_40491# VDD.t1802 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2957 VDAC_P.t1355 C9_P_btm.t325 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2958 C9_N_btm.t538 a_4758_30651.t8 VCM.t59 VSS.t2989 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2959 a_15471_43806# a_14955_43806# a_15376_43806# VSS.t1932 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2960 a_n1827_45412.t2 a_13266_45412# VDD.t914 VDD.t913 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2961 VDAC_N.t691 C5_N_btm.t20 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2962 VDAC_N.t1353 C10_N_btm.t662 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2963 VDAC_P.t691 C9_P_btm.t158 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2964 VDAC_P.t1353 C10_P_btm.t686 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2965 VSS.t720 a_5536_44324# a_n1827_44324.t1 VSS.t719 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X2966 a_12427_42883# a_5542_30651.t7 VSS.t2969 VSS.t2968 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2967 a_14014_46842# a_13427_46756# a_13930_46842# VSS.t1525 sky130_fd_pr__nfet_01v8 ad=0.10795 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2968 VDAC_N.t359 C10_N_btm.t661 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2969 VSS.t3718 C8_N_btm.t269 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2970 VDAC_P.t359 C9_P_btm.t323 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2971 VIN_N.t14 EN_VIN_BSTR_N.t17 a_11730_34132.t2 VSS.t446 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2972 VDAC_N.t1351 C9_N_btm.t353 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2973 VDAC_N.t689 C10_N_btm.t660 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2974 VDAC_N.t1349 C10_N_btm.t659 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2975 VDAC_P.t1351 C10_P_btm.t685 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2976 VDAC_N.t193 C9_N_btm.t352 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2977 VDAC_N.t1347 C7_N_btm.t87 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2978 VDAC_P.t689 C9_P_btm.t322 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2979 a_n2109_42692.t1 a_15187_44868# VSS.t1271 VSS.t1270 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2980 VDAC_P.t1349 C8_P_btm.t163 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2981 VDD.t23 a_9521_45982.t4 a_10079_46532# VDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2982 VDD.t2574 VSS.t3717 VDD.t2573 VDD.t2572 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2983 VDAC_N.t687 C10_N_btm.t658 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2984 VDAC_Ni.t0 a_7754_38636# VSS.t693 sky130_fd_pr__res_high_po_0p35 l=18
X2985 VDAC_P.t193 C10_P_btm.t684 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2986 VSS.t1223 a_1663_45046# a_380_47222# VSS.t1222 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2987 VSS.t382 a_1429_47222.t10 a_1387_44582# VSS.t381 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2988 VDAC_P.t1347 C10_P_btm.t683 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2989 a_22821_39429# a_22400_42718# VSS.t1846 VSS.t1845 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2990 a_6280_46642# a_5382_44582# a_6208_46642# VDD.t2025 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2991 VSS.t3200 VDD.t3169 VSS.t3199 VSS.t3198 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2992 VDAC_N.t1345 C9_N_btm.t351 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2993 VDAC_P.t687 C9_P_btm.t321 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2994 VDD.t1108 a_11427_43566# a_7557_43236.t6 VDD.t1107 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2995 VDAC_P.t1345 C10_P_btm.t682 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X2996 a_6954_46348# a_6235_46124# a_6391_46219# VSS.t2274 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2997 a_558_43262# a_n519_43268# a_396_43640# VDD.t1699 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2998 a_n1827_45412.t6 a_11455_44576.t16 VDD.t2816 VDD.t2815 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2999 VDAC_N.t357 C8_N_btm.t160 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3000 VDAC_P.t357 C10_P_btm.t681 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3001 VDAC_P.t1343 C5_P_btm.t7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3002 a_16513_42718# a_1203_42692.t11 a_16525_42968# VDD.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3003 a_3524_43806# a_2443_43806# a_3177_44048# VDD.t2061 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3004 VDAC_N.t1343 VSS.t3329 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3005 a_9637_43560# a_9304_43494# VSS.t724 VSS.t723 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3006 VDAC_P.t685 C10_P_btm.t680 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3007 VDAC_N.t685 C10_N_btm.t657 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3008 a_3830_44670# a_3882_44324# a_n2103_43780.t4 VSS.t2039 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3009 VDAC_N.t1341 C9_N_btm.t350 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3010 VDAC_P.t1341 C10_P_btm.t679 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3011 a_6661_44716# a_6631_44582# a_6573_44716# VSS.t1505 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X3012 a_19566_45670# a_19555_42718# VSS.t1065 VSS.t1064 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3013 a_15321_46526# a_14757_45982# VDD.t1221 VDD.t1220 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X3014 VDAC_N.t69 C10_N_btm.t656 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3015 DATA[2].t3 a_2351_47614# VSS.t2052 VSS.t2051 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X3016 a_8500_45554# a_8192_44874# a_8416_45554# VDD.t2231 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3017 VDAC_N.t1339 C7_N_btm.t86 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3018 VDAC_N.t683 C10_N_btm.t655 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3019 VSS.t1075 a_8530_39574# a_3754_38470.t0 VSS.t1074 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3020 VSS.t1571 a_10901_42718# a_11183_42718# VSS.t1570 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3021 VDAC_P.t69 C10_P_btm.t678 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3022 VDAC_P.t1339 C10_P_btm.t677 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3023 VDD.t2871 a_n2103_45412.t8 a_n2661_44868# VDD.t2870 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3024 VDAC_N.t1337 C10_N_btm.t654 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3025 VDAC_N.t355 VSS.t3304 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3026 VDAC_P.t683 C9_P_btm.t320 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3027 VDAC_N.t1335 C10_N_btm.t653 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3028 VDAC_N.t681 C8_N_btm.t159 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3029 VDAC_N.t1333 C10_N_btm.t652 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3030 a_18044_45982# a_17927_46195# VDD.t1894 VDD.t1893 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3031 a_n1827_44868.t3 a_8850_45412# a_8798_45758# VSS.t729 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3032 VDAC_N.t191 C9_N_btm.t349 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3033 VDAC_N.t1331 C10_N_btm.t651 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3034 VDAC_P.t1337 C10_P_btm.t676 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3035 VDAC_P.t355 C10_P_btm.t675 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3036 VDAC_P.t1335 C8_P_btm.t162 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3037 VDAC_P.t681 C8_P_btm.t161 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3038 VDAC_N.t679 C10_N_btm.t650 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3039 a_12800_43628# a_12683_43433# VDD.t1486 VDD.t1485 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3040 VDAC_N.t1329 C8_N_btm.t158 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3041 a_n2442_43262.t3 a_n2472_43236# VDD.t2141 VDD.t2140 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3042 a_n2661_43780# a_n1551_44324.t13 VDD.t130 VDD.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3043 a_21540_43236# a_21719_43244# VSS.t1033 VSS.t1032 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3044 VDAC_P.t1333 C5_P_btm.t12 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3045 VDAC_P.t191 C10_P_btm.t674 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3046 C7_P_btm.t0 EN_VIN_BSTR_P.t12 VIN_P.t15 VSS.t554 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3047 VDAC_N.t353 C9_N_btm.t348 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3048 VSS.t3639 C8_P_btm.t12 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3049 a_1209_47588# a_1083_45221# VDD.t836 VDD.t835 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X3050 VDAC_P.t1331 C8_P_btm.t160 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3051 VDAC_N.t1327 C10_N_btm.t649 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3052 VSS.t1427 a_4993_47044# a_6126_46642# VSS.t1426 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3053 VSS.t369 a_n2442_44894.t5 C9_P_btm.t1 VSS.t368 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3054 VDAC_N.t677 C9_N_btm.t347 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3055 VDAC_P.t679 C10_P_btm.t673 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3056 VDD.t2035 START.t0 a_14587_47614# VDD.t2034 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3057 a_17981_45438# a_15730_45670.t20 a_15549_47044.t1 VDD.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3058 VDD.t1710 a_21755_44350# a_22223_44358# VDD.t1709 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3059 a_18348_45758# a_18282_45670# a_12127_46744# VSS.t1765 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3060 VDAC_N.t1325 C7_N_btm.t85 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3061 a_n2074_47070.t1 a_n2104_47044# VSS.t734 VSS.t733 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3062 VSS.t521 a_1203_42692.t10 a_18445_42718# VSS.t520 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3063 VDAC_N.t109 C10_N_btm.t648 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3064 VSS.t3715 C8_P_btm.t11 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3065 a_19437_31459.t3 a_22959_44894# VDD.t2727 VDD.t1286 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3066 VDAC_P.t1329 C10_P_btm.t672 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3067 a_10589_47952# a_n237_45454.t8 VSS.t473 VSS.t472 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X3068 VDAC_N.t1323 C10_N_btm.t647 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3069 VDAC_P.t353 C10_P_btm.t671 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3070 a_10813_46500# a_10595_46904# VSS.t2155 VSS.t2154 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3071 VDAC_P.t1327 C9_P_btm.t319 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3072 VDAC_N.t675 C10_N_btm.t646 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3073 VDAC_N.t1321 C10_N_btm.t645 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3074 VSS.t3222 VDD.t3177 VSS.t3221 VSS.t3220 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3075 a_10069_42718# a_7557_43236.t26 VSS.t232 VSS.t231 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3076 VDD.t616 a_3524_43806# a_3699_43780# VDD.t615 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3077 VDAC_P.t677 C9_P_btm.t318 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3078 VDAC_P.t1325 C10_P_btm.t670 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3079 VDD.t2381 VSS.t3711 VDD.t2380 VDD.t2379 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3080 VDAC_N.t351 C10_N_btm.t644 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3081 a_10905_43236# a_10687_43640# VSS.t2149 VSS.t2148 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3082 VDAC_P.t109 C10_P_btm.t669 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3083 VDAC_P.t1323 C10_P_btm.t668 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3084 VDAC_N.t1319 C9_N_btm.t346 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3085 VSS.t1534 a_7842_44868# a_n2293_46508.t0 VSS.t1533 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X3086 VDAC_P.t675 C10_P_btm.t667 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3087 VDAC_N.t673 C8_N_btm.t157 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3088 VDAC_N.t1317 C10_N_btm.t643 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3089 VDAC_N.t189 C10_N_btm.t642 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3090 VSS.t204 a_4830_43958.t6 a_7227_43806# VSS.t203 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3091 VDAC_N.t1315 C10_N_btm.t641 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3092 VDAC_P.t1321 C9_P_btm.t317 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3093 VDAC_P.t351 C10_P_btm.t666 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3094 a_18796_44728# a_17881_44356# a_18449_44324# VSS.t2682 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3095 VDAC_N.t671 C9_N_btm.t345 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3096 a_4703_44894# a_2587_44868.t28 VSS.t272 VSS.t271 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3097 VDAC_N.t1313 C8_N_btm.t156 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3098 VDAC_P.t1319 C9_P_btm.t316 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3099 a_18319_44868# a_18495_44868# a_18447_44894# VSS.t1736 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X3100 VDAC_P.t673 C7_P_btm.t76 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3101 a_14087_32299.t1 a_22223_43270# VSS.t738 VSS.t737 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3102 VDAC_N.t349 C8_N_btm.t155 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3103 VSS.t2373 VSS.t2374 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3104 VDAC_P.t1317 C4_P_btm.t19 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3105 VSS.t740 a_14819_44582# a_14133_43780# VSS.t739 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X3106 VDAC_P.t189 C7_P_btm.t75 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3107 a_6886_37412# VDAC_Pi.t10 VDD.t3069 VSS.t2971 sky130_fd_pr__nfet_03v3_nvt ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X3108 VCM.t60 a_4758_30651.t9 C9_N_btm.t539 VSS.t2990 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3109 VIN_N.t8 EN_VIN_BSTR_N.t12 C8_N_btm.t3 VSS.t441 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3110 a_17789_43806# a_17623_43806# VSS.t1936 VSS.t1935 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3111 a_15489_43268# a_15323_43268# VSS.t1441 VSS.t1440 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3112 VDAC_P.t1315 C8_P_btm.t159 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3113 VDAC_N.t1311 C10_N_btm.t640 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3114 VDAC_N.t669 C9_N_btm.t343 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3115 VDAC_P.t671 VSS.t3367 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3116 VDAC_N.t1309 C9_N_btm.t342 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3117 VDAC_P.t1313 C10_P_btm.t665 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3118 C10_P_btm.t1059 a_n4515_30659.t7 VREF.t56 VDD.t2993 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3119 VSS.t3543 VDD.t3241 VSS.t3542 VSS.t3541 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3120 VDAC_P.t349 C10_P_btm.t663 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3121 a_12800_43628# a_12683_43433# VSS.t1550 VSS.t1549 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3122 VDAC_N.t33 C9_N_btm.t341 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3123 VDAC_N.t1307 C10_N_btm.t639 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3124 VDAC_N.t667 C10_N_btm.t638 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3125 VDAC_P.t1311 C10_P_btm.t662 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3126 a_n2442_44894.t1 a_n2472_44868# VSS.t742 VSS.t741 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3127 VDAC_N.t1305 C10_N_btm.t637 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3128 C9_P_btm.t10 a_n2467_30659.t9 VREF.t16 VDD.t582 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3129 VDAC_P.t669 C10_P_btm.t661 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3130 VDAC_P.t1309 C10_P_btm.t660 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3131 VDD.t2795 a_22465_38541# a_22521_39947# VDD.t2794 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3132 VDAC_P.t33 C10_P_btm.t659 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3133 DATA[4].t5 a_5847_47614# VDD.t1864 VDD.t1863 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3134 VDAC_P.t1307 C10_P_btm.t658 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3135 a_n193_47098# a_n194_47222# VDD.t976 VDD.t975 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3136 VDD.t3106 a_n2103_44324.t8 a_n2661_43244# VDD.t3027 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3137 VDAC_N.t347 C9_N_btm.t340 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3138 VDAC_N.t1303 C10_N_btm.t636 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3139 a_n2472_47044# a_n2293_47044.t6 VDD.t470 VDD.t469 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3140 VDAC_N.t665 C10_N_btm.t635 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3141 VDAC_P.t667 C10_P_btm.t657 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3142 COMP_P.t3 a_1239_39587# VSS.t1767 VSS.t1766 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3143 VSS.t3602 C10_N_btm.t1070 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3144 VDAC_N.t1301 C10_N_btm.t633 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3145 VDAC_P.t1305 C8_P_btm.t158 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3146 VDAC_P.t347 C10_P_btm.t656 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3147 a_18457_42968# a_13273_44868.t10 VDD.t612 VDD.t611 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3148 VDAC_P.t1303 C10_P_btm.t655 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3149 VDAC_N.t187 C10_N_btm.t632 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3150 VSS.t2078 a_15309_45438# a_15192_46500# VSS.t2077 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3151 a_7372_45670# a_7415_44466# VSS.t1333 VSS.t1332 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X3152 VIN_P.t9 EN_VIN_BSTR_P.t8 C10_P_btm.t8 VSS.t550 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3153 a_9521_45982.t3 a_9343_45982# VDD.t1462 VDD.t1461 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X3154 a_n1429_43262# a_n1459_43236.t8 VSS.t594 VSS.t593 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3155 a_16750_46134# a_1429_47222.t12 VSS.t384 VSS.t383 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0567 ps=0.69 w=0.42 l=0.15
X3156 VDAC_P.t665 C10_P_btm.t654 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3157 VDAC_N.t1299 C5_N_btm.t33 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3158 VDAC_N.t663 C9_N_btm.t339 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3159 VDAC_N.t1297 C8_N_btm.t154 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3160 VDAC_P.t1301 C8_P_btm.t157 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3161 a_4651_44350# a_2755_43494.t14 a_4733_44670# VSS.t512 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3162 VDAC_N.t345 C8_N_btm.t153 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3163 VDAC_N.t1295 C10_N_btm.t631 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3164 VDAC_P.t187 C6_P_btm.t37 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3165 C8_N_btm.t2 EN_VIN_BSTR_N.t8 VIN_N.t7 VSS.t437 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3166 VSS.t1799 a_4527_46830# a_4322_46134# VSS.t1798 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3167 VDAC_N.t661 C10_N_btm.t630 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3168 a_10037_43834# a_n237_45454.t7 VSS.t471 VSS.t470 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X3169 VDAC_P.t1299 C9_P_btm.t315 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3170 VDAC_N.t1293 C10_N_btm.t629 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3171 VDAC_P.t663 VSS.t3366 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3172 a_2209_45982# a_2165_46224# a_2043_45982# VSS.t2589 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3173 a_n2103_44868.t5 a_12651_44576.t16 VDD.t2966 VDD.t2965 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3174 VDAC_N.t107 C10_N_btm.t628 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3175 VDAC_N.t1291 C8_N_btm.t152 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3176 VDAC_P.t1297 C10_P_btm.t653 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3177 VDAC_N.t659 C9_N_btm.t338 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3178 VDAC_P.t345 C9_P_btm.t314 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3179 VDAC_N.t1289 C9_N_btm.t337 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3180 a_7851_46526# a_135_43540.t20 VDD.t2860 VDD.t2859 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3181 VDD.t890 a_n2840_43236# a_n2810_43262.t3 VDD.t889 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3182 a_11269_46904# a_10079_46532# a_11160_46904# VSS.t2253 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3183 VSS.t2432 VSS.t2433 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3184 VDAC_N.t343 C10_N_btm.t627 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3185 VDD.t682 a_22223_43494# a_22223_43270# VDD.t681 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3186 VDD.t1722 a_10596_44324# a_n2661_46508.t0 VDD.t1721 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X3187 VDAC_P.t1295 C10_P_btm.t652 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3188 VDAC_N.t1287 C10_N_btm.t626 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3189 a_n1552_42692# a_n1429_43262# VSS.t954 VSS.t953 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3190 VDAC_P.t661 C10_P_btm.t651 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3191 VDAC_P.t1293 C9_P_btm.t313 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3192 VDAC_N.t657 C10_N_btm.t625 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3193 VDAC_P.t107 C10_P_btm.t650 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3194 VSS.t1507 a_6631_44582# a_6953_43582# VSS.t1506 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3195 VDAC_N.t1285 C9_N_btm.t336 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3196 VDAC_P.t1291 C10_P_btm.t649 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3197 VDAC_P.t659 C9_P_btm.t312 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3198 VDAC_N.t185 C10_N_btm.t624 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3199 VSS.t2371 VSS.t2372 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3200 VDAC_P.t1289 C9_P_btm.t311 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3201 VDAC_P.t343 C10_P_btm.t648 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3202 a_9637_43560# a_9304_43494# VDD.t652 VDD.t651 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3203 VDAC_N.t1283 C10_N_btm.t623 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3204 VREF.t9 a_21020_30659.t5 C7_N_btm.t1 VDD.t255 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3205 VDD.t204 a_4830_43958.t12 a_7227_43806# VDD.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3206 a_1847_45528.t2 a_6091_43780# VSS.t1721 VSS.t1720 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3207 VDD.t1554 a_7311_47614# a_7595_47614# VDD.t1553 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3208 VSS.t2349 VSS.t2350 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3209 VDAC_P.t1287 VSS.t3342 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3210 VDAC_P.t657 C10_P_btm.t647 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3211 VDAC_P.t1285 C10_P_btm.t646 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3212 VSS.t2686 a_22775_42718# a_22465_38541# VSS.t2685 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3213 VDAC_N.t655 C7_N_btm.t84 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3214 VDD.t2158 a_11971_46500# a_n237_45454.t2 VDD.t2157 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3215 a_1387_45670# a_1334_43494.t19 VSS.t400 VSS.t399 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X3216 VDAC_N.t1281 C10_N_btm.t622 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3217 VDAC_N.t341 C3_N_btm.t8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3218 VDAC_N.t1279 C8_N_btm.t151 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3219 VDAC_P.t185 C8_P_btm.t156 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3220 a_15467_47320# a_15437_47044# a_15005_47222# VDD.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
X3221 VSS.t2285 VSS.t2286 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3222 VDAC_N.t653 C9_N_btm.t335 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3223 VDAC_P.t1283 C5_P_btm.t26 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3224 VDAC_N.t1277 C8_N_btm.t150 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3225 VSS.t2293 VSS.t2294 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3226 VDAC_P.t655 C7_P_btm.t74 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3227 a_12545_43268# a_12379_43268# VDD.t1097 VDD.t1096 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3228 VDD.t2674 a_11415_45670# a_9349_46539# VDD.t2673 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X3229 VDAC_N.t67 VSS.t3289 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3230 a_17789_43806# a_17623_43806# VDD.t1884 VDD.t1883 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3231 VDAC_N.t1275 C9_N_btm.t334 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3232 VDAC_P.t1281 C9_P_btm.t310 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3233 a_9335_44324# a_9140_44466# a_9645_44716# VSS.t1110 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X3234 a_4703_44894# a_4322_46134# a_885_44868.t6 VSS.t1822 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3235 VDAC_N.t651 C10_N_btm.t621 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3236 a_n61_46526# a_135_43540.t13 VDD.t2908 VDD.t2907 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3237 VDAC_N.t1273 C9_N_btm.t333 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3238 VDAC_P.t341 C10_P_btm.t645 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3239 a_1161_42968# a_927_42692.t14 VDD.t96 VDD.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3240 a_11507_47833# RST_Z.t2 VSS.t2819 VSS.t2818 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3241 a_5139_44019# a_4651_44350# VSS.t1834 VSS.t1833 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3242 VDAC_P.t1279 C9_P_btm.t309 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3243 a_288_43806# a_171_44019# VSS.t1517 VSS.t1516 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3244 VDD.t2427 VSS.t3631 VDD.t2426 VDD.t2425 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3245 VSS.t256 a_18314_32299.t9 C10_N_btm.t5 VSS.t255 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3246 VDAC_N.t339 C10_N_btm.t618 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3247 a_n2472_47044# a_n2293_47044.t7 VSS.t524 VSS.t105 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3248 VDAC_P.t653 VSS.t3364 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3249 VDAC_P.t1277 C10_P_btm.t644 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3250 a_10337_43268# a_10171_43268# VSS.t2180 VSS.t2179 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3251 VSS.t3183 VDD.t3163 VSS.t3182 VSS.t3181 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3252 VDAC_N.t1271 C8_N_btm.t149 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3253 VSS.t2629 a_n2038_35608# SMPL_ON_P.t3 VSS.t2628 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3254 VDAC_N.t649 C8_N_btm.t148 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3255 a_8150_45144# a_5663_45982# a_8054_45144# VDD.t2690 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3256 VDAC_P.t67 C6_P_btm.t36 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3257 a_12427_46758# a_12699_46616# a_12657_46642# VDD.t1827 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3258 VDAC_N.t1269 VSS.t3269 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3259 a_3895_46526# a_135_43540.t11 VDD.t2906 VDD.t2905 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3260 VDAC_P.t1275 C6_P_btm.t35 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3261 a_3990_30651.t1 a_19187_42718# VSS.t2566 VSS.t2565 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3262 VDD.t472 a_n2293_47044.t8 a_22123_44894# VDD.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3263 VCM.t7 a_3990_30651.t7 C10_P_btm.t0 VSS.t280 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3264 a_20892_30659.t2 a_22959_46534# VDD.t2731 VDD.t1855 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3265 VSS.t1017 a_9943_45046# a_9304_43494# VSS.t1016 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X3266 VDAC_P.t651 C6_P_btm.t34 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3267 a_n53_44363.t1 a_1115_47044# VSS.t1145 VSS.t1144 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3268 VDAC_P.t1273 C9_P_btm.t308 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3269 VSS.t1337 a_16102_47044# a_16046_47070# VSS.t1336 sky130_fd_pr__nfet_01v8 ad=0.258375 pd=1.445 as=0.091 ps=0.93 w=0.65 l=0.15
X3270 VSS.t1375 a_n2840_44868# a_n2810_44894.t0 VSS.t937 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3271 VDAC_P.t339 C10_P_btm.t643 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3272 VDAC_N.t183 C10_N_btm.t617 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3273 VDAC_N.t1267 C5_N_btm.t18 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3274 a_18133_47235# a_4830_43958.t14 VDD.t206 VDD.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3275 a_8862_44482# a_9140_44466# a_9096_44350# VDD.t1049 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X3276 a_18866_46348# a_17789_45982# a_18704_45982# VDD.t1431 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3277 VDAC_N.t647 C6_N_btm.t44 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3278 VDAC_N.t1265 C9_N_btm.t332 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3279 a_14204_44350# a_13725_44350# VSS.t1887 VSS.t1886 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.112125 ps=0.995 w=0.65 l=0.15
X3280 VDAC_P.t1271 C8_P_btm.t155 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3281 VSS.t833 a_n2104_43236# a_n2074_43262.t0 VSS.t832 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3282 a_3830_44670# a_3165_45982# a_4080_44670# VSS.t1466 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3283 VDD.t2755 a_11795_47044# a_10227_47214.t7 VDD.t2754 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3284 a_4733_44350# a_4322_46134# VDD.t1791 VDD.t1790 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3285 VDAC_N.t337 C10_N_btm.t616 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3286 a_3222_30651.t1 a_21303_42718# VSS.t2604 VSS.t2603 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3287 a_10150_47322# a_10467_47212# a_10425_47070# VSS.t2171 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X3288 VDAC_P.t649 C8_P_btm.t154 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3289 a_n2810_45982.t2 a_n2840_45956# VDD.t1596 VDD.t1595 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3290 VDAC_N.t1263 C9_N_btm.t331 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3291 VDAC_P.t1269 C10_P_btm.t642 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3292 VDAC_P.t183 C8_P_btm.t153 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3293 VDD.t1476 a_21847_43806# a_21855_42718# VDD.t1475 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3294 a_6563_45260# a_5655_43780# VDD.t2203 VDD.t2202 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3295 VDAC_P.t1267 C9_P_btm.t307 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3296 VDAC_P.t647 C9_P_btm.t306 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3297 VDAC_N.t645 C10_N_btm.t615 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3298 VDD.t1708 a_49_43236# a_n61_43262# VDD.t1707 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3299 VDAC_N.t1261 C9_N_btm.t330 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3300 VDD.t2791 a_22775_42718# a_22465_38541# VDD.t2790 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3301 a_18796_44728# a_17715_44356# a_18449_44324# VDD.t633 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3302 a_18404_46526# a_18190_46526# VDD.t1065 VDD.t1064 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X3303 VDD.t2777 a_2151_45670# a_1735_46195# VDD.t2776 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X3304 VDAC_N.t105 C10_N_btm.t614 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3305 VDAC_P.t1265 C8_P_btm.t152 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3306 VDAC_N.t1259 C10_N_btm.t613 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3307 C9_P_btm.t4 EN_VIN_BSTR_P.t16 VIN_P.t12 VSS.t558 sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X3308 VDAC_P.t337 C10_P_btm.t641 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3309 VDAC_N.t643 C9_N_btm.t329 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3310 VDAC_N.t1257 C9_N_btm.t328 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3311 a_4091_47070# a_4061_47044# VSS.t1578 VSS.t1577 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3312 VDAC_P.t1263 C9_P_btm.t305 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3313 C10_N_btm.t18 a_22812_30659.t4 VREF.t40 VDD.t516 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3314 a_15589_44350# a_12769_44594.t7 VDD.t55 VDD.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X3315 VDAC_N.t335 C8_N_btm.t147 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3316 VCM.t13 a_3990_30651.t14 C10_N_btm.t13 VSS.t286 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3317 VSS.t2551 VSS.t2552 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3318 a_215_46348# a_n409_45982# a_107_45982# VDD.t979 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3319 VDAC_P.t645 C5_P_btm.t11 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3320 VDAC_P.t1261 C6_P_btm.t33 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3321 VDD.t355 a_n690_43494.t10 a_1431_45982# VDD.t354 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3322 VSS.t2523 VSS.t2524 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3323 VDAC_P.t105 C10_P_btm.t640 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3324 VDAC_N.t1255 C5_N_btm.t17 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3325 VDAC_N.t641 C9_N_btm.t327 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3326 VDAC_N.t1253 C10_N_btm.t611 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3327 a_6673_45136# a_6455_44894# VDD.t872 VDD.t871 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3328 VDAC_N.t181 C7_N_btm.t38 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3329 VDAC_N.t1251 C8_N_btm.t146 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3330 VDAC_P.t1259 C8_P_btm.t151 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3331 VSS.t3457 VDD.t3211 VSS.t3456 VSS.t3455 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3332 VDAC_N.t639 C10_N_btm.t610 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3333 VDAC_N.t1249 C10_N_btm.t609 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3334 a_20647_31459.t1 a_22223_47070# VSS.t2695 VSS.t1136 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3335 VSS.t2401 VSS.t2402 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3336 VDAC_P.t643 C9_P_btm.t304 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3337 VDAC_N.t333 C10_N_btm.t608 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3338 VDAC_P.t1257 C9_P_btm.t303 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3339 VDAC_P.t335 C9_P_btm.t302 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3340 VDAC_P.t1255 C10_P_btm.t639 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3341 VDAC_P.t641 C8_P_btm.t150 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3342 VDAC_N.t1247 C9_N_btm.t326 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3343 VDAC_N.t637 C10_N_btm.t607 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3344 VDAC_P.t1253 C10_P_btm.t638 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3345 VDAC_N.t1245 C10_N_btm.t606 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3346 VDAC_N.t47 C10_N_btm.t605 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3347 a_8609_46232# a_6485_44582.t12 a_8514_46232# VDD.t3016 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X3348 VDAC_P.t181 C10_P_btm.t637 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3349 VDAC_N.t1243 C10_N_btm.t604 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3350 VDAC_N.t635 C7_N_btm.t81 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3351 VDD.t1678 a_16291_44914# a_16211_44582# VDD.t1677 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3352 VDAC_P.t1251 C10_P_btm.t636 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3353 VDAC_N.t1241 C6_N_btm.t65 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3354 VDAC_N.t331 C9_N_btm.t325 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3355 C10_N_btm.t14 a_3990_30651.t16 VCM.t15 VSS.t288 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3356 VDD.t73 a_n1551_45412.t12 a_n2293_44332# VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3357 VDAC_N.t1239 C7_N_btm.t80 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3358 VDD.t2642 VSS.t3561 VDD.t2641 VDD.t2640 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3359 VDAC_P.t639 C6_P_btm.t32 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3360 a_10537_46224# a_10319_45982# VDD.t1490 VDD.t1489 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3361 VSS.t1746 a_16475_45412# a_18845_42746# VSS.t1745 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3362 a_2864_43806# a_2627_42718# VSS.t1414 VSS.t1413 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3363 VSS.t3478 VDD.t3219 VSS.t3477 VSS.t3476 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3364 VDAC_P.t1249 C8_P_btm.t149 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3365 VREF.t11 a_n2467_30659.t4 C9_P_btm.t5 VDD.t577 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3366 a_14819_44582# a_15091_44440# VSS.t761 VSS.t760 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3367 a_2358_46565# a_885_44868.t17 VDD.t2838 VDD.t2837 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3368 VDD.t1540 a_11507_47833# a_11299_47832# VDD.t1539 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3369 VDAC_N.t633 C10_N_btm.t603 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3370 VSS.t1293 a_20283_43262# a_20383_42718# VSS.t1292 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3371 VSS.t590 a_13524_46832.t6 a_16291_46758# VSS.t589 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3372 VDAC_P.t333 C10_P_btm.t635 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3373 VSS.t1344 a_4987_45742# a_4921_45816# VSS.t1343 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3374 VSS.t1410 a_12427_46758# a_10684_45670# VSS.t1409 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X3375 VDAC_N.t1237 C4_N_btm.t4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3376 VDD.t48 a_8727_47222.t16 a_9343_43806# VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X3377 VDAC_N.t179 C8_N_btm.t145 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3378 VDAC_P.t1247 C10_P_btm.t634 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3379 VDAC_N.t1235 C9_N_btm.t324 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3380 VSS.t819 a_571_43566# a_505_43640# VSS.t818 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3381 a_n2833_47874# a_n2497_47846.t7 VDD.t2050 VDD.t2049 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X3382 VSS.t3592 C8_N_btm.t270 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3383 VSS.t2900 a_n2810_43806.t5 C6_P_btm.t70 VSS.t2899 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3384 VDAC_N.t631 C9_N_btm.t323 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3385 VDAC_N.t1233 C10_N_btm.t602 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3386 VSS.t1029 a_22223_47622# a_21788_30659.t1 VSS.t1028 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3387 a_10224_45982# a_9973_46526# VSS.t867 VSS.t866 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3388 VDAC_N.t329 C10_N_btm.t601 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3389 VDAC_P.t637 C10_P_btm.t633 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3390 VDAC_P.t1245 C9_P_btm.t297 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3391 a_1663_46565# a_1412_46794.t9 a_1204_46758# VDD.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3392 VDAC_N.t1231 C10_N_btm.t600 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3393 VSS.t1813 a_12896_47044# a_n2661_47044.t1 VSS.t1812 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X3394 a_22276_45412# a_22455_45420# VSS.t1322 VSS.t1321 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3395 VDAC_N.t629 C10_N_btm.t294 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3396 VDAC_P.t47 C9_P_btm.t296 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3397 a_n1827_44324.t0 a_5536_44324# VSS.t718 VSS.t717 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X3398 VDAC_P.t1243 C9_P_btm.t295 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3399 VDAC_P.t635 C10_P_btm.t632 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3400 VDAC_P.t1241 C10_P_btm.t310 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3401 VSS.t3670 C8_N_btm.t262 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3402 VSS.t1922 a_7754_38470# VSS.t1921 VSS.t1920 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X3403 a_8061_43262# a_6631_44582# VDD.t1443 VDD.t1442 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3404 VSS.t2032 a_4791_42883# a_3576_44364# VSS.t2031 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3405 VSS.t3041 VDD.t3115 VSS.t3040 VSS.t3039 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3406 VDAC_N.t1229 C6_N_btm.t42 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3407 VDAC_P.t331 C7_P_btm.t73 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3408 VDD.t357 a_n690_43494.t12 a_n409_45982# VDD.t356 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3409 VDAC_P.t1239 C9_P_btm.t294 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3410 VDAC_N.t103 C8_N_btm.t142 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3411 VDAC_N.t1227 C10_N_btm.t596 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3412 VDAC_P.t633 C5_P_btm.t23 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3413 VDD.t2900 a_1334_43494.t8 a_6491_44716# VDD.t2899 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X3414 VDAC_P.t1237 C10_P_btm.t628 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3415 a_15139_47730# a_13524_46832.t18 VSS.t606 VSS.t605 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3416 VDAC_P.t179 C7_P_btm.t72 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3417 a_n1085_47874# a_n749_47846# VSS.t952 VSS.t951 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X3418 a_6635_47044# a_4830_43958.t4 VDD.t196 VDD.t195 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X3419 VDAC_P.t1235 C8_P_btm.t148 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3420 a_5700_37509.t15 VDAC_N.t627 a_8912_37509.t21 VDD.t2252 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3421 a_18190_46526# a_18103_46768# a_17786_46658# VDD.t1796 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X3422 VDAC_P.t631 C10_P_btm.t627 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3423 a_14331_43806# a_14077_44133# VSS.t841 VSS.t840 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X3424 a_15329_47044# a_15879_47320# VSS.t1412 VSS.t1411 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258375 ps=1.445 w=0.65 l=0.15
X3425 VSS.t246 a_18314_32299.t4 C10_N_btm.t0 VSS.t245 sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X3426 VSS.t1071 a_12684_45276# a_12436_44868# VSS.t1070 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3427 VSS.t363 a_n1827_45412.t13 a_n2661_44332# VSS.t362 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3428 VDAC_N.t1225 C9_N_btm.t322 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3429 a_10185_47070# a_10150_47322# a_9947_47044# VSS.t755 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3430 VDAC_P.t1233 C10_P_btm.t626 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3431 VDAC_N.t327 C10_N_btm.t594 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3432 a_n73_46904# a_n519_46532# a_n169_46904# VSS.t1134 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3433 a_8416_45554# a_5419_47258# VDD.t1529 VDD.t1528 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X3434 a_9144_45144# a_9096_45276.t3 a_9060_45144# VDD.t532 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3435 VDAC_N.t1223 C9_N_btm.t321 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3436 VDAC_N.t625 C10_N_btm.t593 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3437 VDD.t2499 VSS.t3667 VDD.t2498 VDD.t2342 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3438 VDAC_N.t1221 C10_N_btm.t592 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3439 VDAC_N.t177 C10_N_btm.t591 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3440 VDAC_P.t329 C10_P_btm.t625 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3441 a_2113_38308# a_2113_38308# a_2113_38308# VSS.t2632 sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X3442 VDAC_P.t1231 C10_P_btm.t624 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3443 VDAC_P.t629 C10_P_btm.t623 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3444 VDAC_N.t1219 C10_N_btm.t590 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3445 a_3624_44466# a_3576_44364# a_3540_44466# VDD.t1088 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3446 VDD.t1255 a_2075_42718# a_2252_42718.t2 VDD.t1254 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3447 a_11671_44019# a_11183_44350# VSS.t1021 VSS.t1020 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3448 VDAC_P.t1229 C10_P_btm.t622 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3449 VDAC_N.t623 C7_N_btm.t79 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3450 VDAC_P.t103 C10_P_btm.t621 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3451 VDAC_N.t1217 C10_N_btm.t589 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3452 a_n1123_35174.t3 a_n1732_35090.t15 VSS.t2740 VSS.t2739 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3453 VSS.t3775 C7_P_btm.t5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3454 VDAC_N.t325 C5_N_btm.t32 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3455 VDAC_P.t1227 C8_P_btm.t147 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3456 VDAC_N.t1215 C10_N_btm.t588 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3457 a_10596_44324# a_10447_44403# VSS.t767 VSS.t766 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3458 VDD.t2139 a_n2472_43236# a_n2442_43262.t2 VDD.t2138 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3459 VDAC_N.t621 C8_N_btm.t141 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3460 VDD.t128 a_n1551_44324.t12 a_n2661_43780# VDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3461 VDAC_P.t627 C7_P_btm.t71 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3462 VDAC_P.t1225 C10_P_btm.t620 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3463 VDAC_P.t327 C9_P_btm.t293 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3464 VDAC_N.t1213 C9_N_btm.t320 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3465 VDAC_P.t1223 C10_P_btm.t619 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3466 VSS.t3772 C9_P_btm.t14 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3467 a_n2104_43236# a_n2073_43806# VSS.t829 VSS.t828 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3468 VDAC_N.t65 C9_N_btm.t319 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3469 a_n1459_43236.t4 a_570_44324# a_518_44670# VSS.t1652 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3470 VDAC_P.t625 C10_P_btm.t618 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3471 VDAC_N.t1211 C10_N_btm.t587 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3472 VDAC_N.t619 C10_N_btm.t586 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3473 VDAC_P.t1221 C9_P_btm.t291 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3474 VDAC_N.t1209 C10_N_btm.t585 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3475 C10_N_btm.t7 a_18314_32299.t11 VSS.t260 VSS.t259 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3476 VDD.t1073 a_18704_43806# a_18879_43780# VDD.t1072 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3477 a_4703_44894# a_4322_46134# a_885_44868.t7 VSS.t1820 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3478 VSS.t3053 VDD.t3119 VSS.t3052 VSS.t3051 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3479 VDD.t1950 a_n1085_47874# DATA[0].t4 VDD.t1949 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3480 VDAC_N.t323 C10_N_btm.t584 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3481 a_3895_46526# a_3271_46532# a_3787_46904# VDD.t1621 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3482 VDAC_P.t177 C10_P_btm.t617 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3483 VDAC_N.t1207 C10_N_btm.t583 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3484 VDAC_N.t617 C9_N_btm.t318 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3485 VSS.t2220 a_1431_47070# a_1203_42692.t2 VSS.t2219 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3486 VDAC_N.t1205 C10_N_btm.t582 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3487 VSS.t732 a_n2104_47044# a_n2074_47070.t0 VSS.t731 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3488 VDAC_P.t1219 C10_P_btm.t616 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3489 VSS.t637 a_10227_47214.t44 a_17821_46892# VSS.t636 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X3490 VSS.t1994 a_22591_43806# a_14409_32299.t1 VSS.t1993 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3491 VDAC_N.t175 C10_N_btm.t581 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3492 a_1429_47222.t1 a_15323_44894# VSS.t2122 VSS.t2121 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3493 VDAC_N.t1203 C10_N_btm.t580 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3494 VDAC_P.t623 C8_P_btm.t146 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3495 VDD.t829 a_9159_43262# a_9898_44350# VDD.t828 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X3496 VDAC_P.t1217 C9_P_btm.t290 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3497 VDD.t1909 a_16579_43566# a_16566_43262# VDD.t1908 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3498 EN_COMP.t3 a_n2288_42692# VDD.t700 VDD.t699 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3499 VSS.t966 a_8483_43780# a_6485_44582.t0 VSS.t965 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3500 VDAC_N.t615 C10_N_btm.t579 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3501 VDAC_P.t325 C9_P_btm.t289 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3502 C9_P_btm.t539 a_4758_30651.t11 VCM.t62 VSS.t2992 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3503 a_3699_43780# a_135_43540.t10 VDD.t2904 VDD.t2903 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3504 a_15321_46526# a_15163_45670.t4 VDD.t116 VDD.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3505 VDAC_P.t1215 C10_P_btm.t615 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3506 VDAC_P.t621 C10_P_btm.t614 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3507 VDD.t1602 a_5441_46500# a_5089_47044# VDD.t1601 sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.26 ps=2.52 w=1 l=0.15
X3508 VSS.t999 a_5715_45956# a_5663_45982# VSS.t998 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X3509 a_10384_47436# a_9947_47044# VDD.t1968 VDD.t1967 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3510 VDAC_P.t1213 C9_P_btm.t287 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3511 VSS.t2305 VSS.t2306 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3512 VDAC_P.t5 a_3222_30651.t16 VCM.t37 VSS.t667 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X3513 VDAC_P.t1211 C10_P_btm.t613 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3514 VDAC_N.t1201 C7_N_btm.t78 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3515 VDAC_P.t619 C10_P_btm.t612 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3516 VSS.t3069 VDD.t3125 VSS.t3068 VSS.t3067 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3517 a_19732_46642# a_7208_47044# VDD.t2708 VDD.t2707 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X3518 a_4758_30651.t2 a_16703_42718# VDD.t846 VDD.t845 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3519 VDAC_P.t1209 C10_P_btm.t611 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3520 VDAC_N.t321 C6_N_btm.t41 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3521 VDD.t795 a_2043_43958# a_n60_44618# VDD.t794 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X3522 VDAC_N.t1199 C4_N_btm.t12 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3523 VDAC_N.t613 C10_N_btm.t578 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3524 VDD.t1498 a_16211_43780# a_16198_44172# VDD.t1497 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3525 VDAC_P.t323 C9_P_btm.t286 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3526 VDAC_N.t1197 C10_N_btm.t577 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3527 a_135_43540.t6 a_8391_47044# VDD.t1143 VDD.t1142 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3528 VSS.t236 a_2587_44868.t8 a_4703_44894# VSS.t235 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3529 VDAC_P.t1207 VSS.t3339 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3530 VDAC_N.t101 C9_N_btm.t317 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3531 VSS.t2511 VSS.t2512 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3532 a_n331_42718.t1 a_n501_42718# VDD.t1962 VDD.t1961 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3533 VDD.t403 a_13248_45956.t15 a_15079_46134# VDD.t402 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3534 VDAC_N.t1195 C9_N_btm.t316 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3535 VDAC_P.t617 C10_P_btm.t610 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3536 VDAC_P.t1205 C8_P_btm.t145 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3537 VDAC_P.t175 C10_P_btm.t609 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3538 VDAC_N.t611 C10_N_btm.t576 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3539 VSS.t3162 VDD.t3156 VSS.t3161 VSS.t3160 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3540 a_5569_44048# a_5351_43806# VDD.t857 VDD.t856 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3541 VDAC_N.t1193 C9_N_btm.t315 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3542 VDAC_P.t1203 C8_P_btm.t144 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3543 VDD.t3041 COMP_N.t9 a_n501_42718# VDD.t3040 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3544 VDAC_P.t615 C10_P_btm.t608 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3545 VDAC_N.t319 C10_N_btm.t575 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3546 VDAC_P.t1201 C10_P_btm.t607 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3547 VDAC_N.t1191 C10_N_btm.t574 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3548 VDAC_P.t321 C10_P_btm.t606 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3549 EN_VIN_BSTR_P.t6 a_n1732_35090.t13 w_1375_34946.t17 w_1375_34946.t16 sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3550 VDAC_P.t1199 C10_P_btm.t605 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3551 VDD.t2537 VSS.t3654 VDD.t2536 VDD.t2535 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3552 a_15962_47320# a_15691_47436# a_15879_47320# VDD.t701 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3553 VSS.t304 a_n1827_44324.t8 a_n2293_43244# VSS.t303 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3554 a_283_42692# a_1203_42692.t16 a_1161_42968# VDD.t478 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3555 VSS.t3610 C10_N_btm.t1071 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3556 VDAC_N.t609 C10_N_btm.t572 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3557 VREF.t28 a_21788_30659.t9 C9_N_btm.t10 VDD.t2056 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3558 VDAC_N.t1189 C8_N_btm.t140 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3559 VDAC_N.t173 C10_N_btm.t571 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3560 a_15733_43806# a_15689_44048# a_15567_43806# VSS.t1488 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3561 VSS.t744 a_n2472_44868# a_n2442_44894.t0 VSS.t743 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3562 VDAC_P.t613 C10_P_btm.t604 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3563 VDAC_P.t1197 C10_P_btm.t603 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3564 VDAC_N.t0 a_3222_30651.t4 VCM.t31 VSS.t656 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3565 a_4239_42883# a_2252_42718.t6 VSS.t2980 VSS.t2979 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3566 VDAC_P.t101 C10_P_btm.t602 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3567 VDAC_N.t607 C10_N_btm.t570 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3568 VDAC_P.t1195 C4_P_btm.t12 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3569 VREF.t21 a_n1890_47614.t5 C7_P_btm.t2 VDD.t2039 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3570 a_5485_43262# a_4322_46134# VDD.t1784 VDD.t1783 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3571 a_18401_45982# a_18357_46224# a_18235_45982# VSS.t1495 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3572 VDAC_P.t611 C10_P_btm.t601 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3573 VDAC_P.t1193 C10_P_btm.t600 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3574 a_4791_42883# a_4000_42718.t4 VDD.t259 VDD.t258 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3575 VDD.t2546 VSS.t3651 VDD.t2545 VDD.t2544 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X3576 VDAC_N.t1185 C8_N_btm.t139 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3577 a_3726_37500# a_6886_37412# VSS.t1297 VSS.t1296 sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X3578 VDAC_P.t319 C10_P_btm.t599 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3579 a_14331_44133# a_n1067_42718.t5 a_14331_43806# VSS.t315 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3580 VSS.t1093 a_21197_42718# a_18766_43236# VSS.t1092 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3581 VDAC_P.t1191 C10_P_btm.t598 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3582 a_16579_47320# a_14766_45596.t8 a_15221_47044# VDD.t2881 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.265 ps=2.53 w=1 l=0.15
X3583 VDAC_N.t317 C7_N_btm.t77 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3584 VDAC_P.t609 C9_P_btm.t285 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3585 VDAC_N.t1183 C10_N_btm.t569 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3586 VSS.t799 a_22521_41035# a_22717_37721# VSS.t713 sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3587 VDAC_N.t605 C10_N_btm.t568 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3588 VDAC_N.t1181 C9_N_btm.t313 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3589 VDAC_P.t1189 C10_P_btm.t597 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3590 VDAC_N.t37 C9_N_btm.t312 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3591 a_n169_46904# a_n685_46532# a_n264_46892# VSS.t1640 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3592 VDD.t2184 a_4352_43640# a_4527_43566# VDD.t2183 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3593 VDAC_N.t1179 C9_N_btm.t311 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3594 VDD.t588 a_13273_44868.t16 a_14219_47070# VDD.t587 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3595 VDAC_P.t173 C10_P_btm.t596 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3596 a_n1890_47614.t0 a_n1920_47588# VSS.t2677 VSS.t2676 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3597 VDAC_P.t1187 C7_P_btm.t67 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3598 a_16618_44670# a_6104_45706.t9 a_16868_44670# VSS.t3010 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3599 VDD.t3098 a_6104_45706.t4 a_n2103_44868.t6 VDD.t3097 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3600 VSS.t3096 VDD.t3134 VSS.t3095 VSS.t3094 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X3601 a_1522_45554# a_1334_43494.t15 VDD.t337 VDD.t336 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X3602 VSS.t2942 SMPL.t11 a_18394_35068.t2 VSS.t2941 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3603 VDAC_N.t603 C9_N_btm.t310 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3604 VDAC_P.t607 C10_P_btm.t595 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3605 VDAC_N.t1177 C10_N_btm.t567 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3606 a_21755_44350# a_n2661_46508.t7 VDD.t2651 VDD.t2650 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3607 VDAC_N.t315 VSS.t3301 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3608 VDAC_P.t1185 VSS.t3346 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3609 VDAC_N.t1175 C8_N_btm.t138 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3610 VDAC_N.t601 C10_N_btm.t566 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3611 a_n2661_46508.t1 a_10596_44324# VDD.t1724 VDD.t1723 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3612 a_12461_44350# a_11455_44576.t20 a_12379_44350# VDD.t2823 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3613 VDAC_N.t1173 VSS.t3266 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3614 VREF.t71 a_19921_31459.t4 C2_N_btm.t8 VDD.t3070 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X3615 a_3067_44172# a_135_43540.t34 VDD.t184 VDD.t183 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3616 VDAC_N.t171 C10_N_btm.t565 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3617 VDAC_P.t317 C10_P_btm.t594 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3618 VDAC_P.t1183 C10_P_btm.t593 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3619 VSS.t398 a_1334_43494.t17 a_3089_42718# VSS.t397 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3620 VDAC_N.t1171 C10_N_btm.t564 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3621 VDAC_P.t605 C10_P_btm.t592 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3622 VCM.t49 a_5334_30651.t7 C7_N_btm.t138 VSS.t2936 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X3623 VDD.t1231 a_7961_46500# a_7851_46526# VDD.t1230 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3624 VDD.t2834 a_885_44868.t14 a_1297_45221# VDD.t2833 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X3625 a_647_47070# a_n53_44363.t17 a_284_47222# VSS.t623 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3626 VDAC_P.t1181 C9_P_btm.t284 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3627 VSS.t2468 VSS.t2469 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3628 VDAC_P.t37 C10_P_btm.t591 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3629 VSS.t1295 a_6886_37412# a_4338_37500.t5 VSS.t1294 sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X3630 a_14297_32299.t0 a_22959_43270# VSS.t1455 VSS.t1454 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3631 VSS.t2460 VSS.t2461 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3632 a_n1735_43236.t4 a_2134_44324# a_2082_44670# VSS.t1786 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3633 VDD.t1253 a_2075_42870# a_2075_42718# VDD.t479 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3634 VDAC_P.t1179 C10_P_btm.t590 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3635 VDD.t2405 VSS.t3736 VDD.t2404 VDD.t2403 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3636 VDAC_N.t599 C10_N_btm.t563 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3637 VDAC_N.t1169 C8_N_btm.t137 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3638 a_14757_47614# a_14587_47614# VSS.t1404 VSS.t1403 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3639 VDAC_N.t313 C10_N_btm.t562 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3640 VDAC_P.t603 C9_P_btm.t283 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3641 VDAC_N.t1167 C10_N_btm.t561 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3642 VDAC_P.t1177 C10_P_btm.t589 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3643 VDAC_N.t597 C8_N_btm.t136 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3644 VSS.t2452 VSS.t2453 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3645 VDAC_P.t315 C10_P_btm.t588 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3646 VSS.t1115 a_428_42724# a_n2293_45420.t0 VSS.t1114 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3647 a_7961_44048# a_7743_43806# VSS.t1013 VSS.t1012 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3648 VSS.t2056 a_1488_43236# a_n2661_45420.t1 VSS.t2055 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X3649 VDAC_N.t1165 C8_N_btm.t135 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3650 DATA[5].t5 a_7595_47614# VDD.t1166 VDD.t1165 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3651 VDAC_P.t1175 C9_P_btm.t282 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3652 VDAC_P.t601 C8_P_btm.t143 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3653 VDAC_N.t99 C10_N_btm.t560 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3654 VDD.t2408 VSS.t3647 VDD.t2407 VDD.t2406 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3655 VSS.t3428 VDD.t3200 VSS.t3427 VSS.t3426 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3656 VDAC_P.t1173 VSS.t3345 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3657 VDAC_N.t1163 C9_N_btm.t309 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3658 a_6629_45982# a_5655_43780# VSS.t2246 VSS.t2245 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X3659 a_6491_44716# a_6485_44582.t10 VDD.t3015 VDD.t3014 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X3660 VDAC_P.t171 C7_P_btm.t66 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3661 VSS.t3186 VDD.t3164 VSS.t3185 VSS.t3184 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X3662 a_13661_46298# a_4322_46134# VDD.t1789 VDD.t1788 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3663 a_15468_45412# a_13715_43780# VSS.t1263 VSS.t1262 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3664 a_8727_47222.t3 a_11143_47588# VDD.t1377 VDD.t1376 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3665 VDAC_N.t595 C7_N_btm.t75 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3666 a_14821_43600# a_10251_45454# VSS.t1362 VSS.t1361 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X3667 a_6455_44894# a_6105_44894# a_6360_44894# VDD.t1548 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3668 VDAC_P.t1171 C10_P_btm.t587 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3669 VDD.t1803 a_22400_42718# a_22521_41035# VDD.t1802 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3670 VSS.t129 a_n1551_44324.t8 a_22959_46534# VSS.t128 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3671 a_2082_44670# a_82_45670# a_2332_44670# VSS.t1689 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3672 a_11265_44350# a_10259_42870.t20 a_11183_44350# VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3673 VSS.t780 a_15443_44582# a_15415_44350# VSS.t779 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3674 VSS.t3438 VDD.t3204 VSS.t3437 VSS.t3436 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3675 VDAC_N.t1161 C10_N_btm.t559 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3676 VDD.t1812 a_18689_45412# a_17763_44868# VDD.t1811 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3677 VDAC_P.t599 VSS.t3363 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3678 C0_P_btm.t2 a_134_42718.t5 VCM.t44 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X3679 VDAC_N.t311 C9_N_btm.t308 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3680 a_11834_46309# a_11788_46134# VDD.t1584 VDD.t1583 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3681 VDAC_P.t1169 C9_P_btm.t281 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3682 VDD.t1787 a_4322_46134# a_4993_47044# VDD.t1786 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3683 VDAC_N.t1159 C10_N_btm.t558 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3684 VDAC_P.t313 C10_P_btm.t586 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3685 VDAC_P.t1167 C10_P_btm.t585 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3686 a_18813_43806# a_17623_43806# a_18704_43806# VSS.t1937 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3687 VDAC_P.t597 C8_P_btm.t142 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3688 VDAC_N.t593 C10_N_btm.t557 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3689 VDAC_N.t1157 C10_N_btm.t556 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3690 VDAC_P.t1165 C10_P_btm.t584 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3691 a_9096_44350# a_8659_44324# VDD.t1225 VDD.t1224 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3692 a_85_47070# a_n193_47098# VDD.t676 VDD.t675 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3693 VDAC_N.t169 C10_N_btm.t555 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3694 VDAC_N.t1155 C10_N_btm.t554 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3695 VDAC_P.t99 C10_P_btm.t583 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3696 VDAC_P.t1163 C9_P_btm.t280 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3697 a_14552_43806# a_14301_44035# a_14331_44133# VSS.t1379 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3698 VDD.t2237 a_6235_46124# a_6196_46250# VDD.t2236 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3699 VDAC_N.t591 C10_N_btm.t553 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3700 VDAC_P.t595 C8_P_btm.t141 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3701 C7_P_btm.t138 a_5334_30651.t6 VCM.t48 VSS.t2935 sky130_fd_pr__nfet_01v8_lvt ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X3702 VDAC_N.t1153 C10_N_btm.t552 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3703 VDAC_N.t309 C7_N_btm.t74 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3704 VDAC_N.t1151 C10_N_btm.t551 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3705 VDAC_P.t1161 C9_P_btm.t279 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3706 VDD.t1381 a_22959_43270# a_14297_32299.t3 VDD.t1380 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3707 a_5840_42718.t3 a_5663_42718# VDD.t842 VDD.t841 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3708 VDAC_N.t589 C10_N_btm.t550 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3709 a_22780_40517# EN_COMP.t7 a_22521_40491# VSS.t2693 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3710 VSS.t406 a_1334_43494.t23 a_2075_42870# VSS.t405 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3711 VDD.t713 a_1633_46824# a_1663_46565# VDD.t712 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3712 a_1011_45221# a_829_45221# VDD.t639 VDD.t638 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X3713 VDAC_P.t311 C10_P_btm.t582 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3714 VSS.t2896 a_15549_47044.t12 a_n2497_42870.t0 VSS.t2895 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3715 VDAC_N.t1149 C9_N_btm.t307 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3716 a_n2288_42692# a_n2109_42692.t4 VSS.t2985 VSS.t2984 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3717 VDAC_N.t63 C9_N_btm.t306 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3718 VDAC_P.t1159 C10_P_btm.t581 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3719 w_11534_34010.t17 a_11730_34132.t7 w_11534_34010.t16 w_11534_34010.t10 sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X3720 VDD.t2595 VSS.t3714 VDD.t2594 VDD.t2593 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X3721 a_14194_46348# a_13524_46832.t10 VSS.t601 VSS.t600 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3722 VSS.t2420 VSS.t2421 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3723 VDAC_N.t1147 C8_N_btm.t134 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3724 VDAC_P.t593 C5_P_btm.t22 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3725 VDD.t62 a_1343_38525.t12 a_1736_39043.t0 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3726 VDAC_P.t1157 C10_P_btm.t580 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3727 VSS.t2417 VSS.t2415 a_3726_37500# VSS.t2416 sky130_fd_pr__nfet_01v8_lvt ad=0.589 pd=4.42 as=0.3135 ps=2.23 w=1.9 l=0.15
X3728 a_n2810_45438.t0 a_n2840_45412# VSS.t2107 VSS.t1656 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3729 C10_P_btm.t1078 a_n2810_44894.t10 VSS.t3284 VSS.t3283 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3730 a_7735_42692# a_1203_42692.t28 a_8061_43262# VDD.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3731 VDD.t545 a_13524_46832.t9 a_13427_46756# VDD.t544 sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.1083 ps=1.36 w=0.42 l=0.15
X3732 VIN_P.t0 EN_VIN_BSTR_P.t10 C0_P_btm.t1 VSS.t552 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X3733 VREF.t55 a_n4515_30659.t6 C10_P_btm.t1058 VDD.t2992 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3734 a_4921_45816# a_3731_45444# a_4812_45816# VSS.t2153 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3735 a_17613_44894# a_17763_44868# VSS.t1856 VSS.t1855 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X3736 VDAC_N.t587 VSS.t3254 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3737 VDAC_P.t169 C9_P_btm.t278 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3738 VDAC_N.t1145 C10_N_btm.t549 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3739 VDAC_P.t1155 C10_P_btm.t577 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3740 VDAC_P.t591 C10_P_btm.t576 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3741 VDAC_N.t307 C10_N_btm.t548 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3742 VDAC_N.t1143 C9_N_btm.t305 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3743 VDAC_P.t1153 C10_P_btm.t575 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3744 VDAC_N.t585 C10_N_btm.t547 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3745 VSS.t2397 VSS.t2398 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3746 VDAC_N.t1141 C10_N_btm.t546 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3747 a_16513_42718# a_12651_44576.t20 VSS.t2871 VSS.t2870 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3748 VDAC_N.t167 C10_N_btm.t545 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3749 VSS.t2525 VSS.t2526 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3750 VDD.t1245 a_12623_43780# a_10259_42870.t6 VDD.t1244 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3751 VDAC_P.t309 C10_P_btm.t574 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3752 VDD.t894 a_n447_47044# a_n749_47846# VDD.t893 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3753 VDAC_N.t1139 C10_N_btm.t544 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3754 VDAC_N.t583 VSS.t3253 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3755 VDAC_N.t1137 C10_N_btm.t543 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3756 a_1123_43780# a_948_43806# a_1302_43806# VSS.t856 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3757 VDAC_N.t305 C9_N_btm.t150 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3758 VSS.t328 a_10227_47214.t8 a_10949_43628# VSS.t327 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3759 VDAC_N.t1135 C10_N_btm.t542 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3760 VDAC_N.t581 C8_N_btm.t261 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3761 VDAC_P.t1151 C10_P_btm.t573 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3762 a_5536_44324# a_5387_44403# VSS.t916 VSS.t915 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3763 VDAC_N.t1133 C10_N_btm.t541 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3764 a_n2103_43780.t3 a_1847_45528.t8 VDD.t174 VDD.t173 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3765 VDAC_N.t97 C10_N_btm.t540 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3766 VDAC_P.t589 C10_P_btm.t572 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3767 VDAC_P.t1149 C8_P_btm.t140 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3768 VSS.t215 a_4830_43958.t18 a_9343_45982# VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3769 VDAC_P.t63 C8_P_btm.t139 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3770 VDD.t2984 a_15549_47044.t3 a_15467_47320# VDD.t2983 sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X3771 VDAC_N.t1131 C7_N_btm.t73 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3772 a_10475_43433# a_9987_42968# VDD.t1639 VDD.t1638 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3773 VSS.t63 a_12769_44594.t8 a_17242_43806# VSS.t62 sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X3774 VDAC_P.t1147 C10_P_btm.t571 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3775 VCM.t42 a_3222_30651.t10 VDAC_P.t3 VSS.t662 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3776 VSS.t964 a_8483_43780# a_6485_44582.t2 VSS.t963 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3777 VSS.t798 a_22521_41035# a_22469_41061# VSS.t797 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3778 VDD.t2606 VSS.t3704 VDD.t2605 VDD.t2604 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3779 VDAC_N.t579 C9_N_btm.t304 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3780 a_22609_38426# a_22521_39947# CAL_P.t0 VDD.t2685 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3781 a_11692_46134# a_n53_44363.t11 a_11834_46309# VDD.t558 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3782 VDAC_P.t1145 C2_P_btm.t5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3783 a_20049_43262# a_19771_43600# VSS.t1968 VSS.t1967 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3784 a_15221_47730# a_14766_45596.t10 a_15139_47730# VDD.t2882 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X3785 VSS.t1626 a_1123_43780# a_1581_43806.t3 VSS.t1625 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3786 VDAC_P.t307 C6_P_btm.t30 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3787 a_18044_43806# a_17515_43806# VSS.t1283 VSS.t1282 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3788 VDD.t2439 VSS.t3633 VDD.t2438 VDD.t2437 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X3789 VDAC_N.t1129 C9_N_btm.t303 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3790 VDAC_N.t303 VSS.t3300 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3791 a_7020_44894# a_5939_44894# a_6673_45136# VDD.t1543 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3792 VDAC_P.t1143 C8_P_btm.t138 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3793 VDAC_P.t585 C8_P_btm.t137 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3794 a_948_43806# a_n133_43806# a_601_44048# VDD.t850 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3795 VSS.t578 a_15730_45670.t26 a_16651_46500# VSS.t577 sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X3796 VSS.t2754 a_885_44868.t24 a_2301_45758# VSS.t2753 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3797 VSS.t2631 a_22959_44894# a_19437_31459.t1 VSS.t1122 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3798 VDAC_N.t1127 C9_N_btm.t302 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3799 VDD.t2615 VSS.t3700 VDD.t2614 VDD.t2613 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3800 VSS.t394 a_1429_47222.t22 a_1663_45046# VSS.t393 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3801 VDAC_P.t1141 C10_P_btm.t570 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3802 VDAC_N.t577 C9_N_btm.t301 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3803 VSS.t3579 C7_N_btm.t134 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3804 VDAC_P.t167 C8_P_btm.t136 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3805 VDAC_N.t1125 C10_N_btm.t539 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3806 VDAC_N.t165 C9_N_btm.t300 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3807 a_16291_46758# a_16291_44914# VSS.t1731 VSS.t1730 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X3808 VDAC_P.t1139 C10_P_btm.t569 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3809 a_3221_43806# a_3177_44048# a_3055_43806# VSS.t1219 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3810 a_7839_46904# a_7393_46532# a_7743_46904# VSS.t1278 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3811 a_16576_44868# a_16427_44894# VSS.t2054 VSS.t2053 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3812 VDAC_N.t1123 C10_N_btm.t538 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3813 VDAC_P.t583 C10_P_btm.t568 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3814 VDAC_N.t575 C10_N_btm.t537 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3815 VDAC_P.t1137 C9_P_btm.t277 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3816 VDAC_N.t1121 C8_N_btm.t132 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3817 VDAC_N.t301 C9_N_btm.t299 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3818 VDAC_P.t305 C10_P_btm.t567 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3819 VDAC_P.t1135 C10_P_btm.t566 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3820 VSS.t3630 C9_N_btm.t534 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3821 a_14331_44133# a_14301_44035# a_14259_44133# VDD.t1307 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3822 VDAC_P.t581 C9_P_btm.t276 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3823 VDAC_P.t1133 C10_P_btm.t565 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3824 a_10861_47070# a_10227_47214.t36 VSS.t629 VSS.t628 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X3825 VDAC_P.t97 C6_P_btm.t67 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3826 VDD.t386 a_n237_45454.t5 a_n193_47098# VDD.t385 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3827 a_4812_45816# a_3731_45444# a_4465_45412# VDD.t2116 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3828 VSS.t1757 a_16576_44868# a_n2293_47044.t1 VSS.t1756 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X3829 VSS.t3132 VDD.t3146 VSS.t3131 VSS.t3130 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X3830 VDAC_N.t1119 VSS.t3264 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3831 VDD.t728 a_22521_41035# a_22705_38842# VDD.t642 sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3832 a_n2661_47044.t0 a_12896_47044# VSS.t1815 VSS.t1814 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X3833 VDAC_P.t1131 C10_P_btm.t564 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3834 VDAC_N.t573 C10_N_btm.t536 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3835 VDD.t1313 a_n2833_47874# CLK_DATA.t7 VDD.t1312 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3836 VDD.t2946 a_2424_46794.t9 a_10415_47846# VDD.t2945 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3837 VDAC_N.t1117 C6_N_btm.t40 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3838 VDAC_P.t579 VSS.t3362 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3839 VDAC_N.t45 C9_N_btm.t297 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3840 a_n2840_45412# a_n2661_45420.t4 VSS.t354 VSS.t353 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3841 VDAC_P.t1129 C10_P_btm.t563 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3842 VDAC_P.t303 C9_P_btm.t275 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3843 VDAC_N.t1115 C8_N_btm.t131 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3844 VDAC_N.t571 C10_N_btm.t535 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3845 VSS.t2547 VSS.t2548 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3846 VDAC_P.t1127 C5_P_btm.t21 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3847 VSS.t2242 a_5655_43780# a_8897_44716# VSS.t2241 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X3848 a_n2467_30659.t3 a_n2472_47044# VDD.t2747 VDD.t2746 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3849 VDAC_N.t1113 C9_N_btm.t296 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3850 VDAC_P.t577 C7_P_btm.t64 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3851 a_n2810_44350.t0 a_n2840_44324# VSS.t936 VSS.t935 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3852 VDAC_P.t1125 C8_P_btm.t135 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3853 VDAC_N.t299 C10_N_btm.t534 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3854 VDD.t2676 a_9349_46539# a_9293_46565# VDD.t2675 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X3855 a_5088_37509.t5 VDAC_P.t165 a_8912_37509.t23 VDD.t2250 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3856 VSS.t310 a_17930_32299.t5 C9_N_btm.t1 VSS.t309 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3857 VDAC_N.t1111 C9_N_btm.t295 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3858 VDAC_P.t1123 C9_P_btm.t274 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3859 VDAC_N.t569 C9_N_btm.t294 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3860 VDAC_P.t575 C10_P_btm.t562 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3861 VDAC_P.t1121 C10_P_btm.t561 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3862 VDAC_P.t301 C10_P_btm.t560 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3863 VSS.t112 a_15163_45670.t2 a_15139_47730# VSS.t111 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X3864 VDAC_N.t1109 C9_N_btm.t293 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3865 VDAC_P.t1119 C8_P_btm.t134 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3866 VDAC_P.t573 C10_P_btm.t559 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3867 VDD.t1818 a_18971_44654# a_15730_45670.t5 VDD.t1817 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3868 VDAC_N.t163 C10_N_btm.t533 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3869 VDD.t2152 a_22591_44894# a_17930_32299.t3 VDD.t2151 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3870 a_4005_43236# a_3787_43640# VDD.t721 VDD.t720 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3871 VDAC_N.t1107 C10_N_btm.t1057 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3872 a_10414_43780# a_10844_44364# VDD.t2664 VDD.t2663 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.17575 ps=1.395 w=0.42 l=0.15
X3873 a_21276_30659.t1 a_22959_47070# VSS.t1204 VSS.t1203 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3874 VDAC_P.t1117 C10_P_btm.t558 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3875 VDAC_P.t45 C10_P_btm.t557 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3876 VDD.t609 a_n1735_43236.t13 a_22959_45446# VDD.t538 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3877 VDD.t715 a_7020_44894# a_7195_44868# VDD.t714 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3878 VDAC_N.t567 C8_N_btm.t130 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3879 a_12436_44868# a_2424_46794.t4 VSS.t2851 VSS.t2850 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X3880 VDAC_N.t1105 C8_N_btm.t129 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3881 a_2687_45956# a_2512_45982# a_2866_45982# VSS.t2590 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3882 VDAC_N.t297 C10_N_btm.t531 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3883 a_18541_43582# a_18766_43236# VSS.t1406 VSS.t1405 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3884 VDAC_P.t1115 C10_P_btm.t556 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3885 VSS.t932 a_104_42692# a_134_42718.t0 VSS.t931 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3886 VDAC_P.t571 C10_P_btm.t555 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3887 a_9969_45982# a_9803_45982# VSS.t2579 VSS.t2578 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3888 VSS.t1366 a_10251_45454# a_10197_45776# VSS.t1365 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3889 VDAC_N.t1103 C7_N_btm.t71 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3890 VDAC_N.t565 C10_N_btm.t530 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3891 VDAC_P.t1113 C10_P_btm.t554 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3892 VDAC_N.t1101 C5_N_btm.t16 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3893 VDAC_N.t95 C9_N_btm.t292 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3894 VDAC_P.t299 C8_P_btm.t273 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3895 a_5351_43806# a_5001_43806# a_5256_43806# VDD.t1162 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3896 VDAC_N.t1099 C9_N_btm.t291 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3897 VDD.t2630 VSS.t3570 VDD.t2629 VDD.t2628 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3898 VSS.t3454 VDD.t3210 VSS.t3453 VSS.t3452 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3899 VDAC_N.t563 C8_N_btm.t128 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3900 VDAC_N.t1097 C10_N_btm.t529 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3901 VSS.t352 a_10227_47214.t32 a_18401_45982# VSS.t351 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3902 a_5473_43582# a_1203_42692.t8 a_5485_43262# VDD.t466 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3903 VDAC_N.t295 C10_N_btm.t528 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3904 VDAC_P.t1111 C6_P_btm.t66 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3905 a_12151_46309# a_7208_47044# a_11692_46134# VDD.t2711 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3906 VDAC_P.t569 C10_P_btm.t553 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3907 a_3787_43640# a_3271_43268# a_3692_43628# VSS.t2111 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3908 VDAC_P.t1109 C8_P_btm.t133 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3909 VSS.t869 a_1204_46758# a_n447_47044# VSS.t868 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3910 VDAC_P.t163 C10_P_btm.t552 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3911 VSS.t3669 C9_P_btm.t20 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3912 VDAC_N.t1095 C10_N_btm.t527 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3913 a_7311_47614# a_6951_47070# VSS.t1612 VSS.t1611 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3914 VDAC_P.t1107 C9_P_btm.t273 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3915 VDAC_P.t567 VSS.t3360 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3916 a_18339_44350# a_10227_47214.t30 VDD.t303 VDD.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3917 a_18133_47235# a_4830_43958.t5 VSS.t202 VSS.t201 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3918 VDAC_P.t1105 C9_P_btm.t272 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3919 C9_N_btm.t2 a_17930_32299.t6 VSS.t312 VSS.t311 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3920 VDAC_N.t561 C10_N_btm.t526 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3921 a_13192_47320# a_13144_47452.t4 a_13108_47320# VDD.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3922 VDAC_P.t297 C9_P_btm.t271 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3923 VDAC_N.t1093 C8_N_btm.t127 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3924 VDAC_P.t1103 C9_P_btm.t270 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3925 a_16426_46642# a_16291_44914# VDD.t1674 VDD.t1673 sky130_fd_pr__pfet_01v8_hvt ad=0.05985 pd=0.705 as=0.14825 ps=1.34 w=0.42 l=0.15
X3926 VDAC_N.t161 C9_N_btm.t287 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3927 VDAC_N.t1091 C9_N_btm.t286 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3928 VDAC_N.t559 C10_N_btm.t525 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3929 VDAC_P.t565 C10_P_btm.t551 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3930 VDAC_N.t1089 C10_N_btm.t524 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3931 VDAC_N.t293 C10_N_btm.t523 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3932 a_22733_47833# DEBUG_MUX[3].t0 VDD.t3082 VDD.t3081 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3933 VDAC_P.t1101 C10_P_btm.t550 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3934 VDAC_P.t0 a_3222_30651.t6 VCM.t38 VSS.t658 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3935 VDAC_N.t1087 C9_N_btm.t285 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3936 VDAC_P.t1099 C9_P_btm.t269 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3937 C9_P_btm.t3 a_n2442_44894.t7 VSS.t373 VSS.t372 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3938 a_18879_43780# a_8727_47222.t10 VDD.t79 VDD.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3939 VDAC_N.t557 C10_N_btm.t522 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3940 VSS.t3575 C7_P_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3941 VDAC_P.t563 C9_P_btm.t266 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3942 VDAC_P.t1097 C10_P_btm.t549 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3943 VDAC_N.t1085 C8_N_btm.t126 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3944 VDAC_P.t295 C4_P_btm.t21 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3945 a_14409_32299.t0 a_22591_43806# VSS.t1992 VSS.t1991 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3946 a_6767_44716# a_1847_45528.t10 a_6661_44716# VSS.t166 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X3947 VDAC_P.t1095 C10_P_btm.t548 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3948 VDAC_P.t561 C10_P_btm.t547 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3949 a_16566_43262# a_15489_43268# a_16404_43640# VDD.t1644 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3950 VSS.t1055 a_9863_47874# DEBUG_OUT.t3 VSS.t1054 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3951 VDAC_P.t1093 C10_P_btm.t546 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3952 VDAC_N.t61 C6_N_btm.t39 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3953 VDAC_N.t1083 C9_N_btm.t284 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3954 VDAC_N.t555 C2_N_btm.t2 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3955 VDAC_P.t161 C9_P_btm.t265 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3956 VDAC_N.t29 C10_N_btm.t521 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3957 VDAC_N.t27 C9_N_btm.t283 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3958 VSS.t3102 VDD.t3136 VSS.t3101 VSS.t3100 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3959 VSS.t3012 a_n2103_44324.t4 a_22959_45982# VSS.t674 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3960 VDAC_N.t25 C9_N_btm.t282 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3961 VSS.t2474 VSS.t2475 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3962 a_135_43540.t7 a_8391_47044# VDD.t1149 VDD.t1148 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X3963 VDAC_N.t23 C8_N_btm.t260 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3964 VDAC_P.t1091 C10_P_btm.t545 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3965 VDAC_P.t559 C7_P_btm.t135 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3966 a_15121_43806# a_14955_43806# VSS.t1930 VSS.t1929 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3967 a_15831_42883# a_5142_30651.t7 VSS.t124 VSS.t123 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3968 VDAC_N.t21 C9_N_btm.t281 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3969 a_5542_30651.t2 a_11183_42718# VDD.t656 VDD.t655 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3970 VDAC_P.t1089 C9_P_btm.t264 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3971 VDAC_N.t19 C10_N_btm.t1056 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3972 EN_VIN_BSTR_P.t1 VDD.t3216 a_n283_35174# VSS.t3469 sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.9
X3973 VDAC_N.t17 C10_N_btm.t1054 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3974 a_16198_44172# a_15121_43806# a_16036_43806# VDD.t862 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3975 VDAC_P.t293 C10_P_btm.t544 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3976 a_15079_46134# a_13248_45956.t19 VDD.t407 VDD.t406 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3977 a_5088_37509.t15 VDAC_P.t1087 a_8912_37509.t33 VDD.t2242 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3978 a_4987_45742# a_4812_45816# a_5166_45804# VSS.t1340 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3979 VDAC_P.t557 C9_P_btm.t263 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3980 VDD.t741 a_4465_45412# a_4355_45438# VDD.t740 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3981 a_8850_45412# a_9096_45276.t4 VDD.t534 VDD.t533 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.17575 ps=1.395 w=0.42 l=0.15
X3982 C10_N_btm.t8 a_3990_30651.t4 VCM.t4 VSS.t277 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3983 a_19320_35138# VDD.t3174 EN_VIN_BSTR_N.t5 VSS.t3213 sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.9
X3984 VDD.t2090 a_n2840_47044# a_n2810_47070.t3 VDD.t2089 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3985 VDD.t1178 a_13635_43566# a_13622_43262# VDD.t1177 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3986 a_8912_37509.t35 VDAC_P.t1085 a_5088_37509.t17 VDD.t2243 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3987 a_1488_43236# a_82_45670# VSS.t1688 VSS.t1687 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X3988 VDAC_N.t15 VSS.t3287 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3989 VDAC_P.t61 VSS.t3371 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3990 a_18704_43806# a_17789_43806# a_18357_44048# VSS.t1132 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3991 VDAC_P.t1083 C10_P_btm.t543 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3992 VDAC_P.t555 C9_P_btm.t536 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3993 VDAC_N.t13 C8_N_btm.t125 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3994 VDD.t439 a_7754_40130.t5 a_8912_37509.t1 VDD.t438 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3995 a_215_46348# a_135_43540.t8 VDD.t2902 VDD.t2901 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3996 VDAC_P.t29 C6_P_btm.t64 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3997 VDAC_P.t27 C10_P_btm.t542 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3998 VDAC_P.t25 C6_P_btm.t28 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X3999 VDAC_P.t23 C10_P_btm.t541 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4000 VSS.t3657 C9_P_btm.t18 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4001 VDAC_P.t21 C10_P_btm.t540 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4002 VDAC_P.t19 C10_P_btm.t539 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4003 a_14955_45982# a_n1067_42718.t6 a_15133_45982# VSS.t316 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X4004 VDAC_N.t11 C6_N_btm.t38 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4005 VDAC_N.t10 C9_N_btm.t280 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4006 VSS.t1717 a_6091_43780# a_6025_43806# VSS.t1716 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4007 VDAC_P.t17 C8_P_btm.t272 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4008 VSS.t3003 a_14087_32299.t4 C3_N_btm.t12 VSS.t2880 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4009 a_2973_43582# a_1334_43494.t10 a_2627_43262# VSS.t374 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4010 VDAC_N.t1070 C8_N_btm.t124 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4011 VDAC_N.t2110 C10_N_btm.t1050 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4012 VDAC_N.t158 C9_N_btm.t279 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4013 a_n2833_42692# a_n2497_42870.t9 VDD.t2978 VDD.t2977 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X4014 VDD.t2552 VSS.t3754 VDD.t2551 VDD.t2550 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4015 VDAC_P.t15 C8_P_btm.t270 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4016 VDAC_P.t13 C10_P_btm.t538 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4017 a_14658_46526# a_13248_45956.t26 a_13930_46842# VSS.t492 sky130_fd_pr__nfet_01v8 ad=0.151025 pd=1.285 as=0.1092 ps=1.36 w=0.42 l=0.15
X4018 VDAC_P.t11 C10_P_btm.t537 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4019 a_7981_45956# a_7648_46134# VDD.t1492 VDD.t1491 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4020 a_4812_45816# a_3897_45444# a_4465_45412# VSS.t2159 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4021 VSS.t3587 C8_P_btm.t14 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4022 VDAC_N.t8 C9_N_btm.t278 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4023 VDAC_P.t10 C9_P_btm.t535 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4024 VDAC_P.t1070 C9_P_btm.t534 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4025 VDAC_P.t2110 C10_P_btm.t536 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4026 a_4527_43566# a_135_43540.t28 VDD.t176 VDD.t175 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4027 VDAC_N.t1066 C10_N_btm.t1048 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4028 VSS.t3505 VDD.t3228 VSS.t3504 VSS.t3503 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X4029 VSS.t2385 VSS.t2386 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4030 VDAC_N.t2102 C8_N_btm.t256 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4031 a_1513_47320# a_1429_47222.t8 a_1431_47070# VDD.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4032 a_16868_44670# a_6104_45706.t2 a_16618_44670# VSS.t3006 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4033 VSS.t3511 VDD.t3230 VSS.t3510 VSS.t3509 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4034 VDD.t1174 a_n2288_47588# a_n4515_30659.t2 VDD.t1173 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4035 a_6104_45706.t0 a_16211_43780# VSS.t1563 VSS.t1562 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X4036 VDAC_N.t546 C9_N_btm.t277 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4037 VDAC_N.t2098 C10_N_btm.t1046 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4038 a_18394_35068.t1 SMPL.t10 VSS.t2940 VSS.t2939 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4039 VDD.t1184 a_13635_43566# a_11455_44576.t7 VDD.t1183 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X4040 VSS.t2062 a_12887_47833# a_9551_47203# VSS.t2061 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4041 VDAC_P.t158 C10_P_btm.t535 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4042 VDAC_N.t1062 C8_N_btm.t123 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4043 VDAC_P.t8 C8_P_btm.t266 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4044 VDAC_N.t2094 C8_N_btm.t122 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4045 VDAC_P.t1066 C5_P_btm.t20 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4046 VDAC_P.t2102 C7_P_btm.t134 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4047 VDAC_P.t546 C7_P_btm.t61 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4048 a_12887_47833# CLK.t1 VSS.t2961 VSS.t2960 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4049 a_5441_46500# a_1429_47222.t7 a_5728_46526# VDD.t320 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X4050 VDAC_P.t2098 C10_P_btm.t534 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4051 VDD.t641 a_15437_47044# a_15691_47436# VDD.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4052 VDAC_P.t1062 C10_P_btm.t533 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4053 VDD.t1195 a_16211_44582# a_13715_43780# VDD.t1194 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X4054 VDAC_N.t286 C9_N_btm.t276 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4055 VDAC_N.t2090 C10_N_btm.t1044 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4056 VSS.t3150 VDD.t3152 VSS.t3149 VSS.t3148 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4057 a_11206_38545.t0 CAL_N.t3 a_4338_37500.t0 VDD.t145 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X4058 VDAC_N.t1058 C7_N_btm.t70 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4059 VDD.t57 a_12769_44594.t9 a_20107_43806# VDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4060 VDAC_N.t2086 C10_N_btm.t1042 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4061 VDAC_P.t2094 C9_P_btm.t532 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4062 VDAC_P.t286 C10_P_btm.t532 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4063 VSS.t2339 VSS.t2340 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4064 VDAC_P.t2090 C10_P_btm.t1055 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4065 a_15121_43806# a_14955_43806# VDD.t1879 VDD.t691 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4066 a_6360_44894# a_6243_45107# VSS.t2024 VSS.t2023 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4067 VDAC_P.t1058 C9_P_btm.t530 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4068 VSS.t3522 VDD.t3234 VSS.t3521 VSS.t3520 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4069 VDAC_P.t2086 C9_P_btm.t528 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4070 a_n2103_44868.t3 a_16670_44324# VDD.t1201 VDD.t1200 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4071 DATA[5].t4 a_7595_47614# VDD.t1170 VDD.t1169 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X4072 a_4279_46232# a_2755_43494.t18 VDD.t428 VDD.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4073 VDAC_P.t542 C10_P_btm.t530 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4074 VDAC_P.t2082 C10_P_btm.t529 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4075 VIN_N.t13 EN_VIN_BSTR_N.t18 C1_N_btm.t0 VSS.t444 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X4076 VDAC_N.t542 C10_N_btm.t1040 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4077 VDAC_N.t2082 C9_N_btm.t275 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4078 VDAC_N.t1054 C10_N_btm.t1038 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4079 VDAC_P.t1054 C10_P_btm.t528 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4080 VDD.t1831 a_13991_42883# a_12684_45276# VDD.t1830 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4081 VSS.t1400 a_8483_46830# a_8417_46904# VSS.t1399 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4082 a_n2293_45420.t1 a_428_42724# VSS.t1117 VSS.t1116 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X4083 a_1083_44894# a_829_45221# VSS.t709 VSS.t708 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X4084 a_468_42870# a_927_42692.t8 VDD.t91 VDD.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X4085 a_n2661_45420.t0 a_1488_43236# VSS.t2058 VSS.t2057 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4086 VDD.t1164 a_5916_43806# a_6091_43780# VDD.t1163 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4087 VDAC_N.t2078 C7_N_btm.t69 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4088 a_5088_37509.t19 VDAC_P.t2078 a_8912_37509.t37 VDD.t2248 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4089 VDAC_P.t30 C10_P_btm.t527 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4090 VDAC_N.t30 C6_N_btm.t37 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4091 a_10259_42870.t2 a_12623_43780# VSS.t1306 VSS.t1305 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4092 VDAC_N.t2074 C5_N_btm.t30 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4093 VDAC_N.t1050 C8_N_btm.t252 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4094 VDAC_P.t2074 C8_P_btm.t265 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4095 VDAC_N.t2070 C10_N_btm.t509 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4096 a_4279_46232# a_n2497_47846.t3 a_4061_45956# VDD.t2046 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X4097 VSS.t3540 VDD.t3240 VSS.t3539 VSS.t3538 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4098 VDD.t93 a_927_42692.t9 a_n1459_43236.t0 VDD.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.135 ps=1.27 w=1 l=0.15
X4099 a_8912_37509.t36 VDAC_P.t1050 a_5088_37509.t18 VDD.t2255 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4100 VDAC_N.t538 C9_N_btm.t274 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4101 VDAC_P.t2070 C8_P_btm.t127 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4102 VDAC_P.t538 C10_P_btm.t526 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4103 C10_N_btm.t4 a_18314_32299.t8 VSS.t254 VSS.t253 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4104 a_19037_42718# a_18759_42746# VSS.t1751 VSS.t1750 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X4105 VSS.t1663 a_5089_47044# a_4704_47044# VSS.t1662 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X4106 VDAC_N.t2066 C10_N_btm.t507 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4107 VDAC_P.t2066 C10_P_btm.t525 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4108 a_17763_44868# a_18689_45412# VDD.t1808 VDD.t1807 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4109 VDAC_P.t1046 C10_P_btm.t524 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4110 VDAC_N.t1046 C10_N_btm.t506 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4111 VDAC_P.t2062 C10_P_btm.t523 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4112 a_594_42968# a_546_43100# a_510_42968# VDD.t1764 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4113 VDAC_N.t2062 C8_N_btm.t251 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4114 VDAC_N.t282 C9_N_btm.t273 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4115 VDAC_N.t2058 C10_N_btm.t505 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4116 a_n243_45982# a_n409_45982# VSS.t1039 VSS.t1038 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4117 VSS.t3156 VDD.t3154 VSS.t3155 VSS.t3154 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4118 a_13930_46842# a_13524_46832.t8 a_13848_46842# VSS.t599 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4119 a_468_42870# a_927_42692.t12 VSS.t90 VSS.t89 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4120 C10_P_btm.t2 a_3990_30651.t10 VCM.t10 VSS.t283 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4121 VDAC_N.t1042 C10_N_btm.t504 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4122 VDAC_N.t2054 C8_N_btm.t250 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4123 VDD.t508 a_1053_45123.t3 a_n1551_44324.t7 VDD.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4124 a_20283_43262# a_1203_42692.t18 VDD.t481 VDD.t480 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4125 VDAC_P.t282 C10_P_btm.t521 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4126 a_11971_46500# a_12127_46744# VSS.t1109 VSS.t85 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X4127 VDAC_N.t534 C10_N_btm.t503 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4128 VDAC_P.t2058 C9_P_btm.t526 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4129 VSS.t1130 a_571_46830# a_505_46904# VSS.t1129 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4130 VSS.t380 a_1429_47222.t6 a_n2109_42692.t2 VSS.t379 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4131 VDAC_N.t2050 C9_N_btm.t272 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4132 VDAC_P.t1042 C9_P_btm.t255 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4133 VDAC_P.t2054 C9_P_btm.t522 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4134 a_13113_43236# a_12895_43640# VSS.t1567 VSS.t1566 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4135 VSS.t455 a_n331_42718.t3 a_15393_45982# VSS.t454 sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X4136 a_n2472_45412# a_n2293_45420.t7 VSS.t2785 VSS.t2784 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4137 VSS.t178 a_135_43540.t36 a_3221_43806# VSS.t177 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4138 VSS.t641 a_13273_44868.t15 a_n2497_42870.t6 VSS.t640 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4139 a_10933_47070# a_10554_47436# a_10861_47070# VSS.t1176 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X4140 VDAC_P.t534 C10_P_btm.t520 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4141 a_18348_43262# a_15549_47044.t9 a_18093_43262# VDD.t2986 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4142 a_2075_42870# a_1203_42692.t22 VSS.t534 VSS.t533 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4143 a_7851_46526# a_7227_46532# a_7743_46904# VDD.t1211 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4144 VSS.t2513 VSS.t2514 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4145 VDD.t147 CAL_N.t4 VDD.t147 VDD.t146 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X4146 VDAC_N.t1038 C6_N_btm.t36 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4147 VDAC_P.t2050 C8_P_btm.t126 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4148 a_15155_47320# a_15113_47222# VDD.t1666 VDD.t1665 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4149 VDAC_N.t2046 C6_N_btm.t35 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4150 VDAC_N.t154 C10_N_btm.t502 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4151 VDAC_P.t1038 C10_P_btm.t519 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4152 a_n291_45776# a_n1067_42718.t7 a_n377_45776# VSS.t317 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4153 VDAC_N.t2042 C8_N_btm.t249 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4154 VDAC_P.t2046 C8_P_btm.t262 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4155 VDAC_N.t1034 C10_N_btm.t1030 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4156 VDAC_P.t154 C5_P_btm.t19 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4157 a_663_47874# a_999_47846# VSS.t2010 VSS.t2009 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X4158 VDAC_P.t2042 C10_P_btm.t1054 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4159 VDAC_P.t1034 C8_P_btm.t125 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4160 a_15582_45982# a_14955_45982# VSS.t1665 VSS.t1664 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X4161 VDAC_N.t2038 C10_N_btm.t1027 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4162 VSS.t3546 VDD.t3242 VSS.t3545 VSS.t3544 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4163 a_n2661_45956.t2 a_6126_46642# VDD.t1248 VDD.t1247 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X4164 VDAC_P.t2038 C7_P_btm.t130 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4165 VDD.t2684 a_2512_45982# a_2687_45956# VDD.t2683 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4166 a_n1735_43236.t0 a_1334_43494.t11 VDD.t332 VDD.t331 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4167 VDAC_N.t530 C10_N_btm.t1012 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4168 C10_N_btm.t10 a_3990_30651.t6 VCM.t6 VSS.t279 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4169 VDAC_N.t2034 C9_N_btm.t271 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4170 VDD.t384 a_n2109_47596.t9 a_22455_45420# VDD.t383 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4171 VDAC_N.t1030 C9_N_btm.t270 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4172 VSS.t2399 VSS.t2400 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4173 VDAC_N.t2030 C10_N_btm.t991 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4174 VDAC_N.t278 C10_N_btm.t974 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4175 VDAC_P.t530 C10_P_btm.t1052 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4176 VDAC_N.t2026 VSS.t3314 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4177 a_3800_45982# a_3165_45982# a_3320_46134# VSS.t1465 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4178 a_4509_45804# a_4465_45412# a_4343_45816# VSS.t811 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X4179 VDD.t343 a_1334_43494.t20 a_1659_44440# VDD.t342 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4180 a_13273_44868.t3 a_18879_43780# VSS.t1636 VSS.t1635 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4181 VDD.t1391 a_3165_45982# a_n2103_43780.t0 VDD.t1390 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4182 a_1203_42692.t3 a_1431_47070# VSS.t2222 VSS.t2221 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4183 a_4527_43566# a_4352_43640# a_4706_43628# VSS.t2216 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X4184 VDAC_P.t2034 C10_P_btm.t1050 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4185 VDAC_N.t1026 C10_N_btm.t905 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4186 VDAC_P.t1030 VSS.t3351 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4187 VDAC_P.t2030 C7_P_btm.t60 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4188 VDAC_N.t2022 C4_N_btm.t19 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4189 a_3470_45982# a_1847_45528.t9 VSS.t165 VSS.t164 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X4190 VDD.t52 a_12769_44594.t5 a_12461_44350# VDD.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4191 VDAC_N.t526 C8_N_btm.t248 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4192 VDAC_P.t278 C8_P_btm.t260 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4193 C2_N_btm.t1 EN_VIN_BSTR_N.t10 VIN_N.t10 VSS.t439 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X4194 a_6485_44582.t3 a_8483_43780# VSS.t960 VSS.t959 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4195 VSS.t681 a_13273_44868.t8 a_19168_45758# VSS.t680 sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.08775 ps=0.92 w=0.65 l=0.15
X4196 VDAC_P.t2026 C8_P_btm.t124 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4197 VDAC_N.t2018 C10_N_btm.t892 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4198 VDAC_P.t1026 C10_P_btm.t1048 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4199 a_1581_43806.t0 a_1123_43780# VSS.t1620 VSS.t1619 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4200 VDAC_P.t2022 C10_P_btm.t1046 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4201 VSS.t420 a_n690_43494.t16 a_n133_43806# VSS.t419 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4202 a_2252_42718.t0 a_2075_42718# VSS.t1326 VSS.t1325 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4203 VDAC_N.t1022 C10_N_btm.t772 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4204 a_6707_45776# a_5663_45982# VDD.t2692 VDD.t2691 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4205 VDAC_P.t526 C9_P_btm.t520 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4206 VDAC_P.t2018 C9_P_btm.t252 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4207 VDAC_N.t2014 C9_N_btm.t269 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4208 a_2112_39137# a_1343_38525.t11 VDD.t60 VDD.t58 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4209 a_n1827_44868.t0 a_1412_46794.t4 VDD.t159 VDD.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4210 VDAC_P.t1022 C10_P_btm.t1044 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4211 VDAC_P.t2014 C9_P_btm.t251 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4212 a_8912_37509.t26 VDAC_P.t90 a_5088_37509.t8 VDD.t2246 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4213 a_18445_42718# a_13273_44868.t26 VSS.t650 VSS.t649 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4214 a_n169_46904# a_n519_46532# a_n264_46892# VDD.t1075 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4215 VDD.t489 a_15730_45670.t8 a_14635_44324# VDD.t488 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X4216 VDAC_P.t2010 C10_P_btm.t515 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4217 VDAC_N.t90 C9_N_btm.t268 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4218 VDAC_N.t2010 C10_N_btm.t757 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4219 a_10892_44466# a_10844_44364# a_10808_44466# VDD.t2662 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4220 a_16921_46364# a_13248_45956.t9 VDD.t397 VDD.t396 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4221 VSS.t2713 a_11455_44576.t12 a_11687_45528# VSS.t2712 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4222 a_1663_45046# a_1581_43806.t14 VSS.t2906 VSS.t2905 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X4223 VDAC_N.t1018 C10_N_btm.t619 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4224 VSS.t1632 a_18879_43780# a_13273_44868.t1 VSS.t1631 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X4225 a_17881_44356# a_17715_44356# VDD.t631 VDD.t630 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4226 a_n268_44582# a_n60_44618# a_n126_44716# VSS.t827 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4227 VDAC_P.t1018 C10_P_btm.t1040 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4228 VSS.t3746 C9_N_btm.t525 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4229 VSS.t2950 SMPL.t18 a_n1732_35090.t4 VSS.t2949 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4230 a_13569_43640# a_12379_43268# a_13460_43640# VSS.t1156 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4231 VDAC_N.t2006 C9_N_btm.t266 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4232 a_7000_47222# a_7208_47044# a_7142_47070# VSS.t2610 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4233 VDAC_P.t2006 C8_P_btm.t258 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4234 VDAC_P.t522 C9_P_btm.t250 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4235 VDAC_P.t2002 C10_P_btm.t1038 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4236 VDD.t1315 a_n2833_47874# CLK_DATA.t6 VDD.t1314 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X4237 VDD.t1607 a_15582_45982# a_15962_47320# VDD.t1606 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X4238 VDAC_P.t1014 C10_P_btm.t1036 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4239 VDAC_P.t1998 C9_P_btm.t249 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4240 C5_P_btm.t37 a_n2442_43806.t4 VSS.t2981 VSS.t457 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X4241 a_n2293_47044.t0 a_16576_44868# VSS.t1755 VSS.t1754 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4242 VDAC_P.t274 C9_P_btm.t248 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4243 VDAC_N.t522 C10_N_btm.t612 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4244 VDD.t3105 a_n2103_44324.t7 a_22959_45982# VDD.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4245 VSS.t3712 C7_N_btm.t136 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4246 a_15691_47614# a_15163_45670.t3 VSS.t114 VSS.t113 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4247 VDD.t3018 a_6485_44582.t18 a_n1827_44868.t6 VDD.t3017 sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.135 ps=1.27 w=1 l=0.15
X4248 VSS.t2454 VSS.t2455 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4249 VDAC_P.t1994 C7_P_btm.t128 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4250 VDAC_P.t1010 C10_P_btm.t508 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4251 VDAC_N.t2002 C6_N_btm.t34 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4252 a_10415_47846# a_n237_45454.t20 VDD.t422 VDD.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X4253 VDAC_N.t1014 C10_N_btm.t597 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4254 VDAC_N.t1998 C10_N_btm.t595 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4255 a_7020_44894# a_6105_44894# a_6673_45136# VSS.t1609 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4256 VDAC_N.t274 C8_N_btm.t247 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4257 VDAC_P.t1990 VSS.t3378 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4258 VSS.t3231 VDD.t3180 VSS.t3230 VSS.t3229 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4259 VDD.t1566 a_10623_47307# a_10554_47436# VDD.t1565 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X4260 a_12931_45982# a_13248_45956.t7 a_13181_45982# VSS.t477 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.085225 ps=0.925 w=0.42 l=0.15
X4261 VDAC_P.t518 C8_P_btm.t121 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4262 VDAC_N.t1994 C9_N_btm.t265 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4263 VDAC_N.t1010 C10_N_btm.t519 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4264 VDD.t239 a_2587_44868.t18 a_11265_44350# VDD.t238 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4265 VDAC_P.t1986 C10_P_btm.t507 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4266 VDAC_P.t1006 C10_P_btm.t506 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4267 VDAC_P.t1982 C9_P_btm.t247 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4268 VDAC_N.t1990 C10_N_btm.t518 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4269 VDAC_P.t150 C10_P_btm.t505 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4270 VDAC_N.t518 C7_N_btm.t68 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4271 VDD.t2745 a_n2472_47044# a_n2467_30659.t2 VDD.t2744 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4272 VDAC_P.t1978 C9_P_btm.t512 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4273 VDAC_N.t1986 C10_N_btm.t513 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4274 VDAC_P.t1002 C9_P_btm.t502 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4275 a_601_44048# a_383_43806# VSS.t942 VSS.t941 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4276 VDAC_N.t1006 C10_N_btm.t512 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4277 VSS.t1182 a_10588_45670# a_10383_46697# VSS.t1181 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4278 VDAC_N.t1982 C9_N_btm.t264 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4279 VDAC_P.t1974 C10_P_btm.t504 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4280 VDD.t2810 a_11455_44576.t8 a_13023_44716# VDD.t2809 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X4281 VDAC_N.t150 C10_N_btm.t510 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4282 VDAC_N.t1978 C10_N_btm.t501 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4283 VDD.t373 a_n2661_45956.t9 a_22223_43494# VDD.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4284 a_6025_43806# a_4835_43806# a_5916_43806# VSS.t1005 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4285 a_15730_45670.t6 a_18971_44654# VDD.t1820 VDD.t1819 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4286 VDD.t3073 a_n1925_47044.t4 a_22591_43958# VDD.t3072 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4287 a_n2442_46526.t1 a_n2472_46500# VSS.t1670 VSS.t1669 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4288 a_17930_32299.t2 a_22591_44894# VDD.t2150 VDD.t2149 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4289 VDAC_N.t1002 C10_N_btm.t498 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4290 VDAC_P.t514 C10_P_btm.t503 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4291 VDD.t2396 VSS.t3676 VDD.t2395 VDD.t2394 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4292 a_18541_43582# a_15730_45670.t9 a_n2497_42870.t2 VSS.t563 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4293 VSS.t3108 VDD.t3138 VSS.t3107 VSS.t3106 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4294 a_12545_43268# a_12379_43268# VSS.t1158 VSS.t1157 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4295 a_13181_45982# a_14194_46348# a_14382_46348# VSS.t2609 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.151025 ps=1.285 w=0.42 l=0.15
X4296 a_18348_43262# a_18766_43236# VDD.t1335 VDD.t1334 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4297 VDAC_N.t1974 C10_N_btm.t497 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4298 VSS.t3219 VDD.t3176 VSS.t3218 VSS.t3217 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4299 VDD.t394 a_13248_45956.t6 a_16369_46232# VDD.t393 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
X4300 VDD.t2472 VSS.t3707 VDD.t2471 VDD.t2470 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X4301 VDAC_N.t514 C7_N_btm.t67 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4302 VDAC_N.t1970 C10_N_btm.t495 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4303 VDAC_P.t1970 C10_P_btm.t502 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4304 VDAC_P.t998 C10_P_btm.t1029 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4305 a_10197_45776# a_4908_45956# a_10111_45776# VSS.t1791 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4306 VDAC_N.t998 C10_N_btm.t494 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4307 VDAC_N.t1966 VSS.t3311 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4308 a_6974_31099.t3 a_20383_42718# VDD.t2225 VDD.t2224 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4309 a_16513_46642# a_13524_46832.t24 a_16426_46642# VDD.t555 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.05985 ps=0.705 w=0.42 l=0.15
X4310 VDAC_N.t270 C7_N_btm.t66 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4311 VDAC_P.t1966 C9_P_btm.t499 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4312 VDAC_N.t1962 C10_N_btm.t490 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4313 VDAC_P.t270 C9_P_btm.t452 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4314 VSS.t3773 C9_N_btm.t530 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4315 VDAC_N.t994 C9_N_btm.t524 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4316 VDAC_N.t1958 C9_N_btm.t261 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4317 VDAC_N.t510 C9_N_btm.t260 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4318 COMP_P.t0 a_1239_39587# VSS.t1769 VSS.t1768 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4319 VDD.t349 a_n690_43494.t4 a_n133_43806# VDD.t348 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4320 VDAC_P.t1962 C10_P_btm.t1019 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4321 VDD.t900 a_5839_47070# a_5847_47614# VDD.t899 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4322 VDAC_P.t994 C8_P_btm.t120 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4323 C10_P_btm.t1079 a_n2810_44894.t11 VSS.t3286 VSS.t3285 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X4324 a_18704_43806# a_17623_43806# a_18357_44048# VDD.t1885 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4325 VDAC_P.t1958 C10_P_btm.t993 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4326 a_13108_47320# a_4908_45956# VDD.t1744 VDD.t1743 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X4327 VDAC_N.t1954 C9_N_btm.t259 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4328 VDAC_P.t510 C9_P_btm.t397 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4329 VDAC_N.t990 C9_N_btm.t258 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4330 VDD.t1077 a_22223_46534# a_20163_31459.t2 VDD.t1076 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4331 VSS.t3808 C8_N_btm.t267 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4332 VDAC_P.t1954 VSS.t3386 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4333 VDAC_P.t990 C4_P_btm.t20 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4334 a_1304_44894# a_1053_45123.t8 a_1083_45221# VSS.t582 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4335 a_10467_47212# a_9521_45982.t7 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4336 VSS.t1713 a_6091_43780# a_1847_45528.t1 VSS.t1712 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4337 VDAC_P.t1950 C7_P_btm.t59 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4338 VDAC_P.t58 C10_P_btm.t965 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4339 VDAC_N.t1950 C10_N_btm.t489 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4340 VSS.t3481 VDD.t3220 VSS.t3480 VSS.t3479 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4341 VCM.t23 a_6974_31099.t5 C0_dummy_N_btm.t1 VSS.t306 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4342 VDAC_P.t1946 C10_P_btm.t929 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4343 VDAC_N.t58 C9_N_btm.t257 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4344 VSS.t3209 VDD.t3172 VSS.t3208 VSS.t3207 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4345 VDAC_P.t986 C10_P_btm.t867 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4346 VSS.t3138 VDD.t3148 VSS.t3137 VSS.t3136 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4347 VDAC_P.t1942 C9_P_btm.t377 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4348 a_n2073_43806# a_n2103_43780.t12 VSS.t2928 VSS.t2927 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4349 VDAC_P.t506 C9_P_btm.t350 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4350 a_5088_37509.t0 VSS.t3625 VDAC_Ni.t1 VDD.t2267 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X4351 VDAC_N.t1946 C10_N_btm.t487 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4352 VSS.t1113 a_12833_42718# a_13023_42718# VSS.t1112 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4353 a_13193_44716# a_11455_44576.t10 a_13105_44716# VSS.t2709 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X4354 a_3165_45982# a_2687_45956# VSS.t1461 VSS.t1460 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X4355 a_12121_45956# a_11788_46134# VDD.t1586 VDD.t1585 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4356 VDAC_P.t1938 C10_P_btm.t859 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4357 a_12_45982# a_n105_46195# VDD.t1938 VDD.t1937 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X4358 VDAC_N.t986 C10_N_btm.t486 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4359 VSS.t483 a_13248_45956.t14 a_13151_45956# VSS.t482 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4360 VDAC_P.t982 C10_P_btm.t768 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4361 a_5256_43806# a_5139_44019# VSS.t2060 VSS.t2059 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4362 VDAC_N.t1942 C10_N_btm.t483 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4363 VDAC_N.t506 C10_N_btm.t482 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4364 VCM.t63 a_4758_30651.t13 C9_P_btm.t540 VSS.t2995 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4365 a_14757_43806# a_14331_44133# VDD.t705 VDD.t704 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X4366 a_1057_43806# a_n133_43806# a_948_43806# VSS.t909 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4367 VDAC_N.t1938 C10_N_btm.t480 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4368 VDAC_P.t1934 C10_P_btm.t757 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4369 VSS.t988 a_n2833_42692# SMPL.t2 VSS.t987 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4370 VDAC_P.t266 C10_P_btm.t754 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4371 VSS.t699 a_5129_45956# a_5063_45982# VSS.t698 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4372 VDAC_N.t982 C8_N_btm.t161 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4373 VDAC_N.t1934 C10_N_btm.t479 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4374 a_4833_47070# a_n53_44363.t9 VSS.t618 VSS.t617 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4375 VDAC_N.t266 C8_N_btm.t119 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4376 VDAC_N.t1930 C10_N_btm.t473 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4377 VDAC_P.t1930 C9_P_btm.t298 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4378 VDAC_P.t978 C10_P_btm.t699 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4379 VDD.t3034 a_1736_39587.t3 a_1239_39587# VDD.t3033 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4380 a_8013_47098# a_n237_45454.t14 VSS.t497 VSS.t496 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X4381 VSS.t264 a_2587_44868.t22 a_10333_42718# VSS.t263 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4382 VDAC_P.t1926 C8_P_btm.t252 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4383 VDD.t2266 VSS.t3566 VDD.t2265 VDD.t2264 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4384 VDD.t1519 a_4091_47070# a_4651_47614# VDD.t738 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X4385 VDAC_N.t978 C10_N_btm.t472 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4386 VDD.t1833 a_15468_45412# a_11788_46134# VDD.t1832 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X4387 a_8483_43780# a_5655_43780# VDD.t2209 VDD.t2208 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4388 VSS.t1819 a_4322_46134# a_5626_46846# VSS.t1818 sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X4389 VDAC_N.t1926 C8_N_btm.t118 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4390 a_13101_44894# a_927_42692.t22 a_13013_44894# VSS.t99 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X4391 VDAC_P.t502 C7_P_btm.t126 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4392 VSS.t2972 a_13458_32299.t4 C0_N_btm.t5 VSS.t2706 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4393 a_13819_44350# a_10114_45276.t8 a_13725_44350# VDD.t170 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X4394 VDAC_P.t1922 C5_P_btm.t17 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4395 VDAC_P.t974 C10_P_btm.t629 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4396 VDAC_N.t502 C6_N_btm.t33 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4397 VSS.t3560 C8_P_btm.t9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4398 VDAC_N.t1922 C10_N_btm.t470 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4399 a_491_44172# a_135_43540.t32 VDD.t182 VDD.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X4400 a_n2840_44868# a_n2661_44868# VDD.t849 VDD.t306 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X4401 VDAC_P.t1918 VSS.t3384 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4402 a_18135_47588# DEBUG_MUX[0].t1 VDD.t154 VDD.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X4403 VDAC_N.t974 C10_N_btm.t469 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4404 w_1375_34946.t15 a_n1732_35090.t11 EN_VIN_BSTR_P.t5 w_1375_34946.t14 sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X4405 VDD.t2270 VSS.t3554 VDD.t2269 VDD.t2268 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4406 VDAC_N.t1918 C9_N_btm.t256 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4407 VDAC_P.t146 C10_P_btm.t522 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4408 VSS.t2276 a_n2840_46500# a_n2810_46526.t1 VSS.t2126 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4409 VDAC_N.t146 C10_N_btm.t465 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4410 VSS.t1515 a_6631_44582# a_5419_47258# VSS.t1514 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4411 a_10537_46224# a_10319_45982# VSS.t1554 VSS.t1553 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4412 VDAC_N.t1914 C9_N_btm.t255 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4413 VCM.t29 a_3222_30651.t5 VDAC_N.t1 VSS.t657 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4414 VSS.t711 a_15437_47044# a_15691_47436# VSS.t710 sky130_fd_pr__nfet_01v8 ad=0.1359 pd=1.1 as=0.1113 ps=1.37 w=0.42 l=0.15
X4415 VDAC_P.t1914 C10_P_btm.t517 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4416 VDAC_N.t1910 C10_N_btm.t466 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4417 VDAC_N.t498 C10_N_btm.t464 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4418 VDAC_P.t970 C10_P_btm.t516 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4419 w_11534_34010.t12 a_11730_34132.t4 w_11534_34010.t11 w_11534_34010.t10 sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X4420 VDAC_P.t1910 C9_P_btm.t292 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4421 VDAC_N.t1906 C9_N_btm.t523 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4422 VDAC_N.t966 C10_N_btm.t463 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4423 VDAC_N.t1902 C10_N_btm.t462 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4424 VSS.t2115 a_2471_45046# a_171_44019# VSS.t2114 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X4425 VDAC_P.t498 C9_P_btm.t267 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4426 VDAC_P.t1906 C10_P_btm.t510 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4427 VSS.t2766 a_885_44868.t36 a_829_45221# VSS.t2765 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X4428 VDAC_N.t262 C10_N_btm.t461 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4429 VDAC_P.t966 C10_P_btm.t509 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4430 a_10069_42968# a_10259_42870.t8 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4431 VDAC_P.t1902 C10_P_btm.t500 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4432 VDAC_N.t1898 C8_N_btm.t116 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4433 VSS.t2625 a_n2038_35608# SMPL_ON_P.t2 VSS.t2624 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4434 VDAC_N.t962 C10_N_btm.t460 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4435 VDAC_P.t262 C8_P_btm.t246 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4436 VDAC_N.t1894 C10_N_btm.t459 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4437 VDAC_N.t494 C10_N_btm.t458 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4438 VSS.t2147 a_6635_47044# a_n690_43494.t0 VSS.t2146 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X4439 VSS.t752 a_22223_43494# a_22223_43270# VSS.t751 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4440 VSS.t3 a_10259_42870.t10 a_12636_45758# VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.08775 ps=0.92 w=0.65 l=0.15
X4441 VDAC_P.t1898 C10_P_btm.t499 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4442 a_7648_46892# a_7503_45982# VSS.t1352 VSS.t1351 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4443 VDAC_N.t1890 C10_N_btm.t457 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4444 VDD.t1929 a_11248_47319# a_11186_47436# VDD.t1928 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X4445 VDAC_N.t958 C9_N_btm.t522 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4446 VDAC_P.t962 C9_P_btm.t261 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4447 VDD.t928 a_n2833_42692# SMPL.t6 VDD.t927 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4448 VDAC_N.t1886 C8_N_btm.t115 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4449 a_491_44172# a_n133_43806# a_383_43806# VDD.t851 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4450 VDAC_P.t1894 C9_P_btm.t257 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4451 VSS.t2462 VSS.t2463 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4452 VDAC_P.t494 C5_P_btm.t36 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4453 VDAC_N.t86 C8_N_btm.t114 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4454 VDAC_P.t1890 C6_P_btm.t62 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4455 VDAC_N.t1882 C4_N_btm.t10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4456 a_15468_45412# a_15730_45670.t24 a_15688_45758# VSS.t576 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4457 VDAC_N.t954 C10_N_btm.t456 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4458 VDAC_P.t958 C9_P_btm.t256 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4459 VDD.t1123 a_989_45736# a_1019_45477# VDD.t1122 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4460 VDD.t1726 a_1239_39043# COMP_N.t5 VDD.t1725 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4461 VDAC_N.t1878 C10_N_btm.t455 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4462 a_18822_46526# a_18064_46642# a_18259_46500# VDD.t1801 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X4463 VDAC_N.t490 C8_N_btm.t113 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4464 VDAC_P.t1886 C10_P_btm.t496 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4465 a_10857_46892# a_10813_46500# a_10691_46904# VSS.t1951 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X4466 VDAC_P.t86 C10_P_btm.t495 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4467 VDAC_N.t1874 C9_N_btm.t520 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4468 VDAC_P.t1882 C9_P_btm.t253 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4469 DATA[4].t4 a_5847_47614# VDD.t1866 VDD.t1865 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X4470 VDD.t2621 VSS.t3751 VDD.t2620 VDD.t2619 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4471 VDAC_N.t950 C10_N_btm.t454 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4472 VDAC_N.t1870 C10_N_btm.t453 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4473 VDAC_N.t258 C10_N_btm.t452 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4474 VDD.t1890 a_21540_43236# a_13458_32299.t2 VDD.t1889 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4475 VSS.t2403 VSS.t2404 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4476 VDD.t2612 VSS.t3655 VDD.t2611 VDD.t2610 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4477 VDAC_P.t954 C10_P_btm.t493 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4478 VDAC_N.t1866 C10_N_btm.t451 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4479 a_4355_45438# a_3731_45444# a_4247_45816# VDD.t2117 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4480 VDAC_P.t1878 C10_P_btm.t492 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4481 VDAC_P.t490 C10_P_btm.t488 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4482 VDAC_N.t946 C10_N_btm.t450 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4483 VDAC_P.t1874 C10_P_btm.t487 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4484 VDAC_N.t1862 C9_N_btm.t518 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4485 VDD.t150 CAL_N.t5 VDD.t149 VDD.t148 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=10
X4486 a_6152_46348# a_5715_45956# VDD.t940 VDD.t939 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4487 VDAC_N.t486 C10_N_btm.t449 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4488 VDAC_P.t950 C10_P_btm.t485 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4489 a_19633_43262# a_19191_43262# VSS.t1785 VSS.t1784 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258375 ps=1.445 w=0.65 l=0.15
X4490 VSS.t1475 a_713_47044# a_647_47070# VSS.t1474 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4491 a_1346_46892# a_885_44868.t38 VSS.t2768 VSS.t2767 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4492 a_82_45670# a_847_45956# VDD.t1625 VDD.t1624 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X4493 a_9573_44716# a_5655_43780# VSS.t2238 VSS.t2237 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X4494 VDAC_P.t1870 C8_P_btm.t233 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4495 VDAC_P.t258 C10_P_btm.t484 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4496 VDD.t1137 a_22959_47070# a_21276_30659.t3 VDD.t1136 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4497 VDAC_N.t1858 C7_N_btm.t130 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4498 C10_N_btm.t32 a_22812_30659.t18 VREF.t43 VDD.t530 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4499 a_2675_46565# a_2424_46794.t2 a_2216_46758# VDD.t2942 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X4500 VSS.t1374 a_16921_46364# a_16750_46134# VSS.t1373 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4501 VSS.t3443 VDD.t3206 VSS.t3442 VSS.t3112 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4502 VSS.t1738 a_7429_47044# a_7363_47070# VSS.t1737 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4503 VDAC_P.t1866 C10_P_btm.t481 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4504 VSS.t1957 a_16579_43566# a_12651_44576.t3 VSS.t1956 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4505 a_16670_44324# a_16824_45276# VDD.t1989 VDD.t1988 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.17575 ps=1.395 w=0.42 l=0.15
X4506 VDAC_N.t942 C5_N_btm.t27 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4507 VDAC_N.t1854 C8_N_btm.t112 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4508 VDAC_P.t946 C8_P_btm.t221 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4509 VDAC_P.t1862 C3_P_btm.t9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4510 a_21997_47833# SMPL_ON_N.t8 VDD.t108 VDD.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4511 VDD.t1384 a_2655_42870# a_2627_42718# VDD.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X4512 VDAC_N.t142 C8_N_btm.t111 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4513 VDAC_P.t486 C7_P_btm.t58 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4514 C9_N_btm.t5 a_21788_30659.t4 VREF.t23 VDD.t2051 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4515 a_18845_42746# a_1581_43806.t10 a_18759_42746# VSS.t2875 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4516 a_17156_43806# a_13273_44868.t18 VSS.t643 VSS.t642 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X4517 a_8417_46904# a_7227_46532# a_8308_46904# VSS.t1277 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4518 VDD.t788 a_10537_46224# a_10427_46348# VDD.t787 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4519 VDAC_P.t1858 C10_P_btm.t480 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4520 VDAC_N.t1850 VSS.t3316 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4521 VDD.t2600 VSS.t3591 VDD.t2599 VDD.t2417 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4522 VSS.t2828 a_135_43540.t16 a_93_43628# VSS.t2827 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4523 VDAC_N.t938 C10_N_btm.t447 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4524 VDAC_N.t1846 C9_N_btm.t514 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4525 VDAC_P.t942 C10_P_btm.t478 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4526 VDD.t1924 a_10415_47846# a_9517_46539# VDD.t1923 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X4527 VDAC_N.t482 C10_N_btm.t446 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4528 a_n2840_43780# a_n2661_43780# VDD.t2123 VDD.t2122 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X4529 VDAC_N.t1842 C9_N_btm.t512 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4530 VDAC_P.t1854 C9_P_btm.t246 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4531 VDAC_N.t934 C10_N_btm.t445 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4532 VDAC_P.t142 C10_P_btm.t477 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4533 a_885_44868.t3 a_2587_44868.t24 VDD.t245 VDD.t244 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4534 VDAC_P.t1850 C10_P_btm.t471 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4535 VDAC_N.t1838 C9_N_btm.t510 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4536 VDAC_P.t938 C10_P_btm.t470 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4537 VDAC_P.t1846 C9_P_btm.t241 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4538 VDAC_N.t254 C8_N_btm.t110 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4539 VDAC_N.t1834 C9_N_btm.t249 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4540 VDAC_P.t482 C9_P_btm.t240 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4541 VDAC_P.t1842 VSS.t3381 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4542 VDAC_P.t934 C6_P_btm.t27 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4543 a_7961_44048# a_7743_43806# VDD.t955 VDD.t954 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4544 a_15008_42692# a_15133_43582# VSS.t1256 VSS.t1255 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4545 a_n1551_44324.t6 a_1053_45123.t10 VDD.t514 VDD.t513 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4546 VDD.t2583 VSS.t3671 VDD.t2582 VDD.t2581 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4547 VDAC_N.t930 VSS.t3261 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4548 a_702_45477# a_656_45670# VDD.t963 VDD.t962 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4549 a_4322_46134# a_4527_46830# VDD.t1758 VDD.t1757 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4550 a_49_43236# a_n169_43640# VDD.t719 VDD.t718 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4551 a_n2109_42692.t3 a_9521_45982.t6 VSS.t25 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4552 VSS.t2307 VSS.t2308 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4553 VDAC_N.t1830 C10_N_btm.t444 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4554 VDAC_P.t1838 C10_P_btm.t467 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4555 a_n2497_42870.t4 a_13273_44868.t9 a_18093_43262# VDD.t610 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4556 VDAC_P.t254 C9_P_btm.t238 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4557 VDAC_N.t478 C6_N_btm.t32 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4558 VDAC_N.t1826 C10_N_btm.t443 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4559 a_5896_45670# a_5382_44582# a_6038_45477# VDD.t2024 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4560 VDAC_P.t1834 C9_P_btm.t237 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4561 a_505_46904# a_n685_46532# a_396_46904# VSS.t1639 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4562 a_7418_45477# a_7372_45670# VDD.t680 VDD.t679 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4563 VDAC_N.t926 C8_N_btm.t109 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4564 VDAC_P.t930 C9_P_btm.t234 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4565 VDAC_P.t1830 C8_P_btm.t190 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4566 a_5916_43806# a_5001_43806# a_5569_44048# VSS.t1227 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4567 VSS.t2533 VSS.t2534 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4568 VDAC_P.t478 C5_P_btm.t35 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4569 VDAC_P.t1826 C8_P_btm.t188 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4570 VDAC_N.t1822 C9_N_btm.t508 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4571 VSS.t2379 VSS.t2380 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4572 VDAC_P.t926 C8_P_btm.t175 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4573 a_7694_45982# a_7648_46134# VSS.t1556 VSS.t1555 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4574 VDAC_N.t42 C10_N_btm.t442 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4575 VDAC_N.t1818 C10_N_btm.t441 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4576 VSS.t1978 a_11248_47319# a_11186_47436# VSS.t1977 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X4577 a_1633_46824# a_885_44868.t22 VDD.t2842 VDD.t2841 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4578 VDAC_N.t922 C10_N_btm.t440 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4579 a_7839_43806# a_7393_43806# a_7743_43806# VSS.t1596 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4580 VDAC_P.t1822 C9_P_btm.t233 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4581 VDAC_N.t1814 C9_N_btm.t500 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4582 VDAC_P.t42 C10_P_btm.t468 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4583 VSS.t501 a_n237_45454.t18 a_n291_45776# VSS.t500 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4584 VDAC_P.t1818 C10_P_btm.t466 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4585 VDAC_P.t922 C8_P_btm.t168 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4586 VDAC_P.t1814 C10_P_btm.t465 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4587 VSS.t3282 a_n2810_44894.t9 C10_P_btm.t1077 VSS.t3281 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4588 VSS.t1395 a_2343_47070# a_2351_47614# VSS.t1394 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X4589 a_4461_46904# a_3271_46532# a_4352_46904# VSS.t1681 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4590 VSS.t326 a_n1827_44868.t13 a_n2293_43780# VSS.t303 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4591 a_10245_46532# a_10079_46532# VDD.t2221 VDD.t2220 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4592 a_107_45982# a_n243_45982# a_12_45982# VDD.t2193 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4593 a_2687_45956# a_135_43540.t15 VDD.t2926 VDD.t2925 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4594 a_1387_44582# a_1659_44440# VSS.t1178 VSS.t1177 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4595 VDAC_N.t474 C9_N_btm.t499 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4596 a_999_47846# a_1209_47588# VDD.t1956 VDD.t1955 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4597 a_13654_46032# a_14194_46348# a_14382_46348# VDD.t2703 sky130_fd_pr__pfet_01v8_hvt ad=0.2688 pd=2.12 as=0.092075 ps=0.99 w=0.42 l=0.15
X4598 VDAC_N.t1810 C8_N_btm.t108 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4599 VDAC_P.t474 C3_P_btm.t8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4600 a_4830_43958.t3 a_9395_47044# VDD.t1188 VDD.t1187 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4601 a_22455_45420# a_n2109_47596.t8 VDD.t382 VDD.t381 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4602 a_3540_44466# a_3165_45982# VDD.t1395 VDD.t1394 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X4603 a_13878_32299.t2 a_21908_43236# VDD.t1966 VDD.t1965 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4604 a_15443_44582# a_12651_44576.t12 a_15589_44350# VDD.t2960 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4605 a_95_44716# a_n53_44363.t10 a_n268_44582# VSS.t619 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4606 VDAC_P.t1810 C10_P_btm.t463 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4607 VDAC_N.t918 C6_N_btm.t31 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4608 VDAC_N.t1806 C10_N_btm.t439 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4609 VDAC_N.t250 C4_N_btm.t18 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4610 a_3320_46134# a_3470_45982# VSS.t1595 VSS.t1594 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X4611 a_15744_43628# a_15415_44350# VDD.t711 VDD.t710 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X4612 VDAC_N.t1802 C7_N_btm.t64 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4613 VDAC_N.t914 C9_N_btm.t355 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4614 VDAC_P.t918 C8_P_btm.t129 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4615 VDAC_N.t1798 C8_N_btm.t107 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4616 VDAC_P.t1806 C8_P_btm.t128 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4617 VDAC_N.t470 C10_N_btm.t438 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4618 VSS.t1919 a_7754_38470# a_7754_38470# VSS.t1918 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4619 VDAC_P.t250 C9_P_btm.t231 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4620 VDAC_P.t1802 C10_P_btm.t462 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4621 a_22780_40293# a_22465_38541# a_22521_39947# VSS.t2693 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4622 a_8204_45412# a_8055_45491# a_8500_45554# VDD.t2694 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4623 VDAC_P.t914 C8_P_btm.t122 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4624 VDAC_P.t1798 C10_P_btm.t461 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4625 VDAC_P.t470 C9_P_btm.t230 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4626 VDAC_N.t1794 C10_N_btm.t437 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4627 VDAC_N.t910 C10_N_btm.t436 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4628 VDAC_P.t1794 VSS.t3389 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4629 VDAC_P.t910 C9_P_btm.t226 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4630 VDAC_N.t1790 C9_N_btm.t314 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4631 a_8912_37509.t15 VDAC_N.t138 a_5700_37509.t9 VDD.t2240 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4632 VDAC_P.t1790 C9_P_btm.t225 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4633 VDAC_P.t138 C10_P_btm.t460 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4634 a_16585_46642# a_16555_46616# a_16513_46642# VDD.t1124 sky130_fd_pr__pfet_01v8_hvt ad=0.1215 pd=1.33 as=0.0441 ps=0.63 w=0.42 l=0.15
X4635 VDAC_N.t1786 C10_N_btm.t435 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4636 a_22705_38426# a_22521_40491# a_22609_38426# VDD.t1474 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X4637 a_15376_43806# a_14757_43806# VDD.t1121 VDD.t1120 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X4638 VDAC_N.t906 C9_N_btm.t288 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4639 VDAC_N.t1782 C10_N_btm.t434 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4640 a_8798_45758# a_8850_45412# a_n1827_44868.t2 VSS.t730 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4641 a_560_45670# a_n53_44363.t12 a_702_45477# VDD.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4642 VDAC_N.t466 C10_N_btm.t433 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4643 VDAC_N.t1778 C10_N_btm.t432 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4644 VDD.t1850 a_11252_43640# a_11427_43566# VDD.t1849 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4645 VDAC_P.t1786 C10_P_btm.t459 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4646 VSS.t1744 a_22591_47070# a_21020_30659.t1 VSS.t1743 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4647 VDAC_N.t902 C6_N_btm.t30 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4648 a_2301_45758# a_n53_44363.t16 VSS.t622 VSS.t621 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X4649 VDAC_P.t906 C10_P_btm.t458 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4650 a_10808_44466# a_1053_45123.t7 VDD.t512 VDD.t511 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X4651 VDAC_N.t1774 C9_N_btm.t253 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4652 VDAC_P.t1782 C7_P_btm.t124 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4653 VDAC_N.t246 C9_N_btm.t251 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4654 VDAC_P.t466 C9_P_btm.t223 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4655 VDD.t698 a_n2288_42692# EN_COMP.t2 VDD.t697 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4656 a_6485_44582.t1 a_8483_43780# VSS.t968 VSS.t967 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4657 a_8379_46134# a_1429_47222.t5 VSS.t378 VSS.t377 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X4658 a_n2103_43780.t7 a_3882_44324# VDD.t1991 VDD.t1990 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4659 VDAC_P.t1778 C9_P_btm.t222 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4660 VDAC_N.t1770 C8_N_btm.t106 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4661 VDD.t1359 a_14950_43958# a_17715_44356# VDD.t1358 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4662 VSS.t2517 VSS.t2518 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4663 DATA[2].t7 a_2351_47614# VDD.t2006 VDD.t2005 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4664 VDAC_P.t902 C5_P_btm.t34 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4665 VDAC_P.t1774 C10_P_btm.t457 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4666 VSS.t2291 VSS.t2292 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4667 VDAC_P.t246 C10_P_btm.t456 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4668 a_2684_37794# VDAC_Pi.t9 a_2113_38308# VSS.t2970 sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X4669 VDAC_N.t898 C6_N_btm.t64 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4670 VDAC_N.t1766 C9_N_btm.t250 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4671 a_15877_44670# a_13715_43780# a_15443_44582# VSS.t1261 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4672 VDAC_N.t462 C10_N_btm.t431 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4673 VIN_N.t6 EN_VIN_BSTR_N.t21 C9_N_btm.t4 VSS.t448 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X4674 VDAC_N.t1762 C8_N_btm.t105 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4675 VDAC_P.t1770 VSS.t3387 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4676 VDAC_N.t894 C9_N_btm.t245 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4677 VDAC_P.t898 C8_P_btm.t119 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4678 VDAC_N.t1758 C10_N_btm.t430 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4679 VDAC_N.t82 C9_N_btm.t244 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4680 VDAC_P.t1766 C9_P_btm.t218 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4681 VSS.t2708 a_11455_44576.t9 a_13464_45758# VSS.t2707 sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.08775 ps=0.92 w=0.65 l=0.15
X4682 VSS.t2325 VSS.t2326 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4683 VDAC_N.t1754 C9_N_btm.t242 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4684 VDAC_P.t462 C9_P_btm.t219 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4685 VDAC_N.t890 C10_N_btm.t429 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4686 VDAC_P.t1762 C9_P_btm.t217 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4687 VDAC_N.t1750 C10_N_btm.t428 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4688 DATA[0].t0 a_n1085_47874# VSS.t1998 VSS.t1997 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4689 VDAC_N.t458 C8_N_btm.t104 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4690 VDAC_P.t894 C9_P_btm.t216 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4691 VDAC_N.t1746 C10_N_btm.t427 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4692 a_17821_46892# a_17786_46658# a_17583_46500# VSS.t1576 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X4693 VSS.t3120 VDD.t3142 VSS.t3119 VSS.t3118 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X4694 a_15744_43628# a_15415_44350# VSS.t782 VSS.t781 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4695 a_2055_46348# a_135_43540.t14 VDD.t2924 VDD.t2923 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X4696 a_9475_46565# a_9293_46565# VDD.t3092 VDD.t3091 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4697 VDAC_N.t886 C7_N_btm.t63 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4698 a_6208_46642# a_5784_44364# a_6126_46642# VDD.t919 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4699 a_n2472_44868# a_n2293_44868# VDD.t1423 VDD.t1422 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X4700 VDAC_P.t1758 C7_P_btm.t118 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4701 C9_N_btm.t3 a_17930_32299.t7 VSS.t314 VSS.t313 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4702 a_22223_43494# a_n2661_45956.t8 VDD.t371 VDD.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4703 a_n1435_47614.t1 a_n1605_47614# VDD.t618 VDD.t617 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4704 VDD.t1233 a_284_47222# a_n381_46697# VDD.t1232 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X4705 VDAC_N.t1742 C9_N_btm.t241 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4706 a_n2293_44868# a_n2103_44868.t13 VDD.t2936 VDD.t2873 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4707 VDAC_P.t82 C5_P_btm.t33 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4708 a_571_43566# a_135_43540.t46 VDD.t194 VDD.t193 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4709 VDAC_P.t1754 C6_P_btm.t68 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4710 a_18348_43262# a_15730_45670.t18 VDD.t495 VDD.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4711 a_22591_43958# a_n1925_47044.t8 VDD.t3077 VDD.t3076 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4712 VSS.t1668 a_n2472_46500# a_n2442_46526.t0 VSS.t1667 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4713 VSS.t736 a_22223_43270# a_14087_32299.t0 VSS.t735 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4714 VSS.t2048 a_2351_47614# DATA[2].t1 VSS.t2047 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4715 VSS.t1019 a_19037_42718# a_22223_42718# VSS.t1018 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4716 VDAC_P.t890 C9_P_btm.t215 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4717 a_n268_44582# a_n53_44363.t4 a_n126_44389# VDD.t556 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4718 VDAC_P.t1750 C10_P_btm.t455 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4719 C3_P_btm.t0 EN_VIN_BSTR_P.t21 VIN_P.t6 VSS.t552 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X4720 VDAC_N.t242 C6_N_btm.t63 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4721 a_n2038_35608# a_n1586_35608# VSS.t1389 VSS.t1388 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4722 VDAC_P.t458 C10_P_btm.t454 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4723 VDAC_N.t1738 C9_N_btm.t238 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4724 VDAC_N.t882 C9_N_btm.t237 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4725 VDAC_P.t1746 C8_P_btm.t116 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4726 VSS.t3568 C8_N_btm.t271 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4727 a_16369_46232# a_15328_46134# a_16273_46232# VDD.t1436 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X4728 VDAC_N.t1734 C9_N_btm.t235 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4729 VDAC_N.t454 C10_N_btm.t426 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4730 VDAC_P.t886 C10_P_btm.t453 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4731 a_12623_43780# a_10227_47214.t20 VDD.t293 VDD.t292 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4732 VDAC_P.t1742 C8_P_btm.t115 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4733 VDAC_N.t1730 C9_N_btm.t234 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4734 VDAC_P.t242 C9_P_btm.t214 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4735 VDAC_N.t878 C10_N_btm.t425 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4736 VDAC_P.t1738 C9_P_btm.t213 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4737 VSS.t161 a_10114_45276.t10 a_9943_45046# VSS.t160 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4738 VDD.t2534 VSS.t3653 VDD.t2533 VDD.t2532 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X4739 VDAC_P.t882 C10_P_btm.t452 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4740 a_6631_44582# a_7195_44868# VDD.t2195 VDD.t2194 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X4741 VDAC_P.t1734 C10_P_btm.t451 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4742 VREF.t30 a_21788_30659.t11 C9_N_btm.t12 VDD.t2058 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4743 a_14757_45982# a_14382_46348# VSS.t1285 VSS.t1284 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4744 a_15112_45798# a_15033_46526# a_15040_45798# VSS.t1895 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X4745 a_4514_46526# a_3437_46532# a_4352_46904# VDD.t1828 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X4746 VDAC_P.t454 C10_P_btm.t450 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4747 VDAC_N.t1726 C7_N_btm.t62 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4748 a_3883_43640# a_3437_43268# a_3787_43640# VSS.t1672 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4749 VDAC_N.t134 C10_N_btm.t424 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4750 a_1567_46892# a_n194_47222# a_1204_46758# VSS.t1034 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4751 w_1375_34946.t9 a_n1123_35174.t7 w_1375_34946.t8 w_1375_34946.t5 sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X4752 VDAC_N.t1722 C6_N_btm.t62 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4753 VDAC_N.t874 C9_N_btm.t233 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4754 VDD.t3066 a_n2661_47044.t9 a_22031_45438# VDD.t3065 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4755 VDAC_P.t1730 C7_P_btm.t117 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4756 VDAC_N.t1718 C10_N_btm.t423 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4757 VDAC_P.t878 C9_P_btm.t212 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4758 VDD.t1464 a_9343_45982# a_9521_45982.t2 VDD.t1463 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4759 VDD.t1037 a_20159_47588# a_13248_45956.t3 VDD.t1036 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4760 VDAC_N.t450 C8_N_btm.t102 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4761 VDAC_P.t1726 C7_P_btm.t97 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4762 VDAC_P.t134 C10_P_btm.t449 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4763 VDAC_P.t1722 C7_P_btm.t80 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4764 VDAC_P.t874 C9_P_btm.t211 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4765 VDAC_P.t1718 C10_P_btm.t448 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4766 VDD.t2519 VSS.t3760 VDD.t2518 VDD.t2517 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4767 VDD.t214 a_7557_43236.t12 a_13023_44716# VDD.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X4768 a_1847_45528.t0 a_6091_43780# VSS.t1719 VSS.t1718 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4769 VSS.t2539 VSS.t2540 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4770 VCM.t43 a_3222_30651.t8 VDAC_P.t1 VSS.t660 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4771 VSS.t670 a_3222_30651.t18 a_21027_42718# VSS.t669 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4772 VDAC_N.t1714 C10_N_btm.t422 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4773 VSS.t3057 VDD.t3121 VSS.t3056 VSS.t3055 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4774 VDD.t2513 VSS.t3811 VDD.t2512 VDD.t2287 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4775 VDAC_P.t1714 C10_P_btm.t447 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4776 VDAC_P.t870 C10_P_btm.t446 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4777 VDAC_N.t870 C9_N_btm.t232 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4778 VDAC_N.t1710 C10_N_btm.t421 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4779 VDAC_N.t238 C9_N_btm.t231 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4780 VSS.t2926 a_n2103_43780.t9 a_n2073_43806# VSS.t2925 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4781 VDAC_N.t1706 C10_N_btm.t420 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4782 VDAC_P.t1710 C10_P_btm.t445 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4783 a_2627_43262# a_2755_43494.t23 a_2709_43262# VDD.t433 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4784 VDAC_P.t238 C8_P_btm.t113 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4785 VDAC_N.t866 C10_N_btm.t419 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4786 VSS.t990 a_n2833_42692# SMPL.t0 VSS.t989 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X4787 a_n2810_43262.t2 a_n2840_43236# VDD.t888 VDD.t887 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4788 VDAC_N.t1702 C10_N_btm.t418 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4789 VDAC_P.t1706 C9_P_btm.t210 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4790 VDAC_N.t446 C10_N_btm.t417 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4791 VDAC_N.t1698 C10_N_btm.t416 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4792 VSS.t2813 a_1334_43494.t9 a_6767_44716# VSS.t2812 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X4793 VDAC_P.t866 C10_P_btm.t444 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4794 a_8308_46904# a_7393_46532# a_7961_46500# VSS.t1279 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4795 VDAC_P.t1702 C10_P_btm.t443 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4796 VDAC_P.t446 C8_P_btm.t112 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4797 VDAC_P.t1698 C10_P_btm.t442 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4798 VDD.t2508 VSS.t3599 VDD.t2507 VDD.t2506 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4799 VDAC_N.t862 C10_N_btm.t415 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4800 VDD.t541 a_n1459_43236.t10 a_n1429_43262# VDD.t540 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4801 VSS.t707 a_18879_45956# a_18813_45982# VSS.t706 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4802 a_18530_47070# a_14757_47614# a_18444_47070# VSS.t1496 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X4803 VDAC_N.t1694 C10_N_btm.t414 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4804 a_n99_45438.t0 a_n377_45776# VSS.t2703 VSS.t2702 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X4805 a_9645_44716# a_9266_44350# a_9573_44716# VSS.t2645 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X4806 VDAC_N.t54 C6_N_btm.t27 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4807 a_19274_43262# a_2587_44868.t14 VDD.t237 VDD.t236 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4808 VDD.t2502 VSS.t3695 VDD.t2501 VDD.t2500 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X4809 VDAC_P.t862 C10_P_btm.t441 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4810 VDAC_N.t1690 C7_N_btm.t129 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4811 a_4322_46134# a_4527_46830# VDD.t1752 VDD.t1751 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4812 VDAC_P.t1694 C10_P_btm.t440 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4813 a_2332_44670# a_82_45670# a_2082_44670# VSS.t1691 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4814 VDAC_N.t858 C5_N_btm.t28 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4815 VDD.t1510 a_4061_45956# a_3575_46697# VDD.t1509 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4816 a_n2472_43780# a_n2293_43780# VDD.t1141 VDD.t1140 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X4817 VDAC_P.t54 C8_P_btm.t107 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4818 VDAC_N.t1686 C10_N_btm.t413 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4819 VDD.t1126 a_2645_46824# a_2675_46565# VDD.t1125 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4820 VSS.t392 a_1429_47222.t20 a_1387_45670# VSS.t391 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4821 a_702_45804# a_656_45670# VSS.t1025 VSS.t1024 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4822 a_17531_44894# a_14204_44350# VDD.t1921 VDD.t1920 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.182 ps=1.92 w=0.7 l=0.15
X4823 VDD.t2121 a_4005_46500# a_3895_46526# VDD.t2120 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4824 VDAC_N.t442 C9_N_btm.t230 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4825 VDAC_P.t1690 C8_P_btm.t106 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4826 VDAC_P.t858 C10_P_btm.t439 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4827 VDD.t2186 a_1431_47070# a_1203_42692.t4 VDD.t2185 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X4828 VCM.t5 a_3990_30651.t5 C10_N_btm.t9 VSS.t278 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4829 VREF.t7 a_20405_31459.t4 C4_N_btm.t0 VDD.t172 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X4830 VDAC_P.t1686 C10_P_btm.t438 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4831 VDAC_N.t1682 C10_N_btm.t411 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4832 VSS.t3605 C8_P_btm.t13 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4833 a_107_45982# a_n409_45982# a_12_45982# VSS.t1037 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4834 VDD.t2922 a_7029_44350.t3 a_13819_44350# VDD.t2921 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.16 ps=1.32 w=1 l=0.15
X4835 a_7418_45804# a_7372_45670# VSS.t748 VSS.t747 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4836 VDAC_P.t442 C10_P_btm.t437 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4837 VDAC_N.t854 C10_N_btm.t410 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4838 VDAC_N.t1678 C10_N_btm.t409 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4839 VDAC_P.t1682 C10_P_btm.t436 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4840 VDAC_N.t234 C10_N_btm.t408 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4841 a_7915_45982# a_n53_44363.t8 a_7552_46134# VSS.t616 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4842 VDAC_P.t854 C9_P_btm.t209 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4843 VDAC_N.t1674 C8_N_btm.t101 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4844 VDAC_N.t850 C10_N_btm.t407 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4845 VDAC_N.t1670 C10_N_btm.t406 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4846 a_n264_43628# a_n381_43433# VSS.t1891 VSS.t1890 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4847 a_396_46904# a_n519_46532# a_49_46500# VSS.t1135 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4848 VDAC_P.t1678 C10_P_btm.t435 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4849 VDAC_N.t438 C8_N_btm.t100 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4850 VDAC_N.t1666 C10_N_btm.t405 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4851 VDAC_N.t846 C10_N_btm.t404 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4852 a_14647_43494# a_10251_45454# VDD.t1295 VDD.t1294 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X4853 VDD.t807 a_6673_45136# a_6563_45260# VDD.t806 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4854 VSS.t1200 a_7552_46134# a_7503_45982# VSS.t1199 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4855 VDAC_P.t234 C10_P_btm.t434 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4856 VSS.t3724 C4_P_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4857 VDD.t289 a_10227_47214.t14 a_18404_46526# VDD.t288 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X4858 VDAC_P.t1674 C9_P_btm.t208 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4859 C6_N_btm.t70 a_14601_32299.t4 VSS.t2834 VSS.t2833 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X4860 VSS.t3035 VDD.t3113 VSS.t3034 VSS.t3033 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4861 VDAC_P.t850 C10_P_btm.t433 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4862 VDAC_P.t1670 C10_P_btm.t432 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4863 SMPL_ON_P.t1 a_n2038_35608# VSS.t2627 VSS.t2626 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4864 VDD.t2493 VSS.t3619 VDD.t2492 VDD.t2491 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X4865 VDAC_P.t438 C9_P_btm.t207 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4866 a_n1732_35090.t0 SMPL.t9 VDD.t3045 VDD.t3044 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4867 VSS.t2564 a_19187_42718# a_3990_30651.t0 VSS.t2563 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4868 VDD.t930 a_n2833_42692# SMPL.t7 VDD.t929 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X4869 VDAC_N.t1662 C8_N_btm.t258 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4870 a_4352_46904# a_3437_46532# a_4005_46500# VSS.t1872 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4871 VDAC_P.t1666 C10_P_btm.t431 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4872 VDAC_P.t846 C10_P_btm.t430 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4873 VDAC_N.t130 C6_N_btm.t50 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4874 a_7309_44466# a_6485_44582.t22 VDD.t3022 VDD.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4875 a_12636_45758# a_10259_42870.t9 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4876 a_n2810_44894.t1 a_n2840_44868# VSS.t1376 VSS.t935 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4877 VDAC_N.t1658 C7_N_btm.t60 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4878 a_16177_45982# a_16128_46134# a_16085_45982# VSS.t802 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.2015 ps=1.92 w=0.65 l=0.15
X4879 VDAC_N.t842 C6_N_btm.t58 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4880 VDAC_N.t1654 C10_N_btm.t403 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4881 VSS.t679 a_n1735_43236.t12 a_n1741_42692# VSS.t678 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4882 VSS.t3794 C10_P_btm.t11 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4883 VDAC_P.t1662 C8_P_btm.t104 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4884 VDAC_N.t434 C10_N_btm.t402 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4885 VDAC_P.t130 C10_P_btm.t428 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4886 VDD.t112 a_n2293_46508.t6 a_22031_44350# VDD.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4887 VDAC_N.t1650 C9_N_btm.t229 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4888 VDAC_P.t1658 C10_P_btm.t427 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4889 VDD.t2451 VSS.t3551 VDD.t2450 VDD.t2449 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X4890 VDAC_P.t842 C10_P_btm.t426 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4891 VDD.t614 a_13273_44868.t12 a_15605_45438# VDD.t613 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4892 VDAC_P.t1654 C8_P_btm.t103 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4893 VDAC_N.t838 C9_N_btm.t228 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4894 VSS.t2606 a_21303_42718# a_3222_30651.t0 VSS.t2605 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4895 VDAC_N.t1646 C10_N_btm.t401 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4896 VDD.t2448 VSS.t3556 VDD.t2447 VDD.t2446 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4897 a_571_43566# a_396_43640# a_750_43628# VSS.t2120 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X4898 VDAC_P.t434 C7_P_btm.t68 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4899 SMPL_ON_N.t3 a_21789_35634# VSS.t2663 VSS.t2662 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4900 COMP_N.t6 a_1239_39043# VDD.t1728 VDD.t1727 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4901 VDAC_P.t1650 C10_P_btm.t425 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4902 a_12101_44048# a_11883_43806# VDD.t723 VDD.t722 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4903 VDAC_N.t230 C10_N_btm.t400 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4904 C9_P_btm.t12 a_n2467_30659.t11 VREF.t18 VDD.t584 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4905 VDAC_P.t838 C10_P_btm.t424 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4906 VDAC_N.t1642 C9_N_btm.t227 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4907 VDD.t2445 VSS.t3626 VDD.t2444 VDD.t2443 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4908 VDAC_N.t834 C10_N_btm.t399 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4909 VSS.t976 a_5784_44364# a_5536_44324# VSS.t975 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4910 VDAC_N.t1638 VSS.t3325 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4911 a_8798_45758# a_1412_46794.t2 a_9048_45758# VSS.t148 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4912 VDAC_P.t1646 VSS.t3392 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4913 VDD.t2168 a_11599_42883# a_9096_45276.t1 VDD.t2167 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4914 VDAC_P.t230 C10_P_btm.t423 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4915 VDAC_N.t430 VSS.t3306 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4916 a_10905_43236# a_10687_43640# VDD.t2113 VDD.t2112 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4917 VSS.t186 a_135_43540.t42 a_645_43806# VSS.t185 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4918 VSS.t1580 a_4061_47044# a_4091_47070# VSS.t1579 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4919 VDAC_P.t1642 C10_P_btm.t422 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4920 VDAC_P.t834 C10_P_btm.t421 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4921 a_5916_43806# a_4835_43806# a_5569_44048# VDD.t948 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4922 VSS.t896 a_5663_42718# a_5840_42718.t0 VSS.t895 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4923 VREF.t53 a_n4515_30659.t4 C10_P_btm.t1056 VDD.t2990 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4924 a_5953_45982# a_5918_46234# a_5715_45956# VSS.t995 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X4925 VSS.t3445 VDD.t3207 VSS.t3444 VSS.t3042 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4926 VDAC_P.t1638 C10_P_btm.t419 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4927 a_927_42692.t0 a_4527_43566# VSS.t2209 VSS.t2208 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4928 a_11979_43806# a_11533_43806# a_11883_43806# VSS.t1531 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4929 a_2959_43806# a_2609_43806# a_2864_43806# VDD.t1160 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4930 VDAC_P.t430 C10_P_btm.t418 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4931 a_1597_45982# a_1431_45982# VDD.t689 VDD.t688 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4932 VSS.t2661 a_21789_35634# SMPL_ON_N.t2 VSS.t2660 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4933 VDD.t1239 a_12623_43780# a_10259_42870.t7 VDD.t1238 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X4934 VDAC_N.t1634 C8_N_btm.t257 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4935 VDAC_N.t830 C10_N_btm.t398 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4936 VDAC_P.t1634 C8_P_btm.t269 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4937 VDAC_N.t1630 C10_N_btm.t397 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4938 VDAC_P.t830 C10_P_btm.t417 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4939 VDAC_P.t1630 C10_P_btm.t416 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4940 a_4527_46830# a_4352_46904# a_4706_46892# VSS.t1080 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X4941 VDAC_N.t78 C10_N_btm.t396 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4942 VDAC_N.t1626 C8_N_btm.t98 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4943 a_n2109_47596.t1 a_19520_46500# VSS.t2105 VSS.t2104 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4944 VDAC_P.t78 C9_P_btm.t206 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4945 a_21197_42718# a_21027_42718# VDD.t625 VDD.t624 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4946 VDAC_P.t1626 C9_P_btm.t205 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4947 VSS.t2694 a_22223_47070# a_20647_31459.t0 VSS.t1138 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4948 VSS.t2637 a_22959_46534# a_20892_30659.t0 VSS.t1201 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4949 a_17951_44868# a_12127_46744# VSS.t1108 VSS.t1107 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X4950 a_10595_46904# a_10079_46532# a_10500_46892# VSS.t2254 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4951 a_18247_44172# a_8727_47222.t6 VDD.t75 VDD.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X4952 a_1302_43806# a_135_43540.t30 VSS.t174 VSS.t173 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X4953 VDD.t2436 VSS.t3693 VDD.t2435 VDD.t2434 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X4954 VDAC_N.t826 C9_N_btm.t226 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4955 a_10687_43640# a_10171_43268# a_10592_43628# VSS.t2181 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4956 VDAC_N.t1622 C10_N_btm.t395 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4957 VDAC_N.t426 C7_N_btm.t128 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4958 VSS.t252 a_18314_32299.t7 C10_N_btm.t3 VSS.t251 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4959 VDD.t347 a_1334_43494.t25 a_2157_43262# VDD.t346 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4960 VDD.t455 a_7754_40130.t12 VDD.t454 VDD.t453 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.5
X4961 VDAC_N.t1618 C10_N_btm.t393 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4962 VDAC_P.t826 C10_P_btm.t415 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4963 VDAC_P.t1622 C10_P_btm.t414 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4964 VDAC_P.t426 C10_P_btm.t413 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4965 VDAC_N.t822 C10_N_btm.t392 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4966 VDAC_P.t1618 C9_P_btm.t204 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4967 VCM.t16 a_3990_30651.t18 C10_P_btm.t5 VSS.t291 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4968 VDAC_P.t822 C9_P_btm.t203 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4969 VSS.t2486 VSS.t2487 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4970 VDAC_P.t1614 C10_P_btm.t411 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4971 VSS.t2478 VSS.t2479 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4972 VDAC_N.t1614 C10_N_btm.t391 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4973 VDAC_P.t226 C7_P_btm.t63 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4974 VDAC_N.t226 C10_N_btm.t390 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4975 VDD.t2800 a_15008_42692# a_5142_30651.t2 VDD.t2799 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4976 VDAC_P.t1610 C10_P_btm.t410 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4977 VDAC_N.t1610 C10_N_btm.t389 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4978 a_16291_46758# a_16555_46616# VSS.t1188 VSS.t1187 sky130_fd_pr__nfet_01v8 ad=0.05985 pd=0.705 as=0.0567 ps=0.69 w=0.42 l=0.15
X4979 VDAC_N.t818 C8_N_btm.t255 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4980 VDAC_P.t818 C9_P_btm.t202 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4981 VDAC_N.t1606 C9_N_btm.t225 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4982 VDAC_P.t1606 C10_P_btm.t409 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4983 VDAC_P.t422 C10_P_btm.t408 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4984 VSS.t2458 VSS.t2459 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4985 VDAC_P.t1602 C10_P_btm.t407 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4986 VDAC_N.t422 C9_N_btm.t224 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4987 VDAC_N.t1602 C7_N_btm.t58 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4988 VDAC_P.t814 C8_P_btm.t99 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4989 VDAC_P.t1598 C9_P_btm.t201 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4990 VDAC_P.t126 C9_P_btm.t200 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4991 VDAC_N.t814 C10_N_btm.t1053 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4992 VDD.t593 a_13273_44868.t20 a_15091_44440# VDD.t592 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4993 VDAC_N.t1598 C10_N_btm.t1052 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4994 VSS.t1622 a_1123_43780# a_1057_43806# VSS.t1621 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4995 a_9863_47874# a_10199_47846.t3 VDD.t3094 VDD.t3093 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X4996 a_15251_47320# a_15221_47044# a_15155_47320# VDD.t1877 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X4997 VSS.t2178 a_2216_46758# a_2167_46526# VSS.t2177 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4998 VDAC_P.t1594 C10_P_btm.t406 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X4999 VDAC_N.t126 C9_N_btm.t223 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5000 VDAC_P.t810 C5_P_btm.t32 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5001 a_13023_44716# a_12651_44576.t8 VDD.t2957 VDD.t2956 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X5002 a_134_42718.t1 a_104_42692# VSS.t934 VSS.t933 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X5003 VDAC_P.t1590 C10_P_btm.t405 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5004 a_4700_46134# a_4908_45956# a_4842_45982# VSS.t1788 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5005 a_2617_45144# a_2587_44868.t9 VDD.t229 VDD.t228 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X5006 VDAC_P.t418 C10_P_btm.t404 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5007 VDAC_N.t1594 C10_N_btm.t1049 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5008 a_9547_46565# a_9517_46539# a_9475_46565# VDD.t1925 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X5009 VDAC_N.t810 C10_N_btm.t387 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5010 VDAC_P.t1586 C10_P_btm.t403 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5011 VDAC_P.t806 C10_P_btm.t402 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5012 VDAC_N.t1590 C9_N_btm.t222 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5013 VDD.t435 a_7754_40130.t1 a_7754_40130.t2 VDD.t434 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X5014 a_21788_30659.t2 a_22223_47622# VDD.t969 VDD.t968 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5015 a_8897_44716# a_8862_44482# a_8659_44324# VSS.t2644 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X5016 VSS.t479 a_13248_45956.t10 a_15139_47730# VSS.t478 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X5017 VDAC_N.t418 C10_N_btm.t1047 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5018 VDD.t1824 a_18971_44654# a_15730_45670.t7 VDD.t1823 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X5019 a_6573_44716# a_6485_44582.t24 a_6491_44716# VSS.t2922 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X5020 VSS.t1481 a_3699_43780# a_3633_43806# VSS.t1480 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X5021 a_15589_44350# a_13715_43780# a_15443_44582# VDD.t1197 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X5022 VDAC_P.t1582 C10_P_btm.t401 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5023 VDAC_P.t222 C10_P_btm.t400 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5024 VDAC_N.t1586 C10_N_btm.t1045 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5025 VDAC_N.t806 VSS.t3258 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5026 VDD.t2413 VSS.t3635 VDD.t2412 VDD.t2320 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5027 VDAC_P.t1578 C9_P_btm.t199 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5028 VDAC_N.t1582 C10_N_btm.t386 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5029 VDAC_N.t222 C9_N_btm.t221 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5030 VDAC_N.t1578 C10_N_btm.t1043 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5031 VDAC_N.t802 C8_N_btm.t254 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5032 VDAC_P.t802 C10_P_btm.t399 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5033 a_18530_47070# a_17927_46195# a_18361_47320# VDD.t1895 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X5034 a_n2661_44332# a_n1827_45412.t12 VSS.t361 VSS.t360 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5035 VDAC_N.t1574 C10_N_btm.t385 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5036 a_n2442_43806.t3 a_n2472_43780# VDD.t736 VDD.t735 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5037 VDAC_P.t1574 C8_P_btm.t100 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5038 VDAC_N.t414 C10_N_btm.t1041 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5039 VDAC_P.t414 C8_P_btm.t98 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5040 VDAC_N.t1570 C10_N_btm.t384 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5041 a_13827_46298# a_13151_45956# a_13654_46032# VDD.t1482 sky130_fd_pr__pfet_01v8_hvt ad=0.090125 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X5042 VSS.t1907 a_12436_44868# a_n1741_47596.t0 VSS.t1906 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X5043 VDAC_P.t1570 C10_P_btm.t398 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5044 VDAC_N.t798 C9_N_btm.t220 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5045 a_2866_45982# a_135_43540.t22 VSS.t2776 VSS.t2775 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X5046 VDAC_N.t1566 C9_N_btm.t219 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5047 VDAC_N.t34 C9_N_btm.t218 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5048 a_11550_45554# a_10259_42870.t18 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X5049 VSS.t2418 VSS.t2419 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5050 VDAC_P.t798 C5_P_btm.t31 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5051 a_11335_46830# a_10227_47214.t13 VDD.t287 VDD.t286 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5052 a_3328_44324# a_3179_44403# a_3624_44466# VDD.t621 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5053 VSS.t519 a_1203_42692.t9 a_3541_42718# VSS.t518 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5054 a_7839_47222# a_1412_46794.t3 a_8013_47098# VSS.t149 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X5055 a_11427_43566# a_10227_47214.t12 VDD.t285 VDD.t284 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5056 a_21020_30659.t0 a_22591_47070# VSS.t1742 VSS.t1741 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5057 VDD.t2048 a_n2497_47846.t6 a_4833_47320# VDD.t2047 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X5058 VDAC_P.t1566 C7_P_btm.t136 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5059 VDAC_N.t1562 C10_N_btm.t383 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5060 VDAC_N.t794 C9_N_btm.t217 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5061 VDAC_P.t34 C10_P_btm.t397 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5062 VDAC_P.t1562 C9_P_btm.t198 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5063 VDAC_N.t1558 C9_N_btm.t216 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5064 VDAC_P.t794 C10_P_btm.t396 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5065 VDAC_N.t410 C10_N_btm.t1039 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5066 a_1110_44172# a_33_43806# a_948_43806# VDD.t884 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5067 VDAC_N.t1554 C7_N_btm.t126 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5068 VDD.t510 a_1053_45123.t5 a_9863_43958# VDD.t509 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X5069 a_923_45804# a_n53_44363.t7 a_560_45670# VSS.t615 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X5070 a_3882_44324# a_3576_44364# VDD.t1090 VDD.t1089 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.17575 ps=1.395 w=0.42 l=0.15
X5071 VDAC_N.t790 C10_N_btm.t382 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5072 VSS.t2549 VSS.t2550 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5073 VDAC_N.t1550 C10_N_btm.t381 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5074 VDAC_N.t218 C10_N_btm.t380 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5075 a_7129_44894# a_5939_44894# a_7020_44894# VSS.t1608 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5076 VDAC_P.t1558 C10_P_btm.t395 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5077 VDAC_N.t1546 C10_N_btm.t379 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5078 a_518_44670# a_570_44324# a_n1459_43236.t5 VSS.t1653 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5079 VDAC_N.t786 C9_N_btm.t215 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5080 VDAC_N.t1542 C8_N_btm.t96 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5081 VDAC_P.t410 C10_P_btm.t394 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5082 VDAC_N.t406 C10_N_btm.t378 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5083 VREF.t36 a_22812_30659.t8 C10_N_btm.t22 VDD.t520 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5084 VDAC_N.t1538 C10_N_btm.t377 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5085 VDAC_P.t1554 C10_P_btm.t393 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5086 VDAC_P.t790 C8_P_btm.t97 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5087 VSS.t2124 a_15323_44894# a_1429_47222.t0 VSS.t2123 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5088 C6_P_btm.t72 a_5542_30651.t4 VCM.t50 VSS.t2897 sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X5089 VDAC_N.t782 C7_N_btm.t57 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5090 a_3633_43806# a_2443_43806# a_3524_43806# VSS.t2101 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5091 a_5626_46526# a_5419_47258# VDD.t1531 VDD.t1530 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.3125 ps=1.625 w=1 l=0.15
X5092 a_10333_42718# a_10259_42870.t22 a_9987_42968# VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5093 VDAC_N.t1534 C9_N_btm.t214 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5094 a_10150_47322# a_10428_47338# a_10384_47436# VDD.t2080 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X5095 VDAC_P.t1550 C4_P_btm.t8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5096 SMPL_ON_P.t0 a_n2038_35608# VSS.t2623 VSS.t2622 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5097 VDAC_P.t218 C6_P_btm.t52 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5098 VDAC_N.t122 C10_N_btm.t376 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5099 VDAC_P.t1546 C8_P_btm.t264 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5100 VSS.t2046 a_2351_47614# DATA[2].t0 VSS.t2045 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5101 a_4364_45982# a_4322_46134# a_4061_45956# VSS.t1816 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X5102 VDD.t848 a_16703_42718# a_4758_30651.t3 VDD.t847 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X5103 a_18401_43806# a_18357_44048# a_18235_43806# VSS.t796 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X5104 VDAC_N.t1530 C9_N_btm.t213 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5105 a_16101_43628# a_16057_43236# a_15935_43640# VSS.t1966 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X5106 VDAC_N.t778 C10_N_btm.t375 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5107 VDAC_P.t786 C10_P_btm.t392 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5108 VDD.t2934 a_n2103_44868.t10 a_n2293_44868# VDD.t2870 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5109 a_11415_45670# a_11687_45528# VSS.t1180 VSS.t1179 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5110 VDAC_P.t1542 C10_P_btm.t391 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5111 VDAC_N.t1526 C9_N_btm.t212 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5112 VDAC_N.t402 C10_N_btm.t183 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5113 VSS.t3730 C9_P_btm.t17 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5114 VDAC_P.t406 C10_P_btm.t390 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5115 VDD.t644 a_12427_42883# a_10844_44364# VDD.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5116 a_8912_37509.t14 VDAC_N.t1522 a_5700_37509.t8 VDD.t2243 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X5117 a_3553_42968# a_1847_45528.t22 VDD.t2892 VDD.t2891 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5118 VDAC_N.t774 C9_N_btm.t211 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5119 VDAC_N.t1518 C10_N_btm.t373 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5120 VDAC_P.t1538 C10_P_btm.t389 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5121 VDAC_N.t214 C9_N_btm.t210 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5122 VDAC_N.t1514 C10_N_btm.t372 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5123 VDAC_N.t770 C10_N_btm.t371 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5124 VDAC_P.t782 C10_P_btm.t388 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5125 VDAC_P.t1534 C10_P_btm.t1051 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5126 VDAC_P.t122 C9_P_btm.t533 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5127 VDAC_N.t1510 C8_N_btm.t95 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5128 VDAC_N.t398 C9_N_btm.t209 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5129 a_12427_42883# a_5542_30651.t8 VDD.t3068 VDD.t3067 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5130 VDAC_P.t1530 C10_P_btm.t1049 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5131 VSS.t3607 C8_N_btm.t265 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5132 VSS.t2930 a_n2103_43780.t13 a_22591_45982# VSS.t2929 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5133 VDAC_P.t778 C10_P_btm.t387 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5134 VDAC_P.t1526 C10_P_btm.t1047 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5135 a_5166_45804# a_135_43540.t9 VSS.t2815 VSS.t2814 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X5136 a_n2293_43244# a_n1827_44324.t4 VSS.t300 VSS.t299 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5137 a_14658_46526# a_13248_45956.t22 a_13457_46892# VDD.t411 sky130_fd_pr__pfet_01v8_hvt ad=0.092075 pd=0.99 as=0.1092 ps=1.36 w=0.42 l=0.15
X5138 VDD.t799 a_663_47874# DATA[1].t4 VDD.t798 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X5139 VDAC_N.t1506 C10_N_btm.t370 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5140 a_11730_34132.t1 a_18394_35068.t14 VSS.t198 VSS.t197 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X5141 VDAC_P.t402 C10_P_btm.t1045 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5142 VDAC_N.t766 C10_N_btm.t369 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5143 a_9943_45046# a_7557_43236.t8 VSS.t217 VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X5144 VDD.t1970 a_9947_47044# a_7208_47044# VDD.t1969 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X5145 VDAC_N.t1502 C6_N_btm.t49 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5146 VDAC_N.t74 C9_N_btm.t208 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5147 VCM.t26 a_5923_31099.t5 C4_N_btm.t3 VSS.t2082 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X5148 VDD.t106 a_927_42692.t24 a_1935_44874# VDD.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5149 VDAC_N.t1498 C9_N_btm.t207 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5150 VDAC_P.t1522 C7_P_btm.t133 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5151 VDD.t2313 VSS.t3652 VDD.t2312 VDD.t2311 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5152 VDAC_N.t762 C9_N_btm.t206 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5153 VDAC_P.t774 C9_P_btm.t531 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5154 VDD.t1094 a_3328_44324# a_n2293_45956.t3 VDD.t1093 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X5155 VDAC_N.t1494 C8_N_btm.t92 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5156 VDAC_N.t394 C10_N_btm.t368 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5157 VSS.t302 a_n1827_44324.t7 a_22223_46534# VSS.t301 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5158 VDAC_P.t1518 C10_P_btm.t386 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5159 VDAC_P.t214 C6_P_btm.t58 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5160 VSS.t3757 C4_N_btm.t22 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5161 VDD.t1523 a_n2840_43780# a_n2810_43806.t3 VDD.t881 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5162 a_10251_45454# a_17951_44868# VDD.t1290 VDD.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5163 VDAC_P.t1514 C8_P_btm.t263 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5164 VDAC_N.t1490 C10_N_btm.t367 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5165 VSS.t1749 a_16475_45412# a_16287_45744# VSS.t1748 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5166 VDAC_N.t758 C10_N_btm.t366 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5167 VDAC_P.t770 VSS.t3358 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5168 VDD.t1155 a_3177_44048# a_3067_44172# VDD.t1154 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X5169 VDAC_Ni.t8 a_3754_38470.t9 a_3726_37500# VSS.t2843 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X5170 a_927_42692.t1 a_4527_43566# VSS.t2203 VSS.t2202 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5171 a_13248_45956.t2 a_20159_47588# VDD.t1035 VDD.t1034 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5172 VDAC_P.t1510 C10_P_btm.t385 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5173 VDAC_P.t398 C10_P_btm.t1043 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5174 VDAC_N.t1486 C8_N_btm.t91 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5175 VDAC_N.t210 C9_N_btm.t205 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5176 VDAC_P.t1506 C9_P_btm.t197 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5177 VDAC_P.t766 C10_P_btm.t1042 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5178 a_19566_45670# a_19555_42718# VDD.t1005 VDD.t1004 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5179 VDAC_N.t1482 C10_N_btm.t365 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5180 VDAC_P.t1502 C10_P_btm.t1041 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5181 VDD.t2825 a_11455_44576.t24 a_11687_45528# VDD.t2824 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5182 VDAC_N.t754 C10_N_btm.t364 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5183 VDD.t1128 a_6325_45736# a_6355_45477# VDD.t1127 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5184 VDAC_N.t1478 C10_N_btm.t363 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5185 VDAC_P.t74 C10_P_btm.t384 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5186 VSS.t528 a_1203_42692.t12 a_8969_43582# VSS.t527 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5187 VSS.t2744 a_885_44868.t12 a_1304_44894# VSS.t2743 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X5188 VDAC_N.t390 C10_N_btm.t362 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5189 a_14219_47070# a_13248_45956.t12 VDD.t399 VDD.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5190 VSS.t2817 a_135_43540.t12 a_8005_46892# VSS.t2816 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5191 VSS.t3778 C10_N_btm.t1072 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5192 VSS.t1836 a_11692_46134# a_11248_47319# VSS.t1835 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X5193 VSS.t3496 VDD.t3225 VSS.t3495 VSS.t3494 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5194 VSS.t2333 VSS.t2334 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5195 VDAC_N.t1474 C10_N_btm.t360 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5196 VDD.t2042 a_1651_47044.t3 a_1597_47320# VDD.t2041 sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.135 ps=1.27 w=1 l=0.15
X5197 VDAC_P.t1498 C10_P_btm.t1039 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5198 VDAC_P.t762 C10_P_btm.t383 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5199 VDAC_N.t750 C10_N_btm.t359 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5200 VDD.t1130 a_11017_45736# a_11047_45477# VDD.t1129 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5201 a_13536_43780# a_13715_43780# VSS.t1265 VSS.t1264 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5202 a_18394_35068.t4 SMPL.t16 VSS.t2948 VSS.t2947 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5203 a_2709_43262# a_927_42692.t11 a_2627_43262# VDD.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5204 VDD.t1277 a_7839_47222# a_7760_45956# VDD.t1276 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X5205 VDAC_P.t1494 C8_P_btm.t261 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5206 VSS.t860 a_663_47874# DATA[1].t2 VSS.t859 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X5207 VDD.t2649 a_n2661_46508.t5 a_21755_44350# VDD.t2648 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5208 VDAC_N.t1470 C10_N_btm.t358 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5209 VDAC_Ni.t3 VSS.t3792 a_5088_37509.t2 VDD.t2372 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X5210 VDAC_P.t394 C10_P_btm.t1037 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5211 a_12379_44350# a_2755_43494.t21 a_12461_44350# VDD.t431 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5212 a_18766_43236# a_21197_42718# VDD.t1033 VDD.t1032 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5213 a_11183_44350# a_2755_43494.t9 a_11265_44670# VSS.t508 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X5214 VDAC_N.t118 C7_N_btm.t124 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5215 C9_P_btm.t537 a_4758_30651.t4 VCM.t56 VSS.t2986 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5216 VDAC_N.t1466 C7_N_btm.t112 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5217 VDAC_N.t746 C10_N_btm.t357 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5218 VDAC_P.t1490 C10_P_btm.t382 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5219 VDAC_N.t1462 C5_N_btm.t13 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5220 VDAC_P.t758 C8_P_btm.t94 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5221 VSS.t517 a_1736_39043.t6 a_1239_39043# VSS.t516 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5222 VDAC_N.t386 C9_N_btm.t204 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5223 a_n1459_43236.t1 a_927_42692.t21 VDD.t104 VDD.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5224 a_n2442_45438.t3 a_n2472_45412# VDD.t1378 VDD.t671 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5225 VDAC_N.t1458 C8_N_btm.t90 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5226 VSS.t930 a_22031_45438# a_22959_44358# VSS.t597 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5227 a_19191_43262# a_19003_43262# VSS.t1783 VSS.t1782 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1359 ps=1.1 w=0.65 l=0.15
X5228 VDAC_P.t1486 C7_P_btm.t55 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5229 VDAC_N.t742 VSS.t3255 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5230 VDAC_N.t1454 C10_N_btm.t356 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5231 VDD.t2773 a_n1920_47588# a_n1890_47614.t3 VDD.t2772 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5232 VDD.t1754 a_4527_46830# a_4322_46134# VDD.t1753 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5233 VDAC_P.t210 C9_P_btm.t196 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5234 DATA[3].t4 a_4651_47614# VDD.t1351 VDD.t1350 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X5235 a_1798_45144# a_1581_43806.t8 VDD.t2974 VDD.t2973 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X5236 a_2082_44670# a_2134_44324# a_n1735_43236.t5 VSS.t1787 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5237 VDAC_P.t1482 C10_P_btm.t381 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5238 VDAC_N.t206 C10_N_btm.t355 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5239 VSS.t3451 VDD.t3209 VSS.t3450 VSS.t3449 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5240 VDAC_P.t754 C10_P_btm.t380 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5241 VDAC_N.t1450 C9_N_btm.t203 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5242 a_13524_46832.t1 a_18135_47588# VSS.t1175 VSS.t1174 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5243 VDAC_N.t738 C10_N_btm.t354 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5244 a_11427_43566# a_11252_43640# a_11606_43628# VSS.t1892 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5245 VSS.t2778 a_135_43540.t24 a_93_46892# VSS.t2777 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5246 VDAC_P.t1478 C9_P_btm.t195 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5247 VDD.t1044 a_13561_44350# a_13819_44350# VDD.t1043 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5248 VDAC_N.t1446 C9_N_btm.t202 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5249 VDAC_N.t382 C10_N_btm.t353 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5250 a_13181_45982# a_13151_45956# a_12931_46348# VDD.t1481 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5251 VDAC_P.t390 C10_P_btm.t379 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5252 a_13373_46892# a_12651_44576.t10 VSS.t2861 VSS.t2860 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5253 VDAC_N.t1442 C9_N_btm.t201 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5254 VDAC_P.t1474 C9_P_btm.t525 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5255 VDAC_N.t734 C8_N_btm.t89 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5256 VSS.t3815 C6_P_btm.t1 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5257 a_8912_37509.t20 VDAC_N.t1438 a_5700_37509.t14 VDD.t2255 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X5258 VDAC_N.t50 VSS.t3288 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5259 VDAC_P.t750 C9_P_btm.t193 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5260 VDAC_P.t1470 VSS.t3333 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5261 VDAC_P.t118 C6_P_btm.t65 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5262 VDAC_P.t1466 C10_P_btm.t378 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5263 VDAC_P.t746 C4_P_btm.t7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5264 VDD.t1375 a_11143_47588# a_8727_47222.t2 VDD.t1374 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5265 a_8417_43806# a_7227_43806# a_8308_43806# VSS.t1008 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X5266 VDAC_P.t1462 C10_P_btm.t377 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5267 VDAC_N.t1434 C7_N_btm.t122 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5268 a_14647_43494# a_6104_45706.t8 a_14821_43600# VSS.t3009 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X5269 VDAC_P.t386 C10_P_btm.t376 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5270 VDAC_N.t730 C10_N_btm.t352 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5271 VDD.t2565 VSS.t3684 VDD.t2564 VDD.t2563 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5272 a_4908_45956# a_11335_46830# VDD.t866 VDD.t865 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X5273 a_18061_46892# a_17583_46500# VSS.t877 VSS.t876 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X5274 VDAC_P.t1458 C9_P_btm.t524 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5275 a_11183_44350# a_2755_43494.t10 a_11265_44350# VDD.t424 sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5276 VSS.t21 SMPL_ON_P.t8 a_n1605_47614# VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5277 a_13299_44716# a_10259_42870.t24 a_13193_44716# VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X5278 VDAC_N.t1430 C6_N_btm.t56 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5279 VDAC_N.t378 C9_N_btm.t200 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5280 VDAC_P.t742 C7_P_btm.t132 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5281 VDAC_P.t1454 C9_P_btm.t523 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5282 a_12931_44894# a_1581_43806.t21 VDD.t2915 VDD.t2914 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5283 VDAC_P.t206 C9_P_btm.t192 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5284 VDAC_P.t1450 C9_P_btm.t191 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5285 VDAC_P.t738 C10_P_btm.t375 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5286 VDAC_N.t1426 C10_N_btm.t351 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5287 VDAC_N.t726 C9_N_btm.t199 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5288 a_17671_42883# a_4758_30651.t12 VSS.t2994 VSS.t2993 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5289 VDD.t684 a_18133_47235# a_14950_43958# VDD.t683 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5290 VDAC_P.t1446 C8_P_btm.t259 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5291 VDAC_N.t1422 C9_N_btm.t198 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5292 VDAC_N.t202 VSS.t3296 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5293 a_5334_30651.t3 a_13023_42718# VDD.t1840 VDD.t1839 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5294 a_17881_44356# a_17715_44356# VSS.t701 VSS.t700 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5295 VDAC_P.t382 C10_P_btm.t89 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5296 VDAC_P.t1442 C8_P_btm.t92 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5297 VDAC_N.t1418 C10_N_btm.t350 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5298 VDAC_N.t722 C9_N_btm.t197 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5299 VDAC_P.t734 C10_P_btm.t373 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5300 VDD.t844 a_16513_42718# a_16703_42718# VDD.t843 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X5301 VDAC_P.t1438 C8_P_btm.t91 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5302 VDAC_P.t50 C10_P_btm.t372 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5303 a_6235_46124# a_4830_43958.t7 VDD.t198 VDD.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5304 VDAC_N.t1414 C8_N_btm.t88 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5305 VSS.t2138 a_2167_46526# a_2343_47070# VSS.t2137 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5306 a_13207_44894# a_1581_43806.t17 a_13101_44894# VSS.t2958 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X5307 VSS.t1844 a_22400_42718# a_22780_40517# VSS.t1843 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5308 VDAC_P.t1434 C10_P_btm.t371 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5309 VDAC_N.t374 C8_N_btm.t87 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5310 VDAC_P.t730 C8_P_btm.t90 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5311 VDAC_P.t1430 C3_P_btm.t11 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5312 a_22465_38541# a_22775_42718# VSS.t2688 VSS.t2687 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5313 a_15145_43262# a_11455_44576.t18 VDD.t2820 VDD.t2819 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5314 VDD.t2478 VSS.t3682 VDD.t2477 VDD.t2476 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5315 VSS.t82 a_8727_47222.t8 a_9343_43806# VSS.t81 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X5316 VDAC_P.t378 C10_P_btm.t370 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5317 VDAC_P.t1426 C6_P_btm.t57 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5318 a_5536_44324# a_4993_47044# VSS.t1425 VSS.t1424 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X5319 VDAC_P.t726 C10_P_btm.t369 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5320 a_9048_45758# a_1412_46794.t8 a_8798_45758# VSS.t150 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5321 VSS.t3177 VDD.t3161 VSS.t3176 VSS.t3175 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X5322 VDAC_P.t1422 C10_P_btm.t368 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5323 VDAC_N.t1410 C6_N_btm.t25 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5324 a_18139_43806# a_17789_43806# a_18044_43806# VDD.t1070 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5325 VDAC_P.t202 C10_P_btm.t367 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5326 VDAC_N.t718 C10_N_btm.t349 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5327 a_14382_46348# a_13524_46832.t5 a_13181_45982# VDD.t537 sky130_fd_pr__pfet_01v8_hvt ad=0.092075 pd=0.99 as=0.1092 ps=1.36 w=0.42 l=0.15
X5328 VDAC_N.t1406 C7_N_btm.t111 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5329 VDAC_N.t114 C9_N_btm.t521 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5330 a_19168_45758# a_13273_44868.t24 VSS.t646 VSS.t645 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5331 VDAC_P.t1418 C8_P_btm.t89 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5332 VDAC_N.t1402 C9_N_btm.t196 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5333 a_1204_46758# a_1412_46794.t10 a_1346_46892# VSS.t151 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5334 VDAC_N.t714 C10_N_btm.t348 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5335 a_n2442_44350.t3 a_n2472_44324# VDD.t988 VDD.t735 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5336 VDAC_P.t722 C9_P_btm.t190 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5337 VDAC_N.t1398 C10_N_btm.t347 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5338 VDAC_P.t1414 C9_P_btm.t519 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5339 VDAC_P.t374 C10_P_btm.t366 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5340 VDAC_P.t1410 C10_P_btm.t365 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5341 VSS.t542 a_1203_42692.t26 a_16513_42718# VSS.t541 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5342 C9_N_btm.t9 a_21788_30659.t8 VREF.t27 VDD.t2055 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5343 a_13266_45412# a_13144_47452.t5 VSS.t47 VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.11975 ps=1.045 w=0.42 l=0.15
X5344 VDAC_P.t718 C10_P_btm.t364 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5345 VDAC_P.t1406 C9_P_btm.t188 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5346 VDAC_N.t370 C9_N_btm.t519 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5347 a_10259_42870.t4 a_12623_43780# VDD.t1237 VDD.t1236 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5348 a_14635_44324# a_16074_45046# VDD.t1838 VDD.t1837 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5349 VDAC_P.t114 C10_P_btm.t363 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5350 a_n749_47846# a_n447_47044# VDD.t892 VDD.t891 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5351 VDAC_P.t1402 C9_P_btm.t187 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5352 VDAC_P.t714 C10_P_btm.t362 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5353 a_6563_45260# a_5939_44894# a_6455_44894# VDD.t1546 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5354 VDAC_N.t1394 C10_N_btm.t346 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5355 VDD.t2365 VSS.t3621 VDD.t2364 VDD.t2363 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5356 VDAC_N.t710 C10_N_btm.t345 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5357 VDD.t2067 a_n2840_45412# a_n2810_45438.t3 VDD.t1301 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5358 VSS.t2879 a_17564_32305.t4 C7_N_btm.t137 VSS.t2878 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X5359 VDD.t2886 a_1847_45528.t18 a_n2103_43780.t2 VDD.t2885 sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.135 ps=1.27 w=1 l=0.15
X5360 VDAC_N.t1390 C10_N_btm.t344 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5361 VDAC_N.t198 C7_N_btm.t82 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5362 a_15155_47070# a_15329_47044# VSS.t1119 VSS.t1118 sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X5363 a_20405_31459.t2 a_22959_45982# VDD.t1856 VDD.t1855 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5364 VDAC_N.t1386 C6_N_btm.t54 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5365 VDAC_N.t706 C9_N_btm.t195 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5366 VDAC_N.t1382 C10_N_btm.t343 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5367 VDAC_P.t1398 C10_P_btm.t361 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5368 VDAC_P.t370 C9_P_btm.t186 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5369 VDAC_N.t366 C8_N_btm.t86 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5370 VDAC_N.t1378 C9_N_btm.t517 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5371 VDAC_P.t1394 C5_P_btm.t30 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5372 DATA[3].t2 a_4651_47614# VSS.t1422 VSS.t1421 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5373 VDAC_P.t710 C8_P_btm.t88 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5374 VDAC_P.t1390 C9_P_btm.t185 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5375 a_18879_45956# a_18704_45982# a_19058_45982# VSS.t812 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5376 a_8912_37509.t12 VDAC_N.t702 a_5700_37509.t6 VDD.t2246 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X5377 VSS.t787 a_16651_46500# a_16291_46758# VSS.t786 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.05985 ps=0.705 w=0.42 l=0.15
X5378 VDAC_N.t1374 C9_N_btm.t194 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5379 VSS.t2361 VSS.t2362 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5380 a_4706_43628# a_135_43540.t40 VSS.t184 VSS.t183 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X5381 a_10730_45477# a_10684_45670# VDD.t695 VDD.t694 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X5382 VDAC_P.t198 C10_P_btm.t360 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5383 VDAC_P.t1386 C10_P_btm.t359 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5384 VDAC_N.t70 C0_N_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5385 VSS.t2718 a_11455_44576.t22 a_12747_47070# VSS.t2717 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X5386 a_8470_46526# a_7393_46532# a_8308_46904# VDD.t1212 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5387 a_17073_44056# a_15730_45670.t22 VDD.t500 VDD.t499 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X5388 VDAC_P.t706 C10_P_btm.t358 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5389 VDAC_N.t1370 C9_N_btm.t193 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5390 VDD.t1998 a_16287_45744# a_16111_45412# VDD.t1997 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X5391 VDAC_N.t698 C8_N_btm.t85 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5392 VDAC_N.t1366 C10_N_btm.t342 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5393 a_672_45982# a_n409_45982# a_325_46224# VDD.t980 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X5394 VDAC_N.t362 C8_N_btm.t84 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5395 VDAC_P.t1382 VSS.t3336 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5396 a_22465_38541# a_22775_42718# VDD.t2789 VDD.t2788 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5397 VDAC_N.t1362 C10_N_btm.t341 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5398 VDAC_P.t366 C9_P_btm.t184 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5399 VDAC_N.t694 C9_N_btm.t192 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5400 a_1663_45046# a_1935_44874# VSS.t1221 VSS.t1220 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5401 VDAC_P.t1378 C10_P_btm.t357 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5402 VDAC_N.t1358 C8_N_btm.t83 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5403 VSS.t2411 VSS.t2412 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5404 a_1115_47044# a_n99_45438.t4 VSS.t2091 VSS.t2090 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X5405 a_14601_32299.t1 a_22223_44358# VSS.t1523 VSS.t1522 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5406 VDAC_P.t702 C10_P_btm.t356 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5407 VDAC_P.t1374 C9_P_btm.t183 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5408 VSS.t3537 VDD.t3239 VSS.t3536 VSS.t3535 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5409 VDAC_N.t194 C10_N_btm.t340 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5410 a_14853_45438# a_14766_45596.t3 VDD.t2878 VDD.t2877 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5411 VDAC_N.t1354 C8_N_btm.t82 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5412 VDD.t1946 a_7016_46231# a_6954_46348# VDD.t1945 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X5413 VDAC_N.t690 C10_N_btm.t339 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5414 VDAC_P.t70 C9_P_btm.t182 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5415 a_2905_44894# a_2755_43494.t5 a_2471_45046# VSS.t505 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5416 a_1736_39587.t2 a_1343_38525.t9 VDD.t59 VDD.t58 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X5417 VSS.t3525 VDD.t3235 VSS.t3524 VSS.t3523 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5418 C5_N_btm.t0 EN_VIN_BSTR_N.t14 VIN_N.t2 VSS.t443 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X5419 a_636_42870# a_571_43566# VDD.t753 VDD.t752 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X5420 a_7552_46134# a_7760_45956# a_7694_45982# VSS.t2043 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5421 VDAC_N.t1350 C7_N_btm.t118 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5422 a_3692_46892# a_3575_46697# VDD.t1512 VDD.t1511 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X5423 VDAC_P.t1370 C10_P_btm.t355 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5424 VDAC_P.t698 C7_P_btm.t131 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5425 a_2301_45438# a_1847_45528.t24 VDD.t2896 VDD.t2895 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5426 a_n2442_45982.t1 a_n2472_45956# VSS.t1519 VSS.t1450 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X5427 VDD.t924 a_7000_47222# a_6951_47070# VDD.t923 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X5428 VDAC_N.t358 C6_N_btm.t23 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5429 VDAC_N.t1346 C8_N_btm.t81 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5430 a_3787_43640# a_3437_43268# a_3692_43628# VDD.t1611 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5431 VDAC_P.t1366 C10_P_btm.t354 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5432 VDAC_P.t362 C8_P_btm.t87 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5433 VDAC_N.t686 C10_N_btm.t338 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5434 VDAC_P.t1362 C5_P_btm.t29 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5435 VDAC_P.t694 C10_P_btm.t353 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5436 a_161_44648# a_n172_44582# VDD.t1009 VDD.t1008 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X5437 a_12683_43433# a_12379_44350# VSS.t1548 VSS.t1547 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X5438 VDAC_P.t1358 C8_P_btm.t86 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5439 VDAC_P.t194 C10_P_btm.t352 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5440 a_8391_47044# a_8727_47222.t18 VSS.t51 VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X5441 VSS.t2211 a_4527_43566# a_4461_43640# VSS.t2210 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X5442 a_361_45438# a_83_45776# VDD.t1927 VDD.t1926 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X5443 VDAC_P.t1354 C10_P_btm.t351 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5444 a_15121_46232# a_15328_46134# VDD.t1435 VDD.t1434 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X5445 VSS.t2134 a_8969_43582# a_9343_42718# VSS.t2133 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5446 VDAC_P.t690 C10_P_btm.t350 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5447 VSS.t53 a_8727_47222.t20 a_18401_43806# VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5448 VDAC_N.t1342 C9_N_btm.t513 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5449 VDAC_N.t110 C9_N_btm.t191 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5450 VDAC_N.t1338 C9_N_btm.t511 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5451 VDAC_N.t682 C10_N_btm.t337 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5452 VSS.t80 a_8727_47222.t5 a_16101_43628# VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5453 a_325_46224# a_107_45982# VSS.t692 VSS.t691 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X5454 VDD.t3032 a_n2103_43780.t11 a_22591_45982# VDD.t3031 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X5455 VDAC_N.t1334 C10_N_btm.t336 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5456 w_1375_34946.t7 a_n1123_35174.t5 w_1375_34946.t6 w_1375_34946.t5 sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X5457 a_15730_45670.t4 a_18971_44654# VDD.t1822 VDD.t1821 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5458 VDAC_P.t1350 C10_P_btm.t349 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5459 a_16074_45046# a_16291_44914# VSS.t1726 VSS.t1725 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X5460 VDAC_N.t354 C10_N_btm.t335 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5461 VDAC_P.t358 C9_P_btm.t181 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5462 VDD.t1903 a_18449_44324# a_18339_44350# VDD.t1902 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X5463 VDAC_P.t1346 C9_P_btm.t180 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5464 VSS.t855 a_2043_43958# a_n60_44618# VSS.t854 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X5465 a_6631_42883# a_5840_42718.t7 VSS.t2882 VSS.t2881 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5466 VDD.t734 a_n2472_43780# a_n2442_43806.t2 VDD.t733 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5467 VDD.t882 a_n2840_44324# a_n2810_44350.t3 VDD.t881 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5468 VSS.t2527 VSS.t2528 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5469 VDD.t2136 a_10467_47212# a_10428_47338# VDD.t2135 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5470 a_10588_45670# a_n53_44363.t6 a_10730_45477# VDD.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5471 a_n1741_47596.t1 a_12436_44868# VSS.t1909 VSS.t1908 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X5472 VDAC_N.t1330 C10_N_btm.t334 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5473 a_7842_44868# a_8192_44874# VSS.t2266 VSS.t2265 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5474 VDAC_N.t678 C5_N_btm.t12 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5475 VDAC_P.t686 C7_P_btm.t51 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5476 VDAC_N.t1326 C10_N_btm.t333 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5477 a_2134_44324# a_1736_43276# VDD.t1132 VDD.t1131 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.17575 ps=1.395 w=0.42 l=0.15
X5478 VDAC_N.t190 C10_N_btm.t332 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5479 VDD.t1542 a_5473_43582# a_5663_42718# VDD.t1541 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X5480 a_7029_44350.t0 a_6491_44716# VSS.t1565 VSS.t1564 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X5481 VDAC_P.t1342 VSS.t3334 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5482 VDD.t3013 a_6485_44582.t9 a_6665_43262# VDD.t3012 sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X5483 VDAC_N.t1322 C8_N_btm.t80 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5484 VDAC_P.t110 C8_P_btm.t85 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5485 VDD.t643 a_22469_41061# a_22705_38426# VDD.t642 sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X5486 a_16057_43236# a_15839_43640# VDD.t1647 VDD.t1646 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X5487 VDAC_P.t1338 C7_P_btm.t50 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5488 VDAC_P.t682 C10_P_btm.t348 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5489 VDAC_P.t1334 C9_P_btm.t179 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5490 VDAC_P.t354 C9_P_btm.t178 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5491 a_6091_43780# a_5916_43806# a_6270_43806# VSS.t1228 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5492 VREF.t13 a_n2467_30659.t6 C9_P_btm.t7 VDD.t579 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5493 VDAC_N.t674 C10_N_btm.t331 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5494 VDAC_P.t1330 C10_P_btm.t347 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5495 VSS.t2365 VSS.t2366 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5496 VDAC_N.t1318 C10_N_btm.t330 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5497 VDAC_N.t350 C10_N_btm.t329 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5498 VDAC_P.t678 C9_P_btm.t177 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5499 VDAC_P.t1326 C10_P_btm.t346 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5500 VDAC_N.t1314 C10_N_btm.t328 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5501 VSS.t1614 a_6951_47070# a_7311_47614# VSS.t1613 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5502 VSS.t2164 a_22399_44894# a_22959_43806# VSS.t991 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5503 VSS.t170 a_1847_45528.t12 a_1659_45528# VSS.t169 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5504 VDAC_N.t670 C9_N_btm.t509 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5505 VDAC_N.t1310 C10_N_btm.t327 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5506 a_12896_47044# a_12747_47070# a_13192_47320# VDD.t717 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5507 VDAC_P.t190 C9_P_btm.t176 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5508 VDAC_N.t38 C9_N_btm.t188 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5509 VDD.t1798 a_18103_46768# a_18064_46642# VDD.t1797 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5510 VDAC_N.t1306 C10_N_btm.t326 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5511 VDAC_N.t666 C10_N_btm.t325 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5512 VDAC_P.t1322 C10_P_btm.t345 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5513 VDAC_P.t674 C8_P_btm.t41 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5514 C10_P_btm.t1070 a_n4515_30659.t18 VREF.t67 VDD.t3004 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5515 VSS.t2820 RST_Z.t3 a_7754_39964# VSS.t1074 sky130_fd_pr__nfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.15
X5516 a_14259_44133# a_14077_44133# VDD.t780 VDD.t779 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X5517 VSS.t117 a_15163_45670.t8 a_15112_45798# VSS.t116 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X5518 C10_N_btm.t16 EN_VIN_BSTR_N.t11 VIN_N.t5 VSS.t440 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5519 a_5459_44172# a_5655_43780# VDD.t2199 VDD.t2198 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X5520 VDAC_N.t1302 C7_N_btm.t56 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5521 a_22123_44894# a_n2293_47044.t9 VSS.t526 VSS.t525 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5522 VDAC_P.t1318 C10_P_btm.t343 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5523 VDAC_N.t346 C7_N_btm.t52 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5524 VDAC_N.t1298 C10_N_btm.t324 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5525 VDAC_N.t662 C4_N_btm.t15 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5526 VDAC_P.t350 C8_P_btm.t83 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5527 VDAC_N.t1294 C8_N_btm.t79 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5528 a_20064_35138# VDD.t3189 EN_VIN_BSTR_N.t4 VSS.t3396 sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.9
X5529 VDD.t831 a_325_46224# a_215_46348# VDD.t830 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X5530 VDAC_P.t1314 C8_P_btm.t82 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5531 VDAC_N.t186 C9_N_btm.t507 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5532 a_4352_43640# a_3271_43268# a_4005_43236# VDD.t2072 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X5533 VDAC_P.t670 C10_P_btm.t342 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5534 VDAC_P.t1310 C10_P_btm.t341 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5535 VDAC_N.t1290 C10_N_btm.t323 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5536 VSS.t3243 VDD.t3184 VSS.t3242 VSS.t3241 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X5537 VDAC_P.t38 C10_P_btm.t340 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5538 VDAC_P.t1306 C10_P_btm.t339 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5539 VDAC_P.t666 C8_P_btm.t81 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5540 a_22812_30659.t2 a_22959_47622# VDD.t1706 VDD.t1138 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5541 a_8308_43806# a_7393_43806# a_7961_44048# VSS.t1597 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5542 a_5419_47258# a_6631_44582# VSS.t1511 VSS.t1510 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5543 VDD.t654 a_11183_42718# a_5542_30651.t3 VDD.t653 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X5544 VDAC_P.t1302 C10_P_btm.t338 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5545 VDAC_N.t658 C10_N_btm.t322 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5546 VDAC_P.t346 C10_P_btm.t337 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5547 VDAC_N.t1286 C10_N_btm.t321 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5548 VDD.t1168 a_7595_47614# DATA[5].t6 VDD.t1167 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X5549 VDD.t351 a_n690_43494.t7 a_3731_45444# VDD.t350 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5550 VDD.t1298 a_10251_45454# a_19003_43262# VDD.t1297 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5551 VSS.t1655 a_n2840_45956# a_n2810_45982.t1 VSS.t1654 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5552 VSS.t1007 a_14573_47070# a_14955_45982# VSS.t1006 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X5553 VCM.t55 a_2252_42718.t7 C1_N_btm.t6 VSS.t2831 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X5554 VDAC_N.t342 C9_N_btm.t186 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5555 VDAC_P.t1298 C10_P_btm.t336 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5556 VDD.t595 a_13273_44868.t22 a_19371_46579# VDD.t594 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X5557 a_1297_45221# a_636_42870# a_1083_45221# VDD.t762 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X5558 a_8483_46830# a_8308_46904# a_8662_46892# VSS.t894 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5559 a_10389_45438# a_10111_45776# VDD.t792 VDD.t791 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X5560 a_n2810_47070.t2 a_n2840_47044# VDD.t2092 VDD.t2091 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5561 a_n264_46892# a_n381_46697# VSS.t1304 VSS.t1303 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X5562 VDAC_N.t1282 C10_N_btm.t320 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5563 VSS.t1196 a_1736_43276# a_1488_43236# VSS.t1195 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5564 VDAC_P.t662 C4_P_btm.t13 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5565 VDAC_P.t1294 C9_P_btm.t175 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5566 VDD.t801 a_663_47874# DATA[1].t6 VDD.t800 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5567 VDAC_N.t654 C10_N_btm.t319 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5568 VDAC_P.t186 C10_P_btm.t335 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5569 a_n1459_43236.t2 a_636_42870# VDD.t757 VDD.t756 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5570 VSS.t775 a_4239_42883# a_1736_43276# VSS.t774 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5571 VDAC_P.t1290 C10_P_btm.t334 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5572 VDAC_P.t658 C9_P_btm.t174 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5573 VDAC_P.t1286 C10_P_btm.t333 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5574 VDAC_N.t1278 C8_N_btm.t78 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5575 VDD.t2285 VSS.t3637 VDD.t2284 VDD.t2283 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5576 VSS.t3709 C6_N_btm.t67 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5577 a_6322_46348# a_6196_46250# a_5918_46234# VSS.t1053 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X5578 a_2358_46892# a_885_44868.t20 VSS.t2750 VSS.t2749 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X5579 a_18970_45412# a_19566_45670# VSS.t1041 VSS.t1040 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.11975 ps=1.045 w=0.42 l=0.15
X5580 VSS.t2466 VSS.t2467 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5581 a_12386_45758# a_2424_46794.t3 a_12636_45758# VSS.t2849 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5582 VDAC_N.t106 VSS.t3291 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5583 VDD.t1984 a_4791_42883# a_3576_44364# VDD.t1983 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5584 VDAC_N.t1274 C7_N_btm.t53 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5585 VDD.t233 a_2587_44868.t12 a_2709_43262# VDD.t232 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5586 VDAC_N.t650 C10_N_btm.t318 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5587 VDAC_N.t1270 C10_N_btm.t317 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5588 VDD.t1538 a_22821_39429# a_22521_39947# VDD.t1537 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5589 VDAC_P.t342 C10_P_btm.t332 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5590 VDAC_N.t338 C9_N_btm.t185 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5591 VDAC_N.t1266 C9_N_btm.t184 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5592 VDAC_P.t1282 C10_P_btm.t331 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5593 a_n2293_45956.t2 a_3328_44324# VDD.t1092 VDD.t1091 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X5594 VDAC_P.t654 C8_P_btm.t80 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5595 VDAC_N.t646 C9_N_btm.t183 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5596 VDAC_P.t1278 C9_P_btm.t173 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5597 a_n1920_42692# a_n1741_42692# VDD.t2733 VDD.t2732 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5598 VDAC_P.t106 C10_P_btm.t330 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5599 VDAC_P.t1274 C10_P_btm.t329 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5600 C8_N_btm.t1 a_5142_30651.t9 VCM.t3 VSS.t125 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5601 VDAC_P.t650 C10_P_btm.t328 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5602 VDAC_N.t1262 C9_N_btm.t182 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5603 VDAC_P.t1270 C8_P_btm.t79 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5604 VSS.t2967 a_13878_32299.t4 C2_N_btm.t7 VSS.t298 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X5605 VDAC_N.t182 C10_N_btm.t316 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5606 VSS.t784 a_1633_46824# a_1567_46892# VSS.t783 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5607 VDD.t374 EN_VIN_BSTR_N.t19 w_11534_34010.t9 w_11534_34010.t8 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X5608 VSS.t2205 a_4527_43566# a_927_42692.t3 VSS.t2204 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5609 a_9137_44716# a_8659_44324# VSS.t1291 VSS.t1290 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X5610 VDAC_P.t338 C10_P_btm.t327 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5611 VDAC_N.t1258 C10_N_btm.t315 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5612 VSS.t414 a_n690_43494.t6 a_1431_45982# VSS.t413 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5613 a_16671_47320# a_16703_45982# VDD.t985 VDD.t984 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5614 VDAC_N.t642 C10_N_btm.t314 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5615 a_571_46830# a_396_46904# a_750_46892# VSS.t911 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5616 VSS.t410 a_1334_43494.t27 a_1659_44440# VSS.t409 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5617 VDAC_N.t1254 C8_N_btm.t77 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5618 VDAC_N.t334 VSS.t3302 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5619 VDAC_P.t1266 VSS.t3341 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5620 VDAC_P.t646 C6_P_btm.t63 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5621 C10_P_btm.t6 a_3990_30651.t20 VCM.t18 VSS.t293 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5622 a_1597_47320# a_n1435_47614.t3 a_1513_47320# VDD.t3071 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5623 VDAC_N.t1250 C10_N_btm.t313 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5624 VDAC_P.t1262 C10_P_btm.t326 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5625 VSS.t3044 VDD.t3116 VSS.t3043 VSS.t3042 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5626 VDAC_P.t182 C10_P_btm.t325 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5627 a_16872_45144# a_16824_45276# a_16788_45144# VDD.t1987 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5628 VDD.t552 a_13524_46832.t16 a_15328_46134# VDD.t402 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5629 a_22400_42718# a_22223_42718# VDD.t869 VDD.t667 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X5630 VDAC_N.t638 C10_N_btm.t312 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5631 C4_P_btm.t0 a_n2810_43262.t4 VSS.t147 VSS.t146 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X5632 VDAC_P.t1258 C10_P_btm.t324 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5633 VDAC_N.t1246 C10_N_btm.t311 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5634 a_n1920_47588# a_n1741_47596.t7 VSS.t321 VSS.t320 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X5635 VDAC_N.t66 C10_N_btm.t310 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5636 VDAC_N.t1242 C8_N_btm.t76 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5637 VDAC_P.t642 C10_P_btm.t323 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5638 VDAC_P.t1254 C10_P_btm.t322 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5639 VDAC_N.t634 C10_N_btm.t309 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5640 VDAC_P.t334 C8_P_btm.t78 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5641 VDAC_P.t1250 C10_P_btm.t321 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5642 VDAC_N.t1238 C9_N_btm.t181 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5643 VDAC_N.t330 C10_N_btm.t308 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5644 VDD.t1379 a_n2472_45412# a_n2442_45438.t2 VDD.t673 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5645 a_10730_45804# a_10684_45670# VSS.t765 VSS.t764 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X5646 VDAC_N.t1234 C8_N_btm.t75 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5647 VDAC_P.t638 C9_P_btm.t172 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5648 VDD.t821 a_17583_46500# a_16291_44914# VDD.t820 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X5649 VSS.t2084 START.t1 a_14587_47614# VSS.t2083 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5650 VDAC_P.t1246 C7_P_btm.t48 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5651 VDD.t1203 a_16670_44324# a_n2103_44868.t2 VDD.t1202 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5652 a_16211_43780# a_8727_47222.t12 VDD.t83 VDD.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X5653 VSS.t1269 a_16111_45412# a_15187_44868# VSS.t1268 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X5654 VDAC_N.t630 C9_N_btm.t180 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5655 a_9395_47044# a_9551_47203# VSS.t2030 VSS.t2029 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X5656 a_2645_46824# a_885_44868.t34 VDD.t2854 VDD.t2853 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X5657 VDD.t743 a_18704_45982# a_18879_45956# VDD.t742 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5658 VSS.t3559 C7_P_btm.t8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5659 VDAC_P.t66 C9_P_btm.t171 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5660 VDAC_N.t1230 C9_N_btm.t179 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5661 a_12657_46642# a_10114_45276.t3 a_12562_46642# VDD.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X5662 VDAC_P.t1242 C4_P_btm.t9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5663 a_12833_42718# a_1203_42692.t20 a_12845_42968# VDD.t482 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5664 VDAC_N.t178 C7_N_btm.t51 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5665 VDD.t902 a_9208_43494# a_9159_43262# VDD.t901 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X5666 a_7276_45670# a_6985_45438# a_7418_45804# VSS.t1709 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5667 VDAC_N.t1226 C10_N_btm.t307 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5668 VSS.t2724 a_11455_44576.t26 a_13207_46892# VSS.t2723 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5669 VSS.t3111 VDD.t3139 VSS.t3110 VSS.t3109 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5670 VDAC_P.t634 C10_P_btm.t320 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5671 VSS.t2327 VSS.t2328 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5672 VDAC_P.t1238 C10_P_btm.t319 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5673 VSS.t1312 a_12623_43780# a_10259_42870.t3 VSS.t1311 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5674 VSS.t1161 a_7981_45956# a_7915_45982# VSS.t1160 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X5675 a_n2293_46508.t3 a_7842_44868# VDD.t1472 VDD.t1471 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.315 ps=2.63 w=1 l=0.15
X5676 VDAC_N.t626 C10_N_btm.t306 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5677 VDAC_N.t1222 C9_N_btm.t178 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5678 VDAC_P.t330 C10_P_btm.t318 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5679 VDD.t2260 VSS.t3576 VDD.t2259 VDD.t2258 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X5680 a_3067_44172# a_2443_43806# a_2959_43806# VDD.t2062 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5681 VDAC_P.t1234 C9_P_btm.t170 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5682 VDAC_P.t630 C9_P_btm.t169 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5683 VDAC_P.t1230 C10_P_btm.t317 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5684 a_1203_42692.t7 a_1431_47070# VDD.t2192 VDD.t2191 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.4 ps=1.8 w=1 l=0.15
X5685 VDAC_N.t326 C10_N_btm.t305 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5686 VDAC_P.t178 C7_P_btm.t127 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5687 VDAC_P.t1226 C10_P_btm.t316 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5688 VDAC_N.t1218 C10_N_btm.t304 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5689 VDD.t2073 a_22959_43806# a_17564_32305.t2 VDD.t1062 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X5690 VDAC_P.t626 C10_P_btm.t315 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5691 VDD.t1439 a_6631_44582# a_7569_44466# VDD.t1438 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5692 a_161_44648# a_n172_44582# VSS.t1069 VSS.t1068 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X5693 VDAC_N.t622 C10_N_btm.t303 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5694 VDAC_N.t1214 C10_N_btm.t302 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5695 VSS.t2836 a_14601_32299.t5 C6_N_btm.t71 VSS.t2835 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X5696 VDAC_P.t1222 C10_P_btm.t314 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5697 VDAC_N.t102 C10_N_btm.t301 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5698 VDAC_P.t326 C10_P_btm.t313 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5699 VDAC_P.t1218 C10_P_btm.t312 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5700 VDD.t755 a_636_42870# a_594_42968# VDD.t754 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0567 ps=0.69 w=0.42 l=0.15
X5701 VDAC_N.t1210 C10_N_btm.t300 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5702 VSS.t412 a_n690_43494.t5 a_n409_45982# VSS.t411 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5703 VDAC_P.t622 C8_P_btm.t77 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5704 a_5613_43806# a_5569_44048# a_5447_43806# VSS.t914 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X5705 VDAC_P.t1214 C10_P_btm.t311 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5706 VDAC_N.t618 C7_N_btm.t50 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5707 VSS.t1433 a_14950_43958# a_17715_44356# VSS.t1432 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5708 VDAC_N.t1206 C10_N_btm.t299 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5709 VDAC_P.t102 C9_P_btm.t168 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5710 VDAC_N.t322 C10_N_btm.t298 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5711 VDAC_P.t1210 C10_P_btm.t151 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5712 a_n1551_44324.t0 a_7557_43236.t10 VDD.t212 VDD.t211 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5713 VDD.t476 a_1203_42692.t14 a_20283_43262# VDD.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5714 VDD.t210 a_7557_43236.t9 a_7493_43262# VDD.t209 sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X5715 a_14819_44582# a_15091_44440# a_15049_44466# VDD.t691 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X5716 VDAC_N.t1202 C10_N_btm.t297 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5717 a_n1522_42718.t3 a_n1552_42692# VDD.t2659 VDD.t2658 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X5718 a_18259_46500# a_18064_46642# a_18569_46892# VSS.t1842 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X5719 VSS.t2230 a_7195_44868# a_7129_44894# VSS.t2229 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X5720 VSS.t1368 a_10251_45454# a_16177_45982# VSS.t1367 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X5721 a_n1735_43236.t3 a_82_45670# VDD.t1630 VDD.t1629 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5722 VDAC_P.t618 C10_P_btm.t309 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5723 VDAC_N.t614 C8_N_btm.t74 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5724 VDD.t1508 a_10901_42718# a_11183_42718# VDD.t1507 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X5725 VDAC_P.t1206 C5_P_btm.t28 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5726 C9_P_btm.t6 a_n2467_30659.t5 VREF.t12 VDD.t578 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5727 VDAC_P.t322 C10_P_btm.t308 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5728 a_10554_47436# a_10428_47338# a_10150_47322# VSS.t2118 sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X5729 a_12436_44868# a_12287_44894# a_12732_45144# VDD.t785 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5730 a_4338_37500.t1 a_3754_38470.t10 VDAC_Pi.t0 VSS.t2844 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X5731 VSS.t3766 C9_P_btm.t16 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5732 a_4239_42883# a_2252_42718.t5 VDD.t3080 VDD.t3079 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5733 VSS.t3502 VDD.t3227 VSS.t3501 VSS.t3500 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5734 VDAC_N.t1198 C10_N_btm.t296 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5735 VDD.t39 a_9521_45982.t20 a_17623_45982# VDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5736 VDAC_P.t1202 C10_P_btm.t307 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5737 VDAC_P.t614 C10_P_btm.t306 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5738 VDD.t367 a_n690_43494.t20 a_n685_46532# VDD.t366 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5739 VDAC_N.t174 C9_N_btm.t177 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5740 VDAC_N.t1194 C10_N_btm.t295 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5741 VSS.t3017 VDD.t3107 VSS.t3016 VSS.t3015 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X5742 VDAC_N.t610 C9_N_btm.t176 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5743 VDAC_N.t1190 C10_N_btm.t143 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5744 VSS.t3038 VDD.t3114 VSS.t3037 VSS.t3036 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5745 a_11533_43806# a_11367_43806# VSS.t1675 VSS.t1674 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5746 VDAC_N.t318 C10_N_btm.t293 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5747 VDAC_N.t1186 C10_N_btm.t292 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5748 VDAC_P.t1198 C10_P_btm.t305 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5749 VDAC_N.t606 C10_N_btm.t291 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5750 VDAC_P.t174 C10_P_btm.t304 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5751 VDAC_N.t1182 C10_N_btm.t290 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5752 VDD.t1250 a_6126_46642# a_n2661_45956.t3 VDD.t1249 sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X5753 VDAC_P.t1194 C10_P_btm.t303 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5754 VDAC_N.t46 C9_N_btm.t175 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5755 VDAC_N.t1178 C10_N_btm.t289 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5756 VDD.t339 a_1334_43494.t16 a_n1735_43236.t1 VDD.t338 sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.135 ps=1.27 w=1 l=0.15
X5757 VDAC_P.t610 C9_P_btm.t167 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5758 VDAC_P.t1190 C10_P_btm.t302 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5759 VDAC_N.t602 C10_N_btm.t288 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5760 VDAC_P.t318 C10_P_btm.t301 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5761 VDAC_N.t1174 C7_N_btm.t49 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5762 VDD.t989 a_n2472_44324# a_n2442_44350.t2 VDD.t733 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5763 VDAC_N.t314 C10_N_btm.t287 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5764 VDAC_P.t1186 C8_P_btm.t76 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5765 VDD.t2989 a_15549_47044.t11 a_18361_47320# VDD.t2988 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5766 a_14954_44466# a_12651_44576.t9 VDD.t2959 VDD.t2958 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X5767 VDAC_N.t1170 C7_N_btm.t125 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5768 VDAC_P.t606 C10_P_btm.t300 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5769 VSS.t469 a_n237_45454.t6 a_169_45776# VSS.t468 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X5770 VSS.t2956 a_1581_43806.t15 a_13572_46032# VSS.t2955 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X5771 VDAC_N.t598 C9_N_btm.t174 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5772 VSS.t3608 C0_P_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5773 VSS.t499 a_n237_45454.t16 a_3800_45982# VSS.t498 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5774 VDAC_P.t1182 C9_P_btm.t166 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5775 VDAC_N.t1166 C8_N_btm.t73 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5776 VDAC_P.t46 C5_P_btm.t27 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5777 VSS.t2822 RST_Z.t4 a_8530_39574# VSS.t2821 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5778 a_8005_46892# a_7961_46500# a_7839_46904# VSS.t1300 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X5779 VDAC_P.t1178 C7_P_btm.t125 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5780 a_16102_47044# a_15871_47614# VSS.t1335 VSS.t1334 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X5781 VDAC_N.t170 VSS.t3295 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5782 a_7743_43806# a_7393_43806# a_7648_43806# VDD.t1534 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5783 a_8912_37509.t32 VDAC_P.t602 a_5088_37509.t14 VDD.t2240 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X5784 a_n1085_47874# a_n749_47846# VDD.t896 VDD.t895 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X5785 a_10691_46904# a_10245_46532# a_10595_46904# VSS.t1983 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5786 VDAC_P.t1174 C10_P_btm.t299 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5787 VDAC_N.t1162 C9_N_btm.t173 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5788 VDAC_P.t314 C9_P_btm.t165 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5789 VSS.t2748 a_885_44868.t18 a_3470_45982# VSS.t2747 sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X5790 a_10588_45670# a_10389_45438# a_10730_45804# VSS.t853 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X5791 VDAC_P.t1170 C10_P_btm.t298 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5792 a_10783_43640# a_10337_43268# a_10687_43640# VSS.t1989 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5793 VDAC_N.t594 C9_N_btm.t172 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5794 VSS.t3072 VDD.t3126 VSS.t3071 VSS.t3070 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X5795 VDAC_P.t598 C9_P_btm.t164 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5796 VDAC_N.t1158 C7_N_btm.t47 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5797 VSS.t2884 a_12651_44576.t24 a_16427_44894# VSS.t2883 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X5798 VDAC_N.t310 C10_N_btm.t286 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5799 VSS.t1328 a_2075_42718# a_2252_42718.t1 VSS.t1327 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5800 VDD.t922 a_3320_46134# a_2535_45670# VDD.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X5801 VSS.t2405 VSS.t2406 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5802 VDAC_N.t1154 C10_N_btm.t285 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5803 VDD.t418 a_n237_45454.t17 a_6707_45776# VDD.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X5804 VDAC_P.t1166 C10_P_btm.t297 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5805 a_19679_31459.t0 a_22959_45446# VSS.t1354 VSS.t1353 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5806 VDD.t161 a_1412_46794.t5 a_n1827_44868.t1 VDD.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5807 VSS.t3240 VDD.t3183 VSS.t3239 VSS.t3238 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X5808 VDAC_P.t170 C10_P_btm.t296 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5809 VDAC_N.t590 C8_N_btm.t72 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5810 VDAC_N.t1150 C10_N_btm.t284 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5811 VDAC_N.t98 C9_N_btm.t171 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5812 a_10596_44324# a_10447_44403# a_10892_44466# VDD.t696 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5813 VDD.t549 a_13524_46832.t14 a_16921_46364# VDD.t548 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5814 VDAC_P.t1162 C6_P_btm.t61 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5815 VDAC_P.t594 C10_P_btm.t295 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5816 a_8379_46134# a_8651_45962# VSS.t1316 VSS.t1315 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5817 a_885_44868.t10 a_4322_46134# VDD.t1776 VDD.t1775 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5818 VSS.t1917 a_7754_38470# VSS.t1916 VSS.t1915 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X5819 VSS.t2446 VSS.t2447 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5820 VDAC_N.t1146 C7_N_btm.t123 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5821 a_3754_38470.t2 a_7754_38470# VSS.t693 sky130_fd_pr__res_high_po_0p35 l=18
X5822 VDAC_P.t1158 C10_P_btm.t294 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5823 VDD.t2316 VSS.t3661 VDD.t2315 VDD.t2314 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5824 VDD.t1016 a_11059_45956# a_11046_46348# VDD.t1015 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5825 VDAC_N.t586 C8_N_btm.t71 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5826 VDAC_P.t310 C8_P_btm.t75 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5827 VSS.t1378 a_14647_43494# a_14301_44035# VSS.t1377 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X5828 VDAC_P.t1154 C3_P_btm.t6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5829 VDAC_N.t1142 C9_N_btm.t170 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5830 VDAC_P.t590 C8_P_btm.t74 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5831 a_5839_47070# a_5749_47222# VSS.t2066 VSS.t2065 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5832 VDAC_P.t1150 VSS.t3344 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5833 a_6665_43262# a_2587_44868.t26 VDD.t247 VDD.t246 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X5834 VDAC_N.t306 C10_N_btm.t283 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5835 a_14819_44582# a_12651_44576.t18 VSS.t2867 VSS.t2866 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X5836 VSS.t1518 a_n2472_45956# a_n2442_45982.t0 VSS.t1448 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5837 EN_COMP.t1 a_n2288_42692# VSS.t771 VSS.t770 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X5838 a_2579_46892# a_82_45670# a_2216_46758# VSS.t1686 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X5839 VDD.t2166 a_n1920_42692# a_n1890_42718.t3 VDD.t2165 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5840 VDAC_N.t1138 C9_N_btm.t169 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5841 a_15567_43806# a_15121_43806# a_15471_43806# VSS.t917 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X5842 VDAC_P.t98 C10_P_btm.t293 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5843 VDAC_P.t1146 C10_P_btm.t292 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5844 VDAC_N.t582 C10_N_btm.t282 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5845 VSS.t1391 a_n1586_35608# a_n2038_35608# VSS.t1390 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5846 VDAC_N.t1134 C10_N_btm.t281 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5847 VDAC_N.t166 C9_N_btm.t168 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5848 VSS.t3117 VDD.t3141 VSS.t3116 VSS.t3115 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X5849 VDAC_P.t586 C8_P_btm.t73 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5850 VDAC_P.t1142 C10_P_btm.t291 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5851 VDAC_P.t306 C9_P_btm.t163 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5852 VDAC_P.t1138 C10_P_btm.t290 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5853 a_16670_44324# a_16824_45276# VSS.t2036 VSS.t2035 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.11975 ps=1.045 w=0.42 l=0.15
X5854 VSS.t3441 VDD.t3205 VSS.t3440 VSS.t3439 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X5855 VSS.t3810 C9_N_btm.t533 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5856 a_11533_43806# a_11367_43806# VDD.t1615 VDD.t1614 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5857 a_5918_46234# a_6235_46124# a_6193_45982# VSS.t2271 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X5858 a_4758_30651.t0 a_16703_42718# VSS.t902 VSS.t901 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5859 VDD.t1289 a_17951_44868# a_10251_45454# VDD.t1288 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5860 VDAC_P.t582 C10_P_btm.t289 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5861 VDD.t2457 VSS.t3687 VDD.t2456 VDD.t2455 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X5862 VDD.t574 a_10227_47214.t42 a_17583_46500# VDD.t573 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X5863 VDAC_N.t1130 C9_N_btm.t166 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5864 VDD.t1353 a_4993_47044# a_6280_46642# VDD.t1352 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5865 VDAC_N.t578 C9_N_btm.t165 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5866 VDAC_P.t1134 C9_P_btm.t162 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5867 VDAC_P.t166 C10_P_btm.t288 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5868 VDAC_N.t1126 C8_N_btm.t70 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5869 VDAC_N.t302 C9_N_btm.t164 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5870 VDAC_P.t1130 C9_P_btm.t161 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5871 VSS.t3419 VDD.t3197 VSS.t3418 VSS.t3417 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X5872 a_14470_46526# a_13248_45956.t16 VDD.t405 VDD.t404 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5873 VDD.t1680 a_16291_44914# a_12127_46744# VDD.t1679 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X5874 VDD.t1285 a_22959_45446# a_19679_31459.t2 VDD.t1284 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X5875 VSS.t2295 VSS.t2296 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5876 VDAC_N.t1122 C7_N_btm.t45 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5877 VDAC_N.t574 C10_N_btm.t280 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5878 VDAC_P.t578 C10_P_btm.t287 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5879 VDAC_P.t1126 C9_P_btm.t160 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5880 VDAC_N.t1118 C5_N_btm.t11 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5881 VDAC_N.t62 C9_N_btm.t163 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5882 VDAC_N.t1114 C10_N_btm.t279 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5883 VDAC_P.t302 C7_P_btm.t45 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5884 a_22031_45438# a_n2661_47044.t8 VDD.t3064 VDD.t3063 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5885 VDAC_N.t570 C9_N_btm.t162 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5886 a_n1552_42692# a_n1429_43262# VDD.t898 VDD.t897 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5887 VSS.t538 a_1203_42692.t24 a_283_42692# VSS.t537 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5888 VDAC_N.t1110 C8_N_btm.t69 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5889 VDAC_P.t1122 C9_P_btm.t159 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5890 VDAC_P.t574 C8_P_btm.t72 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5891 VSS.t2952 SMPL.t20 a_18394_35068.t7 VSS.t2951 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5892 VSS.t2509 VSS.t2510 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5893 VDAC_P.t1118 C6_P_btm.t24 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5894 a_18447_44894# a_15730_45670.t10 VSS.t565 VSS.t564 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X5895 VDAC_P.t62 C9_P_btm.t157 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5896 VSS.t2301 VSS.t2302 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5897 VDAC_P.t1114 C8_P_btm.t71 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5898 C3_P_btm.t12 a_5840_42718.t6 VCM.t47 VSS.t126 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X5899 VSS.t962 a_8483_43780# a_8417_43806# VSS.t961 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X5900 VDAC_N.t298 C10_N_btm.t278 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5901 a_8308_43806# a_7227_43806# a_7961_44048# VDD.t950 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X5902 VDAC_N.t1106 C10_N_btm.t277 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5903 VDAC_P.t570 VSS.t3361 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5904 VSS.t994 a_8379_46134# a_7648_46134# VSS.t993 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X5905 VDAC_N.t566 C10_N_btm.t276 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5906 VDD.t2223 a_20383_42718# a_6974_31099.t2 VDD.t2222 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X5907 a_7393_46532# a_7227_46532# VDD.t1209 VDD.t1208 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X5908 VDAC_N.t1102 C8_N_btm.t68 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5909 VSS.t631 a_10227_47214.t38 a_13157_43628# VSS.t630 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X5910 VDAC_P.t1110 C10_P_btm.t286 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5911 VDAC_P.t298 C10_P_btm.t285 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5912 VDAC_P.t1106 C9_P_btm.t156 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5913 VDAC_N.t162 C10_N_btm.t275 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5914 VDAC_N.t1098 C10_N_btm.t274 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5915 VDAC_P.t566 C10_P_btm.t284 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5916 VDAC_N.t562 C10_N_btm.t273 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5917 VSS.t754 a_18133_47235# a_14950_43958# VSS.t753 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5918 VSS.t2367 VSS.t2368 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5919 a_10951_45804# a_n53_44363.t5 a_10588_45670# VSS.t614 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X5920 VDD.t1085 a_1115_47044# a_n53_44363.t2 VDD.t1084 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X5921 VDAC_P.t1102 C10_P_btm.t283 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5922 a_4833_47320# a_4993_47044# VDD.t1357 VDD.t1356 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5923 VDAC_N.t1094 C7_N_btm.t121 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5924 a_17738_32299.t0 a_22959_44358# VSS.t1125 VSS.t1124 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5925 VDD.t392 a_13248_45956.t5 a_13151_45956# VDD.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.1083 ps=1.36 w=0.42 l=0.15
X5926 VDAC_N.t294 C9_N_btm.t161 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5927 VDD.t1816 a_22733_47833# a_15163_45670.t1 VDD.t1815 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X5928 VDAC_P.t162 C2_P_btm.t7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5929 VDAC_P.t1098 C9_P_btm.t155 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5930 VSS.t3081 VDD.t3129 VSS.t3080 VSS.t3079 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X5931 a_21908_43236# a_22087_43244# VDD.t1279 VDD.t1278 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5932 VREF.t34 a_22812_30659.t16 C10_N_btm.t30 VDD.t528 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X5933 VSS.t69 COMP_P.t10 a_n1237_42718# VSS.t68 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5934 VDAC_N.t1090 C10_N_btm.t272 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5935 VDAC_N.t558 C7_N_btm.t43 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5936 C2_P_btm.t3 a_n2074_43262.t4 VSS.t2085 VSS.t297 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X5937 VDAC_N.t1086 C4_N_btm.t8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5938 VDAC_N.t94 C8_N_btm.t67 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5939 VDAC_N.t1082 C9_N_btm.t160 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5940 VDAC_P.t562 C8_P_btm.t70 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5941 VDAC_N.t1080 C9_N_btm.t159 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5942 VDAC_P.t1094 C8_P_btm.t69 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5943 VDAC_N.t2128 C9_N_btm.t158 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5944 VDD.t1862 a_5847_47614# DATA[4].t6 VDD.t1861 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X5945 VDAC_N.t552 C10_N_btm.t271 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5946 VDAC_P.t294 C9_P_btm.t154 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5947 VDAC_N.t2120 C10_N_btm.t270 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5948 VDAC_P.t1090 C9_P_btm.t153 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5949 a_n2840_44324# a_n2661_44332# VDD.t2137 VDD.t2122 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X5950 VDAC_P.t558 C10_P_btm.t282 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5951 VDAC_N.t1072 C10_N_btm.t269 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5952 VSS.t2791 a_n2103_45412.t11 a_22959_47622# VSS.t2790 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5953 VDAC_P.t1086 C10_P_btm.t281 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5954 VDAC_N.t2112 C8_N_btm.t66 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5955 VSS.t1602 a_11507_47833# a_11299_47832# VSS.t1601 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5956 VDAC_N.t288 C9_N_btm.t157 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5957 VDAC_P.t94 C9_P_btm.t152 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5958 VDAC_P.t1082 C9_P_btm.t151 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5959 VSS.t2701 a_15831_42883# a_13144_47452.t0 VSS.t2700 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X5960 a_7557_43236.t2 a_11427_43566# VSS.t1171 VSS.t1170 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5961 VDD.t2375 VSS.t3686 VDD.t2374 VDD.t2373 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5962 VDAC_N.t2104 C9_N_btm.t156 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5963 VDAC_N.t1064 C9_N_btm.t155 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5964 a_18339_44350# a_17715_44356# a_18231_44728# VDD.t632 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X5965 VDD.t2378 VSS.t3564 VDD.t2377 VDD.t2376 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X5966 VDAC_P.t1080 C10_P_btm.t280 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5967 VDD.t2387 VSS.t3688 VDD.t2386 VDD.t2385 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X5968 VDAC_N.t2096 C9_N_btm.t154 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5969 VDAC_P.t2128 C6_P_btm.t59 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5970 a_12895_43640# a_12379_43268# a_12800_43628# VSS.t1159 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X5971 VDD.t1536 a_8308_43806# a_8483_43780# VDD.t1535 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X5972 VDAC_N.t544 C9_N_btm.t153 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5973 VDAC_P.t552 C9_P_btm.t150 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5974 VDAC_P.t2120 C9_P_btm.t149 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5975 VSS.t35 a_9521_45982.t14 a_10079_46532# VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5976 VDAC_P.t1072 C5_P_btm.t24 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5977 VSS.t59 a_12769_44594.t3 a_20107_43806# VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X5978 a_16475_45412# a_16335_47614# VDD.t1421 VDD.t1420 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X5979 VDD.t2390 VSS.t3727 VDD.t2389 VDD.t2388 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X5980 VDAC_P.t2112 C10_P_btm.t279 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5981 a_1947_45982# a_1597_45982# a_1852_45982# VDD.t2679 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X5982 VDAC_P.t288 C9_P_btm.t148 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5983 VSS.t2273 a_6235_46124# a_6196_46250# VSS.t2272 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5984 VSS.t1889 a_n268_44582# a_n381_43433# VSS.t1888 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X5985 VSS.t3699 C7_N_btm.t131 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5986 VDD.t1506 a_7705_45736# a_7735_45477# VDD.t1505 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5987 VDD.t1063 a_22959_44358# a_17738_32299.t2 VDD.t1062 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X5988 VDD.t2094 a_18319_44868# a_12769_44594.t1 VDD.t2093 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X5989 VSS.t2329 VSS.t2330 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5990 VDAC_P.t2104 C9_P_btm.t147 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5991 VDAC_N.t2088 C9_N_btm.t152 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5992 VDAC_N.t1056 C6_N_btm.t20 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5993 a_15033_46526# a_14658_46526# VSS.t1894 VSS.t1893 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X5994 VDAC_P.t1064 C7_P_btm.t123 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5995 VDAC_N.t2080 C10_N_btm.t268 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5996 VDAC_N.t32 C8_N_btm.t65 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5997 VDAC_P.t2096 C10_P_btm.t278 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5998 VDAC_P.t544 C10_P_btm.t277 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X5999 a_22031_44350# a_n2293_46508.t5 VDD.t110 VDD.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6000 VDAC_P.t2088 C8_P_btm.t68 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6001 VDAC_N.t2072 C9_N_btm.t151 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6002 VDAC_P.t1056 C8_P_btm.t67 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6003 VDAC_P.t2080 C10_P_btm.t276 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6004 VSS.t2299 VSS.t2300 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6005 VDAC_P.t32 C9_P_btm.t146 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6006 a_6536_46348# a_6322_46348# VDD.t1028 VDD.t1027 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X6007 VSS.t2283 VSS.t2284 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6008 a_n2810_46526.t0 a_n2840_46500# VSS.t2275 VSS.t2128 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X6009 VDAC_N.t1048 C10_N_btm.t267 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6010 VSS.t200 a_18394_35068.t15 a_11730_34132.t0 VSS.t199 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X6011 VDAC_N.t2064 C9_N_btm.t149 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6012 VDD.t1349 a_4651_47614# DATA[3].t6 VDD.t1348 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X6013 VDAC_N.t536 VSS.t3252 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6014 VDD.t2416 VSS.t3584 VDD.t2415 VDD.t2414 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X6015 a_22521_39947# a_22545_39429# VDD.t2088 VDD.t2087 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X6016 VDAC_P.t2072 C9_P_btm.t145 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6017 VDAC_N.t2056 C10_N_btm.t266 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6018 a_16671_47320# a_15163_45670.t10 a_16579_47320# VDD.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.155 ps=1.31 w=1 l=0.15
X6019 VSS.t2244 a_5655_43780# a_5613_43806# VSS.t2243 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6020 VDAC_N.t1040 C8_N_btm.t64 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6021 a_n1732_35090.t1 SMPL.t12 VDD.t3047 VDD.t3046 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6022 VDAC_N.t2048 C7_N_btm.t117 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6023 VDAC_P.t1048 C6_P_btm.t22 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6024 a_3726_37500# a_3754_38470.t8 VDAC_Ni.t7 VSS.t2842 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X6025 VDD.t2424 VSS.t3739 VDD.t2423 VDD.t2422 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X6026 VDAC_P.t2064 C8_P_btm.t66 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6027 VSS.t3472 VDD.t3217 VSS.t3471 VSS.t3470 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6028 a_10993_45982# a_9803_45982# a_10884_45982# VSS.t2580 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X6029 VSS.t1273 a_15187_44868# a_16750_46134# VSS.t1272 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X6030 VDAC_N.t280 C9_N_btm.t148 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6031 a_2587_44868.t2 a_20107_43806# VSS.t135 VSS.t134 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6032 VDAC_P.t536 C7_P_btm.t43 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6033 VDD.t1651 a_13536_43780# a_2755_43494.t2 VDD.t1650 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X6034 a_n2840_44868# a_n2661_44868# VSS.t906 VSS.t905 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X6035 a_9761_46565# a_n53_44363.t14 a_9547_46565# VDD.t560 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X6036 VDAC_P.t2056 C6_P_btm.t20 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6037 a_6325_45736# a_885_44868.t16 VDD.t2836 VDD.t2835 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X6038 a_5840_42718.t1 a_5663_42718# VSS.t898 VSS.t897 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6039 a_11599_42883# a_5734_30651.t7 VSS.t459 VSS.t458 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6040 VDD.t2347 VSS.t3806 VDD.t2346 VDD.t2345 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6041 VSS.t2586 a_9349_46539# a_9293_46565# VSS.t2585 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X6042 a_11017_45736# a_10684_45670# VDD.t693 VDD.t692 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X6043 VDAC_P.t1040 C10_P_btm.t275 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6044 VDAC_N.t2040 C10_N_btm.t265 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6045 VDAC_N.t1032 C10_N_btm.t264 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6046 VDAC_N.t2032 C7_N_btm.t40 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6047 SMPL_ON_N.t1 a_21789_35634# VSS.t2659 VSS.t2658 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6048 COMP_N.t7 a_1239_39043# VDD.t1730 VDD.t1729 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6049 a_7648_46892# a_7503_45982# VDD.t1283 VDD.t1282 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X6050 VDAC_P.t2048 C8_P_btm.t65 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6051 VDAC_N.t528 C9_N_btm.t147 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6052 VDAC_P.t280 C8_P_btm.t64 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6053 VSS.t3597 C9_N_btm.t532 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6054 VSS.t3640 C10_P_btm.t24 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6055 VDD.t2938 CAL_P.t4 VDD.t2938 VDD.t146 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X6056 a_16788_45144# a_6104_45706.t10 VDD.t3103 VDD.t3102 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X6057 VDAC_N.t2024 C9_N_btm.t145 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6058 a_15328_46134# a_13524_46832.t12 VDD.t546 VDD.t406 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6059 VDAC_N.t1024 C10_N_btm.t263 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6060 VDAC_P.t2040 C9_P_btm.t144 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6061 VDAC_N.t2016 C10_N_btm.t262 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6062 a_750_43628# a_135_43540.t38 VSS.t182 VSS.t181 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X6063 VDAC_P.t1032 C10_P_btm.t274 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6064 VDD.t437 a_7754_40130.t4 a_8912_37509.t0 VDD.t436 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X6065 VDAC_P.t2032 C10_P_btm.t273 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6066 VDAC_N.t152 C9_N_btm.t144 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6067 VDAC_N.t2008 C10_N_btm.t261 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6068 VDAC_P.t528 C9_P_btm.t143 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6069 VDAC_P.t2024 C10_P_btm.t272 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6070 a_n2840_43236# a_n2661_43244# VDD.t620 VDD.t619 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X6071 VSS.t1593 a_5419_47258# a_n2497_47846.t0 VSS.t1592 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6072 VDAC_P.t1024 C10_P_btm.t271 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6073 VDAC_P.t2016 C10_P_btm.t270 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6074 a_7493_43262# a_2587_44868.t20 VDD.t243 VDD.t242 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X6075 VSS.t1896 a_22959_45982# a_20405_31459.t0 VSS.t1355 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X6076 a_5918_46234# a_6196_46250# a_6152_46348# VDD.t992 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X6077 VDD.t1227 a_20283_43262# a_20383_42718# VDD.t1226 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6078 VDAC_P.t152 C10_P_btm.t269 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6079 a_n2074_43262.t3 a_n2104_43236# VDD.t768 VDD.t767 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X6080 VDAC_N.t1016 C7_N_btm.t39 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6081 VDAC_N.t2000 C6_N_btm.t19 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6082 VDAC_N.t520 C9_N_btm.t143 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6083 VDAC_P.t2008 C7_P_btm.t42 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6084 VDAC_N.t1992 C10_N_btm.t260 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6085 a_11455_44576.t3 a_13635_43566# VSS.t1246 VSS.t1245 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6086 VSS.t697 a_18259_46500# a_18190_46526# VSS.t696 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X6087 a_18879_45956# a_10227_47214.t9 VDD.t283 VDD.t282 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6088 VDAC_P.t1016 C9_P_btm.t142 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6089 a_12651_44576.t1 a_16579_43566# VSS.t1959 VSS.t1958 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6090 a_1412_46794.t0 a_8483_46830# VSS.t1402 VSS.t1401 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X6091 VDAC_N.t1008 C9_N_btm.t142 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6092 VDAC_P.t2000 C8_P_btm.t63 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6093 a_13819_44350# a_13469_44894# VDD.t774 VDD.t773 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X6094 VDAC_P.t520 C10_P_btm.t268 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6095 a_5536_44324# a_5387_44403# a_5832_44466# VDD.t860 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6096 VDAC_P.t1992 C9_P_btm.t141 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6097 VDAC_P.t1008 C10_P_btm.t267 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6098 VDAC_N.t1984 C9_N_btm.t141 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6099 VDAC_N.t272 C10_N_btm.t259 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6100 a_13635_43566# a_10227_47214.t22 VDD.t297 VDD.t296 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X6101 VSS.t3723 C0_N_btm.t4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6102 a_2512_45982# a_1431_45982# a_2165_46224# VDD.t687 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X6103 VREF.t57 a_n4515_30659.t8 C10_P_btm.t1060 VDD.t2994 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6104 VSS.t2535 VSS.t2536 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6105 VDAC_N.t1976 C10_N_btm.t258 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6106 a_10475_43433# a_9987_42968# VSS.t1696 VSS.t1695 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X6107 a_9898_44350# a_9179_44592# a_9335_44324# VSS.t2640 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X6108 VDAC_N.t1000 C8_N_btm.t63 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6109 VDAC_P.t1984 C10_P_btm.t265 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6110 VDAC_P.t272 C10_P_btm.t264 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6111 VDAC_N.t1968 C9_N_btm.t140 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6112 VDAC_N.t512 C10_N_btm.t257 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6113 a_4706_46892# a_135_43540.t18 VSS.t2772 VSS.t2771 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X6114 VDAC_N.t1960 C10_N_btm.t256 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6115 VDAC_P.t1976 VSS.t3377 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6116 VDAC_N.t992 C10_N_btm.t255 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6117 VDAC_P.t1000 C10_P_btm.t263 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6118 VDAC_P.t1968 C10_P_btm.t262 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6119 a_15437_47044# a_15139_47730# VDD.t1281 VDD.t1280 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X6120 VDAC_P.t512 C9_P_btm.t140 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6121 VDAC_N.t1952 C8_N_btm.t62 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6122 VDAC_N.t88 C10_N_btm.t254 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6123 a_13469_44894# a_12931_44894# VSS.t2635 VSS.t2634 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X6124 VDAC_P.t1960 C10_P_btm.t261 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6125 VDAC_N.t1944 C10_N_btm.t253 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6126 VDAC_P.t992 C9_P_btm.t139 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6127 VDAC_P.t1952 C10_P_btm.t260 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6128 a_15831_42883# a_5142_30651.t8 VDD.t124 VDD.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X6129 VDAC_N.t984 C10_N_btm.t252 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6130 a_8514_46232# a_1429_47222.t18 VDD.t328 VDD.t327 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X6131 VDAC_P.t88 C9_P_btm.t138 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6132 VDD.t253 a_2587_44868.t32 a_885_44868.t0 VDD.t252 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6133 VDAC_N.t1936 C10_N_btm.t251 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6134 VSS.t226 a_7557_43236.t18 a_13299_44716# VSS.t225 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X6135 DATA[0].t5 a_n1085_47874# VDD.t1948 VDD.t1947 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X6136 VDAC_P.t1944 C10_P_btm.t259 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6137 VDD.t2678 a_9349_46539# a_9761_46565# VDD.t2677 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X6138 a_11883_43806# a_11533_43806# a_11788_43806# VDD.t1465 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6139 VDAC_N.t504 C6_N_btm.t18 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6140 VDD.t1024 a_22591_45982# a_19921_31459.t3 VDD.t1023 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6141 VDD.t2661 a_n1552_42692# a_n1522_42718.t2 VDD.t2660 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X6142 VDAC_N.t1928 C7_N_btm.t37 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6143 VDAC_P.t984 C7_P_btm.t41 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6144 VDAC_P.t1936 C10_P_btm.t258 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6145 VDAC_N.t976 C6_N_btm.t17 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6146 VDAC_P.t504 C8_P_btm.t62 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6147 VDAC_N.t1920 C10_N_btm.t250 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6148 VDD.t126 a_n1551_44324.t10 a_22959_46534# VDD.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6149 VSS.t886 a_9159_43262# a_9898_44350# VSS.t885 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X6150 VDAC_P.t1928 C10_P_btm.t257 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6151 VDAC_P.t976 C8_P_btm.t61 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6152 VSS.t3159 VDD.t3155 VSS.t3158 VSS.t3157 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6153 a_6322_46348# a_6235_46124# a_5918_46234# VDD.t2238 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X6154 VSS.t639 a_13273_44868.t14 a_13207_44894# VSS.t638 sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X6155 VSS.t3779 C7_P_btm.t4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6156 VSS.t2908 a_6485_44582.t11 a_7781_43582# VSS.t2907 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X6157 a_2165_46224# a_1947_45982# VSS.t3000 VSS.t2999 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X6158 VSS.t1986 a_560_45670# a_n105_46195# VSS.t1985 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X6159 VDAC_N.t264 C9_N_btm.t139 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6160 VDAC_N.t1912 C10_N_btm.t249 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6161 VDAC_P.t1920 C10_P_btm.t256 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6162 a_n519_46532# a_n685_46532# VDD.t1580 VDD.t1579 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X6163 VDAC_N.t968 C10_N_btm.t248 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6164 VSS.t1797 a_4527_46830# a_4461_46904# VSS.t1796 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X6165 VDAC_N.t1904 C9_N_btm.t138 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6166 VDAC_P.t264 C9_P_btm.t137 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6167 VDAC_N.t496 C9_N_btm.t137 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6168 VDAC_N.t1896 C10_N_btm.t247 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6169 a_948_43806# a_33_43806# a_601_44048# VSS.t940 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6170 VDD.t445 a_7754_40130.t8 a_8912_37509.t2 VDD.t444 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X6171 a_11143_47588# a_11299_47832# VSS.t1443 VSS.t1442 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X6172 VSS.t1659 a_15192_46500# a_15113_47222# VSS.t1658 sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X6173 VDAC_N.t960 C10_N_btm.t1031 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6174 a_18497_46892# a_10227_47214.t24 VSS.t344 VSS.t343 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X6175 VSS.t39 a_9521_45982.t18 a_11367_43806# VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6176 VDD.t2489 VSS.t3690 VDD.t2488 VDD.t2487 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X6177 a_2043_45982# a_1597_45982# a_1947_45982# VSS.t2588 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6178 VSS.t1711 a_7276_45670# a_7016_46231# VSS.t1710 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X6179 a_10078_45144# a_7557_43236.t22 VDD.t224 VDD.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X6180 a_n2293_43780# a_n1827_44868.t12 VSS.t325 VSS.t299 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6181 a_13654_46032# a_13248_45956.t8 a_13661_46298# VDD.t395 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X6182 VDAC_P.t1912 C9_P_btm.t136 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6183 VDD.t3024 a_6485_44582.t26 a_8699_44894# VDD.t3023 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X6184 VDAC_P.t968 C10_P_btm.t255 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6185 VDAC_P.t1904 C10_P_btm.t254 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6186 VDD.t1190 a_9395_47044# a_4830_43958.t2 VDD.t1189 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X6187 VDAC_P.t496 C9_P_btm.t135 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6188 VDAC_N.t1888 C3_N_btm.t2 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6189 VDAC_P.t1896 C10_P_btm.t253 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6190 a_3541_42718# a_1847_45528.t26 VSS.t2811 VSS.t2810 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6191 VDAC_N.t144 C10_N_btm.t1013 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6192 VDD.t2571 VSS.t3629 VDD.t2570 VDD.t2569 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6193 VDAC_N.t1880 C8_N_btm.t61 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6194 a_169_45776# a_82_45670# a_83_45776# VSS.t1690 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X6195 VDAC_P.t960 C7_P_btm.t40 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6196 VDAC_N.t952 C10_N_btm.t992 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6197 VDD.t648 a_5536_44324# a_n1827_44324.t3 VDD.t647 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X6198 VSS.t3601 C10_P_btm.t31 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6199 VDAC_P.t1888 C9_P_btm.t134 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6200 VDAC_P.t144 C10_P_btm.t252 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6201 VDD.t2639 VSS.t3702 VDD.t2638 VDD.t2637 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X6202 VDAC_N.t1872 C8_N_btm.t60 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6203 VDAC_P.t1880 C10_P_btm.t251 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6204 VDAC_P.t952 C9_P_btm.t133 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6205 VSS.t2022 a_6519_43494# a_6243_45107# VSS.t2021 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X6206 VSS.t435 a_n2661_45956.t7 a_22223_43494# VSS.t434 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6207 VDAC_P.t1872 C9_P_btm.t132 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6208 VDAC_P.t488 C9_P_btm.t131 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6209 VDAC_N.t488 C10_N_btm.t906 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6210 VDAC_N.t1864 C10_N_btm.t773 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6211 VDAC_N.t944 C9_N_btm.t136 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6212 a_n2103_45412.t3 a_18970_45412# a_18918_45758# VSS.t2025 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6213 VDAC_P.t1864 C9_P_btm.t130 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6214 VDAC_N.t1856 C10_N_btm.t620 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6215 VDAC_N.t256 C10_N_btm.t598 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6216 a_396_43640# a_n685_43268# a_49_43236# VDD.t2226 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X6217 VDAC_N.t1848 C9_N_btm.t135 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6218 a_7557_43236.t0 a_11427_43566# VSS.t1165 VSS.t1164 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6219 VDAC_N.t936 C8_N_btm.t59 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6220 a_1947_45982# a_1431_45982# a_1852_45982# VSS.t759 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6221 VDAC_P.t944 C8_P_btm.t60 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6222 a_4049_43628# a_4005_43236# a_3883_43640# VSS.t1724 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X6223 a_4842_46309# a_885_44868.t30 VDD.t2850 VDD.t2849 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X6224 VDAC_P.t1856 C10_P_btm.t250 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6225 VSS.t2912 a_6485_44582.t14 a_8379_46134# VSS.t2911 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6226 VDD.t1993 a_3882_44324# a_n2103_43780.t6 VDD.t1992 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6227 VDAC_P.t256 C10_P_btm.t249 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6228 VDAC_P.t1848 C10_P_btm.t248 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6229 VDAC_N.t1840 C7_N_btm.t36 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6230 a_12448_43806# a_11367_43806# a_12101_44048# VDD.t1613 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X6231 a_n2472_44324# a_n2293_44332# VDD.t2095 VDD.t1140 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X6232 VDAC_N.t480 C10_N_btm.t520 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6233 VDAC_P.t936 C7_P_btm.t39 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6234 VDAC_P.t1840 C10_P_btm.t247 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6235 a_16385_44688# a_15730_45670.t12 VSS.t569 VSS.t568 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X6236 VDD.t2682 a_2165_46224# a_2055_46348# VDD.t2681 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X6237 VDAC_N.t1832 C6_N_btm.t16 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6238 VDAC_P.t480 C10_P_btm.t1030 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6239 VDAC_N.t928 C10_N_btm.t514 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6240 VDAC_N.t1824 C8_N_btm.t241 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6241 VDAC_P.t1832 C8_P_btm.t59 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6242 a_11046_46348# a_9969_45982# a_10884_45982# VDD.t1487 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6243 VDAC_N.t56 C9_N_btm.t134 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6244 VDAC_P.t928 C10_P_btm.t1011 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6245 VDAC_P.t1824 C10_P_btm.t966 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6246 VSS.t2006 a_1209_47588# a_999_47846# VSS.t2005 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6247 a_518_44670# a_636_42870# a_768_44670# VSS.t820 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6248 VDAC_N.t1816 C10_N_btm.t511 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6249 VDAC_N.t920 C8_N_btm.t190 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6250 a_7648_43806# a_7319_43262# VSS.t1980 VSS.t1979 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X6251 VSS.t155 a_10114_45276.t4 a_11415_45670# VSS.t154 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6252 VDD.t1682 a_18495_44868# a_18319_44868# VDD.t1681 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X6253 VDAC_P.t56 C9_P_btm.t129 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6254 a_426_47397# a_380_47222# VDD.t1403 VDD.t1402 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X6255 a_n1827_44868.t4 a_8850_45412# VDD.t660 VDD.t659 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6256 VDAC_P.t1816 C10_P_btm.t868 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6257 VDAC_N.t1808 C9_N_btm.t133 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6258 VSS.t2014 a_21908_43236# a_13878_32299.t0 VSS.t2013 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X6259 VDAC_N.t472 C10_N_btm.t499 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6260 VDAC_P.t920 C10_P_btm.t769 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6261 C0_P_btm.t0 a_n2442_45438.t4 VREF.t6 VDD.t157 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X6262 VDAC_P.t1808 C10_P_btm.t630 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6263 a_13635_43566# a_13460_43640# a_13814_43628# VSS.t842 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X6264 VDAC_N.t1800 C9_N_btm.t132 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6265 VREF.t44 a_22812_30659.t12 C10_N_btm.t26 VDD.t524 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6266 VDAC_N.t912 C9_N_btm.t131 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6267 VSS.t2064 a_5896_45670# a_5749_47222# VSS.t2063 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X6268 VDD.t25 a_9521_45982.t5 a_11367_43806# VDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6269 a_7309_44466# a_6485_44582.t21 VSS.t2919 VSS.t2918 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6270 a_5542_30651.t1 a_11183_42718# VSS.t726 VSS.t725 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6271 a_17583_46500# a_17786_46658# VDD.t1514 VDD.t1513 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X6272 VDAC_N.t1792 C10_N_btm.t496 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6273 VDAC_P.t472 C10_P_btm.t518 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6274 VDAC_P.t1800 C10_P_btm.t511 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6275 VDAC_N.t248 C10_N_btm.t491 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6276 VDAC_P.t912 C9_P_btm.t128 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6277 a_14757_43806# a_14331_44133# VSS.t777 VSS.t776 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X6278 VDAC_N.t1784 C10_N_btm.t488 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6279 VDD.t2082 a_396_43640# a_571_43566# VDD.t2081 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6280 VDAC_P.t1792 C9_P_btm.t127 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6281 C1_P_btm.t6 a_n2810_45438.t4 VREF.t73 VDD.t3087 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X6282 VDAC_N.t904 C8_N_btm.t120 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6283 VDAC_P.t248 C9_P_btm.t126 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6284 VDD.t1473 a_22521_40491# a_22459_39581# VDD.t726 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6285 VSS.t2422 VSS.t2423 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6286 a_12127_46744# a_18282_45670# VDD.t1712 VDD.t1711 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X6287 VDAC_N.t1776 C5_N_btm.t10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6288 a_2471_45046# a_1581_43806.t19 a_2617_45144# VDD.t2911 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6289 VDAC_P.t1784 C10_P_btm.t501 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6290 a_15309_45438# a_14953_45554# VSS.t2076 VSS.t2075 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X6291 VSS.t2413 VSS.t2414 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6292 VDAC_N.t464 C10_N_btm.t484 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6293 VDAC_N.t1768 VSS.t3322 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6294 VDD.t2531 VSS.t3731 VDD.t2530 VDD.t2529 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X6295 a_1700_43378# a_82_45670# VDD.t1632 VDD.t1631 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X6296 VDAC_N.t896 C10_N_btm.t481 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6297 a_6325_45736# a_885_44868.t26 VSS.t2756 VSS.t2755 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6298 VDAC_N.t1760 C10_N_btm.t474 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6299 VDAC_N.t136 C9_N_btm.t130 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6300 VDAC_N.t1752 C9_N_btm.t129 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6301 VDAC_N.t888 C10_N_btm.t471 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6302 VDAC_P.t904 C9_P_btm.t125 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6303 a_10884_45982# a_9969_45982# a_10537_46224# VSS.t1552 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X6304 VDAC_P.t1776 C9_P_btm.t124 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6305 VDAC_N.t1744 C9_N_btm.t128 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6306 VDAC_P.t464 C9_P_btm.t123 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6307 VDAC_P.t1768 C10_P_btm.t497 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6308 a_283_42692# a_927_42692.t25 VSS.t102 VSS.t101 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6309 VDAC_P.t896 C10_P_btm.t494 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6310 VDAC_P.t1760 C8_P_btm.t58 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6311 VDAC_P.t136 C8_P_btm.t57 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6312 a_11017_45736# a_10684_45670# VSS.t763 VSS.t762 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6313 VDAC_N.t456 C10_N_btm.t467 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6314 VDD.t1617 a_12448_43806# a_12623_43780# VDD.t1616 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6315 a_4700_46134# a_3165_45982# a_4842_46309# VDD.t1389 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X6316 VDD.t361 a_n690_43494.t14 a_7227_46532# VDD.t360 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6317 w_11534_34010.t14 a_11730_34132.t5 w_11534_34010.t14 w_11534_34010.t13 sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X6318 a_n2472_44868# a_n2293_44868# VSS.t1492 VSS.t1491 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X6319 a_9943_45046# a_10215_44874# VSS.t1015 VSS.t1014 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6320 VDAC_N.t1736 C10_N_btm.t246 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6321 VDAC_N.t880 C8_N_btm.t117 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6322 VDAC_P.t1752 C1_P_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6323 a_n2833_42692# a_n2497_42870.t8 VSS.t2877 VSS.t2876 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X6324 a_14087_32299.t3 a_22223_43270# VDD.t668 VDD.t667 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X6325 VDD.t670 a_14819_44582# a_14133_43780# VDD.t669 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X6326 VDD.t1756 a_4527_46830# a_4514_46526# VDD.t1755 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6327 VDD.t1145 a_8391_47044# a_135_43540.t4 VDD.t1144 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X6328 VDAC_P.t888 C7_P_btm.t37 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6329 VSS.t1638 a_18879_43780# a_18813_43806# VSS.t1637 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X6330 VSS.t1961 a_16579_43566# a_16513_43640# VSS.t1960 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X6331 EN_VIN_BSTR_N.t2 a_18394_35068.t11 w_11534_34010.t7 w_11534_34010.t6 sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X6332 VDAC_N.t1728 C10_N_btm.t243 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6333 VDAC_P.t1744 C10_P_btm.t489 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6334 a_8912_37509.t34 VDAC_P.t456 a_5088_37509.t16 VDD.t2247 sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X6335 VDAC_N.t240 C7_N_btm.t35 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6336 a_284_47222# a_n53_44363.t18 a_426_47397# VDD.t562 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X6337 a_10623_47307# a_10467_47212# a_10768_47436# VDD.t2133 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X6338 VDAC_N.t1720 C10_N_btm.t242 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6339 a_288_43806# a_171_44019# VDD.t1450 VDD.t1449 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X6340 VDAC_P.t1736 C10_P_btm.t486 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6341 a_n2472_43236# a_n2293_43244# VDD.t1637 VDD.t1636 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X6342 VDAC_N.t872 C10_N_btm.t240 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6343 VDAC_N.t1712 C10_N_btm.t239 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6344 VDD.t1860 a_5847_47614# DATA[4].t7 VDD.t1859 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6345 VDAC_P.t880 C10_P_btm.t482 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6346 VSS.t3171 VDD.t3159 VSS.t3170 VSS.t3169 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6347 VDAC_P.t1728 C10_P_btm.t479 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6348 VDAC_N.t448 C10_N_btm.t235 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6349 a_13105_44716# a_12651_44576.t22 a_13023_44716# VSS.t2872 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X6350 VDAC_N.t1704 C9_N_btm.t127 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6351 VDAC_P.t240 C10_P_btm.t472 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6352 VIN_N.t4 EN_VIN_BSTR_N.t22 C10_N_btm.t17 VSS.t449 sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X6353 a_5734_30651.t2 a_9343_42718# VDD.t2235 VDD.t2234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X6354 VDAC_N.t864 C8_N_btm.t56 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6355 a_14953_45554# a_15033_46526# VDD.t1854 VDD.t1853 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X6356 VDAC_P.t1720 C10_P_btm.t469 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6357 VDAC_N.t1696 VSS.t3321 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6358 VSS.t3425 VDD.t3199 VSS.t3424 VSS.t3423 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6359 VDAC_P.t872 C8_P_btm.t253 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6360 VDAC_N.t80 C10_N_btm.t234 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6361 a_n61_43262# a_n685_43268# a_n169_43640# VDD.t2229 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X6362 a_15192_46500# a_15309_45438# a_15321_46526# VDD.t2030 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X6363 a_7372_45670# a_7415_44466# VDD.t1263 VDD.t1262 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X6364 VDAC_N.t1688 C9_N_btm.t126 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6365 VDAC_P.t1712 C7_P_btm.t36 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6366 VDAC_N.t856 C9_N_btm.t125 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6367 VDAC_P.t448 C9_P_btm.t122 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6368 VDAC_N.t1680 C9_N_btm.t124 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6369 a_n1429_43262# a_n1459_43236.t13 VDD.t543 VDD.t542 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6370 a_4152_45804# a_4035_45609# VDD.t1193 VDD.t1192 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X6371 VDAC_P.t1704 C5_P_btm.t14 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6372 VCM.t39 a_3222_30651.t20 VDAC_P.t7 VSS.t672 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X6373 a_18231_44728# a_17715_44356# a_18136_44716# VSS.t703 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6374 VDD.t2940 CAL_P.t5 VDD.t2939 VDD.t148 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=10
X6375 VSS.t3099 VDD.t3135 VSS.t3098 VSS.t3097 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6376 VDD.t365 a_n690_43494.t18 a_3271_46532# VDD.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6377 VDAC_N.t440 C10_N_btm.t232 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6378 VDD.t1760 a_4527_46830# a_4322_46134# VDD.t1759 sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X6379 VDAC_N.t1672 C9_N_btm.t123 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6380 VDAC_P.t1696 VSS.t3395 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6381 VDAC_N.t848 C10_N_btm.t231 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6382 VDAC_P.t80 C10_P_btm.t245 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6383 a_15133_45982# a_15079_46134# VSS.t1693 VSS.t1692 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6384 VDAC_P.t1688 C9_P_btm.t121 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6385 VDAC_N.t1664 C9_N_btm.t122 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6386 VSS.t1370 a_10251_45454# a_19003_43262# VSS.t1369 sky130_fd_pr__nfet_01v8 ad=0.1359 pd=1.1 as=0.1113 ps=1.37 w=0.42 l=0.15
X6387 VDAC_P.t856 C10_P_btm.t244 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6388 VDAC_N.t232 C10_N_btm.t228 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6389 a_1387_45670# a_1659_45528# VSS.t1878 VSS.t1877 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6390 VDAC_P.t1680 C9_P_btm.t120 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6391 VDAC_P.t440 C10_P_btm.t241 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6392 VDAC_P.t1672 C9_P_btm.t513 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6393 a_n2288_42692# a_n2109_42692.t5 VDD.t3084 VDD.t3083 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X6394 VDAC_Pi.t5 VSS.t3788 a_5700_37509.t17 VDD.t2580 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X6395 VSS.t2363 VSS.t2364 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6396 VSS.t2545 VSS.t2546 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6397 VDAC_P.t848 C10_P_btm.t240 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6398 a_10500_46892# a_10383_46697# VSS.t1103 VSS.t1102 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X6399 VDAC_N.t1656 C10_N_btm.t227 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6400 VDAC_N.t840 C10_N_btm.t225 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6401 VSS.t683 a_13273_44868.t11 a_15091_44440# VSS.t682 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6402 a_325_46224# a_107_45982# VDD.t623 VDD.t622 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X6403 VDAC_N.t1648 C9_N_btm.t501 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6404 VDAC_N.t432 C10_N_btm.t224 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6405 VDAC_P.t1664 C10_P_btm.t238 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6406 a_6519_43494# a_6631_44582# a_6665_43262# VDD.t1444 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6407 VDAC_N.t1640 C10_N_btm.t218 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6408 DATA[4].t1 a_5847_47614# VSS.t1899 VSS.t1898 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6409 a_11606_43628# a_10227_47214.t40 VSS.t633 VSS.t632 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X6410 a_7961_46500# a_7743_46904# VSS.t1299 VSS.t1298 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X6411 VDAC_N.t832 C8_N_btm.t55 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6412 VDAC_P.t232 C9_P_btm.t500 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6413 a_5382_44582# a_4987_45742# VSS.t1342 VSS.t1341 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X6414 VDAC_P.t1656 C8_P_btm.t234 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6415 a_16561_45982# a_16085_45982# VDD.t991 VDD.t990 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.195 ps=1.39 w=1 l=0.15
X6416 VDAC_N.t1632 C10_N_btm.t217 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6417 VDAC_N.t128 C10_N_btm.t215 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6418 VDAC_P.t840 C10_P_btm.t237 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6419 a_2216_46758# a_2424_46794.t8 a_2358_46892# VSS.t2854 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X6420 VDAC_P.t1648 C10_P_btm.t233 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6421 VDD.t3096 a_6104_45706.t3 a_14647_43494# VDD.t3095 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X6422 a_2343_47070# a_2167_46526# VSS.t2136 VSS.t2135 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6423 a_3882_44324# a_3576_44364# VSS.t1151 VSS.t1150 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.11975 ps=1.045 w=0.42 l=0.15
X6424 VDAC_N.t1624 C7_N_btm.t34 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6425 VDAC_N.t824 C10_N_btm.t214 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6426 VSS.t1982 a_7347_43494# a_7319_43262# VSS.t1981 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X6427 VDAC_P.t432 C7_P_btm.t35 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6428 VSS.t2163 a_8204_45412# a_n2103_44324.t1 VSS.t2162 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X6429 VDAC_N.t1616 C9_N_btm.t356 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6430 VCM.t1 a_5142_30651.t5 C8_N_btm.t0 VSS.t121 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X6431 VDAC_P.t1640 C6_P_btm.t19 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6432 VDAC_N.t424 C4_N_btm.t14 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6433 a_3726_37500# CAL_P.t6 a_11206_38545.t4 VDD.t2941 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X6434 a_2587_44868.t3 a_20107_43806# VSS.t139 VSS.t138 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X6435 VDD.t3055 SMPL.t22 a_n1732_35090.t6 VDD.t3054 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6436 VDAC_N.t1608 C10_N_btm.t210 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6437 VDAC_P.t832 C9_P_btm.t398 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6438 VDAC_P.t1632 VSS.t3391 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6439 VDAC_P.t128 C9_P_btm.t351 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6440 VDAC_N.t816 C9_N_btm.t289 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6441 a_n2288_47588# a_n2109_47596.t4 VSS.t461 VSS.t460 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X6442 VDAC_P.t1624 C10_P_btm.t232 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6443 VDAC_N.t1600 C10_N_btm.t211 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6444 VDAC_N.t224 C9_N_btm.t252 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6445 VDAC_P.t824 C9_P_btm.t299 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6446 a_2755_43494.t3 a_13536_43780# VDD.t1649 VDD.t1648 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X6447 a_n1741_42692# a_n1735_43236.t10 VSS.t677 VSS.t676 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6448 a_10595_46904# a_10245_46532# a_10500_46892# VDD.t1934 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6449 VDAC_N.t1592 C9_N_btm.t246 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6450 VDD.t2888 a_1847_45528.t20 a_1659_45528# VDD.t2887 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6451 VDAC_N.t808 C10_N_btm.t209 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6452 VSS.t3804 C10_P_btm.t17 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6453 a_5139_44019# a_4651_44350# VDD.t1793 VDD.t1792 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6454 VDAC_P.t1616 C10_P_btm.t230 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6455 a_10687_43640# a_10337_43268# a_10592_43628# VDD.t1939 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X6456 VDAC_N.t1584 C10_N_btm.t208 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6457 VDD.t2019 a_5749_47222# a_5839_47070# VDD.t2018 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6458 VDAC_N.t416 C10_N_btm.t207 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6459 a_49_46500# a_n169_46904# VSS.t1330 VSS.t1329 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X6460 VDAC_N.t1576 C10_N_btm.t206 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6461 VDAC_P.t424 C10_P_btm.t229 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6462 VSS.t1628 a_10623_47307# a_10554_47436# VSS.t1627 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X6463 VDAC_N.t800 C10_N_btm.t205 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6464 a_12438_45412# a_12684_45276# VDD.t1012 VDD.t1011 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.17575 ps=1.395 w=0.42 l=0.15
X6465 VDAC_P.t1608 C10_P_btm.t226 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6466 VDAC_N.t1568 C9_N_btm.t243 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6467 a_11971_46500# a_12127_46744# VDD.t1046 VDD.t1045 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X6468 VSS.t2665 a_21789_35634# SMPL_ON_N.t0 VSS.t2664 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6469 VSS.t1163 a_11427_43566# a_11361_43640# VSS.t1162 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X6470 VDD.t739 a_4704_47044# a_4035_45609# VDD.t738 sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X6471 VDAC_N.t40 C10_N_btm.t204 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6472 VDAC_N.t1560 C9_N_btm.t239 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6473 VDAC_P.t816 C10_P_btm.t225 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6474 a_8848_44868# a_1412_46794.t11 VSS.t153 VSS.t152 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X6475 VDAC_P.t1600 C9_P_btm.t268 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6476 VDAC_P.t224 C10_P_btm.t223 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6477 VDAC_P.t1592 C8_P_btm.t191 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6478 VDD.t2723 a_n2038_35608# SMPL_ON_P.t5 VDD.t2722 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6479 VDD.t2618 VSS.t3624 VDD.t2617 VDD.t2616 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X6480 a_6038_45477# a_885_44868.t13 VDD.t2832 VDD.t2831 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X6481 VDAC_P.t808 C10_P_btm.t222 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6482 VSS.t3809 C7_N_btm.t132 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6483 VSS.t2732 a_1847_45528.t16 a_3179_44403# VSS.t2731 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X6484 VDAC_P.t1584 C10_P_btm.t216 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6485 a_18569_46892# a_18190_46526# a_18497_46892# VSS.t1126 sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X6486 VDAC_N.t792 C7_N_btm.t32 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6487 VDD.t2948 a_2424_46794.t10 a_n1551_45412.t6 VDD.t2947 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6488 VDD.t2624 VSS.t3685 VDD.t2623 VDD.t2622 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X6489 VDAC_N.t1552 C10_N_btm.t203 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6490 VDAC_P.t416 C10_P_btm.t215 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6491 a_n2497_47846.t2 a_1429_47222.t14 VSS.t388 VSS.t387 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6492 a_4005_46500# a_3787_46904# VSS.t2143 VSS.t2142 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X6493 a_18704_45982# a_17623_45982# a_18357_46224# VDD.t1083 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X6494 VDD.t725 a_18357_44048# a_18247_44172# VDD.t724 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X6495 a_22733_47833# DEBUG_MUX[3].t1 VSS.t2983 VSS.t2982 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6496 VDAC_N.t408 C6_N_btm.t15 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6497 VDAC_N.t1544 C9_N_btm.t236 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6498 VDAC_P.t1576 C7_P_btm.t34 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6499 VDAC_P.t800 C0_P_btm.t4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6500 VDAC_N.t784 C9_N_btm.t118 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6501 VDAC_P.t1568 C9_P_btm.t258 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6502 a_14204_44350# a_13725_44350# VDD.t1844 VDD.t1843 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1725 ps=1.345 w=1 l=0.15
X6503 VDAC_N.t1536 C8_N_btm.t53 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6504 VDD.t770 a_n2104_43236# a_n2074_43262.t2 VDD.t769 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X6505 VDAC_P.t40 C10_P_btm.t212 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6506 VDAC_P.t1560 C7_P_btm.t33 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6507 VDAC_N.t216 VSS.t3298 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6508 C5_P_btm.t0 a_n2074_47070.t4 VREF.t5 VDD.t144 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X6509 a_663_47874# a_999_47846# VDD.t1960 VDD.t1959 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X6510 VDAC_P.t792 C9_P_btm.t254 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6511 VDAC_N.t1528 C10_N_btm.t202 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6512 a_7851_44172# a_5655_43780# VDD.t2205 VDD.t2204 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X6513 VDAC_N.t776 C9_N_btm.t117 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6514 VDAC_P.t1552 C10_P_btm.t213 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6515 a_2587_44868.t6 a_20107_43806# VDD.t142 VDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6516 VDAC_P.t408 C9_P_btm.t242 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6517 a_3699_43780# a_3524_43806# a_3878_43806# VSS.t684 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X6518 VDAC_P.t1544 C10_P_btm.t211 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6519 VDAC_N.t1520 C9_N_btm.t115 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6520 VDAC_P.t784 C9_P_btm.t239 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6521 VDAC_N.t400 C10_N_btm.t201 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6522 VDAC_P.t1536 C10_P_btm.t210 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6523 VDAC_N.t1512 C9_N_btm.t114 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6524 VDAC_N.t768 C10_N_btm.t200 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6525 a_8969_43582# a_6485_44582.t23 VSS.t2921 VSS.t2920 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6526 VSS.t2103 a_19520_46500# a_n2109_47596.t0 VSS.t2102 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X6527 VDAC_P.t216 C10_P_btm.t209 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6528 VDAC_N.t1504 C10_N_btm.t199 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6529 a_3754_39964# a_7754_39964# VSS.t693 sky130_fd_pr__res_high_po_0p35 l=18
X6530 VSS.t3703 C10_N_btm.t1073 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6531 VDD.t315 a_n1827_45412.t11 a_22959_47070# VDD.t314 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6532 VSS.t2438 VSS.t2439 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6533 VSS.t163 a_10114_45276.t11 a_14819_44582# VSS.t162 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6534 VDAC_P.t1528 C10_P_btm.t208 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6535 VDAC_N.t120 C8_N_btm.t52 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6536 VDAC_N.t1496 C9_N_btm.t111 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6537 VSS.t230 a_7557_43236.t24 a_10447_44403# VSS.t229 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X6538 VDAC_P.t776 C6_P_btm.t18 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6539 a_11059_45956# a_10884_45982# a_11238_45982# VSS.t850 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X6540 VDAC_P.t1520 C8_P_btm.t176 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6541 a_18327_44728# a_17881_44356# a_18231_44728# VSS.t2683 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6542 a_570_44324# a_546_43100# VDD.t1763 VDD.t1762 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.17575 ps=1.395 w=0.42 l=0.15
X6543 VDAC_N.t760 VSS.t3257 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6544 a_n107_47098# a_n194_47222# a_n193_47098# VSS.t1035 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X6545 VDAC_N.t1488 C10_N_btm.t197 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6546 VDAC_N.t392 C6_N_btm.t14 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6547 VDAC_N.t1480 C7_N_btm.t31 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6548 VDAC_N.t752 C10_N_btm.t196 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6549 a_5441_46500# a_5382_44582# a_5945_46846# VSS.t2069 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X6550 VDAC_P.t400 C10_P_btm.t207 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6551 VDAC_P.t1512 C6_P_btm.t17 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6552 a_1343_38525.t5 a_1177_38525# VDD.t2767 VDD.t2766 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6553 VDAC_P.t768 C10_P_btm.t206 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6554 VDAC_P.t1504 C8_P_btm.t130 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6555 VDD.t273 a_n1741_47596.t6 a_22399_44894# VDD.t272 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6556 VDAC_P.t120 C8_P_btm.t123 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6557 a_19058_45982# a_10227_47214.t26 VSS.t346 VSS.t345 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X6558 VDAC_N.t1472 C9_N_btm.t110 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6559 VCM.t24 a_5734_30651.t5 C5_N_btm.t1 VSS.t456 sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X6560 VDD.t2636 VSS.t3634 VDD.t2635 VDD.t2634 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6561 a_7556_42692# a_7735_42692# VSS.t1469 VSS.t1468 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X6562 VDAC_P.t1496 C8_P_btm.t117 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6563 a_18803_47070# a_18530_47070# VSS.t1950 VSS.t1949 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X6564 VDAC_N.t208 C10_N_btm.t195 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6565 a_19921_31459.t2 a_22591_45982# VDD.t1022 VDD.t1021 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X6566 VSS.t1063 a_16750_46134# a_16703_45982# VSS.t1062 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.1755 ps=1.84 w=0.65 l=0.15
X6567 VDAC_N.t1464 C9_N_btm.t108 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6568 a_14573_47070# a_14219_47070# VSS.t844 VSS.t843 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X6569 VDAC_P.t760 C10_P_btm.t205 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6570 a_18822_46526# a_18103_46768# a_18259_46500# VSS.t1840 sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X6571 VDAC_P.t1488 C10_P_btm.t204 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6572 VDAC_N.t744 C10_N_btm.t194 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6573 VDAC_N.t1456 C10_N_btm.t193 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6574 VDAC_P.t392 C8_P_btm.t114 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6575 VDAC_P.t1480 C10_P_btm.t203 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6576 VSS.t837 a_14133_43780# a_14552_43806# VSS.t836 sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X6577 VDD.t2890 a_1847_45528.t21 a_2801_42968# VDD.t2889 sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X6578 VSS.t3093 VDD.t3133 VSS.t3092 VSS.t3091 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X6579 VSS.t3114 VDD.t3140 VSS.t3113 VSS.t3112 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6580 a_11252_43640# a_10171_43268# a_10905_43236# VDD.t2147 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X6581 a_15121_46232# a_15079_46134# a_15037_46232# VDD.t1635 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6582 VDAC_N.t384 C9_N_btm.t107 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6583 VDAC_P.t752 C9_P_btm.t235 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6584 VDAC_N.t1448 C8_N_btm.t51 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6585 VSS.t3638 C3_P_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6586 VDAC_P.t1472 C9_P_btm.t232 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6587 a_7182_45260# a_6105_44894# a_7020_44894# VDD.t1547 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6588 VDAC_P.t208 VSS.t3370 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6589 VDAC_P.t1464 C6_P_btm.t16 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6590 VDAC_P.t744 C10_P_btm.t202 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6591 VDAC_N.t736 C5_N_btm.t9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6592 VDAC_P.t1456 C10_P_btm.t201 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6593 VDAC_N.t1440 C7_N_btm.t30 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6594 VDAC_N.t72 C10_N_btm.t192 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6595 VDD.t1750 a_4700_46134# a_4061_47044# VDD.t1749 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X6596 VSS.t1880 a_1387_45670# a_656_45670# VSS.t1879 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X6597 a_1617_44466# a_1429_47222.t16 a_1522_44466# VDD.t325 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X6598 VDAC_N.t1432 C10_N_btm.t191 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6599 VDAC_P.t384 C9_P_btm.t227 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6600 VDD.t118 a_15163_45670.t6 a_15691_47614# VDD.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6601 VDD.t1339 a_12427_46758# a_10684_45670# VDD.t1338 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X6602 VDAC_N.t728 C7_N_btm.t29 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6603 VDAC_N.t1424 C9_N_btm.t106 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6604 VDAC_N.t376 C9_N_btm.t105 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6605 VDAC_P.t1448 C7_P_btm.t32 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6606 a_11788_43806# a_11671_44019# VSS.t1001 VSS.t1000 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X6607 VSS.t416 a_n690_43494.t8 a_3731_45444# VSS.t415 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6608 VDAC_P.t736 C9_P_btm.t224 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6609 VDAC_P.t1440 C9_P_btm.t220 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6610 VSS.t3247 VDD.t3186 VSS.t3246 VSS.t3245 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X6611 VDAC_P.t72 C10_P_btm.t200 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6612 VDAC_N.t1416 C10_N_btm.t190 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6613 VDAC_P.t1432 C9_P_btm.t119 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6614 VDAC_P.t728 C9_P_btm.t114 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6615 VDAC_N.t720 C10_N_btm.t189 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6616 VDAC_P.t1424 C10_P_btm.t199 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6617 VDD.t971 a_22223_47622# a_21788_30659.t3 VDD.t970 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6618 VDAC_P.t376 C8_P_btm.t108 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6619 VDAC_N.t1408 C10_N_btm.t188 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6620 VDD.t2279 VSS.t3567 VDD.t2278 VDD.t2277 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X6621 VDAC_N.t200 C9_N_btm.t104 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6622 a_n690_43494.t3 a_6635_47044# VDD.t2111 VDD.t2110 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6623 VDAC_P.t1416 C10_P_btm.t198 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6624 a_4974_45438# a_3897_45444# a_4812_45816# VDD.t2125 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6625 VDAC_P.t720 C10_P_btm.t197 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6626 a_n1827_44324.t2 a_5536_44324# VDD.t646 VDD.t645 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X6627 VDAC_N.t1400 C9_N_btm.t103 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6628 VDAC_P.t1408 C10_P_btm.t196 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6629 VREF.t33 a_22812_30659.t5 C10_N_btm.t19 VDD.t517 sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=0.35
X6630 VSS.t359 a_n1827_45412.t10 a_22959_47070# VSS.t128 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6631 a_22223_43494# a_n2661_45956.t5 VSS.t433 VSS.t432 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6632 VDAC_P.t200 C10_P_btm.t195 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6633 VDAC_N.t712 C10_N_btm.t187 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6634 w_1375_34946.t1 EN_VIN_BSTR_P.t18 VDD.t487 w_1375_34946.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X6635 CLK_DATA.t5 a_n2833_47874# VDD.t1311 VDD.t1310 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X6636 VDAC_N.t1392 C10_N_btm.t186 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6637 VDAC_N.t368 C8_N_btm.t50 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6638 a_n194_47222# a_571_46830# VSS.t1128 VSS.t1127 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X6639 VDAC_N.t1384 C7_N_btm.t28 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6640 VDD.t1952 a_n1085_47874# DATA[0].t7 VDD.t1951 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X6641 a_6974_31099.t0 a_20383_42718# VSS.t2256 VSS.t2255 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6642 a_5655_43780# a_9343_43806# VDD.t2180 VDD.t2179 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X6643 VDAC_P.t1400 C10_P_btm.t194 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6644 VDAC_N.t704 C8_N_btm.t49 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6645 VDAC_P.t712 C3_P_btm.t10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6646 a_n264_46892# a_n381_46697# VDD.t1235 VDD.t1234 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X6647 a_15317_47730# a_15163_45670.t11 a_15221_47730# VDD.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6648 VDAC_P.t1392 C10_P_btm.t193 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6649 VDAC_P.t368 C10_P_btm.t192 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6650 VDAC_P.t1384 C10_P_btm.t191 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6651 VDD.t1901 a_11160_46904# a_11335_46830# VDD.t1900 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6652 VDAC_N.t1376 C6_N_btm.t13 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6653 VDD.t2162 a_14635_44324# a_15323_44894# VDD.t2161 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X6654 VDAC_N.t112 C8_N_btm.t48 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6655 VDAC_P.t704 C10_P_btm.t190 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6656 VDAC_N.t1368 C10_N_btm.t185 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6657 VDAC_P.t1376 C10_P_btm.t189 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6658 VDAC_N.t696 C8_N_btm.t47 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6659 VDAC_N.t1360 C9_N_btm.t102 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6660 VDD.t823 a_601_44048# a_491_44172# VDD.t822 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X6661 VDAC_P.t112 VSS.t3373 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6662 VDD.t313 a_n1827_45412.t9 a_n2661_44332# VDD.t278 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6663 VDAC_P.t1368 C8_P_btm.t105 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6664 VDAC_N.t360 C9_N_btm.t101 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6665 VREF.t17 a_n2467_30659.t10 C9_P_btm.t11 VDD.t583 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6666 a_13457_46892# a_14470_46526# a_14658_46526# VSS.t2998 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.151025 ps=1.285 w=0.42 l=0.15
X6667 a_6270_43806# a_5655_43780# VSS.t2234 VSS.t2233 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X6668 VDD.t1564 a_1123_43780# a_1110_44172# VDD.t1563 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6669 VDAC_P.t696 C9_P_btm.t113 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6670 VDAC_N.t1352 C10_N_btm.t184 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6671 VDD.t2421 VSS.t3586 VDD.t2420 VDD.t2299 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6672 VDAC_N.t688 C10_N_btm.t91 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6673 VDAC_P.t1360 C9_P_btm.t111 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6674 VDAC_N.t1344 C8_N_btm.t46 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6675 VDAC_P.t360 C9_P_btm.t110 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6676 VDAC_P.t1352 C9_P_btm.t107 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6677 VDAC_N.t192 C10_N_btm.t182 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6678 a_768_44670# a_636_42870# a_518_44670# VSS.t825 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6679 a_11415_45670# a_10259_42870.t12 VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X6680 VDAC_N.t1336 C9_N_btm.t100 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6681 VDAC_N.t680 C7_N_btm.t27 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6682 a_11671_44019# a_11183_44350# VDD.t961 VDD.t960 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X6683 VDAC_P.t688 C7_P_btm.t31 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6684 VSS.t1190 a_2645_46824# a_2579_46892# VSS.t1189 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X6685 VSS.t1398 a_22591_43958# a_22591_43806# VSS.t1397 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6686 VDAC_N.t1328 C9_N_btm.t99 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6687 VDAC_N.t352 C10_N_btm.t181 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6688 VDAC_P.t1344 C10_P_btm.t188 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6689 VSS.t3741 C5_P_btm.t4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6690 VDAC_P.t192 C9_P_btm.t106 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6691 VDAC_P.t1336 C5_P_btm.t13 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6692 VDAC_P.t680 C9_P_btm.t104 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6693 VDAC_P.t1328 C8_P_btm.t101 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6694 VDAC_P.t352 C9_P_btm.t103 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6695 VSS.t2931 a_1736_39587.t4 a_1239_39587# VSS.t516 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6696 VDAC_N.t1320 C4_N_btm.t6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6697 VDAC_P.t1320 C10_P_btm.t187 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6698 VSS.t2028 a_1387_44582# a_n172_44582# VSS.t2027 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X6699 a_n1459_43236.t7 a_570_44324# VDD.t1592 VDD.t1591 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6700 VDAC_N.t672 C10_N_btm.t180 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6701 VDAC_N.t1312 C9_N_btm.t98 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6702 VDAC_P.t672 C10_P_btm.t186 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6703 VSS.t1764 a_21755_44350# a_22223_44358# VSS.t1763 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6704 VDAC_N.t48 C10_N_btm.t179 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6705 VDAC_N.t1304 C8_N_btm.t45 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6706 VDAC_P.t1312 C10_P_btm.t185 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6707 a_15689_44048# a_15471_43806# VDD.t1417 VDD.t1416 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X6708 a_6985_45438# a_6707_45776# VSS.t1584 VSS.t1583 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X6709 VDAC_P.t48 C9_P_btm.t99 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6710 VDAC_N.t664 C9_N_btm.t97 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6711 VDAC_P.t1304 C10_P_btm.t184 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6712 a_12101_44048# a_11883_43806# VSS.t795 VSS.t794 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X6713 VDD.t2715 a_8848_44868# a_n1925_47044.t3 VDD.t2714 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X6714 VSS.t2537 VSS.t2538 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6715 a_383_43806# a_n133_43806# a_288_43806# VSS.t910 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X6716 VDAC_N.t1296 C10_N_btm.t178 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6717 VDD.t2411 VSS.t3756 VDD.t2410 VDD.t2409 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X6718 a_2617_45144# a_2755_43494.t8 a_2471_45046# VDD.t423 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X6719 VDAC_P.t664 C10_P_btm.t90 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6720 a_10227_47214.t2 a_11795_47044# VSS.t2657 VSS.t2656 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6721 VDAC_N.t344 VSS.t3303 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6722 VDAC_P.t1296 C9_P_btm.t98 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6723 a_2627_43262# a_2755_43494.t7 a_2709_43582# VSS.t507 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X6724 a_8662_46892# a_135_43540.t26 VSS.t2780 VSS.t2779 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X6725 VDAC_N.t1288 C8_N_btm.t44 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6726 a_14470_46526# a_13248_45956.t18 VSS.t487 VSS.t486 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6727 VSS.t2375 VSS.t2376 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6728 VDAC_N.t656 C6_N_btm.t12 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6729 a_6038_45804# a_885_44868.t32 VSS.t2764 VSS.t2763 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X6730 VDAC_P.t344 C7_P_btm.t30 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6731 a_9350_43628# a_9304_43494# VSS.t722 VSS.t721 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X6732 VDAC_P.t1288 C8_P_btm.t56 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6733 VDAC_N.t1280 C8_N_btm.t43 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6734 a_2055_46348# a_1431_45982# a_1947_45982# VDD.t690 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X6735 VDAC_P.t656 VSS.t3365 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6736 VDAC_P.t1280 C8_P_btm.t53 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6737 VDAC_P.t184 C7_P_btm.t29 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6738 VDAC_P.t1272 C10_P_btm.t182 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6739 VDD.t629 a_5129_45956# a_5159_46309# VDD.t628 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6740 VDAC_P.t648 C9_P_btm.t96 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6741 VDAC_P.t1264 VSS.t3340 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6742 VDAC_P.t336 C10_P_btm.t181 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6743 a_8912_37509.t10 VDAC_N.t184 a_5700_37509.t4 VDD.t2251 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X6744 a_n2810_43806.t2 a_n2840_43780# VDD.t1522 VDD.t879 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X6745 VSS.t2448 VSS.t2449 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6746 a_18689_45412# a_18879_45956# VSS.t705 VSS.t704 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X6747 VDAC_P.t1256 C10_P_btm.t180 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6748 a_1633_46824# a_885_44868.t15 VSS.t2746 VSS.t2745 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6749 VDAC_N.t1272 C10_N_btm.t177 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6750 VSS.t2207 a_4527_43566# a_927_42692.t2 VSS.t2206 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X6751 VSS.t2042 a_3541_42718# a_3823_42718# VSS.t2041 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6752 VDAC_N.t648 C9_N_btm.t96 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6753 VDAC_N.t1264 C10_N_btm.t176 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6754 VDAC_P.t640 C9_P_btm.t95 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6755 VDAC_N.t336 C9_N_btm.t95 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6756 VDAC_P.t1248 C8_P_btm.t52 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6757 VDAC_P.t104 C10_P_btm.t179 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6758 VSS.t2002 a_n1085_47874# DATA[0].t1 VSS.t2001 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6759 VDD.t263 a_n1827_44324.t6 a_n2293_43244# VDD.t262 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6760 VDAC_N.t1256 C9_N_btm.t94 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6761 VSS.t3769 C10_N_btm.t1074 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6762 VDAC_N.t640 C10_N_btm.t175 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6763 VDD.t1826 a_18971_44654# a_18958_44350# VDD.t1825 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6764 a_16885_46232# a_9521_45982.t8 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.14825 ps=1.34 w=0.42 l=0.15
X6765 VDAC_P.t1240 C8_P_btm.t50 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6766 VDAC_P.t632 C10_P_btm.t178 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6767 VDD.t2562 VSS.t3614 VDD.t2561 VDD.t2366 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6768 VDAC_N.t1248 C10_N_btm.t174 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6769 VDAC_P.t1232 C9_P_btm.t91 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6770 VSS.t371 a_n2442_44894.t6 C9_P_btm.t2 VSS.t370 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X6771 VDAC_P.t328 C9_P_btm.t92 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6772 a_8192_44874# a_8423_42718# VSS.t1216 VSS.t1215 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X6773 a_750_46892# a_135_43540.t17 VSS.t2742 VSS.t2741 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X6774 a_2424_46794.t1 a_11059_45956# VDD.t1014 VDD.t1013 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X6775 VDAC_P.t1224 C10_P_btm.t177 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6776 VDAC_N.t104 C7_N_btm.t26 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6777 VSS.t2464 VSS.t2465 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6778 VDAC_N.t1240 C7_N_btm.t113 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6779 VDAC_N.t632 C6_N_btm.t51 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6780 VDD.t1031 a_21197_42718# a_18766_43236# VDD.t1030 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6781 VDAC_P.t624 C7_P_btm.t28 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6782 VDAC_N.t1232 C10_N_btm.t173 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6783 VDAC_N.t328 C9_N_btm.t93 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6784 VDAC_N.t1224 C9_N_btm.t92 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6785 VSS.t1121 a_15005_47222# a_10199_47846.t0 VSS.t1120 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6786 VDAC_P.t1216 C8_P_btm.t49 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6787 VDAC_P.t176 C8_P_btm.t44 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6788 VREF.t52 a_20647_31459.t4 C5_N_btm.t36 VDD.t2976 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X6789 VDAC_P.t1208 C9_P_btm.t90 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6790 VDAC_P.t616 C10_P_btm.t176 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6791 a_3165_43262# a_2627_43262# VSS.t1101 VSS.t1100 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X6792 VSS.t3398 VDD.t3190 VSS.t3397 VSS.t3201 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6793 VDAC_P.t1200 C9_P_btm.t89 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6794 VDAC_N.t624 C9_N_btm.t91 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6795 VSS.t2783 a_n2293_45420.t6 a_21719_43244# VSS.t2782 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6796 a_19358_43582# a_1581_43806.t16 a_19191_43262# VSS.t2957 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X6797 VDAC_N.t1216 C10_N_btm.t172 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6798 a_5088_37509.t7 VDAC_P.t320 a_8912_37509.t25 VDD.t2241 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X6799 VSS.t2347 VSS.t2348 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6800 VDAC_P.t1192 C10_P_btm.t175 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6801 a_n1890_47614.t2 a_n1920_47588# VDD.t2775 VDD.t2774 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X6802 VDAC_P.t608 C10_P_btm.t174 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6803 VDAC_N.t176 C10_N_btm.t171 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6804 VSS.t2335 VSS.t2336 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6805 VDAC_N.t1208 C10_N_btm.t170 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6806 VDD.t790 a_10884_45982# a_11059_45956# VDD.t789 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X6807 VDAC_P.t1184 C10_P_btm.t173 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6808 a_12991_43640# a_12545_43268# a_12895_43640# VSS.t870 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X6809 VDAC_N.t616 C10_N_btm.t169 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6810 VDAC_N.t1200 C10_N_btm.t168 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6811 VDAC_N.t320 C10_N_btm.t167 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6812 a_n61_43262# a_135_43540.t35 VDD.t186 VDD.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X6813 VSS.t1173 a_18135_47588# a_13524_46832.t0 VSS.t1172 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X6814 VDAC_P.t64 C10_P_btm.t172 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6815 VSS.t262 a_2587_44868.t21 a_4997_44670# VSS.t261 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X6816 VDAC_P.t1176 C9_P_btm.t88 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6817 VDAC_N.t1192 C8_N_btm.t42 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6818 VDAC_P.t600 C9_P_btm.t87 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6819 VDAC_P.t1168 C9_P_btm.t86 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6820 VSS.t1457 a_2655_42870# a_2627_42718# VSS.t1456 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X6821 a_2134_44324# a_1736_43276# VSS.t1198 VSS.t1197 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.11975 ps=1.045 w=0.42 l=0.15
X6822 VDAC_N.t608 C10_N_btm.t166 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6823 VDAC_P.t312 C10_P_btm.t171 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6824 a_7705_45736# a_7372_45670# VDD.t678 VDD.t677 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X6825 a_13097_46348# a_13248_45956.t20 a_13181_45982# VDD.t408 sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6826 VIN_P.t2 EN_VIN_BSTR_P.t20 C5_P_btm.t1 VSS.t561 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X6827 a_13457_46892# a_13427_46756# a_13373_46892# VSS.t1524 sky130_fd_pr__nfet_01v8 ad=0.085225 pd=0.925 as=0.0567 ps=0.69 w=0.42 l=0.15
X6828 VSS.t1308 a_12623_43780# a_10259_42870.t1 VSS.t1307 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X6829 VREF.t48 a_21276_30659.t5 C8_N_btm.t273 VDD.t2931 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6830 VDAC_N.t1184 C9_N_btm.t90 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6831 a_3895_43262# a_135_43540.t45 VDD.t192 VDD.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X6832 VDAC_N.t64 C6_N_btm.t26 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6833 a_14545_44133# a_n1067_42718.t4 a_14331_44133# VDD.t269 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X6834 a_11991_44172# a_10227_47214.t18 VDD.t291 VDD.t290 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X6835 a_n2074_47070.t3 a_n2104_47044# VDD.t664 VDD.t663 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X6836 a_14297_32299.t2 a_22959_43270# VDD.t1383 VDD.t1382 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X6837 a_12732_45144# a_12684_45276# a_12648_45144# VDD.t1010 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6838 VDAC_N.t1176 C7_N_btm.t83 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6839 a_n1735_43236.t7 a_2134_44324# VDD.t1739 VDD.t1738 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6840 VDAC_N.t600 C10_N_btm.t165 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6841 VDAC_N.t1168 C6_N_btm.t10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6842 VDAC_P.t1160 C8_P_btm.t43 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6843 VDAC_N.t312 C9_N_btm.t89 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6844 VDAC_P.t592 C8_P_btm.t42 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6845 VDAC_N.t1160 C9_N_btm.t88 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6846 VDAC_P.t1152 C10_P_btm.t170 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6847 VSS.t2886 a_12651_44576.t26 a_16868_44670# VSS.t2885 sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.08775 ps=0.92 w=0.65 l=0.15
X6848 VDD.t1172 a_7595_47614# DATA[5].t7 VDD.t1171 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6849 VDAC_N.t592 C9_N_btm.t87 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6850 VDD.t2011 a_1488_43236# a_n2661_45420.t3 VDD.t2010 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X6851 VSS.t3783 C9_P_btm.t21 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6852 VDAC_N.t1152 C10_N_btm.t164 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6853 C10_N_btm.t20 a_22812_30659.t6 VREF.t31 VDD.t518 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6854 VDD.t1842 a_13023_42718# a_5334_30651.t2 VDD.t1841 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X6855 VDAC_P.t168 C10_P_btm.t169 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6856 VDD.t1720 a_1239_39587# COMP_P.t5 VDD.t1719 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6857 VDAC_P.t1144 C7_P_btm.t27 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6858 VDAC_N.t168 C9_N_btm.t86 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6859 VDAC_N.t1144 C10_N_btm.t163 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6860 VDAC_Ni.t6 a_3754_38470.t4 a_3726_37500# VSS.t2838 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X6861 a_8912_37509.t9 VDAC_N.t584 a_5700_37509.t3 VDD.t2245 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X6862 VDAC_P.t584 C10_P_btm.t168 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6863 VDAC_N.t1136 C10_N_btm.t162 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6864 VDAC_N.t304 C9_N_btm.t85 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6865 VDAC_N.t1128 C8_N_btm.t40 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6866 VDAC_N.t576 C9_N_btm.t84 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6867 a_15468_45412# a_13715_43780# a_15860_45438# VDD.t1196 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X6868 VDAC_N.t1120 VSS.t3265 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6869 a_22780_41381# COMP_P.t11 a_22521_41035# VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6870 a_18918_45758# a_18970_45412# a_n2103_45412.t2 VSS.t2026 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6871 VDAC_P.t1136 C9_P_btm.t85 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6872 VDAC_P.t304 C10_P_btm.t167 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6873 VSS.t3416 VDD.t3196 VSS.t3415 VSS.t3414 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X6874 VSS.t801 a_16291_46758# a_16128_46134# VSS.t800 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.17875 ps=1.85 w=0.65 l=0.15
X6875 VDAC_N.t96 C10_N_btm.t161 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6876 VDD.t709 a_15443_44582# a_15415_44350# VDD.t708 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X6877 a_5129_45956# a_885_44868.t19 VDD.t2840 VDD.t2839 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X6878 VDAC_P.t1128 C10_P_btm.t166 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6879 VDAC_P.t576 C10_P_btm.t165 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6880 VDAC_P.t1120 C9_P_btm.t84 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6881 a_3089_42718# a_2755_43494.t6 a_2655_42870# VSS.t506 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X6882 VDAC_P.t96 C10_P_btm.t164 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6883 VSS.t3791 C3_N_btm.t10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6884 VSS.t2337 VSS.t2338 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6885 VDAC_N.t1112 C10_N_btm.t160 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6886 a_4993_47044# a_4322_46134# VSS.t1828 VSS.t1827 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6887 VDAC_N.t568 C8_N_btm.t39 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6888 VDAC_N.t1104 C10_N_btm.t159 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6889 VDAC_P.t1112 C7_P_btm.t119 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6890 VDAC_N.t296 C10_N_btm.t158 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6891 VDAC_P.t568 C10_P_btm.t163 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6892 VDAC_N.t1096 C9_N_btm.t83 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6893 VDAC_P.t1104 C10_P_btm.t162 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6894 a_1387_44582# a_1659_44440# a_1617_44466# VDD.t1116 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6895 VDAC_P.t296 C10_P_btm.t161 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6896 VDAC_P.t1096 C8_P_btm.t40 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6897 a_18879_43780# a_18704_43806# a_19058_43806# VSS.t1133 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X6898 a_2587_44868.t5 a_20107_43806# VDD.t140 VDD.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X6899 VDAC_N.t560 C8_N_btm.t38 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6900 VDAC_P.t560 C10_P_btm.t160 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6901 VDAC_P.t1088 C10_P_btm.t159 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6902 VDAC_P.t160 C9_P_btm.t83 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6903 a_10224_45982# a_9973_46526# VDD.t809 VDD.t808 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X6904 VDAC_P.t2132 C10_P_btm.t158 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6905 a_1209_47588# a_1083_45221# VSS.t893 VSS.t892 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X6906 VSS.t3432 VDD.t3202 VSS.t3431 VSS.t3033 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X6907 VDAC_N.t1088 C10_N_btm.t157 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6908 VDAC_P.t1076 C7_P_btm.t98 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6909 DATA[5].t1 a_7595_47614# VSS.t1230 VSS.t1229 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6910 VDAC_N.t160 C10_N_btm.t156 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6911 VDD.t2368 VSS.t3799 VDD.t2367 VDD.t2366 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X6912 VDD.t1323 a_2343_47070# a_2351_47614# VDD.t1322 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X6913 VDD.t604 a_3222_30651.t14 a_21027_42718# VDD.t603 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X6914 a_2801_42968# a_2587_44868.t19 VDD.t241 VDD.t240 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X6915 VDD.t353 a_n690_43494.t9 a_n685_43268# VDD.t352 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6916 VDAC_N.t2132 C10_N_btm.t155 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6917 a_18093_43262# a_15549_47044.t5 a_18348_43262# VDD.t2985 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6918 a_8848_44868# a_8699_44894# VSS.t848 VSS.t847 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6919 VDAC_N.t1076 C10_N_btm.t154 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6920 a_19437_31459.t0 a_22959_44894# VSS.t2630 VSS.t1124 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X6921 a_1083_45221# a_636_42870# a_1083_44894# VSS.t821 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X6922 a_9350_43301# a_9304_43494# VDD.t650 VDD.t649 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X6923 VDAC_N.t2116 C8_N_btm.t37 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6924 VDD.t776 a_14133_43780# a_14545_44133# VDD.t775 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X6925 a_n2810_45438.t2 a_n2840_45412# VDD.t2068 VDD.t1303 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X6926 a_847_45956# a_672_45982# a_1026_45982# VSS.t2187 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X6927 VDD.t707 a_7961_44048# a_7851_44172# VDD.t706 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X6928 VDAC_N.t548 C10_N_btm.t153 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6929 VDAC_P.t2116 C10_P_btm.t157 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6930 VDAC_P.t548 C10_P_btm.t156 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6931 a_4049_46892# a_4005_46500# a_3883_46904# VSS.t2156 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X6932 VDAC_Pi.t8 a_7754_39632# VSS.t693 sky130_fd_pr__res_high_po_0p35 l=18
X6933 a_15389_47730# a_13524_46832.t20 a_15317_47730# VDD.t553 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6934 VDAC_P.t2100 C7_P_btm.t69 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6935 VDAC_N.t2100 C10_N_btm.t152 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6936 a_n2442_43806.t1 a_n2472_43780# VSS.t804 VSS.t803 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X6937 VDAC_N.t1060 C10_N_btm.t151 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6938 VDAC_P.t1060 C10_P_btm.t155 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6939 VREF.t4 a_19437_31459.t4 C0_N_btm.t0 VDD.t143 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X6940 VDAC_N.t2084 C10_N_btm.t150 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6941 VDAC_N.t36 C10_N_btm.t149 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6942 VDAC_N.t2068 C8_N_btm.t36 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6943 VDAC_P.t2084 C10_P_btm.t154 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6944 VDD.t2765 a_1177_38525# a_1343_38525.t4 VDD.t2764 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6945 VDD.t1329 a_8483_46830# a_8470_46526# VDD.t1328 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6946 VDAC_P.t36 C10_P_btm.t153 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6947 VSS.t769 a_n2288_42692# EN_COMP.t0 VSS.t768 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X6948 VDAC_P.t2068 C8_P_btm.t36 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6949 VDAC_P.t1044 C10_P_btm.t152 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6950 VDAC_N.t1044 C10_N_btm.t148 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6951 VDAC_P.t2052 C8_P_btm.t37 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6952 a_22399_44894# a_n1741_47596.t9 VDD.t275 VDD.t274 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6953 VDAC_N.t2052 C7_N_btm.t54 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6954 a_7142_47397# a_885_44868.t23 VDD.t2844 VDD.t2843 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X6955 VDAC_N.t532 C10_N_btm.t147 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6956 VDAC_P.t532 C9_P_btm.t82 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6957 VDAC_N.t2036 C10_N_btm.t146 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6958 VSS.t1212 a_8391_47044# a_135_43540.t1 VSS.t1211 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X6959 VDAC_P.t2036 C10_P_btm.t72 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6960 VSS.t1521 a_22223_44358# a_14601_32299.t0 VSS.t1520 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X6961 a_885_44868.t11 a_4322_46134# VDD.t1780 VDD.t1779 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6962 VDAC_N.t1028 C10_N_btm.t145 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6963 VDAC_P.t1028 C10_P_btm.t150 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6964 VDD.t1874 a_7556_42692# a_5923_31099.t2 VDD.t1873 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X6965 a_12055_45982# a_n53_44363.t20 a_11692_46134# VSS.t624 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X6966 VDAC_N.t2020 C9_N_btm.t82 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6967 VDAC_P.t2020 C10_P_btm.t149 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6968 VSS.t3802 C5_P_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6969 VDD.t727 a_22521_41035# a_22469_41061# VDD.t726 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6970 a_18247_44172# a_17623_43806# a_18139_43806# VDD.t1886 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X6971 a_20049_43262# a_19771_43600# VDD.t1919 VDD.t1918 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X6972 VDD.t441 a_7754_40130.t6 a_11206_38545.t1 VDD.t440 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X6973 a_7754_40130.t3 RST_Z.t5 VDD.t2920 VDD.t2919 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X6974 VDD.t18 a_10259_42870.t26 a_10215_44874# VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6975 VDAC_P.t276 C10_P_btm.t148 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6976 VDAC_N.t276 C10_N_btm.t144 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6977 VDAC_N.t2004 C10_N_btm.t142 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6978 VSS.t3681 C10_P_btm.t15 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6979 a_2385_45438# a_885_44868.t35 a_2301_45438# VDD.t2855 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X6980 VDAC_N.t1012 C10_N_btm.t141 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6981 VDAC_P.t2004 C9_P_btm.t81 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6982 VSS.t2232 a_5655_43780# a_8005_43806# VSS.t2231 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6983 a_6259_45804# a_5382_44582# a_5896_45670# VSS.t2074 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X6984 VDAC_N.t1988 C9_N_btm.t81 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6985 a_9571_43628# a_n53_44363.t23 a_9208_43494# VSS.t625 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X6986 VDAC_P.t1012 C9_P_btm.t80 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6987 VDAC_P.t1988 C9_P_btm.t79 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6988 VREF.t54 a_n4515_30659.t5 C10_P_btm.t1057 VDD.t2991 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X6989 VDAC_N.t516 C9_N_btm.t80 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6990 VDAC_P.t516 C10_P_btm.t146 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6991 VDAC_N.t1972 C10_N_btm.t140 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6992 VDAC_P.t1972 C10_P_btm.t145 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6993 a_10467_47212# a_9521_45982.t21 VSS.t41 VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6994 VDD.t1067 a_571_46830# a_558_46526# VDD.t1066 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X6995 a_9521_45982.t0 a_9343_45982# VSS.t1529 VSS.t1528 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X6996 VSS.t3805 C5_N_btm.t34 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6997 VDAC_P.t996 C10_P_btm.t144 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6998 VDAC_N.t996 C10_N_btm.t139 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X6999 VSS.t7 a_10259_42870.t14 a_12287_44894# VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X7000 VDAC_N.t1956 C10_N_btm.t138 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7001 VDAC_N.t148 VSS.t3294 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7002 w_11534_34010.t15 a_11730_34132.t6 w_11534_34010.t15 w_11534_34010.t13 sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X7003 VDAC_N.t1940 C10_N_btm.t137 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7004 VSS.t3448 VDD.t3208 VSS.t3447 VSS.t3446 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X7005 VDAC_N.t980 C10_N_btm.t136 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7006 a_7842_44868# a_5419_47258# VSS.t1589 VSS.t1588 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X7007 VDAC_N.t1924 C9_N_btm.t79 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7008 VSS.t2117 a_6391_46219# a_6322_46348# VSS.t2116 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X7009 VDAC_N.t500 C9_N_btm.t78 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7010 VDAC_P.t1956 C10_P_btm.t143 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7011 VDAC_N.t1908 C10_N_btm.t135 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7012 VCM.t8 a_3990_30651.t8 C10_N_btm.t11 VSS.t281 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7013 a_13991_42883# a_5334_30651.t5 VSS.t2934 VSS.t2933 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7014 VDAC_P.t148 C9_P_btm.t78 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7015 VDAC_P.t1940 C10_P_btm.t142 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7016 VDAC_P.t980 C10_P_btm.t141 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7017 a_9208_43494# a_n53_44363.t19 a_9350_43301# VDD.t563 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X7018 VDAC_P.t1924 C8_P_btm.t35 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7019 VDAC_P.t500 C10_P_btm.t140 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7020 VDAC_P.t1908 C8_P_btm.t268 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7021 VDAC_N.t964 C10_N_btm.t134 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7022 a_n73_43640# a_n519_43268# a_n169_43640# VSS.t1753 sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X7023 VDAC_N.t1892 C8_N_btm.t35 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7024 VDD.t2419 VSS.t3689 VDD.t2418 VDD.t2417 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7025 C10_P_btm.t1068 a_n4515_30659.t16 VREF.t65 VDD.t3002 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=0.35
X7026 a_n53_44363.t3 a_1115_47044# VDD.t1087 VDD.t1086 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7027 a_17053_46232# a_1429_47222.t17 a_16981_46232# VDD.t326 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7028 VDD.t1052 a_12833_42718# a_13023_42718# VDD.t1051 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7029 a_15962_47320# a_16102_47044# VDD.t1267 VDD.t1266 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7030 a_13654_46032# a_13248_45956.t24 a_13572_46032# VSS.t489 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7031 a_17927_46195# a_10251_45454# VSS.t1364 VSS.t1363 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7032 VDAC_N.t260 C9_N_btm.t77 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7033 VDAC_P.t964 C3_P_btm.t4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7034 VDAC_N.t1876 VSS.t3319 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7035 VDD.t1623 a_847_45956# a_834_46348# VDD.t1622 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X7036 VDAC_P.t1892 C10_P_btm.t138 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7037 a_781_45982# a_n409_45982# a_672_45982# VSS.t1036 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X7038 VDAC_P.t260 C7_P_btm.t57 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7039 a_15471_43806# a_15121_43806# a_15376_43806# VDD.t861 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7040 a_n2810_44350.t2 a_n2840_44324# VDD.t880 VDD.t879 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7041 VSS.t1600 a_22821_39429# a_22876_40293# VSS.t1599 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7042 a_16757_47070# a_16561_45982# a_15221_47044# VSS.t834 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7043 VDAC_P.t1876 C10_P_btm.t137 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7044 VSS.t3460 VDD.t3212 VSS.t3459 VSS.t3458 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X7045 VDAC_N.t948 C10_N_btm.t1051 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7046 VDAC_P.t948 C10_P_btm.t136 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7047 VDAC_N.t1860 C7_N_btm.t25 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7048 a_n2104_47044# a_n1925_47044.t7 VDD.t3075 VDD.t3074 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X7049 a_11795_47044# a_8727_47222.t14 VSS.t86 VSS.t85 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X7050 a_7000_47222# a_5663_45982# a_7142_47397# VDD.t2693 sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X7051 VDD.t859 a_5569_44048# a_5459_44172# VDD.t858 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X7052 VDAC_N.t484 C10_N_btm.t133 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7053 a_21997_47833# SMPL_ON_N.t9 VSS.t104 VSS.t103 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7054 VDAC_N.t1844 C10_N_btm.t132 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7055 VDAC_N.t932 C10_N_btm.t131 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7056 VDAC_P.t1860 C10_P_btm.t135 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7057 VDAC_N.t1828 C8_N_btm.t34 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7058 VDAC_N.t84 C10_N_btm.t130 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7059 VDAC_P.t484 C10_P_btm.t134 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7060 VSS.t1289 a_8659_44324# a_1053_45123.t0 VSS.t1288 sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X7061 VDAC_P.t1844 VSS.t3382 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7062 C9_N_btm.t7 a_21788_30659.t6 VREF.t25 VDD.t2053 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7063 VDAC_N.t1812 C9_N_btm.t76 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7064 VDAC_P.t932 C10_P_btm.t133 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7065 a_4091_47070# a_4061_47044# VDD.t1518 VDD.t1517 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7066 VDD.t2898 a_1847_45528.t27 a_3179_44403# VDD.t2897 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X7067 VDAC_N.t916 VSS.t3259 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7068 a_18103_46768# a_14950_43958# VDD.t1363 VDD.t1362 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7069 a_3895_43262# a_3271_43268# a_3787_43640# VDD.t2069 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X7070 VDD.t1337 a_18766_43236# a_18348_43262# VDD.t1336 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7071 VSS.t1431 a_14950_43958# a_14955_43806# VSS.t1430 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7072 VSS.t1585 a_n2840_43780# a_n2810_43806.t0 VSS.t943 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7073 VDAC_N.t1796 C7_N_btm.t21 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7074 C1_P_btm.t5 a_2252_42718.t4 VCM.t54 VSS.t364 sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X7075 a_18247_46348# a_10227_47214.t45 VDD.t576 VDD.t575 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X7076 VDAC_P.t1828 C10_P_btm.t132 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7077 VSS.t1383 a_n2833_47874# CLK_DATA.t0 VSS.t1382 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7078 DEBUG_OUT.t4 a_9863_47874# VDD.t1001 VDD.t1000 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X7079 VDAC_N.t468 C9_N_btm.t75 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7080 VSS.t3696 C4_P_btm.t4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7081 VDAC_P.t84 C9_P_btm.t77 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7082 a_7705_45736# a_7372_45670# VSS.t750 VSS.t749 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X7083 VDAC_N.t1780 C9_N_btm.t74 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7084 VDAC_P.t1812 C5_P_btm.t9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7085 VDAC_P.t916 C8_P_btm.t267 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7086 VDAC_N.t900 C10_N_btm.t129 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7087 a_5473_43582# a_4322_46134# VSS.t1824 VSS.t1823 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7088 a_20647_31459.t2 a_22223_47070# VDD.t2797 VDD.t968 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7089 VDD.t811 a_1204_46758# a_n447_47044# VDD.t810 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X7090 VSS.t523 a_n2293_47044.t4 a_22123_44894# VSS.t522 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7091 VDAC_P.t1796 VSS.t3390 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7092 VDAC_N.t1764 C9_N_btm.t73 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7093 VDAC_N.t244 C10_N_btm.t128 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7094 VSS.t3697 C10_P_btm.t27 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7095 a_7311_47614# a_6951_47070# VDD.t1550 VDD.t1549 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7096 VDAC_P.t468 C9_P_btm.t76 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7097 VDAC_P.t1780 C10_P_btm.t131 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7098 VSS.t3203 VDD.t3170 VSS.t3202 VSS.t3201 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7099 VDAC_N.t1748 C10_N_btm.t127 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7100 VDAC_P.t900 C8_P_btm.t34 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7101 VDAC_P.t1764 C10_P_btm.t130 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7102 a_1581_43806.t4 a_1123_43780# VDD.t1556 VDD.t1555 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7103 VDAC_P.t244 C9_P_btm.t75 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7104 VDAC_P.t1748 C10_P_btm.t129 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7105 VDAC_P.t884 C9_P_btm.t74 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7106 VDAC_N.t884 C10_N_btm.t126 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7107 VDD.t627 a_18259_46500# a_18190_46526# VDD.t626 sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X7108 a_104_42692# a_283_42692# VSS.t1027 VSS.t1026 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7109 a_93_43628# a_49_43236# a_n73_43640# VSS.t1762 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X7110 a_2165_46224# a_1947_45982# VDD.t3090 VDD.t3089 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X7111 VDAC_N.t1732 C10_N_btm.t125 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7112 VDD.t222 a_7557_43236.t20 a_10447_44403# VDD.t221 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X7113 VDAC_N.t452 C10_N_btm.t124 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7114 VDAC_N.t1716 C10_N_btm.t123 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7115 VDAC_P.t1732 C9_P_btm.t73 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7116 VDAC_P.t452 C10_P_btm.t128 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7117 a_18449_44324# a_18231_44728# VSS.t978 VSS.t977 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X7118 VDAC_P.t1716 C10_P_btm.t127 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7119 a_12386_45758# a_12438_45412# a_n1551_45412.t0 VSS.t814 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7120 VSS.t65 a_1343_38525.t8 a_2113_38308# VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X7121 VDAC_N.t868 C9_N_btm.t72 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7122 VDAC_P.t868 C10_P_btm.t126 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7123 VDAC_N.t1700 C8_N_btm.t33 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7124 VDAC_N.t132 C10_N_btm.t122 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7125 VDD.t461 a_7754_40130.t15 a_8912_37509.t5 VDD.t460 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X7126 a_10227_47214.t1 a_11795_47044# VSS.t2651 VSS.t2650 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X7127 a_3897_45444# a_3731_45444# VDD.t2115 VDD.t2114 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7128 VDAC_N.t1684 C8_N_btm.t253 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7129 a_n2810_45982.t0 a_n2840_45956# VSS.t1657 VSS.t1656 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7130 VDAC_P.t1700 C9_P_btm.t72 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7131 VSS.t1996 a_7016_46231# a_6954_46348# VSS.t1995 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X7132 VIN_P.t7 EN_VIN_BSTR_P.t22 C2_P_btm.t2 VSS.t562 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X7133 C0_P_btm.t5 a_n1522_42718.t4 VSS.t23 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X7134 VDD.t1572 a_18879_43780# a_13273_44868.t5 VDD.t1571 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7135 a_n1925_47044.t2 a_8848_44868# VDD.t2717 VDD.t2716 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X7136 a_17515_43806# a_17242_43806# VDD.t1321 VDD.t1320 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7137 VSS.t3493 VDD.t3224 VSS.t3492 VSS.t3491 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X7138 a_15040_45798# a_14853_45438# a_14953_45554# VSS.t813 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X7139 a_16404_43640# a_15323_43268# a_16057_43236# VDD.t1370 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X7140 DEBUG_OUT.t2 a_9863_47874# VSS.t1061 VSS.t1060 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X7141 VDAC_N.t852 C8_N_btm.t31 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7142 VSS.t2277 VSS.t2278 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7143 a_4733_44670# a_1847_45528.t11 VSS.t168 VSS.t167 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7144 VDAC_N.t1668 C7_N_btm.t22 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7145 VDAC_N.t436 C10_N_btm.t121 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7146 VDAC_P.t132 C7_P_btm.t52 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7147 a_1488_43236# a_1339_43315# VSS.t2176 VSS.t2175 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7148 VDD.t493 a_15730_45670.t16 a_16651_46500# VDD.t492 sky130_fd_pr__pfet_01v8_hvt ad=0.1226 pd=1.32 as=0.1176 ps=1.4 w=0.42 l=0.15
X7149 VDAC_N.t1652 C8_N_btm.t30 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7150 VDAC_P.t1684 C8_P_btm.t33 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7151 VDAC_P.t852 C6_P_btm.t15 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7152 VDAC_N.t836 C4_N_btm.t5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7153 VDD.t759 a_636_42870# a_n1459_43236.t3 VDD.t758 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7154 a_n2109_42692.t0 a_15187_44868# a_15133_45144# VDD.t1206 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7155 VDAC_P.t1668 C8_P_btm.t32 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7156 a_12379_44350# a_2755_43494.t15 a_12461_44670# VSS.t513 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X7157 VDAC_N.t1636 C10_N_btm.t120 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7158 SMPL.t3 a_n2833_42692# VSS.t986 VSS.t985 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X7159 VDAC_P.t436 C9_P_btm.t71 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7160 VDAC_P.t1652 VSS.t3393 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7161 a_16036_43806# a_14955_43806# a_15689_44048# VDD.t1880 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X7162 VDD.t1158 a_1663_45046# a_380_47222# VDD.t1157 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X7163 a_21908_43236# a_22087_43244# VSS.t1348 VSS.t1347 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7164 a_n2104_47044# a_n1925_47044.t9 VSS.t2978 VSS.t2977 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7165 VCM.t57 a_4758_30651.t6 C9_P_btm.t538 VSS.t2987 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7166 VDAC_N.t228 C8_N_btm.t29 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7167 VDAC_P.t836 C10_P_btm.t125 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7168 VDD.t1766 a_12896_47044# a_n2661_47044.t2 VDD.t1765 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X7169 VDAC_P.t1636 C10_P_btm.t124 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7170 VDAC_P.t228 C9_P_btm.t69 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7171 VDAC_N.t1620 C10_N_btm.t1032 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7172 VDAC_N.t820 C10_N_btm.t993 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7173 VSS.t3144 VDD.t3150 VSS.t3143 VSS.t3142 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X7174 VDAC_N.t1604 C9_N_btm.t71 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7175 VDAC_N.t420 C10_N_btm.t774 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7176 VDD.t2516 VSS.t3710 VDD.t2515 VDD.t2514 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X7177 VDAC_P.t1620 C10_P_btm.t123 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7178 a_9973_46526# a_9547_46565# VSS.t2608 VSS.t2607 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X7179 VDAC_P.t820 C10_P_btm.t122 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7180 VDAC_P.t1604 C9_P_btm.t68 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7181 VDAC_P.t420 C10_P_btm.t121 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7182 a_6953_43582# a_2755_43494.t4 a_6519_43494# VSS.t504 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7183 a_n169_43640# a_n685_43268# a_n264_43628# VSS.t2262 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X7184 VDAC_N.t1588 C10_N_btm.t599 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7185 VSS.t3636 C10_N_btm.t1075 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7186 VDAC_N.t804 C10_N_btm.t500 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7187 VDAC_P.t1588 C10_P_btm.t120 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7188 a_13930_46842# a_14470_46526# a_14658_46526# VDD.t3088 sky130_fd_pr__pfet_01v8_hvt ad=0.2688 pd=2.12 as=0.092075 ps=0.99 w=0.42 l=0.15
X7189 VSS.t3499 VDD.t3226 VSS.t3498 VSS.t3497 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7190 VSS.t3280 a_n2810_44894.t8 C10_P_btm.t1076 VSS.t3279 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7191 w_11534_34010.t3 a_18394_35068.t10 EN_VIN_BSTR_N.t1 w_11534_34010.t2 sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X7192 VDAC_N.t1572 C9_N_btm.t70 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7193 VDAC_P.t804 C9_P_btm.t67 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7194 VDAC_N.t52 C9_N_btm.t69 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7195 VSS.t3225 VDD.t3178 VSS.t3224 VSS.t3223 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X7196 VDAC_P.t1572 C9_P_btm.t66 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7197 VDAC_P.t52 C8_P_btm.t31 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7198 a_1597_45982# a_1431_45982# VSS.t757 VSS.t756 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7199 a_7195_44868# a_7020_44894# a_7374_44894# VSS.t785 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X7200 VDD.t457 a_7754_40130.t13 a_3754_38470.t1 VDD.t456 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X7201 a_22609_38426# a_22469_39973# CAL_P.t1 VSS.t2592 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X7202 VDD.t1361 a_14950_43958# a_14955_43806# VDD.t1360 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7203 VDAC_N.t1556 C7_N_btm.t20 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7204 VDAC_N.t788 C10_N_btm.t492 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7205 VDAC_P.t1556 C10_P_btm.t967 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7206 VSS.t503 a_n237_45454.t21 a_n107_47098# VSS.t502 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X7207 VSS.t1761 a_22959_47622# a_22812_30659.t1 VSS.t1760 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7208 VDAC_P.t788 C9_P_btm.t65 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7209 a_9547_46892# a_9293_46565# VSS.t3002 VSS.t3001 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X7210 VDAC_N.t1540 C5_N_btm.t6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7211 VDAC_P.t1540 C7_P_btm.t49 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7212 a_19520_46500# a_19371_46579# VSS.t1091 VSS.t1090 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7213 VDAC_N.t404 C10_N_btm.t485 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7214 a_15329_47044# a_15879_47320# VDD.t1341 VDD.t1340 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7215 VDAC_N.t1524 C9_N_btm.t68 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7216 VDAC_N.t772 C9_N_btm.t67 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7217 VDAC_N.t1508 C8_N_btm.t28 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7218 VDAC_P.t404 C9_P_btm.t64 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7219 VDAC_P.t1524 C7_P_btm.t25 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7220 a_5832_44466# a_5784_44364# a_5748_44466# VDD.t918 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7221 a_16576_44868# a_16427_44894# a_16872_45144# VDD.t2007 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7222 VDAC_P.t772 C9_P_btm.t63 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7223 VDAC_N.t212 C10_N_btm.t475 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7224 VDD.t870 a_22223_42718# a_22400_42718# VDD.t665 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7225 VDAC_N.t1492 C10_N_btm.t468 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7226 VDAC_N.t756 C10_N_btm.t244 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7227 a_15008_42692# a_15133_43582# VDD.t1191 VDD.t474 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X7228 VDAC_P.t1508 C10_P_btm.t770 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7229 VDD.t1325 a_16404_43640# a_16579_43566# VDD.t1324 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X7230 VSS.t873 a_22276_45412# a_18314_32299.t1 VSS.t872 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7231 VSS.t2426 VSS.t2427 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7232 VDAC_N.t1476 C10_N_btm.t241 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7233 VDAC_P.t212 C9_P_btm.t62 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7234 VDD.t551 a_13524_46832.t15 a_14219_47070# VDD.t550 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X7235 VDAC_P.t1492 C10_P_btm.t631 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7236 VDAC_P.t756 C9_P_btm.t61 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7237 VDAC_N.t388 C10_N_btm.t236 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7238 VDAC_N.t1460 C10_N_btm.t233 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7239 VDAC_N.t740 C9_N_btm.t66 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7240 VDD.t2154 a_672_45982# a_847_45956# VDD.t2153 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X7241 VDAC_P.t1476 C10_P_btm.t512 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7242 a_21719_43244# a_n2293_45420.t9 VSS.t2787 VSS.t2786 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7243 VDAC_P.t6 a_3222_30651.t17 VCM.t36 VSS.t668 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7244 SMPL.t5 a_n2833_42692# VDD.t932 VDD.t931 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X7245 VDAC_P.t1460 C10_P_btm.t498 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7246 VSS.t884 a_20064_35138# a_21789_35634# VSS.t883 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7247 VDD.t1496 a_16036_43806# a_16211_43780# VDD.t1495 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X7248 VDAC_P.t740 C4_P_btm.t10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7249 C10_P_btm.t1064 a_n4515_30659.t12 VREF.t61 VDD.t2998 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7250 VDAC_P.t1444 C9_P_btm.t60 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7251 a_11455_44576.t2 a_13635_43566# VSS.t1248 VSS.t1247 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7252 VSS.t2890 a_15549_47044.t6 a_15468_45412# VSS.t2889 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X7253 a_6360_44894# a_6243_45107# VDD.t1974 VDD.t1973 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X7254 VDAC_N.t1444 C7_N_btm.t19 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7255 C8_P_btm.t1 a_n2810_47070.t5 VREF.t1 VDD.t87 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7256 VDAC_N.t116 C7_N_btm.t18 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7257 VDAC_N.t1428 C10_N_btm.t229 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7258 VDAC_P.t116 C6_P_btm.t14 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7259 a_10259_42870.t0 a_12623_43780# VSS.t1310 VSS.t1309 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7260 VDD.t1470 a_7842_44868# a_n2293_46508.t2 VDD.t1469 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X7261 VDAC_N.t724 C8_N_btm.t242 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7262 VDAC_P.t1428 C8_P_btm.t30 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7263 VDAC_P.t724 C8_P_btm.t29 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7264 VDAC_N.t1412 C9_N_btm.t516 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7265 VDAC_P.t1412 C8_P_btm.t28 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7266 a_n1435_47614.t0 a_n1605_47614# VSS.t686 VSS.t685 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7267 VDAC_N.t372 VSS.t3305 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7268 VDD.t2668 a_10414_43780# a_n1551_44324.t5 VDD.t2667 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7269 VDD.t662 a_n2104_47044# a_n2074_47070.t2 VDD.t661 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X7270 VDD.t2190 a_1431_47070# a_1203_42692.t6 VDD.t2189 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7271 VDAC_N.t1396 C10_N_btm.t226 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7272 a_12461_44350# a_12651_44576.t14 VDD.t2962 VDD.t2961 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X7273 a_12648_45144# a_2424_46794.t6 VDD.t2944 VDD.t2943 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X7274 VDAC_N.t708 C9_N_btm.t65 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7275 VDAC_N.t7 a_3222_30651.t21 VCM.t33 VSS.t673 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7276 VDAC_P.t372 C10_P_btm.t483 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7277 VDAC_P.t1396 C10_P_btm.t473 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7278 VSS.t2034 a_17671_42883# a_16824_45276# VSS.t2033 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X7279 VDAC_P.t708 C10_P_btm.t246 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7280 VDD.t2609 VSS.t3816 VDD.t2608 VDD.t2607 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X7281 VDAC_N.t196 C10_N_btm.t219 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7282 VDAC_P.t1380 C9_P_btm.t59 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7283 CAL_N.t2 a_22465_38541# VDD.t2793 VDD.t2792 sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X7284 VDD.t251 a_2587_44868.t31 a_885_44868.t1 VDD.t250 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7285 VREF.t63 a_n4515_30659.t14 C10_P_btm.t1066 VDD.t3000 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7286 C9_N_btm.t540 a_4758_30651.t10 VCM.t61 VSS.t2991 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7287 VDAC_N.t1364 C9_N_btm.t63 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7288 a_n2661_45420.t2 a_1488_43236# VDD.t2009 VDD.t2008 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X7289 VDAC_N.t692 C9_N_btm.t62 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7290 VDD.t2627 VSS.t3733 VDD.t2626 VDD.t2625 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X7291 a_13013_44894# a_4322_46134# a_12931_44894# VSS.t1832 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X7292 VDD.t218 a_7557_43236.t16 a_n1551_44324.t1 VDD.t217 sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.135 ps=1.27 w=1 l=0.15
X7293 VDD.t299 a_10227_47214.t25 a_10768_47436# VDD.t298 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X7294 VSS.t2697 a_15008_42692# a_5142_30651.t0 VSS.t2696 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7295 VDAC_N.t1348 C9_N_btm.t61 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7296 VDAC_P.t196 C7_P_btm.t24 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7297 VDAC_N.t356 C9_N_btm.t60 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7298 VDAC_P.t1364 C3_P_btm.t7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7299 VDD.t1273 a_4987_45742# a_4974_45438# VDD.t1272 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X7300 VDAC_P.t692 C9_P_btm.t58 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7301 VDD.t459 a_7754_40130.t14 a_8912_37509.t4 VDD.t458 sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X7302 a_17242_43806# a_15730_45670.t14 a_17156_43806# VSS.t570 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X7303 a_645_43806# a_601_44048# a_479_43806# VSS.t880 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X7304 VDD.t2289 VSS.t3585 VDD.t2288 VDD.t2287 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7305 a_n2840_43236# a_n2661_43244# VSS.t688 VSS.t687 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7306 VDAC_P.t1348 C6_P_btm.t13 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7307 VDAC_P.t356 C10_P_btm.t239 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7308 VDAC_N.t1332 C9_N_btm.t59 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7309 a_n2442_44894.t2 a_n2472_44868# VDD.t672 VDD.t671 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7310 VDAC_P.t1332 C10_P_btm.t234 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7311 VSS.t3735 C5_N_btm.t35 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7312 VSS.t2389 VSS.t2390 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7313 VDAC_P.t676 C9_P_btm.t57 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7314 VDAC_N.t676 C10_N_btm.t216 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7315 VDAC_N.t1316 C10_N_btm.t212 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7316 a_989_45736# a_656_45670# VDD.t965 VDD.t964 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X7317 VDAC_N.t68 C7_N_btm.t17 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7318 VDAC_N.t1300 C9_N_btm.t502 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7319 VDAC_N.t660 C10_N_btm.t119 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7320 VDAC_P.t1316 C7_P_btm.t20 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7321 VDD.t1345 a_4651_47614# DATA[3].t7 VDD.t1344 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7322 a_17789_45982# a_17623_45982# VDD.t1082 VDD.t1081 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7323 VDAC_N.t1284 C9_N_btm.t290 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7324 VDAC_P.t68 C10_P_btm.t231 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7325 VDAC_P.t1300 C10_P_btm.t227 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7326 VDAC_P.t660 C8_P_btm.t27 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7327 VDAC_P.t1284 C9_P_btm.t514 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7328 VDAC_P.t340 C10_P_btm.t224 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7329 VDAC_P.t1268 C9_P_btm.t399 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7330 VSS.t3737 C10_N_btm.t1076 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7331 VDAC_P.t644 C10_P_btm.t217 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7332 VSS.t2383 VSS.t2384 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7333 VDD.t309 a_n2661_45420.t8 a_21847_43806# VDD.t308 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7334 VDAC_N.t340 C10_N_btm.t115 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7335 a_672_45982# a_n243_45982# a_325_46224# VSS.t2226 sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7336 VDAC_N.t1268 C9_N_btm.t247 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7337 VDAC_N.t644 C9_N_btm.t240 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7338 VDAC_N.t1252 C10_N_btm.t113 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7339 DATA[5].t2 a_7595_47614# VSS.t1234 VSS.t1233 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X7340 VDAC_P.t1252 C10_P_btm.t214 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7341 a_11265_44350# a_11455_44576.t14 VDD.t2814 VDD.t2813 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X7342 VDD.t2460 VSS.t3738 VDD.t2459 VDD.t2458 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X7343 VDAC_N.t180 C10_N_btm.t112 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7344 VSS.t652 a_13273_44868.t28 a_19371_46579# VSS.t651 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X7345 VDAC_P.t180 C8_P_btm.t26 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7346 VDAC_P.t1236 C10_P_btm.t118 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7347 VDAC_N.t1236 C10_N_btm.t108 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7348 VDAC_P.t628 C9_P_btm.t300 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7349 a_18093_43262# a_13273_44868.t17 a_n2497_42870.t5 VDD.t589 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7350 VSS.t2323 VSS.t2324 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7351 VDAC_N.t628 C8_N_btm.t121 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7352 VDAC_P.t1220 C10_P_btm.t117 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7353 VDAC_N.t1220 C6_N_btm.t9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7354 a_2157_43262# a_1203_42692.t17 a_2075_42870# VDD.t479 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7355 VDAC_N.t324 C7_N_btm.t16 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7356 VSS.t350 a_10227_47214.t29 a_12145_43806# VSS.t349 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X7357 a_n519_43268# a_n685_43268# VDD.t2228 VDD.t2227 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7358 DEBUG_OUT.t5 a_9863_47874# VDD.t999 VDD.t998 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7359 VDAC_P.t324 C6_P_btm.t12 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7360 VDAC_N.t1204 C9_N_btm.t119 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7361 VDAC_P.t1204 C8_P_btm.t254 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7362 a_13738_46032# a_4322_46134# VSS.t1826 VSS.t1825 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7363 a_13214_45758# a_13266_45412# a_n1827_45412.t1 VSS.t969 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7364 VDAC_P.t612 C10_P_btm.t114 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7365 VDAC_N.t612 C3_N_btm.t9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7366 VDAC_P.t1188 C10_P_btm.t113 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7367 VDAC_N.t1188 C9_N_btm.t116 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7368 VDAC_N.t100 C8_N_btm.t57 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7369 VDAC_N.t1172 C10_N_btm.t107 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7370 VDAC_N.t596 C10_N_btm.t105 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7371 a_8483_43780# a_8308_43806# a_8662_43806# VSS.t1598 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X7372 a_n2103_45412.t4 a_7208_47044# VDD.t2705 VDD.t2704 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7373 VDAC_N.t1156 C8_N_btm.t54 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7374 VDAC_P.t100 VSS.t3372 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7375 VDAC_P.t1172 C8_P_btm.t192 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7376 VDAC_N.t308 C9_N_btm.t112 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7377 VDAC_P.t596 C9_P_btm.t259 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7378 VDD.t3049 SMPL.t14 a_18394_35068.t3 VDD.t3048 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7379 VSS.t3740 C10_P_btm.t14 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7380 VDAC_N.t1140 C9_N_btm.t109 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7381 VDD.t761 a_636_42870# a_2043_43958# VDD.t760 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X7382 VDAC_N.t580 C10_N_btm.t104 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7383 a_16111_45412# a_1581_43806.t20 VDD.t2913 VDD.t2912 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X7384 VDAC_N.t1124 C10_N_btm.t101 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7385 VDAC_P.t1156 C9_P_btm.t243 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7386 VSS.t806 a_n2472_43780# a_n2442_43806.t0 VSS.t805 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7387 VDAC_N.t164 C10_N_btm.t100 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7388 VDAC_P.t308 C10_P_btm.t111 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7389 VDAC_N.t1108 C8_N_btm.t25 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7390 VSS.t1214 a_8391_47044# a_135_43540.t0 VSS.t1213 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7391 a_15443_44582# a_13273_44868.t21 a_15589_44670# VSS.t644 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X7392 VDAC_P.t1140 C9_P_btm.t236 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7393 VDAC_P.t580 C9_P_btm.t228 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7394 VDAC_N.t564 C10_N_btm.t98 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7395 VDD.t959 a_19037_42718# a_22223_42718# VDD.t681 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7396 VDAC_P.t1124 C10_P_btm.t110 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7397 a_7415_44466# a_1429_47222.t13 VSS.t386 VSS.t385 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7398 VDAC_P.t164 C10_P_btm.t106 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7399 VDAC_N.t1092 C9_N_btm.t55 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7400 VDD.t1415 a_3699_43780# a_3686_44172# VDD.t1414 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X7401 DEBUG_OUT.t0 a_9863_47874# VSS.t1059 VSS.t1058 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7402 VDAC_N.t292 C6_N_btm.t8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7403 VDAC_N.t2124 C7_N_btm.t15 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7404 VDAC_P.t1108 C7_P_btm.t19 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7405 VDD.t1774 a_4322_46134# a_885_44868.t8 VDD.t1773 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7406 VDD.t1020 a_21997_47833# a_1651_47044.t1 VDD.t1019 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7407 a_5923_31099.t3 a_7556_42692# VDD.t1876 VDD.t1875 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7408 a_16555_46616# a_13248_45956.t11 VSS.t481 VSS.t480 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06195 ps=0.715 w=0.42 l=0.15
X7409 VDAC_N.t1068 C6_N_btm.t7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7410 VDAC_N.t2092 C9_N_btm.t54 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7411 VDAC_P.t564 C7_P_btm.t17 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7412 a_13207_46892# a_13524_46832.t17 a_13457_46892# VSS.t604 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.085225 ps=0.925 w=0.42 l=0.15
X7413 VDAC_N.t44 C10_N_btm.t97 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7414 a_7781_43582# a_2755_43494.t11 a_7347_43494# VSS.t509 sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7415 a_6717_44894# a_6673_45136# a_6551_44894# VSS.t865 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X7416 VDAC_P.t1092 C5_P_btm.t8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7417 VSS.t3650 C10_P_btm.t10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7418 VDAC_P.t292 C9_P_btm.t221 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7419 VDAC_P.t2124 C9_P_btm.t115 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7420 VDD.t591 a_13273_44868.t19 a_n2103_45412.t6 VDD.t590 sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.135 ps=1.27 w=1 l=0.15
X7421 VDAC_P.t1068 C8_P_btm.t131 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7422 a_1334_43494.t7 a_3699_43780# VDD.t1413 VDD.t1412 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7423 a_n2661_44868# a_n2103_45412.t10 VSS.t2789 VSS.t2788 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7424 a_22087_43244# a_n2293_45956.t5 VDD.t2952 VDD.t2951 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7425 VDAC_P.t2092 C9_P_btm.t112 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7426 VDAC_P.t44 C10_P_btm.t105 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7427 VDAC_P.t2060 C10_P_btm.t103 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7428 VSS.t3743 C4_N_btm.t21 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7429 VSS.t3516 VDD.t3232 VSS.t3515 VSS.t3514 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X7430 VDAC_N.t2060 C10_N_btm.t92 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7431 VDAC_N.t1036 C9_N_btm.t52 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7432 VDAC_N.t2028 C9_N_btm.t51 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7433 VDAC_P.t1036 C10_P_btm.t102 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7434 a_n1890_42718.t2 a_n1920_42692# VDD.t2164 VDD.t2163 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7435 VDAC_N.t524 C9_N_btm.t48 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7436 VDAC_N.t1996 C10_N_btm.t90 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7437 VDAC_N.t1004 C10_N_btm.t88 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7438 VDAC_P.t2028 C10_P_btm.t99 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7439 VDAC_P.t524 C10_P_btm.t98 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7440 a_9335_44324# a_9179_44592# a_9480_44350# VDD.t2737 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X7441 VDD.t1292 a_10251_45454# a_10111_45776# VDD.t1291 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X7442 VDAC_P.t1996 C10_P_btm.t96 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7443 VDAC_N.t1964 C10_N_btm.t87 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7444 a_17671_42883# a_4758_30651.t5 VDD.t3086 VDD.t3085 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7445 VDD.t958 a_9943_45046# a_9304_43494# VDD.t957 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X7446 C10_P_btm.t1073 a_n2810_44894.t5 VSS.t3274 VSS.t3273 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7447 a_558_46526# a_n519_46532# a_396_46904# VDD.t1074 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X7448 VDAC_P.t1004 VSS.t3350 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7449 VSS.t3749 C10_N_btm.t1077 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7450 VDAC_P.t1964 C10_P_btm.t91 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7451 VSS.t2846 a_n2103_44868.t9 a_22223_47622# VSS.t2845 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7452 VDD.t1302 a_n2840_44868# a_n2810_44894.t2 VDD.t1301 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X7453 VDAC_N.t268 VSS.t3299 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7454 VSS.t904 a_16703_42718# a_4758_30651.t1 VSS.t903 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7455 a_13814_43628# a_10227_47214.t43 VSS.t635 VSS.t634 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X7456 a_7851_44172# a_7227_43806# a_7743_43806# VDD.t953 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X7457 a_10581_45982# a_10537_46224# a_10415_45982# VSS.t849 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X7458 VREF.t46 a_22812_30659.t7 C10_N_btm.t21 VDD.t519 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7459 VDAC_N.t1932 C10_N_btm.t84 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7460 VDAC_N.t972 C6_N_btm.t6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7461 VSS.t972 a_6631_42883# a_5784_44364# VSS.t971 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X7462 VDD.t2481 VSS.t3753 VDD.t2480 VDD.t2479 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X7463 VDAC_N.t1900 C8_N_btm.t24 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7464 VDAC_P.t268 C7_P_btm.t16 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7465 a_9048_45758# a_6485_44582.t17 VSS.t2917 VSS.t2916 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7466 VDAC_P.t1932 C6_P_btm.t53 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7467 VSS.t3487 VDD.t3222 VSS.t3486 VSS.t3485 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X7468 VDAC_P.t972 C8_P_btm.t118 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7469 VDAC_P.t1900 C10_P_btm.t88 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7470 a_9768_46892# a_9517_46539# a_9547_46565# VSS.t1974 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7471 a_15415_46846# a_14766_45596.t5 a_15321_46846# VSS.t2798 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X7472 VDAC_P.t492 C9_P_btm.t108 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7473 VDAC_P.t1868 C10_P_btm.t85 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7474 VDD.t2217 a_5655_43780# a_9480_44350# VDD.t2216 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X7475 a_15005_47222# a_15437_47044# a_15155_47070# VSS.t712 sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X7476 a_22876_40293# a_22545_39429# a_22780_40293# VSS.t2125 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X7477 VDAC_N.t492 C10_N_btm.t82 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7478 VDD.t1119 a_10588_45670# a_10383_46697# VDD.t1118 sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X7479 VDAC_N.t1868 C10_N_btm.t81 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7480 a_18139_45982# a_17789_45982# a_18044_45982# VDD.t1430 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7481 VDAC_N.t940 C10_N_btm.t80 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7482 VDAC_N.t1836 C10_N_btm.t79 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7483 VDAC_N.t140 C10_N_btm.t78 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7484 VDAC_P.t940 C9_P_btm.t105 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7485 VDAC_N.t1804 C9_N_btm.t47 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7486 VDAC_P.t1836 C8_P_btm.t109 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7487 VDD.t745 a_14853_45438# a_14953_45554# VDD.t744 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X7488 a_12895_43640# a_12545_43268# a_12800_43628# VDD.t812 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7489 VDAC_N.t908 C10_N_btm.t77 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7490 a_n2442_46526.t3 a_n2472_46500# VDD.t1609 VDD.t1453 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X7491 VSS.t675 a_n1735_43236.t9 a_22959_45446# VSS.t674 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7492 VDAC_P.t140 C8_P_btm.t102 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7493 a_14103_46576# a_13427_46756# a_13930_46842# VDD.t1460 sky130_fd_pr__pfet_01v8_hvt ad=0.090125 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X7494 VDD.t506 a_15730_45670.t27 a_18348_43262# VDD.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7495 a_2151_45670# a_2535_45670# a_2301_45758# VSS.t1910 sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X7496 VSS.t1250 a_13635_43566# a_13569_43640# VSS.t1249 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X7497 VDAC_P.t1804 C9_P_btm.t100 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7498 a_8912_37509.t8 VDAC_N.t1772 a_5700_37509.t2 VDD.t2247 sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X7499 VDAC_P.t908 C10_P_btm.t86 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7500 VDAC_P.t1772 C9_P_btm.t97 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7501 VDAC_N.t460 C7_N_btm.t14 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7502 VSS.t1381 a_n2833_47874# CLK_DATA.t1 VSS.t1380 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X7503 VDAC_P.t460 C9_P_btm.t93 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7504 VDD.t2371 VSS.t3759 VDD.t2370 VDD.t2369 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X7505 VDD.t1480 a_21855_42718# a_13667_32299.t2 VDD.t1479 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7506 VDAC_P.t1740 C7_P_btm.t15 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7507 VDAC_N.t1740 C0_dummy_N_btm.t2 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7508 a_13561_44350# a_13023_44716# VSS.t1088 VSS.t1087 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X7509 VDAC_P.t876 C10_P_btm.t84 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7510 VDAC_N.t876 C7_N_btm.t13 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7511 VDAC_N.t1708 C10_N_btm.t76 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7512 a_18357_46224# a_18139_45982# VDD.t1425 VDD.t1424 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X7513 VDAC_N.t236 C8_N_btm.t22 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7514 VDAC_P.t1708 C7_P_btm.t14 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7515 VDAC_N.t1676 C9_N_btm.t45 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7516 VDD.t2356 VSS.t3613 VDD.t2355 VDD.t2354 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X7517 VDAC_P.t236 C9_P_btm.t56 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7518 VSS.t3761 C10_P_btm.t28 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7519 a_12_45982# a_n105_46195# VSS.t1988 VSS.t1987 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X7520 VDAC_P.t1676 C10_P_btm.t83 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7521 VDD.t2282 VSS.t3660 VDD.t2281 VDD.t2280 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X7522 VDAC_N.t844 C8_N_btm.t21 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7523 VDAC_P.t844 C10_P_btm.t82 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7524 a_15839_43640# a_15323_43268# a_15744_43628# VSS.t1438 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X7525 a_15376_43806# a_14757_43806# VSS.t1184 VSS.t1183 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X7526 VDAC_P.t1644 C9_P_btm.t51 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7527 a_n2661_43244# a_n2103_44324.t5 VSS.t3013 VSS.t2901 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7528 VDAC_P.t428 C9_P_btm.t50 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7529 VSS.t891 a_468_42870# a_428_42724# VSS.t890 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7530 VDAC_P.t1612 C10_P_btm.t81 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7531 VDAC_N.t1644 C10_N_btm.t75 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7532 VDAC_N.t428 C10_N_btm.t74 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7533 VDAC_N.t1612 C10_N_btm.t73 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7534 VDAC_P.t812 C10_P_btm.t80 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7535 VDAC_P.t1580 C10_P_btm.t79 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7536 VDAC_N.t812 C10_N_btm.t72 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7537 VDD.t2505 VSS.t3662 VDD.t2504 VDD.t2503 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X7538 VDD.t2543 VSS.t3767 VDD.t2542 VDD.t2541 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X7539 VDAC_N.t1580 C10_N_btm.t71 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7540 a_6665_43262# a_2755_43494.t13 a_6519_43494# VDD.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X7541 VDAC_N.t76 C10_N_btm.t70 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7542 VDAC_P.t76 C10_P_btm.t78 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7543 VSS.t1167 a_11427_43566# a_7557_43236.t3 VSS.t1166 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7544 VDAC_P.t1548 C9_P_btm.t48 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7545 VDAC_P.t780 C9_P_btm.t47 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7546 VDD.t2215 a_5655_43780# a_6536_46348# VDD.t2214 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X7547 a_20163_31459.t0 a_22223_46534# VSS.t1137 VSS.t1136 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X7548 a_n1551_45412.t1 a_12438_45412# a_12386_45758# VSS.t815 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7549 C0_dummy_P_btm.t0 EN_VIN_BSTR_P.t17 VIN_P.t3 VSS.t559 sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X7550 VSS.t2428 VSS.t2429 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7551 VDAC_P.t1516 C10_P_btm.t77 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7552 VSS.t308 a_17930_32299.t4 C9_N_btm.t0 VSS.t307 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7553 VDAC_P.t396 C10_P_btm.t76 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7554 VDAC_P.t1484 C10_P_btm.t75 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7555 a_n2103_44324.t0 a_8204_45412# VSS.t2161 VSS.t2160 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X7556 VDAC_N.t1548 C8_N_btm.t20 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7557 a_10245_46532# a_10079_46532# VSS.t2252 VSS.t2251 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7558 VDAC_N.t780 C6_N_btm.t5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7559 VDD.t2310 VSS.t3768 VDD.t2309 VDD.t2308 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X7560 VDAC_N.t1516 C10_N_btm.t69 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7561 VSS.t2440 VSS.t2441 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7562 a_5459_44172# a_4835_43806# a_5351_43806# VDD.t945 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X7563 VSS.t3063 VDD.t3123 VSS.t3062 VSS.t3061 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7564 VDAC_N.t396 C7_N_btm.t12 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7565 VDAC_N.t1484 C10_N_btm.t68 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7566 a_6235_46124# a_4830_43958.t11 VSS.t208 VSS.t207 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7567 VCM.t9 a_3990_30651.t9 C10_P_btm.t1 VSS.t282 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7568 SMPL.t1 a_n2833_42692# VSS.t984 VSS.t983 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7569 VDAC_N.t748 C9_N_btm.t44 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7570 VDAC_P.t748 C8_P_btm.t54 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7571 VDAC_N.t1452 C9_N_btm.t43 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7572 VDAC_P.t1452 C10_P_btm.t74 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7573 VDD.t102 a_927_42692.t19 a_12931_44894# VDD.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X7574 VDAC_P.t204 C10_P_btm.t73 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7575 VDAC_N.t204 C10_N_btm.t67 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7576 a_17721_45144# a_10251_45454# a_17531_44894# VDD.t1293 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.174 ps=1.39 w=1 l=0.15
X7577 a_13524_46832.t2 a_18135_47588# VDD.t1113 VDD.t683 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7578 VDAC_N.t1420 C10_N_btm.t66 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7579 VDAC_N.t716 C9_N_btm.t42 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7580 VSS.t2865 a_12651_44576.t13 a_12699_46616# VSS.t2864 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7581 a_6355_45477# a_6104_45706.t5 a_5896_45670# VDD.t3099 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X7582 VDAC_P.t1420 C8_P_btm.t51 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7583 VDAC_P.t716 C9_P_btm.t44 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7584 a_989_45736# a_656_45670# VSS.t1023 VSS.t1022 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X7585 VDAC_P.t1388 C10_P_btm.t43 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7586 VDD.t359 a_n690_43494.t13 a_3271_43268# VDD.t358 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7587 a_5896_45670# a_6104_45706.t11 a_6038_45804# VSS.t3011 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X7588 VSS.t3665 C9_N_btm.t536 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7589 a_8005_43806# a_7961_44048# a_7839_43806# VSS.t778 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X7590 VDAC_N.t1388 C10_N_btm.t65 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7591 VDAC_P.t364 C10_P_btm.t71 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7592 a_2684_37794# a_1736_39587.t5 a_1736_39043.t1 VSS.t2932 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X7593 a_n2661_47044.t3 a_12896_47044# VDD.t1768 VDD.t1767 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X7594 a_11047_45477# a_10389_45438# a_10588_45670# VDD.t793 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X7595 VDAC_N.t364 C10_N_btm.t64 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7596 a_n2472_43236# a_n2293_43244# VSS.t1694 VSS.t1205 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X7597 a_5728_46526# a_4322_46134# a_5626_46526# VDD.t1785 sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X7598 VDAC_N.t1356 C8_N_btm.t19 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7599 VDAC_N.t684 C9_N_btm.t40 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7600 a_13373_46526# a_12651_44576.t25 VDD.t2982 VDD.t2981 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7601 VDAC_P.t1356 C9_P_btm.t43 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7602 a_5334_30651.t1 a_13023_42718# VSS.t1883 VSS.t1882 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X7603 a_10913_42968# a_7557_43236.t15 VDD.t216 VDD.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X7604 VDAC_P.t684 C6_P_btm.t45 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7605 VDD.t2589 VSS.t3774 VDD.t2588 VDD.t2587 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X7606 VSS.t2112 a_22959_43806# a_17564_32305.t0 VSS.t1452 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7607 a_n1551_45412.t7 a_2424_46794.t11 VDD.t2950 VDD.t2949 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7608 VDAC_N.t1324 C10_N_btm.t63 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7609 VDAC_P.t1324 C10_P_btm.t70 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7610 VDAC_P.t108 C9_P_btm.t41 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7611 a_10813_46500# a_10595_46904# VDD.t2119 VDD.t2118 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X7612 VDAC_P.t1292 C10_P_btm.t69 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7613 a_6631_42883# a_5840_42718.t5 VDD.t2980 VDD.t2979 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X7614 VDAC_P.t652 C9_P_btm.t40 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7615 VDAC_P.t1260 C9_P_btm.t36 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7616 VSS.t2505 VSS.t2506 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7617 a_16981_46232# a_16921_46364# a_16885_46232# VDD.t1300 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X7618 VDD.t2257 a_n2840_46500# a_n2810_46526.t2 VDD.t1597 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X7619 VDAC_N.t108 C7_N_btm.t11 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7620 VSS.t862 a_663_47874# DATA[1].t0 VSS.t861 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7621 VDAC_P.t332 C10_P_btm.t68 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7622 VDAC_N.t1292 C10_N_btm.t62 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7623 VDAC_N.t652 C10_N_btm.t61 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7624 VDD.t1441 a_6631_44582# a_5419_47258# VDD.t1440 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7625 VDD.t265 a_n1827_44324.t9 a_22223_46534# VDD.t264 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7626 a_11834_45982# a_11788_46134# VSS.t1648 VSS.t1647 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X7627 VDAC_P.t1228 C10_P_btm.t67 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7628 a_10612_43806# a_7557_43236.t27 VSS.t234 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7629 VDAC_N.t1260 C10_N_btm.t60 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7630 VDAC_P.t620 C10_P_btm.t66 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7631 C8_P_btm.t275 a_n2810_44350.t5 VSS.t2797 VSS.t2796 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7632 VSS.t1043 a_19566_45670# a_19520_46500# VSS.t1042 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7633 a_21276_30659.t2 a_22959_47070# VDD.t1139 VDD.t1138 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7634 VDAC_N.t332 C9_N_btm.t39 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7635 VDAC_N.t1228 C10_N_btm.t59 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7636 VDAC_P.t1196 C9_P_btm.t35 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7637 VDAC_P.t172 C10_P_btm.t65 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7638 VDAC_N.t620 C8_N_btm.t18 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7639 VDAC_P.t1164 C9_P_btm.t33 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7640 VREF.t58 a_n4515_30659.t9 C10_P_btm.t1061 VDD.t2995 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7641 VDAC_P.t588 C9_P_btm.t32 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7642 a_12651_44576.t0 a_16579_43566# VSS.t1963 VSS.t1962 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7643 VDD.t2725 a_n2038_35608# SMPL_ON_P.t7 VDD.t2724 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7644 a_5748_44466# a_4993_47044# VDD.t1355 VDD.t1354 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X7645 VDAC_P.t1132 C7_P_btm.t13 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7646 VDAC_N.t1196 VSS.t3268 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7647 a_16579_43566# a_8727_47222.t11 VDD.t81 VDD.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7648 a_18314_32299.t0 a_22276_45412# VSS.t875 VSS.t874 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7649 VDD.t3 a_10259_42870.t11 a_n1551_45412.t5 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.135 ps=1.27 w=1 l=0.15
X7650 VDAC_N.t172 C10_N_btm.t58 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7651 VDAC_P.t300 C2_P_btm.t8 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7652 VDAC_N.t1164 C8_N_btm.t17 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7653 a_20159_47588# DEBUG_MUX[1].t1 VSS.t145 VSS.t144 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X7654 a_21789_35634# a_20064_35138# VSS.t882 VSS.t881 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7655 a_1019_45477# a_361_45438# a_560_45670# VDD.t763 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X7656 VSS.t2501 VSS.t2502 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7657 a_15605_45438# a_15730_45670.t23 VDD.t502 VDD.t501 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7658 VDD.t1770 a_4322_46134# a_885_44868.t9 VDD.t1769 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7659 VDAC_N.t588 C10_N_btm.t57 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7660 VDAC_P.t1100 C10_P_btm.t63 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7661 VSS.t1242 a_13635_43566# a_11455_44576.t0 VSS.t1241 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7662 a_560_45670# a_361_45438# a_702_45804# VSS.t826 sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X7663 VDAC_P.t556 C10_P_btm.t62 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7664 VSS.t1955 a_16579_43566# a_12651_44576.t2 VSS.t1954 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X7665 a_1429_47222.t2 a_15323_44894# VDD.t2086 VDD.t2085 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7666 VDAC_N.t1132 C10_N_btm.t1033 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7667 C10_N_btm.t12 a_3990_30651.t11 VCM.t11 VSS.t284 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7668 VDD.t782 a_13460_43640# a_13635_43566# VDD.t781 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X7669 a_13458_32299.t0 a_21540_43236# VSS.t1942 VSS.t1941 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7670 a_6635_47044# a_4830_43958.t8 VSS.t206 VSS.t205 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X7671 VDAC_P.t2108 C10_P_btm.t61 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7672 VDAC_N.t300 C10_N_btm.t775 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7673 VDAC_N.t1100 C10_N_btm.t516 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7674 VDD.t2484 VSS.t3780 VDD.t2483 VDD.t2482 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X7675 VDAC_P.t60 C10_P_btm.t60 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7676 VDAC_P.t2044 C10_P_btm.t59 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7677 VDD.t1405 a_713_47044# a_743_47397# VDD.t1404 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7678 VDD.t942 a_5715_45956# a_5663_45982# VDD.t941 sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X7679 VDAC_P.t1020 C10_P_btm.t58 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7680 a_3878_43806# a_135_43540.t44 VSS.t190 VSS.t189 sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X7681 VDAC_P.t1980 C10_P_btm.t57 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7682 VDAC_N.t556 C8_N_btm.t16 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7683 a_4000_42718.t2 a_3823_42718# VDD.t1643 VDD.t1642 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X7684 VDAC_P.t508 C9_P_btm.t28 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7685 VDAC_N.t2108 C9_N_btm.t38 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7686 VDAC_P.t1916 C8_P_btm.t38 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7687 a_19633_43262# a_19191_43262# VDD.t1735 VDD.t1734 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X7688 VDAC_N.t60 C10_N_btm.t493 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7689 a_14301_47070# a_13273_44868.t30 a_14219_47070# VSS.t653 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7690 a_n377_45776# a_n1067_42718.t3 VDD.t268 VDD.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7691 VDAC_P.t956 C10_P_btm.t1032 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7692 VDAC_N.t2044 C10_N_btm.t476 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7693 C10_N_btm.t24 a_22812_30659.t10 VREF.t37 VDD.t522 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7694 VDAC_N.t1020 C10_N_btm.t245 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7695 VDAC_P.t1852 C10_P_btm.t771 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7696 a_885_44868.t2 a_2587_44868.t30 VDD.t249 VDD.t248 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7697 VDAC_P.t252 C10_P_btm.t513 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7698 VDAC_N.t1980 C9_N_btm.t37 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7699 a_n4515_30659.t1 a_n2288_47588# VSS.t1238 VSS.t1237 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7700 VSS.t2186 a_22591_44894# a_17930_32299.t0 VSS.t2185 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7701 VDAC_P.t1788 C5_P_btm.t16 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7702 VDD.t1913 a_16579_43566# a_12651_44576.t7 VDD.t1912 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7703 VDAC_N.t508 C9_N_btm.t36 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7704 VDAC_N.t1916 C5_N_btm.t19 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7705 VSS.t1780 a_1239_39043# COMP_N.t1 VSS.t1770 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7706 a_8850_45412# a_9096_45276.t5 VSS.t588 VSS.t587 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.11975 ps=1.045 w=0.42 l=0.15
X7707 VDD.t69 a_n1551_45412.t10 a_22591_47070# VDD.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7708 VSS.t532 a_1203_42692.t21 a_15133_43582# VSS.t531 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7709 a_12623_43780# a_12448_43806# a_12802_43806# VSS.t1677 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X7710 a_18139_45982# a_17623_45982# a_18044_45982# VSS.t1142 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X7711 VDAC_N.t956 C10_N_btm.t237 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7712 a_16291_46758# a_16651_46500# a_16585_46642# VDD.t716 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1215 ps=1.33 w=0.42 l=0.15
X7713 VDAC_N.t1852 C9_N_btm.t35 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7714 VDAC_P.t892 C10_P_btm.t491 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7715 VSS.t2353 VSS.t2354 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7716 VDAC_N.t252 C10_N_btm.t230 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7717 VDAC_P.t1724 C9_P_btm.t29 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7718 VDD.t1261 a_49_46500# a_n61_46526# VDD.t1260 sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X7719 VDAC_P.t444 C9_P_btm.t27 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7720 VDAC_N.t1788 C9_N_btm.t34 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7721 VSS.t1854 a_18689_45412# a_17927_46195# VSS.t1853 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7722 VDAC_N.t892 C10_N_btm.t220 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7723 VDD.t703 a_4239_42883# a_1736_43276# VDD.t702 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7724 VSS.t2236 a_5655_43780# a_6717_44894# VSS.t2235 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X7725 VDAC_N.t1724 C9_N_btm.t33 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7726 VDAC_P.t1660 C9_P_btm.t26 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7727 DATA[4].t2 a_5847_47614# VSS.t1901 VSS.t1900 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X7728 VDAC_P.t828 C10_P_btm.t474 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7729 VDAC_P.t1596 C9_P_btm.t515 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7730 VDAC_P.t124 C8_P_btm.t25 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7731 VDAC_N.t444 C10_N_btm.t213 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7732 a_2801_42968# a_2755_43494.t19 a_2655_42870# VDD.t429 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X7733 VDD.t674 a_n2472_44868# a_n2442_44894.t3 VDD.t673 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X7734 VSS.t3781 C10_N_btm.t1078 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7735 VSS.t2317 VSS.t2318 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7736 VSS.t2321 VSS.t2322 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7737 VDAC_P.t1532 C10_P_btm.t243 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7738 VDAC_N.t1660 C10_N_btm.t114 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7739 VDAC_N.t828 C9_N_btm.t32 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7740 VDAC_N.t1596 C10_N_btm.t109 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7741 VSS.t290 a_3990_30651.t17 a_19555_42718# VSS.t289 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X7742 VDAC_N.t124 C10_N_btm.t106 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7743 VDAC_N.t1532 C10_N_btm.t102 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7744 VDAC_P.t764 C10_P_btm.t235 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7745 VDAC_N.t764 C10_N_btm.t99 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7746 VDAC_N.t1468 C10_N_btm.t93 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7747 VDAC_N.t380 C7_N_btm.t114 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7748 VDAC_P.t1468 C10_P_btm.t228 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7749 VDAC_P.t380 C9_P_btm.t301 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7750 VDAC_P.t1404 C8_P_btm.t22 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7751 VDAC_N.t1404 C10_N_btm.t89 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7752 a_n2293_44332# a_n1551_45412.t8 VSS.t72 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7753 VDD.t2273 VSS.t3784 VDD.t2272 VDD.t2271 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X7754 a_21847_43806# a_n2661_45420.t9 VDD.t311 VDD.t310 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7755 VDAC_N.t700 C8_N_btm.t15 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7756 a_15947_43262# a_8727_47222.t15 VDD.t43 VDD.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X7757 VDAC_P.t700 C10_P_btm.t218 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7758 a_10768_47436# a_10554_47436# VDD.t1115 VDD.t1114 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X7759 VDAC_N.t1340 C7_N_btm.t55 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7760 VDAC_P.t1340 C10_P_btm.t119 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7761 VDAC_P.t188 C6_P_btm.t25 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7762 VSS.t1079 a_11059_45956# a_10993_45982# VSS.t1078 sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X7763 a_2621_45982# a_1431_45982# a_2512_45982# VSS.t758 sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X7764 VDAC_N.t188 C9_N_btm.t31 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7765 VDAC_P.t1276 C7_P_btm.t12 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7766 VSS.t342 a_10227_47214.t23 a_10581_45982# VSS.t341 sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X7767 VDAC_N.t1276 VSS.t3270 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7768 VDAC_N.t636 C10_N_btm.t85 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7769 a_7493_43262# a_2755_43494.t16 a_7347_43494# VDD.t426 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X7770 VDAC_P.t636 C10_P_btm.t115 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7771 DATA[2].t5 a_2351_47614# VDD.t2000 VDD.t1999 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X7772 VDAC_N.t1212 C10_N_btm.t56 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7773 VDAC_P.t1212 C9_P_btm.t244 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7774 VDAC_N.t316 C7_N_btm.t23 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7775 a_n1827_45412.t0 a_13266_45412# a_13214_45758# VSS.t970 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7776 VDAC_N.t1148 C9_N_btm.t30 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7777 VSS.t3618 C10_P_btm.t21 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7778 VDAC_N.t572 C10_N_btm.t53 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7779 VDAC_N.t1084 C9_N_btm.t29 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7780 a_22276_45412# a_22455_45420# VDD.t1252 VDD.t1251 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X7781 VDAC_N.t2076 C10_N_btm.t52 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7782 VDAC_P.t316 C10_P_btm.t112 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7783 VDAC_N.t2134 C8_N_btm.t14 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7784 VDAC_N.t92 C10_N_btm.t50 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7785 a_n169_43640# a_n519_43268# a_n264_43628# VDD.t1700 sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X7786 a_11991_44172# a_11367_43806# a_11883_43806# VDD.t1612 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X7787 VDAC_P.t1148 VSS.t3343 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7788 VDAC_N.t554 C9_N_btm.t28 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7789 VSS.t3674 C6_P_btm.t3 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7790 VDAC_P.t572 C10_P_btm.t107 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7791 VDAC_P.t1084 C8_P_btm.t21 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7792 a_18394_35068.t6 SMPL.t19 VDD.t3053 VDD.t3052 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7793 VDAC_P.t2076 C10_P_btm.t104 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7794 a_2043_43958# a_n237_45454.t22 VDD.t317 VDD.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X7795 VSS.t3531 VDD.t3237 VSS.t3530 VSS.t3529 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X7796 a_7639_45804# a_n99_45438.t5 a_7276_45670# VSS.t2092 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7797 VDAC_P.t2134 C10_P_btm.t100 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7798 VSS.t1169 a_11427_43566# a_7557_43236.t1 VSS.t1168 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X7799 VDD.t410 a_13248_45956.t21 a_15389_47730# VDD.t409 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X7800 a_15879_47320# a_15691_47436# VSS.t773 VSS.t772 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1359 ps=1.1 w=0.65 l=0.15
X7801 C10_N_btm.t6 a_18314_32299.t10 VSS.t258 VSS.t257 sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7802 a_13464_45758# a_11455_44576.t15 VSS.t2715 VSS.t2714 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7803 VDAC_N.t1052 C7_N_btm.t10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7804 VDAC_N.t2012 C10_N_btm.t49 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7805 VDAC_P.t92 C10_P_btm.t97 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7806 VSS.t808 a_7309_44466# a_7415_44466# VSS.t807 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7807 VDAC_N.t28 C9_N_btm.t503 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7808 VDAC_P.t554 C7_P_btm.t120 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7809 VSS.t76 a_n1551_45412.t13 a_22591_47070# VSS.t75 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X7810 VSS.t1281 a_18803_47070# a_18822_46526# VSS.t1280 sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X7811 VDAC_P.t1052 C4_P_btm.t16 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7812 VDAC_P.t2012 C9_P_btm.t229 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7813 a_16579_43566# a_16404_43640# a_16758_43628# VSS.t1396 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X7814 VDAC_N.t2130 C9_N_btm.t248 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7815 C10_P_btm.t3 a_3990_30651.t12 VCM.t12 VSS.t285 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7816 a_3686_44172# a_2609_43806# a_3524_43806# VDD.t1159 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X7817 VDAC_P.t28 C8_P_btm.t19 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7818 VDAC_N.t1564 C10_N_btm.t45 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7819 a_9947_47044# a_10150_47322# VDD.t686 VDD.t685 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X7820 a_15321_46846# a_14757_45982# VSS.t1287 VSS.t1286 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X7821 a_16211_44582# a_16291_44914# a_16385_44688# VSS.t1727 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X7822 VDAC_N.t988 C9_N_btm.t120 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7823 VDAC_P.t2130 C10_P_btm.t92 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7824 a_5351_43806# a_4835_43806# a_5256_43806# VSS.t1002 sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X7825 VDAC_P.t1564 C10_P_btm.t87 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7826 VDAC_P.t988 C9_P_btm.t116 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7827 VSS.t1650 a_12121_45956# a_12055_45982# VSS.t1649 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X7828 VDAC_P.t26 C10_P_btm.t55 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7829 VDAC_N.t26 C9_N_btm.t113 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7830 a_9987_42968# a_2755_43494.t17 a_10069_42718# VSS.t514 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X7831 VDAC_P.t1078 C8_P_btm.t18 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7832 VDAC_P.t540 C10_P_btm.t54 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7833 VSS.t2806 a_14766_45596.t11 a_15221_47044# VSS.t2805 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.17225 ps=1.83 w=0.65 l=0.15
X7834 VSS.t2793 a_n2103_45412.t12 a_n2661_44868# VSS.t2792 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7835 VDAC_N.t1078 C10_N_btm.t44 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7836 VDAC_P.t1884 C10_P_btm.t51 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7837 VDAC_N.t540 C10_N_btm.t42 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7838 VDAC_P.t24 C10_P_btm.t50 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7839 VDD.t658 a_8850_45412# a_n1827_44868.t5 VDD.t657 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7840 VREF.t66 a_n4515_30659.t17 C10_P_btm.t1069 VDD.t3003 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7841 VDAC_P.t2126 C9_P_btm.t109 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7842 VSS.t3620 C10_N_btm.t1058 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7843 VDAC_P.t1308 C10_P_btm.t47 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7844 VDAC_N.t1884 C8_N_btm.t13 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7845 VDAC_N.t24 C9_N_btm.t56 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7846 a_2151_45670# a_n53_44363.t22 a_2385_45438# VDD.t566 sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X7847 a_93_46892# a_49_46500# a_n73_46904# VSS.t1331 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X7848 a_2645_46824# a_885_44868.t28 VSS.t2760 VSS.t2759 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X7849 VSS.t1192 a_6325_45736# a_6259_45804# VSS.t1191 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X7850 a_3754_39466# a_7754_39632# VSS.t693 sky130_fd_pr__res_high_po_0p35 l=18
X7851 a_10111_45776# a_4908_45956# VDD.t1748 VDD.t1747 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7852 EN_VIN_BSTR_P.t3 a_n1732_35090.t9 w_1375_34946.t11 w_1375_34946.t10 sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X7853 VSS.t1194 a_11017_45736# a_10951_45804# VSS.t1193 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X7854 VSS.t3141 VDD.t3149 VSS.t3140 VSS.t3139 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X7855 a_n2442_43262.t0 a_n2472_43236# VSS.t2173 VSS.t803 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X7856 a_n2661_43780# a_n1551_44324.t11 VSS.t133 VSS.t132 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7857 VDAC_N.t2126 C8_N_btm.t243 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7858 VDAC_N.t1308 C10_N_btm.t38 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7859 a_18136_44716# a_17531_44894# VDD.t1922 VDD.t1070 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X7860 VSS.t728 a_11183_42718# a_5542_30651.t0 VSS.t727 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X7861 a_4704_47044# a_5089_47044# a_4833_47320# VDD.t1603 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X7862 VDAC_N.t476 C6_N_btm.t52 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7863 VDAC_N.t22 C7_N_btm.t6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7864 VDAC_N.t290 C10_N_btm.t37 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7865 VDAC_P.t476 C7_P_btm.t70 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7866 C10_P_btm.t1062 a_n4515_30659.t10 VREF.t59 VDD.t2996 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X7867 VDAC_P.t22 C10_P_btm.t42 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7868 VDAC_P.t290 C6_P_btm.t9 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7869 VDAC_N.t4 a_3222_30651.t12 VCM.t30 VSS.t664 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7870 VDAC_P.t9 C8_P_btm.t255 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7871 VDAC_P.t12 C9_P_btm.t101 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7872 a_13536_43780# a_13715_43780# VDD.t1199 VDD.t1198 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X7873 VSS.t219 a_7557_43236.t11 a_13848_46842# VSS.t218 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X7874 VDAC_P.t14 C8_P_btm.t132 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7875 VDD.t2827 a_11455_44576.t27 a_n1827_45412.t7 VDD.t2826 sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.135 ps=1.27 w=1 l=0.15
X7876 VSS.t3129 VDD.t3145 VSS.t3128 VSS.t3127 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X7877 VDAC_N.t12 C10_N_btm.t35 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7878 a_15549_47044.t2 a_15730_45670.t11 VSS.t567 VSS.t566 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7879 a_570_44324# a_546_43100# VSS.t1811 VSS.t1810 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.11975 ps=1.045 w=0.42 l=0.15
X7880 VDAC_N.t14 C9_N_btm.t53 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7881 VDAC_P.t16 VSS.t3375 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7882 VDAC_P.t18 C10_P_btm.t40 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7883 VDAC_P.t20 C10_P_btm.t39 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7884 a_10795_43262# a_10227_47214.t28 VDD.t301 VDD.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X7885 a_1784_43378# a_1736_43276# a_1700_43378# VDD.t1133 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7886 VDAC_P.t796 C10_P_btm.t36 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7887 VDAC_N.t16 C10_N_btm.t34 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7888 VDAC_N.t18 C10_N_btm.t1034 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7889 VDAC_N.t20 C10_N_btm.t517 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7890 VDAC_P.t1820 C10_P_btm.t35 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7891 a_22609_38842# a_22469_39973# CAL_N.t1 VSS.t2592 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X7892 VSS.t3800 C10_P_btm.t30 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7893 VDD.t1814 a_17763_44868# a_17721_45144# VDD.t1813 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7894 VDAC_N.t796 C7_N_btm.t7 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7895 VDAC_N.t1820 C10_N_btm.t477 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7896 a_16111_45412# a_16287_45744# a_16239_45804# VSS.t2044 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X7897 a_5700_37509.t1 VDAC_N.t284 a_8912_37509.t7 VDD.t2244 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X7898 a_10554_47436# a_10467_47212# a_10150_47322# VDD.t2134 sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X7899 VDAC_N.t1180 C9_N_btm.t49 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7900 VSS.t3801 C0_dummy_P_btm.t2 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7901 VDAC_P.t284 C9_P_btm.t94 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7902 VDAC_P.t1180 C8_P_btm.t110 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7903 a_11415_45670# a_11687_45528# a_11645_45554# VDD.t1117 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7904 a_8912_37509.t31 VDAC_P.t668 a_5088_37509.t13 VDD.t2251 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X7905 VSS.t511 a_2755_43494.t12 a_4364_45982# VSS.t510 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7906 VDAC_P.t1436 C10_P_btm.t33 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7907 DATA[2].t2 a_2351_47614# VSS.t2050 VSS.t2049 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7908 VDD.t1608 a_n2472_46500# a_n2442_46526.t2 VDD.t1451 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X7909 VDD.t666 a_22223_43270# a_14087_32299.t2 VDD.t665 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7910 VDD.t2402 VSS.t3680 VDD.t2401 VDD.t2400 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X7911 a_10901_42718# a_1203_42692.t27 a_10913_42968# VDD.t483 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X7912 VDAC_P.t412 C10_P_btm.t32 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7913 VDAC_N.t668 C1_N_btm.t1 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7914 VDAC_N.t1436 C7_N_btm.t5 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7915 VDAC_N.t412 C10_N_btm.t238 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7916 VDAC_N.t1692 C10_N_btm.t221 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7917 VDAC_P.t1692 C9_P_btm.t52 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7918 VDAC_N.t924 C9_N_btm.t46 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7919 VDAC_N.t1948 C8_N_btm.t58 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7920 VDAC_P.t924 VSS.t3354 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7921 a_n1067_42718.t0 a_n1237_42718# VSS.t2647 VSS.t2646 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X7922 VDAC_N.t156 C9_N_btm.t24 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7923 VDAC_P.t1948 C7_P_btm.t53 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7924 VDAC_N.t1116 C9_N_btm.t23 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7925 a_n2038_35608# a_n1586_35608# VDD.t1317 VDD.t1316 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7926 VDAC_P.t156 C9_P_btm.t49 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7927 VDAC_P.t1116 C10_P_btm.t1033 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7928 VDD.t208 a_4830_43958.t17 a_9343_45982# VDD.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X7929 VSS.t1186 a_989_45736# a_923_45804# VSS.t1185 sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X7930 VDAC_P.t604 C9_P_btm.t45 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7931 VDAC_N.t604 C10_N_btm.t118 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7932 VSS.t3468 VDD.t3215 VSS.t3467 VSS.t3466 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X7933 VDAC_N.t1244 C10_N_btm.t110 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7934 VDAC_P.t1244 C9_P_btm.t42 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7935 a_9480_44350# a_9266_44350# VDD.t2741 VDD.t2740 sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X7936 a_4061_45956# a_n2497_47846.t8 VSS.t2097 VSS.t2096 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X7937 VDAC_N.t348 C10_N_btm.t103 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7938 VDAC_N.t1372 C8_N_btm.t26 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7939 VDAC_N.t732 C9_N_btm.t21 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7940 VDAC_P.t348 C9_P_btm.t37 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7941 VDD.t3036 a_1736_39587.t6 a_1736_39043.t2 VDD.t3035 sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X7942 VDAC_P.t1372 C9_P_btm.t34 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7943 VSS.t88 a_927_42692.t10 a_1935_44874# VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7944 VDAC_N.t1500 C9_N_btm.t20 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7945 VDD.t2233 a_9343_42718# a_5734_30651.t3 VDD.t2232 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7946 a_7981_45956# a_7648_46134# VSS.t1558 VSS.t1557 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X7947 VDAC_N.t220 C10_N_btm.t94 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7948 a_18136_44716# a_17531_44894# VSS.t1971 VSS.t1970 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X7949 a_85_47070# a_n193_47098# VSS.t746 VSS.t745 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X7950 VDAC_N.t1628 C10_N_btm.t86 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7951 VDAC_P.t732 C10_P_btm.t514 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7952 VSS.t3014 a_n2103_44324.t9 a_n2661_43244# VSS.t2847 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7953 VSS.t1708 a_13536_43780# a_2755_43494.t0 VSS.t1707 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7954 VDAC_P.t1500 C10_P_btm.t475 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7955 a_22400_42718# a_22223_42718# VSS.t927 VSS.t926 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X7956 VDAC_N.t860 C8_N_btm.t23 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7957 a_1203_42692.t5 a_1431_47070# VDD.t2188 VDD.t2187 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7958 VDAC_P.t220 C7_P_btm.t26 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7959 VCM.t53 a_5542_30651.t9 C6_P_btm.t73 VSS.t2899 sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X7960 VDD.t2726 a_22959_44894# a_19437_31459.t2 VDD.t1284 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X7961 VDD.t152 CAL_N.t6 VDD.t152 VDD.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X7962 VDAC_P.t1628 C10_P_btm.t236 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7963 VDAC_P.t860 C4_P_btm.t11 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7964 VDAC_P.t1756 C10_P_btm.t219 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7965 VDAC_P.t2122 C10_P_btm.t116 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7966 a_5700_37509.t10 VDAC_N.t1756 a_8912_37509.t16 VDD.t2241 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X7967 VDAC_N.t2122 C7_N_btm.t4 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7968 a_18020_46526# a_17583_46500# VDD.t819 VDD.t818 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7969 VDAC_N.t1074 C6_N_btm.t43 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7970 VDD.t2037 EN_OFFSET_CAL.t1 a_16335_47614# VDD.t2036 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X7971 a_3437_46532# a_3271_46532# VDD.t1619 VDD.t1618 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7972 VDAC_N.t2118 C10_N_btm.t532 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7973 VDAC_N.t550 C9_N_btm.t17 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7974 VDAC_P.t1074 C10_P_btm.t108 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7975 VDAC_P.t2118 C7_P_btm.t21 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7976 VDAC_N.t2114 C8_N_btm.t10 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7977 VDAC_P.t550 C10_P_btm.t101 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7978 VSS.t428 a_n690_43494.t22 a_n685_43268# VSS.t427 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7979 VDAC_P.t2114 C8_P_btm.t55 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7980 VDAC_N.t9 C9_N_btm.t16 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7981 VSS.t3475 VDD.t3218 VSS.t3474 VSS.t3473 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7982 VDAC_N.t1380 VSS.t3331 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7983 VDD.t1702 a_16576_44868# a_n2293_47044.t2 VDD.t1701 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X7984 VSS.t3078 VDD.t3128 VSS.t3077 VSS.t3076 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X7985 VSS.t544 a_1203_42692.t30 a_12833_42718# VSS.t543 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7986 a_16868_44670# a_12651_44576.t11 VSS.t2863 VSS.t2862 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7987 VDD.t3057 SMPL.t23 a_n1732_35090.t7 VDD.t3056 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7988 VDAC_N.t970 C9_N_btm.t14 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7989 VDAC_P.t388 C10_P_btm.t93 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7990 VSS.t944 a_n2840_43236# a_n2810_43262.t0 VSS.t943 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X7991 VSS.t1775 a_10596_44324# a_n2661_46508.t2 VSS.t1774 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X7992 VDAC_P.t864 C9_P_btm.t30 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7993 a_16555_46616# a_13248_45956.t13 VDD.t401 VDD.t400 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1226 ps=1.32 w=0.42 l=0.15
X7994 VDAC_N.t1187 VSS.t3267 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7995 VSS.t950 a_n447_47044# a_n749_47846# VSS.t949 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7996 VDAC_N.t693 C9_N_btm.t13 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X7997 VDD.t277 a_n1827_44868.t9 a_22223_47070# VDD.t276 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X7998 VSS.t43 a_9521_45982.t22 a_17623_45982# VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7999 VDAC_N.t1371 C8_N_btm.t133 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8000 a_n99_45438.t1 a_n377_45776# VDD.t2806 VDD.t2805 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X8001 VDAC_N.t1417 C7_N_btm.t65 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8002 VDAC_P.t450 C6_P_btm.t6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8003 a_14373_47070# a_13248_45956.t27 a_14301_47070# VSS.t493 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X8004 VDD.t200 a_4830_43958.t9 a_5939_44894# VDD.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8005 VDAC_P.t95 C7_P_btm.t18 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8006 C8_P_btm.t4 a_5142_30651.t4 VCM.t0 VSS.t120 sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8007 a_11186_47436# a_10428_47338# a_10623_47307# VDD.t2079 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X8008 VDAC_N.t93 C9_N_btm.t504 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8009 VREF.t29 a_21788_30659.t10 C9_N_btm.t11 VDD.t2057 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X8010 a_15155_47070# a_15549_47044.t4 a_15005_47222# VSS.t2888 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.13325 ps=1.06 w=0.65 l=0.15
X8011 VSS.t1914 a_7754_38470# a_6886_37412# VSS.t1913 sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X8012 VSS.t3550 C7_P_btm.t6 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8013 VDD.t2822 a_11455_44576.t19 a_13207_46526# VDD.t2821 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8014 VDAC_P.t587 C6_P_btm.t60 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8015 VDAC_P.t65 C9_P_btm.t25 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8016 VDAC_P.t1367 C9_P_btm.t516 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8017 VDAC_P.t2115 C10_P_btm.t531 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8018 VDAC_P.t2106 C9_P_btm.t262 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8019 a_4465_45412# a_4247_45816# VSS.t1965 VSS.t1964 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X8020 VDAC_N.t2106 C9_N_btm.t262 sky130_fd_pr__cap_mim_m3_1 l=1 w=1
X8021 VDD.t1018 a_4352_46904# a_4527_46830# VDD.t1017 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X8022 a_12427_46758# a_11455_44576.t11 VSS.t2711 VSS.t2710 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
R0 a_n2661_46508.n6 a_n2661_46508.n5 642.619
R1 a_n2661_46508.n1 a_n2661_46508.t9 276.464
R2 a_n2661_46508.n4 a_n2661_46508.n1 236.27
R3 a_n2661_46508.n4 a_n2661_46508.n3 217.331
R4 a_n2661_46508.n2 a_n2661_46508.t5 212.081
R5 a_n2661_46508.n3 a_n2661_46508.t7 212.081
R6 a_n2661_46508.n5 a_n2661_46508.n0 210.234
R7 a_n2661_46508.n1 a_n2661_46508.t4 196.131
R8 a_n2661_46508.n2 a_n2661_46508.t8 139.78
R9 a_n2661_46508.n3 a_n2661_46508.t6 139.78
R10 a_n2661_46508.n3 a_n2661_46508.n2 61.346
R11 a_n2661_46508.t0 a_n2661_46508.n6 26.5955
R12 a_n2661_46508.n6 a_n2661_46508.t1 26.5955
R13 a_n2661_46508.n0 a_n2661_46508.t2 24.9236
R14 a_n2661_46508.n0 a_n2661_46508.t3 24.9236
R15 a_n2661_46508.n5 a_n2661_46508.n4 13.863
R16 VSS.n1222 VSS.n977 1.0384e+06
R17 VSS.n4627 VSS.n4626 394812
R18 VSS.n4624 VSS.t101 142422
R19 VSS.n4657 VSS.n4656 117646
R20 VSS.n4629 VSS.n4628 90524.6
R21 VSS.n4798 VSS.n476 70183.6
R22 VSS.n4657 VSS.n476 55036.1
R23 VSS.n4626 VSS.t3469 52759.4
R24 VSS.n1222 VSS.t2660 46648.6
R25 VSS.n4656 VSS.n1238 39376.9
R26 VSS.n177 VSS.t1845 35131.5
R27 VSS.n1223 VSS.n976 27943.1
R28 VSS.n4661 VSS.n942 27875.5
R29 VSS.n1149 VSS.n1142 27875.5
R30 VSS.n4661 VSS.n4660 27736.4
R31 VSS.n1151 VSS.n1142 27736.4
R32 VSS.n943 VSS.n942 27701.7
R33 VSS.n1149 VSS.n1143 27701.7
R34 VSS.n4660 VSS.n943 27562.6
R35 VSS.n1151 VSS.n1143 27562.6
R36 VSS.n4626 VSS.n1238 23080.8
R37 VSS.n1223 VSS.n1222 22838.1
R38 VSS.n1106 VSS.n1105 20879.2
R39 VSS.n1072 VSS.n306 19062.6
R40 VSS.n1072 VSS.n307 19062.6
R41 VSS.n4984 VSS.n306 19062.6
R42 VSS.n4984 VSS.n307 19062.6
R43 VSS.n4799 VSS.n4798 17268.8
R44 VSS.n1235 VSS.n1234 14988.8
R45 VSS.n4631 VSS.n4624 11901.6
R46 VSS.n4590 VSS.n4589 9192.33
R47 VSS.n4590 VSS.n475 9165.36
R48 VSS.n4798 VSS.n4797 8906.03
R49 VSS.n1185 VSS.n1108 8690.32
R50 VSS.n4658 VSS.n1238 8669.31
R51 VSS.n1105 VSS.n1018 7785.2
R52 VSS.t3446 VSS.t3051 7754.79
R53 VSS.n1091 VSS.n1034 6361.94
R54 VSS.n1091 VSS.n1035 6361.94
R55 VSS.t1074 VSS.n949 6285.71
R56 VSS.t3532 VSS.t3449 6203.83
R57 VSS.n1055 VSS.n1054 6153.48
R58 VSS.t2821 VSS.t1915 6029.23
R59 VSS.n1039 VSS.n1034 5446.47
R60 VSS.n1041 VSS.n1035 5446.47
R61 VSS.t3021 VSS.t3091 5428.35
R62 VSS.n1104 VSS.n1019 5342.18
R63 VSS.n1104 VSS.n1023 5342.18
R64 VSS.n1023 VSS.n1020 5342.18
R65 VSS.n1020 VSS.n1019 5342.18
R66 VSS.n4647 VSS.n1250 4345.59
R67 VSS.n4619 VSS.n1250 4345.59
R68 VSS.n4593 VSS.n1257 4345.59
R69 VSS.n4613 VSS.n1257 4345.59
R70 VSS.n1211 VSS.n990 4345.59
R71 VSS.n995 VSS.n990 4345.59
R72 VSS.n1197 VSS.n1005 4345.59
R73 VSS.n1008 VSS.n1005 4345.59
R74 VSS.n1022 VSS.n949 4280.65
R75 VSS.t3423 VSS.n3828 4265.13
R76 VSS.n4971 VSS.n352 4154.38
R77 VSS.n4947 VSS.n352 4154.38
R78 VSS.t73 VSS.t3048 3911.11
R79 VSS.t3497 VSS.n5354 3795.76
R80 VSS.n4994 VSS.n297 3743
R81 VSS.n297 VSS.n296 3743
R82 VSS.n4987 VSS.n4986 3743
R83 VSS.n4986 VSS.n303 3743
R84 VSS.n1064 VSS.n1049 3685.06
R85 VSS.n1056 VSS.n1049 3685.06
R86 VSS.n1064 VSS.n1050 3685.06
R87 VSS.n1056 VSS.n1050 3685.06
R88 VSS.n4586 VSS.t3455 3655.3
R89 VSS.t3500 VSS.t3121 3489.66
R90 VSS.n1236 VSS.n949 3439.63
R91 VSS.t2139 VSS.t1886 3144.06
R92 VSS.n1258 VSS.n464 3128.82
R93 VSS.n1258 VSS.n1254 3128.82
R94 VSS.n1253 VSS.n463 3128.82
R95 VSS.n4618 VSS.n1253 3128.82
R96 VSS.n1208 VSS.n991 3128.82
R97 VSS.n1208 VSS.n994 3128.82
R98 VSS.n1002 VSS.n1000 3128.82
R99 VSS.n1002 VSS.n998 3128.82
R100 VSS.t3103 VSS.t427 3118.77
R101 VSS.t3399 VSS.t3210 3101.92
R102 VSS.t3076 VSS.t3399 3101.92
R103 VSS.t3449 VSS.t3479 3101.92
R104 VSS.t3106 VSS.t3532 3101.92
R105 VSS.n2313 VSS.t1861 3101.92
R106 VSS.t3526 VSS.t3544 3101.92
R107 VSS.t3494 VSS.t3103 3101.92
R108 VSS.n1183 VSS.n1016 3082.34
R109 VSS.n1187 VSS.n1016 3082.34
R110 VSS.n4633 VSS.n1239 3082.34
R111 VSS.n4654 VSS.n1239 3082.34
R112 VSS.t3184 VSS.t3458 3036
R113 VSS.n4942 VSS.n369 2914.44
R114 VSS.n4968 VSS.n353 2885.47
R115 VSS.n4949 VSS.n369 2885.47
R116 VSS.n4968 VSS.n351 2821.74
R117 VSS.t3461 VSS.t2585 2731.03
R118 VSS.n3231 VSS.t3509 2714.18
R119 VSS.t3073 VSS.n3690 2714.18
R120 VSS.t3235 VSS.n2313 2714.18
R121 VSS.n2258 VSS.t3439 2714.18
R122 VSS.t3118 VSS.t3142 2698.67
R123 VSS.t3172 VSS.t3036 2698.67
R124 VSS.t3082 VSS.t3482 2698.67
R125 VSS.n1192 VSS.n1010 2690.47
R126 VSS.n1192 VSS.n1011 2690.47
R127 VSS.n1246 VSS.n1244 2690.47
R128 VSS.n4650 VSS.n1244 2690.47
R129 VSS.n1227 VSS.n1224 2549.41
R130 VSS.n1227 VSS.n951 2549.41
R131 VSS.n1232 VSS.n952 2549.41
R132 VSS.n976 VSS.n952 2549.41
R133 VSS.t1845 VSS.t2166 2438.55
R134 VSS.t3544 VSS.t140 2410.73
R135 VSS.n5354 VSS.n5353 2402.01
R136 VSS.n5353 VSS.n5352 2402.01
R137 VSS.n5352 VSS.n5351 2402.01
R138 VSS.t3482 VSS.t1235 2398
R139 VSS.t3458 VSS.t2047 2398
R140 VSS.t3169 VSS.t863 2398
R141 VSS.t3055 VSS.t144 2372.33
R142 VSS.t3142 VSS.t142 2372.33
R143 VSS.t1739 VSS.t3055 2368.67
R144 VSS.t3036 VSS.t2960 2368.67
R145 VSS.t3479 VSS.t2964 2360.15
R146 VSS.t3210 VSS.t429 2343.29
R147 VSS.t2977 VSS.t3076 2343.29
R148 VSS.t3198 VSS.t1272 2343.29
R149 VSS.t3248 VSS.t3021 2326.44
R150 VSS.t3091 VSS.t3235 2326.44
R151 VSS.t3064 VSS.t3136 2326.44
R152 VSS.t3506 VSS.t3538 2326.44
R153 VSS.n4587 VSS.n4586 2294.92
R154 VSS.n4588 VSS.n4587 2294.92
R155 VSS.n4589 VSS.n4588 2294.92
R156 VSS.n5351 VSS.n5350 2258.84
R157 VSS.n1234 VSS.n177 2210.13
R158 VSS.n4585 VSS.t3169 2192.67
R159 VSS.n4676 VSS.n4675 2187.94
R160 VSS.n911 VSS.n909 2187.94
R161 VSS.t156 VSS.t1087 2174.71
R162 VSS.n4677 VSS.n616 2166.4
R163 VSS.n908 VSS.n770 2166.4
R164 VSS.n4796 VSS.n545 2160.03
R165 VSS.t1574 VSS.t1678 2149.43
R166 VSS.n1090 VSS.n1040 2126.44
R167 VSS.n1090 VSS.n1043 2126.44
R168 VSS.t1282 VSS.t3223 2098.85
R169 VSS.t1770 VSS.t516 2065.13
R170 VSS.n4591 VSS.n475 2048.11
R171 VSS.t1068 VSS.t1652 2031.42
R172 VSS.n4797 VSS.n478 2013.99
R173 VSS.n1105 VSS.t2821 2011.15
R174 VSS.t2077 VSS.t710 1980.84
R175 VSS.n4990 VSS.n298 1970
R176 VSS.n4990 VSS.n302 1970
R177 VSS.t3244 VSS.n1247 1966.78
R178 VSS.t1201 VSS.t3042 1963.98
R179 VSS.t3085 VSS.t2128 1963.98
R180 VSS.t1355 VSS.t3058 1963.98
R181 VSS.t3201 VSS.t1656 1963.98
R182 VSS.t1122 VSS.t3145 1963.98
R183 VSS.t935 VSS.t3033 1963.98
R184 VSS.t1452 VSS.t3112 1963.98
R185 VSS.t3178 VSS.t945 1963.98
R186 VSS.t301 VSS.t3500 1955.56
R187 VSS.t417 VSS.t3187 1955.56
R188 VSS.t3070 VSS.t2759 1955.56
R189 VSS.n3690 VSS.t411 1955.56
R190 VSS.t2731 VSS.t3214 1955.56
R191 VSS.t3207 VSS.t1888 1955.56
R192 VSS.n3231 VSS.t3106 1938.7
R193 VSS.t3181 VSS.n3230 1938.7
R194 VSS.t3061 VSS.t3506 1938.7
R195 VSS.t2693 VSS.t1537 1930.27
R196 VSS.t1791 VSS.t2578 1921.84
R197 VSS.t1062 VSS.t1050 1904.98
R198 VSS.t1747 VSS.t1784 1888.12
R199 VSS.n4958 VSS.n363 1877.29
R200 VSS.n1112 VSS.n1111 1857.31
R201 VSS.n1111 VSS.n1015 1857.31
R202 VSS.n4623 VSS.n4622 1857.31
R203 VSS.n4622 VSS.n1240 1857.31
R204 VSS.n140 VSS.t3541 1855.33
R205 VSS.t1284 VSS.t2609 1854.41
R206 VSS.n4628 VSS.t3054 1803.53
R207 VSS.n4958 VSS.n364 1784.59
R208 VSS.n4994 VSS.n298 1773
R209 VSS.n4987 VSS.n298 1773
R210 VSS.n302 VSS.n296 1773
R211 VSS.n303 VSS.n302 1773
R212 VSS.t1576 VSS.t878 1753.26
R213 VSS.t3160 VSS.t1904 1723.33
R214 VSS.t2040 VSS.t689 1719.54
R215 VSS.t955 VSS.t3094 1697.67
R216 VSS.t3541 VSS.t1489 1694
R217 VSS.n1237 VSS.n1236 1645.72
R218 VSS.t480 VSS.t488 1643.68
R219 VSS.t1572 VSS.t2150 1635.25
R220 VSS.t566 VSS.t1140 1618.39
R221 VSS.t2792 VSS.t360 1618.39
R222 VSS.t109 VSS.t2557 1618.39
R223 VSS.t132 VSS.t303 1618.39
R224 VSS.t299 VSS.t2847 1618.39
R225 VSS.t678 VSS.t593 1618.39
R226 VSS.t1915 VSS.n1019 1615.98
R227 VSS.t973 VSS.t2069 1609.96
R228 VSS.t2962 VSS.t874 1609.96
R229 VSS.t739 VSS.t2194 1609.96
R230 VSS.t1941 VSS.t1092 1609.96
R231 VSS.n1235 VSS.n950 1607.72
R232 VSS.t1827 VSS.t1341 1601.53
R233 VSS.t2784 VSS.t2788 1601.53
R234 VSS.t2901 VSS.t1491 1601.53
R235 VSS.t1428 VSS.t1392 1601.53
R236 VSS.t3426 VSS.t2259 1601.53
R237 VSS.t828 VSS.t676 1601.53
R238 VSS.t1743 VSS.t128 1593.1
R239 VSS.t1336 VSS.t1411 1593.1
R240 VSS.t105 VSS.t733 1593.1
R241 VSS.t2559 VSS.t1669 1593.1
R242 VSS.t1083 VSS.t674 1593.1
R243 VSS.t1268 VSS.t1262 1593.1
R244 VSS.t353 VSS.t1450 1593.1
R245 VSS.t2185 VSS.t597 1593.1
R246 VSS.t741 VSS.t905 1593.1
R247 VSS.t1993 VSS.t991 1593.1
R248 VSS.t1205 VSS.t830 1593.1
R249 VSS.t687 VSS.t803 1593.1
R250 VSS.t651 VSS.t1436 1584.67
R251 VSS.t612 VSS.t604 1584.67
R252 VSS.t609 VSS.t600 1584.67
R253 VSS.t600 VSS.t1825 1584.67
R254 VSS.t0 VSS.t2849 1584.67
R255 VSS.t220 VSS.t1315 1584.67
R256 VSS.t979 VSS.t1460 1584.67
R257 VSS.t2555 VSS.t3248 1584.67
R258 VSS.t2716 VSS.t508 1584.67
R259 VSS.t2807 VSS.t1466 1584.67
R260 VSS.t3538 VSS.t130 1584.67
R261 VSS.t1245 VSS.t842 1584.67
R262 VSS.t967 VSS.t1598 1584.67
R263 VSS.t1718 VSS.t1228 1584.67
R264 VSS.t1881 VSS.t2868 1576.25
R265 VSS.t218 VSS.t1525 1567.82
R266 VSS.t3232 VSS.t1020 1567.82
R267 VSS.t10 VSS.t3523 1567.82
R268 VSS.t1288 VSS.t3064 1567.82
R269 VSS.n1078 VSS.n1048 1564.22
R270 VSS.n1080 VSS.n1048 1564.22
R271 VSS.n1080 VSS.n1047 1564.22
R272 VSS.n1078 VSS.n1047 1564.22
R273 VSS.t50 VSS.t1401 1559.39
R274 VSS.t922 VSS.t40 1550.96
R275 VSS.t34 VSS.t2017 1550.96
R276 VSS.t2063 VSS.t998 1550.96
R277 VSS.t2862 VSS.t2053 1550.96
R278 VSS.n2836 VSS.t3061 1550.96
R279 VSS.t599 VSS.t3485 1542.53
R280 VSS.n59 VSS.t3160 1518
R281 VSS.n1228 VSS.n953 1494.88
R282 VSS.n1228 VSS.n957 1494.88
R283 VSS.n5354 VSS.t3042 1483.52
R284 VSS.n4586 VSS.t3085 1483.52
R285 VSS.n5353 VSS.t3058 1483.52
R286 VSS.n4587 VSS.t3201 1483.52
R287 VSS.n5352 VSS.t3145 1483.52
R288 VSS.n4588 VSS.t3033 1483.52
R289 VSS.n5351 VSS.t3112 1483.52
R290 VSS.t3488 VSS.t824 1483.52
R291 VSS.n4589 VSS.t3178 1483.52
R292 VSS.n5350 VSS.t3517 1460.74
R293 VSS.n4799 VSS.n475 1460.58
R294 VSS.t2916 VSS.t3124 1458.24
R295 VSS.t1737 VSS.t2751 1416.09
R296 VSS.t2759 VSS.t1189 1416.09
R297 VSS.t1645 VSS.t1649 1416.09
R298 VSS.t888 VSS.t1068 1416.09
R299 VSS.t2156 VSS.t1871 1399.23
R300 VSS.t849 VSS.t1551 1399.23
R301 VSS.t1488 VSS.t917 1399.23
R302 VSS.t685 VSS.t1999 1393.33
R303 VSS.n4940 VSS.n366 1390.59
R304 VSS.n4940 VSS.n4939 1390.59
R305 VSS.n4971 VSS.n351 1390.59
R306 VSS.n4947 VSS.n4942 1390.59
R307 VSS.n4955 VSS.n356 1390.59
R308 VSS.n4955 VSS.n359 1390.59
R309 VSS.n360 VSS.n357 1390.59
R310 VSS.n361 VSS.n360 1390.59
R311 VSS.t3094 VSS.t1415 1386
R312 VSS.t2680 VSS.t1877 1373.95
R313 VSS.t2005 VSS.t3133 1364
R314 VSS.t1174 VSS.t3529 1356.67
R315 VSS.t2061 VSS.t3466 1356.67
R316 VSS.t3115 VSS.t2818 1356.67
R317 VSS.t1183 VSS.t531 1340.23
R318 VSS.t3514 VSS.t2023 1323.37
R319 VSS.t1590 VSS.t1660 1306.51
R320 VSS.t2739 VSS.n1257 1301.15
R321 VSS.t2998 VSS.t492 1289.66
R322 VSS.t3226 VSS.t649 1284.62
R323 VSS.t504 VSS.t1714 1281.23
R324 VSS.t2605 VSS.t1539 1281.19
R325 VSS.t2745 VSS.t2088 1264.37
R326 VSS.t2678 VSS.t2588 1264.37
R327 VSS.n3828 VSS.t1090 1255.94
R328 VSS.t329 VSS.t920 1255.94
R329 VSS.t2019 VSS.t335 1255.94
R330 VSS.t2775 VSS.t1458 1255.94
R331 VSS.t333 VSS.t1867 1255.94
R332 VSS.t77 VSS.t1637 1255.94
R333 VSS.t2239 VSS.t961 1255.94
R334 VSS.t2233 VSS.t1716 1255.94
R335 VSS.n1361 VSS.t2175 1255.94
R336 VSS.t173 VSS.t1621 1255.94
R337 VSS.t778 VSS.t2907 1247.51
R338 VSS.n1071 VSS.n1070 1239.46
R339 VSS.t815 VSS.n3059 1239.08
R340 VSS.t1549 VSS.t1313 1239.08
R341 VSS.t2609 VSS.t3417 1230.65
R342 VSS.n1510 VSS.t62 1230.65
R343 VSS.n1183 VSS.n1112 1225.03
R344 VSS.n1187 VSS.n1015 1225.03
R345 VSS.n4633 VSS.n4623 1225.03
R346 VSS.n4654 VSS.n1240 1225.03
R347 VSS.n4647 VSS.n463 1216.76
R348 VSS.n4812 VSS.n463 1216.76
R349 VSS.n4812 VSS.n464 1216.76
R350 VSS.n4593 VSS.n464 1216.76
R351 VSS.n4619 VSS.n4618 1216.76
R352 VSS.n4618 VSS.n4617 1216.76
R353 VSS.n4617 VSS.n1254 1216.76
R354 VSS.n4613 VSS.n1254 1216.76
R355 VSS.n1211 VSS.n991 1216.76
R356 VSS.n1201 VSS.n991 1216.76
R357 VSS.n1201 VSS.n1000 1216.76
R358 VSS.n1197 VSS.n1000 1216.76
R359 VSS.n995 VSS.n994 1216.76
R360 VSS.n1204 VSS.n994 1216.76
R361 VSS.n1204 VSS.n998 1216.76
R362 VSS.n1008 VSS.n998 1216.76
R363 VSS.n1040 VSS.n1039 1210.97
R364 VSS.n1043 VSS.n1041 1210.97
R365 VSS.n4585 VSS.n4584 1198.25
R366 VSS.n5745 VSS.n19 1198.25
R367 VSS.n5699 VSS.n37 1198.25
R368 VSS.n5654 VSS.n59 1198.25
R369 VSS.n5609 VSS.n79 1198.25
R370 VSS.n138 VSS.n99 1198.25
R371 VSS.n139 VSS.n116 1198.25
R372 VSS.n5469 VSS.n140 1198.25
R373 VSS.n5424 VSS.n158 1198.25
R374 VSS.n5356 VSS.n5355 1198.25
R375 VSS.n4057 VSS.n4056 1198.25
R376 VSS.n4240 VSS.n4239 1198.25
R377 VSS.n4242 VSS.n4241 1198.25
R378 VSS.n3870 VSS.n3869 1198.25
R379 VSS.n3690 VSS.n3689 1198.25
R380 VSS.n3628 VSS.n2954 1198.25
R381 VSS.n3345 VSS.n3081 1198.25
R382 VSS.n3229 VSS.n3228 1198.25
R383 VSS.n2257 VSS.n2211 1198.25
R384 VSS.n2258 VSS.n2233 1198.25
R385 VSS.n2312 VSS.n2287 1198.25
R386 VSS.n2736 VSS.n2735 1198.25
R387 VSS.n2738 VSS.n2737 1198.25
R388 VSS.n2835 VSS.n2834 1198.25
R389 VSS.n2356 VSS.n2355 1198.25
R390 VSS.n2000 VSS.n1361 1198.25
R391 VSS.n1742 VSS.n1488 1198.25
R392 VSS.n1576 VSS.n1575 1198.25
R393 VSS.n4936 VSS.n4935 1198.25
R394 VSS.n4997 VSS.n4996 1198.25
R395 VSS.n5038 VSS.n274 1198.25
R396 VSS.n1066 VSS.n254 1198.25
R397 VSS.n5178 VSS.n5177 1198.25
R398 VSS.n5180 VSS.n5179 1198.25
R399 VSS.n1017 VSS.n212 1198.25
R400 VSS.n5274 VSS.n196 1198.25
R401 VSS.n5348 VSS.n5347 1198.25
R402 VSS.n4815 VSS.n4814 1198.25
R403 VSS.n4492 VSS.n4491 1197.79
R404 VSS.n2068 VSS.n2067 1197.79
R405 VSS.n4624 VSS.t1766 1196.93
R406 VSS.n3918 VSS.n3828 1196.86
R407 VSS.n2902 VSS.n2836 1196.86
R408 VSS.n1843 VSS.n1436 1196.63
R409 VSS.n3232 VSS.n3231 1196.22
R410 VSS.n4353 VSS.n3715 1194.5
R411 VSS.n4295 VSS.n3737 1194.5
R412 VSS.n4112 VSS.n3780 1194.5
R413 VSS.n4055 VSS.n4054 1194.5
R414 VSS.n3565 VSS.n2981 1194.5
R415 VSS.n3512 VSS.n3005 1194.5
R416 VSS.n3453 VSS.n3033 1194.5
R417 VSS.n3400 VSS.n3059 1194.5
R418 VSS.n3230 VSS.n3107 1194.5
R419 VSS.n2503 VSS.n2259 1194.5
R420 VSS.n2406 VSS.n2313 1194.5
R421 VSS.n1945 VSS.n1385 1194.5
R422 VSS.n1887 VSS.n1411 1194.5
R423 VSS.n1792 VSS.n1462 1194.5
R424 VSS.n1685 VSS.n1510 1194.5
R425 VSS.n1625 VSS.t1967 1194.5
R426 VSS.n3869 VSS.t1138 1188.51
R427 VSS.n3780 VSS.t85 1188.51
R428 VSS.n2355 VSS.t1520 1188.51
R429 VSS.n1575 VSS.t735 1188.51
R430 VSS.t58 VSS.t1967 1188.51
R431 VSS.t2799 VSS.n139 1188
R432 VSS.n5350 VSS.n177 1186.35
R433 VSS.n158 VSS.t3118 1180.67
R434 VSS.t3529 VSS.n140 1180.67
R435 VSS.n138 VSS.t3115 1180.67
R436 VSS.n79 VSS.t3082 1180.67
R437 VSS.n37 VSS.t3184 1180.67
R438 VSS.t3133 VSS.n19 1180.67
R439 VSS.n4055 VSS.t878 1180.08
R440 VSS.t387 VSS.t1798 1180.08
R441 VSS.t1321 VSS.n3229 1180.08
R442 VSS.t1006 VSS.n3081 1180.08
R443 VSS.n3033 VSS.t1526 1180.08
R444 VSS.t1710 VSS.n3005 1180.08
R445 VSS.t1969 VSS.n2312 1180.08
R446 VSS.n2312 VSS.t2035 1180.08
R447 VSS.n2737 VSS.t167 1180.08
R448 VSS.t203 VSS.n1411 1180.08
R449 VSS.t2945 VSS.n4799 1167.23
R450 VSS.t3024 VSS.n4055 1163.22
R451 VSS.t3100 VSS.n3780 1163.22
R452 VSS.t1127 VSS.t1470 1163.22
R453 VSS.t1341 VSS.t2761 1163.22
R454 VSS.t1684 VSS.t1022 1163.22
R455 VSS.n4056 VSS.t1893 1146.36
R456 VSS.n2835 VSS.t87 1146.36
R457 VSS.t1594 VSS.t3151 1137.93
R458 VSS.t1064 VSS.n196 1112.88
R459 VSS.t1329 VSS.t2777 1112.64
R460 VSS.t691 VSS.t187 1112.64
R461 VSS.t977 VSS.t626 1112.64
R462 VSS.t1939 VSS.t52 1112.64
R463 VSS.t1430 VSS.t3009 1112.64
R464 VSS.t30 VSS.t579 1112.64
R465 VSS.t912 VSS.t2243 1112.64
R466 VSS.t520 VSS.t2875 1085.4
R467 VSS.t2154 VSS.t1176 1078.93
R468 VSS.t1951 VSS.t1627 1078.93
R469 VSS.t3473 VSS.t644 1078.93
R470 VSS.t2177 VSS.t2223 1062.07
R471 VSS.t762 VSS.t1078 1062.07
R472 VSS.t2593 VSS.t1160 1062.07
R473 VSS.n1224 VSS.n957 1054.53
R474 VSS.n1232 VSS.n953 1054.53
R475 VSS.n953 VSS.n951 1054.53
R476 VSS.n976 VSS.n957 1054.53
R477 VSS.t1686 VSS.t2854 1053.64
R478 VSS.t624 VSS.t2612 1053.64
R479 VSS.t2765 VSS.t97 1053.64
R480 VSS.t1379 VSS.t315 1053.64
R481 VSS.t1615 VSS.t1613 1037.67
R482 VSS.n1234 VSS.n1233 1037.11
R483 VSS.t2581 VSS.t850 1036.78
R484 VSS.t1516 VSS.t2827 1036.78
R485 VSS.t1081 VSS.t2725 1026.67
R486 VSS.t2086 VSS.t1334 1026.67
R487 VSS.t2083 VSS.t3172 1019.33
R488 VSS.t1842 VSS.t1947 1011.49
R489 VSS.t1964 VSS.n2981 1011.49
R490 VSS.t1782 VSS.t1369 1011.49
R491 VSS.t212 VSS.t2216 1011.49
R492 VSS.n4490 VSS.n4423 1010.52
R493 VSS.t3045 VSS.t2590 994.636
R494 VSS.t3109 VSS.t2684 994.636
R495 VSS.t164 VSS.t979 986.207
R496 VSS.n3878 VSS.n3841 983.718
R497 VSS.t3420 VSS.t2853 982.668
R498 VSS.n364 VSS.n351 979.207
R499 VSS.t1962 VSS.t3166 977.779
R500 VSS.t3163 VSS.t2870 968.619
R501 VSS.n4939 VSS.n363 961.823
R502 VSS.n364 VSS.n361 961.823
R503 VSS.t903 VSS.t3547 958.314
R504 VSS.t2993 VSS.t3226 954.88
R505 VSS.t123 VSS.t3163 954.88
R506 VSS.t2771 VSS.n3737 952.49
R507 VSS.t1765 VSS.t1497 952.49
R508 VSS.t749 VSS.t2043 952.49
R509 VSS.t183 VSS.n1385 952.49
R510 VSS.t149 VSS.t1298 944.062
R511 VSS.t2065 VSS.t1818 935.633
R512 VSS.n3005 VSS.t1995 935.633
R513 VSS.t1987 VSS.t2702 935.633
R514 VSS.t1535 VSS.t1332 927.203
R515 VSS.t2607 VSS.t2583 918.774
R516 VSS.t1279 VSS.t1277 918.774
R517 VSS.t2769 VSS.t981 918.774
R518 VSS.t1040 VSS.t680 918.774
R519 VSS.t1647 VSS.t1835 918.774
R520 VSS.t702 VSS.t2682 918.774
R521 VSS.t1111 VSS.t2643 918.774
R522 VSS.t1150 VSS.t2729 918.774
R523 VSS.t2114 VSS.t1689 918.774
R524 VSS.t1888 VSS.t1066 918.774
R525 VSS.t2182 VSS.t1990 918.774
R526 VSS.t721 VSS.t957 918.774
R527 VSS.t1008 VSS.t1597 918.774
R528 VSS.t2101 VSS.t1224 918.774
R529 VSS.n4949 VSS.n366 915.471
R530 VSS.n4953 VSS.n366 915.471
R531 VSS.n4953 VSS.n356 915.471
R532 VSS.n4963 VSS.n356 915.471
R533 VSS.n4963 VSS.n357 915.471
R534 VSS.n357 VSS.n353 915.471
R535 VSS.n4939 VSS.n365 915.471
R536 VSS.n365 VSS.n359 915.471
R537 VSS.n4962 VSS.n359 915.471
R538 VSS.n4962 VSS.n361 915.471
R539 VSS.n1039 VSS.n1038 915.471
R540 VSS.n1041 VSS.n1038 915.471
R541 VSS.t745 VSS.t502 910.346
R542 VSS.t1975 VSS.t468 910.346
R543 VSS.t2702 VSS.t500 910.346
R544 VSS.t505 VSS.t1197 910.346
R545 VSS.t1967 VSS.t339 910.346
R546 VSS.t470 VSS.t2616 910.346
R547 VSS.n1075 VSS.n1074 903.087
R548 VSS.t2144 VSS.t1319 901.917
R549 VSS.t2575 VSS.t2179 901.917
R550 VSS.n1148 VSS.n1147 894.395
R551 VSS.n946 VSS.n944 894.212
R552 VSS.t654 VSS.t1664 893.487
R553 VSS.t489 VSS.t1792 893.487
R554 VSS.t2245 VSS.t2755 893.487
R555 VSS.t1705 VSS.t871 893.487
R556 VSS.n4942 VSS.n363 886.5
R557 VSS.t704 VSS.t2615 885.058
R558 VSS.t915 VSS.t210 885.058
R559 VSS.t3455 VSS.t1384 880
R560 VSS.t1837 VSS.t1853 876.629
R561 VSS.t2075 VSS.t316 876.629
R562 VSS.t2955 VSS.t2707 876.629
R563 VSS.n1462 VSS.t349 876.629
R564 VSS.n1152 VSS.n1141 871.289
R565 VSS.n948 VSS.n947 871.111
R566 VSS.n1070 VSS.n310 870.4
R567 VSS.t3523 VSS.t766 868.199
R568 VSS.t3491 VSS.t1227 868.199
R569 VSS.n1146 VSS.n1144 867.322
R570 VSS.n4663 VSS.n940 867.322
R571 VSS.n4649 VSS.n1248 862.899
R572 VSS.t620 VSS.n4240 859.77
R573 VSS.t1818 VSS.t1590 859.77
R574 VSS.t947 VSS.t1641 859.77
R575 VSS.n4622 VSS.n1245 856.985
R576 VSS.t1760 VSS.t3497 854.333
R577 VSS.t1972 VSS.t3004 854.333
R578 VSS.t1394 VSS.t3079 854.333
R579 VSS.t843 VSS.t486 851.341
R580 VSS.t233 VSS.t1989 851.341
R581 VSS.t816 VSS.t940 851.341
R582 VSS.t1444 VSS.t3420 850.668
R583 VSS.n1153 VSS.n1140 850.336
R584 VSS.n4662 VSS.n941 850.336
R585 VSS.t3466 VSS.n138 843.333
R586 VSS.t2717 VSS.t1869 842.913
R587 VSS.t1345 VSS.t1300 842.913
R588 VSS.t1359 VSS.t700 842.913
R589 VSS.t644 VSS.t56 842.913
R590 VSS.t273 VSS.t2716 842.913
R591 VSS.n2257 VSS.t2645 842.913
R592 VSS.t1564 VSS.t1608 842.913
R593 VSS.t222 VSS.t241 842.913
R594 VSS.t95 VSS.t2099 842.913
R595 VSS.t696 VSS.t1841 834.484
R596 VSS.t1298 VSS.t1279 834.484
R597 VSS.t1510 VSS.t205 834.484
R598 VSS.t1872 VSS.t2142 834.484
R599 VSS.t1498 VSS.t1493 834.484
R600 VSS.t2116 VSS.t1053 834.484
R601 VSS.t1879 VSS.t1684 834.484
R602 VSS.t1643 VSS.t1111 834.484
R603 VSS.t928 VSS.t1609 834.484
R604 VSS.t918 VSS.t1486 834.484
R605 VSS.t871 VSS.t1566 834.484
R606 VSS.t1530 VSS.t794 834.484
R607 VSS.t1990 VSS.t2148 834.484
R608 VSS.t1597 VSS.t1012 834.484
R609 VSS.t1227 VSS.t912 834.484
R610 VSS.t940 VSS.t941 834.484
R611 VSS.n1112 VSS.n1010 833.155
R612 VSS.n1015 VSS.n1011 833.155
R613 VSS.n4623 VSS.n1246 833.155
R614 VSS.n4650 VSS.n1240 833.155
R615 VSS.t2613 VSS.t2102 826.054
R616 VSS.t591 VSS.t3024 826.054
R617 VSS.t800 VSS.t1730 826.054
R618 VSS.t1789 VSS.t1812 826.054
R619 VSS.t1317 VSS.t1426 826.054
R620 VSS.t36 VSS.t1062 826.054
R621 VSS.t993 VSS.t2162 826.054
R622 VSS.t1763 VSS.t522 826.054
R623 VSS.t564 VSS.t2130 826.054
R624 VSS.t2850 VSS.t1906 826.054
R625 VSS.t583 VSS.t1774 826.054
R626 VSS.t1588 VSS.t1533 826.054
R627 VSS.t1605 VSS.t3514 826.054
R628 VSS.t1462 VSS.t1154 826.054
R629 VSS.t751 VSS.t2858 826.054
R630 VSS.t357 VSS.t1032 826.054
R631 VSS.t604 VSS.t1524 817.625
R632 VSS.t2710 VSS.t1409 817.625
R633 VSS.t477 VSS.t1545 817.625
R634 VSS.t1754 VSS.t2883 817.625
R635 VSS.t1776 VSS.t229 817.625
R636 VSS.t2620 VSS.t2914 817.625
R637 VSS.t3018 VSS.t1424 817.625
R638 VSS.t2070 VSS.t717 817.625
R639 VSS.t1152 VSS.t2731 817.625
R640 VSS.t1222 VSS.t2905 817.625
R641 VSS.t2057 VSS.t407 817.625
R642 VSS.t1839 VSS.t876 809.196
R643 VSS.t2583 VSS.t1974 809.196
R644 VSS.t1274 VSS.t1278 809.196
R645 VSS.t1796 VSS.t1681 809.196
R646 VSS.t1189 VSS.t1686 809.196
R647 VSS.t151 VSS.t2767 809.196
R648 VSS.t1144 VSS.t1127 809.196
R649 VSS.t1474 VSS.t623 809.196
R650 VSS.t706 VSS.t1143 809.196
R651 VSS.t1497 VSS.t1142 809.196
R652 VSS.t1272 VSS.t383 809.196
R653 VSS.t454 VSS.t1503 809.196
R654 VSS.t2801 VSS.t1284 809.196
R655 VSS.t1160 VSS.t616 809.196
R656 VSS.t1709 VSS.t747 809.196
R657 VSS.t698 VSS.t1464 809.196
R658 VSS.t1458 VSS.t758 809.196
R659 VSS.t1185 VSS.t615 809.196
R660 VSS.t3470 VSS.t71 809.196
R661 VSS.t362 VSS.t3470 809.196
R662 VSS.t1867 VSS.t702 809.196
R663 VSS.t2683 VSS.t703 809.196
R664 VSS.t1855 VSS.t1371 809.196
R665 VSS.t2192 VSS.t682 809.196
R666 VSS.t835 VSS.t1106 809.196
R667 VSS.t1106 VSS.t156 809.196
R668 VSS.t1832 VSS.t1547 809.196
R669 VSS.t229 VSS.t8 809.196
R670 VSS.t2640 VSS.t1110 809.196
R671 VSS.t1607 VSS.t1610 809.196
R672 VSS.t271 VSS.t2070 809.196
R673 VSS.t582 VSS.t2743 809.196
R674 VSS.t619 VSS.t888 809.196
R675 VSS.t1066 VSS.t827 809.196
R676 VSS.t1094 VSS.t3526 809.196
R677 VSS.t1960 VSS.t1439 809.196
R678 VSS.t1701 VSS.t1438 809.196
R679 VSS.t836 VSS.t1379 809.196
R680 VSS.t870 VSS.t1159 809.196
R681 VSS.t1313 VSS.t1676 809.196
R682 VSS.t1716 VSS.t1005 809.196
R683 VSS.t1226 VSS.t1002 809.196
R684 VSS.t2210 VSS.t2110 809.196
R685 VSS.t1621 VSS.t909 809.196
R686 VSS.t818 VSS.t2261 809.196
R687 VSS.t1753 VSS.t2262 809.196
R688 VSS.t128 VSS.t1203 800.766
R689 VSS.t75 VSS.t1741 800.766
R690 VSS.t1136 VSS.t301 800.766
R691 VSS.t1280 VSS.t1840 800.766
R692 VSS.t85 VSS.t2190 800.766
R693 VSS.t1351 VSS.t1274 800.766
R694 VSS.t205 VSS.t2146 800.766
R695 VSS.t1680 VSS.t1574 800.766
R696 VSS.t1640 VSS.t1303 800.766
R697 VSS.t731 VSS.t2977 800.766
R698 VSS.t1667 VSS.t105 800.766
R699 VSS.t2126 VSS.t2559 800.766
R700 VSS.t674 VSS.t1353 800.766
R701 VSS.t2152 VSS.t1257 800.766
R702 VSS.t1037 VSS.t1987 800.766
R703 VSS.t1448 VSS.t2784 800.766
R704 VSS.t1654 VSS.t353 800.766
R705 VSS.t597 VSS.t1124 800.766
R706 VSS.t2023 VSS.t1607 800.766
R707 VSS.t1491 VSS.t743 800.766
R708 VSS.t905 VSS.t937 800.766
R709 VSS.t991 VSS.t1454 800.766
R710 VSS.t1347 VSS.t2013 800.766
R711 VSS.t1032 VSS.t1943 800.766
R712 VSS.t1938 VSS.t1282 800.766
R713 VSS.t1673 VSS.t1000 800.766
R714 VSS.t1011 VSS.t1979 800.766
R715 VSS.t1002 VSS.t2059 800.766
R716 VSS.t2098 VSS.t1413 800.766
R717 VSS.t2262 VSS.t1890 800.766
R718 VSS.t805 VSS.t1205 800.766
R719 VSS.t943 VSS.t687 800.766
R720 VSS.t2257 VSS.t3220 800.312
R721 VSS.t3220 VSS.t669 796.878
R722 VSS.t3408 VSS.t1292 796.878
R723 VSS.t1750 VSS.t2561 796.878
R724 VSS.n1017 VSS.t2033 796.878
R725 VSS.t1401 VSS.t3461 792.337
R726 VSS.t2095 VSS.t617 792.337
R727 VSS.t2135 VSS.t2177 792.337
R728 VSS.t2929 VSS.t464 792.337
R729 VSS.t3509 VSS.t1040 792.337
R730 VSS.t28 VSS.t3190 792.337
R731 VSS.t1933 VSS.t2975 792.337
R732 VSS.t318 VSS.t1763 792.337
R733 VSS.t2823 VSS.t835 792.337
R734 VSS.t1397 VSS.t2786 792.337
R735 VSS.t432 VSS.t751 792.337
R736 VSS.t2616 VSS.t723 792.337
R737 VSS.t2925 VSS.t828 792.337
R738 VSS.t3148 VSS.t2133 791.59
R739 VSS.t3547 VSS.n1017 790.009
R740 VSS.t529 VSS.t58 783.909
R741 VSS.n1248 VSS.n1247 777.385
R742 VSS.t3121 VSS.t3446 775.48
R743 VSS.t3051 VSS.t3423 775.48
R744 VSS.t2598 VSS.t1089 775.48
R745 VSS.t3048 VSS.t3073 775.48
R746 VSS.t779 VSS.t2192 775.48
R747 VSS.t682 VSS.t1270 775.48
R748 VSS.t1087 VSS.t2634 775.48
R749 VSS.t225 VSS.t638 775.48
R750 VSS.t15 VSS.t2958 775.48
R751 VSS.t1547 VSS.t60 775.48
R752 VSS.t2721 VSS.t6 775.48
R753 VSS.t3439 VSS.t3232 775.48
R754 VSS.t1020 VSS.t273 775.48
R755 VSS.t8 VSS.t26 775.48
R756 VSS.t2914 VSS.t1288 775.48
R757 VSS.n2836 VSS.t3207 775.48
R758 VSS.t241 VSS.t1981 775.48
R759 VSS.n1411 VSS.t3193 775.48
R760 VSS.t1100 VSS.t237 775.48
R761 VSS.t854 VSS.n1361 775.48
R762 VSS.t636 VSS.t1576 767.051
R763 VSS.t911 VSS.t2741 767.051
R764 VSS.t2025 VSS.t706 767.051
R765 VSS.t850 VSS.t331 767.051
R766 VSS.t1340 VSS.t2814 767.051
R767 VSS.t2590 VSS.t2775 767.051
R768 VSS.t2187 VSS.t179 767.051
R769 VSS.t2684 VSS.t333 767.051
R770 VSS.t785 VSS.t2249 767.051
R771 VSS.t1133 VSS.t77 767.051
R772 VSS.t1396 VSS.t54 767.051
R773 VSS.t842 VSS.t634 767.051
R774 VSS.t1677 VSS.t347 767.051
R775 VSS.t1000 VSS.t1892 767.051
R776 VSS.t1892 VSS.t632 767.051
R777 VSS.t1598 VSS.t2239 767.051
R778 VSS.t1228 VSS.t2233 767.051
R779 VSS.t2216 VSS.t183 767.051
R780 VSS.t189 VSS.t2111 767.051
R781 VSS.t856 VSS.t173 767.051
R782 VSS.t2120 VSS.t181 767.051
R783 VSS.n1023 VSS.t1920 761.157
R784 VSS.t3039 VSS.t651 758.621
R785 VSS.t3011 VSS.t2247 758.621
R786 VSS.t1460 VSS.t3045 758.621
R787 VSS.t2035 VSS.t3127 758.621
R788 VSS.t1305 VSS.t870 758.621
R789 VSS.t723 VSS.n1436 758.621
R790 VSS.t577 VSS.t480 750.192
R791 VSS.t413 VSS.t1879 750.192
R792 VSS.t1886 VSS.t3476 750.192
R793 VSS.t1332 VSS.t2227 750.192
R794 VSS.t201 VSS.t753 741.763
R795 VSS.t2864 VSS.t2717 741.763
R796 VSS.t2194 VSS.t2139 741.763
R797 VSS.t2709 VSS.t2872 741.763
R798 VSS.t99 VSS.t1832 741.763
R799 VSS.t2922 VSS.t1505 741.763
R800 VSS.t38 VSS.t2182 741.763
R801 VSS.t492 VSS.t843 733.333
R802 VSS.t2090 VSS.t868 733.333
R803 VSS.t587 VSS.t214 733.333
R804 VSS.t1989 VSS.t580 733.333
R805 VSS.t1224 VSS.t2108 733.333
R806 VSS.n992 VSS.t881 731.062
R807 VSS.t3244 VSS.n4649 729.404
R808 VSS.n1195 VSS.t3396 729.404
R809 VSS.t834 VSS.t1044 724.904
R810 VSS.t1666 VSS.t1336 724.904
R811 VSS.t2656 VSS.t2654 724.904
R812 VSS.t2654 VSS.t2650 724.904
R813 VSS.t1209 VSS.t1213 724.904
R814 VSS.t2889 VSS.t576 724.904
R815 VSS.t576 VSS.t654 724.904
R816 VSS.t2274 VSS.t494 724.904
R817 VSS.t510 VSS.t1816 724.904
R818 VSS.t140 VSS.t134 724.904
R819 VSS.t134 VSS.t136 724.904
R820 VSS.t1407 VSS.t563 724.904
R821 VSS.t2891 VSS.t640 724.904
R822 VSS.t3229 VSS.t1008 724.904
R823 VSS.t684 VSS.t1672 724.904
R824 VSS.t910 VSS.t790 724.904
R825 VSS.t1076 VSS.t2581 716.476
R826 VSS.t2763 VSS.t995 716.476
R827 VSS.t2027 VSS.t892 716.476
R828 VSS.t83 VSS.t1703 716.476
R829 VSS.n5179 VSS.t3217 709.346
R830 VSS.t1768 VSS.t1770 708.047
R831 VSS.t1772 VSS.t1768 708.047
R832 VSS.t1766 VSS.t1772 708.047
R833 VSS.t1599 VSS.t2125 708.047
R834 VSS.t1843 VSS.t2693 708.047
R835 VSS.t1203 VSS.t1201 708.047
R836 VSS.t1138 VSS.t1136 708.047
R837 VSS.t1090 VSS.t1042 708.047
R838 VSS.t1042 VSS.t2613 708.047
R839 VSS.t2102 VSS.t2104 708.047
R840 VSS.t1436 VSS.t1837 708.047
R841 VSS.t1853 VSS.t1363 708.047
R842 VSS.t876 VSS.t209 708.047
R843 VSS.t488 VSS.t591 708.047
R844 VSS.t1730 VSS.t589 708.047
R845 VSS.t772 VSS.t1666 708.047
R846 VSS.t484 VSS.t490 708.047
R847 VSS.t1120 VSS.t1722 708.047
R848 VSS.n4056 VSS.t2998 708.047
R849 VSS.t12 VSS.t218 708.047
R850 VSS.t1525 VSS.t599 708.047
R851 VSS.t1524 VSS.t2860 708.047
R852 VSS.t2860 VSS.t2723 708.047
R853 VSS.t788 VSS.t44 708.047
R854 VSS.t44 VSS.t1789 708.047
R855 VSS.t1812 VSS.t1814 708.047
R856 VSS.t1869 VSS.t158 708.047
R857 VSS.t158 VSS.t2710 708.047
R858 VSS.t1251 VSS.t1253 708.047
R859 VSS.t1514 VSS.t1510 708.047
R860 VSS.t2146 VSS.t2144 708.047
R861 VSS.t1319 VSS.t1317 708.047
R862 VSS.t2072 VSS.t973 708.047
R863 VSS.t1592 VSS.t387 708.047
R864 VSS.t1798 VSS.t1802 708.047
R865 VSS.t1678 VSS.t417 708.047
R866 VSS.t2223 VSS.t2221 708.047
R867 VSS.t2219 VSS.t2217 708.047
R868 VSS.t1146 VSS.t1144 708.047
R869 VSS.t949 VSS.t947 708.047
R870 VSS.t733 VSS.t731 708.047
R871 VSS.t1669 VSS.t1667 708.047
R872 VSS.t2128 VSS.t2126 708.047
R873 VSS.t1353 VSS.t1355 708.047
R874 VSS.t874 VSS.t872 708.047
R875 VSS.t2964 VSS.t2962 708.047
R876 VSS.t680 VSS.t645 708.047
R877 VSS.t2615 VSS.t2611 708.047
R878 VSS.t1849 VSS.t1851 708.047
R879 VSS.t1140 VSS.t42 708.047
R880 VSS.t383 VSS.t1373 708.047
R881 VSS.t475 VSS.t1501 708.047
R882 VSS.t607 VSS.t602 708.047
R883 VSS.t1664 VSS.t1875 708.047
R884 VSS.t1503 VSS.t2075 708.047
R885 VSS.t1793 VSS.t969 708.047
R886 VSS.t969 VSS.t970 708.047
R887 VSS.t2909 VSS.t401 708.047
R888 VSS.t2 VSS.t0 708.047
R889 VSS.t2852 VSS.t814 708.047
R890 VSS.t814 VSS.t815 708.047
R891 VSS.t1179 VSS.t154 708.047
R892 VSS.t154 VSS.t4 708.047
R893 VSS.t2578 VSS.t28 708.047
R894 VSS.t1526 VSS.t1528 708.047
R895 VSS.t2923 VSS.t2916 708.047
R896 VSS.t148 VSS.t150 708.047
R897 VSS.t150 VSS.t730 708.047
R898 VSS.t730 VSS.t729 708.047
R899 VSS.t1315 VSS.t2911 708.047
R900 VSS.t2263 VSS.t993 708.047
R901 VSS.t2162 VSS.t2160 708.047
R902 VSS.t207 VSS.t2272 708.047
R903 VSS.t1830 VSS.t1827 708.047
R904 VSS.t1465 VSS.t1594 708.047
R905 VSS.t2747 VSS.t164 708.047
R906 VSS.t2753 VSS.t2727 708.047
R907 VSS.t1877 VSS.t391 708.047
R908 VSS.t71 VSS.t73 708.047
R909 VSS.t360 VSS.t362 708.047
R910 VSS.t2788 VSS.t2792 708.047
R911 VSS.t1450 VSS.t1448 708.047
R912 VSS.t1656 VSS.t1654 708.047
R913 VSS.t1124 VSS.t1122 708.047
R914 VSS.t522 VSS.t525 708.047
R915 VSS.t107 VSS.t109 708.047
R916 VSS.t2557 VSS.t2555 708.047
R917 VSS.t1861 VSS.t1865 708.047
R918 VSS.t1865 VSS.t1859 708.047
R919 VSS.t1859 VSS.t1863 708.047
R920 VSS.t1357 VSS.t1359 708.047
R921 VSS.t700 VSS.t1432 708.047
R922 VSS.t1371 VSS.t1969 708.047
R923 VSS.t2885 VSS.t2862 708.047
R924 VSS.t1266 VSS.t1267 708.047
R925 VSS.t1756 VSS.t1754 708.047
R926 VSS.t1727 VSS.t568 708.047
R927 VSS.t572 VSS.t1881 708.047
R928 VSS.t2123 VSS.t2121 708.047
R929 VSS.t1270 VSS.t379 708.047
R930 VSS.t162 VSS.t2866 708.047
R931 VSS.t845 VSS.t1070 708.047
R932 VSS.t766 VSS.t2571 708.047
R933 VSS.t2571 VSS.t583 708.047
R934 VSS.t1774 VSS.t1776 708.047
R935 VSS.t26 VSS.t2641 708.047
R936 VSS.t1014 VSS.t160 708.047
R937 VSS.t160 VSS.t216 708.047
R938 VSS.t847 VSS.t585 708.047
R939 VSS.t2265 VSS.t2596 708.047
R940 VSS.t2596 VSS.t1588 708.047
R941 VSS.t1533 VSS.t1535 708.047
R942 VSS.t1508 VSS.t385 708.047
R943 VSS.t385 VSS.t807 708.047
R944 VSS.t2918 VSS.t2229 708.047
R945 VSS.t210 VSS.t1605 708.047
R946 VSS.t975 VSS.t915 708.047
R947 VSS.t1424 VSS.t975 708.047
R948 VSS.t717 VSS.t719 708.047
R949 VSS.t235 VSS.t271 708.047
R950 VSS.t239 VSS.t235 708.047
R951 VSS.t1822 VSS.t1821 708.047
R952 VSS.t1466 VSS.t1467 708.047
R953 VSS.t1467 VSS.t2039 708.047
R954 VSS.t2039 VSS.t2040 708.047
R955 VSS.t1148 VSS.t1462 708.047
R956 VSS.t1154 VSS.t1152 708.047
R957 VSS.t1689 VSS.t1691 708.047
R958 VSS.t1691 VSS.t1787 708.047
R959 VSS.t1787 VSS.t1786 708.047
R960 VSS.t393 VSS.t1220 708.047
R961 VSS.t381 VSS.t1177 708.047
R962 VSS.t91 VSS.t381 708.047
R963 VSS.t825 VSS.t820 708.047
R964 VSS.t1653 VSS.t825 708.047
R965 VSS.t1652 VSS.t1653 708.047
R966 VSS.t130 VSS.t132 708.047
R967 VSS.t303 VSS.t299 708.047
R968 VSS.t2847 VSS.t2901 708.047
R969 VSS.t743 VSS.t741 708.047
R970 VSS.t937 VSS.t935 708.047
R971 VSS.t1454 VSS.t1452 708.047
R972 VSS.t2858 VSS.t2856 708.047
R973 VSS.t2013 VSS.t2015 708.047
R974 VSS.t355 VSS.t357 708.047
R975 VSS.t1943 VSS.t1941 708.047
R976 VSS.t1092 VSS.t1094 708.047
R977 VSS.t1631 VSS.t1629 708.047
R978 VSS.t1935 VSS.t1428 708.047
R979 VSS.t1956 VSS.t1962 708.047
R980 VSS.t531 VSS.t2719 708.047
R981 VSS.t1929 VSS.t1430 708.047
R982 VSS.t1247 VSS.t1241 708.047
R983 VSS.t1307 VSS.t1309 708.047
R984 VSS.t1157 VSS.t32 708.047
R985 VSS.t1168 VSS.t1164 708.047
R986 VSS.t1166 VSS.t1170 708.047
R987 VSS.t2576 VSS.t2575 708.047
R988 VSS.t2179 VSS.t30 708.047
R989 VSS.t579 VSS.t470 708.047
R990 VSS.t963 VSS.t959 708.047
R991 VSS.t1009 VSS.t203 708.047
R992 VSS.t535 VSS.t1823 708.047
R993 VSS.t2206 VSS.t2202 708.047
R994 VSS.t2202 VSS.t2204 708.047
R995 VSS.t1484 VSS.t1482 708.047
R996 VSS.t2099 VSS.t425 708.047
R997 VSS.t907 VSS.t419 708.047
R998 VSS.t593 VSS.t595 708.047
R999 VSS.t676 VSS.t678 708.047
R1000 VSS.t803 VSS.t805 708.047
R1001 VSS.t945 VSS.t943 708.047
R1002 VSS.n1193 VSS.t3396 705.898
R1003 VSS.t2009 VSS.t2007 700.333
R1004 VSS.t1085 VSS.t462 699.617
R1005 VSS.t645 VSS.t704 699.617
R1006 VSS.t2183 VSS.t2973 699.617
R1007 VSS.t322 VSS.t1522 699.617
R1008 VSS.t2682 VSS.t1728 699.617
R1009 VSS.t1991 VSS.t2782 699.617
R1010 VSS.t434 VSS.t737 699.617
R1011 VSS.t939 VSS.t1752 699.617
R1012 VSS.t2927 VSS.t832 699.617
R1013 VSS.t113 VSS.t1349 696.668
R1014 VSS.t2093 VSS.t1237 696.668
R1015 VSS.t1601 VSS.t1442 693
R1016 VSS.t460 VSS.t2676 693
R1017 VSS.t2652 VSS.t2188 691.188
R1018 VSS.t3245 VSS.t36 691.188
R1019 VSS.t2707 VSS.t1546 691.188
R1020 VSS.t2714 VSS.t489 691.188
R1021 VSS.t1792 VSS.t482 691.188
R1022 VSS.t3436 VSS.t624 691.188
R1023 VSS.t315 VSS.t1243 691.188
R1024 VSS.t1225 VSS.t374 691.188
R1025 VSS.t2982 VSS.t2790 689.333
R1026 VSS.t2845 VSS.t103 689.333
R1027 VSS.t919 VSS.t113 689.333
R1028 VSS.t320 VSS.t20 689.333
R1029 VSS.t1426 VSS.t3405 682.76
R1030 VSS.t2067 VSS.t389 682.76
R1031 VSS.t689 VSS.t3411 682.76
R1032 VSS.t1707 VSS.t1156 682.76
R1033 VSS.t2951 VSS.n977 681.093
R1034 VSS.t3079 VSS.n19 674.668
R1035 VSS.t1399 VSS.t1207 674.331
R1036 VSS.t1545 VSS.t1072 674.331
R1037 VSS.t3010 VSS.t2037 674.331
R1038 VSS.t3006 VSS.t3007 674.331
R1039 VSS.t1197 VSS.t100 674.331
R1040 VSS.t2905 VSS.t409 674.331
R1041 VSS.t547 VSS.t138 674.331
R1042 VSS.t1132 VSS.t571 674.331
R1043 VSS.t1562 VSS.t1960 674.331
R1044 VSS.t1264 VSS.t1249 674.331
R1045 VSS.t1724 VSS.t684 674.331
R1046 VSS.t2893 VSS.t696 665.9
R1047 VSS.t1129 VSS.t2079 665.9
R1048 VSS.t1639 VSS.t1472 665.9
R1049 VSS.t1135 VSS.t1301 665.9
R1050 VSS.t1825 VSS.t46 665.9
R1051 VSS.t1343 VSS.t1788 665.9
R1052 VSS.t2153 VSS.t2757 665.9
R1053 VSS.t2159 VSS.t1794 665.9
R1054 VSS.t1682 VSS.t826 665.9
R1055 VSS.t1036 VSS.t1024 665.9
R1056 VSS.t2226 VSS.t1985 665.9
R1057 VSS.t403 VSS.t2114 665.9
R1058 VSS.t1413 VSS.t507 665.9
R1059 VSS.n1054 VSS.t693 665.087
R1060 VSS.t2142 VSS.t1579 657.471
R1061 VSS.t917 VSS.t1440 657.471
R1062 VSS.n1436 VSS.t1046 657.471
R1063 VSS.t1541 VSS.t1018 649.181
R1064 VSS.t2563 VSS.t289 649.181
R1065 VSS.t1187 VSS.t118 649.043
R1066 VSS.t2849 VSS.t3027 649.043
R1067 VSS.t764 VSS.t341 649.043
R1068 VSS.t2887 VSS.t2850 649.043
R1069 VSS.t1290 VSS.t152 649.043
R1070 VSS.t1559 VSS.t1702 649.043
R1071 VSS.t694 VSS.t2601 645.745
R1072 VSS.t541 VSS.t899 645.745
R1073 VSS.t1695 VSS.t223 644.237
R1074 VSS.t786 VSS.t834 640.614
R1075 VSS.t1493 VSS.t574 640.614
R1076 VSS.t756 VSS.t399 640.614
R1077 VSS.t2868 VSS.t1261 640.614
R1078 VSS.t508 VSS.t10 640.614
R1079 VSS.t2873 VSS.t505 640.614
R1080 VSS.t339 VSS.t3157 640.614
R1081 VSS.n1488 VSS.t1361 640.614
R1082 VSS.t1651 VSS.t1305 640.614
R1083 VSS.t1674 VSS.t1162 640.614
R1084 VSS.t2148 VSS.t2573 640.614
R1085 VSS.t81 VSS.t721 640.614
R1086 VSS.t1012 VSS.t545 640.614
R1087 VSS.t1506 VSS.t504 640.614
R1088 VSS.t507 VSS.t95 640.614
R1089 VSS.t3520 VSS.t1884 635.67
R1090 VSS.t3204 VSS.t2700 633.957
R1091 VSS.t3217 VSS.t2933 633.957
R1092 VSS.t1873 VSS.t3520 633.957
R1093 VSS.t920 VSS.t1977 632.184
R1094 VSS.t1102 VSS.t2019 632.184
R1095 VSS.t216 VSS.t885 632.184
R1096 VSS.t2181 VSS.t581 632.184
R1097 VSS.t2214 VSS.t1504 632.184
R1098 VSS.n196 VSS.t3408 632.006
R1099 VSS.t2253 VSS.t2170 623.755
R1100 VSS.t2254 VSS.t2171 623.755
R1101 VSS.t1211 VSS.t894 623.755
R1102 VSS.t1142 VSS.t1732 623.755
R1103 VSS.t1052 VSS.t2598 623.755
R1104 VSS.t2634 VSS.t225 623.755
R1105 VSS.t3452 VSS.t1643 623.755
R1106 VSS.t2235 VSS.t2812 623.755
R1107 VSS.t1164 VSS.t1531 623.755
R1108 VSS.n1221 VSS.t883 618.003
R1109 VSS.t1995 VSS.t1583 615.327
R1110 VSS.t1016 VSS.t2640 615.327
R1111 VSS.t2729 VSS.t3503 615.327
R1112 VSS.t632 VSS.t1674 615.327
R1113 VSS.t610 VSS.t493 606.898
R1114 VSS.t493 VSS.t653 606.898
R1115 VSS.t2069 VSS.t474 606.898
R1116 VSS.t1871 VSS.t3402 606.898
R1117 VSS.t2777 VSS.t1331 606.898
R1118 VSS.t1895 VSS.t813 606.898
R1119 VSS.t1089 VSS.t2245 606.898
R1120 VSS.t175 VSS.t811 606.898
R1121 VSS.t171 VSS.t2589 606.898
R1122 VSS.t187 VSS.t887 606.898
R1123 VSS.t760 VSS.t24 606.898
R1124 VSS.t2645 VSS.t2237 606.898
R1125 VSS.t152 VSS.t2241 606.898
R1126 VSS.t3166 VSS.t1396 606.898
R1127 VSS.t349 VSS.t1532 606.898
R1128 VSS.t2243 VSS.t914 606.898
R1129 VSS.t1478 VSS.t792 606.898
R1130 VSS.t2773 VSS.t1724 606.898
R1131 VSS.t1217 VSS.t423 606.898
R1132 VSS.t177 VSS.t1219 606.898
R1133 VSS.t185 VSS.t880 606.898
R1134 VSS.t2827 VSS.t1762 606.898
R1135 VSS.t2610 VSS.t421 598.467
R1136 VSS.t375 VSS.t151 598.467
R1137 VSS.t2712 VSS.t1647 598.467
R1138 VSS.t2599 VSS.t377 598.467
R1139 VSS.t1199 VSS.t1709 598.467
R1140 VSS.t498 VSS.t415 598.467
R1141 VSS.t703 VSS.t1107 598.467
R1142 VSS.t1970 VSS.t1357 598.467
R1143 VSS.t513 VSS.t1908 598.467
R1144 VSS.t395 VSS.t265 598.467
R1145 VSS.t1810 VSS.t582 598.467
R1146 VSS.n4969 VSS.t2670 597.412
R1147 VSS.t1456 VSS.t1327 591.211
R1148 VSS.t1927 VSS.t1286 590.038
R1149 VSS.t1470 VSS.t911 590.038
R1150 VSS.t851 VSS.t2577 590.038
R1151 VSS.t2761 VSS.t1340 590.038
R1152 VSS.n2954 VSS.t759 590.038
R1153 VSS.t759 VSS.t169 590.038
R1154 VSS.t1022 VSS.t2187 590.038
R1155 VSS.t1863 VSS.t3109 590.038
R1156 VSS.t840 VSS.t1247 590.038
R1157 VSS.t838 VSS.t1245 590.038
R1158 VSS.t589 VSS.t2805 581.61
R1159 VSS.t1207 VSS.t2779 581.61
R1160 VSS.n4241 VSS.t2610 581.61
R1161 VSS.t2137 VSS.t2749 581.61
R1162 VSS.t1303 VSS.t949 581.61
R1163 VSS.t827 VSS.t3139 581.61
R1164 VSS.t1405 VSS.t1937 581.61
R1165 VSS.t54 VSS.t1562 581.61
R1166 VSS.t634 VSS.t1264 581.61
R1167 VSS.n1107 VSS.n1106 575.024
R1168 VSS.t1949 VSS.t1842 573.181
R1169 VSS.t115 VSS.t2888 573.181
R1170 VSS.t337 VSS.t628 573.181
R1171 VSS.t621 VSS.t2999 573.181
R1172 VSS.t275 VSS.t1833 573.181
R1173 VSS.t1560 VSS.t79 573.181
R1174 VSS.t2204 VSS.t1003 573.181
R1175 VSS.t2208 VSS.t212 573.181
R1176 VSS.n1253 VSS.n461 565.554
R1177 VSS.n1259 VSS.n1258 565.554
R1178 VSS.t1363 VSS.t1280 564.751
R1179 VSS.t1722 VSS.t1658 564.751
R1180 VSS.t614 VSS.t1552 564.751
R1181 VSS.n4797 VSS.n477 562.729
R1182 VSS.t2739 VSS.t2949 561.201
R1183 VSS.t2939 VSS.t199 561.201
R1184 VSS.n316 VSS.t3641 557.02
R1185 VSS.n311 VSS.t3728 557.013
R1186 VSS.n316 VSS.t3692 556.54
R1187 VSS.n314 VSS.t3625 556.54
R1188 VSS.n315 VSS.t3798 556.54
R1189 VSS.n313 VSS.t3649 556.54
R1190 VSS.n312 VSS.t3792 556.54
R1191 VSS.n311 VSS.t3788 556.54
R1192 VSS.t1278 VSS.t1345 556.322
R1193 VSS.t1275 VSS.t1737 556.322
R1194 VSS.t783 VSS.t2996 556.322
R1195 VSS.t1191 VSS.t2271 556.322
R1196 VSS.t2074 VSS.t996 556.322
R1197 VSS.t1110 VSS.n2257 556.322
R1198 VSS.t1932 VSS.t1434 556.322
R1199 VSS.n1066 VSS.t231 555.14
R1200 VSS.n5178 VSS.t3175 551.713
R1201 VSS.t209 VSS.t636 547.894
R1202 VSS.t812 VSS.t2026 547.894
R1203 VSS.t1910 VSS.t2587 547.894
R1204 VSS.t2618 VSS.t2644 547.894
R1205 VSS.t2249 VSS.t2918 547.894
R1206 VSS.t1966 VSS.t918 547.894
R1207 VSS.t1377 VSS.t836 547.894
R1208 VSS.t2141 VSS.t233 547.894
R1209 VSS.t1890 VSS.t3426 547.894
R1210 VSS.t1060 VSS.n79 542.668
R1211 VSS.t496 VSS.t2816 539.465
R1212 VSS.t2158 VSS.t2096 539.465
R1213 VSS.t568 VSS.t1725 539.465
R1214 VSS.t1703 VSS.t1560 539.465
R1215 VSS.t1361 VSS.t776 539.465
R1216 VSS.t630 VSS.t1311 539.465
R1217 VSS.t1104 VSS.t2576 539.465
R1218 VSS.n1071 VSS.n1069 538.28
R1219 VSS.t1080 VSS.t809 531.034
R1220 VSS.t1945 VSS.t566 531.034
R1221 VSS.t820 VSS.t2765 531.034
R1222 VSS.t1633 VSS.t2957 531.034
R1223 VSS.t1635 VSS.t1782 531.034
R1224 VSS.t1617 VSS.t2055 531.034
R1225 VSS.t1623 VSS.t2057 531.034
R1226 VSS.n318 VSS.t2488 526.735
R1227 VSS.n322 VSS.t2415 526.552
R1228 VSS.n3715 VSS.t2219 522.606
R1229 VSS.t1035 VSS.t1640 522.606
R1230 VSS.t2903 VSS.t802 522.606
R1231 VSS.t1690 VSS.t1037 522.606
R1232 VSS.t1046 VSS.t2212 522.606
R1233 VSS.t1611 VSS.n59 520.668
R1234 VSS.n5355 VSS.t1028 517
R1235 VSS.t1581 VSS.n37 517
R1236 VSS.t951 VSS.n4585 517
R1237 VSS.t1984 VSS.t2119 514.177
R1238 VSS.t1983 VSS.t2118 514.177
R1239 VSS.t1257 VSS.t1572 514.177
R1240 VSS.t1629 VSS.t267 514.177
R1241 VSS.t48 VSS.t781 514.177
R1242 VSS.n5355 VSS.t1857 513.333
R1243 VSS.t1098 VSS.n158 513.333
R1244 VSS.n139 VSS.t1403 513.333
R1245 VSS.t197 VSS.t446 509.325
R1246 VSS.t1952 VSS.t2168 505.748
R1247 VSS.t2251 VSS.t755 505.748
R1248 VSS.t116 VSS.t1692 505.748
R1249 VSS.t1261 VSS.t3473 505.748
R1250 VSS.t1820 VSS.t261 505.748
R1251 VSS.t512 VSS.t1822 505.748
R1252 VSS.t1712 VSS.t2021 505.748
R1253 VSS.t423 VSS.t177 505.748
R1254 VSS.t824 VSS.t405 505.748
R1255 VSS.t466 VSS.t533 505.748
R1256 VSS.t1762 VSS.t907 505.748
R1257 VSS.t996 VSS.t3011 497.318
R1258 VSS.t811 VSS.t510 497.318
R1259 VSS.t1131 VSS.t647 497.318
R1260 VSS.t1338 VSS.t2101 497.318
R1261 VSS.t445 VSS.n950 490.298
R1262 VSS.t552 VSS.n1237 490.298
R1263 VSS.t1804 VSS.t2095 488.889
R1264 VSS.t345 VSS.t2025 488.889
R1265 VSS.t1552 VSS.t853 488.889
R1266 VSS.t2237 VSS.t3452 488.889
R1267 VSS.t2812 VSS.t928 488.889
R1268 VSS.t1596 VSS.t509 488.889
R1269 VSS.t2111 VSS.t1480 488.889
R1270 VSS.t16 VSS.t2968 486.604
R1271 VSS.t1215 VSS.t3148 485.212
R1272 VSS.n1067 VSS.t2971 482.099
R1273 VSS.t19 VSS.n1075 482.099
R1274 VSS.t3001 VSS.t2029 480.461
R1275 VSS.t3535 VSS.t1872 480.461
R1276 VSS.t1365 VSS.t866 480.461
R1277 VSS.t1476 VSS.t1671 480.461
R1278 VSS.t539 VSS.t1570 479.752
R1279 VSS.t458 VSS.t3175 476.325
R1280 VSS.t1118 VSS.t2798 472.031
R1281 VSS.t574 VSS.t351 472.031
R1282 VSS.t1050 VSS.t1748 472.031
R1283 VSS.t2866 VSS.n2259 472.031
R1284 VSS.n2736 VSS.t2229 472.031
R1285 VSS.t1505 VSS.t865 472.031
R1286 VSS.t3139 VSS.t619 472.031
R1287 VSS.t2573 VSS.t327 472.031
R1288 VSS.t959 VSS.t527 472.031
R1289 VSS.t965 VSS.t2920 472.031
R1290 VSS.t545 VSS.t2231 472.031
R1291 VSS.t914 VSS.t535 472.031
R1292 VSS.t1219 VSS.t1100 472.031
R1293 VSS.t1553 VSS.t764 463.603
R1294 VSS.t2160 VSS.t1557 463.603
R1295 VSS.t2043 VSS.t1568 463.603
R1296 VSS.t1555 VSS.t2092 463.603
R1297 VSS.t93 VSS.t821 463.603
R1298 VSS.t1979 VSS.t222 463.603
R1299 VSS.t421 VSS.t2595 455.173
R1300 VSS.t1579 VSS.t191 455.173
R1301 VSS.t1034 VSS.t375 455.173
R1302 VSS.t1193 VSS.t2580 455.173
R1303 VSS.t2092 VSS.t1199 455.173
R1304 VSS.t821 VSS.t1810 455.173
R1305 VSS.n1018 VSS.t3204 452.337
R1306 VSS.t199 VSS.n992 451.998
R1307 VSS.t197 VSS.n1209 451.998
R1308 VSS.n1209 VSS.t446 451.998
R1309 VSS.t343 VSS.t2893 446.743
R1310 VSS.t1495 VSS.t1765 446.743
R1311 VSS.t1259 VSS.t572 446.743
R1312 VSS.t796 VSS.t2891 446.743
R1313 VSS.t327 VSS.t227 446.743
R1314 VSS.t2704 VSS.t3015 439.368
R1315 VSS.t2798 VSS.t712 438.315
R1316 VSS.t1681 VSS.t3535 438.315
R1317 VSS.t1748 VSS.t475 438.315
R1318 VSS.t1501 VSS.t2044 438.315
R1319 VSS.t167 VSS.t1817 438.315
R1320 VSS.t1220 VSS.n2835 438.315
R1321 VSS.t1720 VSS.t243 438.315
R1322 VSS.t2110 VSS.t1476 438.315
R1323 VSS.t1918 VSS.n1021 431.373
R1324 VSS.t1915 VSS.t1911 431.373
R1325 VSS.t1911 VSS.t1918 431.373
R1326 VSS.t872 VSS.t3433 429.885
R1327 VSS.t1603 VSS.t3238 423.147
R1328 VSS.t1662 VSS.t1800 421.457
R1329 VSS.t502 VSS.t1134 421.457
R1330 VSS.t468 VSS.t2225 421.457
R1331 VSS.t865 VSS.t166 421.457
R1332 VSS.t625 VSS.t2214 421.457
R1333 VSS.t70 VSS.n5348 417.125
R1334 VSS.t1958 VSS.t642 413.027
R1335 VSS.t1625 VSS.t1195 413.027
R1336 VSS.t1619 VSS.t1687 413.027
R1337 VSS.n3869 VSS.t75 404.599
R1338 VSS.n3229 VSS.t2929 404.599
R1339 VSS.t1038 VSS.t317 404.599
R1340 VSS.n2355 VSS.t1933 404.599
R1341 VSS.t6 VSS.n2258 404.599
R1342 VSS.n2737 VSS.t1150 404.599
R1343 VSS.t3214 VSS.t2873 404.599
R1344 VSS.n1575 VSS.t1397 404.599
R1345 VSS.t957 VSS.t963 404.599
R1346 VSS.t3193 VSS.t1506 404.599
R1347 VSS.t2913 VSS.t1720 404.599
R1348 VSS.t425 VSS.t3488 404.599
R1349 VSS.t533 VSS.t854 404.599
R1350 VSS.t1954 VSS.t570 396.17
R1351 VSS.t472 VSS.t1972 396
R1352 VSS.t3517 VSS.t2689 387.808
R1353 VSS.t1947 VSS.t1126 387.74
R1354 VSS.t2585 VSS.t1251 387.74
R1355 VSS.t1800 VSS.t1423 387.74
R1356 VSS.t3187 VSS.t3070 387.74
R1357 VSS.t623 VSS.t1129 387.74
R1358 VSS.n3230 VSS.t3198 387.74
R1359 VSS.t3190 VSS.n3033 387.74
R1360 VSS.t1464 VSS.t1343 387.74
R1361 VSS.t615 VSS.t1682 387.74
R1362 VSS.t1953 VSS.t564 387.74
R1363 VSS.t1745 VSS.t1750 370.961
R1364 VSS.t712 VSS.t115 370.882
R1365 VSS.t429 VSS.n4492 370.882
R1366 VSS.t3433 VSS.t1321 370.882
R1367 VSS.t2044 VSS.t1367 370.882
R1368 VSS.n3081 VSS.t2801 370.882
R1369 VSS.t758 VSS.t1910 370.882
R1370 VSS.t1725 VSS.t1259 370.882
R1371 VSS.t1821 VSS.t1829 370.882
R1372 VSS.t1784 VSS.t1631 370.882
R1373 VSS.t1931 VSS.t1966 370.882
R1374 VSS.t776 VSS.t1377 370.882
R1375 VSS.t1512 VSS.t778 370.882
R1376 VSS.t880 VSS.t818 370.882
R1377 VSS.t427 VSS.n2068 370.882
R1378 VSS.n1084 VSS.n1083 369.245
R1379 VSS.n1065 VSS.t2416 366.668
R1380 VSS.n1055 VSS.t2489 366.668
R1381 VSS.t2660 VSS.t2658 365.579
R1382 VSS.t2658 VSS.t2664 365.579
R1383 VSS.t2664 VSS.t2662 365.579
R1384 VSS.t881 VSS.t883 365.579
R1385 VSS.n4936 VSS.t3015 364.034
R1386 VSS.t3067 VSS.t1743 362.452
R1387 VSS.t1053 VSS.t1191 362.452
R1388 VSS.t97 VSS.t708 362.452
R1389 VSS.t1334 VSS.t2803 359.334
R1390 VSS.t1349 VSS.t478 359.334
R1391 VSS.n1188 VSS.n1014 356.894
R1392 VSS.n4653 VSS.n1241 356.894
R1393 VSS.t3004 VSS.t1056 355.668
R1394 VSS.t1233 VSS.t1615 355.668
R1395 VSS.t1900 VSS.t955 355.668
R1396 VSS.t1419 VSS.t1581 355.668
R1397 VSS.t2051 VSS.t1394 355.668
R1398 VSS.t859 VSS.t2009 355.668
R1399 VSS.t2003 VSS.t951 355.668
R1400 VSS.t1380 VSS.t2093 355.668
R1401 VSS.t1577 VSS.t2156 354.024
R1402 VSS.t1078 VSS.t1193 354.024
R1403 VSS.t2580 VSS.t614 354.024
R1404 VSS.t1557 VSS.t2593 354.024
R1405 VSS.t1392 VSS.n1510 354.024
R1406 VSS.n1085 VSS.n1032 353.882
R1407 VSS.n1087 VSS.n1084 353.882
R1408 VSS.n3944 VSS.n3943 352
R1409 VSS.n3447 VSS.n3445 352
R1410 VSS.n1987 VSS.n1986 352
R1411 VSS.t111 VSS.t2799 352
R1412 VSS.t2790 VSS.t1758 348.334
R1413 VSS.t1030 VSS.t2845 348.334
R1414 VSS.t144 VSS.t1096 348.334
R1415 VSS.t142 VSS.t1172 348.334
R1416 VSS.t1442 VSS.t1446 348.334
R1417 VSS.t2674 VSS.t320 348.334
R1418 VSS.t1239 VSS.t460 348.334
R1419 VSS.n1103 VSS.n1102 347.404
R1420 VSS.n1103 VSS.n1024 347.301
R1421 VSS.t1741 VSS.t3067 345.594
R1422 VSS.t351 VSS.t1734 345.594
R1423 VSS.t853 VSS.t1553 345.594
R1424 VSS.t1568 VSS.t1555 345.594
R1425 VSS.n2259 VSS.t739 345.594
R1426 VSS.t708 VSS.t93 345.594
R1427 VSS.t1468 VSS.t3130 338.885
R1428 VSS.t3414 VSS.t971 338.885
R1429 VSS.n5349 VSS.t1599 337.166
R1430 VSS.t2217 VSS.t2745 337.166
R1431 VSS.n4492 VSS.t1641 337.166
R1432 VSS.t1181 VSS.t849 337.166
R1433 VSS.t626 VSS.t1736 337.166
R1434 VSS.t2883 VSS.t1727 337.166
R1435 VSS.t1608 VSS.n2736 337.166
R1436 VSS.t1829 VSS.t1820 337.166
R1437 VSS.n2068 VSS.t2259 337.166
R1438 VSS.n1182 VSS.n1014 333.628
R1439 VSS.n4634 VSS.n1241 333.628
R1440 VSS.n1184 VSS.t3251 332.024
R1441 VSS.t3244 VSS.n1245 330.818
R1442 VSS.n1245 VSS.t3054 330.818
R1443 VSS.t1126 VSS.t1496 328.736
R1444 VSS.t2029 VSS.t620 328.736
R1445 VSS.t52 VSS.t2895 328.736
R1446 VSS.t1018 VSS.t926 326.308
R1447 VSS.t1539 VSS.t1543 326.308
R1448 VSS.t2601 VSS.t2603 326.308
R1449 VSS.t1292 VSS.t2255 326.308
R1450 VSS.t2561 VSS.t2565 326.308
R1451 VSS.t899 VSS.t901 326.308
R1452 VSS.n1235 VSS.n478 324.589
R1453 VSS.t727 VSS.t2200 323.832
R1454 VSS.t1857 VSS.t2982 322.668
R1455 VSS.t103 VSS.t1081 322.668
R1456 VSS.t2725 VSS.t1739 322.668
R1457 VSS.t1489 VSS.t2086 322.668
R1458 VSS.t1403 VSS.t2083 322.668
R1459 VSS.t2960 VSS.t2061 322.668
R1460 VSS.t2818 VSS.t1601 322.668
R1461 VSS.t20 VSS.t685 322.668
R1462 VSS.t1112 VSS.t543 322.118
R1463 VSS.t514 VSS.t14 322.118
R1464 VSS.t1286 VSS.t1118 320.307
R1465 VSS.t1893 VSS.t1120 320.307
R1466 VSS.t2119 VSS.t2154 320.307
R1467 VSS.t1627 VSS.t1983 320.307
R1468 VSS.t1253 VSS.t3001 320.307
R1469 VSS.t1423 VSS.t1804 320.307
R1470 VSS.t2577 VSS.t1365 320.307
R1471 VSS.t62 VSS.t1954 320.307
R1472 VSS.t509 VSS.t1011 320.307
R1473 VSS.t1056 VSS.t1058 315.334
R1474 VSS.t1058 VSS.t1054 315.334
R1475 VSS.t1054 VSS.t1060 315.334
R1476 VSS.t1235 VSS.t1229 315.334
R1477 VSS.t1229 VSS.t1231 315.334
R1478 VSS.t1231 VSS.t1233 315.334
R1479 VSS.t1904 VSS.t1898 315.334
R1480 VSS.t1898 VSS.t1902 315.334
R1481 VSS.t1902 VSS.t1900 315.334
R1482 VSS.t1415 VSS.t1421 315.334
R1483 VSS.t1421 VSS.t1417 315.334
R1484 VSS.t1417 VSS.t1419 315.334
R1485 VSS.t2047 VSS.t2049 315.334
R1486 VSS.t2049 VSS.t2045 315.334
R1487 VSS.t2045 VSS.t2051 315.334
R1488 VSS.t857 VSS.t859 315.334
R1489 VSS.t861 VSS.t857 315.334
R1490 VSS.t863 VSS.t861 315.334
R1491 VSS.t1997 VSS.t2003 315.334
R1492 VSS.t2001 VSS.t1997 315.334
R1493 VSS.t1999 VSS.t2001 315.334
R1494 VSS.t1386 VSS.t1380 315.334
R1495 VSS.t1382 VSS.t1386 315.334
R1496 VSS.t1384 VSS.t1382 315.334
R1497 VSS.n1185 VSS.n1184 315.283
R1498 VSS.t1920 VSS.n1022 314.286
R1499 VSS.n1191 VSS.n1190 312.094
R1500 VSS.n4651 VSS.n1243 312.094
R1501 VSS.t647 VSS.t1938 311.877
R1502 VSS.t570 VSS.t1958 311.877
R1503 VSS.t1480 VSS.t1338 311.877
R1504 VSS.n1195 VSS.n1194 309.702
R1505 VSS.t1758 VSS.t1760 308
R1506 VSS.t1028 VSS.t1030 308
R1507 VSS.t1096 VSS.t1098 308
R1508 VSS.t1172 VSS.t1174 308
R1509 VSS.t478 VSS.t605 308
R1510 VSS.t605 VSS.t111 308
R1511 VSS.t1446 VSS.t1444 308
R1512 VSS.t2853 VSS.t472 308
R1513 VSS.t1613 VSS.t1611 308
R1514 VSS.t2007 VSS.t2005 308
R1515 VSS.t2676 VSS.t2674 308
R1516 VSS.t1237 VSS.t1239 308
R1517 VSS.n3818 VSS.t1281 307.536
R1518 VSS.n4418 VSS.t1304 307.536
R1519 VSS.n3681 VSS.t1988 307.536
R1520 VSS.n3633 VSS.t2681 307.536
R1521 VSS.n3578 VSS.t1258 307.536
R1522 VSS.n3443 VSS.t867 307.536
R1523 VSS.n2446 VSS.t1971 307.536
R1524 VSS.n1984 VSS.t1414 307.536
R1525 VSS.n1967 VSS.t1339 307.536
R1526 VSS.n1934 VSS.t2060 307.536
R1527 VSS.n1883 VSS.t1980 307.536
R1528 VSS.n1829 VSS.t1105 307.536
R1529 VSS.n1454 VSS.t1001 307.536
R1530 VSS.n1466 VSS.t1550 307.536
R1531 VSS.n1728 VSS.t782 307.536
R1532 VSS.n3728 VSS.t1575 307.08
R1533 VSS.n4195 VSS.t1352 306.372
R1534 VSS.n4131 VSS.t1978 304.238
R1535 VSS.n4153 VSS.t1103 304.238
R1536 VSS.n3511 VSS.t1996 304.238
R1537 VSS.n3269 VSS.t1946 304.238
R1538 VSS.n2593 VSS.t886 304.238
R1539 VSS.n2667 VSS.t2024 304.238
R1540 VSS.n2061 VSS.t1891 304.238
R1541 VSS.n1337 VSS.t1517 304.238
R1542 VSS.n1734 VSS.t1184 304.238
R1543 VSS.n1672 VSS.t1283 304.238
R1544 VSS.t617 VSS.t1080 303.449
R1545 VSS.n3737 VSS.t1796 303.449
R1546 VSS.t802 VSS.t1268 303.449
R1547 VSS.t500 VSS.t1038 303.449
R1548 VSS.t317 VSS.t411 303.449
R1549 VSS.t1714 VSS.t2913 303.449
R1550 VSS.n1385 VSS.t2210 303.449
R1551 VSS.t1482 VSS.t2773 303.449
R1552 VSS.t669 VSS.t694 302.264
R1553 VSS.t289 VSS.t1064 302.264
R1554 VSS.t2033 VSS.t2993 302.264
R1555 VSS.t506 VSS.t2809 297.983
R1556 VSS.t537 VSS.t1806 297.127
R1557 VSS.t2170 VSS.t1984 295.019
R1558 VSS.t2118 VSS.t2254 295.019
R1559 VSS.t642 VSS.t1956 295.019
R1560 VSS.t2175 VSS.t1625 295.019
R1561 VSS.t1195 VSS.t1619 295.019
R1562 VSS.t1687 VSS.t1617 295.019
R1563 VSS.n1086 VSS.n1038 292.5
R1564 VSS.t1074 VSS.n1038 292.5
R1565 VSS.n1092 VSS.n1091 292.5
R1566 VSS.n1091 VSS.t1074 292.5
R1567 VSS.n1090 VSS.n1089 292.5
R1568 VSS.t1074 VSS.n1090 292.5
R1569 VSS.n4943 VSS.n365 292.5
R1570 VSS.t2932 VSS.n365 292.5
R1571 VSS.n4962 VSS.n4961 292.5
R1572 VSS.t515 VSS.n4962 292.5
R1573 VSS.n4950 VSS.n4949 292.5
R1574 VSS.n4949 VSS.t64 292.5
R1575 VSS.n4953 VSS.n4952 292.5
R1576 VSS.t2932 VSS.n4953 292.5
R1577 VSS.n4964 VSS.n4963 292.5
R1578 VSS.n4963 VSS.t515 292.5
R1579 VSS.n4966 VSS.n353 292.5
R1580 VSS.n353 VSS.t66 292.5
R1581 VSS.n4606 VSS.t2623 292.252
R1582 VSS.n980 VSS.t2661 292.252
R1583 VSS.n1054 VSS.t3238 291.257
R1584 VSS.n1094 VSS.n1093 290.296
R1585 VSS.n4004 VSS.t1894 290.289
R1586 VSS.n3079 VSS.t1285 290.289
R1587 VSS.n1168 VSS.t2952 289.26
R1588 VSS.n473 VSS.t2946 289.188
R1589 VSS.t1543 VSS.t1541 288.526
R1590 VSS.t2603 VSS.t2605 288.526
R1591 VSS.t2255 VSS.t2257 288.526
R1592 VSS.t2565 VSS.t2563 288.526
R1593 VSS.t2875 VSS.t1745 288.526
R1594 VSS.t649 VSS.t520 288.526
R1595 VSS.t901 VSS.t903 288.526
R1596 VSS.t2870 VSS.t541 288.526
R1597 VSS.n3388 VSS.t1 287.534
R1598 VSS.n3069 VSS.t2715 287.534
R1599 VSS.n3243 VSS.t646 287.534
R1600 VSS.n1823 VSS.t234 287.534
R1601 VSS.t1802 VSS.t1662 286.591
R1602 VSS.t1134 VSS.t1035 286.591
R1603 VSS.t1367 VSS.t2903 286.591
R1604 VSS.t2225 VSS.t1690 286.591
R1605 VSS.t1438 VSS.t48 286.591
R1606 VSS.t2212 VSS.t625 286.591
R1607 VSS.n330 VSS.t1771 286.433
R1608 VSS.n330 VSS.t1780 286.433
R1609 VSS.t2803 VSS.t919 286
R1610 VSS.n337 VSS.t1767 285.481
R1611 VSS.n337 VSS.t1778 285.481
R1612 VSS.n2812 VSS.t98 285.315
R1613 VSS.n2464 VSS.t2863 284.683
R1614 VSS.t693 VSS.t3414 283.93
R1615 VSS.t663 VSS.t448 283.789
R1616 VSS.t667 VSS.t558 283.789
R1617 VSS.n3464 VSS.t2917 283.182
R1618 VSS.n2747 VSS.t2808 283.182
R1619 VSS.n2788 VSS.t404 283.182
R1620 VSS.n4621 VSS.n4620 282.353
R1621 VSS.n4614 VSS.n1256 282.353
R1622 VSS.n1007 VSS.n1006 282.353
R1623 VSS.n996 VSS.n988 282.353
R1624 VSS.n4609 VSS.t2629 282.327
R1625 VSS.n978 VSS.t2663 282.327
R1626 VSS.n1093 VSS.n1032 281.771
R1627 VSS.n1173 VSS.t2940 281.13
R1628 VSS.n4803 VSS.t2950 281.13
R1629 VSS.n4281 VSS.t1799 280.822
R1630 VSS.n2413 VSS.t1862 280.822
R1631 VSS.n2002 VSS.t1626 280.822
R1632 VSS.n1946 VSS.t1477 280.822
R1633 VSS.n1932 VSS.t2207 280.822
R1634 VSS.n1895 VSS.t1715 280.822
R1635 VSS.n1852 VSS.t964 280.822
R1636 VSS.n1796 VSS.t1169 280.822
R1637 VSS.n1773 VSS.t1308 280.822
R1638 VSS.n1484 VSS.t1244 280.822
R1639 VSS.n1687 VSS.t1955 280.822
R1640 VSS.n1637 VSS.t1632 280.822
R1641 VSS.n1022 VSS.n1021 279.366
R1642 VSS.n1194 VSS.n1193 279.012
R1643 VSS.n2501 VSS.t25 278.589
R1644 VSS.t1496 VSS.t343 278.161
R1645 VSS.t2895 VSS.t796 278.161
R1646 VSS.t181 VSS.t185 278.161
R1647 VSS.n1665 VSS.t2896 277.952
R1648 VSS.t1074 VSS.n1036 277.193
R1649 VSS.n3197 VSS.t3621 276.101
R1650 VSS.n964 VSS.t1600 274.812
R1651 VSS.n4348 VSS.t2224 272.728
R1652 VSS.t341 VSS.t1181 269.733
R1653 VSS.t2096 VSS.t2152 269.733
R1654 VSS.t1736 VSS.t1953 269.733
R1655 VSS.t807 VSS.t785 269.733
R1656 VSS.t1439 VSS.t1559 269.733
R1657 VSS.t243 VSS.t1712 269.733
R1658 VSS.n3174 VSS.t3554 269.44
R1659 VSS.t2082 VSS.t2880 266.053
R1660 VSS.t2880 VSS.t298 266.053
R1661 VSS.t298 VSS.t2831 266.053
R1662 VSS.t2831 VSS.t2706 266.053
R1663 VSS.t2706 VSS.t306 266.053
R1664 VSS.t306 VSS.t441 266.053
R1665 VSS.t442 VSS.t443 266.053
R1666 VSS.t443 VSS.t447 266.053
R1667 VSS.t447 VSS.t439 266.053
R1668 VSS.t556 VSS.t562 266.053
R1669 VSS.t561 VSS.t556 266.053
R1670 VSS.t553 VSS.t561 266.053
R1671 VSS.t305 VSS.t557 266.053
R1672 VSS.t22 VSS.t305 266.053
R1673 VSS.t364 VSS.t22 266.053
R1674 VSS.t297 VSS.t364 266.053
R1675 VSS.t126 VSS.t297 266.053
R1676 VSS.t146 VSS.t126 266.053
R1677 VSS.n3893 VSS.t3705 265.473
R1678 VSS.n4467 VSS.t3790 265.298
R1679 VSS.t449 VSS.t2878 264.786
R1680 VSS.t551 VSS.t2825 264.786
R1681 VSS.n1111 VSS.n1110 264.755
R1682 VSS.t2936 VSS.t2835 263.519
R1683 VSS.t456 VSS.t2082 263.519
R1684 VSS.t436 VSS.t442 263.519
R1685 VSS.t439 VSS.t444 263.519
R1686 VSS.t562 VSS.t559 263.519
R1687 VSS.t554 VSS.t553 263.519
R1688 VSS.t457 VSS.t146 263.519
R1689 VSS.t2935 VSS.t2897 263.519
R1690 VSS.n3840 VSS.t3556 262.798
R1691 VSS.n3852 VSS.t3811 262.784
R1692 VSS.n3853 VSS.t3635 262.784
R1693 VSS.n4443 VSS.t3589 262.784
R1694 VSS.n4444 VSS.t3701 262.784
R1695 VSS.n3140 VSS.t3677 262.784
R1696 VSS.n3141 VSS.t3750 262.784
R1697 VSS.n2088 VSS.t3586 262.784
R1698 VSS.n2089 VSS.t3799 262.784
R1699 VSS.n2341 VSS.t3616 262.784
R1700 VSS.n2342 VSS.t3573 262.784
R1701 VSS.n2854 VSS.t3614 262.784
R1702 VSS.n2855 VSS.t3689 262.784
R1703 VSS.n2164 VSS.t3734 262.784
R1704 VSS.n1561 VSS.t3713 262.784
R1705 VSS.n1562 VSS.t3797 262.784
R1706 VSS.n1279 VSS.t3591 262.784
R1707 VSS.n1280 VSS.t3760 262.784
R1708 VSS.n4560 VSS.t3624 262.719
R1709 VSS.n5719 VSS.t3710 262.719
R1710 VSS.n70 VSS.t3793 262.719
R1711 VSS.n5542 VSS.t3687 262.719
R1712 VSS.n149 VSS.t3733 262.719
R1713 VSS.n5410 VSS.t3626 262.719
R1714 VSS.n3832 VSS.t3664 262.719
R1715 VSS.n3911 VSS.t3685 262.719
R1716 VSS.n4334 VSS.t3693 262.719
R1717 VSS.n4429 VSS.t3763 262.719
R1718 VSS.n3165 VSS.t3570 262.719
R1719 VSS.n3182 VSS.t3706 262.719
R1720 VSS.n2075 VSS.t3637 262.719
R1721 VSS.n2574 VSS.t3738 262.719
R1722 VSS.n2525 VSS.t3682 262.719
R1723 VSS.n2306 VSS.t3774 262.719
R1724 VSS.n2316 VSS.t3762 262.719
R1725 VSS.n2401 VSS.t3598 262.719
R1726 VSS.n2175 VSS.t3577 262.719
R1727 VSS.n2160 VSS.t3645 262.719
R1728 VSS.n1608 VSS.t3599 262.719
R1729 VSS.n1310 VSS.t3668 262.719
R1730 VSS.n4983 VSS.n308 262.551
R1731 VSS.t2168 VSS.t329 261.303
R1732 VSS.t335 VSS.t2251 261.303
R1733 VSS.t1734 VSS.t1495 261.303
R1734 VSS.t2587 VSS.t621 261.303
R1735 VSS.n4097 VSS.t2865 259.51
R1736 VSS.n2952 VSS.t170 259.51
R1737 VSS.n3474 VSS.t221 259.51
R1738 VSS.n3410 VSS.t2713 259.51
R1739 VSS.n3346 VSS.t2802 259.51
R1740 VSS.n2219 VSS.t9 259.51
R1741 VSS.n2265 VSS.t683 259.51
R1742 VSS.n2796 VSS.t88 259.51
R1743 VSS.n4511 VSS.t3667 259.082
R1744 VSS.n5740 VSS.t3806 259.082
R1745 VSS.n5588 VSS.t3578 259.082
R1746 VSS.n5365 VSS.t3585 259.082
R1747 VSS.n3865 VSS.t3736 259.082
R1748 VSS.n4300 VSS.t3671 259.082
R1749 VSS.n4328 VSS.t3563 259.082
R1750 VSS.n3588 VSS.t3596 259.082
R1751 VSS.n3405 VSS.t3700 259.082
R1752 VSS.n3222 VSS.t3595 259.082
R1753 VSS.n2487 VSS.t3622 259.082
R1754 VSS.n2778 VSS.t3752 259.082
R1755 VSS.n1991 VSS.t3771 259.082
R1756 VSS.n1892 VSS.t3566 259.082
R1757 VSS.n1698 VSS.t3652 259.082
R1758 VSS.n1631 VSS.t3708 259.082
R1759 VSS.n4823 VSS.t3768 259.082
R1760 VSS.n5033 VSS.t3629 259.082
R1761 VSS.n5041 VSS.t3676 259.082
R1762 VSS.n5277 VSS.t3654 259.082
R1763 VSS.n5291 VSS.t3634 259.082
R1764 VSS.n5332 VSS.t3576 259.082
R1765 VSS.n416 VSS.t3747 259.082
R1766 VSS.n2833 VSS.t410 258.623
R1767 VSS.n4042 VSS.t1045 256.815
R1768 VSS.n2185 VSS.t2919 255.326
R1769 VSS.n1110 VSS.t3396 254.388
R1770 VSS.n1110 VSS.t3251 254.388
R1771 VSS.t64 VSS.n4938 254.28
R1772 VSS.t515 VSS.n358 254.28
R1773 VSS.n2904 VSS.t3751 253.029
R1774 VSS.t2595 VSS.t1275 252.875
R1775 VSS.t191 VSS.t1577 252.875
R1776 VSS.t2996 VSS.t1034 252.875
R1777 VSS.t1472 VSS.t1135 252.875
R1778 VSS.t2271 VSS.t2074 252.875
R1779 VSS.t2757 VSS.t2159 252.875
R1780 VSS.t1024 VSS.t2226 252.875
R1781 VSS.t2662 VSS.n1221 252.423
R1782 VSS.n3375 VSS.t483 251.821
R1783 VSS.t2700 VSS.t123 248.9
R1784 VSS.n4079 VSS.t613 248.069
R1785 VSS.n4948 VSS.n4941 246.233
R1786 VSS.t2691 VSS.t1847 244.893
R1787 VSS.t1658 VSS.t1927 244.445
R1788 VSS.t100 VSS.t395 244.445
R1789 VSS.t1434 VSS.t1183 244.445
R1790 VSS.n4993 VSS.n299 243.306
R1791 VSS.n4508 VSS.t1385 243.286
R1792 VSS.n4546 VSS.t2000 243.286
R1793 VSS.n5765 VSS.t864 243.286
R1794 VSS.n26 VSS.t2048 243.286
R1795 VSS.n42 VSS.t1416 243.286
R1796 VSS.n51 VSS.t1905 243.286
R1797 VSS.n5640 VSS.t1236 243.286
R1798 VSS.n5608 VSS.t1061 243.286
R1799 VSS.n4209 VSS.t1210 243.286
R1800 VSS.n5329 VSS.t2690 243.286
R1801 VSS.n413 VSS.t986 243.286
R1802 VSS.t2632 VSS.t66 243.014
R1803 VSS.n5511 VSS.t2800 242.965
R1804 VSS.n972 VSS.t714 242.945
R1805 VSS.n972 VSS.t799 241.695
R1806 VSS.n5179 VSS.t2698 241.589
R1807 VSS.t2269 VSS.n1066 241.589
R1808 VSS.n1671 VSS.t648 241.054
R1809 VSS.n1618 VSS.t141 240.583
R1810 VSS.n123 VSS.t114 240.575
R1811 VSS.n2434 VSS.t1729 240.575
R1812 VSS.t715 VSS.n5178 239.875
R1813 VSS.n1057 VSS.n1051 239.843
R1814 VSS.t2932 VSS.t2633 239.796
R1815 VSS.n3103 VSS.t1273 239.668
R1816 VSS.n1063 VSS.n1051 239.435
R1817 VSS.n4122 VSS.t2651 239.4
R1818 VSS.n90 VSS.t1445 238.856
R1819 VSS.n144 VSS.t1175 238.856
R1820 VSS.n5423 VSS.t1099 238.856
R1821 VSS.n4120 VSS.t2189 238.856
R1822 VSS.n4374 VSS.t1145 238.856
R1823 VSS.n2447 VSS.t1360 238.856
R1824 VSS.n1844 VSS.t2213 238.856
R1825 VSS.n4065 VSS.t487 238.311
R1826 VSS.n3579 VSS.t499 237.332
R1827 VSS.n3306 VSS.t1749 237.327
R1828 VSS.n3986 VSS.t787 237.226
R1829 VSS.n1068 VSS.t2080 236.633
R1830 VSS.n4970 VSS.n4969 236.577
R1831 VSS.n3456 VSS.t1527 236.554
R1832 VSS.t1840 VSS.t1949 236.016
R1833 VSS.t2888 VSS.t2077 236.016
R1834 VSS.t809 VSS.t2771 236.016
R1835 VSS.t2999 VSS.t2753 236.016
R1836 VSS.t79 VSS.t1931 236.016
R1837 VSS.t1566 VSS.t1307 236.016
R1838 VSS.t794 VSS.n1462 236.016
R1839 VSS.t527 VSS.t965 236.016
R1840 VSS.t2920 VSS.t967 236.016
R1841 VSS.t2231 VSS.t1512 236.016
R1842 VSS.t407 VSS.t856 236.016
R1843 VSS.n4232 VSS.t1252 235.607
R1844 VSS.n3756 VSS.t2145 235.607
R1845 VSS.n3362 VSS.t601 235.014
R1846 VSS.n2979 VSS.t511 234.239
R1847 VSS.n1694 VSS.t643 234.239
R1848 VSS.n4042 VSS.n3985 231.494
R1849 VSS.n3996 VSS.t2078 230.977
R1850 VSS.n4283 VSS.t1663 230.977
R1851 VSS.n3962 VSS.t2894 230.488
R1852 VSS.n2247 VSS.t157 227.68
R1853 VSS.t486 VSS.t610 227.587
R1854 VSS.n4241 VSS.t2769 227.587
R1855 VSS.t2854 VSS.t2137 227.587
R1856 VSS.t866 VSS.t1791 227.587
R1857 VSS.t3151 VSS.t2747 227.587
R1858 VSS.t1637 VSS.t1405 227.587
R1859 VSS.t640 VSS.t1131 227.587
R1860 VSS.t1671 VSS.t1478 227.587
R1861 VSS.n4161 VSS.t2018 226.882
R1862 VSS.n3706 VSS.t1128 226.882
R1863 VSS.n2944 VSS.t1685 226.882
R1864 VSS.n2989 VSS.t1342 226.882
R1865 VSS.n2991 VSS.t999 226.882
R1866 VSS.n3244 VSS.t705 226.882
R1867 VSS.n2201 VSS.t1289 226.882
R1868 VSS.n2649 VSS.t2228 226.882
R1869 VSS.n2021 VSS.t817 226.882
R1870 VSS.n3417 VSS.t1077 226.216
R1871 VSS.n3836 VSS.t3052 223.662
R1872 VSS.n2310 VSS.t3110 223.662
R1873 VSS.n2172 VSS.t3413 223.504
R1874 VSS.n3894 VSS.t3123 223.438
R1875 VSS.n2408 VSS.t3237 223.438
R1876 VSS.n3978 VSS.t879 223.315
R1877 VSS.n4123 VSS.t923 223.315
R1878 VSS.n4222 VSS.t1402 223.315
R1879 VSS.n3601 VSS.t1461 223.315
R1880 VSS.n1705 VSS.t1563 223.315
R1881 VSS.n1538 VSS.t3528 222.784
R1882 VSS.n2628 VSS.t3653 221.958
R1883 VSS.t1323 VSS.n4936 221.903
R1884 VSS.t926 VSS.t924 221.327
R1885 VSS.n2070 VSS.t3594 220.952
R1886 VSS.n2232 VSS.t3688 220.952
R1887 VSS.n3917 VSS.t3425 220.02
R1888 VSS.n3109 VSS.t3199 219.972
R1889 VSS.n2775 VSS.t3215 219.31
R1890 VSS.t1044 VSS.t577 219.157
R1891 VSS.t2026 VSS.t345 219.157
R1892 VSS.t1551 VSS.t851 219.157
R1893 VSS.t2755 VSS.t2116 219.157
R1894 VSS.t2588 VSS.n2954 219.157
R1895 VSS.t2241 VSS.t2618 219.157
R1896 VSS.t1823 VSS.t1226 219.157
R1897 VSS.t2261 VSS.t939 219.157
R1898 VSS.n3111 VSS.t3561 218.607
R1899 VSS.n3106 VSS.t3795 218.607
R1900 VSS.n3288 VSS.t3246 218.428
R1901 VSS.n5617 VSS.t3813 218.308
R1902 VSS.n5561 VSS.t3683 218.308
R1903 VSS.n5526 VSS.t3552 218.308
R1904 VSS.n5432 VSS.t3695 218.308
R1905 VSS.n4108 VSS.t3711 218.308
R1906 VSS.n4224 VSS.t3753 218.308
R1907 VSS.n4314 VSS.t3553 218.308
R1908 VSS.n4484 VSS.t3786 218.308
R1909 VSS.n3471 VSS.t3632 218.308
R1910 VSS.n3454 VSS.t3673 218.308
R1911 VSS.n3394 VSS.t3780 218.308
R1912 VSS.n2608 VSS.t3661 218.308
R1913 VSS.n2459 VSS.t3729 218.308
R1914 VSS.n2716 VSS.t3767 218.308
R1915 VSS.n2675 VSS.t3814 218.308
R1916 VSS.n2748 VSS.t3686 218.308
R1917 VSS.n2062 VSS.t3660 218.308
R1918 VSS.n4873 VSS.t3571 218.308
R1919 VSS.n238 VSS.t3666 218.308
R1920 VSS.n230 VSS.t3684 218.308
R1921 VSS.n222 VSS.t3704 218.308
R1922 VSS.n214 VSS.t3551 218.308
R1923 VSS.n5237 VSS.t3584 218.308
R1924 VSS.n455 VSS.t3725 218.308
R1925 VSS.n2908 VSS.t3141 217.953
R1926 VSS.n2629 VSS.t3065 217.934
R1927 VSS.t1296 VSS.t2416 217.285
R1928 VSS.t2489 VSS.t1294 217.285
R1929 VSS.n2122 VSS.t3049 216.959
R1930 VSS.n1326 VSS.t3104 216.933
R1931 VSS.n1189 VSS.n1013 216.847
R1932 VSS.n4652 VSS.n1242 216.847
R1933 VSS.n2121 VSS.t3471 216.632
R1934 VSS.n2387 VSS.t3092 216.632
R1935 VSS.n3882 VSS.t3122 216.579
R1936 VSS.n2838 VSS.t3507 215.407
R1937 VSS.n2631 VSS.t3137 215.407
R1938 VSS.n1191 VSS.n1012 214.589
R1939 VSS.n1114 VSS.n1013 214.589
R1940 VSS.n4642 VSS.n1242 214.589
R1941 VSS.n4644 VSS.n1243 214.589
R1942 VSS.n4558 VSS.t3171 214.456
R1943 VSS.n4564 VSS.t3170 214.456
R1944 VSS.n4510 VSS.t3457 214.456
R1945 VSS.n4513 VSS.t3456 214.456
R1946 VSS.n5726 VSS.t3460 214.456
R1947 VSS.n32 VSS.t3459 214.456
R1948 VSS.n20 VSS.t3081 214.456
R1949 VSS.n5739 VSS.t3080 214.456
R1950 VSS.n17 VSS.t3134 214.456
R1951 VSS.n16 VSS.t3135 214.456
R1952 VSS.n5700 VSS.t3185 214.456
R1953 VSS.n34 VSS.t3186 214.456
R1954 VSS.n5589 VSS.t3422 214.456
R1955 VSS.n5586 VSS.t3421 214.456
R1956 VSS.n5618 VSS.t3084 214.456
R1957 VSS.n5611 VSS.t3083 214.456
R1958 VSS.n68 VSS.t3484 214.456
R1959 VSS.n74 VSS.t3483 214.456
R1960 VSS.n5655 VSS.t3161 214.456
R1961 VSS.n5669 VSS.t3162 214.456
R1962 VSS.n45 VSS.t3095 214.456
R1963 VSS.n44 VSS.t3096 214.456
R1964 VSS.n5471 VSS.t3542 214.456
R1965 VSS.n5486 VSS.t3543 214.456
R1966 VSS.n5527 VSS.t3174 214.456
R1967 VSS.n5520 VSS.t3173 214.456
R1968 VSS.n5548 VSS.t3038 214.456
R1969 VSS.n5529 VSS.t3037 214.456
R1970 VSS.n5562 VSS.t3468 214.456
R1971 VSS.n101 VSS.t3467 214.456
R1972 VSS.n5568 VSS.t3116 214.456
R1973 VSS.n96 VSS.t3117 214.456
R1974 VSS.n5416 VSS.t3057 214.456
R1975 VSS.n5397 VSS.t3056 214.456
R1976 VSS.n5433 VSS.t3120 214.456
R1977 VSS.n5426 VSS.t3119 214.456
R1978 VSS.n5451 VSS.t3144 214.456
R1979 VSS.n153 VSS.t3143 214.456
R1980 VSS.n5463 VSS.t3530 214.456
R1981 VSS.n141 VSS.t3531 214.456
R1982 VSS.n5363 VSS.t3499 214.456
R1983 VSS.n5364 VSS.t3498 214.456
R1984 VSS.n3867 VSS.t3069 214.456
R1985 VSS.n3846 VSS.t3068 214.456
R1986 VSS.n3852 VSS.t3044 214.456
R1987 VSS.n3852 VSS.t3043 214.456
R1988 VSS.n3853 VSS.t3445 214.456
R1989 VSS.n3853 VSS.t3444 214.456
R1990 VSS.n4431 VSS.t3401 214.456
R1991 VSS.n4428 VSS.t3077 214.456
R1992 VSS.n4425 VSS.t3400 214.456
R1993 VSS.n4483 VSS.t3212 214.456
R1994 VSS.n4425 VSS.t3211 214.456
R1995 VSS.n4340 VSS.t3072 214.456
R1996 VSS.n3723 VSS.t3189 214.456
R1997 VSS.n4327 VSS.t3188 214.456
R1998 VSS.n4320 VSS.t3071 214.456
R1999 VSS.n4315 VSS.t3404 214.456
R2000 VSS.n3730 VSS.t3403 214.456
R2001 VSS.n4301 VSS.t3537 214.456
R2002 VSS.n3735 VSS.t3536 214.456
R2003 VSS.n3750 VSS.t3407 214.456
R2004 VSS.n4256 VSS.t3406 214.456
R2005 VSS.n4223 VSS.t3463 214.456
R2006 VSS.n4173 VSS.t3462 214.456
R2007 VSS.n3781 VSS.t3102 214.456
R2008 VSS.n4105 VSS.t3101 214.456
R2009 VSS.n4087 VSS.t3487 214.456
R2010 VSS.n4072 VSS.t3486 214.456
R2011 VSS.n3983 VSS.t3026 214.456
R2012 VSS.n3977 VSS.t3025 214.456
R2013 VSS.n3940 VSS.t3041 214.456
R2014 VSS.n3922 VSS.t3040 214.456
R2015 VSS.n3830 VSS.t3053 214.456
R2016 VSS.n3899 VSS.t3424 214.456
R2017 VSS.n3890 VSS.t3448 214.456
R2018 VSS.n3884 VSS.t3447 214.456
R2019 VSS.n3840 VSS.t3502 214.456
R2020 VSS.n3840 VSS.t3501 214.456
R2021 VSS.n4461 VSS.t3078 214.456
R2022 VSS.n4443 VSS.t3087 214.456
R2023 VSS.n4443 VSS.t3086 214.456
R2024 VSS.n4444 VSS.t3197 214.456
R2025 VSS.n4444 VSS.t3196 214.456
R2026 VSS.n3113 VSS.t3182 214.456
R2027 VSS.n3110 VSS.t3183 214.456
R2028 VSS.n3105 VSS.t3200 214.456
R2029 VSS.n3304 VSS.t3247 214.456
R2030 VSS.n3350 VSS.t3418 214.456
R2031 VSS.n3076 VSS.t3419 214.456
R2032 VSS.n3395 VSS.t3029 214.456
R2033 VSS.n3062 VSS.t3028 214.456
R2034 VSS.n3055 VSS.t3438 214.456
R2035 VSS.n3404 VSS.t3437 214.456
R2036 VSS.n3455 VSS.t3192 214.456
R2037 VSS.n3034 VSS.t3191 214.456
R2038 VSS.n3472 VSS.t3126 214.456
R2039 VSS.n3465 VSS.t3125 214.456
R2040 VSS.n3589 VSS.t3153 214.456
R2041 VSS.n3583 VSS.t3152 214.456
R2042 VSS.n3592 VSS.t3046 214.456
R2043 VSS.n3612 VSS.t3047 214.456
R2044 VSS.n3221 VSS.t3435 214.456
R2045 VSS.n3157 VSS.t3434 214.456
R2046 VSS.n3161 VSS.t3480 214.456
R2047 VSS.n3167 VSS.t3481 214.456
R2048 VSS.n3164 VSS.t3450 214.456
R2049 VSS.n3195 VSS.t3533 214.456
R2050 VSS.n3171 VSS.t3451 214.456
R2051 VSS.n3176 VSS.t3534 214.456
R2052 VSS.n3188 VSS.t3107 214.456
R2053 VSS.n3236 VSS.t3510 214.456
R2054 VSS.n3238 VSS.t3108 214.456
R2055 VSS.n3127 VSS.t3511 214.456
R2056 VSS.n3140 VSS.t3430 214.456
R2057 VSS.n3140 VSS.t3429 214.456
R2058 VSS.n3141 VSS.t3060 214.456
R2059 VSS.n3141 VSS.t3059 214.456
R2060 VSS.n2088 VSS.t3203 214.456
R2061 VSS.n2088 VSS.t3202 214.456
R2062 VSS.n2089 VSS.t3398 214.456
R2063 VSS.n2089 VSS.t3397 214.456
R2064 VSS.n2078 VSS.t3472 214.456
R2065 VSS.n2124 VSS.t3050 214.456
R2066 VSS.n2070 VSS.t3075 214.456
R2067 VSS.n2070 VSS.t3074 214.456
R2068 VSS.n2583 VSS.t3525 214.456
R2069 VSS.n2226 VSS.t3524 214.456
R2070 VSS.n2607 VSS.t3454 214.456
R2071 VSS.n2604 VSS.t3453 214.456
R2072 VSS.n2324 VSS.t3249 214.456
R2073 VSS.n2320 VSS.t3250 214.456
R2074 VSS.n2322 VSS.t3022 214.456
R2075 VSS.n2385 VSS.t3023 214.456
R2076 VSS.n2400 VSS.t3093 214.456
R2077 VSS.n2388 VSS.t3236 214.456
R2078 VSS.n2303 VSS.t3111 214.456
R2079 VSS.n2284 VSS.t3129 214.456
R2080 VSS.n2456 VSS.t3128 214.456
R2081 VSS.n2270 VSS.t3475 214.456
R2082 VSS.n2486 VSS.t3474 214.456
R2083 VSS.n2531 VSS.t3478 214.456
R2084 VSS.n2511 VSS.t3477 214.456
R2085 VSS.n2230 VSS.t3233 214.456
R2086 VSS.n2232 VSS.t3441 214.456
R2087 VSS.n2232 VSS.t3440 214.456
R2088 VSS.n2228 VSS.t3234 214.456
R2089 VSS.n2341 VSS.t3465 214.456
R2090 VSS.n2341 VSS.t3464 214.456
R2091 VSS.n2342 VSS.t3147 214.456
R2092 VSS.n2342 VSS.t3146 214.456
R2093 VSS.n2164 VSS.t3063 214.456
R2094 VSS.n2164 VSS.t3062 214.456
R2095 VSS.n2897 VSS.t3539 214.456
R2096 VSS.n2891 VSS.t3508 214.456
R2097 VSS.n2846 VSS.t3540 214.456
R2098 VSS.n2854 VSS.t3035 214.456
R2099 VSS.n2854 VSS.t3034 214.456
R2100 VSS.n2855 VSS.t3432 214.456
R2101 VSS.n2855 VSS.t3431 214.456
R2102 VSS.n2905 VSS.t3208 214.456
R2103 VSS.n2155 VSS.t3140 214.456
R2104 VSS.n2779 VSS.t3216 214.456
R2105 VSS.n2180 VSS.t3412 214.456
R2106 VSS.n2749 VSS.t3505 214.456
R2107 VSS.n2741 VSS.t3504 214.456
R2108 VSS.n2677 VSS.t3020 214.456
R2109 VSS.n2706 VSS.t3019 214.456
R2110 VSS.n2715 VSS.t3516 214.456
R2111 VSS.n2665 VSS.t3515 214.456
R2112 VSS.n2195 VSS.t3138 214.456
R2113 VSS.n2628 VSS.t3066 214.456
R2114 VSS.n2903 VSS.t3209 214.456
R2115 VSS.n1893 VSS.t3195 214.456
R2116 VSS.n1409 VSS.t3194 214.456
R2117 VSS.n1909 VSS.t3492 214.456
R2118 VSS.n1395 VSS.t3493 214.456
R2119 VSS.n1992 VSS.t3490 214.456
R2120 VSS.n1989 VSS.t3489 214.456
R2121 VSS.n1332 VSS.t3428 214.456
R2122 VSS.n2059 VSS.t3427 214.456
R2123 VSS.n1630 VSS.t3159 214.456
R2124 VSS.n1629 VSS.t3158 214.456
R2125 VSS.n1511 VSS.t3225 214.456
R2126 VSS.n1673 VSS.t3224 214.456
R2127 VSS.n1503 VSS.t3168 214.456
R2128 VSS.n1696 VSS.t3167 214.456
R2129 VSS.n1864 VSS.t3230 214.456
R2130 VSS.n1423 VSS.t3231 214.456
R2131 VSS.n1593 VSS.t3527 214.456
R2132 VSS.n1607 VSS.t3545 214.456
R2133 VSS.n1617 VSS.t3546 214.456
R2134 VSS.n1561 VSS.t3443 214.456
R2135 VSS.n1561 VSS.t3442 214.456
R2136 VSS.n1562 VSS.t3114 214.456
R2137 VSS.n1562 VSS.t3113 214.456
R2138 VSS.n1279 VSS.t3180 214.456
R2139 VSS.n1279 VSS.t3179 214.456
R2140 VSS.n1280 VSS.t3513 214.456
R2141 VSS.n1280 VSS.t3512 214.456
R2142 VSS.n1303 VSS.t3496 214.456
R2143 VSS.n1324 VSS.t3495 214.456
R2144 VSS.n1318 VSS.t3105 214.456
R2145 VSS.n4872 VSS.t3017 214.456
R2146 VSS.n372 VSS.t3016 214.456
R2147 VSS.n4822 VSS.t3156 214.456
R2148 VSS.n390 VSS.t3155 214.456
R2149 VSS.n5010 VSS.t3239 214.456
R2150 VSS.n289 VSS.t3240 214.456
R2151 VSS.n5040 VSS.t3090 214.456
R2152 VSS.n272 VSS.t3089 214.456
R2153 VSS.n5032 VSS.t3032 214.456
R2154 VSS.n276 VSS.t3031 214.456
R2155 VSS.n5024 VSS.t3415 214.456
R2156 VSS.n281 VSS.t3416 214.456
R2157 VSS.n266 VSS.t3131 214.456
R2158 VSS.n267 VSS.t3132 214.456
R2159 VSS.n240 VSS.t3177 214.456
R2160 VSS.n5118 VSS.t3176 214.456
R2161 VSS.n5069 VSS.t3149 214.456
R2162 VSS.n260 VSS.t3150 214.456
R2163 VSS.n5133 VSS.t3521 214.456
R2164 VSS.n5132 VSS.t3522 214.456
R2165 VSS.n5334 VSS.t3519 214.456
R2166 VSS.n5331 VSS.t3518 214.456
R2167 VSS.n5290 VSS.t3222 214.456
R2168 VSS.n5293 VSS.t3221 214.456
R2169 VSS.n5276 VSS.t3410 214.456
R2170 VSS.n194 VSS.t3409 214.456
R2171 VSS.n5236 VSS.t3228 214.456
R2172 VSS.n208 VSS.t3227 214.456
R2173 VSS.n216 VSS.t3549 214.456
R2174 VSS.n5223 VSS.t3548 214.456
R2175 VSS.n224 VSS.t3165 214.456
R2176 VSS.n5205 VSS.t3164 214.456
R2177 VSS.n231 VSS.t3206 214.456
R2178 VSS.n5192 VSS.t3205 214.456
R2179 VSS.n5142 VSS.t3218 214.456
R2180 VSS.n5144 VSS.t3219 214.456
R2181 VSS.n415 VSS.t3099 214.456
R2182 VSS.n418 VSS.t3098 214.456
R2183 VSS.n454 VSS.t3243 214.456
R2184 VSS.n395 VSS.t3242 214.456
R2185 VSS.t3088 VSS.t1923 213.406
R2186 VSS.t2881 VSS.t3030 212.49
R2187 VSS.t560 VSS.n461 211.828
R2188 VSS.t2737 VSS.n1259 211.828
R2189 VSS.t2735 VSS.n461 211.828
R2190 VSS.n1259 VSS.t549 211.828
R2191 VSS.n2552 VSS.n2235 211.109
R2192 VSS.n1644 VSS.n1643 211.062
R2193 VSS.t710 VSS.t484 210.728
R2194 VSS.t2612 VSS.t2712 210.728
R2195 VSS.t169 VSS.t2680 210.728
R2196 VSS.n2692 VSS.n2682 210.51
R2197 VSS.n1757 VSS.n1483 210.099
R2198 VSS.t1499 VSS.t70 209.909
R2199 VSS.n1098 VSS.t2822 209.686
R2200 VSS.n3970 VSS.n3969 209.254
R2201 VSS.n4390 VSS.n4388 209.254
R2202 VSS.n3648 VSS.n2942 209.254
R2203 VSS.n3556 VSS.n2987 209.254
R2204 VSS.n2995 VSS.n2994 209.254
R2205 VSS.n3250 VSS.n3124 209.254
R2206 VSS.n2205 VSS.n2204 209.254
R2207 VSS.n2033 VSS.n2032 209.254
R2208 VSS.n1350 VSS.n1349 209.254
R2209 VSS.n1961 VSS.n1960 209.254
R2210 VSS.n1712 VSS.n1499 209.254
R2211 VSS.n1524 VSS.n1523 209.254
R2212 VSS.n3928 VSS.n3825 208.719
R2213 VSS.n3931 VSS.n3930 208.719
R2214 VSS.n3789 VSS.n3788 208.719
R2215 VSS.n4099 VSS.n3787 208.719
R2216 VSS.n3487 VSS.n3016 208.719
R2217 VSS.n3018 VSS.n3017 208.719
R2218 VSS.n2619 VSS.n2203 208.719
R2219 VSS.n2622 VSS.n2621 208.719
R2220 VSS.n2585 VSS.n2584 208.719
R2221 VSS.n2581 VSS.n2221 208.719
R2222 VSS.n2550 VSS.n2236 208.719
R2223 VSS.n2471 VSS.n2280 208.719
R2224 VSS.n2278 VSS.n2277 208.719
R2225 VSS.n2699 VSS.n2678 208.719
R2226 VSS.n2704 VSS.n2674 208.719
R2227 VSS.n2770 VSS.n2174 208.719
R2228 VSS.n2764 VSS.n2763 208.719
R2229 VSS.n2014 VSS.n1352 208.719
R2230 VSS.n2009 VSS.n1355 208.719
R2231 VSS.n4858 VSS.n377 208.719
R2232 VSS.n4837 VSS.n4836 208.719
R2233 VSS.n4064 VSS.n4063 208.553
R2234 VSS.n3743 VSS.n3742 207.965
R2235 VSS.n4354 VSS.n3714 207.965
R2236 VSS.n4366 VSS.n3711 207.965
R2237 VSS.n2416 VSS.n2415 207.965
R2238 VSS.n2007 VSS.n1356 207.965
R2239 VSS.n1952 VSS.n1382 207.965
R2240 VSS.n1391 VSS.n1390 207.965
R2241 VSS.n1901 VSS.n1406 207.965
R2242 VSS.n1857 VSS.n1429 207.965
R2243 VSS.n1457 VSS.n1456 207.965
R2244 VSS.n1778 VSS.n1470 207.965
R2245 VSS.n1693 VSS.n1506 207.965
R2246 VSS.n982 VSS.n981 207.213
R2247 VSS.n1169 VSS.n1167 207.213
R2248 VSS.n335 VSS.n327 207.213
R2249 VSS.n335 VSS.n328 207.213
R2250 VSS.n4008 VSS.n4003 207.213
R2251 VSS.n4070 VSS.n3801 207.213
R2252 VSS.n3368 VSS.n3072 207.213
R2253 VSS.n2697 VSS.n2679 207.213
R2254 VSS.n474 VSS.n472 207.213
R2255 VSS.n4604 VSS.n4603 207.213
R2256 VSS.n1466 VSS.n1465 206.823
R2257 VSS.n345 VSS.n344 206.333
R2258 VSS.n3423 VSS.n3045 205.661
R2259 VSS.n1109 VSS.t245 205.24
R2260 VSS.n4520 VSS.n4519 205.078
R2261 VSS.n4551 VSS.n4550 205.078
R2262 VSS.n5763 VSS.n10 205.078
R2263 VSS.n5732 VSS.n25 205.078
R2264 VSS.n5693 VSS.n41 205.078
R2265 VSS.n5675 VSS.n50 205.078
R2266 VSS.n66 VSS.n65 205.078
R2267 VSS.n82 VSS.n81 205.078
R2268 VSS.n1619 VSS.n1535 205.078
R2269 VSS.n5340 VSS.n5327 205.078
R2270 VSS.n424 VSS.n412 205.078
R2271 VSS.n5596 VSS.n87 204.457
R2272 VSS.n4202 VSS.n4184 204.457
R2273 VSS.n4411 VSS.n4410 204.457
R2274 VSS.n3682 VSS.n2133 204.457
R2275 VSS.n3674 VSS.n2137 204.457
R2276 VSS.n3517 VSS.n3002 204.457
R2277 VSS.n3437 VSS.n3436 204.457
R2278 VSS.n2478 VSS.n2276 204.457
R2279 VSS.n1998 VSS.n1363 204.457
R2280 VSS.n1837 VSS.n1836 204.457
R2281 VSS.n5256 VSS.n5255 204.457
R2282 VSS.n4120 VSS.n3778 204.06
R2283 VSS.n4506 VSS.n4505 203.619
R2284 VSS.n4554 VSS.n4553 203.619
R2285 VSS.n12 VSS.n11 203.619
R2286 VSS.n23 VSS.n22 203.619
R2287 VSS.n39 VSS.n38 203.619
R2288 VSS.n48 VSS.n47 203.619
R2289 VSS.n5646 VSS.n64 203.619
R2290 VSS.n5602 VSS.n84 203.619
R2291 VSS.n5580 VSS.n92 203.619
R2292 VSS.n5457 VSS.n146 203.619
R2293 VSS.n161 VSS.n160 203.619
R2294 VSS.n4116 VSS.n4114 203.619
R2295 VSS.n4116 VSS.n4115 203.619
R2296 VSS.n4168 VSS.n4167 203.619
R2297 VSS.n4217 VSS.n4176 203.619
R2298 VSS.n4250 VSS.n4249 203.619
R2299 VSS.n2445 VSS.n2295 203.619
R2300 VSS.n1434 VSS.n1433 203.619
R2301 VSS.n1621 VSS.n1534 203.619
R2302 VSS.n5342 VSS.n5326 203.619
R2303 VSS.n410 VSS.n409 203.619
R2304 VSS.n4130 VSS.n3773 203.526
R2305 VSS.n4155 VSS.n3766 203.526
R2306 VSS.n4215 VSS.n4177 203.526
R2307 VSS.n4294 VSS.n3738 203.526
R2308 VSS.n3611 VSS.n2961 203.526
R2309 VSS.n2428 VSS.n2305 203.526
R2310 VSS.n2655 VSS.n2187 203.526
R2311 VSS.n1944 VSS.n1386 203.526
R2312 VSS.n1911 VSS.n1402 203.526
R2313 VSS.n1425 VSS.n1424 203.526
R2314 VSS.n1809 VSS.n1453 203.526
R2315 VSS.n1766 VSS.n1478 203.526
R2316 VSS.n1704 VSS.n1502 203.526
R2317 VSS.n1003 VSS.n997 203.294
R2318 VSS.n4615 VSS.n1255 203.294
R2319 VSS.n1252 VSS.n1251 203.294
R2320 VSS.n1207 VSS.n1206 203.294
R2321 VSS.n3339 VSS.n3085 203.214
R2322 VSS.n4372 VSS.n3709 202.959
R2323 VSS.n2479 VSS.n2275 202.349
R2324 VSS.t40 VSS.t1952 202.299
R2325 VSS.t755 VSS.t34 202.299
R2326 VSS.t3402 VSS.t1680 202.299
R2327 VSS.t995 VSS.t2063 202.299
R2328 VSS.t1107 VSS.t1970 202.299
R2329 VSS.t261 VSS.t275 202.299
R2330 VSS.t1817 VSS.t512 202.299
R2331 VSS.t2743 VSS.t2027 202.299
R2332 VSS.t2021 VSS.t1718 202.299
R2333 VSS.t405 VSS.t466 202.299
R2334 VSS.n3083 VSS.n3082 202.067
R2335 VSS.n1199 VSS.n1003 201.036
R2336 VSS.n1255 VSS.n466 201.036
R2337 VSS.n4645 VSS.n4621 201.036
R2338 VSS.n4595 VSS.n1256 201.036
R2339 VSS.n1252 VSS.n465 201.036
R2340 VSS.n1207 VSS.n989 201.036
R2341 VSS.n1006 VSS.n1004 201.036
R2342 VSS.n1213 VSS.n988 201.036
R2343 VSS.n4214 VSS.n4178 200.812
R2344 VSS.n5668 VSS.n5667 200.692
R2345 VSS.n5485 VSS.n5484 200.692
R2346 VSS.n4086 VSS.n4085 200.692
R2347 VSS.n3939 VSS.n3938 200.692
R2348 VSS.n3303 VSS.n3302 200.692
R2349 VSS.n3361 VSS.n3360 200.692
R2350 VSS.n3610 VSS.n3609 200.692
R2351 VSS.n2887 VSS.n2842 200.692
R2352 VSS.n2641 VSS.n2640 200.692
R2353 VSS.n1921 VSS.n1920 200.692
R2354 VSS.n342 VSS.n341 200.516
R2355 VSS.n120 VSS.n119 200.516
R2356 VSS.n4036 VSS.n3989 200.516
R2357 VSS.n4092 VSS.n3793 200.516
R2358 VSS.n3785 VSS.n3784 200.516
R2359 VSS.n3740 VSS.n3739 200.516
R2360 VSS.n3634 VSS.n2950 200.516
R2361 VSS.n3480 VSS.n3022 200.516
R2362 VSS.n3479 VSS.n3023 200.516
R2363 VSS.n3051 VSS.n3050 200.516
R2364 VSS.n2614 VSS.n2207 200.516
R2365 VSS.n2592 VSS.n2216 200.516
R2366 VSS.n2545 VSS.n2239 200.516
R2367 VSS.n2500 VSS.n2262 200.516
R2368 VSS.n2466 VSS.n2283 200.516
R2369 VSS.n2189 VSS.n2188 200.516
R2370 VSS.n2671 VSS.n2670 200.516
R2371 VSS.n2833 VSS.n2800 200.516
R2372 VSS.n2828 VSS.n2805 200.516
R2373 VSS.n4847 VSS.n4835 200.516
R2374 VSS.n126 VSS.n125 200.231
R2375 VSS.n3092 VSS.n3091 200.231
R2376 VSS.n2440 VSS.n2299 200.231
R2377 VSS.n2499 VSS.n2263 200.127
R2378 VSS.n1746 VSS.n1743 200.105
R2379 VSS.n1627 VSS.n1626 199.921
R2380 VSS.n4503 VSS.n4502 199.739
R2381 VSS.n4500 VSS.n4499 199.739
R2382 VSS.n4540 VSS.n4539 199.739
R2383 VSS.n5575 VSS.n95 199.739
R2384 VSS.n104 VSS.n103 199.739
R2385 VSS.n5518 VSS.n115 199.739
R2386 VSS.n129 VSS.n128 199.739
R2387 VSS.n5395 VSS.n170 199.739
R2388 VSS.n5389 VSS.n173 199.739
R2389 VSS.n5384 VSS.n176 199.739
R2390 VSS.n5377 VSS.n5358 199.739
R2391 VSS.n5372 VSS.n5361 199.739
R2392 VSS.n3858 VSS.n3848 199.739
R2393 VSS.n3858 VSS.n3850 199.739
R2394 VSS.n3877 VSS.n3875 199.739
R2395 VSS.n3877 VSS.n3876 199.739
R2396 VSS.n3967 VSS.n3813 199.739
R2397 VSS.n3792 VSS.n3791 199.739
R2398 VSS.n4128 VSS.n3775 199.739
R2399 VSS.n4139 VSS.n4138 199.739
R2400 VSS.n4146 VSS.n4145 199.739
R2401 VSS.n3764 VSS.n3763 199.739
R2402 VSS.n4163 VSS.n4162 199.739
R2403 VSS.n4182 VSS.n4181 199.739
R2404 VSS.n4190 VSS.n4189 199.739
R2405 VSS.n4244 VSS.n4243 199.739
R2406 VSS.n4347 VSS.n4346 199.739
R2407 VSS.n4372 VSS.n4371 199.739
R2408 VSS.n4404 VSS.n4403 199.739
R2409 VSS.n3696 VSS.n3695 199.739
R2410 VSS.n4491 VSS.n4422 199.739
R2411 VSS.n4442 VSS.n4440 199.739
R2412 VSS.n4442 VSS.n4441 199.739
R2413 VSS.n4438 VSS.n4436 199.739
R2414 VSS.n4438 VSS.n4437 199.739
R2415 VSS.n3684 VSS.n2132 199.739
R2416 VSS.n3668 VSS.n3667 199.739
R2417 VSS.n3666 VSS.n2141 199.739
R2418 VSS.n3635 VSS.n2947 199.739
R2419 VSS.n3622 VSS.n2958 199.739
R2420 VSS.n3580 VSS.n2974 199.739
R2421 VSS.n3562 VSS.n2983 199.739
R2422 VSS.n3538 VSS.n2993 199.739
R2423 VSS.n3524 VSS.n2999 199.739
R2424 VSS.n3503 VSS.n3010 199.739
R2425 VSS.n3412 VSS.n3053 199.739
R2426 VSS.n3135 VSS.n3134 199.739
R2427 VSS.n3139 VSS.n3137 199.739
R2428 VSS.n3139 VSS.n3138 199.739
R2429 VSS.n2095 VSS.n2086 199.739
R2430 VSS.n2095 VSS.n2094 199.739
R2431 VSS.n2101 VSS.n2082 199.739
R2432 VSS.n2101 VSS.n2083 199.739
R2433 VSS.n2591 VSS.n2218 199.739
R2434 VSS.n2494 VSS.n2267 199.739
R2435 VSS.n2448 VSS.n2292 199.739
R2436 VSS.n2301 VSS.n2300 199.739
R2437 VSS.n2362 VSS.n2330 199.739
R2438 VSS.n2354 VSS.n2333 199.739
R2439 VSS.n2347 VSS.n2337 199.739
R2440 VSS.n2347 VSS.n2339 199.739
R2441 VSS.n2862 VSS.n2860 199.739
R2442 VSS.n2862 VSS.n2861 199.739
R2443 VSS.n2870 VSS.n2868 199.739
R2444 VSS.n2870 VSS.n2869 199.739
R2445 VSS.n2729 VSS.n2662 199.739
R2446 VSS.n2067 VSS.n1331 199.739
R2447 VSS.n2054 VSS.n1336 199.739
R2448 VSS.n2030 VSS.n1346 199.739
R2449 VSS.n1954 VSS.n1381 199.739
R2450 VSS.n1938 VSS.n1389 199.739
R2451 VSS.n1885 VSS.n1412 199.739
R2452 VSS.n1442 VSS.n1441 199.739
R2453 VSS.n1790 VSS.n1464 199.739
R2454 VSS.n1472 VSS.n1471 199.739
R2455 VSS.n1490 VSS.n1489 199.739
R2456 VSS.n1493 VSS.n1492 199.739
R2457 VSS.n1722 VSS.n1721 199.739
R2458 VSS.n1714 VSS.n1713 199.739
R2459 VSS.n1517 VSS.n1516 199.739
R2460 VSS.n1587 VSS.n1548 199.739
R2461 VSS.n1582 VSS.n1551 199.739
R2462 VSS.n1574 VSS.n1554 199.739
R2463 VSS.n1567 VSS.n1557 199.739
R2464 VSS.n1567 VSS.n1559 199.739
R2465 VSS.n1278 VSS.n1276 199.739
R2466 VSS.n1278 VSS.n1277 199.739
R2467 VSS.n1274 VSS.n1272 199.739
R2468 VSS.n1274 VSS.n1273 199.739
R2469 VSS.n1270 VSS.n1269 199.739
R2470 VSS.n393 VSS.n392 199.739
R2471 VSS.n388 VSS.n387 199.739
R2472 VSS.n4867 VSS.n4866 199.739
R2473 VSS.n4880 VSS.n4879 199.739
R2474 VSS.n4904 VSS.n4893 199.739
R2475 VSS.n4896 VSS.n4895 199.739
R2476 VSS.n5003 VSS.n5002 199.739
R2477 VSS.n5016 VSS.n286 199.739
R2478 VSS.n278 VSS.n277 199.739
R2479 VSS.n5049 VSS.n5048 199.739
R2480 VSS.n5062 VSS.n5061 199.739
R2481 VSS.n5075 VSS.n257 199.739
R2482 VSS.n5105 VSS.n245 199.739
R2483 VSS.n5111 VSS.n242 199.739
R2484 VSS.n5124 VSS.n5123 199.739
R2485 VSS.n5164 VSS.n5129 199.739
R2486 VSS.n5151 VSS.n5135 199.739
R2487 VSS.n5185 VSS.n233 199.739
R2488 VSS.n5198 VSS.n226 199.739
R2489 VSS.n218 VSS.n217 199.739
R2490 VSS.n5231 VSS.n5230 199.739
R2491 VSS.n5262 VSS.n202 199.739
R2492 VSS.n5268 VSS.n199 199.739
R2493 VSS.n5284 VSS.n5283 199.739
R2494 VSS.n5298 VSS.n188 199.739
R2495 VSS.n185 VSS.n184 199.739
R2496 VSS.n5312 VSS.n5311 199.739
R2497 VSS.n5319 VSS.n5318 199.739
R2498 VSS.n449 VSS.n399 199.739
R2499 VSS.n401 VSS.n400 199.739
R2500 VSS.n404 VSS.n403 199.739
R2501 VSS.n407 VSS.n406 199.739
R2502 VSS.n3461 VSS.n3030 199.662
R2503 VSS.n5348 VSS.t797 199.144
R2504 VSS.n3118 VSS.n3117 199.052
R2505 VSS.n4037 VSS.n3988 198.964
R2506 VSS.n3320 VSS.n3090 198.964
R2507 VSS.n2544 VSS.n2240 198.964
R2508 VSS.n2493 VSS.n2268 198.964
R2509 VSS.n2449 VSS.n2289 198.964
R2510 VSS.n2692 VSS.n2683 198.964
R2511 VSS.n1978 VSS.n1373 198.964
R2512 VSS.n1902 VSS.n1405 198.964
R2513 VSS.n1884 VSS.n1415 198.964
R2514 VSS.n1657 VSS.n1522 198.964
R2515 VSS.n4923 VSS.n4884 198.964
R2516 VSS.n250 VSS.n249 198.964
R2517 VSS.n2889 VSS.n2888 198.696
R2518 VSS.n3636 VSS.n2946 198.654
R2519 VSS.n3481 VSS.n3020 198.654
R2520 VSS.n3417 VSS.n3049 198.654
R2521 VSS.n2648 VSS.n2647 198.654
R2522 VSS.n2803 VSS.n2802 198.654
R2523 VSS.n5505 VSS.n122 198.475
R2524 VSS.n3991 VSS.n3990 198.475
R2525 VSS.t3285 VSS.n4657 197.639
R2526 VSS.n3748 VSS.n3747 197.288
R2527 VSS.n3921 VSS.n3920 197.219
R2528 VSS.n4002 VSS.n4001 197.219
R2529 VSS.n4261 VSS.n3752 197.219
R2530 VSS.n3294 VSS.n3102 197.219
R2531 VSS.n2575 VSS.n2573 197.219
R2532 VSS.n2519 VSS.n2518 197.219
R2533 VSS.n2761 VSS.n2177 197.219
R2534 VSS.n1358 VSS.n1357 197.219
R2535 VSS.n2560 VSS.n2559 196.981
R2536 VSS.n3866 VSS.n3845 196.442
R2537 VSS.n3961 VSS.n3815 196.442
R2538 VSS.n3999 VSS.n3998 196.442
R2539 VSS.n3733 VSS.n3732 196.442
R2540 VSS.n3726 VSS.n3725 196.442
R2541 VSS.n4434 VSS.n4433 196.442
R2542 VSS.n3276 VSS.n3112 196.442
R2543 VSS.n3564 VSS.n2982 196.442
R2544 VSS.n3008 VSS.n3007 196.442
R2545 VSS.n3509 VSS.n3006 196.442
R2546 VSS.n3430 VSS.n3042 196.442
R2547 VSS.n3040 VSS.n3039 196.442
R2548 VSS.n3383 VSS.n3382 196.442
R2549 VSS.n3258 VSS.n3120 196.442
R2550 VSS.n3223 VSS.n3158 196.442
R2551 VSS.n2606 VSS.n2210 196.442
R2552 VSS.n2825 VSS.n2807 196.442
R2553 VSS.n2910 VSS.n2162 196.442
R2554 VSS.n2048 VSS.n2047 196.442
R2555 VSS.n1971 VSS.n1970 196.442
R2556 VSS.n1972 VSS.n1969 196.442
R2557 VSS.n1399 VSS.n1398 196.442
R2558 VSS.n1421 VSS.n1420 196.442
R2559 VSS.n1851 VSS.n1432 196.442
R2560 VSS.n1818 VSS.n1449 196.442
R2561 VSS.n1811 VSS.n1452 196.442
R2562 VSS.n1460 VSS.n1459 196.442
R2563 VSS.n1476 VSS.n1475 196.442
R2564 VSS.n1745 VSS.n1744 196.442
R2565 VSS.n1680 VSS.n1513 196.442
R2566 VSS.n1663 VSS.n1519 196.442
R2567 VSS.n1592 VSS.n1591 196.442
R2568 VSS.n4106 VSS.n3783 195.752
R2569 VSS.n2214 VSS.n2213 195.752
R2570 VSS.n2502 VSS.n2260 195.752
R2571 VSS.n2826 VSS.n2806 195.752
R2572 VSS.n2789 VSS.n2787 195.667
R2573 VSS.n3754 VSS.n3753 195.612
R2574 VSS.n3100 VSS.n3099 195.612
R2575 VSS.n2194 VSS.n2193 195.612
R2576 VSS.n4801 VSS.n4800 195
R2577 VSS.n1171 VSS.n1170 195
R2578 VSS.n4240 VSS.t1974 193.87
R2579 VSS.t894 VSS.t50 193.87
R2580 VSS.t331 VSS.t762 193.87
R2581 VSS.t267 VSS.t1633 193.87
R2582 VSS.t1074 VSS.n1037 192.364
R2583 VSS.n2970 VSS.n2968 190.761
R2584 VSS.n3594 VSS.n3593 190.601
R2585 VSS.n55 VSS.n54 190.399
R2586 VSS.n133 VSS.n132 190.399
R2587 VSS.n3797 VSS.n3796 190.399
R2588 VSS.n3823 VSS.n3822 190.399
R2589 VSS.n3295 VSS.n3098 190.399
R2590 VSS.n3359 VSS.n3358 190.399
R2591 VSS.n2964 VSS.n2963 190.399
R2592 VSS.n2637 VSS.n2196 190.399
R2593 VSS.n1919 VSS.n1918 190.399
R2594 VSS.n2198 VSS.n2197 189.99
R2595 VSS.n3332 VSS.n3331 189.8
R2596 VSS.n2713 VSS.n2669 189.481
R2597 VSS.n2509 VSS.n2254 189.407
R2598 VSS.n3943 VSS.n3942 189.201
R2599 VSS.n3447 VSS.n3446 189.201
R2600 VSS.n1987 VSS.n1367 189.201
R2601 VSS.n4655 VSS.t3054 187.067
R2602 VSS.n1186 VSS.t3251 187.067
R2603 VSS.n1002 VSS.n999 186.341
R2604 VSS.t474 VSS.t2067 185.441
R2605 VSS.t2221 VSS.n3715 185.441
R2606 VSS.t2767 VSS.t2090 185.441
R2607 VSS.t214 VSS.t2923 185.441
R2608 VSS.t1583 VSS.t2274 185.441
R2609 VSS.t2130 VSS.t2683 185.441
R2610 VSS.t885 VSS.t1016 185.441
R2611 VSS.t166 VSS.t2235 185.441
R2612 VSS.t1610 VSS.t2922 185.441
R2613 VSS.t419 VSS.t1753 185.441
R2614 VSS.n3952 VSS.n3951 185
R2615 VSS.n3954 VSS.n3953 185
R2616 VSS.n4028 VSS.n4027 185
R2617 VSS.n4030 VSS.n4029 185
R2618 VSS.n4387 VSS.n4386 185
R2619 VSS.n4385 VSS.n4384 185
R2620 VSS.n3646 VSS.n3645 185
R2621 VSS.n3644 VSS.n3643 185
R2622 VSS.n3620 VSS.n3619 185
R2623 VSS.n2972 VSS.n2971 185
R2624 VSS.n3571 VSS.n2977 185
R2625 VSS.n3573 VSS.n3572 185
R2626 VSS.n3554 VSS.n3553 185
R2627 VSS.n3552 VSS.n3551 185
R2628 VSS.n3526 VSS.n2997 185
R2629 VSS.n3528 VSS.n3527 185
R2630 VSS.n3496 VSS.n3012 185
R2631 VSS.n3498 VSS.n3497 185
R2632 VSS.n3488 VSS.n3014 185
R2633 VSS.n3490 VSS.n3489 185
R2634 VSS.n3329 VSS.n3328 185
R2635 VSS.n3327 VSS.n3326 185
R2636 VSS.n3313 VSS.n3312 185
R2637 VSS.n1642 VSS.n1641 185
R2638 VSS.n1640 VSS.n1639 185
R2639 VSS.n1077 VSS.n1045 183.341
R2640 VSS.n1077 VSS.n1076 183.341
R2641 VSS.t924 VSS.t797 180.306
R2642 VSS.n1079 VSS.t2971 178.808
R2643 VSS.n1079 VSS.t19 178.808
R2644 VSS.n4656 VSS.n4655 177.636
R2645 VSS.n1186 VSS.n1185 177.636
R2646 VSS.t1977 VSS.t2253 177.012
R2647 VSS.t2171 VSS.t1102 177.012
R2648 VSS.t2751 VSS.t1351 177.012
R2649 VSS.t1732 VSS.t1945 177.012
R2650 VSS.t1692 VSS.t1895 177.012
R2651 VSS.t401 VSS.t2 177.012
R2652 VSS.t747 VSS.t207 177.012
R2653 VSS.t1816 VSS.t2158 177.012
R2654 VSS.t2957 VSS.t1635 177.012
R2655 VSS.t2055 VSS.t1623 177.012
R2656 VSS.n4937 VSS.t2810 176.053
R2657 VSS.n1101 VSS.n1025 172.139
R2658 VSS.t14 VSS.t263 171.34
R2659 VSS.n1021 VSS.t1913 169.477
R2660 VSS.n4957 VSS.t18 168.983
R2661 VSS.t2816 VSS.t149 168.583
R2662 VSS.t1301 VSS.t1329 168.583
R2663 VSS.t1794 VSS.t1964 168.583
R2664 VSS.t2727 VSS.t171 168.583
R2665 VSS.t1985 VSS.t691 168.583
R2666 VSS.t1309 VSS.t630 168.583
R2667 VSS.t581 VSS.t1104 168.583
R2668 VSS.t1504 VSS.t81 168.583
R2669 VSS.t3030 VSS.n274 168.526
R2670 VSS.n4937 VSS.t397 168.012
R2671 VSS.n970 VSS.t2167 167.112
R2672 VSS.n970 VSS.t1846 166.275
R2673 VSS.n1226 VSS.n955 165.648
R2674 VSS.n1226 VSS.n1225 165.648
R2675 VSS.n1231 VSS.n954 165.648
R2676 VSS.n960 VSS.t798 165.571
R2677 VSS.n1938 VSS.t2209 164.097
R2678 VSS.t3130 VSS.n1073 163.947
R2679 VSS.n1060 VSS.n1059 163.742
R2680 VSS.t438 VSS.n999 162.889
R2681 VSS.t195 VSS.n999 162.889
R2682 VSS.t1255 VSS.t2696 162.774
R2683 VSS.t1882 VSS.t1112 162.774
R2684 VSS.t1570 VSS.t725 162.774
R2685 VSS.t2133 VSS.t2267 162.774
R2686 VSS.n5757 VSS.t2008 162.471
R2687 VSS.n61 VSS.t1614 162.471
R2688 VSS.n4020 VSS.t485 162.471
R2689 VSS.n4248 VSS.t1511 162.471
R2690 VSS.n4267 VSS.t2068 162.471
R2691 VSS.n4308 VSS.t1578 162.471
R2692 VSS.n3718 VSS.t2138 162.471
R2693 VSS.n3691 VSS.t948 162.471
R2694 VSS.n3088 VSS.t603 162.471
R2695 VSS.n3256 VSS.t1852 162.471
R2696 VSS.n2364 VSS.t108 162.471
R2697 VSS.n2363 VSS.t523 162.471
R2698 VSS.n2874 VSS.t3013 162.471
R2699 VSS.n2874 VSS.t2902 162.471
R2700 VSS.n2848 VSS.t300 162.471
R2701 VSS.n2848 VSS.t325 162.471
R2702 VSS.n1588 VSS.t356 162.471
R2703 VSS.n1549 VSS.t2859 162.471
R2704 VSS.n1619 VSS.t548 161.558
R2705 VSS.n2991 VSS.t1831 160.858
R2706 VSS.n4288 VSS.t1805 160.8
R2707 VSS.n2422 VSS.t1864 160.8
R2708 VSS.n1353 VSS.t1624 160.8
R2709 VSS.n1379 VSS.t1483 160.8
R2710 VSS.n1903 VSS.t1719 160.8
R2711 VSS.n1427 VSS.t968 160.8
R2712 VSS.n1803 VSS.t1171 160.8
R2713 VSS.n1468 VSS.t1306 160.8
R2714 VSS.n1759 VSS.t1246 160.8
R2715 VSS.n1697 VSS.t1963 160.8
R2716 VSS.n1650 VSS.t1636 160.8
R2717 VSS.t2611 VSS.t812 160.154
R2718 VSS.t3127 VSS.t2885 160.154
R2719 VSS.t2644 VSS.t2620 160.154
R2720 VSS.t571 VSS.t1939 160.154
R2721 VSS.t227 VSS.t2141 160.154
R2722 VSS.t2059 VSS.t2206 160.154
R2723 VSS.n14 VSS.t2006 160.017
R2724 VSS.n5653 VSS.t1612 160.017
R2725 VSS.n3993 VSS.t491 160.017
R2726 VSS.n3544 VSS.t1828 160.017
R2727 VSS.n3122 VSS.t1850 160.017
R2728 VSS.n2366 VSS.t110 160.017
R2729 VSS.n2876 VSS.t3014 160.017
R2730 VSS.n2881 VSS.t304 160.017
R2731 VSS.n4417 VSS.t950 160.017
R2732 VSS.n3319 VSS.t608 160.017
R2733 VSS.n2365 VSS.t526 160.017
R2734 VSS.n2876 VSS.t2848 160.017
R2735 VSS.n2881 VSS.t326 160.017
R2736 VSS.n1590 VSS.t358 160.017
R2737 VSS.n1621 VSS.t530 159.243
R2738 VSS.n4244 VSS.t1515 158.583
R2739 VSS.n3135 VSS.t465 158.583
R2740 VSS.n2354 VSS.t2976 158.583
R2741 VSS.n1574 VSS.t2787 158.583
R2742 VSS.n4347 VSS.t2136 158.583
R2743 VSS.n2362 VSS.t319 158.583
R2744 VSS.n1587 VSS.t2857 158.583
R2745 VSS.n1582 VSS.t433 158.583
R2746 VSS.n1270 VSS.t2926 158.583
R2747 VSS.t2809 VSS.t269 158.501
R2748 VSS.n965 VSS.t2591 158.361
R2749 VSS.n965 VSS.t1538 158.361
R2750 VSS.n331 VSS.t517 158.361
R2751 VSS.n331 VSS.t2931 158.361
R2752 VSS.n3748 VSS.t2066 158.186
R2753 VSS.t263 VSS.t1695 157.632
R2754 VSS.n2331 VSS.t323 157.291
R2755 VSS.n1580 VSS.t435 157.291
R2756 VSS.n1297 VSS.t2928 157.291
R2757 VSS.n3215 VSS.t2963 157.291
R2758 VSS.n3152 VSS.t463 157.291
R2759 VSS.n2080 VSS.t2789 157.291
R2760 VSS.n2077 VSS.t361 157.291
R2761 VSS.n2073 VSS.t72 157.291
R2762 VSS.n2367 VSS.t2558 157.291
R2763 VSS.n2335 VSS.t2974 157.291
R2764 VSS.n2847 VSS.t133 157.291
R2765 VSS.n1601 VSS.t1093 157.291
R2766 VSS.n1555 VSS.t2783 157.291
R2767 VSS.n1305 VSS.t677 157.291
R2768 VSS.n1312 VSS.t594 157.291
R2769 VSS.n4598 VSS.t1389 157.291
R2770 VSS.n987 VSS.t884 157.291
R2771 VSS.n3949 VSS.t1364 156.915
R2772 VSS.n4280 VSS.t388 156.915
R2773 VSS.n4864 VSS.t538 156.915
R2774 VSS.n4909 VSS.t519 156.915
R2775 VSS.n5100 VSS.t540 156.915
R2776 VSS.n5127 VSS.t544 156.915
R2777 VSS.n5211 VSS.t542 156.915
R2778 VSS.n5248 VSS.t521 156.915
R2779 VSS.n1999 VSS.t534 156.915
R2780 VSS.n1926 VSS.t536 156.915
R2781 VSS.n4956 VSS.t2970 156.108
R2782 VSS.n340 VSS.t2671 155.376
R2783 VSS.n3213 VSS.t2965 155.286
R2784 VSS.n2107 VSS.t2793 155.286
R2785 VSS.n2113 VSS.t363 155.286
R2786 VSS.n2119 VSS.t74 155.286
R2787 VSS.n2372 VSS.t2556 155.286
R2788 VSS.n2843 VSS.t131 155.286
R2789 VSS.n1541 VSS.t1095 155.286
R2790 VSS.n1267 VSS.t679 155.286
R2791 VSS.n1265 VSS.t596 155.286
R2792 VSS.n4597 VSS.t1391 155.286
R2793 VSS.n1215 VSS.t882 155.286
R2794 VSS.n4303 VSS.t1580 155.286
R2795 VSS.n4526 VSS.t1238 154.561
R2796 VSS.n4532 VSS.t2677 154.561
R2797 VSS.n5382 VSS.t1029 154.561
R2798 VSS.n5370 VSS.t1761 154.561
R2799 VSS.n3851 VSS.t2637 154.561
R2800 VSS.n3851 VSS.t1202 154.561
R2801 VSS.n3843 VSS.t1139 154.561
R2802 VSS.n3843 VSS.t2694 154.561
R2803 VSS.n4447 VSS.t2275 154.561
R2804 VSS.n4447 VSS.t2129 154.561
R2805 VSS.n4453 VSS.t1670 154.561
R2806 VSS.n4453 VSS.t2648 154.561
R2807 VSS.n3144 VSS.t1356 154.561
R2808 VSS.n3144 VSS.t1896 154.561
R2809 VSS.n2087 VSS.t2107 154.561
R2810 VSS.n2087 VSS.t1657 154.561
R2811 VSS.n2097 VSS.t1451 154.561
R2812 VSS.n2097 VSS.t1519 154.561
R2813 VSS.n2492 VSS.t2124 154.561
R2814 VSS.n2340 VSS.t1123 154.561
R2815 VSS.n2340 VSS.t2631 154.561
R2816 VSS.n2858 VSS.t936 154.561
R2817 VSS.n2858 VSS.t1376 154.561
R2818 VSS.n2866 VSS.t1049 154.561
R2819 VSS.n2866 VSS.t742 154.561
R2820 VSS.n1771 VSS.t1706 154.561
R2821 VSS.n1589 VSS.t2016 154.561
R2822 VSS.n1560 VSS.t1453 154.561
R2823 VSS.n1560 VSS.t2112 154.561
R2824 VSS.n1283 VSS.t946 154.561
R2825 VSS.n1283 VSS.t1586 154.561
R2826 VSS.n1289 VSS.t2173 154.561
R2827 VSS.n1289 VSS.t804 154.561
R2828 VSS.n4828 VSS.t934 154.561
R2829 VSS.n4929 VSS.t1328 154.561
R2830 VSS.n4902 VSS.t1700 154.561
R2831 VSS.n5018 VSS.t896 154.561
R2832 VSS.n5046 VSS.t1924 154.561
R2833 VSS.n5077 VSS.t2270 154.561
R2834 VSS.n5107 VSS.t728 154.561
R2835 VSS.n5130 VSS.t1885 154.561
R2836 VSS.n5181 VSS.t2699 154.561
R2837 VSS.n5217 VSS.t904 154.561
R2838 VSS.n5264 VSS.t2564 154.561
R2839 VSS.n190 VSS.t2258 154.561
R2840 VSS.n5305 VSS.t2606 154.561
R2841 VSS.n180 VSS.t1542 154.561
R2842 VSS.n178 VSS.t925 154.561
R2843 VSS.n442 VSS.t2570 154.561
R2844 VSS.n436 VSS.t2199 154.561
R2845 VSS.n430 VSS.t771 154.561
R2846 VSS.n3945 VSS.t1854 154.131
R2847 VSS.n3115 VSS.t1733 154.131
R2848 VSS.n1364 VSS.t406 154.131
R2849 VSS.n1393 VSS.t1824 154.131
R2850 VSS.n1876 VSS.t1513 154.131
R2851 VSS.n4860 VSS.t102 154.131
R2852 VSS.n4911 VSS.t2811 154.131
R2853 VSS.n247 VSS.t224 154.131
R2854 VSS.n5170 VSS.t17 154.131
R2855 VSS.n220 VSS.t2871 154.131
R2856 VSS.n5244 VSS.t650 154.131
R2857 VSS.n1490 VSS.t2720 153.399
R2858 VSS.n4619 VSS.n1249 152.596
R2859 VSS.n4617 VSS.n462 152.596
R2860 VSS.n4613 VSS.n4612 152.596
R2861 VSS.n3271 VSS.t567 152.381
R2862 VSS.n1871 VSS.t546 152.381
R2863 VSS.n1430 VSS.t528 152.381
R2864 VSS.n1735 VSS.t532 152.381
R2865 VSS.n5667 VSS.n5666 152
R2866 VSS.n5484 VSS.n5483 152
R2867 VSS.n3938 VSS.n3937 152
R2868 VSS.n4085 VSS.n4084 152
R2869 VSS.n3609 VSS.n3608 152
R2870 VSS.n3360 VSS.n3075 152
R2871 VSS.n3302 VSS.n3301 152
R2872 VSS.n2887 VSS.n2886 152
R2873 VSS.n2640 VSS.n2639 152
R2874 VSS.n1920 VSS.n1397 152
R2875 VSS.n4629 VSS.n4627 151.964
R2876 VSS.t2088 VSS.t783 151.725
R2877 VSS.t970 VSS.t477 151.725
R2878 VSS.t1440 VSS.t1932 151.725
R2879 VSS.t2907 VSS.t1596 151.725
R2880 VSS.t237 VSS.t1225 151.725
R2881 VSS.n966 VSS.t1844 150.922
R2882 VSS.n962 VSS.t1848 150.922
R2883 VSS.t2080 VSS.t1215 150.897
R2884 VSS.t2933 VSS.t1873 150.78
R2885 VSS.t2968 VSS.t715 150.78
R2886 VSS.t2200 VSS.t458 150.78
R2887 VSS.t1325 VSS.t1323 150.577
R2888 VSS.n3582 VSS.n2972 150.4
R2889 VSS.n3860 VSS.t1744 150.376
R2890 VSS.n4459 VSS.t734 150.376
R2891 VSS.n3159 VSS.t875 150.376
R2892 VSS.n3150 VSS.t1084 150.376
R2893 VSS.n2357 VSS.t1521 150.376
R2894 VSS.n2349 VSS.t2186 150.376
R2895 VSS.n1599 VSS.t1942 150.376
R2896 VSS.n1552 VSS.t736 150.376
R2897 VSS.n1569 VSS.t1994 150.376
R2898 VSS.n1295 VSS.t831 150.376
R2899 VSS.n4276 VSS.t1593 150.101
R2900 VSS.n1859 VSS.t2921 150.101
R2901 VSS.t985 VSS.t3097 149.534
R2902 VSS.n1074 VSS.n274 148.376
R2903 VSS.t2737 VSS.t3241 148.287
R2904 VSS.n4049 VSS.t592 147.411
R2905 VSS.n976 VSS.n975 146.25
R2906 VSS.n1225 VSS.n1224 146.25
R2907 VSS.n1224 VSS.n1223 146.25
R2908 VSS.n4614 VSS.n4613 146.25
R2909 VSS.n4617 VSS.n4616 146.25
R2910 VSS.n4620 VSS.n4619 146.25
R2911 VSS.n4647 VSS.n4646 146.25
R2912 VSS.n4648 VSS.n4647 146.25
R2913 VSS.n4812 VSS.n4811 146.25
R2914 VSS.n4813 VSS.n4812 146.25
R2915 VSS.n4594 VSS.n4593 146.25
R2916 VSS.n4593 VSS.n1260 146.25
R2917 VSS.n1088 VSS.n1043 146.25
R2918 VSS.n1043 VSS.n1042 146.25
R2919 VSS.n1044 VSS.n1040 146.25
R2920 VSS.n1040 VSS.n1036 146.25
R2921 VSS.n1047 VSS.n1045 146.25
R2922 VSS.n1067 VSS.n1047 146.25
R2923 VSS.n1076 VSS.n1048 146.25
R2924 VSS.n1075 VSS.n1048 146.25
R2925 VSS.n955 VSS.n951 146.25
R2926 VSS.n1233 VSS.n951 146.25
R2927 VSS.n1232 VSS.n1231 146.25
R2928 VSS.n1233 VSS.n1232 146.25
R2929 VSS.n1008 VSS.n1007 146.25
R2930 VSS.n1009 VSS.n1008 146.25
R2931 VSS.n1205 VSS.n1204 146.25
R2932 VSS.n1204 VSS.n1203 146.25
R2933 VSS.n996 VSS.n995 146.25
R2934 VSS.n995 VSS.n993 146.25
R2935 VSS.n1212 VSS.n1211 146.25
R2936 VSS.n1211 VSS.n1210 146.25
R2937 VSS.n1201 VSS.n1200 146.25
R2938 VSS.n1202 VSS.n1201 146.25
R2939 VSS.n1198 VSS.n1197 146.25
R2940 VSS.n1197 VSS.n1196 146.25
R2941 VSS.n4797 VSS.n4796 146.038
R2942 VSS.t269 VSS.t1456 145.821
R2943 VSS.n4916 VSS.t398 145.212
R2944 VSS.n5083 VSS.t232 145.212
R2945 VSS.n2552 VSS.t2722 145.212
R2946 VSS.n2484 VSS.t2869 145.212
R2947 VSS.n2184 VSS.t168 145.212
R2948 VSS.n1985 VSS.t96 145.212
R2949 VSS.n1877 VSS.t2908 145.212
R2950 VSS.t3154 VSS.t933 145.172
R2951 VSS.t2668 VSS.t2670 144.659
R2952 VSS.t2672 VSS.t2668 144.659
R2953 VSS.t2696 VSS.t2698 143.925
R2954 VSS.t1884 VSS.t1882 143.925
R2955 VSS.t543 VSS.t16 143.925
R2956 VSS.t725 VSS.t727 143.925
R2957 VSS.t223 VSS.t539 143.925
R2958 VSS.t2267 VSS.t2269 143.925
R2959 VSS.n2646 VSS.t1536 143.299
R2960 VSS.t653 VSS.t12 143.296
R2961 VSS.t2779 VSS.t1211 143.296
R2962 VSS.t2079 VSS.t1639 143.296
R2963 VSS.t1788 VSS.t2153 143.296
R2964 VSS.t826 VSS.t1036 143.296
R2965 VSS.t1937 VSS.t1407 143.296
R2966 VSS.n2777 VSS.t2874 142.821
R2967 VSS.n2566 VSS.t11 142.821
R2968 VSS.n1891 VSS.t1507 142.821
R2969 VSS.n2509 VSS.n2508 140.8
R2970 VSS.n1189 VSS.n1188 140.048
R2971 VSS.n4653 VSS.n4652 140.048
R2972 VSS.n4254 VSS.t1320 139.548
R2973 VSS.n1099 VSS.n1098 139.548
R2974 VSS.t1806 VSS.t2704 139.081
R2975 VSS.n4950 VSS.n368 139.06
R2976 VSS.t2689 VSS.t2687 138.964
R2977 VSS.t2687 VSS.t2685 138.964
R2978 VSS.n1089 VSS.n1044 138.166
R2979 VSS.n1089 VSS.n1088 138.166
R2980 VSS.t2589 VSS.t2678 134.867
R2981 VSS.t1728 VSS.t977 134.867
R2982 VSS.t1833 VSS.t239 134.867
R2983 VSS.t1003 VSS.t2208 134.867
R2984 VSS.n1210 VSS.t199 133.925
R2985 VSS.n1210 VSS.t197 133.925
R2986 VSS.n1202 VSS.t446 133.925
R2987 VSS.t438 VSS.n1202 133.925
R2988 VSS.n1196 VSS.t195 133.925
R2989 VSS.n1196 VSS.t193 133.925
R2990 VSS.t1327 VSS.t1325 133.142
R2991 VSS.n4967 VSS.n4966 133.026
R2992 VSS.t101 VSS.t537 132.76
R2993 VSS.t2949 VSS.t2953 132.048
R2994 VSS.t2943 VSS.t2945 132.048
R2995 VSS.t2947 VSS.t2951 132.048
R2996 VSS.t2941 VSS.t2939 132.048
R2997 VSS.t231 VSS.t514 130.219
R2998 VSS.n4611 VSS.n4610 130
R2999 VSS.n1221 VSS.n1220 130
R3000 VSS.n1102 VSS.n1101 129.748
R3001 VSS.n1099 VSS.n1024 129.385
R3002 VSS.n1059 VSS.n299 128.982
R3003 VSS.n4992 VSS.n4991 128
R3004 VSS.n4991 VSS.n301 128
R3005 VSS.t2805 VSS.t1187 126.438
R3006 VSS.t2749 VSS.t2135 126.438
R3007 VSS.t1851 VSS.t1498 126.438
R3008 VSS.t3124 VSS.t148 126.438
R3009 VSS.t1249 VSS.t1707 126.438
R3010 VSS.n1060 VSS.n1057 126.291
R3011 VSS.n1233 VSS.t713 125.01
R3012 VSS.n1063 VSS.n1062 124.236
R3013 VSS.n16 VSS.t3600 121.927
R3014 VSS.n34 VSS.t3633 121.927
R3015 VSS.n44 VSS.t3714 121.927
R3016 VSS.n96 VSS.t3564 121.927
R3017 VSS.n141 VSS.t3680 121.927
R3018 VSS.n3127 VSS.t3651 121.927
R3019 VSS.n1423 VSS.t3731 121.927
R3020 VSS.n289 VSS.t3612 121.927
R3021 VSS.n281 VSS.t3719 121.927
R3022 VSS.n267 VSS.t3816 121.927
R3023 VSS.n260 VSS.t3759 121.927
R3024 VSS.n5132 VSS.t3613 121.927
R3025 VSS.n5144 VSS.t3784 121.927
R3026 VSS.t245 VSS.t259 121.624
R3027 VSS.t259 VSS.t249 121.624
R3028 VSS.t249 VSS.t257 121.624
R3029 VSS.t257 VSS.t251 121.624
R3030 VSS.t255 VSS.t253 121.624
R3031 VSS.t247 VSS.t255 121.624
R3032 VSS.t307 VSS.t247 121.624
R3033 VSS.t313 VSS.t307 121.624
R3034 VSS.t309 VSS.t313 121.624
R3035 VSS.t311 VSS.t309 121.624
R3036 VSS.t452 VSS.t311 121.624
R3037 VSS.t450 VSS.t452 121.624
R3038 VSS.t2878 VSS.t450 121.624
R3039 VSS.t440 VSS.t449 121.624
R3040 VSS.t448 VSS.t440 121.624
R3041 VSS.t659 VSS.t663 121.624
R3042 VSS.t671 VSS.t659 121.624
R3043 VSS.t673 VSS.t671 121.624
R3044 VSS.t657 VSS.t673 121.624
R3045 VSS.t656 VSS.t657 121.624
R3046 VSS.t665 VSS.t656 121.624
R3047 VSS.t664 VSS.t665 121.624
R3048 VSS.t281 VSS.t664 121.624
R3049 VSS.t279 VSS.t281 121.624
R3050 VSS.t286 VSS.t279 121.624
R3051 VSS.t288 VSS.t286 121.624
R3052 VSS.t292 VSS.t288 121.624
R3053 VSS.t284 VSS.t292 121.624
R3054 VSS.t278 VSS.t284 121.624
R3055 VSS.t277 VSS.t278 121.624
R3056 VSS.t2990 VSS.t277 121.624
R3057 VSS.t2989 VSS.t2990 121.624
R3058 VSS.t2988 VSS.t2989 121.624
R3059 VSS.t2991 VSS.t121 121.624
R3060 VSS.t121 VSS.t125 121.624
R3061 VSS.t125 VSS.t2936 121.624
R3062 VSS.t2835 VSS.t2833 121.624
R3063 VSS.t2833 VSS.t456 121.624
R3064 VSS.t441 VSS.t437 121.624
R3065 VSS.t437 VSS.t436 121.624
R3066 VSS.t555 VSS.t554 121.624
R3067 VSS.t557 VSS.t555 121.624
R3068 VSS.t2899 VSS.t457 121.624
R3069 VSS.t2897 VSS.t2899 121.624
R3070 VSS.t122 VSS.t2935 121.624
R3071 VSS.t120 VSS.t122 121.624
R3072 VSS.t2987 VSS.t120 121.624
R3073 VSS.t2986 VSS.t2995 121.624
R3074 VSS.t2995 VSS.t2992 121.624
R3075 VSS.t2992 VSS.t294 121.624
R3076 VSS.t294 VSS.t285 121.624
R3077 VSS.t285 VSS.t291 121.624
R3078 VSS.t291 VSS.t283 121.624
R3079 VSS.t283 VSS.t280 121.624
R3080 VSS.t280 VSS.t287 121.624
R3081 VSS.t287 VSS.t282 121.624
R3082 VSS.t282 VSS.t293 121.624
R3083 VSS.t293 VSS.t660 121.624
R3084 VSS.t660 VSS.t658 121.624
R3085 VSS.t658 VSS.t662 121.624
R3086 VSS.t662 VSS.t661 121.624
R3087 VSS.t661 VSS.t666 121.624
R3088 VSS.t666 VSS.t668 121.624
R3089 VSS.t668 VSS.t672 121.624
R3090 VSS.t672 VSS.t667 121.624
R3091 VSS.t558 VSS.t550 121.624
R3092 VSS.t550 VSS.t551 121.624
R3093 VSS.t2825 VSS.t2794 121.624
R3094 VSS.t2794 VSS.t2796 121.624
R3095 VSS.t2796 VSS.t370 121.624
R3096 VSS.t370 VSS.t372 121.624
R3097 VSS.t372 VSS.t368 121.624
R3098 VSS.t368 VSS.t366 121.624
R3099 VSS.t366 VSS.t3275 121.624
R3100 VSS.t3275 VSS.t3273 121.624
R3101 VSS.t3273 VSS.t3281 121.624
R3102 VSS.t3283 VSS.t3277 121.624
R3103 VSS.t3277 VSS.t3271 121.624
R3104 VSS.t3271 VSS.t3279 121.624
R3105 VSS.t3279 VSS.t3285 121.624
R3106 VSS.n5349 VSS.t2691 121.102
R3107 VSS.t397 VSS.t506 120.462
R3108 VSS.n1068 VSS.n1067 119.96
R3109 VSS.t770 VSS.t2876 118.38
R3110 VSS.t2666 VSS.t2672 118.24
R3111 VSS.n977 VSS.t2592 118.064
R3112 VSS.t1649 VSS.t3436 118.008
R3113 VSS.t2958 VSS.t2709 118.008
R3114 VSS.t1702 VSS.t83 118.008
R3115 VSS.t1243 VSS.t840 118.008
R3116 VSS.t1241 VSS.t838 118.008
R3117 VSS.t374 VSS.t2098 118.008
R3118 VSS.n4021 VSS.n3995 117.889
R3119 VSS.n1651 VSS.n1527 117.889
R3120 VSS.n2713 VSS.n2712 117.334
R3121 VSS.t68 VSS.t953 117.135
R3122 VSS.n4651 VSS.n4650 117.001
R3123 VSS.n4650 VSS.t3244 117.001
R3124 VSS.n4643 VSS.n1246 117.001
R3125 VSS.t3244 VSS.n1246 117.001
R3126 VSS.n360 VSS.n354 117.001
R3127 VSS.n360 VSS.n358 117.001
R3128 VSS.n4955 VSS.n4954 117.001
R3129 VSS.n4956 VSS.n4955 117.001
R3130 VSS.n4940 VSS.n367 117.001
R3131 VSS.n4941 VSS.n4940 117.001
R3132 VSS.n4972 VSS.n4971 117.001
R3133 VSS.n4971 VSS.n4970 117.001
R3134 VSS.n4947 VSS.n4946 117.001
R3135 VSS.n4948 VSS.n4947 117.001
R3136 VSS.n1229 VSS.n1228 117.001
R3137 VSS.n1228 VSS.t2165 117.001
R3138 VSS.n1227 VSS.n1226 117.001
R3139 VSS.t2165 VSS.n1227 117.001
R3140 VSS.n954 VSS.n952 117.001
R3141 VSS.t2165 VSS.n952 117.001
R3142 VSS.n1190 VSS.n1011 117.001
R3143 VSS.n1011 VSS.t3396 117.001
R3144 VSS.n1113 VSS.n1010 117.001
R3145 VSS.n1010 VSS.t3396 117.001
R3146 VSS.n4263 VSS.t3562 116.734
R3147 VSS.n1681 VSS.t3691 116.734
R3148 VSS.n1319 VSS.t3707 116.734
R3149 VSS.n2229 VSS.t3619 115.885
R3150 VSS.n4993 VSS.n4992 115.201
R3151 VSS.n4992 VSS.n300 115.201
R3152 VSS.n2533 VSS.n2246 114.377
R3153 VSS.n2660 VSS.n2659 114.377
R3154 VSS.n2244 VSS.n2243 114.376
R3155 VSS.t3244 VSS.t890 113.397
R3156 VSS.n3369 VSS.n3071 113.195
R3157 VSS.n2785 VSS.n2784 113.195
R3158 VSS.n2819 VSS.n2810 113.195
R3159 VSS.n2971 VSS.n2970 111.43
R3160 VSS.n3242 VSS.n3129 110.584
R3161 VSS.n3462 VSS.n3029 109.684
R3162 VSS.n3065 VSS.n3064 109.684
R3163 VSS.n2458 VSS.n2286 109.684
R3164 VSS.n2740 VSS.n2739 109.684
R3165 VSS.n1447 VSS.n1446 109.684
R3166 VSS.t3097 VSS.n4590 109.657
R3167 VSS.t1841 VSS.t201 109.579
R3168 VSS.t2723 VSS.t788 109.579
R3169 VSS.t2911 VSS.t2599 109.579
R3170 VSS.t377 VSS.t2263 109.579
R3171 VSS.t2150 VSS.t498 109.579
R3172 VSS.t415 VSS.t1465 109.579
R3173 VSS.t1906 VSS.t513 109.579
R3174 VSS.t265 VSS.t403 109.579
R3175 VSS.t32 VSS.t1530 109.579
R3176 VSS.t1752 VSS.t910 109.579
R3177 VSS.n309 VSS.n300 108.8
R3178 VSS.n1052 VSS.t1296 108.642
R3179 VSS.t1294 VSS.n1052 108.642
R3180 VSS.n2243 VSS.t639 108.505
R3181 VSS.n2246 VSS.t226 108.505
R3182 VSS.n2659 VSS.t2813 108.505
R3183 VSS.n4989 VSS.t2837 105.632
R3184 VSS.n4985 VSS.t2843 105.632
R3185 VSS.n2956 VSS.n2955 105.097
R3186 VSS.n3095 VSS.n3094 102.678
R3187 VSS.n1616 VSS.t3702 102.379
R3188 VSS.n3890 VSS.t3690 102.353
R3189 VSS.n323 VSS.t1075 102.332
R3190 VSS.n4063 VSS.t611 101.43
R3191 VSS.t2125 VSS.t1843 101.15
R3192 VSS.t2650 VSS.t922 101.15
R3193 VSS.t316 VSS.t116 101.15
R3194 VSS.t4 VSS.t1076 101.15
R3195 VSS.t616 VSS.t749 101.15
R3196 VSS.n2981 VSS.t175 101.15
R3197 VSS.t379 VSS.t760 101.15
R3198 VSS.t24 VSS.t162 101.15
R3199 VSS.t2641 VSS.t1014 101.15
R3200 VSS.t892 VSS.t91 101.15
R3201 VSS.t2719 VSS.t1929 101.15
R3202 VSS.t1676 VSS.t1157 101.15
R3203 VSS.t792 VSS.t1484 101.15
R3204 VSS.t2108 VSS.t1217 101.15
R3205 VSS.n3969 VSS.t637 100.001
R3206 VSS.n3773 VSS.t330 100.001
R3207 VSS.n3766 VSS.t336 100.001
R3208 VSS.n4177 VSS.t2780 100.001
R3209 VSS.n3738 VSS.t2772 100.001
R3210 VSS.n4388 VSS.t2742 100.001
R3211 VSS.n2942 VSS.t180 100.001
R3212 VSS.n2961 VSS.t2776 100.001
R3213 VSS.n2987 VSS.t2815 100.001
R3214 VSS.n2994 VSS.t2248 100.001
R3215 VSS.n3045 VSS.t332 100.001
R3216 VSS.n3124 VSS.t346 100.001
R3217 VSS.n2204 VSS.t2242 100.001
R3218 VSS.n2305 VSS.t334 100.001
R3219 VSS.n2187 VSS.t2250 100.001
R3220 VSS.n2032 VSS.t182 100.001
R3221 VSS.n1349 VSS.t174 100.001
R3222 VSS.n1960 VSS.t190 100.001
R3223 VSS.n1386 VSS.t184 100.001
R3224 VSS.n1402 VSS.t2234 100.001
R3225 VSS.n1424 VSS.t2240 100.001
R3226 VSS.n1453 VSS.t633 100.001
R3227 VSS.n1465 VSS.t348 100.001
R3228 VSS.n1478 VSS.t635 100.001
R3229 VSS.n1499 VSS.t84 100.001
R3230 VSS.n1502 VSS.t55 100.001
R3231 VSS.n1523 VSS.t78 100.001
R3232 VSS.n4170 VSS.t3002 99.9005
R3233 VSS.n4187 VSS.t1738 99.9005
R3234 VSS.n3720 VSS.t1190 99.9005
R3235 VSS.n4357 VSS.t784 99.9005
R3236 VSS.n3046 VSS.t1194 99.9005
R3237 VSS.n2811 VSS.t709 99.9005
R3238 VSS.n2157 VSS.t889 99.9005
R3239 VSS.n1438 VSS.t1047 99.9005
R3240 VSS.n1481 VSS.t841 99.9005
R3241 VSS.n3058 VSS.t1650 99.7996
R3242 VSS.n4047 VSS.t3662 99.7825
R3243 VSS.n2379 VSS.t3754 99.7825
R3244 VSS.n2839 VSS.t3717 99.7825
R3245 VSS.n2123 VSS.t3583 98.8619
R3246 VSS.n2384 VSS.t3569 98.5139
R3247 VSS.t2970 VSS.t2932 98.1717
R3248 VSS.n1078 VSS.n1077 97.5005
R3249 VSS.n1079 VSS.n1078 97.5005
R3250 VSS.n1081 VSS.n1080 97.5005
R3251 VSS.n1080 VSS.n1079 97.5005
R3252 VSS.n1074 VSS.n1065 97.3256
R3253 VSS.n4386 VSS.n4385 97.1434
R3254 VSS.n3489 VSS.n3488 97.1434
R3255 VSS.n3497 VSS.n3496 97.1434
R3256 VSS.n3527 VSS.n3526 97.1434
R3257 VSS.n3553 VSS.n3552 97.1434
R3258 VSS.n3645 VSS.n3644 97.1434
R3259 VSS.n1230 VSS.n1229 97.1299
R3260 VSS.n1229 VSS.n956 97.1299
R3261 VSS.n1190 VSS.n1189 95.2476
R3262 VSS.n4652 VSS.n4651 95.2476
R3263 VSS.t490 VSS.t772 92.7208
R3264 VSS.t729 VSS.t220 92.7208
R3265 VSS.t3503 VSS.t2807 92.7208
R3266 VSS.t1786 VSS.t87 92.7208
R3267 VSS.t1177 VSS.t1222 92.7208
R3268 VSS.t781 VSS.t1488 92.7208
R3269 VSS.n1093 VSS.n1092 90.9607
R3270 VSS.n4954 VSS.n355 90.3534
R3271 VSS.n4954 VSS.n362 90.3534
R3272 VSS.n4965 VSS.n354 90.3534
R3273 VSS.n4960 VSS.n354 90.3534
R3274 VSS.n4951 VSS.n367 90.3534
R3275 VSS.n4944 VSS.n367 90.3534
R3276 VSS.t253 VSS.n1108 89.9516
R3277 VSS.n1150 VSS.t2991 89.9516
R3278 VSS.n4659 VSS.t2987 89.9516
R3279 VSS.t1388 VSS.n4611 88.474
R3280 VSS.n4814 VSS.t2937 87.2279
R3281 VSS.t1925 VSS.t1468 87.0113
R3282 VSS.t897 VSS.t1603 87.0113
R3283 VSS.n3593 VSS.t165 85.7148
R3284 VSS.n974 VSS.n954 85.0829
R3285 VSS.n4800 VSS.t2943 84.888
R3286 VSS.n1170 VSS.t2947 84.888
R3287 VSS.n4195 VSS.n4187 84.6851
R3288 VSS.n3423 VSS.n3046 84.6851
R3289 VSS.n2812 VSS.n2811 84.6851
R3290 VSS.n1843 VSS.n1438 84.6851
R3291 VSS.n1757 VSS.n1481 84.6851
R3292 VSS.t118 VSS.t786 84.2917
R3293 VSS.t1660 VSS.t1592 84.2917
R3294 VSS.t1143 VSS.t1849 84.2917
R3295 VSS.t494 VSS.t1052 84.2917
R3296 VSS.t1267 VSS.t1756 84.2917
R3297 VSS.t3476 VSS.t2823 84.2917
R3298 VSS.t1531 VSS.t1166 84.2917
R3299 VSS.t961 VSS.t3229 84.2917
R3300 VSS.n3085 VSS.t117 83.899
R3301 VSS.n4938 VSS.n4937 83.6874
R3302 VSS.n1061 VSS.n1050 83.5719
R3303 VSS.n1052 VSS.n1050 83.5719
R3304 VSS.n1051 VSS.n1049 83.5719
R3305 VSS.n1052 VSS.n1049 83.5719
R3306 VSS.n304 VSS.n303 83.5719
R3307 VSS.n4988 VSS.n303 83.5719
R3308 VSS.n1058 VSS.n296 83.5719
R3309 VSS.n4995 VSS.n296 83.5719
R3310 VSS.n4994 VSS.n4993 83.5719
R3311 VSS.n4995 VSS.n4994 83.5719
R3312 VSS.n4987 VSS.n300 83.5719
R3313 VSS.n4988 VSS.n4987 83.5719
R3314 VSS.n4945 VSS.n368 83.1211
R3315 VSS.n4233 VSS.n4170 82.5518
R3316 VSS.n3721 VSS.n3720 82.5518
R3317 VSS.n4358 VSS.n4357 82.5518
R3318 VSS.n2921 VSS.n2157 82.5518
R3319 VSS.n1686 VSS.n1509 81.965
R3320 VSS.n4641 VSS.n4634 81.2805
R3321 VSS.n1182 VSS.n1181 81.2805
R3322 VSS.n4643 VSS.n4642 80.9605
R3323 VSS.n4644 VSS.n4643 80.9605
R3324 VSS.n1113 VSS.n1012 80.9605
R3325 VSS.n1114 VSS.n1113 80.9605
R3326 VSS.t971 VSS.t2881 80.6
R3327 VSS.n975 VSS.n974 80.5652
R3328 VSS.n4620 VSS.n1251 79.0593
R3329 VSS.n4616 VSS.n1251 79.0593
R3330 VSS.n4616 VSS.n4615 79.0593
R3331 VSS.n4615 VSS.n4614 79.0593
R3332 VSS.n1206 VSS.n996 79.0593
R3333 VSS.n1206 VSS.n1205 79.0593
R3334 VSS.n1205 VSS.n997 79.0593
R3335 VSS.n1007 VSS.n997 79.0593
R3336 VSS.n1085 VSS.n1044 78.6829
R3337 VSS.n1088 VSS.n1087 78.6829
R3338 VSS.n3058 VSS.t1646 77.6313
R3339 VSS.n4967 VSS.n350 77.418
R3340 VSS.n4170 VSS.t2586 77.0434
R3341 VSS.n4187 VSS.t2752 77.0434
R3342 VSS.n3720 VSS.t2760 77.0434
R3343 VSS.n4357 VSS.t2746 77.0434
R3344 VSS.n3046 VSS.t763 77.0434
R3345 VSS.n2811 VSS.t2766 77.0434
R3346 VSS.n2157 VSS.t1069 77.0434
R3347 VSS.n1438 VSS.t724 77.0434
R3348 VSS.n1481 VSS.t839 77.0434
R3349 VSS.t1923 VSS.t1925 76.9364
R3350 VSS.t895 VSS.t897 76.9364
R3351 VSS.n4359 VSS.n4356 76.6108
R3352 VSS.t2829 VSS.n4625 76.5626
R3353 VSS.n3402 VSS.n3058 76.0226
R3354 VSS.t1814 VSS.t2864 75.8626
R3355 VSS.t1875 VSS.t454 75.8626
R3356 VSS.t60 VSS.t845 75.8626
R3357 VSS.t1609 VSS.t1564 75.8626
R3358 VSS.t580 VSS.t2181 75.8626
R3359 VSS.t790 VSS.t1516 75.8626
R3360 VSS.n993 VSS.t199 75.456
R3361 VSS.t197 VSS.n993 75.456
R3362 VSS.n1203 VSS.t446 75.456
R3363 VSS.n1203 VSS.t438 75.456
R3364 VSS.n1009 VSS.t195 75.456
R3365 VSS.t193 VSS.n1009 75.456
R3366 VSS.n4162 VSS.t2584 74.2862
R3367 VSS.n4243 VSS.t2770 74.2862
R3368 VSS.n4346 VSS.t2750 74.2862
R3369 VSS.n4371 VSS.t2768 74.2862
R3370 VSS.n4403 VSS.t1473 74.2862
R3371 VSS.n2141 VSS.t1025 74.2862
R3372 VSS.n2983 VSS.t2758 74.2862
R3373 VSS.n2993 VSS.t2764 74.2862
R3374 VSS.n3006 VSS.t748 74.2862
R3375 VSS.n3010 VSS.t1556 74.2862
R3376 VSS.n3039 VSS.t765 74.2862
R3377 VSS.n3053 VSS.t1648 74.2862
R3378 VSS.n2807 VSS.t2744 74.2862
R3379 VSS.n2162 VSS.t1067 74.2862
R3380 VSS.n1432 VSS.t722 74.2862
R3381 VSS.n1744 VSS.t837 74.2862
R3382 VSS.t2165 VSS.t713 74.0798
R3383 VSS.t2165 VSS.t2592 74.0798
R3384 VSS.n1082 VSS.n1045 73.4123
R3385 VSS.n1076 VSS.n1046 73.4123
R3386 VSS.n2199 VSS.n2198 73.1434
R3387 VSS.n1024 VSS.n1019 73.1255
R3388 VSS.n1102 VSS.n1023 73.1255
R3389 VSS.n1057 VSS.n1056 73.1255
R3390 VSS.n1056 VSS.n1055 73.1255
R3391 VSS.n1064 VSS.n1063 73.1255
R3392 VSS.n1065 VSS.n1064 73.1255
R3393 VSS.n4991 VSS.n4990 73.1255
R3394 VSS.n4990 VSS.n4989 73.1255
R3395 VSS.n4986 VSS.n305 73.1255
R3396 VSS.n4986 VSS.n4985 73.1255
R3397 VSS.n299 VSS.n297 73.1255
R3398 VSS.n1053 VSS.n297 73.1255
R3399 VSS.n4968 VSS.n4967 73.1255
R3400 VSS.n4969 VSS.n4968 73.1255
R3401 VSS.n369 VSS.n368 73.1255
R3402 VSS.n4938 VSS.n369 73.1255
R3403 VSS.n87 VSS.t473 72.8576
R3404 VSS.n3815 VSS.t344 72.8576
R3405 VSS.n4138 VSS.t338 72.8576
R3406 VSS.n4145 VSS.t629 72.8576
R3407 VSS.n4181 VSS.t2817 72.8576
R3408 VSS.n4184 VSS.t497 72.8576
R3409 VSS.n3732 VSS.t192 72.8576
R3410 VSS.n3695 VSS.t2778 72.8576
R3411 VSS.n4410 VSS.t503 72.8576
R3412 VSS.n2133 VSS.t501 72.8576
R3413 VSS.n2137 VSS.t469 72.8576
R3414 VSS.n3667 VSS.t188 72.8576
R3415 VSS.n2958 VSS.t172 72.8576
R3416 VSS.n2982 VSS.t176 72.8576
R3417 VSS.n2999 VSS.t2246 72.8576
R3418 VSS.n3002 VSS.t495 72.8576
R3419 VSS.n3436 VSS.t1366 72.8576
R3420 VSS.n3042 VSS.t342 72.8576
R3421 VSS.n3120 VSS.t352 72.8576
R3422 VSS.n2210 VSS.t2238 72.8576
R3423 VSS.n2276 VSS.t569 72.8576
R3424 VSS.n2300 VSS.t627 72.8576
R3425 VSS.n2662 VSS.t2236 72.8576
R3426 VSS.n2047 VSS.t2828 72.8576
R3427 VSS.n1346 VSS.t186 72.8576
R3428 VSS.n1363 VSS.t467 72.8576
R3429 VSS.n1970 VSS.t178 72.8576
R3430 VSS.n1381 VSS.t2774 72.8576
R3431 VSS.n1398 VSS.t2244 72.8576
R3432 VSS.n1420 VSS.t2232 72.8576
R3433 VSS.n1626 VSS.t340 72.8576
R3434 VSS.n1836 VSS.t471 72.8576
R3435 VSS.n1449 VSS.t328 72.8576
R3436 VSS.n1459 VSS.t350 72.8576
R3437 VSS.n1471 VSS.t631 72.8576
R3438 VSS.n1743 VSS.t1362 72.8576
R3439 VSS.n1721 VSS.t49 72.8576
R3440 VSS.n1713 VSS.t80 72.8576
R3441 VSS.n1519 VSS.t53 72.8576
R3442 VSS.n5255 VSS.t1746 72.8576
R3443 VSS.t515 VSS.t18 72.4219
R3444 VSS.n3969 VSS.t877 70.0005
R3445 VSS.n3773 VSS.t921 70.0005
R3446 VSS.n3766 VSS.t2020 70.0005
R3447 VSS.n4177 VSS.t1400 70.0005
R3448 VSS.n3738 VSS.t1797 70.0005
R3449 VSS.n4388 VSS.t1130 70.0005
R3450 VSS.n2942 VSS.t1683 70.0005
R3451 VSS.n2961 VSS.t1459 70.0005
R3452 VSS.n2987 VSS.t1344 70.0005
R3453 VSS.n2994 VSS.t997 70.0005
R3454 VSS.n3045 VSS.t1079 70.0005
R3455 VSS.n3124 VSS.t707 70.0005
R3456 VSS.n2204 VSS.t1291 70.0005
R3457 VSS.n2305 VSS.t1868 70.0005
R3458 VSS.n2187 VSS.t2230 70.0005
R3459 VSS.n2032 VSS.t819 70.0005
R3460 VSS.n1349 VSS.t1622 70.0005
R3461 VSS.n1960 VSS.t1481 70.0005
R3462 VSS.n1386 VSS.t2211 70.0005
R3463 VSS.n1402 VSS.t1717 70.0005
R3464 VSS.n1424 VSS.t962 70.0005
R3465 VSS.n1453 VSS.t1163 70.0005
R3466 VSS.n1465 VSS.t1314 70.0005
R3467 VSS.n1478 VSS.t1250 70.0005
R3468 VSS.n1499 VSS.t1561 70.0005
R3469 VSS.n1502 VSS.t1961 70.0005
R3470 VSS.n1523 VSS.t1638 70.0005
R3471 VSS.t2031 VSS.t2844 69.7693
R3472 VSS.n1185 VSS.n1109 69.6809
R3473 VSS.n4658 VSS.t3283 69.6809
R3474 VSS.n1230 VSS.n955 68.5181
R3475 VSS.n1231 VSS.n1230 68.5181
R3476 VSS.n975 VSS.n956 68.5181
R3477 VSS.n1225 VSS.n956 68.5181
R3478 VSS.n1509 VSS.t1393 68.4925
R3479 VSS.n1509 VSS.t63 68.4925
R3480 VSS.n3995 VSS.t711 68.1564
R3481 VSS.n1527 VSS.t1370 68.1564
R3482 VSS.t89 VSS.n4631 67.9133
R3483 VSS.t753 VSS.t1839 67.4335
R3484 VSS.t1300 VSS.t496 67.4335
R3485 VSS.t868 VSS.t1146 67.4335
R3486 VSS.t1331 VSS.t745 67.4335
R3487 VSS.t1835 VSS.t1179 67.4335
R3488 VSS.t1528 VSS.t587 67.4335
R3489 VSS.t391 VSS.t756 67.4335
R3490 VSS.t399 VSS.t413 67.4335
R3491 VSS.t887 VSS.t1975 67.4335
R3492 VSS.t525 VSS.t107 67.4335
R3493 VSS.t2227 VSS.t1508 67.4335
R3494 VSS.t3157 VSS.t1747 67.4335
R3495 VSS.t3009 VSS.n1488 67.4335
R3496 VSS.t1311 VSS.t1651 67.4335
R3497 VSS.t1532 VSS.t1168 67.4335
R3498 VSS.t1162 VSS.t38 67.4335
R3499 VSS.t1981 VSS.t1009 67.4335
R3500 VSS.t909 VSS.t816 67.4335
R3501 VSS.t941 VSS.t2120 67.4335
R3502 VSS.n4646 VSS.n4645 67.2005
R3503 VSS.n4646 VSS.n465 67.2005
R3504 VSS.n4811 VSS.n465 67.2005
R3505 VSS.n4594 VSS.n466 67.2005
R3506 VSS.n4595 VSS.n4594 67.2005
R3507 VSS.n1213 VSS.n1212 67.2005
R3508 VSS.n1212 VSS.n989 67.2005
R3509 VSS.n1200 VSS.n1199 67.2005
R3510 VSS.n1199 VSS.n1198 67.2005
R3511 VSS.n1198 VSS.n1004 67.2005
R3512 VSS.n4810 VSS.n466 66.8805
R3513 VSS.n1001 VSS.n989 66.8805
R3514 VSS.n3328 VSS.n3327 66.462
R3515 VSS.t2685 VSS.n5349 66.251
R3516 VSS.n4654 VSS.n4653 65.0005
R3517 VSS.n4655 VSS.n4654 65.0005
R3518 VSS.n4634 VSS.n4633 65.0005
R3519 VSS.n4633 VSS.n4632 65.0005
R3520 VSS.n1188 VSS.n1187 65.0005
R3521 VSS.n1187 VSS.n1186 65.0005
R3522 VSS.n1183 VSS.n1182 65.0005
R3523 VSS.n1184 VSS.n1183 65.0005
R3524 VSS.n4029 VSS.n4028 64.6159
R3525 VSS.n1641 VSS.n1640 64.6159
R3526 VSS.n1068 VSS.n1037 64.5278
R3527 VSS.n4356 VSS.t2218 63.9215
R3528 VSS.n4356 VSS.t2089 63.9215
R3529 VSS.n4630 VSS.n4629 63.7794
R3530 VSS.n2905 VSS.n2904 63.5738
R3531 VSS.n3953 VSS.n3952 62.7697
R3532 VSS.n3572 VSS.n3571 62.7697
R3533 VSS.t2735 VSS.n1249 62.7648
R3534 VSS.t549 VSS.n462 62.7648
R3535 VSS.t2733 VSS.n1249 62.7648
R3536 VSS.t560 VSS.n462 62.7648
R3537 VSS.n4612 VSS.t2739 62.7647
R3538 VSS.n4612 VSS.t2737 62.7647
R3539 VSS.t2844 VSS.t2841 62.5968
R3540 VSS.t2839 VSS.t2840 62.5968
R3541 VSS.n3029 VSS.t588 61.6309
R3542 VSS.n3064 VSS.t1073 61.6309
R3543 VSS.n3071 VSS.t47 61.6309
R3544 VSS.n3129 VSS.t1041 61.6309
R3545 VSS.n2286 VSS.t2036 61.6309
R3546 VSS.n2739 VSS.t1151 61.6309
R3547 VSS.n2784 VSS.t1198 61.6309
R3548 VSS.n2810 VSS.t1811 61.6309
R3549 VSS.n1446 VSS.t2574 61.6309
R3550 VSS.n4386 VSS.t1475 61.4291
R3551 VSS.n3488 VSS.t1161 61.4291
R3552 VSS.n3496 VSS.t1569 61.4291
R3553 VSS.n3526 VSS.t1192 61.4291
R3554 VSS.n3553 VSS.t699 61.4291
R3555 VSS.n3645 VSS.t1186 61.4291
R3556 VSS.t822 VSS.t1116 61.0597
R3557 VSS.n3815 VSS.t697 60.5809
R3558 VSS.n4138 VSS.t2155 60.5809
R3559 VSS.n4145 VSS.t1628 60.5809
R3560 VSS.n4181 VSS.t1299 60.5809
R3561 VSS.n3732 VSS.t2143 60.5809
R3562 VSS.n3695 VSS.t1330 60.5809
R3563 VSS.n3667 VSS.t692 60.5809
R3564 VSS.n2958 VSS.t3000 60.5809
R3565 VSS.n2982 VSS.t1965 60.5809
R3566 VSS.n2999 VSS.t2117 60.5809
R3567 VSS.n3042 VSS.t1554 60.5809
R3568 VSS.n3120 VSS.t1494 60.5809
R3569 VSS.n2210 VSS.t1644 60.5809
R3570 VSS.n2300 VSS.t978 60.5809
R3571 VSS.n2662 VSS.t929 60.5809
R3572 VSS.n2047 VSS.t791 60.5809
R3573 VSS.n1346 VSS.t942 60.5809
R3574 VSS.n1970 VSS.t1218 60.5809
R3575 VSS.n1381 VSS.t793 60.5809
R3576 VSS.n1398 VSS.t913 60.5809
R3577 VSS.n1420 VSS.t1013 60.5809
R3578 VSS.n1449 VSS.t2149 60.5809
R3579 VSS.n1459 VSS.t795 60.5809
R3580 VSS.n1471 VSS.t1567 60.5809
R3581 VSS.n1721 VSS.t1487 60.5809
R3582 VSS.n1713 VSS.t1704 60.5809
R3583 VSS.n1519 VSS.t1940 60.5809
R3584 VSS.t2876 VSS.t989 60.4366
R3585 VSS.n4951 VSS.n4950 59.4829
R3586 VSS.n4952 VSS.n4951 59.4829
R3587 VSS.n4952 VSS.n355 59.4829
R3588 VSS.n4964 VSS.n355 59.4829
R3589 VSS.n4965 VSS.n4964 59.4829
R3590 VSS.n4966 VSS.n4965 59.4829
R3591 VSS.n1086 VSS.n1085 59.4829
R3592 VSS.n1087 VSS.n1086 59.4829
R3593 VSS.t931 VSS.t1026 59.1905
R3594 VSS.t953 VSS.t2567 59.1905
R3595 VSS.t2984 VSS.t768 59.1905
R3596 VSS.n4274 VSS.t1591 59.0774
R3597 VSS.t2104 VSS.t3039 59.0043
R3598 VSS.t1411 VSS.t800 59.0043
R3599 VSS.t2741 VSS.t1474 59.0043
R3600 VSS.t602 VSS.t2889 59.0043
R3601 VSS.t3417 VSS.t609 59.0043
R3602 VSS.t3027 VSS.t2852 59.0043
R3603 VSS.t2814 VSS.t698 59.0043
R3604 VSS.t179 VSS.t1185 59.0043
R3605 VSS.t1070 VSS.t2887 59.0043
R3606 VSS.t585 VSS.t1290 59.0043
R3607 VSS.t2015 VSS.t355 59.0043
R3608 VSS.n125 VSS.t2804 58.5719
R3609 VSS.n3091 VSS.t2904 58.5719
R3610 VSS.n3117 VSS.t575 58.5719
R3611 VSS.n2275 VSS.t1726 58.5719
R3612 VSS.n2299 VSS.t565 58.5719
R3613 VSS.n4632 VSS.t1114 57.9444
R3614 VSS.t774 VSS.t2979 57.3805
R3615 VSS.t2843 VSS.t2041 56.7284
R3616 VSS.n4274 VSS.t1661 56.3082
R3617 VSS.t693 VSS.t895 55.8706
R3618 VSS.n4505 VSS.t1381 55.7148
R3619 VSS.n4553 VSS.t2004 55.7148
R3620 VSS.n11 VSS.t860 55.7148
R3621 VSS.n22 VSS.t2052 55.7148
R3622 VSS.n38 VSS.t1420 55.7148
R3623 VSS.n47 VSS.t1901 55.7148
R3624 VSS.n64 VSS.t1234 55.7148
R3625 VSS.n84 VSS.t1057 55.7148
R3626 VSS.n4114 VSS.t2653 55.7148
R3627 VSS.n4176 VSS.t1212 55.7148
R3628 VSS.n1534 VSS.t139 55.7148
R3629 VSS.n5326 VSS.t2692 55.7148
R3630 VSS.n409 VSS.t990 55.7148
R3631 VSS.t2011 VSS.t2937 54.8292
R3632 VSS.t2810 VSS.t518 54.7723
R3633 VSS.n321 VSS.t2417 53.7941
R3634 VSS.t3241 VSS.t549 53.5831
R3635 VSS.t989 VSS.t983 53.5831
R3636 VSS.t987 VSS.t985 53.5831
R3637 VSS.n92 VSS.t1447 52.8576
R3638 VSS.n122 VSS.t479 52.8576
R3639 VSS.n146 VSS.t1173 52.8576
R3640 VSS.n160 VSS.t1097 52.8576
R3641 VSS.n3825 VSS.t2614 52.8576
R3642 VSS.n3990 VSS.t1731 52.8576
R3643 VSS.n3788 VSS.t1790 52.8576
R3644 VSS.n4115 VSS.t2191 52.8576
R3645 VSS.n4167 VSS.t1254 52.8576
R3646 VSS.n4249 VSS.t2147 52.8576
R3647 VSS.n3753 VSS.t1427 52.8576
R3648 VSS.n3709 VSS.t1147 52.8576
R3649 VSS.n3030 VSS.t1529 52.8576
R3650 VSS.n3017 VSS.t1587 52.8576
R3651 VSS.n3099 VSS.t37 52.8576
R3652 VSS.n2203 VSS.t153 52.8576
R3653 VSS.n2221 VSS.t584 52.8576
R3654 VSS.n2236 VSS.t2851 52.8576
R3655 VSS.n2280 VSS.t3008 52.8576
R3656 VSS.n2295 VSS.t1358 52.8576
R3657 VSS.n2193 VSS.t1589 52.8576
R3658 VSS.n2674 VSS.t1425 52.8576
R3659 VSS.n2763 VSS.t1463 52.8576
R3660 VSS.n1355 VSS.t1688 52.8576
R3661 VSS.n1433 VSS.t2215 52.8576
R3662 VSS.n4836 VSS.t823 52.8576
R3663 VSS.t1808 VSS.t822 52.3369
R3664 VSS.t890 VSS.t1808 52.3369
R3665 VSS.t933 VSS.t931 52.3369
R3666 VSS.t2624 VSS.t2622 52.3369
R3667 VSS.t768 VSS.t770 52.3369
R3668 VSS.t3281 VSS.n4658 51.9441
R3669 VSS.n4960 VSS.n350 51.7539
R3670 VSS.n4502 VSS.t461 51.4291
R3671 VSS.n4499 VSS.t321 51.4291
R3672 VSS.n176 VSS.t2846 51.4291
R3673 VSS.n5361 VSS.t2791 51.4291
R3674 VSS.n3845 VSS.t76 51.4291
R3675 VSS.n3848 VSS.t359 51.4291
R3676 VSS.n3850 VSS.t129 51.4291
R3677 VSS.n3875 VSS.t324 51.4291
R3678 VSS.n3876 VSS.t302 51.4291
R3679 VSS.n3783 VSS.t2711 51.4291
R3680 VSS.n4440 VSS.t2966 51.4291
R3681 VSS.n4441 VSS.t2560 51.4291
R3682 VSS.n4436 VSS.t524 51.4291
R3683 VSS.n4437 VSS.t106 51.4291
R3684 VSS.n4433 VSS.t2978 51.4291
R3685 VSS.n2946 VSS.t400 51.4291
R3686 VSS.n3020 VSS.t378 51.4291
R3687 VSS.n3049 VSS.t5 51.4291
R3688 VSS.n3158 VSS.t1322 51.4291
R3689 VSS.n3134 VSS.t2930 51.4291
R3690 VSS.n3137 VSS.t3012 51.4291
R3691 VSS.n3138 VSS.t675 51.4291
R3692 VSS.n2086 VSS.t431 51.4291
R3693 VSS.n2094 VSS.t354 51.4291
R3694 VSS.n2082 VSS.t2855 51.4291
R3695 VSS.n2083 VSS.t2785 51.4291
R3696 VSS.n2213 VSS.t217 51.4291
R3697 VSS.n2260 VSS.t2867 51.4291
R3698 VSS.n2267 VSS.t2193 51.4291
R3699 VSS.n2330 VSS.t1764 51.4291
R3700 VSS.n2333 VSS.t1934 51.4291
R3701 VSS.n2337 VSS.t598 51.4291
R3702 VSS.n2339 VSS.t930 51.4291
R3703 VSS.n2860 VSS.t906 51.4291
R3704 VSS.n2861 VSS.t2172 51.4291
R3705 VSS.n2868 VSS.t1492 51.4291
R3706 VSS.n2869 VSS.t2132 51.4291
R3707 VSS.n2647 VSS.t1509 51.4291
R3708 VSS.n2802 VSS.t2906 51.4291
R3709 VSS.n2806 VSS.t92 51.4291
R3710 VSS.n1475 VSS.t1265 51.4291
R3711 VSS.n1591 VSS.t1033 51.4291
R3712 VSS.n1548 VSS.t1348 51.4291
R3713 VSS.n1551 VSS.t752 51.4291
R3714 VSS.n1554 VSS.t1398 51.4291
R3715 VSS.n1557 VSS.t2164 51.4291
R3716 VSS.n1559 VSS.t992 51.4291
R3717 VSS.n1276 VSS.t2157 51.4291
R3718 VSS.n1277 VSS.t688 51.4291
R3719 VSS.n1272 VSS.t1206 51.4291
R3720 VSS.n1273 VSS.t1694 51.4291
R3721 VSS.n1269 VSS.t829 51.4291
R3722 VSS.n387 VSS.t1027 51.4291
R3723 VSS.n4879 VSS.t1324 51.4291
R3724 VSS.n4893 VSS.t2042 51.4291
R3725 VSS.n286 VSS.t1604 51.4291
R3726 VSS.n5048 VSS.t1469 51.4291
R3727 VSS.n257 VSS.t2134 51.4291
R3728 VSS.n245 VSS.t1571 51.4291
R3729 VSS.n5129 VSS.t1113 51.4291
R3730 VSS.n233 VSS.t1256 51.4291
R3731 VSS.n217 VSS.t900 51.4291
R3732 VSS.n202 VSS.t2562 51.4291
R3733 VSS.n5283 VSS.t1293 51.4291
R3734 VSS.n184 VSS.t2602 51.4291
R3735 VSS.n5311 VSS.t1540 51.4291
R3736 VSS.n5318 VSS.t1019 51.4291
R3737 VSS.n400 VSS.t954 51.4291
R3738 VSS.n403 VSS.t2639 51.4291
R3739 VSS.n406 VSS.t2985 51.4291
R3740 VSS.t193 VSS.n1195 51.2802
R3741 VSS.t1213 VSS.t1399 50.5752
R3742 VSS.t981 VSS.t1514 50.5752
R3743 VSS.t2247 VSS.t2763 50.5752
R3744 VSS.t998 VSS.t1830 50.5752
R3745 VSS.t2856 VSS.t1347 50.5752
R3746 VSS.t136 VSS.t547 50.5752
R3747 VSS.t563 VSS.t1132 50.5752
R3748 VSS.t3223 VSS.t1935 50.5752
R3749 VSS.t1005 VSS.t3491 50.5752
R3750 VSS.n4975 VSS.t65 50.3389
R3751 VSS.n348 VSS.t67 49.813
R3752 VSS.n305 VSS.n304 49.6897
R3753 VSS.n318 VSS.t2490 49.2941
R3754 VSS.n4959 VSS.n4958 48.7505
R3755 VSS.n4958 VSS.n4957 48.7505
R3756 VSS.n352 VSS.n349 48.7505
R3757 VSS.n4957 VSS.n352 48.7505
R3758 VSS.n1073 VSS.n1068 48.5434
R3759 VSS.t1699 VSS.t2838 48.2518
R3760 VSS.n1115 VSS.t2972 47.7249
R3761 VSS.n917 VSS.t23 47.7249
R3762 VSS.n1030 VSS.t1912 47.2331
R3763 VSS.n1029 VSS.t1919 47.2331
R3764 VSS.n1028 VSS.t1914 47.2331
R3765 VSS.n1121 VSS.t2836 47.1624
R3766 VSS.n1118 VSS.t2781 47.1624
R3767 VSS.n1117 VSS.t3003 47.1624
R3768 VSS.n1116 VSS.t2967 47.1624
R3769 VSS.n1115 VSS.t2832 47.1624
R3770 VSS.n923 VSS.t2898 47.1624
R3771 VSS.n920 VSS.t147 47.1624
R3772 VSS.n919 VSS.t127 47.1624
R3773 VSS.n918 VSS.t2085 47.1624
R3774 VSS.n917 VSS.t365 47.1624
R3775 VSS.n4800 VSS.t2953 47.1602
R3776 VSS.n1170 VSS.t2941 47.1602
R3777 VSS.n4946 VSS.n349 46.6799
R3778 VSS.n4275 VSS.n4274 46.2505
R3779 VSS.n4983 VSS.n4982 46.1526
R3780 VSS.n4628 VSS.t3469 46.0361
R3781 VSS.n4945 VSS.n4944 45.7304
R3782 VSS.n3985 VSS.t481 45.7148
R3783 VSS.t2979 VSS.t2839 44.9916
R3784 VSS.t2622 VSS.t2984 44.2373
R3785 VSS.n3930 VSS.t2105 44.0005
R3786 VSS.n3787 VSS.t1815 44.0005
R3787 VSS.n3016 VSS.t2161 44.0005
R3788 VSS.n2621 VSS.t2621 44.0005
R3789 VSS.n2584 VSS.t1777 44.0005
R3790 VSS.n2235 VSS.t1909 44.0005
R3791 VSS.n2277 VSS.t1755 44.0005
R3792 VSS.n2678 VSS.t718 44.0005
R3793 VSS.n2174 VSS.t1153 44.0005
R3794 VSS.n1352 VSS.t2058 44.0005
R3795 VSS.n377 VSS.t1115 44.0005
R3796 VSS.n1033 VSS.n1025 43.6225
R3797 VSS.n320 VSS.n319 43.373
R3798 VSS.n1026 VSS.t1917 42.7588
R3799 VSS.n1027 VSS.t1922 42.7178
R3800 VSS.n1027 VSS.t1921 42.6544
R3801 VSS.n1026 VSS.t1916 42.6361
R3802 VSS.t3485 VSS.t612 42.1461
R3803 VSS.t1409 VSS.t3100 42.1461
R3804 VSS.t46 VSS.t2955 42.1461
R3805 VSS.t56 VSS.t2123 42.1461
R3806 VSS.t1908 VSS.t2721 42.1461
R3807 VSS.t2643 VSS.t847 42.1461
R3808 VSS.t3136 VSS.t2265 42.1461
R3809 VSS.t1369 VSS.t1133 42.1461
R3810 VSS.t1672 VSS.t189 42.1461
R3811 VSS.n4982 VSS.n310 42.0061
R3812 VSS.n1253 VSS.n1252 41.7862
R3813 VSS.n1258 VSS.n1255 41.7862
R3814 VSS.n1257 VSS.n1256 41.7862
R3815 VSS.n4621 VSS.n1250 41.7862
R3816 VSS.n1250 VSS.n1248 41.7862
R3817 VSS.n1208 VSS.n1207 41.7862
R3818 VSS.n1209 VSS.n1208 41.7862
R3819 VSS.n1003 VSS.n1002 41.7862
R3820 VSS.n1006 VSS.n1005 41.7862
R3821 VSS.n1194 VSS.n1005 41.7862
R3822 VSS.n990 VSS.n988 41.7862
R3823 VSS.n992 VSS.n990 41.7862
R3824 VSS.n3995 VSS.t773 41.6479
R3825 VSS.n1527 VSS.t1783 41.6479
R3826 VSS.n4029 VSS.t1412 41.539
R3827 VSS.n3953 VSS.t1950 41.539
R3828 VSS.n3952 VSS.t1948 41.539
R3829 VSS.n3572 VSS.t2097 41.539
R3830 VSS.n3571 VSS.t1573 41.539
R3831 VSS.n1640 VSS.t1785 41.539
R3832 VSS.n961 VSS.n960 41.3146
R3833 VSS.n4596 VSS.n4595 40.7382
R3834 VSS.n1214 VSS.n1213 40.7382
R3835 VSS.n4028 VSS.t1337 40.6159
R3836 VSS.n3327 VSS.t655 40.6159
R3837 VSS.n3328 VSS.t1876 40.6159
R3838 VSS.n1641 VSS.t268 40.6159
R3839 VSS.n4519 VSS.t1387 40.0005
R3840 VSS.n4519 VSS.t1383 40.0005
R3841 VSS.n4505 VSS.t2094 40.0005
R3842 VSS.n4550 VSS.t1998 40.0005
R3843 VSS.n4550 VSS.t2002 40.0005
R3844 VSS.n4553 VSS.t952 40.0005
R3845 VSS.n10 VSS.t858 40.0005
R3846 VSS.n10 VSS.t862 40.0005
R3847 VSS.n11 VSS.t2010 40.0005
R3848 VSS.n22 VSS.t1395 40.0005
R3849 VSS.n25 VSS.t2050 40.0005
R3850 VSS.n25 VSS.t2046 40.0005
R3851 VSS.n38 VSS.t1582 40.0005
R3852 VSS.n41 VSS.t1422 40.0005
R3853 VSS.n41 VSS.t1418 40.0005
R3854 VSS.n47 VSS.t956 40.0005
R3855 VSS.n50 VSS.t1899 40.0005
R3856 VSS.n50 VSS.t1903 40.0005
R3857 VSS.n64 VSS.t1616 40.0005
R3858 VSS.n65 VSS.t1230 40.0005
R3859 VSS.n65 VSS.t1232 40.0005
R3860 VSS.n81 VSS.t1059 40.0005
R3861 VSS.n81 VSS.t1055 40.0005
R3862 VSS.n84 VSS.t3005 40.0005
R3863 VSS.n92 VSS.t1443 40.0005
R3864 VSS.n146 VSS.t143 40.0005
R3865 VSS.n160 VSS.t145 40.0005
R3866 VSS.n4114 VSS.t86 40.0005
R3867 VSS.n4115 VSS.t1109 40.0005
R3868 VSS.n3778 VSS.t2657 40.0005
R3869 VSS.n3778 VSS.t2655 40.0005
R3870 VSS.n4167 VSS.t2030 40.0005
R3871 VSS.n4176 VSS.t51 40.0005
R3872 VSS.n4178 VSS.t1208 40.0005
R3873 VSS.n4178 VSS.t1214 40.0005
R3874 VSS.n4249 VSS.t206 40.0005
R3875 VSS.n3709 VSS.t2091 40.0005
R3876 VSS.n3030 VSS.t215 40.0005
R3877 VSS.n2295 VSS.t1108 40.0005
R3878 VSS.n1433 VSS.t82 40.0005
R3879 VSS.n1534 VSS.t59 40.0005
R3880 VSS.n1535 VSS.t135 40.0005
R3881 VSS.n1535 VSS.t137 40.0005
R3882 VSS.n5326 VSS.t1500 40.0005
R3883 VSS.n5327 VSS.t2688 40.0005
R3884 VSS.n5327 VSS.t2686 40.0005
R3885 VSS.n409 VSS.t2877 40.0005
R3886 VSS.n412 VSS.t984 40.0005
R3887 VSS.n412 VSS.t988 40.0005
R3888 VSS.n1236 VSS.n1235 39.2749
R3889 VSS.n1016 VSS.n1014 39.0005
R3890 VSS.n1106 VSS.n1016 39.0005
R3891 VSS.n4622 VSS.n1242 39.0005
R3892 VSS.n1244 VSS.n1243 39.0005
R3893 VSS.n1247 VSS.n1244 39.0005
R3894 VSS.n1104 VSS.n1103 39.0005
R3895 VSS.t1918 VSS.n1104 39.0005
R3896 VSS.n1100 VSS.n1020 39.0005
R3897 VSS.t1918 VSS.n1020 39.0005
R3898 VSS.n1241 VSS.n1239 39.0005
R3899 VSS.n4625 VSS.n1239 39.0005
R3900 VSS.n1192 VSS.n1191 39.0005
R3901 VSS.n1193 VSS.n1192 39.0005
R3902 VSS.n1111 VSS.n1013 39.0005
R3903 VSS.n4001 VSS.t1659 38.7697
R3904 VSS.n3747 VSS.t390 38.7697
R3905 VSS.n3747 VSS.t1819 38.7697
R3906 VSS.n3739 VSS.t810 38.7697
R3907 VSS.n2243 VSS.t2635 38.7697
R3908 VSS.n2246 VSS.t1088 38.7697
R3909 VSS.n2518 VSS.t1887 38.7697
R3910 VSS.n2659 VSS.t1565 38.7697
R3911 VSS.n119 VSS.t606 38.5719
R3912 VSS.n119 VSS.t112 38.5719
R3913 VSS.n4385 VSS.t1471 38.5719
R3914 VSS.n3942 VSS.t1437 38.5719
R3915 VSS.n3942 VSS.t1838 38.5719
R3916 VSS.n3920 VSS.t1091 38.5719
R3917 VSS.n3920 VSS.t1043 38.5719
R3918 VSS.n3930 VSS.t652 38.5719
R3919 VSS.n3985 VSS.t578 38.5719
R3920 VSS.n3989 VSS.t1188 38.5719
R3921 VSS.n3989 VSS.t590 38.5719
R3922 VSS.n3801 VSS.t13 38.5719
R3923 VSS.n3801 VSS.t219 38.5719
R3924 VSS.n3791 VSS.t2861 38.5719
R3925 VSS.n3791 VSS.t2724 38.5719
R3926 VSS.n3793 VSS.t789 38.5719
R3927 VSS.n3793 VSS.t45 38.5719
R3928 VSS.n3787 VSS.t2718 38.5719
R3929 VSS.n3784 VSS.t1870 38.5719
R3930 VSS.n3784 VSS.t159 38.5719
R3931 VSS.n3775 VSS.t41 38.5719
R3932 VSS.n3775 VSS.t2169 38.5719
R3933 VSS.n3763 VSS.t2252 38.5719
R3934 VSS.n3763 VSS.t35 38.5719
R3935 VSS.n4189 VSS.t1276 38.5719
R3936 VSS.n4189 VSS.t422 38.5719
R3937 VSS.n3752 VSS.t2073 38.5719
R3938 VSS.n3752 VSS.t974 38.5719
R3939 VSS.n3725 VSS.t1679 38.5719
R3940 VSS.n3725 VSS.t418 38.5719
R3941 VSS.n4422 VSS.t1642 38.5719
R3942 VSS.n4422 VSS.t430 38.5719
R3943 VSS.n3112 VSS.t1141 38.5719
R3944 VSS.n3112 VSS.t43 38.5719
R3945 VSS.n3446 VSS.t2579 38.5719
R3946 VSS.n3446 VSS.t29 38.5719
R3947 VSS.n3489 VSS.t1558 38.5719
R3948 VSS.n3497 VSS.t750 38.5719
R3949 VSS.n3527 VSS.t2756 38.5719
R3950 VSS.n3552 VSS.t2762 38.5719
R3951 VSS.n2971 VSS.t1595 38.5719
R3952 VSS.n2970 VSS.t2748 38.5719
R3953 VSS.n3644 VSS.t1023 38.5719
R3954 VSS.n2132 VSS.t1039 38.5719
R3955 VSS.n2132 VSS.t412 38.5719
R3956 VSS.n2947 VSS.t757 38.5719
R3957 VSS.n2947 VSS.t414 38.5719
R3958 VSS.n2950 VSS.t1878 38.5719
R3959 VSS.n2950 VSS.t392 38.5719
R3960 VSS.n2974 VSS.t2151 38.5719
R3961 VSS.n2974 VSS.t416 38.5719
R3962 VSS.n3007 VSS.t208 38.5719
R3963 VSS.n3007 VSS.t2273 38.5719
R3964 VSS.n3016 VSS.t2594 38.5719
R3965 VSS.n3022 VSS.t2600 38.5719
R3966 VSS.n3022 VSS.t2264 38.5719
R3967 VSS.n3023 VSS.t1316 38.5719
R3968 VSS.n3023 VSS.t2912 38.5719
R3969 VSS.n3050 VSS.t1180 38.5719
R3970 VSS.n3050 VSS.t155 38.5719
R3971 VSS.n3382 VSS.t2910 38.5719
R3972 VSS.n3382 VSS.t402 38.5719
R3973 VSS.n3072 VSS.t1826 38.5719
R3974 VSS.n3072 VSS.t2956 38.5719
R3975 VSS.n3102 VSS.t384 38.5719
R3976 VSS.n3102 VSS.t1374 38.5719
R3977 VSS.n2621 VSS.t2915 38.5719
R3978 VSS.n2207 VSS.t848 38.5719
R3979 VSS.n2207 VSS.t586 38.5719
R3980 VSS.n2216 VSS.t1015 38.5719
R3981 VSS.n2216 VSS.t161 38.5719
R3982 VSS.n2218 VSS.t27 38.5719
R3983 VSS.n2218 VSS.t2642 38.5719
R3984 VSS.n2584 VSS.t230 38.5719
R3985 VSS.n2573 VSS.t767 38.5719
R3986 VSS.n2573 VSS.t2572 38.5719
R3987 VSS.n2235 VSS.t7 38.5719
R3988 VSS.n2239 VSS.t846 38.5719
R3989 VSS.n2239 VSS.t1071 38.5719
R3990 VSS.n2262 VSS.t761 38.5719
R3991 VSS.n2262 VSS.t163 38.5719
R3992 VSS.n2277 VSS.t2884 38.5719
R3993 VSS.n2283 VSS.t2054 38.5719
R3994 VSS.n2283 VSS.t2038 38.5719
R3995 VSS.n2292 VSS.t701 38.5719
R3996 VSS.n2292 VSS.t1433 38.5719
R3997 VSS.n2669 VSS.t1606 38.5719
R3998 VSS.n2669 VSS.t211 38.5719
R3999 VSS.n2197 VSS.t2266 38.5719
R4000 VSS.n2197 VSS.t2597 38.5719
R4001 VSS.n2188 VSS.t386 38.5719
R4002 VSS.n2188 VSS.t808 38.5719
R4003 VSS.n2670 VSS.t916 38.5719
R4004 VSS.n2670 VSS.t976 38.5719
R4005 VSS.n2678 VSS.t2071 38.5719
R4006 VSS.n2174 VSS.t2732 38.5719
R4007 VSS.n2177 VSS.t690 38.5719
R4008 VSS.n2177 VSS.t1149 38.5719
R4009 VSS.n2800 VSS.t1221 38.5719
R4010 VSS.n2800 VSS.t394 38.5719
R4011 VSS.n2805 VSS.t1178 38.5719
R4012 VSS.n2805 VSS.t382 38.5719
R4013 VSS.n1367 VSS.t2100 38.5719
R4014 VSS.n1367 VSS.t426 38.5719
R4015 VSS.n1331 VSS.t2260 38.5719
R4016 VSS.n1331 VSS.t428 38.5719
R4017 VSS.n1336 VSS.t908 38.5719
R4018 VSS.n1336 VSS.t420 38.5719
R4019 VSS.n1352 VSS.t408 38.5719
R4020 VSS.n1357 VSS.t2176 38.5719
R4021 VSS.n1357 VSS.t1196 38.5719
R4022 VSS.n1969 VSS.t2109 38.5719
R4023 VSS.n1969 VSS.t424 38.5719
R4024 VSS.n1389 VSS.t1004 38.5719
R4025 VSS.n1389 VSS.t213 38.5719
R4026 VSS.n1412 VSS.t1010 38.5719
R4027 VSS.n1412 VSS.t204 38.5719
R4028 VSS.n1441 VSS.t2180 38.5719
R4029 VSS.n1441 VSS.t31 38.5719
R4030 VSS.n1452 VSS.t1675 38.5719
R4031 VSS.n1452 VSS.t39 38.5719
R4032 VSS.n1464 VSS.t1158 38.5719
R4033 VSS.n1464 VSS.t33 38.5719
R4034 VSS.n1489 VSS.t1930 38.5719
R4035 VSS.n1489 VSS.t1431 38.5719
R4036 VSS.n1492 VSS.t1441 38.5719
R4037 VSS.n1492 VSS.t1435 38.5719
R4038 VSS.n1513 VSS.t1936 38.5719
R4039 VSS.n1513 VSS.t1429 38.5719
R4040 VSS.n4835 VSS.t1809 38.5719
R4041 VSS.n4835 VSS.t891 38.5719
R4042 VSS.n377 VSS.t90 38.5719
R4043 VSS.n4642 VSS.n4641 37.7605
R4044 VSS.n1181 VSS.n1114 37.7605
R4045 VSS.n1120 VSS.n1119 37.2624
R4046 VSS.n922 VSS.n921 37.2624
R4047 VSS.t1116 VSS.t3054 36.1376
R4048 VSS.n3998 VSS.t1119 36.0005
R4049 VSS.n3998 VSS.t1928 36.0005
R4050 VSS.n2955 VSS.t2728 36.0005
R4051 VSS.n2955 VSS.t2679 36.0005
R4052 VSS.n3082 VSS.t1693 36.0005
R4053 VSS.n3094 VSS.t1051 36.0005
R4054 VSS.n3094 VSS.t476 36.0005
R4055 VSS.n2289 VSS.t1856 36.0005
R4056 VSS.n1053 VSS.t2031 35.863
R4057 VSS.n3594 VSS.n3591 35.4914
R4058 VSS.n4666 VSS.n937 35.0505
R4059 VSS.n1157 VSS.n1156 35.0505
R4060 VSS.n3029 VSS.t2924 34.8099
R4061 VSS.n3064 VSS.t3 34.8099
R4062 VSS.n3071 VSS.t2708 34.8099
R4063 VSS.n3129 VSS.t681 34.8099
R4064 VSS.n2286 VSS.t2886 34.8099
R4065 VSS.n2739 VSS.t2730 34.8099
R4066 VSS.n2784 VSS.t396 34.8099
R4067 VSS.n2810 VSS.t94 34.8099
R4068 VSS.n1446 VSS.t228 34.8099
R4069 VSS.n4010 VSS.n4009 34.6358
R4070 VSS.n4364 VSS.n3712 34.6358
R4071 VSS.n335 VSS.n329 34.6358
R4072 VSS.n336 VSS.n335 34.6358
R4073 VSS.n4538 VSS.n4537 34.6358
R4074 VSS.n4545 VSS.n4544 34.6358
R4075 VSS.n4544 VSS.n4497 34.6358
R4076 VSS.n5681 VSS.n5680 34.6358
R4077 VSS.n5648 VSS.n5647 34.6358
R4078 VSS.n5597 VSS.n85 34.6358
R4079 VSS.n5601 VSS.n85 34.6358
R4080 VSS.n5594 VSS.n88 34.6358
R4081 VSS.n5595 VSS.n5594 34.6358
R4082 VSS.n5579 VSS.n93 34.6358
R4083 VSS.n5555 VSS.n5554 34.6358
R4084 VSS.n5513 VSS.n5512 34.6358
R4085 VSS.n5499 VSS.n5498 34.6358
R4086 VSS.n5500 VSS.n5499 34.6358
R4087 VSS.n5493 VSS.n5492 34.6358
R4088 VSS.n5494 VSS.n5493 34.6358
R4089 VSS.n5390 VSS.n171 34.6358
R4090 VSS.n5394 VSS.n171 34.6358
R4091 VSS.n5388 VSS.n174 34.6358
R4092 VSS.n5376 VSS.n5359 34.6358
R4093 VSS.n3960 VSS.n3959 34.6358
R4094 VSS.n3963 VSS.n3812 34.6358
R4095 VSS.n3971 VSS.n3968 34.6358
R4096 VSS.n3975 VSS.n3810 34.6358
R4097 VSS.n3976 VSS.n3975 34.6358
R4098 VSS.n4015 VSS.n4014 34.6358
R4099 VSS.n4014 VSS.n4013 34.6358
R4100 VSS.n4058 VSS.n3804 34.6358
R4101 VSS.n4062 VSS.n3804 34.6358
R4102 VSS.n4069 VSS.n3802 34.6358
R4103 VSS.n4094 VSS.n4093 34.6358
R4104 VSS.n4124 VSS.n3774 34.6358
R4105 VSS.n4136 VSS.n3771 34.6358
R4106 VSS.n4137 VSS.n4136 34.6358
R4107 VSS.n4140 VSS.n4137 34.6358
R4108 VSS.n4144 VSS.n3769 34.6358
R4109 VSS.n4148 VSS.n4147 34.6358
R4110 VSS.n4148 VSS.n3767 34.6358
R4111 VSS.n4152 VSS.n3767 34.6358
R4112 VSS.n4231 VSS.n4230 34.6358
R4113 VSS.n4213 VSS.n4179 34.6358
R4114 VSS.n4208 VSS.n4207 34.6358
R4115 VSS.n4204 VSS.n4203 34.6358
R4116 VSS.n4201 VSS.n4185 34.6358
R4117 VSS.n4197 VSS.n4185 34.6358
R4118 VSS.n4197 VSS.n4196 34.6358
R4119 VSS.n4287 VSS.n4286 34.6358
R4120 VSS.n4353 VSS.n3716 34.6358
R4121 VSS.n4360 VSS.n4355 34.6358
R4122 VSS.n4365 VSS.n4364 34.6358
R4123 VSS.n4367 VSS.n3708 34.6358
R4124 VSS.n4389 VSS.n3698 34.6358
R4125 VSS.n4402 VSS.n3698 34.6358
R4126 VSS.n4409 VSS.n4408 34.6358
R4127 VSS.n4412 VSS.n3693 34.6358
R4128 VSS.n4416 VSS.n3693 34.6358
R4129 VSS.n3688 VSS.n2130 34.6358
R4130 VSS.n3676 VSS.n3675 34.6358
R4131 VSS.n3676 VSS.n2135 34.6358
R4132 VSS.n3680 VSS.n2135 34.6358
R4133 VSS.n3673 VSS.n2138 34.6358
R4134 VSS.n3649 VSS.n2142 34.6358
R4135 VSS.n3665 VSS.n2142 34.6358
R4136 VSS.n3627 VSS.n3626 34.6358
R4137 VSS.n3614 VSS.n2959 34.6358
R4138 VSS.n3570 VSS.n3569 34.6358
R4139 VSS.n3557 VSS.n2985 34.6358
R4140 VSS.n3561 VSS.n2985 34.6358
R4141 VSS.n3533 VSS.n3532 34.6358
R4142 VSS.n3534 VSS.n3533 34.6358
R4143 VSS.n3519 VSS.n3518 34.6358
R4144 VSS.n3519 VSS.n3000 34.6358
R4145 VSS.n3523 VSS.n3000 34.6358
R4146 VSS.n3516 VSS.n3003 34.6358
R4147 VSS.n3512 VSS.n3510 34.6358
R4148 VSS.n3505 VSS.n3504 34.6358
R4149 VSS.n3495 VSS.n3494 34.6358
R4150 VSS.n3486 VSS.n3485 34.6358
R4151 VSS.n3478 VSS.n3025 34.6358
R4152 VSS.n3461 VSS.n3031 34.6358
R4153 VSS.n3442 VSS.n3037 34.6358
R4154 VSS.n3435 VSS.n3434 34.6358
R4155 VSS.n3438 VSS.n3435 34.6358
R4156 VSS.n3424 VSS.n3043 34.6358
R4157 VSS.n3428 VSS.n3043 34.6358
R4158 VSS.n3429 VSS.n3428 34.6358
R4159 VSS.n3418 VSS.n3047 34.6358
R4160 VSS.n3422 VSS.n3047 34.6358
R4161 VSS.n3400 VSS.n3060 34.6358
R4162 VSS.n3384 VSS.n3381 34.6358
R4163 VSS.n3376 VSS.n3067 34.6358
R4164 VSS.n3380 VSS.n3067 34.6358
R4165 VSS.n3381 VSS.n3380 34.6358
R4166 VSS.n3338 VSS.n3086 34.6358
R4167 VSS.n3311 VSS.n3310 34.6358
R4168 VSS.n3263 VSS.n3262 34.6358
R4169 VSS.n3264 VSS.n3263 34.6358
R4170 VSS.n3248 VSS.n3125 34.6358
R4171 VSS.n3249 VSS.n3248 34.6358
R4172 VSS.n2623 VSS.n2620 34.6358
R4173 VSS.n2598 VSS.n2597 34.6358
R4174 VSS.n2599 VSS.n2598 34.6358
R4175 VSS.n2549 VSS.n2237 34.6358
R4176 VSS.n2538 VSS.n2537 34.6358
R4177 VSS.n2539 VSS.n2538 34.6358
R4178 VSS.n2539 VSS.n2241 34.6358
R4179 VSS.n2543 VSS.n2241 34.6358
R4180 VSS.n2503 VSS.n2255 34.6358
R4181 VSS.n2507 VSS.n2255 34.6358
R4182 VSS.n2483 VSS.n2273 34.6358
R4183 VSS.n2470 VSS.n2281 34.6358
R4184 VSS.n2473 VSS.n2472 34.6358
R4185 VSS.n2477 VSS.n2476 34.6358
R4186 VSS.n2451 VSS.n2450 34.6358
R4187 VSS.n2444 VSS.n2297 34.6358
R4188 VSS.n2439 VSS.n2438 34.6358
R4189 VSS.n2654 VSS.n2653 34.6358
R4190 VSS.n2728 VSS.n2727 34.6358
R4191 VSS.n2727 VSS.n2663 34.6358
R4192 VSS.n2723 VSS.n2663 34.6358
R4193 VSS.n2723 VSS.n2722 34.6358
R4194 VSS.n2696 VSS.n2680 34.6358
R4195 VSS.n2691 VSS.n2690 34.6358
R4196 VSS.n2690 VSS.n2684 34.6358
R4197 VSS.n2686 VSS.n2684 34.6358
R4198 VSS.n2790 VSS.n2786 34.6358
R4199 VSS.n2794 VSS.n2168 34.6358
R4200 VSS.n2795 VSS.n2794 34.6358
R4201 VSS.n2824 VSS.n2808 34.6358
R4202 VSS.n2820 VSS.n2808 34.6358
R4203 VSS.n2814 VSS.n2813 34.6358
R4204 VSS.n2813 VSS.n2154 34.6358
R4205 VSS.n2927 VSS.n2154 34.6358
R4206 VSS.n2053 VSS.n2052 34.6358
R4207 VSS.n2031 VSS.n1339 34.6358
R4208 VSS.n2045 VSS.n1339 34.6358
R4209 VSS.n2046 VSS.n2045 34.6358
R4210 VSS.n2049 VSS.n2046 34.6358
R4211 VSS.n2029 VSS.n1347 34.6358
R4212 VSS.n2020 VSS.n2019 34.6358
R4213 VSS.n2016 VSS.n2015 34.6358
R4214 VSS.n1979 VSS.n1371 34.6358
R4215 VSS.n1983 VSS.n1371 34.6358
R4216 VSS.n1977 VSS.n1374 34.6358
R4217 VSS.n1973 VSS.n1968 34.6358
R4218 VSS.n1966 VSS.n1377 34.6358
R4219 VSS.n1959 VSS.n1958 34.6358
R4220 VSS.n1962 VSS.n1959 34.6358
R4221 VSS.n1947 VSS.n1945 34.6358
R4222 VSS.n1951 VSS.n1383 34.6358
R4223 VSS.n1939 VSS.n1387 34.6358
R4224 VSS.n1943 VSS.n1387 34.6358
R4225 VSS.n1900 VSS.n1407 34.6358
R4226 VSS.n1878 VSS.n1417 34.6358
R4227 VSS.n1882 VSS.n1417 34.6358
R4228 VSS.n1859 VSS.n1858 34.6358
R4229 VSS.n1850 VSS.n1849 34.6358
R4230 VSS.n1842 VSS.n1439 34.6358
R4231 VSS.n1835 VSS.n1834 34.6358
R4232 VSS.n1838 VSS.n1835 34.6358
R4233 VSS.n1824 VSS.n1444 34.6358
R4234 VSS.n1828 VSS.n1444 34.6358
R4235 VSS.n1812 VSS.n1450 34.6358
R4236 VSS.n1816 VSS.n1450 34.6358
R4237 VSS.n1817 VSS.n1816 34.6358
R4238 VSS.n1798 VSS.n1797 34.6358
R4239 VSS.n1802 VSS.n1801 34.6358
R4240 VSS.n1792 VSS.n1791 34.6358
R4241 VSS.n1780 VSS.n1779 34.6358
R4242 VSS.n1784 VSS.n1783 34.6358
R4243 VSS.n1785 VSS.n1784 34.6358
R4244 VSS.n1760 VSS.n1758 34.6358
R4245 VSS.n1764 VSS.n1479 34.6358
R4246 VSS.n1765 VSS.n1764 34.6358
R4247 VSS.n1751 VSS.n1486 34.6358
R4248 VSS.n1752 VSS.n1751 34.6358
R4249 VSS.n1753 VSS.n1752 34.6358
R4250 VSS.n1737 VSS.n1736 34.6358
R4251 VSS.n1727 VSS.n1495 34.6358
R4252 VSS.n1719 VSS.n1497 34.6358
R4253 VSS.n1720 VSS.n1719 34.6358
R4254 VSS.n1723 VSS.n1720 34.6358
R4255 VSS.n1706 VSS.n1500 34.6358
R4256 VSS.n1710 VSS.n1500 34.6358
R4257 VSS.n1711 VSS.n1710 34.6358
R4258 VSS.n1692 VSS.n1507 34.6358
R4259 VSS.n1658 VSS.n1520 34.6358
R4260 VSS.n1662 VSS.n1520 34.6358
R4261 VSS.n1653 VSS.n1652 34.6358
R4262 VSS.n1649 VSS.n1528 34.6358
R4263 VSS.n1625 VSS.n1532 34.6358
R4264 VSS.n4834 VSS.n4833 34.6358
R4265 VSS.n4857 VSS.n378 34.6358
R4266 VSS.n4846 VSS.n4845 34.6358
R4267 VSS.n4924 VSS.n4882 34.6358
R4268 VSS.n4928 VSS.n4882 34.6358
R4269 VSS.n4918 VSS.n4917 34.6358
R4270 VSS.n4918 VSS.n4885 34.6358
R4271 VSS.n4922 VSS.n4885 34.6358
R4272 VSS.n4915 VSS.n4888 34.6358
R4273 VSS.n4908 VSS.n4891 34.6358
R4274 VSS.n4897 VSS.n295 34.6358
R4275 VSS.n5001 VSS.n293 34.6358
R4276 VSS.n5012 VSS.n285 34.6358
R4277 VSS.n5071 VSS.n256 34.6358
R4278 VSS.n5082 VSS.n5081 34.6358
R4279 VSS.n5089 VSS.n5088 34.6358
R4280 VSS.n5088 VSS.n5087 34.6358
R4281 VSS.n5087 VSS.n252 34.6358
R4282 VSS.n5095 VSS.n5094 34.6358
R4283 VSS.n5094 VSS.n5093 34.6358
R4284 VSS.n5101 VSS.n244 34.6358
R4285 VSS.n5172 VSS.n5171 34.6358
R4286 VSS.n5194 VSS.n225 34.6358
R4287 VSS.n5229 VSS.n5228 34.6358
R4288 VSS.n5254 VSS.n204 34.6358
R4289 VSS.n5250 VSS.n204 34.6358
R4290 VSS.n5250 VSS.n5249 34.6358
R4291 VSS.n5258 VSS.n201 34.6358
R4292 VSS.n5258 VSS.n5257 34.6358
R4293 VSS.n5270 VSS.n195 34.6358
R4294 VSS.n5270 VSS.n5269 34.6358
R4295 VSS.n5300 VSS.n5299 34.6358
R4296 VSS.n5310 VSS.n182 34.6358
R4297 VSS.n5306 VSS.n182 34.6358
R4298 VSS.n5346 VSS.n5324 34.6358
R4299 VSS.n448 VSS.n447 34.6358
R4300 VSS.n3618 VSS.n2959 34.3716
R4301 VSS.n54 VSS.t3647 34.2973
R4302 VSS.n132 VSS.t3631 34.2973
R4303 VSS.n3796 VSS.t3567 34.2973
R4304 VSS.n3822 VSS.t3787 34.2973
R4305 VSS.n3098 VSS.t3756 34.2973
R4306 VSS.n3359 VSS.t3727 34.2973
R4307 VSS.n2963 VSS.t3642 34.2973
R4308 VSS.n2888 VSS.t3739 34.2973
R4309 VSS.n2196 VSS.t3655 34.2973
R4310 VSS.n1919 VSS.t3588 34.2973
R4311 VSS.n3485 VSS.n3018 34.2593
R4312 VSS.n2620 VSS.n2619 34.2593
R4313 VSS.n2551 VSS.n2550 34.2593
R4314 VSS.n2472 VSS.n2471 34.2593
R4315 VSS.n2010 VSS.n2009 34.2593
R4316 VSS.n1853 VSS.n1430 34.2593
R4317 VSS.n4837 VSS.n378 34.2593
R4318 VSS.n1054 VSS.t295 33.9068
R4319 VSS.n4007 VSS.n4004 33.8829
R4320 VSS.n4100 VSS.n4099 33.8829
R4321 VSS.n4367 VSS.n4366 33.8829
R4322 VSS.n3510 VSS.n3509 33.8829
R4323 VSS.n3505 VSS.n3008 33.8829
R4324 VSS.n3434 VSS.n3040 33.8829
R4325 VSS.n3150 VSS.n3149 33.8829
R4326 VSS.n2476 VSS.n2278 33.8829
R4327 VSS.n2349 VSS.n2348 33.8829
R4328 VSS.n2698 VSS.n2697 33.8829
R4329 VSS.n2015 VSS.n2014 33.8829
R4330 VSS.n1812 VSS.n1811 33.8829
R4331 VSS.n1569 VSS.n1568 33.8829
R4332 VSS.n1295 VSS.n1294 33.8829
R4333 VSS.n4859 VSS.n4858 33.8829
R4334 VSS.t2188 VSS.t2656 33.717
R4335 VSS.t1176 VSS.t337 33.717
R4336 VSS.t628 VSS.t1951 33.717
R4337 VSS.t2017 VSS.t2607 33.717
R4338 VSS.t1277 VSS.t1209 33.717
R4339 VSS.t1072 VSS.t2909 33.717
R4340 VSS.t2272 VSS.t1710 33.717
R4341 VSS.t1432 VSS.t1855 33.717
R4342 VSS.t2053 VSS.t3010 33.717
R4343 VSS.t2037 VSS.t3006 33.717
R4344 VSS.t3007 VSS.t1266 33.717
R4345 VSS.t638 VSS.t15 33.717
R4346 VSS.t2872 VSS.t99 33.717
R4347 VSS.t409 VSS.t393 33.717
R4348 VSS.t138 VSS.t529 33.717
R4349 VSS.t595 VSS.t3494 33.717
R4350 VSS.t983 VSS.n4591 33.6454
R4351 VSS.n4539 VSS.t686 33.462
R4352 VSS.n4539 VSS.t21 33.462
R4353 VSS.n95 VSS.t2819 33.462
R4354 VSS.n95 VSS.t1602 33.462
R4355 VSS.n103 VSS.t2961 33.462
R4356 VSS.n103 VSS.t2062 33.462
R4357 VSS.n115 VSS.t1404 33.462
R4358 VSS.n115 VSS.t2084 33.462
R4359 VSS.n128 VSS.t1490 33.462
R4360 VSS.n128 VSS.t2087 33.462
R4361 VSS.n170 VSS.t2726 33.462
R4362 VSS.n170 VSS.t1740 33.462
R4363 VSS.n173 VSS.t104 33.462
R4364 VSS.n173 VSS.t1082 33.462
R4365 VSS.n5358 VSS.t2983 33.462
R4366 VSS.n5358 VSS.t1858 33.462
R4367 VSS.n3813 VSS.t202 33.462
R4368 VSS.n3813 VSS.t754 33.462
R4369 VSS.n2254 VSS.t2195 33.462
R4370 VSS.n2254 VSS.t2140 33.462
R4371 VSS.n392 VSS.t2012 33.462
R4372 VSS.n392 VSS.t2938 33.462
R4373 VSS.n4866 VSS.t2705 33.462
R4374 VSS.n4866 VSS.t1807 33.462
R4375 VSS.n4895 VSS.t2980 33.462
R4376 VSS.n4895 VSS.t775 33.462
R4377 VSS.n5002 VSS.t296 33.462
R4378 VSS.n5002 VSS.t2032 33.462
R4379 VSS.n277 VSS.t2882 33.462
R4380 VSS.n277 VSS.t972 33.462
R4381 VSS.n5061 VSS.t1216 33.462
R4382 VSS.n5061 VSS.t2081 33.462
R4383 VSS.n242 VSS.t459 33.462
R4384 VSS.n242 VSS.t2201 33.462
R4385 VSS.n5123 VSS.t2969 33.462
R4386 VSS.n5123 VSS.t716 33.462
R4387 VSS.n5135 VSS.t2934 33.462
R4388 VSS.n5135 VSS.t1874 33.462
R4389 VSS.n226 VSS.t124 33.462
R4390 VSS.n226 VSS.t2701 33.462
R4391 VSS.n5230 VSS.t2994 33.462
R4392 VSS.n5230 VSS.t2034 33.462
R4393 VSS.n199 VSS.t1065 33.462
R4394 VSS.n199 VSS.t290 33.462
R4395 VSS.n188 VSS.t695 33.462
R4396 VSS.n188 VSS.t670 33.462
R4397 VSS.n399 VSS.t2647 33.462
R4398 VSS.n399 VSS.t69 33.462
R4399 VSS.n3331 VSS.t1665 33.2313
R4400 VSS.n3153 VSS.n3152 33.1299
R4401 VSS.n2361 VSS.n2331 33.1299
R4402 VSS.n2353 VSS.n2335 33.1299
R4403 VSS.n1581 VSS.n1580 33.1299
R4404 VSS.n1573 VSS.n1555 33.1299
R4405 VSS.n1298 VSS.n1297 33.1299
R4406 VSS.n4251 VSS.n3756 32.7534
R4407 VSS.n2559 VSS.t274 32.3082
R4408 VSS.n2240 VSS.t61 32.3082
R4409 VSS.n2268 VSS.t57 32.3082
R4410 VSS.n2683 VSS.t262 32.3082
R4411 VSS.n2787 VSS.t266 32.3082
R4412 VSS.n1373 VSS.t238 32.3082
R4413 VSS.n1405 VSS.t244 32.3082
R4414 VSS.n1415 VSS.t242 32.3082
R4415 VSS.n4884 VSS.t270 32.3082
R4416 VSS.n249 VSS.t264 32.3082
R4417 VSS.n309 VSS.n305 32.1808
R4418 VSS.n3333 VSS.n3332 32.0005
R4419 VSS.n2006 VSS.n1358 32.0005
R4420 VSS.n1770 VSS.n1476 32.0005
R4421 VSS.n4645 VSS.n4644 32.0005
R4422 VSS.n1012 VSS.n1004 32.0005
R4423 VSS.n4273 VSS.n4272 31.8805
R4424 VSS.t251 VSS.n1108 31.6734
R4425 VSS.n1150 VSS.t2988 31.6734
R4426 VSS.n4659 VSS.t2986 31.6734
R4427 VSS.n1666 VSS.n1665 31.624
R4428 VSS.n4995 VSS.t2840 31.2987
R4429 VSS.n4988 VSS.t2842 31.2987
R4430 VSS.n3463 VSS.n3462 31.2476
R4431 VSS.n3387 VSS.n3065 31.2476
R4432 VSS.n2827 VSS.n2826 31.2476
R4433 VSS.n1822 VSS.n1447 31.2476
R4434 VSS.t1390 VSS.t2569 31.1531
R4435 VSS.t2628 VSS.t2196 31.1531
R4436 VSS.t2626 VSS.t2198 31.1531
R4437 VSS.n3990 VSS.t801 31.1434
R4438 VSS.n3388 VSS.n3387 30.8711
R4439 VSS.n3370 VSS.n3069 30.8711
R4440 VSS.n1823 VSS.n1822 30.8711
R4441 VSS.n3955 VSS.n3950 30.7665
R4442 VSS.n4015 VSS.n3996 30.4946
R4443 VSS.n4071 VSS.n4070 30.4946
R4444 VSS.n4122 VSS.n4121 30.4946
R4445 VSS.n3262 VSS.n3118 30.4946
R4446 VSS.n3312 VSS.t1502 30.462
R4447 VSS.n3312 VSS.t1368 30.462
R4448 VSS.n3619 VSS.t622 30.462
R4449 VSS.n3619 VSS.t2754 30.462
R4450 VSS.t2733 VSS.n4648 29.907
R4451 VSS.n4648 VSS.t2735 29.907
R4452 VSS.t2735 VSS.t2011 29.907
R4453 VSS.n4814 VSS.t560 29.907
R4454 VSS.t560 VSS.n4813 29.907
R4455 VSS.n4813 VSS.t549 29.907
R4456 VSS.t2739 VSS.n1260 29.907
R4457 VSS.n3444 VSS.n3443 29.7417
R4458 VSS.n1968 VSS.n1967 29.7417
R4459 VSS.n1830 VSS.n1829 29.7417
R4460 VSS.n1808 VSS.n1454 29.7417
R4461 VSS.n1789 VSS.n1466 29.7417
R4462 VSS.n1729 VSS.n1728 29.7417
R4463 VSS.n310 VSS.n309 29.2561
R4464 VSS.n345 VSS.n343 28.9887
R4465 VSS.n2788 VSS.n2168 28.9887
R4466 VSS.n4502 VSS.t1240 28.7917
R4467 VSS.n4499 VSS.t2675 28.7917
R4468 VSS.n176 VSS.t1031 28.7917
R4469 VSS.n5361 VSS.t1759 28.7917
R4470 VSS.n3845 VSS.t1742 28.7917
R4471 VSS.n3848 VSS.t1204 28.7917
R4472 VSS.n3850 VSS.t2636 28.7917
R4473 VSS.n3875 VSS.t2695 28.7917
R4474 VSS.n3876 VSS.t1137 28.7917
R4475 VSS.n4440 VSS.t2127 28.7917
R4476 VSS.n4441 VSS.t2276 28.7917
R4477 VSS.n4436 VSS.t2649 28.7917
R4478 VSS.n4437 VSS.t1668 28.7917
R4479 VSS.n4433 VSS.t732 28.7917
R4480 VSS.n3158 VSS.t873 28.7917
R4481 VSS.n3134 VSS.t1086 28.7917
R4482 VSS.n3137 VSS.t1897 28.7917
R4483 VSS.n3138 VSS.t1354 28.7917
R4484 VSS.n2086 VSS.t1655 28.7917
R4485 VSS.n2094 VSS.t2106 28.7917
R4486 VSS.n2082 VSS.t1518 28.7917
R4487 VSS.n2083 VSS.t1449 28.7917
R4488 VSS.n2267 VSS.t2122 28.7917
R4489 VSS.n2330 VSS.t1523 28.7917
R4490 VSS.n2333 VSS.t2184 28.7917
R4491 VSS.n2337 VSS.t2630 28.7917
R4492 VSS.n2339 VSS.t1125 28.7917
R4493 VSS.n2860 VSS.t1375 28.7917
R4494 VSS.n2861 VSS.t938 28.7917
R4495 VSS.n2868 VSS.t744 28.7917
R4496 VSS.n2869 VSS.t1048 28.7917
R4497 VSS.n1475 VSS.t1708 28.7917
R4498 VSS.n1591 VSS.t1944 28.7917
R4499 VSS.n1548 VSS.t2014 28.7917
R4500 VSS.n1551 VSS.t738 28.7917
R4501 VSS.n1554 VSS.t1992 28.7917
R4502 VSS.n1557 VSS.t2113 28.7917
R4503 VSS.n1559 VSS.t1455 28.7917
R4504 VSS.n1276 VSS.t1585 28.7917
R4505 VSS.n1277 VSS.t944 28.7917
R4506 VSS.n1272 VSS.t806 28.7917
R4507 VSS.n1273 VSS.t2174 28.7917
R4508 VSS.n1269 VSS.t833 28.7917
R4509 VSS.n387 VSS.t932 28.7917
R4510 VSS.n4879 VSS.t1326 28.7917
R4511 VSS.n4893 VSS.t1698 28.7917
R4512 VSS.n286 VSS.t898 28.7917
R4513 VSS.n5048 VSS.t1926 28.7917
R4514 VSS.n257 VSS.t2268 28.7917
R4515 VSS.n245 VSS.t726 28.7917
R4516 VSS.n5129 VSS.t1883 28.7917
R4517 VSS.n233 VSS.t2697 28.7917
R4518 VSS.n217 VSS.t902 28.7917
R4519 VSS.n202 VSS.t2566 28.7917
R4520 VSS.n5283 VSS.t2256 28.7917
R4521 VSS.n184 VSS.t2604 28.7917
R4522 VSS.n5311 VSS.t1544 28.7917
R4523 VSS.n5318 VSS.t927 28.7917
R4524 VSS.n400 VSS.t2568 28.7917
R4525 VSS.n403 VSS.t2197 28.7917
R4526 VSS.n406 VSS.t769 28.7917
R4527 VSS.n3988 VSS.t119 28.6159
R4528 VSS.n3988 VSS.t2806 28.6159
R4529 VSS.n3090 VSS.t1263 28.6159
R4530 VSS.n3090 VSS.t2890 28.6159
R4531 VSS.n3783 VSS.t1410 28.3801
R4532 VSS.n2946 VSS.t1880 28.3801
R4533 VSS.n3020 VSS.t994 28.3801
R4534 VSS.n3049 VSS.t2582 28.3801
R4535 VSS.n2213 VSS.t1017 28.3801
R4536 VSS.n2260 VSS.t740 28.3801
R4537 VSS.n2647 VSS.t1333 28.3801
R4538 VSS.n2802 VSS.t1223 28.3801
R4539 VSS.n2806 VSS.t2028 28.3801
R4540 VSS.n3825 VSS.t2103 28.3166
R4541 VSS.n3788 VSS.t1813 28.3166
R4542 VSS.n3017 VSS.t2163 28.3166
R4543 VSS.n3099 VSS.t1063 28.3166
R4544 VSS.n2203 VSS.t2619 28.3166
R4545 VSS.n2221 VSS.t1775 28.3166
R4546 VSS.n2236 VSS.t1907 28.3166
R4547 VSS.n2280 VSS.t1757 28.3166
R4548 VSS.n2193 VSS.t1534 28.3166
R4549 VSS.n2674 VSS.t720 28.3166
R4550 VSS.n2763 VSS.t1155 28.3166
R4551 VSS.n1355 VSS.t2056 28.3166
R4552 VSS.n4546 VSS.n4545 28.2358
R4553 VSS.n5758 VSS.n5757 28.2358
R4554 VSS.n5648 VSS.n61 28.2358
R4555 VSS.n4020 VSS.n4019 28.2358
R4556 VSS.n4209 VSS.n4208 28.2358
R4557 VSS.n3324 VSS.n3088 28.2358
R4558 VSS.n3257 VSS.n3256 28.2358
R4559 VSS.n2874 VSS.n2850 28.2358
R4560 VSS.t2638 VSS.t2628 28.0379
R4561 VSS.n4289 VSS.n4288 27.8593
R4562 VSS.n2013 VSS.n1353 27.8593
R4563 VSS.n1958 VSS.n1379 27.8593
R4564 VSS.n1903 VSS.n1403 27.8593
R4565 VSS.n1862 VSS.n1427 27.8593
R4566 VSS.n1804 VSS.n1803 27.8593
R4567 VSS.n1783 VSS.n1468 27.8593
R4568 VSS.n1759 VSS.n1479 27.8593
R4569 VSS.n3959 VSS.n3816 27.6711
R4570 VSS.n3574 VSS.n3570 27.6711
R4571 VSS.n122 VSS.t1350 27.5691
R4572 VSS.n3753 VSS.t1318 27.5691
R4573 VSS.n4836 VSS.t1117 27.5691
R4574 VSS.n4233 VSS.n4232 27.4829
R4575 VSS.n4293 VSS.n3740 27.4829
R4576 VSS.n2734 VSS.n2660 27.4829
R4577 VSS.n1657 VSS.n1656 27.4829
R4578 VSS.n4131 VSS.n3771 27.1064
R4579 VSS.n4153 VSS.n4152 27.1064
R4580 VSS.n4355 VSS.n4354 27.1064
R4581 VSS.n3511 VSS.n3003 27.1064
R4582 VSS.n3375 VSS.n3374 27.1064
R4583 VSS.n3269 VSS.n3268 27.1064
R4584 VSS.n1734 VSS.n1733 27.1064
R4585 VSS.n4025 VSS.n3993 26.7299
R4586 VSS.n4417 VSS.n4416 26.7299
R4587 VSS.n3545 VSS.n3544 26.7299
R4588 VSS.n3319 VSS.n3318 26.7299
R4589 VSS.n3251 VSS.n3122 26.7299
R4590 VSS.n3106 VSS.n3105 26.7039
R4591 VSS.n3111 VSS.n3110 26.7039
R4592 VSS.n5398 VSS.n5396 26.6009
R4593 VSS.n2927 VSS.n2926 26.6009
R4594 VSS.n4026 VSS.n4025 26.3813
R4595 VSS.n2785 VSS.n2170 26.3534
R4596 VSS.n2820 VSS.n2819 26.3534
R4597 VSS.n5550 VSS.n5549 26.314
R4598 VSS.n5456 VSS.n147 26.314
R4599 VSS.n5418 VSS.n5417 26.314
R4600 VSS.n2103 VSS.n2102 26.314
R4601 VSS.n4459 VSS.n4458 26.1349
R4602 VSS.n4098 VSS.n4097 25.977
R4603 VSS.n4280 VSS.n3745 25.977
R4604 VSS.n3632 VSS.n2952 25.977
R4605 VSS.n3474 VSS.n3025 25.977
R4606 VSS.n3411 VSS.n3410 25.977
R4607 VSS.n2590 VSS.n2219 25.977
R4608 VSS.n2498 VSS.n2265 25.977
R4609 VSS.n2796 VSS.n2166 25.977
R4610 VSS.n1927 VSS.n1926 25.977
R4611 VSS.n4864 VSS.n375 25.977
R4612 VSS.n4910 VSS.n4909 25.977
R4613 VSS.n5100 VSS.n5099 25.977
R4614 VSS.n5169 VSS.n5127 25.977
R4615 VSS.n5211 VSS.n5210 25.977
R4616 VSS.n5248 VSS.n206 25.977
R4617 VSS.n4063 VSS.t844 25.9346
R4618 VSS.n3593 VSS.t980 25.9346
R4619 VSS.n1516 VSS.t2892 25.8467
R4620 VSS.n1516 VSS.t641 25.8467
R4621 VSS.n1522 VSS.t1406 25.8467
R4622 VSS.n1522 VSS.t1408 25.8467
R4623 VSS.n4296 VSS.n4295 25.7355
R4624 VSS.n5738 VSS.n5737 25.7355
R4625 VSS.n5590 VSS.n88 25.7355
R4626 VSS.n4304 VSS.n4302 25.7355
R4627 VSS.n2780 VSS.n2170 25.7355
R4628 VSS.n1896 VSS.n1894 25.7355
R4629 VSS.n1887 VSS.n1886 25.7355
R4630 VSS.n1703 VSS.n1702 25.7355
R4631 VSS.n1636 VSS.n1530 25.7355
R4632 VSS.n4821 VSS.n4820 25.7355
R4633 VSS.n5031 VSS.n5030 25.7355
R4634 VSS.n5282 VSS.n192 25.7355
R4635 VSS.n5294 VSS.n187 25.7355
R4636 VSS.n5682 VSS.n5681 25.6926
R4637 VSS.n5612 VSS.n5610 25.6926
R4638 VSS.n5556 VSS.n5555 25.6926
R4639 VSS.n5521 VSS.n5519 25.6926
R4640 VSS.n5472 VSS.n5470 25.6926
R4641 VSS.n5427 VSS.n5425 25.6926
R4642 VSS.n3923 VSS.n3919 25.6926
R4643 VSS.n3979 VSS.n3976 25.6926
R4644 VSS.n4073 VSS.n4071 25.6926
R4645 VSS.n4113 VSS.n4112 25.6926
R4646 VSS.n4230 VSS.n4171 25.6926
R4647 VSS.n4221 VSS.n4174 25.6926
R4648 VSS.n4255 VSS.n4254 25.6926
R4649 VSS.n3466 VSS.n3463 25.6926
R4650 VSS.n3396 VSS.n3060 25.6926
R4651 VSS.n2613 VSS.n2208 25.6926
R4652 VSS.n2722 VSS.n2721 25.6926
R4653 VSS.n2058 VSS.n1334 25.6926
R4654 VSS.n1908 VSS.n1403 25.6926
R4655 VSS.n1863 VSS.n1862 25.6926
R4656 VSS.n1685 VSS.n1684 25.6926
R4657 VSS.n4871 VSS.n373 25.6926
R4658 VSS.n5012 VSS.n5011 25.6926
R4659 VSS.n5026 VSS.n5025 25.6926
R4660 VSS.n5060 VSS.n264 25.6926
R4661 VSS.n5071 VSS.n5070 25.6926
R4662 VSS.n5113 VSS.n5112 25.6926
R4663 VSS.n5119 VSS.n236 25.6926
R4664 VSS.n5153 VSS.n5152 25.6926
R4665 VSS.n5141 VSS.n235 25.6926
R4666 VSS.n5187 VSS.n5186 25.6926
R4667 VSS.n5194 VSS.n5193 25.6926
R4668 VSS.n5200 VSS.n5199 25.6926
R4669 VSS.n5235 VSS.n210 25.6926
R4670 VSS.n5243 VSS.n5242 25.6926
R4671 VSS.n453 VSS.n397 25.6926
R4672 VSS.n4973 VSS.n349 25.6576
R4673 VSS.n4520 VSS.n4518 25.6005
R4674 VSS.n4527 VSS.n4526 25.6005
R4675 VSS.n4533 VSS.n4532 25.6005
R4676 VSS.n4551 VSS.n4495 25.6005
R4677 VSS.n5764 VSS.n5763 25.6005
R4678 VSS.n5732 VSS.n5731 25.6005
R4679 VSS.n5693 VSS.n5692 25.6005
R4680 VSS.n5675 VSS.n5674 25.6005
R4681 VSS.n5641 VSS.n66 25.6005
R4682 VSS.n5607 VSS.n82 25.6005
R4683 VSS.n5383 VSS.n5382 25.6005
R4684 VSS.n5371 VSS.n5370 25.6005
R4685 VSS.n3857 VSS.n3851 25.6005
R4686 VSS.n3874 VSS.n3843 25.6005
R4687 VSS.n4448 VSS.n4447 25.6005
R4688 VSS.n4454 VSS.n4453 25.6005
R4689 VSS.n3145 VSS.n3144 25.6005
R4690 VSS.n2087 VSS.n2085 25.6005
R4691 VSS.n2097 VSS.n2081 25.6005
R4692 VSS.n2502 VSS.n2501 25.6005
R4693 VSS.n2346 VSS.n2340 25.6005
R4694 VSS.n2859 VSS.n2858 25.6005
R4695 VSS.n2867 VSS.n2866 25.6005
R4696 VSS.n1771 VSS.n1770 25.6005
R4697 VSS.n1566 VSS.n1560 25.6005
R4698 VSS.n1284 VSS.n1283 25.6005
R4699 VSS.n1290 VSS.n1289 25.6005
R4700 VSS.n4829 VSS.n4828 25.6005
R4701 VSS.n4930 VSS.n4929 25.6005
R4702 VSS.n4903 VSS.n4902 25.6005
R4703 VSS.n5018 VSS.n5017 25.6005
R4704 VSS.n5047 VSS.n5046 25.6005
R4705 VSS.n5077 VSS.n5076 25.6005
R4706 VSS.n5107 VSS.n5106 25.6005
R4707 VSS.n5163 VSS.n5130 25.6005
R4708 VSS.n5181 VSS.n232 25.6005
R4709 VSS.n5217 VSS.n5216 25.6005
R4710 VSS.n5264 VSS.n5263 25.6005
R4711 VSS.n5285 VSS.n190 25.6005
R4712 VSS.n5305 VSS.n5304 25.6005
R4713 VSS.n5313 VSS.n180 25.6005
R4714 VSS.n5320 VSS.n178 25.6005
R4715 VSS.n5340 VSS.n5339 25.6005
R4716 VSS.n443 VSS.n442 25.6005
R4717 VSS.n437 VSS.n436 25.6005
R4718 VSS.n431 VSS.n430 25.6005
R4719 VSS.n424 VSS.n423 25.6005
R4720 VSS.n3860 VSS.n3859 25.5964
R4721 VSS.n2699 VSS.n2698 25.5564
R4722 VSS.n1062 VSS.n1046 25.4945
R4723 VSS.n125 VSS.t1335 25.4291
R4724 VSS.n4162 VSS.t2608 25.4291
R4725 VSS.n4243 VSS.t982 25.4291
R4726 VSS.n4346 VSS.t2178 25.4291
R4727 VSS.n4371 VSS.t869 25.4291
R4728 VSS.n4403 VSS.t1302 25.4291
R4729 VSS.n2141 VSS.t1986 25.4291
R4730 VSS.n2983 VSS.t1795 25.4291
R4731 VSS.n2993 VSS.t2064 25.4291
R4732 VSS.n3006 VSS.t1711 25.4291
R4733 VSS.n3010 VSS.t1200 25.4291
R4734 VSS.n3039 VSS.t1182 25.4291
R4735 VSS.n3053 VSS.t1836 25.4291
R4736 VSS.n3091 VSS.t1269 25.4291
R4737 VSS.n2299 VSS.t2131 25.4291
R4738 VSS.n2807 VSS.t893 25.4291
R4739 VSS.n2162 VSS.t1889 25.4291
R4740 VSS.n1432 VSS.t958 25.4291
R4741 VSS.n1744 VSS.t777 25.4291
R4742 VSS.n3272 VSS.n3271 25.3161
R4743 VSS.n616 VSS.n548 25.3005
R4744 VSS.n616 VSS.n615 25.3005
R4745 VSS.n788 VSS.n770 25.3005
R4746 VSS.n855 VSS.n770 25.3005
R4747 VSS.n4675 VSS.n617 25.2897
R4748 VSS.n911 VSS.n910 25.2897
R4749 VSS.t3405 VSS.t2072 25.2879
R4750 VSS.t389 VSS.t2065 25.2879
R4751 VSS.t813 VSS.t1006 25.2879
R4752 VSS.t2121 VSS.t779 25.2879
R4753 VSS.t3411 VSS.t1148 25.2879
R4754 VSS.t1156 VSS.t1705 25.2879
R4755 VSS.n3565 VSS.n2979 25.224
R4756 VSS.n5756 VSS.n14 25.224
R4757 VSS.n5757 VSS.n5756 25.224
R4758 VSS.n5652 VSS.n61 25.224
R4759 VSS.n5653 VSS.n5652 25.224
R4760 VSS.n3950 VSS.n3949 25.224
R4761 VSS.n4248 VSS.n3758 25.224
R4762 VSS.n4268 VSS.n4267 25.224
R4763 VSS.n4308 VSS.n4307 25.224
R4764 VSS.n4345 VSS.n3718 25.224
R4765 VSS.n3544 VSS.n3543 25.224
R4766 VSS.n3255 VSS.n3122 25.224
R4767 VSS.n3256 VSS.n3255 25.224
R4768 VSS.n2876 VSS.n2875 25.224
R4769 VSS.n2875 VSS.n2874 25.224
R4770 VSS.n2881 VSS.n2880 25.224
R4771 VSS.n2880 VSS.n2848 25.224
R4772 VSS.n1586 VSS.n1549 25.224
R4773 VSS.n4865 VSS.n4864 25.224
R4774 VSS.n4909 VSS.n4908 25.224
R4775 VSS.n5101 VSS.n5100 25.224
R4776 VSS.n5165 VSS.n5127 25.224
R4777 VSS.n5212 VSS.n5211 25.224
R4778 VSS.n5249 VSS.n5248 25.224
R4779 VSS.n4675 VSS.n4674 25.1992
R4780 VSS.n912 VSS.n911 25.1992
R4781 VSS.n5488 VSS.n5487 24.9894
R4782 VSS.n3614 VSS.n3613 24.9894
R4783 VSS.n3367 VSS.n3073 24.9894
R4784 VSS.n3307 VSS.n3305 24.9894
R4785 VSS.n981 VSS.t2659 24.9236
R4786 VSS.n981 VSS.t2665 24.9236
R4787 VSS.n1167 VSS.t2948 24.9236
R4788 VSS.n1167 VSS.t2942 24.9236
R4789 VSS.n328 VSS.t1769 24.9236
R4790 VSS.n328 VSS.t1773 24.9236
R4791 VSS.n327 VSS.t1781 24.9236
R4792 VSS.n327 VSS.t1779 24.9236
R4793 VSS.n341 VSS.t2669 24.9236
R4794 VSS.n341 VSS.t2673 24.9236
R4795 VSS.n344 VSS.t2667 24.9236
R4796 VSS.n344 VSS.t2830 24.9236
R4797 VSS.n4001 VSS.t1287 24.9236
R4798 VSS.n4003 VSS.t1723 24.9236
R4799 VSS.n4003 VSS.t1121 24.9236
R4800 VSS.n3742 VSS.t1803 24.9236
R4801 VSS.n3742 VSS.t1801 24.9236
R4802 VSS.n3739 VSS.t618 24.9236
R4803 VSS.n3714 VSS.t2222 24.9236
R4804 VSS.n3714 VSS.t2220 24.9236
R4805 VSS.n3711 VSS.t2997 24.9236
R4806 VSS.n3711 VSS.t376 24.9236
R4807 VSS.n3082 VSS.t1007 24.9236
R4808 VSS.n3331 VSS.t455 24.9236
R4809 VSS.n2559 VSS.t1021 24.9236
R4810 VSS.n2240 VSS.t1548 24.9236
R4811 VSS.n2518 VSS.t2824 24.9236
R4812 VSS.n2263 VSS.t1271 24.9236
R4813 VSS.n2263 VSS.t380 24.9236
R4814 VSS.n2268 VSS.t780 24.9236
R4815 VSS.n2289 VSS.t1372 24.9236
R4816 VSS.n2415 VSS.t1866 24.9236
R4817 VSS.n2415 VSS.t1860 24.9236
R4818 VSS.n2679 VSS.t272 24.9236
R4819 VSS.n2679 VSS.t236 24.9236
R4820 VSS.n2683 VSS.t1834 24.9236
R4821 VSS.n2682 VSS.t240 24.9236
R4822 VSS.n2682 VSS.t276 24.9236
R4823 VSS.n2787 VSS.t2115 24.9236
R4824 VSS.n1356 VSS.t1620 24.9236
R4825 VSS.n1356 VSS.t1618 24.9236
R4826 VSS.n1373 VSS.t1101 24.9236
R4827 VSS.n1382 VSS.t1479 24.9236
R4828 VSS.n1382 VSS.t1485 24.9236
R4829 VSS.n1390 VSS.t2203 24.9236
R4830 VSS.n1390 VSS.t2205 24.9236
R4831 VSS.n1405 VSS.t2022 24.9236
R4832 VSS.n1406 VSS.t1721 24.9236
R4833 VSS.n1406 VSS.t1713 24.9236
R4834 VSS.n1415 VSS.t1982 24.9236
R4835 VSS.n1643 VSS.t1630 24.9236
R4836 VSS.n1643 VSS.t1634 24.9236
R4837 VSS.n1429 VSS.t960 24.9236
R4838 VSS.n1429 VSS.t966 24.9236
R4839 VSS.n1456 VSS.t1165 24.9236
R4840 VSS.n1456 VSS.t1167 24.9236
R4841 VSS.n1470 VSS.t1310 24.9236
R4842 VSS.n1470 VSS.t1312 24.9236
R4843 VSS.n1483 VSS.t1248 24.9236
R4844 VSS.n1483 VSS.t1242 24.9236
R4845 VSS.n1506 VSS.t1959 24.9236
R4846 VSS.n1506 VSS.t1957 24.9236
R4847 VSS.n4884 VSS.t1457 24.9236
R4848 VSS.n249 VSS.t1696 24.9236
R4849 VSS.n472 VSS.t2954 24.9236
R4850 VSS.n472 VSS.t2944 24.9236
R4851 VSS.n4603 VSS.t2627 24.9236
R4852 VSS.n4603 VSS.t2625 24.9236
R4853 VSS.t2646 VSS.t2737 24.9226
R4854 VSS.n4531 VSS.n4503 24.8476
R4855 VSS.n4537 VSS.n4500 24.8476
R4856 VSS.n5384 VSS.n174 24.8476
R4857 VSS.n5372 VSS.n5359 24.8476
R4858 VSS.n3859 VSS.n3858 24.8476
R4859 VSS.n3878 VSS.n3877 24.8476
R4860 VSS.n4130 VSS.n4129 24.8476
R4861 VSS.n4156 VSS.n4155 24.8476
R4862 VSS.n4161 VSS.n4160 24.8476
R4863 VSS.n4216 VSS.n4215 24.8476
R4864 VSS.n4294 VSS.n4293 24.8476
R4865 VSS.n4383 VSS.n3706 24.8476
R4866 VSS.n4452 VSS.n4442 24.8476
R4867 VSS.n4458 VSS.n4438 24.8476
R4868 VSS.n3642 VSS.n2944 24.8476
R4869 VSS.n3550 VSS.n2989 24.8476
R4870 VSS.n3539 VSS.n2991 24.8476
R4871 VSS.n3244 VSS.n3125 24.8476
R4872 VSS.n3149 VSS.n3139 24.8476
R4873 VSS.n2096 VSS.n2095 24.8476
R4874 VSS.n2102 VSS.n2101 24.8476
R4875 VSS.n2614 VSS.n2613 24.8476
R4876 VSS.n2466 VSS.n2465 24.8476
R4877 VSS.n2348 VSS.n2347 24.8476
R4878 VSS.n2862 VSS.n2852 24.8476
R4879 VSS.n2870 VSS.n2850 24.8476
R4880 VSS.n2655 VSS.n2654 24.8476
R4881 VSS.n2711 VSS.n2671 24.8476
R4882 VSS.n2021 VSS.n1347 24.8476
R4883 VSS.n1944 VSS.n1943 24.8476
R4884 VSS.n1809 VSS.n1808 24.8476
R4885 VSS.n1766 VSS.n1765 24.8476
R4886 VSS.n1704 VSS.n1703 24.8476
R4887 VSS.n1651 VSS.n1650 24.8476
R4888 VSS.n1587 VSS.n1586 24.8476
R4889 VSS.n1568 VSS.n1567 24.8476
R4890 VSS.n1288 VSS.n1278 24.8476
R4891 VSS.n1294 VSS.n1274 24.8476
R4892 VSS.n4847 VSS.n4834 24.8476
R4893 VSS.n4833 VSS.n388 24.8476
R4894 VSS.n4934 VSS.n4880 24.8476
R4895 VSS.n4904 VSS.n4891 24.8476
R4896 VSS.n5016 VSS.n285 24.8476
R4897 VSS.n5049 VSS.n268 24.8476
R4898 VSS.n5075 VSS.n256 24.8476
R4899 VSS.n5105 VSS.n244 24.8476
R4900 VSS.n5165 VSS.n5164 24.8476
R4901 VSS.n5186 VSS.n5185 24.8476
R4902 VSS.n5212 VSS.n218 24.8476
R4903 VSS.n5262 VSS.n201 24.8476
R4904 VSS.n5284 VSS.n5282 24.8476
R4905 VSS.n5300 VSS.n185 24.8476
R4906 VSS.n5312 VSS.n5310 24.8476
R4907 VSS.n5319 VSS.n5317 24.8476
R4908 VSS.n447 VSS.n401 24.8476
R4909 VSS.n441 VSS.n404 24.8476
R4910 VSS.n435 VSS.n407 24.8476
R4911 VSS.t1697 VSS.n4988 24.7782
R4912 VSS.n4276 VSS.n3745 24.5331
R4913 VSS.n4521 VSS.n4520 24.4711
R4914 VSS.n4525 VSS.n4506 24.4711
R4915 VSS.n4552 VSS.n4551 24.4711
R4916 VSS.n4554 VSS.n4493 24.4711
R4917 VSS.n5763 VSS.n5762 24.4711
R4918 VSS.n5758 VSS.n12 24.4711
R4919 VSS.n5737 VSS.n23 24.4711
R4920 VSS.n5733 VSS.n5732 24.4711
R4921 VSS.n5698 VSS.n39 24.4711
R4922 VSS.n5694 VSS.n5693 24.4711
R4923 VSS.n5680 VSS.n48 24.4711
R4924 VSS.n5676 VSS.n5675 24.4711
R4925 VSS.n5647 VSS.n5646 24.4711
R4926 VSS.n5645 VSS.n66 24.4711
R4927 VSS.n5603 VSS.n82 24.4711
R4928 VSS.n5602 VSS.n5601 24.4711
R4929 VSS.n5580 VSS.n5579 24.4711
R4930 VSS.n5512 VSS.n5511 24.4711
R4931 VSS.n5457 VSS.n5456 24.4711
R4932 VSS.n5418 VSS.n161 24.4711
R4933 VSS.n4116 VSS.n4113 24.4711
R4934 VSS.n4238 VSS.n4168 24.4711
R4935 VSS.n4217 VSS.n4174 24.4711
R4936 VSS.n3268 VSS.n3115 24.4711
R4937 VSS.n3264 VSS.n3115 24.4711
R4938 VSS.n2445 VSS.n2444 24.4711
R4939 VSS.n1997 VSS.n1364 24.4711
R4940 VSS.n1931 VSS.n1393 24.4711
R4941 VSS.n1927 VSS.n1393 24.4711
R4942 VSS.n1876 VSS.n1875 24.4711
R4943 VSS.n1849 VSS.n1434 24.4711
R4944 VSS.n1621 VSS.n1532 24.4711
R4945 VSS.n1620 VSS.n1619 24.4711
R4946 VSS.n4860 VSS.n4859 24.4711
R4947 VSS.n4860 VSS.n375 24.4711
R4948 VSS.n4911 VSS.n4888 24.4711
R4949 VSS.n4911 VSS.n4910 24.4711
R4950 VSS.n5095 VSS.n247 24.4711
R4951 VSS.n5099 VSS.n247 24.4711
R4952 VSS.n5171 VSS.n5170 24.4711
R4953 VSS.n5170 VSS.n5169 24.4711
R4954 VSS.n5210 VSS.n220 24.4711
R4955 VSS.n5244 VSS.n5243 24.4711
R4956 VSS.n5244 VSS.n206 24.4711
R4957 VSS.n5342 VSS.n5324 24.4711
R4958 VSS.n5341 VSS.n5340 24.4711
R4959 VSS.n429 VSS.n410 24.4711
R4960 VSS.n425 VSS.n424 24.4711
R4961 VSS.n3325 VSS.n3324 24.3177
R4962 VSS.n4521 VSS.n4506 24.0946
R4963 VSS.n4526 VSS.n4525 24.0946
R4964 VSS.n4532 VSS.n4531 24.0946
R4965 VSS.n4554 VSS.n4552 24.0946
R4966 VSS.n5762 VSS.n12 24.0946
R4967 VSS.n5733 VSS.n23 24.0946
R4968 VSS.n5694 VSS.n39 24.0946
R4969 VSS.n5676 VSS.n48 24.0946
R4970 VSS.n5646 VSS.n5645 24.0946
R4971 VSS.n5603 VSS.n5602 24.0946
R4972 VSS.n5581 VSS.n5580 24.0946
R4973 VSS.n5504 VSS.n123 24.0946
R4974 VSS.n5458 VSS.n5457 24.0946
R4975 VSS.n5422 VSS.n161 24.0946
R4976 VSS.n4041 VSS.n3986 24.0946
R4977 VSS.n4116 VSS.n3777 24.0946
R4978 VSS.n4121 VSS.n4120 24.0946
R4979 VSS.n4234 VSS.n4168 24.0946
R4980 VSS.n4217 VSS.n4216 24.0946
R4981 VSS.n4251 VSS.n4250 24.0946
R4982 VSS.n4453 VSS.n4452 24.0946
R4983 VSS.n3637 VSS.n3636 24.0946
R4984 VSS.n3482 VSS.n3481 24.0946
R4985 VSS.n3418 VSS.n3417 24.0946
R4986 VSS.n2097 VSS.n2096 24.0946
R4987 VSS.n2622 VSS.n2201 24.0946
R4988 VSS.n2484 VSS.n2483 24.0946
R4989 VSS.n2866 VSS.n2852 24.0946
R4990 VSS.n1845 VSS.n1434 24.0946
R4991 VSS.n1772 VSS.n1771 24.0946
R4992 VSS.n1621 VSS.n1620 24.0946
R4993 VSS.n1289 VSS.n1288 24.0946
R4994 VSS.n4929 VSS.n4928 24.0946
R4995 VSS.n4916 VSS.n4915 24.0946
R4996 VSS.n4902 VSS.n4901 24.0946
R4997 VSS.n5083 VSS.n5082 24.0946
R4998 VSS.n5107 VSS.n241 24.0946
R4999 VSS.n5264 VSS.n198 24.0946
R5000 VSS.n5306 VSS.n5305 24.0946
R5001 VSS.n5317 VSS.n180 24.0946
R5002 VSS.n5342 VSS.n5341 24.0946
R5003 VSS.n442 VSS.n441 24.0946
R5004 VSS.n436 VSS.n435 24.0946
R5005 VSS.n430 VSS.n429 24.0946
R5006 VSS.n425 VSS.n410 24.0946
R5007 VSS.n3117 VSS.t1735 24.0005
R5008 VSS.n2275 VSS.t573 24.0005
R5009 VSS.n1018 VSS.t1255 23.988
R5010 VSS.n4584 VSS.n4493 23.7181
R5011 VSS.n5699 VSS.n5698 23.7181
R5012 VSS.n5610 VSS.n5609 23.7181
R5013 VSS.n5574 VSS.n5573 23.7181
R5014 VSS.n5517 VSS.n116 23.7181
R5015 VSS.n5513 VSS.n116 23.7181
R5016 VSS.n5505 VSS.n5504 23.7181
R5017 VSS.n5470 VSS.n5469 23.7181
R5018 VSS.n5425 VSS.n5424 23.7181
R5019 VSS.n5378 VSS.n5356 23.7181
R5020 VSS.n3919 VSS.n3918 23.7181
R5021 VSS.n4057 VSS.n3806 23.7181
R5022 VSS.n4058 VSS.n4057 23.7181
R5023 VSS.n4239 VSS.n3761 23.7181
R5024 VSS.n4239 VSS.n4238 23.7181
R5025 VSS.n4242 VSS.n3760 23.7181
R5026 VSS.n4268 VSS.n3748 23.7181
R5027 VSS.n3689 VSS.n3688 23.7181
R5028 VSS.n3628 VSS.n3627 23.7181
R5029 VSS.n3345 VSS.n3344 23.7181
R5030 VSS.n2599 VSS.n2211 23.7181
R5031 VSS.n2593 VSS.n2214 23.7181
R5032 VSS.n2556 VSS.n2233 23.7181
R5033 VSS.n2557 VSS.n2556 23.7181
R5034 VSS.n2451 VSS.n2287 23.7181
R5035 VSS.n2735 VSS.n2734 23.7181
R5036 VSS.n2796 VSS.n2795 23.7181
R5037 VSS.n2834 VSS.n2166 23.7181
R5038 VSS.n1327 VSS.n1261 23.7181
R5039 VSS.n2001 VSS.n2000 23.7181
R5040 VSS.n1747 VSS.n1742 23.7181
R5041 VSS.n1742 VSS.n1741 23.7181
R5042 VSS.n1670 VSS.n1517 23.7181
R5043 VSS.n4816 VSS.n4815 23.7181
R5044 VSS.n4935 VSS.n4934 23.7181
R5045 VSS.n4997 VSS.n295 23.7181
R5046 VSS.n4997 VSS.n293 23.7181
R5047 VSS.n5004 VSS.n291 23.7181
R5048 VSS.n5053 VSS.n268 23.7181
R5049 VSS.n5063 VSS.n262 23.7181
R5050 VSS.n5081 VSS.n254 23.7181
R5051 VSS.n5177 VSS.n236 23.7181
R5052 VSS.n5177 VSS.n5176 23.7181
R5053 VSS.n5150 VSS.n5137 23.7181
R5054 VSS.n5180 VSS.n235 23.7181
R5055 VSS.n5228 VSS.n212 23.7181
R5056 VSS.n5274 VSS.n195 23.7181
R5057 VSS.n5347 VSS.n5346 23.7181
R5058 VSS.n1143 VSS.n1141 23.4005
R5059 VSS.n1143 VSS.n950 23.4005
R5060 VSS.n1142 VSS.n1140 23.4005
R5061 VSS.n1142 VSS.n1109 23.4005
R5062 VSS.n947 VSS.n943 23.4005
R5063 VSS.n1237 VSS.n943 23.4005
R5064 VSS.n4662 VSS.n4661 23.4005
R5065 VSS.n4661 VSS.n476 23.4005
R5066 VSS.n4097 VSS.n3789 23.3417
R5067 VSS.n1871 VSS.n1870 23.3417
R5068 VSS.n1123 VSS.n1121 23.1134
R5069 VSS.n925 VSS.n923 23.1134
R5070 VSS.n4649 VSS.t3154 23.0535
R5071 VSS.n2357 VSS.n2356 22.9652
R5072 VSS.n1576 VSS.n1552 22.9652
R5073 VSS.n5510 VSS.n120 22.9652
R5074 VSS.n4100 VSS.n3785 22.9652
R5075 VSS.n4129 VSS.n4128 22.9652
R5076 VSS.n4156 VSS.n3764 22.9652
R5077 VSS.n4163 VSS.n3761 22.9652
R5078 VSS.n4194 VSS.n4190 22.9652
R5079 VSS.n4347 VSS.n4345 22.9652
R5080 VSS.n4372 VSS.n3708 22.9652
R5081 VSS.n4404 VSS.n4402 22.9652
R5082 VSS.n3684 VSS.n3683 22.9652
R5083 VSS.n3666 VSS.n3665 22.9652
R5084 VSS.n3562 VSS.n3561 22.9652
R5085 VSS.n3538 VSS.n3537 22.9652
R5086 VSS.n3503 VSS.n3502 22.9652
R5087 VSS.n3479 VSS.n3478 22.9652
R5088 VSS.n3445 VSS.n3444 22.9652
R5089 VSS.n3412 VSS.n3411 22.9652
R5090 VSS.n3340 VSS.n3339 22.9652
R5091 VSS.n3340 VSS.n3083 22.9652
R5092 VSS.n2653 VSS.n2189 22.9652
R5093 VSS.n2692 VSS.n2691 22.9652
R5094 VSS.n2054 VSS.n2053 22.9652
R5095 VSS.n1979 VSS.n1978 22.9652
R5096 VSS.n1938 VSS.n1937 22.9652
R5097 VSS.n1830 VSS.n1442 22.9652
R5098 VSS.n1790 VSS.n1789 22.9652
R5099 VSS.n1737 VSS.n1490 22.9652
R5100 VSS.n1729 VSS.n1493 22.9652
R5101 VSS.n4923 VSS.n4922 22.9652
R5102 VSS.n5089 VSS.n250 22.9652
R5103 VSS.n1178 VSS.t194 22.6141
R5104 VSS.n1159 VSS.t196 22.6141
R5105 VSS.n4806 VSS.t2740 22.6141
R5106 VSS.n4636 VSS.t2734 22.6141
R5107 VSS.n4637 VSS.t2736 22.6141
R5108 VSS.n468 VSS.t2738 22.6141
R5109 VSS.n1160 VSS.t198 22.6141
R5110 VSS.n1165 VSS.t200 22.6141
R5111 VSS.n4009 VSS.n4008 22.5887
R5112 VSS.n2735 VSS.n2185 22.5887
R5113 VSS.n1084 VSS.n1035 22.5005
R5114 VSS.n1042 VSS.n1035 22.5005
R5115 VSS.n1034 VSS.n1032 22.5005
R5116 VSS.n1036 VSS.n1034 22.5005
R5117 VSS.n1072 VSS.n1071 22.5005
R5118 VSS.n1073 VSS.n1072 22.5005
R5119 VSS.n4984 VSS.n4983 22.5005
R5120 VSS.n4985 VSS.n4984 22.5005
R5121 VSS.n87 VSS.t1973 22.3257
R5122 VSS.n4184 VSS.t1346 22.3257
R5123 VSS.n4410 VSS.t746 22.3257
R5124 VSS.n2133 VSS.t2703 22.3257
R5125 VSS.n2137 VSS.t1976 22.3257
R5126 VSS.n3002 VSS.t1584 22.3257
R5127 VSS.n3436 VSS.t852 22.3257
R5128 VSS.n2276 VSS.t1260 22.3257
R5129 VSS.n1363 VSS.t855 22.3257
R5130 VSS.n1626 VSS.t1968 22.3257
R5131 VSS.n1836 VSS.t2617 22.3257
R5132 VSS.n1743 VSS.t1378 22.3257
R5133 VSS.n5255 VSS.t1751 22.3257
R5134 VSS.n4391 VSS.n4387 22.2496
R5135 VSS.n3647 VSS.n3646 22.2496
R5136 VSS.n3555 VSS.n3554 22.2496
R5137 VSS.n3532 VSS.n2997 22.2496
R5138 VSS.n3502 VSS.n3012 22.2496
R5139 VSS.n3494 VSS.n3014 22.2496
R5140 VSS.n962 VSS.n961 22.2123
R5141 VSS.n330 VSS.n329 22.2123
R5142 VSS.n337 VSS.n336 22.2123
R5143 VSS.n4540 VSS.n4538 22.2123
R5144 VSS.n4540 VSS.n4497 22.2123
R5145 VSS.n5575 VSS.n93 22.2123
R5146 VSS.n5575 VSS.n5574 22.2123
R5147 VSS.n5554 VSS.n104 22.2123
R5148 VSS.n5550 VSS.n104 22.2123
R5149 VSS.n5519 VSS.n5518 22.2123
R5150 VSS.n5518 VSS.n5517 22.2123
R5151 VSS.n5492 VSS.n129 22.2123
R5152 VSS.n5488 VSS.n129 22.2123
R5153 VSS.n5396 VSS.n5395 22.2123
R5154 VSS.n5390 VSS.n5389 22.2123
R5155 VSS.n5395 VSS.n5394 22.2123
R5156 VSS.n5389 VSS.n5388 22.2123
R5157 VSS.n5378 VSS.n5377 22.2123
R5158 VSS.n5377 VSS.n5376 22.2123
R5159 VSS.n3967 VSS.n3812 22.2123
R5160 VSS.n3968 VSS.n3967 22.2123
R5161 VSS.n4021 VSS.n3993 22.2123
R5162 VSS.n3569 VSS.n2979 22.2123
R5163 VSS.n3369 VSS.n3368 22.2123
R5164 VSS.n2508 VSS.n2507 22.2123
R5165 VSS.n1671 VSS.n1670 22.2123
R5166 VSS.n4816 VSS.n393 22.2123
R5167 VSS.n4820 VSS.n393 22.2123
R5168 VSS.n4867 VSS.n4865 22.2123
R5169 VSS.n4867 VSS.n373 22.2123
R5170 VSS.n4901 VSS.n4896 22.2123
R5171 VSS.n4897 VSS.n4896 22.2123
R5172 VSS.n5003 VSS.n5001 22.2123
R5173 VSS.n5004 VSS.n5003 22.2123
R5174 VSS.n5026 VSS.n278 22.2123
R5175 VSS.n5030 VSS.n278 22.2123
R5176 VSS.n5062 VSS.n5060 22.2123
R5177 VSS.n5063 VSS.n5062 22.2123
R5178 VSS.n5111 VSS.n241 22.2123
R5179 VSS.n5112 VSS.n5111 22.2123
R5180 VSS.n5176 VSS.n5124 22.2123
R5181 VSS.n5172 VSS.n5124 22.2123
R5182 VSS.n5152 VSS.n5151 22.2123
R5183 VSS.n5151 VSS.n5150 22.2123
R5184 VSS.n5198 VSS.n225 22.2123
R5185 VSS.n5199 VSS.n5198 22.2123
R5186 VSS.n5231 VSS.n5229 22.2123
R5187 VSS.n5231 VSS.n210 22.2123
R5188 VSS.n5268 VSS.n198 22.2123
R5189 VSS.n5269 VSS.n5268 22.2123
R5190 VSS.n5298 VSS.n187 22.2123
R5191 VSS.n5299 VSS.n5298 22.2123
R5192 VSS.n449 VSS.n397 22.2123
R5193 VSS.n449 VSS.n448 22.2123
R5194 VSS.n4036 VSS.n4035 21.8358
R5195 VSS.n4286 VSS.n3743 21.8358
R5196 VSS.n3582 VSS.n3581 21.8358
R5197 VSS.n3579 VSS.n3578 21.8358
R5198 VSS.n2008 VSS.n2007 21.8358
R5199 VSS.n1953 VSS.n1952 21.8358
R5200 VSS.n1937 VSS.n1391 21.8358
R5201 VSS.n1858 VSS.n1857 21.8358
R5202 VSS.n1801 VSS.n1457 21.8358
R5203 VSS.n1779 VSS.n1778 21.8358
R5204 VSS.n3085 VSS.t2076 21.795
R5205 VSS.n3456 VSS.n3031 21.6128
R5206 VSS.n4649 VSS.t2733 21.5216
R5207 VSS.t295 VSS.n1053 21.518
R5208 VSS.n4973 VSS.n4972 21.5165
R5209 VSS.n5506 VSS.n120 21.4593
R5210 VSS.n5494 VSS.n126 21.4593
R5211 VSS.n4064 VSS.n4062 21.4593
R5212 VSS.n4128 VSS.n3774 21.4593
R5213 VSS.n4160 VSS.n3764 21.4593
R5214 VSS.n4190 VSS.n3760 21.4593
R5215 VSS.n4244 VSS.n3758 21.4593
R5216 VSS.n4349 VSS.n4347 21.4593
R5217 VSS.n4360 VSS.n4359 21.4593
R5218 VSS.n4373 VSS.n4372 21.4593
R5219 VSS.n4405 VSS.n4404 21.4593
R5220 VSS.n4491 VSS.n4490 21.4593
R5221 VSS.n3684 VSS.n2130 21.4593
R5222 VSS.n3669 VSS.n3666 21.4593
R5223 VSS.n3637 VSS.n2944 21.4593
R5224 VSS.n3581 VSS.n3580 21.4593
R5225 VSS.n3563 VSS.n3562 21.4593
R5226 VSS.n3545 VSS.n2989 21.4593
R5227 VSS.n3543 VSS.n2991 21.4593
R5228 VSS.n3539 VSS.n3538 21.4593
R5229 VSS.n3504 VSS.n3503 21.4593
R5230 VSS.n3416 VSS.n3051 21.4593
R5231 VSS.n3344 VSS.n3083 21.4593
R5232 VSS.n3339 VSS.n3338 21.4593
R5233 VSS.n3318 VSS.n3092 21.4593
R5234 VSS.n2591 VSS.n2590 21.4593
R5235 VSS.n2537 VSS.n2244 21.4593
R5236 VSS.n2544 VSS.n2543 21.4593
R5237 VSS.n2499 VSS.n2498 21.4593
R5238 VSS.n2440 VSS.n2297 21.4593
R5239 VSS.n2730 VSS.n2660 21.4593
R5240 VSS.n2712 VSS.n2711 21.4593
R5241 VSS.n2692 VSS.n2680 21.4593
R5242 VSS.n2833 VSS.n2832 21.4593
R5243 VSS.n2828 VSS.n2827 21.4593
R5244 VSS.n2067 VSS.n1261 21.4593
R5245 VSS.n2054 VSS.n1334 21.4593
R5246 VSS.n2021 VSS.n2020 21.4593
R5247 VSS.n1978 VSS.n1977 21.4593
R5248 VSS.n1939 VSS.n1938 21.4593
R5249 VSS.n1904 VSS.n1902 21.4593
R5250 VSS.n1886 VSS.n1885 21.4593
R5251 VSS.n1834 VSS.n1442 21.4593
R5252 VSS.n1791 VSS.n1790 21.4593
R5253 VSS.n1741 VSS.n1490 21.4593
R5254 VSS.n1733 VSS.n1493 21.4593
R5255 VSS.n4924 VSS.n4923 21.4593
R5256 VSS.n5093 VSS.n250 21.4593
R5257 VSS.n2594 VSS.n2592 21.4593
R5258 VSS.n974 VSS.n973 21.3456
R5259 VSS.n1042 VSS.n1037 21.309
R5260 VSS.t2567 VSS.t1390 21.1843
R5261 VSS.t2569 VSS.t1388 21.1843
R5262 VSS.t2196 VSS.t2626 21.1843
R5263 VSS.t2198 VSS.t2624 21.1843
R5264 VSS.n4348 VSS.n3716 21.0829
R5265 VSS.n4625 VSS.t2666 20.8811
R5266 VSS.n1644 VSS.n1528 20.7295
R5267 VSS.n4195 VSS.n4194 20.7064
R5268 VSS.n3424 VSS.n3423 20.7064
R5269 VSS.n2818 VSS.n2812 20.7064
R5270 VSS.n1757 VSS.n1756 20.7064
R5271 VSS.n1666 VSS.n1517 20.7064
R5272 VSS.n2465 VSS.n2464 20.6347
R5273 VSS.n3961 VSS.n3960 20.3299
R5274 VSS.n4307 VSS.n3733 20.3299
R5275 VSS.n4418 VSS.n3691 20.3299
R5276 VSS.n3565 VSS.n3564 20.3299
R5277 VSS.n3431 VSS.n3430 20.3299
R5278 VSS.n3376 VSS.n3375 20.3299
R5279 VSS.n3259 VSS.n3258 20.3299
R5280 VSS.n2876 VSS.n2848 20.3299
R5281 VSS.n1971 VSS.n1374 20.3299
R5282 VSS.n1875 VSS.n1421 20.3299
R5283 VSS.n1819 VSS.n1818 20.3299
R5284 VSS.n1795 VSS.n1460 20.3299
R5285 VSS.n1664 VSS.n1663 20.3299
R5286 VSS.n4610 VSS.n4592 20.3039
R5287 VSS.n4608 VSS.n4604 20.3039
R5288 VSS.n983 VSS.n982 20.3039
R5289 VSS.n1220 VSS.n979 20.3039
R5290 VSS.n4985 VSS.t518 20.2139
R5291 VSS.n5765 VSS.n9 20.2009
R5292 VSS.n1074 VSS.t3088 20.1504
R5293 VSS.n4518 VSS.n4508 19.9534
R5294 VSS.n4546 VSS.n4495 19.9534
R5295 VSS.n5765 VSS.n5764 19.9534
R5296 VSS.n5731 VSS.n26 19.9534
R5297 VSS.n5692 VSS.n42 19.9534
R5298 VSS.n5674 VSS.n51 19.9534
R5299 VSS.n5641 VSS.n5640 19.9534
R5300 VSS.n5608 VSS.n5607 19.9534
R5301 VSS.n5581 VSS.n90 19.9534
R5302 VSS.n5511 VSS.n5510 19.9534
R5303 VSS.n5500 VSS.n123 19.9534
R5304 VSS.n5458 VSS.n144 19.9534
R5305 VSS.n5423 VSS.n5422 19.9534
R5306 VSS.n4042 VSS.n4041 19.9534
R5307 VSS.n4120 VSS.n3777 19.9534
R5308 VSS.n4209 VSS.n4179 19.9534
R5309 VSS.n4374 VSS.n4373 19.9534
R5310 VSS.n3243 VSS.n3242 19.9534
R5311 VSS.n2435 VSS.n2434 19.9534
R5312 VSS.n1845 VSS.n1844 19.9534
R5313 VSS.n5339 VSS.n5329 19.9534
R5314 VSS.n423 VSS.n413 19.9534
R5315 VSS.t2739 VSS.t68 19.9382
R5316 VSS.n4591 VSS.t987 19.9382
R5317 VSS.n5727 VSS.n26 19.914
R5318 VSS.n5640 VSS.n5639 19.914
R5319 VSS.n4341 VSS.n3718 19.914
R5320 VSS.n4599 VSS.n4597 19.8626
R5321 VSS.n1216 VSS.n1215 19.8626
R5322 VSS.n4527 VSS.n4503 19.577
R5323 VSS.n4533 VSS.n4500 19.577
R5324 VSS.n5384 VSS.n5383 19.577
R5325 VSS.n5372 VSS.n5371 19.577
R5326 VSS.n3858 VSS.n3857 19.577
R5327 VSS.n3877 VSS.n3874 19.577
R5328 VSS.n3945 VSS.n3818 19.577
R5329 VSS.n4013 VSS.n3999 19.577
R5330 VSS.n4065 VSS.n3802 19.577
R5331 VSS.n4093 VSS.n4092 19.577
R5332 VSS.n4448 VSS.n4442 19.577
R5333 VSS.n4454 VSS.n4438 19.577
R5334 VSS.n3374 VSS.n3069 19.577
R5335 VSS.n3370 VSS.n3369 19.577
R5336 VSS.n3153 VSS.n3135 19.577
R5337 VSS.n3145 VSS.n3139 19.577
R5338 VSS.n2095 VSS.n2085 19.577
R5339 VSS.n2101 VSS.n2081 19.577
R5340 VSS.n2615 VSS.n2614 19.577
R5341 VSS.n2545 VSS.n2237 19.577
R5342 VSS.n2466 VSS.n2281 19.577
R5343 VSS.n2362 VSS.n2361 19.577
R5344 VSS.n2354 VSS.n2353 19.577
R5345 VSS.n2347 VSS.n2346 19.577
R5346 VSS.n2862 VSS.n2859 19.577
R5347 VSS.n2870 VSS.n2867 19.577
R5348 VSS.n2786 VSS.n2785 19.577
R5349 VSS.n2819 VSS.n2818 19.577
R5350 VSS.n1824 VSS.n1823 19.577
R5351 VSS.n1686 VSS.n1685 19.577
R5352 VSS.n1582 VSS.n1581 19.577
R5353 VSS.n1574 VSS.n1573 19.577
R5354 VSS.n1567 VSS.n1566 19.577
R5355 VSS.n1284 VSS.n1278 19.577
R5356 VSS.n1290 VSS.n1274 19.577
R5357 VSS.n1298 VSS.n1270 19.577
R5358 VSS.n4829 VSS.n388 19.577
R5359 VSS.n4847 VSS.n4846 19.577
R5360 VSS.n4930 VSS.n4880 19.577
R5361 VSS.n4904 VSS.n4903 19.577
R5362 VSS.n5017 VSS.n5016 19.577
R5363 VSS.n5049 VSS.n5047 19.577
R5364 VSS.n5076 VSS.n5075 19.577
R5365 VSS.n5106 VSS.n5105 19.577
R5366 VSS.n5164 VSS.n5163 19.577
R5367 VSS.n5185 VSS.n232 19.577
R5368 VSS.n5216 VSS.n218 19.577
R5369 VSS.n5263 VSS.n5262 19.577
R5370 VSS.n5285 VSS.n5284 19.577
R5371 VSS.n5304 VSS.n185 19.577
R5372 VSS.n5313 VSS.n5312 19.577
R5373 VSS.n5320 VSS.n5319 19.577
R5374 VSS.n443 VSS.n401 19.577
R5375 VSS.n437 VSS.n404 19.577
R5376 VSS.n431 VSS.n407 19.577
R5377 VSS.n4599 VSS.n4598 19.4212
R5378 VSS.n1216 VSS.n987 19.4212
R5379 VSS.n4514 VSS.n4508 19.3355
R5380 VSS.n5335 VSS.n5329 19.3355
R5381 VSS.n419 VSS.n413 19.3355
R5382 VSS.n4267 VSS.n4266 19.2926
R5383 VSS.n4309 VSS.n4308 19.2926
R5384 VSS.n1674 VSS.n1671 19.2926
R5385 VSS.n4065 VSS.n4064 19.2005
R5386 VSS.n1652 VSS.n1651 19.2005
R5387 VSS.n2533 VSS.n2532 19.161
R5388 VSS.n983 VSS.n978 18.9798
R5389 VSS.n4996 VSS.t2841 18.9098
R5390 VSS.n3402 VSS.n3401 18.8449
R5391 VSS.n2364 VSS.n2363 18.824
R5392 VSS.n2002 VSS.n2001 18.824
R5393 VSS.n1947 VSS.n1946 18.824
R5394 VSS.n1932 VSS.n1931 18.824
R5395 VSS.n1896 VSS.n1895 18.824
R5396 VSS.n1796 VSS.n1795 18.824
R5397 VSS.n1773 VSS.n1772 18.824
R5398 VSS.n1753 VSS.n1484 18.824
R5399 VSS.n1688 VSS.n1687 18.824
R5400 VSS.n1637 VSS.n1636 18.824
R5401 VSS.n4609 VSS.n4608 18.7591
R5402 VSS.n1594 VSS.n1590 18.695
R5403 VSS.n5670 VSS.n51 18.5894
R5404 VSS.n3333 VSS.n3086 18.4476
R5405 VSS.n2450 VSS.n2449 18.4476
R5406 VSS.n2363 VSS.n2362 18.4476
R5407 VSS.n1582 VSS.n1549 18.4476
R5408 VSS.n4031 VSS.n3991 18.4197
R5409 VSS.n1627 VSS.n1625 18.1919
R5410 VSS.n5498 VSS.n126 18.0711
R5411 VSS.n4250 VSS.n4248 18.0711
R5412 VSS.n3634 VSS.n3633 18.0711
R5413 VSS.n2479 VSS.n2273 18.0711
R5414 VSS.n2440 VSS.n2439 18.0711
R5415 VSS.n1884 VSS.n1883 18.0711
R5416 VSS.n1852 VSS.n1851 18.0711
R5417 VSS.n1746 VSS.n1745 18.0711
R5418 VSS.n1173 VSS.n1172 17.9205
R5419 VSS.n4803 VSS.n4802 17.9205
R5420 VSS.n3314 VSS.n3092 17.8069
R5421 VSS.n2368 VSS.n2366 17.7867
R5422 VSS.n4970 VSS.t66 17.7035
R5423 VSS.n3220 VSS.n3219 17.7007
R5424 VSS.n3970 VSS.n3810 17.6946
R5425 VSS.n4391 VSS.n4390 17.6946
R5426 VSS.n3648 VSS.n3647 17.6946
R5427 VSS.n3556 VSS.n3555 17.6946
R5428 VSS.n3537 VSS.n2995 17.6946
R5429 VSS.n3250 VSS.n3249 17.6946
R5430 VSS.n2618 VSS.n2205 17.6946
R5431 VSS.n2034 VSS.n2033 17.6946
R5432 VSS.n2016 VSS.n1350 17.6946
R5433 VSS.n1962 VSS.n1961 17.6946
R5434 VSS.n1712 VSS.n1711 17.6946
R5435 VSS.n1653 VSS.n1524 17.6946
R5436 VSS.n5620 VSS.n5619 17.6577
R5437 VSS.n5530 VSS.n5528 17.6577
R5438 VSS.n5435 VSS.n5434 17.6577
R5439 VSS.n2751 VSS.n2750 17.6577
R5440 VSS.n5688 VSS.n42 17.3181
R5441 VSS.n5609 VSS.n5608 17.3181
R5442 VSS.n4272 VSS.n3748 17.3181
R5443 VSS.n3310 VSS.n3095 17.3181
R5444 VSS.n2366 VSS.n2365 17.3181
R5445 VSS.n2904 VSS.n2903 17.2527
R5446 VSS.n1100 VSS.n1099 17.1349
R5447 VSS.n1101 VSS.n1100 17.119
R5448 VSS.n2882 VSS.n2881 17.0835
R5449 VSS.n1172 VSS.n1171 17.0672
R5450 VSS.n4802 VSS.n4801 17.0672
R5451 VSS.n3287 VSS.n3286 16.9936
R5452 VSS.n3288 VSS.n3287 16.9936
R5453 VSS.n3280 VSS.n3109 16.9936
R5454 VSS.n3280 VSS.n3279 16.9936
R5455 VSS.n5506 VSS.n5505 16.9417
R5456 VSS.n4289 VSS.n3740 16.9417
R5457 VSS.n3417 VSS.n3416 16.9417
R5458 VSS.n3401 VSS.n3400 16.9417
R5459 VSS.n2832 VSS.n2803 16.9417
R5460 VSS.n1658 VSS.n1657 16.9417
R5461 VSS.t2190 VSS.t2652 16.8587
R5462 VSS.t42 VSS.t3181 16.8587
R5463 VSS.t1373 VSS.t3245 16.8587
R5464 VSS.t1546 VSS.t2714 16.8587
R5465 VSS.t482 VSS.t1793 16.8587
R5466 VSS.n3059 VSS.t1645 16.8587
R5467 VSS.t1486 VSS.t1701 16.8587
R5468 VSS.t1159 VSS.t1677 16.8587
R5469 VSS.t347 VSS.t1549 16.8587
R5470 VSS.t1170 VSS.t1673 16.8587
R5471 VSS.n4035 VSS.n3991 16.5652
R5472 VSS.n4491 VSS.n3691 16.5652
R5473 VSS.n2775 VSS.n2774 16.5522
R5474 VSS.n1302 VSS.n1270 16.5257
R5475 VSS.n1695 VSS.n1694 16.3238
R5476 VSS.t1114 VSS.t3054 16.1999
R5477 VSS.n1589 VSS.n1588 16.1887
R5478 VSS.n1062 VSS.n1061 16.1856
R5479 VSS.n1058 VSS.n301 16.1856
R5480 VSS.n304 VSS.n301 16.1856
R5481 VSS.n1137 VSS.t246 16.1734
R5482 VSS.n4667 VSS.t3286 16.1734
R5483 VSS.n1059 VSS.n1058 16.1529
R5484 VSS.t1847 VSS.t1499 16.1473
R5485 VSS.n4972 VSS.n350 16.126
R5486 VSS.n1061 VSS.n1060 16.0673
R5487 VSS.n5752 VSS.n14 15.8123
R5488 VSS.n5654 VSS.n5653 15.8123
R5489 VSS.n4282 VSS.n4281 15.8123
R5490 VSS.n2365 VSS.n2364 15.8123
R5491 VSS.n2003 VSS.n2002 15.8123
R5492 VSS.n1946 VSS.n1383 15.8123
R5493 VSS.n1933 VSS.n1932 15.8123
R5494 VSS.n1895 VSS.n1407 15.8123
R5495 VSS.n1853 VSS.n1852 15.8123
R5496 VSS.n1797 VSS.n1796 15.8123
R5497 VSS.n1774 VSS.n1773 15.8123
R5498 VSS.n1756 VSS.n1484 15.8123
R5499 VSS.n1747 VSS.n1746 15.8123
R5500 VSS.n1687 VSS.n1507 15.8123
R5501 VSS.n2434 VSS.n2433 15.7728
R5502 VSS.n5708 VSS.n5707 15.6833
R5503 VSS.n1926 VSS.n1925 15.5776
R5504 VSS.n1993 VSS.n1364 15.5708
R5505 VSS.n5206 VSS.n220 15.5279
R5506 VSS.n343 VSS.n342 15.4358
R5507 VSS.n4584 VSS.n4583 15.3963
R5508 VSS.n3332 VSS.n3330 15.3605
R5509 VSS.n4946 VSS.n4945 15.2301
R5510 VSS.n2585 VSS.n2219 15.2173
R5511 VSS.n5585 VSS.n90 15.1944
R5512 VSS.n5370 VSS.n5369 15.1944
R5513 VSS.n2492 VSS.n2491 15.1944
R5514 VSS.n4828 VSS.n4827 15.1944
R5515 VSS.n5046 VSS.n270 15.1944
R5516 VSS.n5289 VSS.n190 15.1944
R5517 VSS.n5462 VSS.n144 15.1514
R5518 VSS.n5218 VSS.n5217 15.1514
R5519 VSS.n966 VSS.n964 15.0593
R5520 VSS.n3346 VSS.n3345 15.0593
R5521 VSS.n3306 VSS.n3095 15.0593
R5522 VSS.n2447 VSS.n2446 15.0593
R5523 VSS.n1688 VSS.n1686 15.0593
R5524 VSS.n2561 VSS.n2560 14.9303
R5525 VSS.n5745 VSS.n5744 14.8179
R5526 VSS.n3870 VSS.n3868 14.8179
R5527 VSS.n3410 VSS.n3409 14.8179
R5528 VSS.n3228 VSS.n3133 14.8179
R5529 VSS.n5038 VSS.n273 14.8179
R5530 VSS.n5039 VSS.n5038 14.8179
R5531 VSS.n5275 VSS.n5274 14.8179
R5532 VSS.n5746 VSS.n5745 14.775
R5533 VSS.n5701 VSS.n5699 14.775
R5534 VSS.n5656 VSS.n5654 14.775
R5535 VSS.n5567 VSS.n99 14.775
R5536 VSS.n5563 VSS.n99 14.775
R5537 VSS.n4043 VSS.n4042 14.775
R5538 VSS.n3474 VSS.n3473 14.775
R5539 VSS.n2603 VSS.n2211 14.775
R5540 VSS.n2455 VSS.n2287 14.775
R5541 VSS.n2742 VSS.n2738 14.775
R5542 VSS.n4935 VSS.n370 14.775
R5543 VSS.n5224 VSS.n212 14.775
R5544 VSS.n4815 VSS.n460 14.775
R5545 VSS.n1082 VSS.n1081 14.7155
R5546 VSS.n1081 VSS.n1046 14.7155
R5547 VSS.n3681 VSS.n3680 14.6829
R5548 VSS.n3633 VSS.n3632 14.6829
R5549 VSS.n3443 VSS.n3442 14.6829
R5550 VSS.n1984 VSS.n1983 14.6829
R5551 VSS.n1967 VSS.n1966 14.6829
R5552 VSS.n1934 VSS.n1933 14.6829
R5553 VSS.n1883 VSS.n1882 14.6829
R5554 VSS.n1829 VSS.n1828 14.6829
R5555 VSS.n1804 VSS.n1454 14.6829
R5556 VSS.n1785 VSS.n1466 14.6829
R5557 VSS.n1728 VSS.n1727 14.6829
R5558 VSS.n1619 VSS.n1618 14.6829
R5559 VSS.n1590 VSS.n1589 14.6829
R5560 VSS.n3346 VSS.n3079 14.6388
R5561 VSS.n4941 VSS.t2633 14.4848
R5562 VSS.n2230 VSS.n2229 14.3889
R5563 VSS.t2837 VSS.t1699 14.3455
R5564 VSS.n2533 VSS.n2244 14.3064
R5565 VSS.n2000 VSS.n1999 14.3064
R5566 VSS.n1872 VSS.n1421 14.3064
R5567 VSS.n1792 VSS.n1460 14.3064
R5568 VSS.n3564 VSS.n3563 14.3064
R5569 VSS.n3430 VSS.n3429 14.3064
R5570 VSS.n3258 VSS.n3257 14.3064
R5571 VSS.n2049 VSS.n2048 14.3064
R5572 VSS.n1818 VSS.n1817 14.3064
R5573 VSS.n1663 VSS.n1662 14.3064
R5574 VSS.n2646 VSS.n2191 14.0717
R5575 VSS.n2067 VSS.n2066 14.022
R5576 VSS.n4019 VSS.n3996 13.9299
R5577 VSS.n4283 VSS.n4282 13.9299
R5578 VSS.n3320 VSS.n3319 13.9299
R5579 VSS.n3228 VSS.n3135 13.9299
R5580 VSS.n2494 VSS.n2265 13.9299
R5581 VSS.n2493 VSS.n2492 13.9299
R5582 VSS.n2356 VSS.n2354 13.9299
R5583 VSS.n1877 VSS.n1876 13.9299
R5584 VSS.n1576 VSS.n1574 13.9299
R5585 VSS.n936 VSS.n916 13.6992
R5586 VSS.n1135 VSS.n1134 13.6984
R5587 VSS.n1133 VSS.n1132 13.6984
R5588 VSS.n1131 VSS.n1130 13.6984
R5589 VSS.n1129 VSS.n1128 13.6984
R5590 VSS.n1127 VSS.n1126 13.6984
R5591 VSS.n1125 VSS.n1124 13.6984
R5592 VSS.n1123 VSS.n1122 13.6984
R5593 VSS.n935 VSS.n934 13.6984
R5594 VSS.n933 VSS.n932 13.6984
R5595 VSS.n931 VSS.n930 13.6984
R5596 VSS.n929 VSS.n928 13.6984
R5597 VSS.n927 VSS.n926 13.6984
R5598 VSS.n925 VSS.n924 13.6984
R5599 VSS.n4303 VSS.n3733 13.5534
R5600 VSS.n4349 VSS.n4348 13.5534
R5601 VSS.n1972 VSS.n1971 13.5534
R5602 VSS.n4088 VSS.n3792 13.3188
R5603 VSS.n5424 VSS.n5423 13.177
R5604 VSS.n5382 VSS.n5356 13.177
R5605 VSS.n3870 VSS.n3843 13.177
R5606 VSS.n2552 VSS.n2233 13.177
R5607 VSS.n2545 VSS.n2544 13.177
R5608 VSS.n2648 VSS.n2646 13.177
R5609 VSS.n2738 VSS.n2184 13.177
R5610 VSS.n1588 VSS.n1587 13.177
R5611 VSS.n5018 VSS.n283 13.177
R5612 VSS.n5077 VSS.n254 13.177
R5613 VSS.n5159 VSS.n5130 13.177
R5614 VSS.n5181 VSS.n5180 13.177
R5615 VSS.n5347 VSS.n178 13.177
R5616 VSS.n4957 VSS.n4956 12.8754
R5617 VSS.n4677 VSS.n4676 12.8005
R5618 VSS.n909 VSS.n908 12.8005
R5619 VSS.n5469 VSS.n5468 12.8005
R5620 VSS.n3945 VSS.n3944 12.8005
R5621 VSS.n3962 VSS.n3961 12.8005
R5622 VSS.n3689 VSS.n2069 12.8005
R5623 VSS.n3628 VSS.n2952 12.8005
R5624 VSS.n2449 VSS.n2448 12.8005
R5625 VSS.n2902 VSS.n2165 12.8005
R5626 VSS.n2048 VSS.n1337 12.8005
R5627 VSS.n2007 VSS.n2006 12.8005
R5628 VSS.n1952 VSS.n1951 12.8005
R5629 VSS.n1901 VSS.n1900 12.8005
R5630 VSS.n1857 VSS.n1856 12.8005
R5631 VSS.n1798 VSS.n1457 12.8005
R5632 VSS.n1778 VSS.n1777 12.8005
R5633 VSS.n1693 VSS.n1692 12.8005
R5634 VSS.n4104 VSS.n3785 12.5161
R5635 VSS.n2448 VSS.n2447 12.424
R5636 VSS.n2828 VSS.n2803 12.424
R5637 VSS.n1986 VSS.n1985 12.424
R5638 VSS.n4996 VSS.n4995 12.3894
R5639 VSS.n3895 VSS.n3894 12.3514
R5640 VSS.n2409 VSS.n2408 12.3514
R5641 VSS.n3895 VSS.n3836 12.1268
R5642 VSS.n2409 VSS.n2310 12.1268
R5643 VSS.n4037 VSS.n3986 12.0476
R5644 VSS.n4008 VSS.n4007 12.0476
R5645 VSS.n4244 VSS.n4242 12.0476
R5646 VSS.n2834 VSS.n2833 12.0476
R5647 VSS.n2774 VSS.n2172 11.9177
R5648 VSS.n4384 VSS.n4383 11.7085
R5649 VSS.n3643 VSS.n3642 11.7085
R5650 VSS.n3551 VSS.n3550 11.7085
R5651 VSS.n3528 VSS.n3525 11.7085
R5652 VSS.n3498 VSS.n3495 11.7085
R5653 VSS.n4092 VSS.n3792 11.6711
R5654 VSS.n3480 VSS.n3479 11.6711
R5655 VSS.n3320 VSS.n3088 11.6711
R5656 VSS.n2649 VSS.n2189 11.6711
R5657 VSS.n2592 VSS.n2591 11.2946
R5658 VSS.n2500 VSS.n2499 11.2946
R5659 VSS.n358 VSS.t2632 11.266
R5660 VSS.n1174 VSS.n1173 11.0072
R5661 VSS.n4804 VSS.n4803 11.0072
R5662 VSS.n3490 VSS.n3487 10.9555
R5663 VSS.n971 VSS.n970 10.9545
R5664 VSS.n4374 VSS.n3706 10.9181
R5665 VSS.n2552 VSS.n2551 10.9181
R5666 VSS.n2686 VSS.n2184 10.9181
R5667 VSS.n1878 VSS.n1877 10.9181
R5668 VSS.n4917 VSS.n4916 10.9181
R5669 VSS.n5083 VSS.n252 10.9181
R5670 VSS.n3578 VSS.n3577 10.8136
R5671 VSS.n2122 VSS.n2069 10.7135
R5672 VSS.n2629 VSS.n2627 10.7135
R5673 VSS.n3389 VSS.n3388 10.6338
R5674 VSS.n2707 VSS.n2671 10.6338
R5675 VSS.n1327 VSS.n1326 10.5983
R5676 VSS.n2123 VSS.n2122 10.5718
R5677 VSS.n969 VSS.n968 10.5541
R5678 VSS.n2627 VSS.n2201 10.5417
R5679 VSS.n2384 VSS.n2383 10.522
R5680 VSS.n2906 VSS.n2902 10.4353
R5681 VSS.n319 VSS.t1297 10.4216
R5682 VSS.n319 VSS.t1295 10.4216
R5683 VSS.n3403 VSS.n3402 10.2793
R5684 VSS.n1094 VSS.t2820 10.219
R5685 VSS.n4196 VSS.n4195 10.1652
R5686 VSS.n3423 VSS.n3422 10.1652
R5687 VSS.n2814 VSS.n2812 10.1652
R5688 VSS.n1902 VSS.n1901 10.1652
R5689 VSS.n1844 VSS.n1843 10.1652
R5690 VSS.n1843 VSS.n1842 10.1652
R5691 VSS.n1758 VSS.n1757 10.1652
R5692 VSS.n1638 VSS.n1637 10.1373
R5693 VSS.n1119 VSS.t2834 9.9005
R5694 VSS.n1119 VSS.t2959 9.9005
R5695 VSS.n921 VSS.t2981 9.9005
R5696 VSS.n921 VSS.t2900 9.9005
R5697 VSS.n4510 VSS.n4509 9.83768
R5698 VSS.n5367 VSS.n5364 9.83768
R5699 VSS.n5331 VSS.n5330 9.83768
R5700 VSS.n415 VSS.n414 9.83768
R5701 VSS.n4021 VSS.n4020 9.78874
R5702 VSS.n4002 VSS.n3999 9.78874
R5703 VSS.n4132 VSS.n4130 9.78874
R5704 VSS.n4155 VSS.n4154 9.78874
R5705 VSS.n4295 VSS.n4294 9.78874
R5706 VSS.n3635 VSS.n3634 9.78874
R5707 VSS.n3412 VSS.n3051 9.78874
R5708 VSS.n2656 VSS.n2655 9.78874
R5709 VSS.n1945 VSS.n1944 9.78874
R5710 VSS.n1885 VSS.n1884 9.78874
R5711 VSS.n1810 VSS.n1809 9.78874
R5712 VSS.n1767 VSS.n1766 9.78874
R5713 VSS.n973 VSS.n971 9.48661
R5714 VSS.n4656 VSS.t3469 9.43244
R5715 VSS.n5597 VSS.n5596 9.41227
R5716 VSS.n4215 VSS.n4214 9.41227
R5717 VSS.n4202 VSS.n4201 9.41227
R5718 VSS.n4281 VSS.n4280 9.41227
R5719 VSS.n4411 VSS.n4409 9.41227
R5720 VSS.n3674 VSS.n3673 9.41227
R5721 VSS.n3517 VSS.n3516 9.41227
R5722 VSS.n3438 VSS.n3437 9.41227
R5723 VSS.n1837 VSS.n1439 9.41227
R5724 VSS.n1694 VSS.n1693 9.41227
R5725 VSS.n5257 VSS.n5256 9.41227
R5726 VSS.t3244 VSS.t1026 9.34629
R5727 VSS.n968 VSS.n964 9.32264
R5728 VSS.n1172 VSS.n1166 9.3005
R5729 VSS.n963 VSS.n962 9.3005
R5730 VSS.n961 VSS.n958 9.3005
R5731 VSS.n336 VSS.n326 9.3005
R5732 VSS.n335 VSS.n334 9.3005
R5733 VSS.n333 VSS.n329 9.3005
R5734 VSS.n338 VSS.n337 9.3005
R5735 VSS.n343 VSS.n339 9.3005
R5736 VSS.n5367 VSS.n5366 9.3005
R5737 VSS.n5369 VSS.n5368 9.3005
R5738 VSS.n5370 VSS.n5362 9.3005
R5739 VSS.n5371 VSS.n5360 9.3005
R5740 VSS.n5373 VSS.n5372 9.3005
R5741 VSS.n5374 VSS.n5359 9.3005
R5742 VSS.n5376 VSS.n5375 9.3005
R5743 VSS.n5377 VSS.n5357 9.3005
R5744 VSS.n5379 VSS.n5378 9.3005
R5745 VSS.n5382 VSS.n5381 9.3005
R5746 VSS.n5383 VSS.n175 9.3005
R5747 VSS.n5385 VSS.n5384 9.3005
R5748 VSS.n5386 VSS.n174 9.3005
R5749 VSS.n5388 VSS.n5387 9.3005
R5750 VSS.n5389 VSS.n172 9.3005
R5751 VSS.n5391 VSS.n5390 9.3005
R5752 VSS.n5392 VSS.n171 9.3005
R5753 VSS.n5394 VSS.n5393 9.3005
R5754 VSS.n5395 VSS.n169 9.3005
R5755 VSS.n5396 VSS.n168 9.3005
R5756 VSS.n5399 VSS.n5398 9.3005
R5757 VSS.n5400 VSS.n167 9.3005
R5758 VSS.n5402 VSS.n5401 9.3005
R5759 VSS.n5403 VSS.n166 9.3005
R5760 VSS.n5405 VSS.n5404 9.3005
R5761 VSS.n5406 VSS.n165 9.3005
R5762 VSS.n5408 VSS.n5407 9.3005
R5763 VSS.n5409 VSS.n164 9.3005
R5764 VSS.n5412 VSS.n5411 9.3005
R5765 VSS.n5413 VSS.n163 9.3005
R5766 VSS.n5415 VSS.n5414 9.3005
R5767 VSS.n5417 VSS.n162 9.3005
R5768 VSS.n5419 VSS.n5418 9.3005
R5769 VSS.n5420 VSS.n161 9.3005
R5770 VSS.n5422 VSS.n5421 9.3005
R5771 VSS.n5423 VSS.n159 9.3005
R5772 VSS.n5424 VSS.n157 9.3005
R5773 VSS.n5425 VSS.n156 9.3005
R5774 VSS.n5428 VSS.n5427 9.3005
R5775 VSS.n5429 VSS.n155 9.3005
R5776 VSS.n5431 VSS.n5430 9.3005
R5777 VSS.n5434 VSS.n154 9.3005
R5778 VSS.n5436 VSS.n5435 9.3005
R5779 VSS.n5438 VSS.n5437 9.3005
R5780 VSS.n5439 VSS.n152 9.3005
R5781 VSS.n5441 VSS.n5440 9.3005
R5782 VSS.n5442 VSS.n151 9.3005
R5783 VSS.n5444 VSS.n5443 9.3005
R5784 VSS.n5445 VSS.n150 9.3005
R5785 VSS.n5447 VSS.n5446 9.3005
R5786 VSS.n5449 VSS.n5448 9.3005
R5787 VSS.n5450 VSS.n148 9.3005
R5788 VSS.n5453 VSS.n5452 9.3005
R5789 VSS.n5454 VSS.n147 9.3005
R5790 VSS.n5456 VSS.n5455 9.3005
R5791 VSS.n5457 VSS.n145 9.3005
R5792 VSS.n5459 VSS.n5458 9.3005
R5793 VSS.n5460 VSS.n144 9.3005
R5794 VSS.n5462 VSS.n5461 9.3005
R5795 VSS.n5464 VSS.n143 9.3005
R5796 VSS.n5466 VSS.n5465 9.3005
R5797 VSS.n5469 VSS.n137 9.3005
R5798 VSS.n5470 VSS.n136 9.3005
R5799 VSS.n5473 VSS.n5472 9.3005
R5800 VSS.n5474 VSS.n135 9.3005
R5801 VSS.n5476 VSS.n5475 9.3005
R5802 VSS.n5477 VSS.n134 9.3005
R5803 VSS.n5479 VSS.n5478 9.3005
R5804 VSS.n5482 VSS.n5481 9.3005
R5805 VSS.n5480 VSS.n131 9.3005
R5806 VSS.n5487 VSS.n130 9.3005
R5807 VSS.n5489 VSS.n5488 9.3005
R5808 VSS.n5490 VSS.n129 9.3005
R5809 VSS.n5492 VSS.n5491 9.3005
R5810 VSS.n5493 VSS.n127 9.3005
R5811 VSS.n5495 VSS.n5494 9.3005
R5812 VSS.n5496 VSS.n126 9.3005
R5813 VSS.n5498 VSS.n5497 9.3005
R5814 VSS.n5499 VSS.n124 9.3005
R5815 VSS.n5501 VSS.n5500 9.3005
R5816 VSS.n5502 VSS.n123 9.3005
R5817 VSS.n5504 VSS.n5503 9.3005
R5818 VSS.n5505 VSS.n121 9.3005
R5819 VSS.n5507 VSS.n5506 9.3005
R5820 VSS.n5508 VSS.n120 9.3005
R5821 VSS.n5510 VSS.n5509 9.3005
R5822 VSS.n5511 VSS.n118 9.3005
R5823 VSS.n5512 VSS.n117 9.3005
R5824 VSS.n5514 VSS.n5513 9.3005
R5825 VSS.n5515 VSS.n116 9.3005
R5826 VSS.n5517 VSS.n5516 9.3005
R5827 VSS.n5518 VSS.n114 9.3005
R5828 VSS.n5519 VSS.n113 9.3005
R5829 VSS.n5522 VSS.n5521 9.3005
R5830 VSS.n5523 VSS.n112 9.3005
R5831 VSS.n5525 VSS.n5524 9.3005
R5832 VSS.n5528 VSS.n111 9.3005
R5833 VSS.n5531 VSS.n5530 9.3005
R5834 VSS.n5532 VSS.n110 9.3005
R5835 VSS.n5534 VSS.n5533 9.3005
R5836 VSS.n5535 VSS.n109 9.3005
R5837 VSS.n5537 VSS.n5536 9.3005
R5838 VSS.n5538 VSS.n108 9.3005
R5839 VSS.n5540 VSS.n5539 9.3005
R5840 VSS.n5541 VSS.n107 9.3005
R5841 VSS.n5544 VSS.n5543 9.3005
R5842 VSS.n5545 VSS.n106 9.3005
R5843 VSS.n5547 VSS.n5546 9.3005
R5844 VSS.n5549 VSS.n105 9.3005
R5845 VSS.n5551 VSS.n5550 9.3005
R5846 VSS.n5552 VSS.n104 9.3005
R5847 VSS.n5554 VSS.n5553 9.3005
R5848 VSS.n5555 VSS.n102 9.3005
R5849 VSS.n5557 VSS.n5556 9.3005
R5850 VSS.n5559 VSS.n5558 9.3005
R5851 VSS.n5560 VSS.n100 9.3005
R5852 VSS.n5564 VSS.n5563 9.3005
R5853 VSS.n5565 VSS.n99 9.3005
R5854 VSS.n5567 VSS.n5566 9.3005
R5855 VSS.n5569 VSS.n98 9.3005
R5856 VSS.n5571 VSS.n5570 9.3005
R5857 VSS.n5574 VSS.n94 9.3005
R5858 VSS.n5576 VSS.n5575 9.3005
R5859 VSS.n5577 VSS.n93 9.3005
R5860 VSS.n5579 VSS.n5578 9.3005
R5861 VSS.n5580 VSS.n91 9.3005
R5862 VSS.n5582 VSS.n5581 9.3005
R5863 VSS.n5583 VSS.n90 9.3005
R5864 VSS.n5585 VSS.n5584 9.3005
R5865 VSS.n5587 VSS.n89 9.3005
R5866 VSS.n5591 VSS.n5590 9.3005
R5867 VSS.n5592 VSS.n88 9.3005
R5868 VSS.n5594 VSS.n5593 9.3005
R5869 VSS.n5595 VSS.n86 9.3005
R5870 VSS.n5598 VSS.n5597 9.3005
R5871 VSS.n5599 VSS.n85 9.3005
R5872 VSS.n5601 VSS.n5600 9.3005
R5873 VSS.n5602 VSS.n83 9.3005
R5874 VSS.n5604 VSS.n5603 9.3005
R5875 VSS.n5605 VSS.n82 9.3005
R5876 VSS.n5607 VSS.n5606 9.3005
R5877 VSS.n5608 VSS.n80 9.3005
R5878 VSS.n5609 VSS.n78 9.3005
R5879 VSS.n5610 VSS.n77 9.3005
R5880 VSS.n5613 VSS.n5612 9.3005
R5881 VSS.n5614 VSS.n76 9.3005
R5882 VSS.n5616 VSS.n5615 9.3005
R5883 VSS.n5619 VSS.n75 9.3005
R5884 VSS.n5621 VSS.n5620 9.3005
R5885 VSS.n5623 VSS.n5622 9.3005
R5886 VSS.n5624 VSS.n73 9.3005
R5887 VSS.n5626 VSS.n5625 9.3005
R5888 VSS.n5627 VSS.n72 9.3005
R5889 VSS.n5629 VSS.n5628 9.3005
R5890 VSS.n5630 VSS.n71 9.3005
R5891 VSS.n5632 VSS.n5631 9.3005
R5892 VSS.n5634 VSS.n5633 9.3005
R5893 VSS.n5635 VSS.n69 9.3005
R5894 VSS.n5637 VSS.n5636 9.3005
R5895 VSS.n5639 VSS.n5638 9.3005
R5896 VSS.n5640 VSS.n67 9.3005
R5897 VSS.n5642 VSS.n5641 9.3005
R5898 VSS.n5643 VSS.n66 9.3005
R5899 VSS.n5645 VSS.n5644 9.3005
R5900 VSS.n5646 VSS.n63 9.3005
R5901 VSS.n5647 VSS.n62 9.3005
R5902 VSS.n5649 VSS.n5648 9.3005
R5903 VSS.n5650 VSS.n61 9.3005
R5904 VSS.n5652 VSS.n5651 9.3005
R5905 VSS.n5653 VSS.n60 9.3005
R5906 VSS.n5654 VSS.n58 9.3005
R5907 VSS.n5657 VSS.n5656 9.3005
R5908 VSS.n5658 VSS.n57 9.3005
R5909 VSS.n5660 VSS.n5659 9.3005
R5910 VSS.n5661 VSS.n56 9.3005
R5911 VSS.n5663 VSS.n5662 9.3005
R5912 VSS.n5665 VSS.n5664 9.3005
R5913 VSS.n53 VSS.n52 9.3005
R5914 VSS.n5671 VSS.n5670 9.3005
R5915 VSS.n5672 VSS.n51 9.3005
R5916 VSS.n5674 VSS.n5673 9.3005
R5917 VSS.n5675 VSS.n49 9.3005
R5918 VSS.n5677 VSS.n5676 9.3005
R5919 VSS.n5678 VSS.n48 9.3005
R5920 VSS.n5680 VSS.n5679 9.3005
R5921 VSS.n5681 VSS.n46 9.3005
R5922 VSS.n5683 VSS.n5682 9.3005
R5923 VSS.n5685 VSS.n5684 9.3005
R5924 VSS.n5686 VSS.n43 9.3005
R5925 VSS.n5690 VSS.n42 9.3005
R5926 VSS.n5692 VSS.n5691 9.3005
R5927 VSS.n5693 VSS.n40 9.3005
R5928 VSS.n5695 VSS.n5694 9.3005
R5929 VSS.n5696 VSS.n39 9.3005
R5930 VSS.n5698 VSS.n5697 9.3005
R5931 VSS.n5699 VSS.n36 9.3005
R5932 VSS.n5702 VSS.n5701 9.3005
R5933 VSS.n5703 VSS.n35 9.3005
R5934 VSS.n5705 VSS.n5704 9.3005
R5935 VSS.n5709 VSS.n5708 9.3005
R5936 VSS.n5711 VSS.n5710 9.3005
R5937 VSS.n5712 VSS.n31 9.3005
R5938 VSS.n5714 VSS.n5713 9.3005
R5939 VSS.n5715 VSS.n30 9.3005
R5940 VSS.n5717 VSS.n5716 9.3005
R5941 VSS.n5718 VSS.n29 9.3005
R5942 VSS.n5721 VSS.n5720 9.3005
R5943 VSS.n5722 VSS.n28 9.3005
R5944 VSS.n5724 VSS.n5723 9.3005
R5945 VSS.n5725 VSS.n27 9.3005
R5946 VSS.n5728 VSS.n5727 9.3005
R5947 VSS.n5729 VSS.n26 9.3005
R5948 VSS.n5731 VSS.n5730 9.3005
R5949 VSS.n5732 VSS.n24 9.3005
R5950 VSS.n5734 VSS.n5733 9.3005
R5951 VSS.n5735 VSS.n23 9.3005
R5952 VSS.n5737 VSS.n5736 9.3005
R5953 VSS.n5738 VSS.n21 9.3005
R5954 VSS.n5742 VSS.n5741 9.3005
R5955 VSS.n5744 VSS.n5743 9.3005
R5956 VSS.n5745 VSS.n18 9.3005
R5957 VSS.n5747 VSS.n5746 9.3005
R5958 VSS.n5749 VSS.n5748 9.3005
R5959 VSS.n5750 VSS.n15 9.3005
R5960 VSS.n5754 VSS.n14 9.3005
R5961 VSS.n5756 VSS.n5755 9.3005
R5962 VSS.n5757 VSS.n13 9.3005
R5963 VSS.n5759 VSS.n5758 9.3005
R5964 VSS.n5760 VSS.n12 9.3005
R5965 VSS.n5762 VSS.n5761 9.3005
R5966 VSS.n5763 VSS.n5 9.3005
R5967 VSS.n5764 VSS.n6 9.3005
R5968 VSS.n5766 VSS.n5765 9.3005
R5969 VSS.n4565 VSS.n9 9.3005
R5970 VSS.n4567 VSS.n4566 9.3005
R5971 VSS.n4568 VSS.n4563 9.3005
R5972 VSS.n4570 VSS.n4569 9.3005
R5973 VSS.n4571 VSS.n4562 9.3005
R5974 VSS.n4573 VSS.n4572 9.3005
R5975 VSS.n4574 VSS.n4561 9.3005
R5976 VSS.n4576 VSS.n4575 9.3005
R5977 VSS.n4578 VSS.n4577 9.3005
R5978 VSS.n4579 VSS.n4559 9.3005
R5979 VSS.n4581 VSS.n4580 9.3005
R5980 VSS.n4583 VSS.n4582 9.3005
R5981 VSS.n4584 VSS.n4557 9.3005
R5982 VSS.n4556 VSS.n4493 9.3005
R5983 VSS.n4555 VSS.n4554 9.3005
R5984 VSS.n4552 VSS.n4494 9.3005
R5985 VSS.n4551 VSS.n4549 9.3005
R5986 VSS.n4548 VSS.n4495 9.3005
R5987 VSS.n4547 VSS.n4546 9.3005
R5988 VSS.n4545 VSS.n4496 9.3005
R5989 VSS.n4544 VSS.n4543 9.3005
R5990 VSS.n4542 VSS.n4497 9.3005
R5991 VSS.n4541 VSS.n4540 9.3005
R5992 VSS.n4538 VSS.n4498 9.3005
R5993 VSS.n4537 VSS.n4536 9.3005
R5994 VSS.n4535 VSS.n4500 9.3005
R5995 VSS.n4534 VSS.n4533 9.3005
R5996 VSS.n4532 VSS.n4501 9.3005
R5997 VSS.n4531 VSS.n4530 9.3005
R5998 VSS.n4529 VSS.n4503 9.3005
R5999 VSS.n4528 VSS.n4527 9.3005
R6000 VSS.n4526 VSS.n4504 9.3005
R6001 VSS.n4525 VSS.n4524 9.3005
R6002 VSS.n4523 VSS.n4506 9.3005
R6003 VSS.n4522 VSS.n4521 9.3005
R6004 VSS.n4520 VSS.n4507 9.3005
R6005 VSS.n4518 VSS.n4517 9.3005
R6006 VSS.n4516 VSS.n4508 9.3005
R6007 VSS.n4515 VSS.n4514 9.3005
R6008 VSS.n4512 VSS.n4509 9.3005
R6009 VSS.n5380 VSS.n5356 9.3005
R6010 VSS.n4469 VSS.n4468 9.3005
R6011 VSS.n4471 VSS.n4470 9.3005
R6012 VSS.n4472 VSS.n4430 9.3005
R6013 VSS.n4474 VSS.n4473 9.3005
R6014 VSS.n4476 VSS.n4475 9.3005
R6015 VSS.n4477 VSS.n4427 9.3005
R6016 VSS.n4479 VSS.n4478 9.3005
R6017 VSS.n4480 VSS.n4426 9.3005
R6018 VSS.n4466 VSS.n4432 9.3005
R6019 VSS.n4465 VSS.n4464 9.3005
R6020 VSS.n4463 VSS.n4462 9.3005
R6021 VSS.n4460 VSS.n4435 9.3005
R6022 VSS.n4456 VSS.n4438 9.3005
R6023 VSS.n4453 VSS.n4439 9.3005
R6024 VSS.n4450 VSS.n4442 9.3005
R6025 VSS.n4449 VSS.n4448 9.3005
R6026 VSS.n4452 VSS.n4451 9.3005
R6027 VSS.n4455 VSS.n4454 9.3005
R6028 VSS.n4458 VSS.n4457 9.3005
R6029 VSS.n4482 VSS.n4481 9.3005
R6030 VSS.n4485 VSS.n4424 9.3005
R6031 VSS.n4487 VSS.n4486 9.3005
R6032 VSS.n4488 VSS.n4423 9.3005
R6033 VSS.n3857 VSS.n3856 9.3005
R6034 VSS.n3858 VSS.n3849 9.3005
R6035 VSS.n3859 VSS.n3847 9.3005
R6036 VSS.n3862 VSS.n3861 9.3005
R6037 VSS.n3864 VSS.n3863 9.3005
R6038 VSS.n3868 VSS.n3844 9.3005
R6039 VSS.n3872 VSS.n3843 9.3005
R6040 VSS.n3874 VSS.n3873 9.3005
R6041 VSS.n3877 VSS.n3842 9.3005
R6042 VSS.n3879 VSS.n3878 9.3005
R6043 VSS.n3883 VSS.n3839 9.3005
R6044 VSS.n3886 VSS.n3885 9.3005
R6045 VSS.n3887 VSS.n3838 9.3005
R6046 VSS.n3889 VSS.n3888 9.3005
R6047 VSS.n3896 VSS.n3895 9.3005
R6048 VSS.n3898 VSS.n3897 9.3005
R6049 VSS.n3900 VSS.n3835 9.3005
R6050 VSS.n3902 VSS.n3901 9.3005
R6051 VSS.n3903 VSS.n3834 9.3005
R6052 VSS.n3905 VSS.n3904 9.3005
R6053 VSS.n3906 VSS.n3833 9.3005
R6054 VSS.n3908 VSS.n3907 9.3005
R6055 VSS.n3910 VSS.n3909 9.3005
R6056 VSS.n3912 VSS.n3831 9.3005
R6057 VSS.n3914 VSS.n3913 9.3005
R6058 VSS.n3916 VSS.n3915 9.3005
R6059 VSS.n3918 VSS.n3829 9.3005
R6060 VSS.n3919 VSS.n3827 9.3005
R6061 VSS.n3924 VSS.n3923 9.3005
R6062 VSS.n3925 VSS.n3826 9.3005
R6063 VSS.n3927 VSS.n3926 9.3005
R6064 VSS.n3929 VSS.n3824 9.3005
R6065 VSS.n3933 VSS.n3932 9.3005
R6066 VSS.n3936 VSS.n3935 9.3005
R6067 VSS.n3934 VSS.n3821 9.3005
R6068 VSS.n3820 VSS.n3819 9.3005
R6069 VSS.n3946 VSS.n3945 9.3005
R6070 VSS.n3947 VSS.n3818 9.3005
R6071 VSS.n3949 VSS.n3948 9.3005
R6072 VSS.n3950 VSS.n3817 9.3005
R6073 VSS.n3956 VSS.n3955 9.3005
R6074 VSS.n3957 VSS.n3816 9.3005
R6075 VSS.n3959 VSS.n3958 9.3005
R6076 VSS.n3960 VSS.n3814 9.3005
R6077 VSS.n3964 VSS.n3963 9.3005
R6078 VSS.n3965 VSS.n3812 9.3005
R6079 VSS.n3967 VSS.n3966 9.3005
R6080 VSS.n3968 VSS.n3811 9.3005
R6081 VSS.n3972 VSS.n3971 9.3005
R6082 VSS.n3973 VSS.n3810 9.3005
R6083 VSS.n3975 VSS.n3974 9.3005
R6084 VSS.n3976 VSS.n3809 9.3005
R6085 VSS.n3980 VSS.n3979 9.3005
R6086 VSS.n3981 VSS.n3807 9.3005
R6087 VSS.n4054 VSS.n4053 9.3005
R6088 VSS.n4052 VSS.n3808 9.3005
R6089 VSS.n4051 VSS.n4050 9.3005
R6090 VSS.n4048 VSS.n3982 9.3005
R6091 VSS.n4046 VSS.n4045 9.3005
R6092 VSS.n4044 VSS.n4043 9.3005
R6093 VSS.n4042 VSS.n3984 9.3005
R6094 VSS.n4041 VSS.n4040 9.3005
R6095 VSS.n4039 VSS.n3986 9.3005
R6096 VSS.n4038 VSS.n4037 9.3005
R6097 VSS.n4036 VSS.n3987 9.3005
R6098 VSS.n4035 VSS.n4034 9.3005
R6099 VSS.n4033 VSS.n3991 9.3005
R6100 VSS.n4032 VSS.n4031 9.3005
R6101 VSS.n4026 VSS.n3992 9.3005
R6102 VSS.n4025 VSS.n4024 9.3005
R6103 VSS.n4023 VSS.n3993 9.3005
R6104 VSS.n4022 VSS.n4021 9.3005
R6105 VSS.n4020 VSS.n3994 9.3005
R6106 VSS.n4019 VSS.n4018 9.3005
R6107 VSS.n4017 VSS.n3996 9.3005
R6108 VSS.n4016 VSS.n4015 9.3005
R6109 VSS.n4014 VSS.n3997 9.3005
R6110 VSS.n4013 VSS.n4012 9.3005
R6111 VSS.n4011 VSS.n4010 9.3005
R6112 VSS.n4009 VSS.n4000 9.3005
R6113 VSS.n4007 VSS.n4006 9.3005
R6114 VSS.n4005 VSS.n3806 9.3005
R6115 VSS.n4057 VSS.n3805 9.3005
R6116 VSS.n4059 VSS.n4058 9.3005
R6117 VSS.n4060 VSS.n3804 9.3005
R6118 VSS.n4062 VSS.n4061 9.3005
R6119 VSS.n4064 VSS.n3803 9.3005
R6120 VSS.n4066 VSS.n4065 9.3005
R6121 VSS.n4067 VSS.n3802 9.3005
R6122 VSS.n4069 VSS.n4068 9.3005
R6123 VSS.n4071 VSS.n3800 9.3005
R6124 VSS.n4074 VSS.n4073 9.3005
R6125 VSS.n4075 VSS.n3799 9.3005
R6126 VSS.n4077 VSS.n4076 9.3005
R6127 VSS.n4078 VSS.n3798 9.3005
R6128 VSS.n4081 VSS.n4080 9.3005
R6129 VSS.n4083 VSS.n4082 9.3005
R6130 VSS.n3795 VSS.n3794 9.3005
R6131 VSS.n4089 VSS.n4088 9.3005
R6132 VSS.n4090 VSS.n3792 9.3005
R6133 VSS.n4092 VSS.n4091 9.3005
R6134 VSS.n4093 VSS.n3790 9.3005
R6135 VSS.n4095 VSS.n4094 9.3005
R6136 VSS.n4097 VSS.n4096 9.3005
R6137 VSS.n4098 VSS.n3786 9.3005
R6138 VSS.n4101 VSS.n4100 9.3005
R6139 VSS.n4102 VSS.n3785 9.3005
R6140 VSS.n4104 VSS.n4103 9.3005
R6141 VSS.n4107 VSS.n3782 9.3005
R6142 VSS.n4110 VSS.n4109 9.3005
R6143 VSS.n4112 VSS.n4111 9.3005
R6144 VSS.n4113 VSS.n3779 9.3005
R6145 VSS.n4117 VSS.n4116 9.3005
R6146 VSS.n4118 VSS.n3777 9.3005
R6147 VSS.n4120 VSS.n4119 9.3005
R6148 VSS.n4121 VSS.n3776 9.3005
R6149 VSS.n4125 VSS.n4124 9.3005
R6150 VSS.n4126 VSS.n3774 9.3005
R6151 VSS.n4128 VSS.n4127 9.3005
R6152 VSS.n4129 VSS.n3772 9.3005
R6153 VSS.n4133 VSS.n4132 9.3005
R6154 VSS.n4134 VSS.n3771 9.3005
R6155 VSS.n4136 VSS.n4135 9.3005
R6156 VSS.n4137 VSS.n3770 9.3005
R6157 VSS.n4141 VSS.n4140 9.3005
R6158 VSS.n4142 VSS.n3769 9.3005
R6159 VSS.n4144 VSS.n4143 9.3005
R6160 VSS.n4147 VSS.n3768 9.3005
R6161 VSS.n4149 VSS.n4148 9.3005
R6162 VSS.n4150 VSS.n3767 9.3005
R6163 VSS.n4152 VSS.n4151 9.3005
R6164 VSS.n4154 VSS.n3765 9.3005
R6165 VSS.n4157 VSS.n4156 9.3005
R6166 VSS.n4158 VSS.n3764 9.3005
R6167 VSS.n4160 VSS.n4159 9.3005
R6168 VSS.n4161 VSS.n3762 9.3005
R6169 VSS.n4164 VSS.n4163 9.3005
R6170 VSS.n4165 VSS.n3761 9.3005
R6171 VSS.n4239 VSS.n4166 9.3005
R6172 VSS.n4238 VSS.n4237 9.3005
R6173 VSS.n4236 VSS.n4168 9.3005
R6174 VSS.n4235 VSS.n4234 9.3005
R6175 VSS.n4231 VSS.n4169 9.3005
R6176 VSS.n4230 VSS.n4229 9.3005
R6177 VSS.n4228 VSS.n4171 9.3005
R6178 VSS.n4227 VSS.n4226 9.3005
R6179 VSS.n4225 VSS.n4172 9.3005
R6180 VSS.n4221 VSS.n4220 9.3005
R6181 VSS.n4219 VSS.n4174 9.3005
R6182 VSS.n4218 VSS.n4217 9.3005
R6183 VSS.n4216 VSS.n4175 9.3005
R6184 VSS.n4213 VSS.n4212 9.3005
R6185 VSS.n4211 VSS.n4179 9.3005
R6186 VSS.n4210 VSS.n4209 9.3005
R6187 VSS.n4208 VSS.n4180 9.3005
R6188 VSS.n4207 VSS.n4206 9.3005
R6189 VSS.n4205 VSS.n4204 9.3005
R6190 VSS.n4203 VSS.n4183 9.3005
R6191 VSS.n4201 VSS.n4200 9.3005
R6192 VSS.n4199 VSS.n4185 9.3005
R6193 VSS.n4198 VSS.n4197 9.3005
R6194 VSS.n4196 VSS.n4186 9.3005
R6195 VSS.n4195 VSS.n4188 9.3005
R6196 VSS.n4194 VSS.n4193 9.3005
R6197 VSS.n4192 VSS.n4190 9.3005
R6198 VSS.n4191 VSS.n3760 9.3005
R6199 VSS.n4242 VSS.n3759 9.3005
R6200 VSS.n4245 VSS.n4244 9.3005
R6201 VSS.n4246 VSS.n3758 9.3005
R6202 VSS.n4248 VSS.n4247 9.3005
R6203 VSS.n4250 VSS.n3757 9.3005
R6204 VSS.n4252 VSS.n4251 9.3005
R6205 VSS.n4254 VSS.n4253 9.3005
R6206 VSS.n4255 VSS.n3755 9.3005
R6207 VSS.n4258 VSS.n4257 9.3005
R6208 VSS.n4260 VSS.n4259 9.3005
R6209 VSS.n4262 VSS.n3751 9.3005
R6210 VSS.n4264 VSS.n4263 9.3005
R6211 VSS.n4266 VSS.n4265 9.3005
R6212 VSS.n4267 VSS.n3749 9.3005
R6213 VSS.n4269 VSS.n4268 9.3005
R6214 VSS.n4270 VSS.n3748 9.3005
R6215 VSS.n4272 VSS.n4271 9.3005
R6216 VSS.n4273 VSS.n3746 9.3005
R6217 VSS.n4277 VSS.n4276 9.3005
R6218 VSS.n4278 VSS.n3745 9.3005
R6219 VSS.n4280 VSS.n4279 9.3005
R6220 VSS.n4282 VSS.n3744 9.3005
R6221 VSS.n4284 VSS.n4283 9.3005
R6222 VSS.n4286 VSS.n4285 9.3005
R6223 VSS.n4287 VSS.n3741 9.3005
R6224 VSS.n4290 VSS.n4289 9.3005
R6225 VSS.n4291 VSS.n3740 9.3005
R6226 VSS.n4293 VSS.n4292 9.3005
R6227 VSS.n4295 VSS.n3736 9.3005
R6228 VSS.n4297 VSS.n4296 9.3005
R6229 VSS.n4299 VSS.n4298 9.3005
R6230 VSS.n4302 VSS.n3734 9.3005
R6231 VSS.n4305 VSS.n4304 9.3005
R6232 VSS.n4307 VSS.n4306 9.3005
R6233 VSS.n4308 VSS.n3731 9.3005
R6234 VSS.n4310 VSS.n4309 9.3005
R6235 VSS.n4312 VSS.n4311 9.3005
R6236 VSS.n4313 VSS.n3729 9.3005
R6237 VSS.n4317 VSS.n4316 9.3005
R6238 VSS.n4319 VSS.n4318 9.3005
R6239 VSS.n4321 VSS.n3727 9.3005
R6240 VSS.n4323 VSS.n4322 9.3005
R6241 VSS.n4325 VSS.n4324 9.3005
R6242 VSS.n4326 VSS.n3724 9.3005
R6243 VSS.n4330 VSS.n4329 9.3005
R6244 VSS.n4332 VSS.n4331 9.3005
R6245 VSS.n4333 VSS.n3722 9.3005
R6246 VSS.n4336 VSS.n4335 9.3005
R6247 VSS.n4338 VSS.n4337 9.3005
R6248 VSS.n4339 VSS.n3719 9.3005
R6249 VSS.n4342 VSS.n4341 9.3005
R6250 VSS.n4343 VSS.n3718 9.3005
R6251 VSS.n4345 VSS.n4344 9.3005
R6252 VSS.n4347 VSS.n3717 9.3005
R6253 VSS.n4350 VSS.n4349 9.3005
R6254 VSS.n4351 VSS.n3716 9.3005
R6255 VSS.n4353 VSS.n4352 9.3005
R6256 VSS.n4355 VSS.n3713 9.3005
R6257 VSS.n4361 VSS.n4360 9.3005
R6258 VSS.n4362 VSS.n3712 9.3005
R6259 VSS.n4364 VSS.n4363 9.3005
R6260 VSS.n4365 VSS.n3710 9.3005
R6261 VSS.n4368 VSS.n4367 9.3005
R6262 VSS.n4369 VSS.n3708 9.3005
R6263 VSS.n4372 VSS.n4370 9.3005
R6264 VSS.n4373 VSS.n3707 9.3005
R6265 VSS.n4375 VSS.n4374 9.3005
R6266 VSS.n4376 VSS.n3706 9.3005
R6267 VSS.n4383 VSS.n4382 9.3005
R6268 VSS.n4377 VSS.n3705 9.3005
R6269 VSS.n4392 VSS.n4391 9.3005
R6270 VSS.n4389 VSS.n3699 9.3005
R6271 VSS.n4400 VSS.n3698 9.3005
R6272 VSS.n4402 VSS.n4401 9.3005
R6273 VSS.n4404 VSS.n3697 9.3005
R6274 VSS.n4406 VSS.n4405 9.3005
R6275 VSS.n4408 VSS.n4407 9.3005
R6276 VSS.n4409 VSS.n3694 9.3005
R6277 VSS.n4413 VSS.n4412 9.3005
R6278 VSS.n4414 VSS.n3693 9.3005
R6279 VSS.n4416 VSS.n4415 9.3005
R6280 VSS.n4417 VSS.n3692 9.3005
R6281 VSS.n4419 VSS.n4418 9.3005
R6282 VSS.n4420 VSS.n3691 9.3005
R6283 VSS.n4491 VSS.n4421 9.3005
R6284 VSS.n4490 VSS.n4489 9.3005
R6285 VSS.n3871 VSS.n3870 9.3005
R6286 VSS.n2101 VSS.n2100 9.3005
R6287 VSS.n2098 VSS.n2097 9.3005
R6288 VSS.n2095 VSS.n2093 9.3005
R6289 VSS.n2092 VSS.n2085 9.3005
R6290 VSS.n2096 VSS.n2084 9.3005
R6291 VSS.n2099 VSS.n2081 9.3005
R6292 VSS.n2102 VSS.n2079 9.3005
R6293 VSS.n2104 VSS.n2103 9.3005
R6294 VSS.n2106 VSS.n2105 9.3005
R6295 VSS.n2108 VSS.n2076 9.3005
R6296 VSS.n2110 VSS.n2109 9.3005
R6297 VSS.n2112 VSS.n2111 9.3005
R6298 VSS.n2114 VSS.n2074 9.3005
R6299 VSS.n2116 VSS.n2115 9.3005
R6300 VSS.n2118 VSS.n2117 9.3005
R6301 VSS.n2120 VSS.n2072 9.3005
R6302 VSS.n3146 VSS.n3145 9.3005
R6303 VSS.n3147 VSS.n3139 9.3005
R6304 VSS.n3149 VSS.n3148 9.3005
R6305 VSS.n3151 VSS.n3136 9.3005
R6306 VSS.n3154 VSS.n3153 9.3005
R6307 VSS.n3155 VSS.n3135 9.3005
R6308 VSS.n3226 VSS.n3133 9.3005
R6309 VSS.n3225 VSS.n3224 9.3005
R6310 VSS.n3220 VSS.n3156 9.3005
R6311 VSS.n3219 VSS.n3218 9.3005
R6312 VSS.n3217 VSS.n3216 9.3005
R6313 VSS.n3214 VSS.n3160 9.3005
R6314 VSS.n3212 VSS.n3211 9.3005
R6315 VSS.n3210 VSS.n3162 9.3005
R6316 VSS.n3209 VSS.n3208 9.3005
R6317 VSS.n3207 VSS.n3163 9.3005
R6318 VSS.n3206 VSS.n3205 9.3005
R6319 VSS.n3204 VSS.n3203 9.3005
R6320 VSS.n3202 VSS.n3166 9.3005
R6321 VSS.n3201 VSS.n3200 9.3005
R6322 VSS.n3199 VSS.n3198 9.3005
R6323 VSS.n3196 VSS.n3168 9.3005
R6324 VSS.n3194 VSS.n3193 9.3005
R6325 VSS.n3192 VSS.n3169 9.3005
R6326 VSS.n3191 VSS.n3190 9.3005
R6327 VSS.n3189 VSS.n3170 9.3005
R6328 VSS.n3187 VSS.n3186 9.3005
R6329 VSS.n3185 VSS.n3172 9.3005
R6330 VSS.n3184 VSS.n3183 9.3005
R6331 VSS.n3181 VSS.n3173 9.3005
R6332 VSS.n3180 VSS.n3179 9.3005
R6333 VSS.n3178 VSS.n3177 9.3005
R6334 VSS.n3175 VSS.n3132 9.3005
R6335 VSS.n3233 VSS.n3232 9.3005
R6336 VSS.n3235 VSS.n3234 9.3005
R6337 VSS.n3237 VSS.n3130 9.3005
R6338 VSS.n3240 VSS.n3239 9.3005
R6339 VSS.n3243 VSS.n3126 9.3005
R6340 VSS.n3245 VSS.n3244 9.3005
R6341 VSS.n3246 VSS.n3125 9.3005
R6342 VSS.n3248 VSS.n3247 9.3005
R6343 VSS.n3249 VSS.n3123 9.3005
R6344 VSS.n3252 VSS.n3251 9.3005
R6345 VSS.n3253 VSS.n3122 9.3005
R6346 VSS.n3255 VSS.n3254 9.3005
R6347 VSS.n3256 VSS.n3121 9.3005
R6348 VSS.n3257 VSS.n3119 9.3005
R6349 VSS.n3260 VSS.n3259 9.3005
R6350 VSS.n3262 VSS.n3261 9.3005
R6351 VSS.n3263 VSS.n3116 9.3005
R6352 VSS.n3265 VSS.n3264 9.3005
R6353 VSS.n3266 VSS.n3115 9.3005
R6354 VSS.n3268 VSS.n3267 9.3005
R6355 VSS.n3270 VSS.n3114 9.3005
R6356 VSS.n3273 VSS.n3272 9.3005
R6357 VSS.n3275 VSS.n3274 9.3005
R6358 VSS.n3277 VSS.n3108 9.3005
R6359 VSS.n3281 VSS.n3280 9.3005
R6360 VSS.n3282 VSS.n3107 9.3005
R6361 VSS.n3284 VSS.n3283 9.3005
R6362 VSS.n3287 VSS.n3104 9.3005
R6363 VSS.n3290 VSS.n3289 9.3005
R6364 VSS.n3292 VSS.n3291 9.3005
R6365 VSS.n3293 VSS.n3101 9.3005
R6366 VSS.n3297 VSS.n3296 9.3005
R6367 VSS.n3300 VSS.n3299 9.3005
R6368 VSS.n3298 VSS.n3097 9.3005
R6369 VSS.n3305 VSS.n3096 9.3005
R6370 VSS.n3308 VSS.n3307 9.3005
R6371 VSS.n3310 VSS.n3309 9.3005
R6372 VSS.n3311 VSS.n3093 9.3005
R6373 VSS.n3315 VSS.n3314 9.3005
R6374 VSS.n3316 VSS.n3092 9.3005
R6375 VSS.n3318 VSS.n3317 9.3005
R6376 VSS.n3319 VSS.n3089 9.3005
R6377 VSS.n3321 VSS.n3320 9.3005
R6378 VSS.n3322 VSS.n3088 9.3005
R6379 VSS.n3324 VSS.n3323 9.3005
R6380 VSS.n3325 VSS.n3087 9.3005
R6381 VSS.n3335 VSS.n3334 9.3005
R6382 VSS.n3336 VSS.n3086 9.3005
R6383 VSS.n3338 VSS.n3337 9.3005
R6384 VSS.n3339 VSS.n3084 9.3005
R6385 VSS.n3341 VSS.n3340 9.3005
R6386 VSS.n3342 VSS.n3083 9.3005
R6387 VSS.n3344 VSS.n3343 9.3005
R6388 VSS.n3345 VSS.n3080 9.3005
R6389 VSS.n3347 VSS.n3346 9.3005
R6390 VSS.n3349 VSS.n3348 9.3005
R6391 VSS.n3351 VSS.n3078 9.3005
R6392 VSS.n3353 VSS.n3352 9.3005
R6393 VSS.n3354 VSS.n3077 9.3005
R6394 VSS.n3356 VSS.n3355 9.3005
R6395 VSS.n3357 VSS.n3074 9.3005
R6396 VSS.n3364 VSS.n3363 9.3005
R6397 VSS.n3365 VSS.n3073 9.3005
R6398 VSS.n3367 VSS.n3366 9.3005
R6399 VSS.n3369 VSS.n3070 9.3005
R6400 VSS.n3371 VSS.n3370 9.3005
R6401 VSS.n3372 VSS.n3069 9.3005
R6402 VSS.n3374 VSS.n3373 9.3005
R6403 VSS.n3375 VSS.n3068 9.3005
R6404 VSS.n3377 VSS.n3376 9.3005
R6405 VSS.n3378 VSS.n3067 9.3005
R6406 VSS.n3380 VSS.n3379 9.3005
R6407 VSS.n3381 VSS.n3066 9.3005
R6408 VSS.n3385 VSS.n3384 9.3005
R6409 VSS.n3387 VSS.n3386 9.3005
R6410 VSS.n3388 VSS.n3063 9.3005
R6411 VSS.n3390 VSS.n3389 9.3005
R6412 VSS.n3392 VSS.n3391 9.3005
R6413 VSS.n3393 VSS.n3061 9.3005
R6414 VSS.n3397 VSS.n3396 9.3005
R6415 VSS.n3398 VSS.n3060 9.3005
R6416 VSS.n3400 VSS.n3399 9.3005
R6417 VSS.n3057 VSS.n3056 9.3005
R6418 VSS.n3407 VSS.n3406 9.3005
R6419 VSS.n3409 VSS.n3408 9.3005
R6420 VSS.n3410 VSS.n3054 9.3005
R6421 VSS.n3411 VSS.n3052 9.3005
R6422 VSS.n3413 VSS.n3412 9.3005
R6423 VSS.n3414 VSS.n3051 9.3005
R6424 VSS.n3416 VSS.n3415 9.3005
R6425 VSS.n3417 VSS.n3048 9.3005
R6426 VSS.n3419 VSS.n3418 9.3005
R6427 VSS.n3420 VSS.n3047 9.3005
R6428 VSS.n3422 VSS.n3421 9.3005
R6429 VSS.n3423 VSS.n3044 9.3005
R6430 VSS.n3425 VSS.n3424 9.3005
R6431 VSS.n3426 VSS.n3043 9.3005
R6432 VSS.n3428 VSS.n3427 9.3005
R6433 VSS.n3429 VSS.n3041 9.3005
R6434 VSS.n3432 VSS.n3431 9.3005
R6435 VSS.n3434 VSS.n3433 9.3005
R6436 VSS.n3435 VSS.n3038 9.3005
R6437 VSS.n3439 VSS.n3438 9.3005
R6438 VSS.n3440 VSS.n3037 9.3005
R6439 VSS.n3442 VSS.n3441 9.3005
R6440 VSS.n3443 VSS.n3036 9.3005
R6441 VSS.n3444 VSS.n3035 9.3005
R6442 VSS.n3450 VSS.n3449 9.3005
R6443 VSS.n3452 VSS.n3451 9.3005
R6444 VSS.n3453 VSS.n3032 9.3005
R6445 VSS.n3458 VSS.n3457 9.3005
R6446 VSS.n3459 VSS.n3031 9.3005
R6447 VSS.n3461 VSS.n3460 9.3005
R6448 VSS.n3463 VSS.n3028 9.3005
R6449 VSS.n3467 VSS.n3466 9.3005
R6450 VSS.n3468 VSS.n3027 9.3005
R6451 VSS.n3470 VSS.n3469 9.3005
R6452 VSS.n3473 VSS.n3026 9.3005
R6453 VSS.n3475 VSS.n3474 9.3005
R6454 VSS.n3476 VSS.n3025 9.3005
R6455 VSS.n3478 VSS.n3477 9.3005
R6456 VSS.n3479 VSS.n3024 9.3005
R6457 VSS.n3480 VSS.n3021 9.3005
R6458 VSS.n3481 VSS.n3019 9.3005
R6459 VSS.n3483 VSS.n3482 9.3005
R6460 VSS.n3485 VSS.n3484 9.3005
R6461 VSS.n3486 VSS.n3015 9.3005
R6462 VSS.n3492 VSS.n3491 9.3005
R6463 VSS.n3494 VSS.n3493 9.3005
R6464 VSS.n3495 VSS.n3013 9.3005
R6465 VSS.n3500 VSS.n3499 9.3005
R6466 VSS.n3502 VSS.n3501 9.3005
R6467 VSS.n3503 VSS.n3011 9.3005
R6468 VSS.n3504 VSS.n3009 9.3005
R6469 VSS.n3506 VSS.n3505 9.3005
R6470 VSS.n3508 VSS.n3507 9.3005
R6471 VSS.n3510 VSS.n3004 9.3005
R6472 VSS.n3513 VSS.n3512 9.3005
R6473 VSS.n3514 VSS.n3003 9.3005
R6474 VSS.n3516 VSS.n3515 9.3005
R6475 VSS.n3518 VSS.n3001 9.3005
R6476 VSS.n3520 VSS.n3519 9.3005
R6477 VSS.n3521 VSS.n3000 9.3005
R6478 VSS.n3523 VSS.n3522 9.3005
R6479 VSS.n3525 VSS.n2998 9.3005
R6480 VSS.n3530 VSS.n3529 9.3005
R6481 VSS.n3532 VSS.n3531 9.3005
R6482 VSS.n3533 VSS.n2996 9.3005
R6483 VSS.n3535 VSS.n3534 9.3005
R6484 VSS.n3537 VSS.n3536 9.3005
R6485 VSS.n3538 VSS.n2992 9.3005
R6486 VSS.n3540 VSS.n3539 9.3005
R6487 VSS.n3541 VSS.n2991 9.3005
R6488 VSS.n3543 VSS.n3542 9.3005
R6489 VSS.n3544 VSS.n2990 9.3005
R6490 VSS.n3546 VSS.n3545 9.3005
R6491 VSS.n3547 VSS.n2989 9.3005
R6492 VSS.n3550 VSS.n3549 9.3005
R6493 VSS.n3548 VSS.n2988 9.3005
R6494 VSS.n3555 VSS.n2986 9.3005
R6495 VSS.n3558 VSS.n3557 9.3005
R6496 VSS.n3559 VSS.n2985 9.3005
R6497 VSS.n3561 VSS.n3560 9.3005
R6498 VSS.n3562 VSS.n2984 9.3005
R6499 VSS.n3563 VSS.n2980 9.3005
R6500 VSS.n3566 VSS.n3565 9.3005
R6501 VSS.n3567 VSS.n2979 9.3005
R6502 VSS.n3569 VSS.n3568 9.3005
R6503 VSS.n3570 VSS.n2978 9.3005
R6504 VSS.n3575 VSS.n3574 9.3005
R6505 VSS.n3577 VSS.n3576 9.3005
R6506 VSS.n3578 VSS.n2976 9.3005
R6507 VSS.n3579 VSS.n2975 9.3005
R6508 VSS.n3580 VSS.n2973 9.3005
R6509 VSS.n3581 VSS.n2969 9.3005
R6510 VSS.n3585 VSS.n3584 9.3005
R6511 VSS.n3587 VSS.n3586 9.3005
R6512 VSS.n3590 VSS.n2967 9.3005
R6513 VSS.n3597 VSS.n3596 9.3005
R6514 VSS.n3598 VSS.n2966 9.3005
R6515 VSS.n3600 VSS.n3599 9.3005
R6516 VSS.n3602 VSS.n2965 9.3005
R6517 VSS.n3604 VSS.n3603 9.3005
R6518 VSS.n3607 VSS.n3606 9.3005
R6519 VSS.n3605 VSS.n2962 9.3005
R6520 VSS.n3613 VSS.n2960 9.3005
R6521 VSS.n3615 VSS.n3614 9.3005
R6522 VSS.n3616 VSS.n2959 9.3005
R6523 VSS.n3618 VSS.n3617 9.3005
R6524 VSS.n3621 VSS.n2957 9.3005
R6525 VSS.n3624 VSS.n3623 9.3005
R6526 VSS.n3626 VSS.n3625 9.3005
R6527 VSS.n3627 VSS.n2953 9.3005
R6528 VSS.n3629 VSS.n3628 9.3005
R6529 VSS.n3630 VSS.n2952 9.3005
R6530 VSS.n3632 VSS.n3631 9.3005
R6531 VSS.n3633 VSS.n2951 9.3005
R6532 VSS.n3634 VSS.n2949 9.3005
R6533 VSS.n3635 VSS.n2948 9.3005
R6534 VSS.n3636 VSS.n2945 9.3005
R6535 VSS.n3638 VSS.n3637 9.3005
R6536 VSS.n3639 VSS.n2944 9.3005
R6537 VSS.n3642 VSS.n3641 9.3005
R6538 VSS.n3640 VSS.n2943 9.3005
R6539 VSS.n3647 VSS.n2941 9.3005
R6540 VSS.n3650 VSS.n3649 9.3005
R6541 VSS.n3654 VSS.n2142 9.3005
R6542 VSS.n3665 VSS.n3664 9.3005
R6543 VSS.n3666 VSS.n2140 9.3005
R6544 VSS.n3670 VSS.n3669 9.3005
R6545 VSS.n3671 VSS.n2138 9.3005
R6546 VSS.n3673 VSS.n3672 9.3005
R6547 VSS.n3675 VSS.n2136 9.3005
R6548 VSS.n3677 VSS.n3676 9.3005
R6549 VSS.n3678 VSS.n2135 9.3005
R6550 VSS.n3680 VSS.n3679 9.3005
R6551 VSS.n3681 VSS.n2134 9.3005
R6552 VSS.n3683 VSS.n2131 9.3005
R6553 VSS.n3685 VSS.n3684 9.3005
R6554 VSS.n3686 VSS.n2130 9.3005
R6555 VSS.n3688 VSS.n3687 9.3005
R6556 VSS.n3689 VSS.n2129 9.3005
R6557 VSS.n2128 VSS.n2069 9.3005
R6558 VSS.n3228 VSS.n3227 9.3005
R6559 VSS.n2902 VSS.n2901 9.3005
R6560 VSS.n2899 VSS.n2898 9.3005
R6561 VSS.n2896 VSS.n2837 9.3005
R6562 VSS.n2895 VSS.n2894 9.3005
R6563 VSS.n2893 VSS.n2892 9.3005
R6564 VSS.n2890 VSS.n2840 9.3005
R6565 VSS.n2844 VSS.n2841 9.3005
R6566 VSS.n2881 VSS.n2845 9.3005
R6567 VSS.n2877 VSS.n2876 9.3005
R6568 VSS.n2871 VSS.n2870 9.3005
R6569 VSS.n2866 VSS.n2865 9.3005
R6570 VSS.n2863 VSS.n2862 9.3005
R6571 VSS.n2859 VSS.n2853 9.3005
R6572 VSS.n2864 VSS.n2852 9.3005
R6573 VSS.n2867 VSS.n2851 9.3005
R6574 VSS.n2872 VSS.n2850 9.3005
R6575 VSS.n2874 VSS.n2873 9.3005
R6576 VSS.n2875 VSS.n2849 9.3005
R6577 VSS.n2878 VSS.n2848 9.3005
R6578 VSS.n2880 VSS.n2879 9.3005
R6579 VSS.n2883 VSS.n2882 9.3005
R6580 VSS.n2885 VSS.n2884 9.3005
R6581 VSS.n2909 VSS.n2161 9.3005
R6582 VSS.n2912 VSS.n2911 9.3005
R6583 VSS.n2914 VSS.n2913 9.3005
R6584 VSS.n2915 VSS.n2159 9.3005
R6585 VSS.n2917 VSS.n2916 9.3005
R6586 VSS.n2918 VSS.n2158 9.3005
R6587 VSS.n2920 VSS.n2919 9.3005
R6588 VSS.n2922 VSS.n2156 9.3005
R6589 VSS.n2924 VSS.n2923 9.3005
R6590 VSS.n2926 VSS.n2925 9.3005
R6591 VSS.n2346 VSS.n2345 9.3005
R6592 VSS.n2347 VSS.n2338 9.3005
R6593 VSS.n2348 VSS.n2336 9.3005
R6594 VSS.n2351 VSS.n2350 9.3005
R6595 VSS.n2353 VSS.n2352 9.3005
R6596 VSS.n2354 VSS.n2334 9.3005
R6597 VSS.n2359 VSS.n2358 9.3005
R6598 VSS.n2361 VSS.n2360 9.3005
R6599 VSS.n2362 VSS.n2329 9.3005
R6600 VSS.n2363 VSS.n2328 9.3005
R6601 VSS.n2364 VSS.n2327 9.3005
R6602 VSS.n2365 VSS.n2326 9.3005
R6603 VSS.n2366 VSS.n2325 9.3005
R6604 VSS.n2369 VSS.n2368 9.3005
R6605 VSS.n2371 VSS.n2370 9.3005
R6606 VSS.n2373 VSS.n2323 9.3005
R6607 VSS.n2375 VSS.n2374 9.3005
R6608 VSS.n2377 VSS.n2376 9.3005
R6609 VSS.n2378 VSS.n2321 9.3005
R6610 VSS.n2381 VSS.n2380 9.3005
R6611 VSS.n2383 VSS.n2382 9.3005
R6612 VSS.n2390 VSS.n2389 9.3005
R6613 VSS.n2391 VSS.n2318 9.3005
R6614 VSS.n2393 VSS.n2392 9.3005
R6615 VSS.n2394 VSS.n2317 9.3005
R6616 VSS.n2396 VSS.n2395 9.3005
R6617 VSS.n2398 VSS.n2397 9.3005
R6618 VSS.n2399 VSS.n2315 9.3005
R6619 VSS.n2403 VSS.n2402 9.3005
R6620 VSS.n2404 VSS.n2314 9.3005
R6621 VSS.n2406 VSS.n2405 9.3005
R6622 VSS.n2407 VSS.n2311 9.3005
R6623 VSS.n2410 VSS.n2409 9.3005
R6624 VSS.n2412 VSS.n2411 9.3005
R6625 VSS.n2414 VSS.n2309 9.3005
R6626 VSS.n2418 VSS.n2417 9.3005
R6627 VSS.n2419 VSS.n2308 9.3005
R6628 VSS.n2421 VSS.n2420 9.3005
R6629 VSS.n2423 VSS.n2307 9.3005
R6630 VSS.n2425 VSS.n2424 9.3005
R6631 VSS.n2427 VSS.n2426 9.3005
R6632 VSS.n2429 VSS.n2304 9.3005
R6633 VSS.n2431 VSS.n2430 9.3005
R6634 VSS.n2433 VSS.n2432 9.3005
R6635 VSS.n2434 VSS.n2302 9.3005
R6636 VSS.n2436 VSS.n2435 9.3005
R6637 VSS.n2438 VSS.n2437 9.3005
R6638 VSS.n2439 VSS.n2298 9.3005
R6639 VSS.n2441 VSS.n2440 9.3005
R6640 VSS.n2442 VSS.n2297 9.3005
R6641 VSS.n2444 VSS.n2443 9.3005
R6642 VSS.n2445 VSS.n2296 9.3005
R6643 VSS.n2446 VSS.n2294 9.3005
R6644 VSS.n2447 VSS.n2293 9.3005
R6645 VSS.n2448 VSS.n2291 9.3005
R6646 VSS.n2449 VSS.n2290 9.3005
R6647 VSS.n2450 VSS.n2288 9.3005
R6648 VSS.n2452 VSS.n2451 9.3005
R6649 VSS.n2453 VSS.n2287 9.3005
R6650 VSS.n2455 VSS.n2454 9.3005
R6651 VSS.n2457 VSS.n2285 9.3005
R6652 VSS.n2461 VSS.n2460 9.3005
R6653 VSS.n2463 VSS.n2462 9.3005
R6654 VSS.n2465 VSS.n2282 9.3005
R6655 VSS.n2467 VSS.n2466 9.3005
R6656 VSS.n2468 VSS.n2281 9.3005
R6657 VSS.n2470 VSS.n2469 9.3005
R6658 VSS.n2472 VSS.n2279 9.3005
R6659 VSS.n2474 VSS.n2473 9.3005
R6660 VSS.n2476 VSS.n2475 9.3005
R6661 VSS.n2477 VSS.n2274 9.3005
R6662 VSS.n2480 VSS.n2479 9.3005
R6663 VSS.n2481 VSS.n2273 9.3005
R6664 VSS.n2483 VSS.n2482 9.3005
R6665 VSS.n2484 VSS.n2272 9.3005
R6666 VSS.n2485 VSS.n2271 9.3005
R6667 VSS.n2489 VSS.n2488 9.3005
R6668 VSS.n2491 VSS.n2490 9.3005
R6669 VSS.n2492 VSS.n2269 9.3005
R6670 VSS.n2493 VSS.n2266 9.3005
R6671 VSS.n2495 VSS.n2494 9.3005
R6672 VSS.n2496 VSS.n2265 9.3005
R6673 VSS.n2498 VSS.n2497 9.3005
R6674 VSS.n2499 VSS.n2264 9.3005
R6675 VSS.n2500 VSS.n2261 9.3005
R6676 VSS.n2501 VSS.n2256 9.3005
R6677 VSS.n2504 VSS.n2503 9.3005
R6678 VSS.n2505 VSS.n2255 9.3005
R6679 VSS.n2507 VSS.n2506 9.3005
R6680 VSS.n2253 VSS.n2252 9.3005
R6681 VSS.n2513 VSS.n2512 9.3005
R6682 VSS.n2514 VSS.n2251 9.3005
R6683 VSS.n2516 VSS.n2515 9.3005
R6684 VSS.n2517 VSS.n2250 9.3005
R6685 VSS.n2521 VSS.n2520 9.3005
R6686 VSS.n2522 VSS.n2249 9.3005
R6687 VSS.n2524 VSS.n2523 9.3005
R6688 VSS.n2526 VSS.n2248 9.3005
R6689 VSS.n2528 VSS.n2527 9.3005
R6690 VSS.n2530 VSS.n2529 9.3005
R6691 VSS.n2532 VSS.n2245 9.3005
R6692 VSS.n2534 VSS.n2533 9.3005
R6693 VSS.n2535 VSS.n2244 9.3005
R6694 VSS.n2537 VSS.n2536 9.3005
R6695 VSS.n2538 VSS.n2242 9.3005
R6696 VSS.n2540 VSS.n2539 9.3005
R6697 VSS.n2541 VSS.n2241 9.3005
R6698 VSS.n2543 VSS.n2542 9.3005
R6699 VSS.n2544 VSS.n2238 9.3005
R6700 VSS.n2546 VSS.n2545 9.3005
R6701 VSS.n2547 VSS.n2237 9.3005
R6702 VSS.n2549 VSS.n2548 9.3005
R6703 VSS.n2551 VSS.n2234 9.3005
R6704 VSS.n2553 VSS.n2552 9.3005
R6705 VSS.n2554 VSS.n2233 9.3005
R6706 VSS.n2556 VSS.n2555 9.3005
R6707 VSS.n2562 VSS.n2561 9.3005
R6708 VSS.n2564 VSS.n2563 9.3005
R6709 VSS.n2565 VSS.n2225 9.3005
R6710 VSS.n2568 VSS.n2567 9.3005
R6711 VSS.n2569 VSS.n2224 9.3005
R6712 VSS.n2571 VSS.n2570 9.3005
R6713 VSS.n2572 VSS.n2223 9.3005
R6714 VSS.n2577 VSS.n2576 9.3005
R6715 VSS.n2578 VSS.n2222 9.3005
R6716 VSS.n2580 VSS.n2579 9.3005
R6717 VSS.n2582 VSS.n2220 9.3005
R6718 VSS.n2587 VSS.n2586 9.3005
R6719 VSS.n2588 VSS.n2219 9.3005
R6720 VSS.n2590 VSS.n2589 9.3005
R6721 VSS.n2591 VSS.n2217 9.3005
R6722 VSS.n2592 VSS.n2215 9.3005
R6723 VSS.n2595 VSS.n2594 9.3005
R6724 VSS.n2597 VSS.n2596 9.3005
R6725 VSS.n2598 VSS.n2212 9.3005
R6726 VSS.n2600 VSS.n2599 9.3005
R6727 VSS.n2601 VSS.n2211 9.3005
R6728 VSS.n2603 VSS.n2602 9.3005
R6729 VSS.n2605 VSS.n2209 9.3005
R6730 VSS.n2610 VSS.n2609 9.3005
R6731 VSS.n2611 VSS.n2208 9.3005
R6732 VSS.n2613 VSS.n2612 9.3005
R6733 VSS.n2614 VSS.n2206 9.3005
R6734 VSS.n2616 VSS.n2615 9.3005
R6735 VSS.n2618 VSS.n2617 9.3005
R6736 VSS.n2620 VSS.n2202 9.3005
R6737 VSS.n2624 VSS.n2623 9.3005
R6738 VSS.n2625 VSS.n2201 9.3005
R6739 VSS.n2627 VSS.n2626 9.3005
R6740 VSS.n2633 VSS.n2632 9.3005
R6741 VSS.n2635 VSS.n2634 9.3005
R6742 VSS.n2638 VSS.n2192 9.3005
R6743 VSS.n2643 VSS.n2642 9.3005
R6744 VSS.n2644 VSS.n2191 9.3005
R6745 VSS.n2646 VSS.n2645 9.3005
R6746 VSS.n2648 VSS.n2190 9.3005
R6747 VSS.n2650 VSS.n2649 9.3005
R6748 VSS.n2651 VSS.n2189 9.3005
R6749 VSS.n2653 VSS.n2652 9.3005
R6750 VSS.n2654 VSS.n2186 9.3005
R6751 VSS.n2657 VSS.n2656 9.3005
R6752 VSS.n2735 VSS.n2658 9.3005
R6753 VSS.n2734 VSS.n2733 9.3005
R6754 VSS.n2732 VSS.n2660 9.3005
R6755 VSS.n2731 VSS.n2730 9.3005
R6756 VSS.n2728 VSS.n2661 9.3005
R6757 VSS.n2727 VSS.n2726 9.3005
R6758 VSS.n2725 VSS.n2663 9.3005
R6759 VSS.n2724 VSS.n2723 9.3005
R6760 VSS.n2722 VSS.n2664 9.3005
R6761 VSS.n2721 VSS.n2720 9.3005
R6762 VSS.n2719 VSS.n2718 9.3005
R6763 VSS.n2717 VSS.n2666 9.3005
R6764 VSS.n2672 VSS.n2668 9.3005
R6765 VSS.n2711 VSS.n2710 9.3005
R6766 VSS.n2709 VSS.n2671 9.3005
R6767 VSS.n2708 VSS.n2707 9.3005
R6768 VSS.n2705 VSS.n2673 9.3005
R6769 VSS.n2703 VSS.n2702 9.3005
R6770 VSS.n2701 VSS.n2700 9.3005
R6771 VSS.n2698 VSS.n2676 9.3005
R6772 VSS.n2696 VSS.n2695 9.3005
R6773 VSS.n2694 VSS.n2680 9.3005
R6774 VSS.n2693 VSS.n2692 9.3005
R6775 VSS.n2691 VSS.n2681 9.3005
R6776 VSS.n2690 VSS.n2689 9.3005
R6777 VSS.n2688 VSS.n2684 9.3005
R6778 VSS.n2687 VSS.n2686 9.3005
R6779 VSS.n2685 VSS.n2184 9.3005
R6780 VSS.n2738 VSS.n2183 9.3005
R6781 VSS.n2743 VSS.n2742 9.3005
R6782 VSS.n2744 VSS.n2182 9.3005
R6783 VSS.n2746 VSS.n2745 9.3005
R6784 VSS.n2750 VSS.n2181 9.3005
R6785 VSS.n2752 VSS.n2751 9.3005
R6786 VSS.n2754 VSS.n2753 9.3005
R6787 VSS.n2755 VSS.n2179 9.3005
R6788 VSS.n2757 VSS.n2756 9.3005
R6789 VSS.n2758 VSS.n2178 9.3005
R6790 VSS.n2760 VSS.n2759 9.3005
R6791 VSS.n2762 VSS.n2176 9.3005
R6792 VSS.n2766 VSS.n2765 9.3005
R6793 VSS.n2768 VSS.n2767 9.3005
R6794 VSS.n2769 VSS.n2173 9.3005
R6795 VSS.n2772 VSS.n2771 9.3005
R6796 VSS.n2774 VSS.n2773 9.3005
R6797 VSS.n2776 VSS.n2171 9.3005
R6798 VSS.n2781 VSS.n2780 9.3005
R6799 VSS.n2782 VSS.n2170 9.3005
R6800 VSS.n2785 VSS.n2783 9.3005
R6801 VSS.n2786 VSS.n2169 9.3005
R6802 VSS.n2791 VSS.n2790 9.3005
R6803 VSS.n2792 VSS.n2168 9.3005
R6804 VSS.n2794 VSS.n2793 9.3005
R6805 VSS.n2795 VSS.n2167 9.3005
R6806 VSS.n2797 VSS.n2796 9.3005
R6807 VSS.n2798 VSS.n2166 9.3005
R6808 VSS.n2834 VSS.n2799 9.3005
R6809 VSS.n2833 VSS.n2801 9.3005
R6810 VSS.n2832 VSS.n2831 9.3005
R6811 VSS.n2830 VSS.n2803 9.3005
R6812 VSS.n2829 VSS.n2828 9.3005
R6813 VSS.n2827 VSS.n2804 9.3005
R6814 VSS.n2824 VSS.n2823 9.3005
R6815 VSS.n2822 VSS.n2808 9.3005
R6816 VSS.n2821 VSS.n2820 9.3005
R6817 VSS.n2819 VSS.n2809 9.3005
R6818 VSS.n2818 VSS.n2817 9.3005
R6819 VSS.n2816 VSS.n2812 9.3005
R6820 VSS.n2815 VSS.n2814 9.3005
R6821 VSS.n2813 VSS.n2150 9.3005
R6822 VSS.n2154 VSS.n2151 9.3005
R6823 VSS.n2928 VSS.n2927 9.3005
R6824 VSS.n2356 VSS.n2332 9.3005
R6825 VSS.n1300 VSS.n1270 9.3005
R6826 VSS.n1296 VSS.n1271 9.3005
R6827 VSS.n1292 VSS.n1274 9.3005
R6828 VSS.n1289 VSS.n1275 9.3005
R6829 VSS.n1286 VSS.n1278 9.3005
R6830 VSS.n1285 VSS.n1284 9.3005
R6831 VSS.n1288 VSS.n1287 9.3005
R6832 VSS.n1291 VSS.n1290 9.3005
R6833 VSS.n1294 VSS.n1293 9.3005
R6834 VSS.n1299 VSS.n1298 9.3005
R6835 VSS.n1302 VSS.n1301 9.3005
R6836 VSS.n1304 VSS.n1268 9.3005
R6837 VSS.n1307 VSS.n1306 9.3005
R6838 VSS.n1309 VSS.n1308 9.3005
R6839 VSS.n1311 VSS.n1266 9.3005
R6840 VSS.n1314 VSS.n1313 9.3005
R6841 VSS.n1316 VSS.n1315 9.3005
R6842 VSS.n1317 VSS.n1264 9.3005
R6843 VSS.n1320 VSS.n1319 9.3005
R6844 VSS.n1321 VSS.n1263 9.3005
R6845 VSS.n1323 VSS.n1322 9.3005
R6846 VSS.n1325 VSS.n1262 9.3005
R6847 VSS.n1566 VSS.n1565 9.3005
R6848 VSS.n1567 VSS.n1558 9.3005
R6849 VSS.n1568 VSS.n1556 9.3005
R6850 VSS.n1571 VSS.n1570 9.3005
R6851 VSS.n1573 VSS.n1572 9.3005
R6852 VSS.n1574 VSS.n1553 9.3005
R6853 VSS.n1579 VSS.n1578 9.3005
R6854 VSS.n1581 VSS.n1550 9.3005
R6855 VSS.n1583 VSS.n1582 9.3005
R6856 VSS.n1584 VSS.n1549 9.3005
R6857 VSS.n1586 VSS.n1585 9.3005
R6858 VSS.n1587 VSS.n1547 9.3005
R6859 VSS.n1588 VSS.n1546 9.3005
R6860 VSS.n1589 VSS.n1545 9.3005
R6861 VSS.n1590 VSS.n1544 9.3005
R6862 VSS.n1595 VSS.n1594 9.3005
R6863 VSS.n1596 VSS.n1543 9.3005
R6864 VSS.n1598 VSS.n1597 9.3005
R6865 VSS.n1600 VSS.n1542 9.3005
R6866 VSS.n1603 VSS.n1602 9.3005
R6867 VSS.n1605 VSS.n1604 9.3005
R6868 VSS.n1606 VSS.n1540 9.3005
R6869 VSS.n1610 VSS.n1609 9.3005
R6870 VSS.n1611 VSS.n1539 9.3005
R6871 VSS.n1614 VSS.n1613 9.3005
R6872 VSS.n1619 VSS.n1536 9.3005
R6873 VSS.n1620 VSS.n1533 9.3005
R6874 VSS.n1622 VSS.n1621 9.3005
R6875 VSS.n1623 VSS.n1532 9.3005
R6876 VSS.n1625 VSS.n1624 9.3005
R6877 VSS.n1628 VSS.n1531 9.3005
R6878 VSS.n1633 VSS.n1632 9.3005
R6879 VSS.n1634 VSS.n1530 9.3005
R6880 VSS.n1636 VSS.n1635 9.3005
R6881 VSS.n1638 VSS.n1529 9.3005
R6882 VSS.n1646 VSS.n1645 9.3005
R6883 VSS.n1647 VSS.n1528 9.3005
R6884 VSS.n1649 VSS.n1648 9.3005
R6885 VSS.n1651 VSS.n1526 9.3005
R6886 VSS.n1652 VSS.n1525 9.3005
R6887 VSS.n1654 VSS.n1653 9.3005
R6888 VSS.n1656 VSS.n1655 9.3005
R6889 VSS.n1657 VSS.n1521 9.3005
R6890 VSS.n1659 VSS.n1658 9.3005
R6891 VSS.n1660 VSS.n1520 9.3005
R6892 VSS.n1662 VSS.n1661 9.3005
R6893 VSS.n1664 VSS.n1518 9.3005
R6894 VSS.n1667 VSS.n1666 9.3005
R6895 VSS.n1668 VSS.n1517 9.3005
R6896 VSS.n1670 VSS.n1669 9.3005
R6897 VSS.n1671 VSS.n1515 9.3005
R6898 VSS.n1675 VSS.n1674 9.3005
R6899 VSS.n1676 VSS.n1514 9.3005
R6900 VSS.n1678 VSS.n1677 9.3005
R6901 VSS.n1679 VSS.n1512 9.3005
R6902 VSS.n1682 VSS.n1681 9.3005
R6903 VSS.n1684 VSS.n1683 9.3005
R6904 VSS.n1685 VSS.n1508 9.3005
R6905 VSS.n1689 VSS.n1688 9.3005
R6906 VSS.n1690 VSS.n1507 9.3005
R6907 VSS.n1692 VSS.n1691 9.3005
R6908 VSS.n1694 VSS.n1505 9.3005
R6909 VSS.n1695 VSS.n1504 9.3005
R6910 VSS.n1700 VSS.n1699 9.3005
R6911 VSS.n1702 VSS.n1701 9.3005
R6912 VSS.n1703 VSS.n1501 9.3005
R6913 VSS.n1707 VSS.n1706 9.3005
R6914 VSS.n1708 VSS.n1500 9.3005
R6915 VSS.n1710 VSS.n1709 9.3005
R6916 VSS.n1711 VSS.n1498 9.3005
R6917 VSS.n1716 VSS.n1715 9.3005
R6918 VSS.n1717 VSS.n1497 9.3005
R6919 VSS.n1719 VSS.n1718 9.3005
R6920 VSS.n1720 VSS.n1496 9.3005
R6921 VSS.n1724 VSS.n1723 9.3005
R6922 VSS.n1725 VSS.n1495 9.3005
R6923 VSS.n1727 VSS.n1726 9.3005
R6924 VSS.n1728 VSS.n1494 9.3005
R6925 VSS.n1730 VSS.n1729 9.3005
R6926 VSS.n1731 VSS.n1493 9.3005
R6927 VSS.n1733 VSS.n1732 9.3005
R6928 VSS.n1736 VSS.n1491 9.3005
R6929 VSS.n1738 VSS.n1737 9.3005
R6930 VSS.n1739 VSS.n1490 9.3005
R6931 VSS.n1741 VSS.n1740 9.3005
R6932 VSS.n1742 VSS.n1487 9.3005
R6933 VSS.n1748 VSS.n1747 9.3005
R6934 VSS.n1749 VSS.n1486 9.3005
R6935 VSS.n1751 VSS.n1750 9.3005
R6936 VSS.n1752 VSS.n1485 9.3005
R6937 VSS.n1754 VSS.n1753 9.3005
R6938 VSS.n1756 VSS.n1755 9.3005
R6939 VSS.n1757 VSS.n1482 9.3005
R6940 VSS.n1758 VSS.n1480 9.3005
R6941 VSS.n1761 VSS.n1760 9.3005
R6942 VSS.n1762 VSS.n1479 9.3005
R6943 VSS.n1764 VSS.n1763 9.3005
R6944 VSS.n1765 VSS.n1477 9.3005
R6945 VSS.n1768 VSS.n1767 9.3005
R6946 VSS.n1770 VSS.n1769 9.3005
R6947 VSS.n1771 VSS.n1474 9.3005
R6948 VSS.n1772 VSS.n1473 9.3005
R6949 VSS.n1775 VSS.n1774 9.3005
R6950 VSS.n1777 VSS.n1776 9.3005
R6951 VSS.n1779 VSS.n1469 9.3005
R6952 VSS.n1781 VSS.n1780 9.3005
R6953 VSS.n1783 VSS.n1782 9.3005
R6954 VSS.n1784 VSS.n1467 9.3005
R6955 VSS.n1786 VSS.n1785 9.3005
R6956 VSS.n1787 VSS.n1466 9.3005
R6957 VSS.n1789 VSS.n1788 9.3005
R6958 VSS.n1790 VSS.n1463 9.3005
R6959 VSS.n1791 VSS.n1461 9.3005
R6960 VSS.n1793 VSS.n1792 9.3005
R6961 VSS.n1795 VSS.n1794 9.3005
R6962 VSS.n1797 VSS.n1458 9.3005
R6963 VSS.n1799 VSS.n1798 9.3005
R6964 VSS.n1801 VSS.n1800 9.3005
R6965 VSS.n1802 VSS.n1455 9.3005
R6966 VSS.n1805 VSS.n1804 9.3005
R6967 VSS.n1806 VSS.n1454 9.3005
R6968 VSS.n1808 VSS.n1807 9.3005
R6969 VSS.n1810 VSS.n1451 9.3005
R6970 VSS.n1813 VSS.n1812 9.3005
R6971 VSS.n1814 VSS.n1450 9.3005
R6972 VSS.n1816 VSS.n1815 9.3005
R6973 VSS.n1817 VSS.n1448 9.3005
R6974 VSS.n1820 VSS.n1819 9.3005
R6975 VSS.n1822 VSS.n1821 9.3005
R6976 VSS.n1823 VSS.n1445 9.3005
R6977 VSS.n1825 VSS.n1824 9.3005
R6978 VSS.n1826 VSS.n1444 9.3005
R6979 VSS.n1828 VSS.n1827 9.3005
R6980 VSS.n1829 VSS.n1443 9.3005
R6981 VSS.n1831 VSS.n1830 9.3005
R6982 VSS.n1832 VSS.n1442 9.3005
R6983 VSS.n1834 VSS.n1833 9.3005
R6984 VSS.n1835 VSS.n1440 9.3005
R6985 VSS.n1839 VSS.n1838 9.3005
R6986 VSS.n1840 VSS.n1439 9.3005
R6987 VSS.n1842 VSS.n1841 9.3005
R6988 VSS.n1843 VSS.n1437 9.3005
R6989 VSS.n1844 VSS.n1435 9.3005
R6990 VSS.n1846 VSS.n1845 9.3005
R6991 VSS.n1847 VSS.n1434 9.3005
R6992 VSS.n1849 VSS.n1848 9.3005
R6993 VSS.n1850 VSS.n1431 9.3005
R6994 VSS.n1854 VSS.n1853 9.3005
R6995 VSS.n1856 VSS.n1855 9.3005
R6996 VSS.n1858 VSS.n1428 9.3005
R6997 VSS.n1860 VSS.n1859 9.3005
R6998 VSS.n1862 VSS.n1861 9.3005
R6999 VSS.n1863 VSS.n1426 9.3005
R7000 VSS.n1866 VSS.n1865 9.3005
R7001 VSS.n1868 VSS.n1867 9.3005
R7002 VSS.n1873 VSS.n1872 9.3005
R7003 VSS.n1875 VSS.n1874 9.3005
R7004 VSS.n1876 VSS.n1419 9.3005
R7005 VSS.n1877 VSS.n1418 9.3005
R7006 VSS.n1879 VSS.n1878 9.3005
R7007 VSS.n1880 VSS.n1417 9.3005
R7008 VSS.n1882 VSS.n1881 9.3005
R7009 VSS.n1883 VSS.n1416 9.3005
R7010 VSS.n1884 VSS.n1414 9.3005
R7011 VSS.n1885 VSS.n1413 9.3005
R7012 VSS.n1886 VSS.n1410 9.3005
R7013 VSS.n1888 VSS.n1887 9.3005
R7014 VSS.n1890 VSS.n1889 9.3005
R7015 VSS.n1894 VSS.n1408 9.3005
R7016 VSS.n1897 VSS.n1896 9.3005
R7017 VSS.n1898 VSS.n1407 9.3005
R7018 VSS.n1900 VSS.n1899 9.3005
R7019 VSS.n1902 VSS.n1404 9.3005
R7020 VSS.n1905 VSS.n1904 9.3005
R7021 VSS.n1906 VSS.n1403 9.3005
R7022 VSS.n1908 VSS.n1907 9.3005
R7023 VSS.n1910 VSS.n1401 9.3005
R7024 VSS.n1913 VSS.n1912 9.3005
R7025 VSS.n1914 VSS.n1400 9.3005
R7026 VSS.n1916 VSS.n1915 9.3005
R7027 VSS.n1917 VSS.n1396 9.3005
R7028 VSS.n1923 VSS.n1922 9.3005
R7029 VSS.n1925 VSS.n1924 9.3005
R7030 VSS.n1926 VSS.n1394 9.3005
R7031 VSS.n1928 VSS.n1927 9.3005
R7032 VSS.n1929 VSS.n1393 9.3005
R7033 VSS.n1931 VSS.n1930 9.3005
R7034 VSS.n1933 VSS.n1392 9.3005
R7035 VSS.n1935 VSS.n1934 9.3005
R7036 VSS.n1937 VSS.n1936 9.3005
R7037 VSS.n1938 VSS.n1388 9.3005
R7038 VSS.n1940 VSS.n1939 9.3005
R7039 VSS.n1941 VSS.n1387 9.3005
R7040 VSS.n1943 VSS.n1942 9.3005
R7041 VSS.n1945 VSS.n1384 9.3005
R7042 VSS.n1948 VSS.n1947 9.3005
R7043 VSS.n1949 VSS.n1383 9.3005
R7044 VSS.n1951 VSS.n1950 9.3005
R7045 VSS.n1953 VSS.n1380 9.3005
R7046 VSS.n1956 VSS.n1955 9.3005
R7047 VSS.n1958 VSS.n1957 9.3005
R7048 VSS.n1959 VSS.n1378 9.3005
R7049 VSS.n1963 VSS.n1962 9.3005
R7050 VSS.n1964 VSS.n1377 9.3005
R7051 VSS.n1966 VSS.n1965 9.3005
R7052 VSS.n1967 VSS.n1376 9.3005
R7053 VSS.n1968 VSS.n1375 9.3005
R7054 VSS.n1974 VSS.n1973 9.3005
R7055 VSS.n1975 VSS.n1374 9.3005
R7056 VSS.n1977 VSS.n1976 9.3005
R7057 VSS.n1978 VSS.n1372 9.3005
R7058 VSS.n1980 VSS.n1979 9.3005
R7059 VSS.n1981 VSS.n1371 9.3005
R7060 VSS.n1983 VSS.n1982 9.3005
R7061 VSS.n1984 VSS.n1370 9.3005
R7062 VSS.n1985 VSS.n1369 9.3005
R7063 VSS.n1368 VSS.n1366 9.3005
R7064 VSS.n1990 VSS.n1365 9.3005
R7065 VSS.n1994 VSS.n1993 9.3005
R7066 VSS.n1995 VSS.n1364 9.3005
R7067 VSS.n1997 VSS.n1996 9.3005
R7068 VSS.n1999 VSS.n1362 9.3005
R7069 VSS.n2000 VSS.n1360 9.3005
R7070 VSS.n2001 VSS.n1359 9.3005
R7071 VSS.n2004 VSS.n2003 9.3005
R7072 VSS.n2006 VSS.n2005 9.3005
R7073 VSS.n2008 VSS.n1354 9.3005
R7074 VSS.n2011 VSS.n2010 9.3005
R7075 VSS.n2013 VSS.n2012 9.3005
R7076 VSS.n2015 VSS.n1351 9.3005
R7077 VSS.n2017 VSS.n2016 9.3005
R7078 VSS.n2019 VSS.n2018 9.3005
R7079 VSS.n2020 VSS.n1348 9.3005
R7080 VSS.n2022 VSS.n2021 9.3005
R7081 VSS.n2023 VSS.n1347 9.3005
R7082 VSS.n2029 VSS.n2028 9.3005
R7083 VSS.n2035 VSS.n2034 9.3005
R7084 VSS.n2031 VSS.n1340 9.3005
R7085 VSS.n2043 VSS.n1339 9.3005
R7086 VSS.n2045 VSS.n2044 9.3005
R7087 VSS.n2046 VSS.n1338 9.3005
R7088 VSS.n2050 VSS.n2049 9.3005
R7089 VSS.n2052 VSS.n2051 9.3005
R7090 VSS.n2053 VSS.n1335 9.3005
R7091 VSS.n2055 VSS.n2054 9.3005
R7092 VSS.n2056 VSS.n1334 9.3005
R7093 VSS.n2058 VSS.n2057 9.3005
R7094 VSS.n2060 VSS.n1333 9.3005
R7095 VSS.n2064 VSS.n2063 9.3005
R7096 VSS.n2066 VSS.n2065 9.3005
R7097 VSS.n2067 VSS.n1330 9.3005
R7098 VSS.n1329 VSS.n1261 9.3005
R7099 VSS.n1328 VSS.n1327 9.3005
R7100 VSS.n1577 VSS.n1576 9.3005
R7101 VSS.n417 VSS.n414 9.3005
R7102 VSS.n420 VSS.n419 9.3005
R7103 VSS.n5333 VSS.n5330 9.3005
R7104 VSS.n5336 VSS.n5335 9.3005
R7105 VSS.n5337 VSS.n5329 9.3005
R7106 VSS.n5339 VSS.n5338 9.3005
R7107 VSS.n5340 VSS.n5328 9.3005
R7108 VSS.n5341 VSS.n5325 9.3005
R7109 VSS.n5343 VSS.n5342 9.3005
R7110 VSS.n5344 VSS.n5324 9.3005
R7111 VSS.n5346 VSS.n5345 9.3005
R7112 VSS.n5347 VSS.n5323 9.3005
R7113 VSS.n5322 VSS.n178 9.3005
R7114 VSS.n5321 VSS.n5320 9.3005
R7115 VSS.n5319 VSS.n179 9.3005
R7116 VSS.n5317 VSS.n5316 9.3005
R7117 VSS.n5315 VSS.n180 9.3005
R7118 VSS.n5314 VSS.n5313 9.3005
R7119 VSS.n5312 VSS.n181 9.3005
R7120 VSS.n5310 VSS.n5309 9.3005
R7121 VSS.n5308 VSS.n182 9.3005
R7122 VSS.n5307 VSS.n5306 9.3005
R7123 VSS.n5305 VSS.n183 9.3005
R7124 VSS.n5304 VSS.n5303 9.3005
R7125 VSS.n5302 VSS.n185 9.3005
R7126 VSS.n5301 VSS.n5300 9.3005
R7127 VSS.n5299 VSS.n186 9.3005
R7128 VSS.n5298 VSS.n5297 9.3005
R7129 VSS.n5296 VSS.n187 9.3005
R7130 VSS.n5295 VSS.n5294 9.3005
R7131 VSS.n5292 VSS.n189 9.3005
R7132 VSS.n5289 VSS.n5288 9.3005
R7133 VSS.n5287 VSS.n190 9.3005
R7134 VSS.n5286 VSS.n5285 9.3005
R7135 VSS.n5284 VSS.n191 9.3005
R7136 VSS.n5282 VSS.n5281 9.3005
R7137 VSS.n5280 VSS.n192 9.3005
R7138 VSS.n5279 VSS.n5278 9.3005
R7139 VSS.n5275 VSS.n193 9.3005
R7140 VSS.n5274 VSS.n5273 9.3005
R7141 VSS.n5272 VSS.n195 9.3005
R7142 VSS.n5271 VSS.n5270 9.3005
R7143 VSS.n5269 VSS.n197 9.3005
R7144 VSS.n5268 VSS.n5267 9.3005
R7145 VSS.n5266 VSS.n198 9.3005
R7146 VSS.n5265 VSS.n5264 9.3005
R7147 VSS.n5263 VSS.n200 9.3005
R7148 VSS.n5262 VSS.n5261 9.3005
R7149 VSS.n5260 VSS.n201 9.3005
R7150 VSS.n5259 VSS.n5258 9.3005
R7151 VSS.n5257 VSS.n203 9.3005
R7152 VSS.n5254 VSS.n5253 9.3005
R7153 VSS.n5252 VSS.n204 9.3005
R7154 VSS.n5251 VSS.n5250 9.3005
R7155 VSS.n5249 VSS.n205 9.3005
R7156 VSS.n5248 VSS.n5247 9.3005
R7157 VSS.n5246 VSS.n206 9.3005
R7158 VSS.n5245 VSS.n5244 9.3005
R7159 VSS.n5243 VSS.n207 9.3005
R7160 VSS.n5242 VSS.n5241 9.3005
R7161 VSS.n5240 VSS.n5239 9.3005
R7162 VSS.n5238 VSS.n209 9.3005
R7163 VSS.n5235 VSS.n5234 9.3005
R7164 VSS.n5233 VSS.n210 9.3005
R7165 VSS.n5232 VSS.n5231 9.3005
R7166 VSS.n5229 VSS.n211 9.3005
R7167 VSS.n5228 VSS.n5227 9.3005
R7168 VSS.n5226 VSS.n212 9.3005
R7169 VSS.n5225 VSS.n5224 9.3005
R7170 VSS.n5222 VSS.n213 9.3005
R7171 VSS.n5221 VSS.n5220 9.3005
R7172 VSS.n5219 VSS.n5218 9.3005
R7173 VSS.n5217 VSS.n215 9.3005
R7174 VSS.n5216 VSS.n5215 9.3005
R7175 VSS.n5214 VSS.n218 9.3005
R7176 VSS.n5213 VSS.n5212 9.3005
R7177 VSS.n5211 VSS.n219 9.3005
R7178 VSS.n5210 VSS.n5209 9.3005
R7179 VSS.n5208 VSS.n220 9.3005
R7180 VSS.n5207 VSS.n5206 9.3005
R7181 VSS.n5204 VSS.n221 9.3005
R7182 VSS.n5203 VSS.n5202 9.3005
R7183 VSS.n5201 VSS.n5200 9.3005
R7184 VSS.n5199 VSS.n223 9.3005
R7185 VSS.n5198 VSS.n5197 9.3005
R7186 VSS.n5196 VSS.n225 9.3005
R7187 VSS.n5195 VSS.n5194 9.3005
R7188 VSS.n5193 VSS.n227 9.3005
R7189 VSS.n5191 VSS.n5190 9.3005
R7190 VSS.n5189 VSS.n228 9.3005
R7191 VSS.n5188 VSS.n5187 9.3005
R7192 VSS.n5186 VSS.n229 9.3005
R7193 VSS.n5185 VSS.n5184 9.3005
R7194 VSS.n5183 VSS.n232 9.3005
R7195 VSS.n5182 VSS.n5181 9.3005
R7196 VSS.n5180 VSS.n234 9.3005
R7197 VSS.n5139 VSS.n235 9.3005
R7198 VSS.n5141 VSS.n5140 9.3005
R7199 VSS.n5143 VSS.n5138 9.3005
R7200 VSS.n5147 VSS.n5146 9.3005
R7201 VSS.n5150 VSS.n5149 9.3005
R7202 VSS.n5151 VSS.n5136 9.3005
R7203 VSS.n5152 VSS.n5134 9.3005
R7204 VSS.n5154 VSS.n5153 9.3005
R7205 VSS.n5156 VSS.n5155 9.3005
R7206 VSS.n5157 VSS.n5131 9.3005
R7207 VSS.n5161 VSS.n5130 9.3005
R7208 VSS.n5163 VSS.n5162 9.3005
R7209 VSS.n5164 VSS.n5128 9.3005
R7210 VSS.n5166 VSS.n5165 9.3005
R7211 VSS.n5167 VSS.n5127 9.3005
R7212 VSS.n5169 VSS.n5168 9.3005
R7213 VSS.n5170 VSS.n5126 9.3005
R7214 VSS.n5171 VSS.n5125 9.3005
R7215 VSS.n5173 VSS.n5172 9.3005
R7216 VSS.n5174 VSS.n5124 9.3005
R7217 VSS.n5176 VSS.n5175 9.3005
R7218 VSS.n5177 VSS.n5122 9.3005
R7219 VSS.n5121 VSS.n236 9.3005
R7220 VSS.n5120 VSS.n5119 9.3005
R7221 VSS.n5117 VSS.n237 9.3005
R7222 VSS.n5116 VSS.n5115 9.3005
R7223 VSS.n5114 VSS.n5113 9.3005
R7224 VSS.n5112 VSS.n239 9.3005
R7225 VSS.n5111 VSS.n5110 9.3005
R7226 VSS.n5109 VSS.n241 9.3005
R7227 VSS.n5108 VSS.n5107 9.3005
R7228 VSS.n5106 VSS.n243 9.3005
R7229 VSS.n5105 VSS.n5104 9.3005
R7230 VSS.n5103 VSS.n244 9.3005
R7231 VSS.n5102 VSS.n5101 9.3005
R7232 VSS.n5100 VSS.n246 9.3005
R7233 VSS.n5099 VSS.n5098 9.3005
R7234 VSS.n5097 VSS.n247 9.3005
R7235 VSS.n5096 VSS.n5095 9.3005
R7236 VSS.n5094 VSS.n248 9.3005
R7237 VSS.n5093 VSS.n5092 9.3005
R7238 VSS.n5091 VSS.n250 9.3005
R7239 VSS.n5090 VSS.n5089 9.3005
R7240 VSS.n5088 VSS.n251 9.3005
R7241 VSS.n5087 VSS.n5086 9.3005
R7242 VSS.n5085 VSS.n252 9.3005
R7243 VSS.n5084 VSS.n5083 9.3005
R7244 VSS.n5082 VSS.n253 9.3005
R7245 VSS.n5081 VSS.n5080 9.3005
R7246 VSS.n5079 VSS.n254 9.3005
R7247 VSS.n5078 VSS.n5077 9.3005
R7248 VSS.n5076 VSS.n255 9.3005
R7249 VSS.n5075 VSS.n5074 9.3005
R7250 VSS.n5073 VSS.n256 9.3005
R7251 VSS.n5072 VSS.n5071 9.3005
R7252 VSS.n5070 VSS.n258 9.3005
R7253 VSS.n5068 VSS.n5067 9.3005
R7254 VSS.n5066 VSS.n259 9.3005
R7255 VSS.n5064 VSS.n5063 9.3005
R7256 VSS.n5062 VSS.n263 9.3005
R7257 VSS.n5060 VSS.n5059 9.3005
R7258 VSS.n5058 VSS.n264 9.3005
R7259 VSS.n5057 VSS.n5056 9.3005
R7260 VSS.n5055 VSS.n265 9.3005
R7261 VSS.n5051 VSS.n268 9.3005
R7262 VSS.n5050 VSS.n5049 9.3005
R7263 VSS.n5047 VSS.n269 9.3005
R7264 VSS.n5046 VSS.n5045 9.3005
R7265 VSS.n5044 VSS.n270 9.3005
R7266 VSS.n5043 VSS.n5042 9.3005
R7267 VSS.n5039 VSS.n271 9.3005
R7268 VSS.n5038 VSS.n5037 9.3005
R7269 VSS.n5036 VSS.n273 9.3005
R7270 VSS.n5035 VSS.n5034 9.3005
R7271 VSS.n5031 VSS.n275 9.3005
R7272 VSS.n5030 VSS.n5029 9.3005
R7273 VSS.n5028 VSS.n278 9.3005
R7274 VSS.n5027 VSS.n5026 9.3005
R7275 VSS.n5025 VSS.n279 9.3005
R7276 VSS.n5023 VSS.n5022 9.3005
R7277 VSS.n5021 VSS.n280 9.3005
R7278 VSS.n5019 VSS.n5018 9.3005
R7279 VSS.n5017 VSS.n284 9.3005
R7280 VSS.n5016 VSS.n5015 9.3005
R7281 VSS.n5014 VSS.n285 9.3005
R7282 VSS.n5013 VSS.n5012 9.3005
R7283 VSS.n5011 VSS.n287 9.3005
R7284 VSS.n5009 VSS.n5008 9.3005
R7285 VSS.n5007 VSS.n288 9.3005
R7286 VSS.n5005 VSS.n5004 9.3005
R7287 VSS.n5003 VSS.n292 9.3005
R7288 VSS.n5001 VSS.n5000 9.3005
R7289 VSS.n4999 VSS.n293 9.3005
R7290 VSS.n4998 VSS.n4997 9.3005
R7291 VSS.n295 VSS.n294 9.3005
R7292 VSS.n4898 VSS.n4897 9.3005
R7293 VSS.n4899 VSS.n4896 9.3005
R7294 VSS.n4901 VSS.n4900 9.3005
R7295 VSS.n4902 VSS.n4894 9.3005
R7296 VSS.n4903 VSS.n4892 9.3005
R7297 VSS.n4905 VSS.n4904 9.3005
R7298 VSS.n4906 VSS.n4891 9.3005
R7299 VSS.n4908 VSS.n4907 9.3005
R7300 VSS.n4909 VSS.n4890 9.3005
R7301 VSS.n4910 VSS.n4889 9.3005
R7302 VSS.n4912 VSS.n4911 9.3005
R7303 VSS.n4913 VSS.n4888 9.3005
R7304 VSS.n4915 VSS.n4914 9.3005
R7305 VSS.n4916 VSS.n4887 9.3005
R7306 VSS.n4917 VSS.n4886 9.3005
R7307 VSS.n4919 VSS.n4918 9.3005
R7308 VSS.n4920 VSS.n4885 9.3005
R7309 VSS.n4922 VSS.n4921 9.3005
R7310 VSS.n4923 VSS.n4883 9.3005
R7311 VSS.n4925 VSS.n4924 9.3005
R7312 VSS.n4926 VSS.n4882 9.3005
R7313 VSS.n4928 VSS.n4927 9.3005
R7314 VSS.n4929 VSS.n4881 9.3005
R7315 VSS.n4931 VSS.n4930 9.3005
R7316 VSS.n4932 VSS.n4880 9.3005
R7317 VSS.n4934 VSS.n4933 9.3005
R7318 VSS.n4935 VSS.n4878 9.3005
R7319 VSS.n4877 VSS.n370 9.3005
R7320 VSS.n4876 VSS.n4875 9.3005
R7321 VSS.n4874 VSS.n371 9.3005
R7322 VSS.n4871 VSS.n4870 9.3005
R7323 VSS.n4869 VSS.n373 9.3005
R7324 VSS.n4868 VSS.n4867 9.3005
R7325 VSS.n4865 VSS.n374 9.3005
R7326 VSS.n4864 VSS.n4863 9.3005
R7327 VSS.n4862 VSS.n375 9.3005
R7328 VSS.n4861 VSS.n4860 9.3005
R7329 VSS.n4859 VSS.n376 9.3005
R7330 VSS.n4857 VSS.n4856 9.3005
R7331 VSS.n379 VSS.n378 9.3005
R7332 VSS.n4845 VSS.n4844 9.3005
R7333 VSS.n4846 VSS.n385 9.3005
R7334 VSS.n4848 VSS.n4847 9.3005
R7335 VSS.n4834 VSS.n386 9.3005
R7336 VSS.n4833 VSS.n4832 9.3005
R7337 VSS.n4831 VSS.n388 9.3005
R7338 VSS.n4830 VSS.n4829 9.3005
R7339 VSS.n4828 VSS.n389 9.3005
R7340 VSS.n4827 VSS.n4826 9.3005
R7341 VSS.n4825 VSS.n4824 9.3005
R7342 VSS.n4821 VSS.n391 9.3005
R7343 VSS.n4820 VSS.n4819 9.3005
R7344 VSS.n4818 VSS.n393 9.3005
R7345 VSS.n4817 VSS.n4816 9.3005
R7346 VSS.n460 VSS.n459 9.3005
R7347 VSS.n458 VSS.n457 9.3005
R7348 VSS.n456 VSS.n396 9.3005
R7349 VSS.n453 VSS.n452 9.3005
R7350 VSS.n451 VSS.n397 9.3005
R7351 VSS.n450 VSS.n449 9.3005
R7352 VSS.n448 VSS.n398 9.3005
R7353 VSS.n447 VSS.n446 9.3005
R7354 VSS.n445 VSS.n401 9.3005
R7355 VSS.n444 VSS.n443 9.3005
R7356 VSS.n442 VSS.n402 9.3005
R7357 VSS.n441 VSS.n440 9.3005
R7358 VSS.n439 VSS.n404 9.3005
R7359 VSS.n438 VSS.n437 9.3005
R7360 VSS.n436 VSS.n405 9.3005
R7361 VSS.n435 VSS.n434 9.3005
R7362 VSS.n433 VSS.n407 9.3005
R7363 VSS.n432 VSS.n431 9.3005
R7364 VSS.n430 VSS.n408 9.3005
R7365 VSS.n429 VSS.n428 9.3005
R7366 VSS.n427 VSS.n410 9.3005
R7367 VSS.n426 VSS.n425 9.3005
R7368 VSS.n424 VSS.n411 9.3005
R7369 VSS.n423 VSS.n422 9.3005
R7370 VSS.n421 VSS.n413 9.3005
R7371 VSS.n4815 VSS.n394 9.3005
R7372 VSS.n4596 VSS.n469 9.3005
R7373 VSS.n4600 VSS.n4599 9.3005
R7374 VSS.n4601 VSS.n4592 9.3005
R7375 VSS.n4610 VSS.n4602 9.3005
R7376 VSS.n4608 VSS.n4607 9.3005
R7377 VSS.n4802 VSS.n471 9.3005
R7378 VSS.n984 VSS.n983 9.3005
R7379 VSS.n1220 VSS.n1219 9.3005
R7380 VSS.n1218 VSS.n979 9.3005
R7381 VSS.n1217 VSS.n1216 9.3005
R7382 VSS.n1214 VSS.n986 9.3005
R7383 VSS.n1616 VSS.n1615 9.29365
R7384 VSS.n4745 VSS.n545 9.25132
R7385 VSS.n545 VSS.n544 9.25132
R7386 VSS.n2229 VSS.n2228 8.90485
R7387 VSS.n1145 VSS.n1139 8.88145
R7388 VSS.n945 VSS.n939 8.88145
R7389 VSS.n1070 VSS.n307 8.86414
R7390 VSS.t693 VSS.n307 8.86414
R7391 VSS.n1069 VSS.n306 8.86414
R7392 VSS.t693 VSS.n306 8.86414
R7393 VSS.n1154 VSS.n1139 8.8249
R7394 VSS.n945 VSS.n938 8.8249
R7395 VSS.n3595 VSS.n3594 8.8005
R7396 VSS.n3401 VSS.n3057 8.79436
R7397 VSS.n2636 VSS.n2198 8.67847
R7398 VSS.n4283 VSS.n3743 8.65932
R7399 VSS.n4944 VSS.n4943 8.64324
R7400 VSS.n4943 VSS.n362 8.64324
R7401 VSS.n4961 VSS.n4960 8.64324
R7402 VSS.n332 VSS.n331 8.58762
R7403 VSS.n1145 VSS.n1138 8.54514
R7404 VSS.n4664 VSS.n939 8.54514
R7405 VSS.n3329 VSS.n3326 8.53383
R7406 VSS.t462 VSS.t1083 8.42962
R7407 VSS.t464 VSS.t1085 8.42962
R7408 VSS.t1262 VSS.t607 8.42962
R7409 VSS.t2973 VSS.t2185 8.42962
R7410 VSS.t2975 VSS.t2183 8.42962
R7411 VSS.t1520 VSS.t322 8.42962
R7412 VSS.t1522 VSS.t318 8.42962
R7413 VSS.t719 VSS.t3018 8.42962
R7414 VSS.t2782 VSS.t1993 8.42962
R7415 VSS.t2786 VSS.t1991 8.42962
R7416 VSS.t735 VSS.t434 8.42962
R7417 VSS.t737 VSS.t432 8.42962
R7418 VSS.t832 VSS.t2925 8.42962
R7419 VSS.t830 VSS.t2927 8.42962
R7420 VSS.n967 VSS.n965 8.32651
R7421 VSS.n4030 VSS.n4027 8.2968
R7422 VSS.n1642 VSS.n1639 8.2968
R7423 VSS.n4163 VSS.n4161 8.28285
R7424 VSS.n1705 VSS.n1704 8.28285
R7425 VSS.n4665 VSS.n938 8.2471
R7426 VSS.n1155 VSS.n1154 8.24672
R7427 VSS.n4568 VSS.n4567 8.23546
R7428 VSS.n4569 VSS.n4568 8.23546
R7429 VSS.n4569 VSS.n4562 8.23546
R7430 VSS.n4573 VSS.n4562 8.23546
R7431 VSS.n4574 VSS.n4573 8.23546
R7432 VSS.n4575 VSS.n4574 8.23546
R7433 VSS.n4579 VSS.n4578 8.23546
R7434 VSS.n4580 VSS.n4579 8.23546
R7435 VSS.n5712 VSS.n5711 8.23546
R7436 VSS.n5713 VSS.n5712 8.23546
R7437 VSS.n5713 VSS.n30 8.23546
R7438 VSS.n5717 VSS.n30 8.23546
R7439 VSS.n5718 VSS.n5717 8.23546
R7440 VSS.n5720 VSS.n5718 8.23546
R7441 VSS.n5724 VSS.n28 8.23546
R7442 VSS.n5725 VSS.n5724 8.23546
R7443 VSS.n5624 VSS.n5623 8.23546
R7444 VSS.n5625 VSS.n5624 8.23546
R7445 VSS.n5625 VSS.n72 8.23546
R7446 VSS.n5629 VSS.n72 8.23546
R7447 VSS.n5630 VSS.n5629 8.23546
R7448 VSS.n5631 VSS.n5630 8.23546
R7449 VSS.n5635 VSS.n5634 8.23546
R7450 VSS.n5636 VSS.n5635 8.23546
R7451 VSS.n5534 VSS.n110 8.23546
R7452 VSS.n5535 VSS.n5534 8.23546
R7453 VSS.n5536 VSS.n5535 8.23546
R7454 VSS.n5536 VSS.n108 8.23546
R7455 VSS.n5540 VSS.n108 8.23546
R7456 VSS.n5541 VSS.n5540 8.23546
R7457 VSS.n5543 VSS.n106 8.23546
R7458 VSS.n5547 VSS.n106 8.23546
R7459 VSS.n5439 VSS.n5438 8.23546
R7460 VSS.n5440 VSS.n5439 8.23546
R7461 VSS.n5440 VSS.n151 8.23546
R7462 VSS.n5444 VSS.n151 8.23546
R7463 VSS.n5445 VSS.n5444 8.23546
R7464 VSS.n5446 VSS.n5445 8.23546
R7465 VSS.n5450 VSS.n5449 8.23546
R7466 VSS.n5452 VSS.n5450 8.23546
R7467 VSS.n5402 VSS.n167 8.23546
R7468 VSS.n5403 VSS.n5402 8.23546
R7469 VSS.n5404 VSS.n5403 8.23546
R7470 VSS.n5404 VSS.n165 8.23546
R7471 VSS.n5408 VSS.n165 8.23546
R7472 VSS.n5409 VSS.n5408 8.23546
R7473 VSS.n5411 VSS.n163 8.23546
R7474 VSS.n5415 VSS.n163 8.23546
R7475 VSS.n4322 VSS.n4321 8.23546
R7476 VSS.n4339 VSS.n4338 8.23546
R7477 VSS.n4466 VSS.n4465 8.23546
R7478 VSS.n2115 VSS.n2114 8.23546
R7479 VSS.n2109 VSS.n2108 8.23546
R7480 VSS.n2565 VSS.n2564 8.23546
R7481 VSS.n2567 VSS.n2565 8.23546
R7482 VSS.n2571 VSS.n2224 8.23546
R7483 VSS.n2572 VSS.n2571 8.23546
R7484 VSS.n2576 VSS.n2572 8.23546
R7485 VSS.n2580 VSS.n2222 8.23546
R7486 VSS.n2512 VSS.n2251 8.23546
R7487 VSS.n2516 VSS.n2251 8.23546
R7488 VSS.n2517 VSS.n2516 8.23546
R7489 VSS.n2520 VSS.n2517 8.23546
R7490 VSS.n2524 VSS.n2249 8.23546
R7491 VSS.n2527 VSS.n2526 8.23546
R7492 VSS.n2417 VSS.n2414 8.23546
R7493 VSS.n2421 VSS.n2308 8.23546
R7494 VSS.n2424 VSS.n2423 8.23546
R7495 VSS.n2430 VSS.n2429 8.23546
R7496 VSS.n2407 VSS.n2406 8.23546
R7497 VSS.n2755 VSS.n2754 8.23546
R7498 VSS.n2756 VSS.n2755 8.23546
R7499 VSS.n2756 VSS.n2178 8.23546
R7500 VSS.n2760 VSS.n2178 8.23546
R7501 VSS.n2765 VSS.n2762 8.23546
R7502 VSS.n2769 VSS.n2768 8.23546
R7503 VSS.n2923 VSS.n2922 8.23546
R7504 VSS.n2920 VSS.n2158 8.23546
R7505 VSS.n2916 VSS.n2158 8.23546
R7506 VSS.n2916 VSS.n2915 8.23546
R7507 VSS.n2915 VSS.n2914 8.23546
R7508 VSS.n1598 VSS.n1543 8.23546
R7509 VSS.n4961 VSS.n4959 8.20563
R7510 VSS.n2582 VSS.n2581 8.14595
R7511 VSS.n2714 VSS.n2713 8.10717
R7512 VSS.n4611 VSS.t2638 8.10019
R7513 VSS.n3954 VSS.n3951 8.05976
R7514 VSS.n3573 VSS.n2977 8.05976
R7515 VSS.n4325 VSS.n3726 8.05644
R7516 VSS.n3214 VSS.n3213 8.05644
R7517 VSS.n2119 VSS.n2118 8.05644
R7518 VSS.n2113 VSS.n2112 8.05644
R7519 VSS.n2107 VSS.n2106 8.05644
R7520 VSS.n2771 VSS.n2770 8.05644
R7521 VSS.n2910 VSS.n2909 8.05644
R7522 VSS.n1600 VSS.n1599 8.05644
R7523 VSS.n1602 VSS.n1541 8.05644
R7524 VSS.n1313 VSS.n1265 8.05644
R7525 VSS.n1306 VSS.n1267 8.05644
R7526 VSS.t64 VSS.n4948 8.04732
R7527 VSS.n2510 VSS.n2509 7.97427
R7528 VSS.n4139 VSS.n3769 7.90638
R7529 VSS.n4146 VSS.n4144 7.90638
R7530 VSS.n4204 VSS.n4182 7.90638
R7531 VSS.n4359 VSS.n4358 7.90638
R7532 VSS.n4408 VSS.n3696 7.90638
R7533 VSS.n3668 VSS.n2138 7.90638
R7534 VSS.n3623 VSS.n3622 7.90638
R7535 VSS.n3524 VSS.n3523 7.90638
R7536 VSS.n2438 VSS.n2301 7.90638
R7537 VSS.n2729 VSS.n2728 7.90638
R7538 VSS.n2034 VSS.n2030 7.90638
R7539 VSS.n1955 VSS.n1954 7.90638
R7540 VSS.n1934 VSS.n1391 7.90638
R7541 VSS.n1777 VSS.n1472 7.90638
R7542 VSS.n1722 VSS.n1495 7.90638
R7543 VSS.n1714 VSS.n1497 7.90638
R7544 VSS.n3215 VSS.n3214 7.87742
R7545 VSS.n2118 VSS.n2073 7.87742
R7546 VSS.n1602 VSS.n1601 7.87742
R7547 VSS.n1313 VSS.n1312 7.87742
R7548 VSS.n1306 VSS.n1305 7.87742
R7549 VSS.n3621 VSS.n3620 7.76768
R7550 VSS.n3313 VSS.n3311 7.76768
R7551 VSS.n4567 VSS.n4564 7.6984
R7552 VSS.n4580 VSS.n4558 7.6984
R7553 VSS.n5711 VSS.n32 7.6984
R7554 VSS.n5726 VSS.n5725 7.6984
R7555 VSS.n5623 VSS.n74 7.6984
R7556 VSS.n5636 VSS.n68 7.6984
R7557 VSS.n5529 VSS.n110 7.6984
R7558 VSS.n5548 VSS.n5547 7.6984
R7559 VSS.n5438 VSS.n153 7.6984
R7560 VSS.n5452 VSS.n5451 7.6984
R7561 VSS.n5397 VSS.n167 7.6984
R7562 VSS.n5416 VSS.n5415 7.6984
R7563 VSS.n4321 VSS.n4320 7.6984
R7564 VSS.n4340 VSS.n4339 7.6984
R7565 VSS.n4462 VSS.n4461 7.6984
R7566 VSS.n3216 VSS.n3161 7.6984
R7567 VSS.n2106 VSS.n2078 7.6984
R7568 VSS.n2564 VSS.n2226 7.6984
R7569 VSS.n2583 VSS.n2582 7.6984
R7570 VSS.n2512 VSS.n2511 7.6984
R7571 VSS.n2531 VSS.n2530 7.6984
R7572 VSS.n2430 VSS.n2303 7.6984
R7573 VSS.n2754 VSS.n2180 7.6984
R7574 VSS.n2923 VSS.n2155 7.6984
R7575 VSS.n1304 VSS.n1303 7.6984
R7576 VSS.n3918 VSS.n3917 7.65267
R7577 VSS.n4462 VSS.n4434 7.60889
R7578 VSS.n2762 VSS.n2761 7.60889
R7579 VSS.n1592 VSS.n1543 7.60889
R7580 VSS.n3943 VSS.n3941 7.6005
R7581 VSS.n3448 VSS.n3447 7.6005
R7582 VSS.n1988 VSS.n1987 7.6005
R7583 VSS.n4132 VSS.n4131 7.52991
R7584 VSS.n4154 VSS.n4153 7.52991
R7585 VSS.n4354 VSS.n4353 7.52991
R7586 VSS.n3512 VSS.n3511 7.52991
R7587 VSS.n3270 VSS.n3269 7.52991
R7588 VSS.n2594 VSS.n2593 7.52991
R7589 VSS.n2052 VSS.n1337 7.52991
R7590 VSS.n1083 VSS.n1033 7.26779
R7591 VSS.n3285 VSS.n3106 7.23528
R7592 VSS.n3278 VSS.n3111 7.23528
R7593 VSS.n346 VSS.n345 7.16275
R7594 VSS.n1735 VSS.n1734 7.15344
R7595 VSS.n3212 VSS.n3162 7.15139
R7596 VSS.n332 VSS.n330 7.15034
R7597 VSS.n2406 VSS.n2314 7.11268
R7598 VSS.n967 VSS.n966 7.02466
R7599 VSS.n4316 VSS.n3728 7.00731
R7600 VSS.n4335 VSS.n3721 6.98232
R7601 VSS.n2519 VSS.n2249 6.98232
R7602 VSS.n2922 VSS.n2921 6.98232
R7603 VSS.n4326 VSS.n4325 6.90655
R7604 VSS.n4333 VSS.n4332 6.90655
R7605 VSS.n1606 VSS.n1605 6.88949
R7606 VSS.n1317 VSS.n1316 6.88949
R7607 VSS.n4288 VSS.n4287 6.77697
R7608 VSS.n2010 VSS.n1353 6.77697
R7609 VSS.n1955 VSS.n1379 6.77697
R7610 VSS.n1904 VSS.n1903 6.77697
R7611 VSS.n1859 VSS.n1427 6.77697
R7612 VSS.n1803 VSS.n1802 6.77697
R7613 VSS.n1780 VSS.n1468 6.77697
R7614 VSS.n1760 VSS.n1759 6.77697
R7615 VSS.n1650 VSS.n1649 6.77697
R7616 VSS.n1628 VSS.n1627 6.75062
R7617 VSS.n2972 VSS.n2968 6.7205
R7618 VSS.n2567 VSS.n2566 6.71379
R7619 VSS.n342 VSS.n340 6.67472
R7620 VSS.n2423 VSS.n2422 6.62428
R7621 VSS.n1618 VSS.n1617 6.6092
R7622 VSS.n4796 VSS.n4795 6.57154
R7623 VSS.n3591 VSS.n3590 6.53554
R7624 VSS.t2838 VSS.t1697 6.52095
R7625 VSS.n5596 VSS.n5595 6.4005
R7626 VSS.n4203 VSS.n4202 6.4005
R7627 VSS.n4412 VSS.n4411 6.4005
R7628 VSS.n3683 VSS.n3682 6.4005
R7629 VSS.n3675 VSS.n3674 6.4005
R7630 VSS.n3518 VSS.n3517 6.4005
R7631 VSS.n3437 VSS.n3037 6.4005
R7632 VSS.n3244 VSS.n3243 6.4005
R7633 VSS.n2494 VSS.n2493 6.4005
R7634 VSS.n2478 VSS.n2477 6.4005
R7635 VSS.n2907 VSS.n2906 6.4005
R7636 VSS.n1998 VSS.n1997 6.4005
R7637 VSS.n1838 VSS.n1837 6.4005
R7638 VSS.n5256 VSS.n5254 6.4005
R7639 VSS.n2530 VSS.n2247 6.26623
R7640 VSS.n5750 VSS.n5749 6.26433
R7641 VSS.n5705 VSS.n35 6.26433
R7642 VSS.n5686 VSS.n5685 6.26433
R7643 VSS.n5660 VSS.n57 6.26433
R7644 VSS.n5661 VSS.n5660 6.26433
R7645 VSS.n5616 VSS.n76 6.26433
R7646 VSS.n5570 VSS.n5569 6.26433
R7647 VSS.n5560 VSS.n5559 6.26433
R7648 VSS.n5525 VSS.n112 6.26433
R7649 VSS.n5476 VSS.n135 6.26433
R7650 VSS.n5477 VSS.n5476 6.26433
R7651 VSS.n5465 VSS.n5464 6.26433
R7652 VSS.n5431 VSS.n155 6.26433
R7653 VSS.n3927 VSS.n3826 6.26433
R7654 VSS.n4054 VSS.n3807 6.26433
R7655 VSS.n4054 VSS.n3808 6.26433
R7656 VSS.n4050 VSS.n3808 6.26433
R7657 VSS.n4077 VSS.n3799 6.26433
R7658 VSS.n4078 VSS.n4077 6.26433
R7659 VSS.n4109 VSS.n4107 6.26433
R7660 VSS.n4226 VSS.n4225 6.26433
R7661 VSS.n4263 VSS.n4262 6.26433
R7662 VSS.n4313 VSS.n4312 6.26433
R7663 VSS.n3600 VSS.n2966 6.26433
R7664 VSS.n3470 VSS.n3027 6.26433
R7665 VSS.n3453 VSS.n3452 6.26433
R7666 VSS.n3393 VSS.n3392 6.26433
R7667 VSS.n3352 VSS.n3351 6.26433
R7668 VSS.n3352 VSS.n3077 6.26433
R7669 VSS.n3293 VSS.n3292 6.26433
R7670 VSS.n3284 VSS.n3107 6.26433
R7671 VSS.n2718 VSS.n2717 6.26433
R7672 VSS.n2746 VSS.n2182 6.26433
R7673 VSS.n1912 VSS.n1400 6.26433
R7674 VSS.n1678 VSS.n1514 6.26433
R7675 VSS.n1679 VSS.n1678 6.26433
R7676 VSS.n4875 VSS.n4874 6.26433
R7677 VSS.n5009 VSS.n288 6.26433
R7678 VSS.n5023 VSS.n280 6.26433
R7679 VSS.n5056 VSS.n5055 6.26433
R7680 VSS.n5068 VSS.n259 6.26433
R7681 VSS.n5117 VSS.n5116 6.26433
R7682 VSS.n5157 VSS.n5156 6.26433
R7683 VSS.n5146 VSS.n5143 6.26433
R7684 VSS.n5191 VSS.n228 6.26433
R7685 VSS.n5204 VSS.n5203 6.26433
R7686 VSS.n5222 VSS.n5221 6.26433
R7687 VSS.n5239 VSS.n5238 6.26433
R7688 VSS.n457 VSS.n456 6.26433
R7689 VSS.n474 VSS.n473 6.21883
R7690 VSS.n4606 VSS.n4604 6.21725
R7691 VSS.n982 VSS.n980 6.21725
R7692 VSS.n1169 VSS.n1168 6.20545
R7693 VSS.n3929 VSS.n3928 6.19624
R7694 VSS.n4261 VSS.n4260 6.19624
R7695 VSS.n2704 VSS.n2703 6.19624
R7696 VSS.n4049 VSS.n4048 6.12816
R7697 VSS.n3277 VSS.n3276 6.12816
R7698 VSS.n2372 VSS.n2371 6.12816
R7699 VSS.n1681 VSS.n1680 6.12816
R7700 VSS.n3190 VSS.n3189 6.0286
R7701 VSS.n3949 VSS.n3818 6.02403
R7702 VSS.n1985 VSS.n1984 6.02403
R7703 VSS.n4676 VSS.n478 6.0005
R7704 VSS.n909 VSS.n478 6.0005
R7705 VSS.n3601 VSS.n3600 5.99199
R7706 VSS.n4513 VSS.n4512 5.98311
R7707 VSS.n5741 VSS.n5739 5.98311
R7708 VSS.n5587 VSS.n5586 5.98311
R7709 VSS.n5366 VSS.n5363 5.98311
R7710 VSS.n3864 VSS.n3846 5.98311
R7711 VSS.n4299 VSS.n3735 5.98311
R7712 VSS.n3406 VSS.n3404 5.98311
R7713 VSS.n3224 VSS.n3157 5.98311
R7714 VSS.n2488 VSS.n2486 5.98311
R7715 VSS.n1990 VSS.n1989 5.98311
R7716 VSS.n1890 VSS.n1409 5.98311
R7717 VSS.n1632 VSS.n1629 5.98311
R7718 VSS.n4824 VSS.n390 5.98311
R7719 VSS.n5034 VSS.n276 5.98311
R7720 VSS.n5042 VSS.n272 5.98311
R7721 VSS.n5278 VSS.n194 5.98311
R7722 VSS.n5293 VSS.n5292 5.98311
R7723 VSS.n5334 VSS.n5333 5.98311
R7724 VSS.n418 VSS.n417 5.98311
R7725 VSS.n2428 VSS.n2427 5.90819
R7726 VSS.t2041 VSS.t2842 5.86891
R7727 VSS.n5749 VSS.n17 5.85582
R7728 VSS.n5700 VSS.n35 5.85582
R7729 VSS.n5685 VSS.n45 5.85582
R7730 VSS.n5655 VSS.n57 5.85582
R7731 VSS.n5611 VSS.n76 5.85582
R7732 VSS.n5569 VSS.n5568 5.85582
R7733 VSS.n5559 VSS.n101 5.85582
R7734 VSS.n5520 VSS.n112 5.85582
R7735 VSS.n5471 VSS.n135 5.85582
R7736 VSS.n5464 VSS.n5463 5.85582
R7737 VSS.n5426 VSS.n155 5.85582
R7738 VSS.n3977 VSS.n3807 5.85582
R7739 VSS.n4046 VSS.n3983 5.85582
R7740 VSS.n4072 VSS.n3799 5.85582
R7741 VSS.n4226 VSS.n4173 5.85582
R7742 VSS.n4257 VSS.n4256 5.85582
R7743 VSS.n4263 VSS.n3750 5.85582
R7744 VSS.n4312 VSS.n3730 5.85582
R7745 VSS.n3592 VSS.n2966 5.85582
R7746 VSS.n3452 VSS.n3034 5.85582
R7747 VSS.n3392 VSS.n3062 5.85582
R7748 VSS.n3351 VSS.n3350 5.85582
R7749 VSS.n3292 VSS.n3103 5.85582
R7750 VSS.n3275 VSS.n3113 5.85582
R7751 VSS.n2605 VSS.n2604 5.85582
R7752 VSS.n2457 VSS.n2456 5.85582
R7753 VSS.n2371 VSS.n2324 5.85582
R7754 VSS.n2706 VSS.n2705 5.85582
R7755 VSS.n2060 VSS.n2059 5.85582
R7756 VSS.n1910 VSS.n1909 5.85582
R7757 VSS.n1865 VSS.n1864 5.85582
R7758 VSS.n1681 VSS.n1511 5.85582
R7759 VSS.n4875 VSS.n372 5.85582
R7760 VSS.n5010 VSS.n5009 5.85582
R7761 VSS.n5024 VSS.n5023 5.85582
R7762 VSS.n5056 VSS.n266 5.85582
R7763 VSS.n5069 VSS.n5068 5.85582
R7764 VSS.n5118 VSS.n5117 5.85582
R7765 VSS.n5156 VSS.n5133 5.85582
R7766 VSS.n5143 VSS.n5142 5.85582
R7767 VSS.n5192 VSS.n5191 5.85582
R7768 VSS.n5205 VSS.n5204 5.85582
R7769 VSS.n5223 VSS.n5222 5.85582
R7770 VSS.n5239 VSS.n208 5.85582
R7771 VSS.n457 VSS.n395 5.85582
R7772 VSS.n4482 VSS.n4426 5.80542
R7773 VSS.n3921 VSS.n3826 5.78773
R7774 VSS.n2408 VSS.n2407 5.72917
R7775 VSS.n5662 VSS.n5661 5.65809
R7776 VSS.n5478 VSS.n5477 5.65809
R7777 VSS.n3932 VSS.n3929 5.65809
R7778 VSS.n3603 VSS.n3602 5.65809
R7779 VSS.n3356 VSS.n3077 5.65809
R7780 VSS.n1916 VSS.n1400 5.65809
R7781 VSS.n2460 VSS.n2458 5.65156
R7782 VSS.n2740 VSS.n2182 5.65156
R7783 VSS.n2121 VSS.n2120 5.63966
R7784 VSS.n2412 VSS.n2310 5.63966
R7785 VSS.n2771 VSS.n2172 5.63966
R7786 VSS.n2909 VSS.n2908 5.63966
R7787 VSS.n3232 VSS.n3131 5.5878
R7788 VSS.n4260 VSS.n3754 5.58348
R7789 VSS.n3296 VSS.n3294 5.52192
R7790 VSS.n3286 VSS.n3105 5.51774
R7791 VSS.n3279 VSS.n3110 5.51774
R7792 VSS.n1148 VSS.n1146 5.48621
R7793 VSS.n944 VSS.n940 5.48621
R7794 VSS.n973 VSS.n972 5.438
R7795 VSS.n1645 VSS.n1644 5.37692
R7796 VSS.n2374 VSS.n2373 5.37524
R7797 VSS.n2560 VSS.n2558 5.35702
R7798 VSS.n4010 VSS.n4002 5.27109
R7799 VSS.n4234 VSS.n4233 5.27109
R7800 VSS.n4358 VSS.n3712 5.27109
R7801 VSS.n4418 VSS.n4417 5.27109
R7802 VSS.n4106 VSS.n4105 5.24305
R7803 VSS.n3464 VSS.n3027 5.24305
R7804 VSS.n322 VSS.n321 5.22706
R7805 VSS.n1152 VSS.n1151 5.22371
R7806 VSS.n1151 VSS.n1150 5.22371
R7807 VSS.n1149 VSS.n1148 5.22371
R7808 VSS.n1150 VSS.n1149 5.22371
R7809 VSS.n4660 VSS.n948 5.22371
R7810 VSS.n4660 VSS.n4659 5.22371
R7811 VSS.n944 VSS.n942 5.22371
R7812 VSS.n4659 VSS.n942 5.22371
R7813 VSS.n2416 VSS.n2308 5.19211
R7814 VSS.n1699 VSS.n1697 5.14833
R7815 VSS.n3854 VSS.n3852 5.13108
R7816 VSS.n3854 VSS.n3853 5.13108
R7817 VSS.n4445 VSS.n4443 5.13108
R7818 VSS.n4445 VSS.n4444 5.13108
R7819 VSS.n3142 VSS.n3140 5.13108
R7820 VSS.n3142 VSS.n3141 5.13108
R7821 VSS.n2090 VSS.n2088 5.13108
R7822 VSS.n2090 VSS.n2089 5.13108
R7823 VSS.n2343 VSS.n2341 5.13108
R7824 VSS.n2343 VSS.n2342 5.13108
R7825 VSS.n2856 VSS.n2854 5.13108
R7826 VSS.n2856 VSS.n2855 5.13108
R7827 VSS.n2165 VSS.n2164 5.13108
R7828 VSS.n1563 VSS.n1561 5.13108
R7829 VSS.n1563 VSS.n1562 5.13108
R7830 VSS.n1281 VSS.n1279 5.13108
R7831 VSS.n1281 VSS.n1280 5.13108
R7832 VSS.n1028 VSS.n1027 5.11682
R7833 VSS.n1031 VSS.n1030 5.063
R7834 VSS.n2125 VSS.n2124 5.04614
R7835 VSS.n2386 VSS.n2385 5.04614
R7836 VSS.n4080 VSS.n4079 5.04533
R7837 VSS.n2385 VSS.n2384 5.03813
R7838 VSS.n1260 VSS.t2646 4.98492
R7839 VSS.n3620 VSS.n3618 4.94085
R7840 VSS.n3314 VSS.n3313 4.94085
R7841 VSS.n2061 VSS.n2060 4.90263
R7842 VSS.n2789 VSS.n2788 4.89462
R7843 VSS.n5667 VSS.n54 4.85762
R7844 VSS.n5484 VSS.n132 4.85762
R7845 VSS.n4085 VSS.n3796 4.85762
R7846 VSS.n3938 VSS.n3822 4.85762
R7847 VSS.n3302 VSS.n3098 4.85762
R7848 VSS.n3360 VSS.n3359 4.85762
R7849 VSS.n3609 VSS.n2963 4.85762
R7850 VSS.n2888 VSS.n2887 4.85762
R7851 VSS.n2640 VSS.n2196 4.85762
R7852 VSS.n1920 VSS.n1919 4.85762
R7853 VSS.n4729 VSS.t2431 4.80635
R7854 VSS.n479 VSS.t2378 4.80635
R7855 VSS.n4512 VSS.n4511 4.8005
R7856 VSS.n5741 VSS.n5740 4.8005
R7857 VSS.n5588 VSS.n5587 4.8005
R7858 VSS.n5366 VSS.n5365 4.8005
R7859 VSS.n3865 VSS.n3864 4.8005
R7860 VSS.n4300 VSS.n4299 4.8005
R7861 VSS.n3588 VSS.n3587 4.8005
R7862 VSS.n3406 VSS.n3405 4.8005
R7863 VSS.n2488 VSS.n2487 4.8005
R7864 VSS.n1991 VSS.n1990 4.8005
R7865 VSS.n1699 VSS.n1698 4.8005
R7866 VSS.n1632 VSS.n1631 4.8005
R7867 VSS.n4824 VSS.n4823 4.8005
R7868 VSS.n5034 VSS.n5033 4.8005
R7869 VSS.n5042 VSS.n5041 4.8005
R7870 VSS.n5278 VSS.n5277 4.8005
R7871 VSS.n5292 VSS.n5291 4.8005
R7872 VSS.n5333 VSS.n5332 4.8005
R7873 VSS.n417 VSS.n416 4.8005
R7874 VSS.n320 VSS.n318 4.79738
R7875 VSS.n3855 VSS.n3851 4.75748
R7876 VSS.n3144 VSS.n3143 4.75748
R7877 VSS.n2344 VSS.n2340 4.75748
R7878 VSS.n1564 VSS.n1560 4.75748
R7879 VSS.n4447 VSS.n4446 4.75739
R7880 VSS.n2091 VSS.n2087 4.75739
R7881 VSS.n2858 VSS.n2857 4.75739
R7882 VSS.n1283 VSS.n1282 4.75739
R7883 VSS.n2124 VSS.n2123 4.75419
R7884 VSS.n3901 VSS.n3900 4.67352
R7885 VSS.n3901 VSS.n3834 4.67352
R7886 VSS.n3905 VSS.n3834 4.67352
R7887 VSS.n3906 VSS.n3905 4.67352
R7888 VSS.n3907 VSS.n3906 4.67352
R7889 VSS.n3913 VSS.n3912 4.67352
R7890 VSS.n4478 VSS.n4477 4.67352
R7891 VSS.n4477 VSS.n4476 4.67352
R7892 VSS.n4473 VSS.n4472 4.67352
R7893 VSS.n4472 VSS.n4471 4.67352
R7894 VSS.n3187 VSS.n3172 4.67352
R7895 VSS.n3183 VSS.n3172 4.67352
R7896 VSS.n3181 VSS.n3180 4.67352
R7897 VSS.n3180 VSS.n3177 4.67352
R7898 VSS.n3194 VSS.n3169 4.67352
R7899 VSS.n3208 VSS.n3207 4.67352
R7900 VSS.n3207 VSS.n3206 4.67352
R7901 VSS.n3203 VSS.n3202 4.67352
R7902 VSS.n3202 VSS.n3201 4.67352
R7903 VSS.n2393 VSS.n2318 4.67352
R7904 VSS.n2394 VSS.n2393 4.67352
R7905 VSS.n2395 VSS.n2394 4.67352
R7906 VSS.n2399 VSS.n2398 4.67352
R7907 VSS.n2402 VSS.n2399 4.67352
R7908 VSS.n2907 VSS.n2163 4.62124
R7909 VSS.n2560 VSS.n2227 4.62124
R7910 VSS.n1612 VSS.n1538 4.62124
R7911 VSS.n1618 VSS.n1537 4.62124
R7912 VSS.n2908 VSS.n2907 4.6085
R7913 VSS.n615 VSS.n614 4.57739
R7914 VSS.n614 VSS.n548 4.57739
R7915 VSS.n855 VSS.n854 4.57739
R7916 VSS.n854 VSS.n788 4.57739
R7917 VSS.n3898 VSS.n3836 4.55559
R7918 VSS.n2389 VSS.n2387 4.55559
R7919 VSS.n3682 VSS.n3681 4.51815
R7920 VSS.n5775 VSS.n3 4.51401
R7921 VSS.n8 VSS.n7 4.51401
R7922 VSS.n4381 VSS.n4380 4.51401
R7923 VSS.n4399 VSS.n4398 4.51401
R7924 VSS.n3657 VSS.n3651 4.51401
R7925 VSS.n3661 VSS.n2139 4.51401
R7926 VSS.n2937 VSS.n2148 4.51401
R7927 VSS.n2153 VSS.n2152 4.51401
R7928 VSS.n2027 VSS.n2026 4.51401
R7929 VSS.n2042 VSS.n2041 4.51401
R7930 VSS.n4855 VSS.n4854 4.51401
R7931 VSS.n4850 VSS.n4849 4.51401
R7932 VSS.n4674 VSS.n4673 4.5005
R7933 VSS.n635 VSS.n617 4.5005
R7934 VSS.n910 VSS.n768 4.5005
R7935 VSS.n913 VSS.n912 4.5005
R7936 VSS.n5774 VSS.n5773 4.5005
R7937 VSS.n5772 VSS.n5771 4.5005
R7938 VSS.n5768 VSS.n5767 4.5005
R7939 VSS.n4378 VSS.n3703 4.5005
R7940 VSS.n4394 VSS.n4393 4.5005
R7941 VSS.n3704 VSS.n3700 4.5005
R7942 VSS.n3656 VSS.n3655 4.5005
R7943 VSS.n3652 VSS.n2143 4.5005
R7944 VSS.n3663 VSS.n3662 4.5005
R7945 VSS.n2936 VSS.n2935 4.5005
R7946 VSS.n2934 VSS.n2933 4.5005
R7947 VSS.n2930 VSS.n2929 4.5005
R7948 VSS.n2024 VSS.n1344 4.5005
R7949 VSS.n2037 VSS.n2036 4.5005
R7950 VSS.n1345 VSS.n1341 4.5005
R7951 VSS.n4838 VSS.n380 4.5005
R7952 VSS.n4842 VSS.n4841 4.5005
R7953 VSS.n4843 VSS.n384 4.5005
R7954 VSS.n2667 VSS.n2665 4.49412
R7955 VSS.n1911 VSS.n1910 4.49412
R7956 VSS.n1865 VSS.n1425 4.49412
R7957 VSS.n1673 VSS.n1672 4.49412
R7958 VSS.n2413 VSS.n2412 4.47602
R7959 VSS.n1098 VSS.n1097 4.43994
R7960 VSS.n2776 VSS.n2775 4.38311
R7961 VSS.n3900 VSS.n3899 4.36875
R7962 VSS.n3913 VSS.n3830 4.36875
R7963 VSS.n4478 VSS.n4428 4.36875
R7964 VSS.n4471 VSS.n4431 4.36875
R7965 VSS.n3188 VSS.n3187 4.36875
R7966 VSS.n3177 VSS.n3176 4.36875
R7967 VSS.n3195 VSS.n3194 4.36875
R7968 VSS.n3171 VSS.n3169 4.36875
R7969 VSS.n3208 VSS.n3164 4.36875
R7970 VSS.n3201 VSS.n3167 4.36875
R7971 VSS.n2388 VSS.n2318 4.36875
R7972 VSS.n4384 VSS.n3705 4.35795
R7973 VSS.n3643 VSS.n2943 4.35795
R7974 VSS.n3551 VSS.n2988 4.35795
R7975 VSS.n3529 VSS.n3528 4.35795
R7976 VSS.n3499 VSS.n3498 4.35795
R7977 VSS.n3491 VSS.n3490 4.35795
R7978 VSS.n2632 VSS.n2199 4.35795
R7979 VSS.n3223 VSS.n3222 4.31354
R7980 VSS.n3883 VSS.n3882 4.29369
R7981 VSS.n5751 VSS.n5750 4.28986
R7982 VSS.n5706 VSS.n5705 4.28986
R7983 VSS.n5687 VSS.n5686 4.28986
R7984 VSS.n5570 VSS.n97 4.28986
R7985 VSS.n5465 VSS.n142 4.28986
R7986 VSS.n3289 VSS.n3288 4.28986
R7987 VSS.n3109 VSS.n3107 4.28986
R7988 VSS.n2632 VSS.n2631 4.28986
R7989 VSS.n1869 VSS.n1868 4.28986
R7990 VSS.n290 VSS.n288 4.28986
R7991 VSS.n282 VSS.n280 4.28986
R7992 VSS.n5055 VSS.n5054 4.28986
R7993 VSS.n261 VSS.n259 4.28986
R7994 VSS.n5158 VSS.n5157 4.28986
R7995 VSS.n5146 VSS.n5145 4.28986
R7996 VSS.n1185 VSS.n1107 4.18141
R7997 VSS.n4070 VSS.n4069 4.14168
R7998 VSS.n3368 VSS.n3367 4.14168
R7999 VSS.n3259 VSS.n3118 4.14168
R8000 VSS.n2446 VSS.n2445 4.14168
R8001 VSS.n4575 VSS.n4560 4.11798
R8002 VSS.n4578 VSS.n4560 4.11798
R8003 VSS.n5720 VSS.n5719 4.11798
R8004 VSS.n5719 VSS.n28 4.11798
R8005 VSS.n5631 VSS.n70 4.11798
R8006 VSS.n5634 VSS.n70 4.11798
R8007 VSS.n5542 VSS.n5541 4.11798
R8008 VSS.n5543 VSS.n5542 4.11798
R8009 VSS.n5446 VSS.n149 4.11798
R8010 VSS.n5449 VSS.n149 4.11798
R8011 VSS.n5410 VSS.n5409 4.11798
R8012 VSS.n5411 VSS.n5410 4.11798
R8013 VSS.n4334 VSS.n4333 4.11798
R8014 VSS.n4335 VSS.n4334 4.11798
R8015 VSS.n2112 VSS.n2075 4.11798
R8016 VSS.n2574 VSS.n2222 4.11798
R8017 VSS.n2525 VSS.n2524 4.11798
R8018 VSS.n2526 VSS.n2525 4.11798
R8019 VSS.n2424 VSS.n2306 4.11798
R8020 VSS.n2427 VSS.n2306 4.11798
R8021 VSS.n2768 VSS.n2175 4.11798
R8022 VSS.n2914 VSS.n2160 4.11798
R8023 VSS.n2911 VSS.n2160 4.11798
R8024 VSS.n1311 VSS.n1310 4.11798
R8025 VSS.n1310 VSS.n1309 4.11798
R8026 VSS.n4275 VSS.n4273 4.07962
R8027 VSS.n5752 VSS.n5751 4.07323
R8028 VSS.n5707 VSS.n5706 4.07323
R8029 VSS.n5688 VSS.n5687 4.07323
R8030 VSS.n5573 VSS.n97 4.07323
R8031 VSS.n5468 VSS.n142 4.07323
R8032 VSS.n3242 VSS.n3128 4.07323
R8033 VSS.n2838 VSS.n2165 4.07323
R8034 VSS.n2630 VSS.n2629 4.07323
R8035 VSS.n2631 VSS.n2630 4.07323
R8036 VSS.n1870 VSS.n1869 4.07323
R8037 VSS.n291 VSS.n290 4.07323
R8038 VSS.n283 VSS.n282 4.07323
R8039 VSS.n5054 VSS.n5053 4.07323
R8040 VSS.n262 VSS.n261 4.07323
R8041 VSS.n5159 VSS.n5158 4.07323
R8042 VSS.n5145 VSS.n5137 4.07323
R8043 VSS.n4729 VSS.t3299 4.03712
R8044 VSS.n4730 VSS.t3266 4.03712
R8045 VSS.n4731 VSS.t3310 4.03712
R8046 VSS.n4732 VSS.t3306 4.03712
R8047 VSS.n4733 VSS.t3323 4.03712
R8048 VSS.n4734 VSS.t3259 4.03712
R8049 VSS.n4735 VSS.t3269 4.03712
R8050 VSS.n4736 VSS.t3290 4.03712
R8051 VSS.n4737 VSS.t3261 4.03712
R8052 VSS.n4738 VSS.t3293 4.03712
R8053 VSS.n4739 VSS.t3303 4.03712
R8054 VSS.n4740 VSS.t3330 4.03712
R8055 VSS.n4741 VSS.t3267 4.03712
R8056 VSS.n4742 VSS.t3314 4.03712
R8057 VSS.n4743 VSS.t3315 4.03712
R8058 VSS.n4744 VSS.t3321 4.03712
R8059 VSS.n4694 VSS.t3309 4.03712
R8060 VSS.n4693 VSS.t3291 4.03712
R8061 VSS.n4692 VSS.t3322 4.03712
R8062 VSS.n4691 VSS.t3294 4.03712
R8063 VSS.n4690 VSS.t3311 4.03712
R8064 VSS.n4689 VSS.t3258 4.03712
R8065 VSS.n4688 VSS.t3297 4.03712
R8066 VSS.n4687 VSS.t3304 4.03712
R8067 VSS.n4686 VSS.t3253 4.03712
R8068 VSS.n4685 VSS.t3308 4.03712
R8069 VSS.n4684 VSS.t3307 4.03712
R8070 VSS.n4683 VSS.t3328 4.03712
R8071 VSS.n4682 VSS.t3329 4.03712
R8072 VSS.n4681 VSS.t3254 4.03712
R8073 VSS.n4680 VSS.t3318 4.03712
R8074 VSS.n4679 VSS.t3320 4.03712
R8075 VSS.n547 VSS.t3319 4.03712
R8076 VSS.n618 VSS.t3270 4.03712
R8077 VSS.n619 VSS.t3313 4.03712
R8078 VSS.n620 VSS.t3295 4.03712
R8079 VSS.n621 VSS.t3298 4.03712
R8080 VSS.n622 VSS.t3300 4.03712
R8081 VSS.n623 VSS.t3316 4.03712
R8082 VSS.n624 VSS.t3255 4.03712
R8083 VSS.n625 VSS.t3326 4.03712
R8084 VSS.n626 VSS.t3289 4.03712
R8085 VSS.n627 VSS.t3312 4.03712
R8086 VSS.n628 VSS.t3260 4.03712
R8087 VSS.n629 VSS.t3324 4.03712
R8088 VSS.n630 VSS.t3305 4.03712
R8089 VSS.n631 VSS.t3331 4.03712
R8090 VSS.n632 VSS.t3296 4.03712
R8091 VSS.n633 VSS.t2300 4.03712
R8092 VSS.n4761 VSS.t3325 4.03712
R8093 VSS.n4760 VSS.t3263 4.03712
R8094 VSS.n4759 VSS.t3301 4.03712
R8095 VSS.n4758 VSS.t3257 4.03712
R8096 VSS.n4757 VSS.t3327 4.03712
R8097 VSS.n4756 VSS.t3288 4.03712
R8098 VSS.n4755 VSS.t3317 4.03712
R8099 VSS.n4754 VSS.t3287 4.03712
R8100 VSS.n4753 VSS.t3265 4.03712
R8101 VSS.n4752 VSS.t3292 4.03712
R8102 VSS.n4751 VSS.t3302 4.03712
R8103 VSS.n4750 VSS.t3252 4.03712
R8104 VSS.n4749 VSS.t3262 4.03712
R8105 VSS.n4748 VSS.t3264 4.03712
R8106 VSS.n4747 VSS.t3268 4.03712
R8107 VSS.n4746 VSS.t3256 4.03712
R8108 VSS.n891 VSS.t3355 4.03712
R8109 VSS.n892 VSS.t3354 4.03712
R8110 VSS.n893 VSS.t3349 4.03712
R8111 VSS.n894 VSS.t3388 4.03712
R8112 VSS.n895 VSS.t3373 4.03712
R8113 VSS.n896 VSS.t3372 4.03712
R8114 VSS.n897 VSS.t3387 4.03712
R8115 VSS.n898 VSS.t3336 4.03712
R8116 VSS.n899 VSS.t3377 4.03712
R8117 VSS.n900 VSS.t3339 4.03712
R8118 VSS.n901 VSS.t3378 4.03712
R8119 VSS.n902 VSS.t3342 4.03712
R8120 VSS.n903 VSS.t3356 4.03712
R8121 VSS.n904 VSS.t3394 4.03712
R8122 VSS.n905 VSS.t3338 4.03712
R8123 VSS.n906 VSS.t3352 4.03712
R8124 VSS.n787 VSS.t3389 4.03712
R8125 VSS.n786 VSS.t3360 4.03712
R8126 VSS.n785 VSS.t3366 4.03712
R8127 VSS.n784 VSS.t3361 4.03712
R8128 VSS.n783 VSS.t3358 4.03712
R8129 VSS.n782 VSS.t3375 4.03712
R8130 VSS.n781 VSS.t3393 4.03712
R8131 VSS.n780 VSS.t3391 4.03712
R8132 VSS.n779 VSS.t3368 4.03712
R8133 VSS.n778 VSS.t3374 4.03712
R8134 VSS.n777 VSS.t3367 4.03712
R8135 VSS.n776 VSS.t3357 4.03712
R8136 VSS.n775 VSS.t3376 4.03712
R8137 VSS.n774 VSS.t3384 4.03712
R8138 VSS.n773 VSS.t3363 4.03712
R8139 VSS.n772 VSS.t3395 4.03712
R8140 VSS.n771 VSS.t2328 4.03712
R8141 VSS.n479 VSS.t3381 4.03712
R8142 VSS.n480 VSS.t3380 4.03712
R8143 VSS.n481 VSS.t3364 4.03712
R8144 VSS.n482 VSS.t3382 4.03712
R8145 VSS.n483 VSS.t3369 4.03712
R8146 VSS.n484 VSS.t3392 4.03712
R8147 VSS.n485 VSS.t3348 4.03712
R8148 VSS.n486 VSS.t3346 4.03712
R8149 VSS.n487 VSS.t3350 4.03712
R8150 VSS.n488 VSS.t3359 4.03712
R8151 VSS.n489 VSS.t3333 4.03712
R8152 VSS.n490 VSS.t3383 4.03712
R8153 VSS.n491 VSS.t3371 4.03712
R8154 VSS.n492 VSS.t3343 4.03712
R8155 VSS.n493 VSS.t3337 4.03712
R8156 VSS.n494 VSS.t3341 4.03712
R8157 VSS.n543 VSS.t3353 4.03712
R8158 VSS.n542 VSS.t3386 4.03712
R8159 VSS.n541 VSS.t3347 4.03712
R8160 VSS.n540 VSS.t3345 4.03712
R8161 VSS.n539 VSS.t3370 4.03712
R8162 VSS.n538 VSS.t3365 4.03712
R8163 VSS.n537 VSS.t3362 4.03712
R8164 VSS.n536 VSS.t3385 4.03712
R8165 VSS.n535 VSS.t3344 4.03712
R8166 VSS.n534 VSS.t3335 4.03712
R8167 VSS.n533 VSS.t3390 4.03712
R8168 VSS.n532 VSS.t3351 4.03712
R8169 VSS.n531 VSS.t3379 4.03712
R8170 VSS.n530 VSS.t3334 4.03712
R8171 VSS.n529 VSS.t3332 4.03712
R8172 VSS.n528 VSS.t3340 4.03712
R8173 VSS.n2764 VSS.n2175 4.02847
R8174 VSS.n3881 VSS.n3841 3.9839
R8175 VSS.n4762 VSS.t2342 3.98193
R8176 VSS.n4696 VSS.t2441 3.98193
R8177 VSS.n889 VSS.t2437 3.98193
R8178 VSS.n527 VSS.t2548 3.98193
R8179 VSS.n4467 VSS.n4466 3.97459
R8180 VSS.n3885 VSS.n3838 3.96548
R8181 VSS.n3889 VSS.n3838 3.96548
R8182 VSS.n4486 VSS.n4485 3.96548
R8183 VSS.n1614 VSS.n1539 3.96548
R8184 VSS.n1323 VSS.n1263 3.96548
R8185 VSS.n1319 VSS.n1263 3.96548
R8186 VSS.n4763 VSS.t2396 3.92851
R8187 VSS.n4764 VSS.t2485 3.92851
R8188 VSS.n4765 VSS.t2425 3.92851
R8189 VSS.n4766 VSS.t2433 3.92851
R8190 VSS.n4767 VSS.t2473 3.92851
R8191 VSS.n4768 VSS.t2318 3.92851
R8192 VSS.n4769 VSS.t2304 3.92851
R8193 VSS.n4770 VSS.t2504 3.92851
R8194 VSS.n4771 VSS.t2364 3.92851
R8195 VSS.n4772 VSS.t2522 3.92851
R8196 VSS.n4773 VSS.t2348 3.92851
R8197 VSS.n4774 VSS.t2435 3.92851
R8198 VSS.n4775 VSS.t2427 3.92851
R8199 VSS.n4776 VSS.t2366 3.92851
R8200 VSS.n4777 VSS.t2506 3.92851
R8201 VSS.n4778 VSS.t2510 3.92851
R8202 VSS.n4779 VSS.t2398 3.92851
R8203 VSS.n4780 VSS.t2423 3.92851
R8204 VSS.n4781 VSS.t2534 3.92851
R8205 VSS.n4782 VSS.t2314 3.92851
R8206 VSS.n4783 VSS.t2487 3.92851
R8207 VSS.n4784 VSS.t2286 3.92851
R8208 VSS.n4785 VSS.t2362 3.92851
R8209 VSS.n4786 VSS.t2469 3.92851
R8210 VSS.n4787 VSS.t2356 3.92851
R8211 VSS.n4788 VSS.t2463 3.92851
R8212 VSS.n4789 VSS.t2290 3.92851
R8213 VSS.n4790 VSS.t2496 3.92851
R8214 VSS.n4791 VSS.t2374 3.92851
R8215 VSS.n4792 VSS.t2520 3.92851
R8216 VSS.n4793 VSS.t2306 3.92851
R8217 VSS.n4794 VSS.t2445 3.92851
R8218 VSS.n4728 VSS.t2502 3.92851
R8219 VSS.n4727 VSS.t2410 3.92851
R8220 VSS.n4726 VSS.t2360 3.92851
R8221 VSS.n4725 VSS.t2376 3.92851
R8222 VSS.n4724 VSS.t2392 3.92851
R8223 VSS.n4723 VSS.t2278 3.92851
R8224 VSS.n4722 VSS.t2532 3.92851
R8225 VSS.n4721 VSS.t2429 3.92851
R8226 VSS.n4720 VSS.t2447 3.92851
R8227 VSS.n4719 VSS.t2382 3.92851
R8228 VSS.n4718 VSS.t2368 3.92851
R8229 VSS.n4717 VSS.t2400 3.92851
R8230 VSS.n4716 VSS.t2538 3.92851
R8231 VSS.n4715 VSS.t2459 3.92851
R8232 VSS.n4714 VSS.t2282 3.92851
R8233 VSS.n4713 VSS.t2412 3.92851
R8234 VSS.n4712 VSS.t2453 3.92851
R8235 VSS.n4711 VSS.t2406 3.92851
R8236 VSS.n4710 VSS.t2340 3.92851
R8237 VSS.n4709 VSS.t2477 3.92851
R8238 VSS.n4708 VSS.t2404 3.92851
R8239 VSS.n4707 VSS.t2451 3.92851
R8240 VSS.n4706 VSS.t2544 3.92851
R8241 VSS.n4705 VSS.t2512 3.92851
R8242 VSS.n4704 VSS.t2492 3.92851
R8243 VSS.n4703 VSS.t2475 3.92851
R8244 VSS.n4702 VSS.t2408 3.92851
R8245 VSS.n4701 VSS.t2481 3.92851
R8246 VSS.n4700 VSS.t2530 3.92851
R8247 VSS.n4699 VSS.t2394 3.92851
R8248 VSS.n4698 VSS.t2449 3.92851
R8249 VSS.n4697 VSS.t2358 3.92851
R8250 VSS.n857 VSS.t2554 3.92851
R8251 VSS.n858 VSS.t2308 3.92851
R8252 VSS.n859 VSS.t2498 3.92851
R8253 VSS.n860 VSS.t2316 3.92851
R8254 VSS.n861 VSS.t2350 3.92851
R8255 VSS.n862 VSS.t2457 3.92851
R8256 VSS.n863 VSS.t2386 3.92851
R8257 VSS.n864 VSS.t2508 3.92851
R8258 VSS.n865 VSS.t2443 3.92851
R8259 VSS.n866 VSS.t2312 3.92851
R8260 VSS.n867 VSS.t2346 3.92851
R8261 VSS.n868 VSS.t2439 3.92851
R8262 VSS.n869 VSS.t2500 3.92851
R8263 VSS.n870 VSS.t2384 3.92851
R8264 VSS.n871 VSS.t2334 3.92851
R8265 VSS.n872 VSS.t2322 3.92851
R8266 VSS.n873 VSS.t2284 3.92851
R8267 VSS.n874 VSS.t2471 3.92851
R8268 VSS.n875 VSS.t2546 3.92851
R8269 VSS.n876 VSS.t2326 3.92851
R8270 VSS.n877 VSS.t2336 3.92851
R8271 VSS.n878 VSS.t2550 3.92851
R8272 VSS.n879 VSS.t2402 3.92851
R8273 VSS.n880 VSS.t2302 3.92851
R8274 VSS.n881 VSS.t2526 3.92851
R8275 VSS.n882 VSS.t2414 3.92851
R8276 VSS.n883 VSS.t2380 3.92851
R8277 VSS.n884 VSS.t2320 3.92851
R8278 VSS.n885 VSS.t2479 3.92851
R8279 VSS.n886 VSS.t2294 3.92851
R8280 VSS.n887 VSS.t2332 3.92851
R8281 VSS.n888 VSS.t2461 3.92851
R8282 VSS.n495 VSS.t2514 3.92851
R8283 VSS.n496 VSS.t2296 3.92851
R8284 VSS.n497 VSS.t2524 3.92851
R8285 VSS.n498 VSS.t2528 3.92851
R8286 VSS.n499 VSS.t2494 3.92851
R8287 VSS.n500 VSS.t2292 3.92851
R8288 VSS.n501 VSS.t2465 3.92851
R8289 VSS.n502 VSS.t2455 3.92851
R8290 VSS.n503 VSS.t2330 3.92851
R8291 VSS.n504 VSS.t2354 3.92851
R8292 VSS.n505 VSS.t2467 3.92851
R8293 VSS.n506 VSS.t2390 3.92851
R8294 VSS.n507 VSS.t2540 3.92851
R8295 VSS.n508 VSS.t2338 3.92851
R8296 VSS.n509 VSS.t2542 3.92851
R8297 VSS.n510 VSS.t2536 3.92851
R8298 VSS.n511 VSS.t2344 3.92851
R8299 VSS.n512 VSS.t2298 3.92851
R8300 VSS.n513 VSS.t2324 3.92851
R8301 VSS.n514 VSS.t2516 3.92851
R8302 VSS.n515 VSS.t2372 3.92851
R8303 VSS.n516 VSS.t2483 3.92851
R8304 VSS.n517 VSS.t2310 3.92851
R8305 VSS.n518 VSS.t2352 3.92851
R8306 VSS.n519 VSS.t2288 3.92851
R8307 VSS.n520 VSS.t2421 3.92851
R8308 VSS.n521 VSS.t2388 3.92851
R8309 VSS.n522 VSS.t2552 3.92851
R8310 VSS.n523 VSS.t2419 3.92851
R8311 VSS.n524 VSS.t2370 3.92851
R8312 VSS.n525 VSS.t2518 3.92851
R8313 VSS.n526 VSS.t2280 3.92851
R8314 VSS.n1083 VSS.n1082 3.91766
R8315 VSS.n2071 VSS.n2070 3.90948
R8316 VSS.n2557 VSS.n2232 3.90948
R8317 VSS.n3636 VSS.n3635 3.76521
R8318 VSS.n2649 VSS.n2648 3.76521
R8319 VSS.n2077 VSS.n2075 3.75994
R8320 VSS.n2414 VSS.n2413 3.75994
R8321 VSS.n4329 VSS.n4327 3.7575
R8322 VSS.n4631 VSS.n4630 3.73795
R8323 VSS.n3885 VSS.n3884 3.7069
R8324 VSS.n4486 VSS.n4425 3.7069
R8325 VSS.n3237 VSS.n3236 3.7069
R8326 VSS.n3238 VSS.n3237 3.7069
R8327 VSS.n1609 VSS.n1607 3.7069
R8328 VSS.n1324 VSS.n1323 3.7069
R8329 VSS.n1319 VSS.n1318 3.7069
R8330 VSS.n2606 VSS.n2605 3.6771
R8331 VSS.n3239 VSS.n3128 3.56523
R8332 VSS.n3587 VSS.n2968 3.54833
R8333 VSS.n2778 VSS.n2777 3.54833
R8334 VSS.n1892 VSS.n1891 3.54833
R8335 VSS.n614 VSS.n613 3.51847
R8336 VSS.n854 VSS.n853 3.51847
R8337 VSS.n5665 VSS.n55 3.50735
R8338 VSS.n5482 VSS.n133 3.50735
R8339 VSS.n3936 VSS.n3823 3.50735
R8340 VSS.n4083 VSS.n3797 3.50735
R8341 VSS.n3607 VSS.n2964 3.50735
R8342 VSS.n3358 VSS.n3357 3.50735
R8343 VSS.n2638 VSS.n2637 3.50735
R8344 VSS.n1918 VSS.n1917 3.50735
R8345 VSS.n2575 VSS.n2574 3.49141
R8346 VSS.n2378 VSS.n2377 3.44377
R8347 VSS.n2896 VSS.n2895 3.44377
R8348 VSS.n7 VSS.n0 3.43925
R8349 VSS.n5776 VSS.n5775 3.43925
R8350 VSS.n4398 VSS.n4397 3.43925
R8351 VSS.n4380 VSS.n4379 3.43925
R8352 VSS.n3661 VSS.n3660 3.43925
R8353 VSS.n3658 VSS.n3657 3.43925
R8354 VSS.n2152 VSS.n2146 3.43925
R8355 VSS.n2938 VSS.n2937 3.43925
R8356 VSS.n2041 VSS.n2040 3.43925
R8357 VSS.n2026 VSS.n2025 3.43925
R8358 VSS.n4851 VSS.n4850 3.43925
R8359 VSS.n4854 VSS.n4853 3.43925
R8360 VSS.n4981 VSS.n308 3.42526
R8361 VSS.n701 VSS.n635 3.41856
R8362 VSS.n768 VSS.n767 3.41856
R8363 VSS.n4673 VSS.n4672 3.4105
R8364 VSS.n914 VSS.n913 3.4105
R8365 VSS.n4 VSS.n2 3.4105
R8366 VSS.n5770 VSS.n5769 3.4105
R8367 VSS.n3702 VSS.n3701 3.4105
R8368 VSS.n4396 VSS.n4395 3.4105
R8369 VSS.n3653 VSS.n2940 3.4105
R8370 VSS.n2145 VSS.n2144 3.4105
R8371 VSS.n2149 VSS.n2147 3.4105
R8372 VSS.n2932 VSS.n2931 3.4105
R8373 VSS.n1343 VSS.n1342 3.4105
R8374 VSS.n2039 VSS.n2038 3.4105
R8375 VSS.n4839 VSS.n381 3.4105
R8376 VSS.n4840 VSS.n383 3.4105
R8377 VSS.n2898 VSS.n2838 3.40077
R8378 VSS.n3462 VSS.n3461 3.38874
R8379 VSS.n2597 VSS.n2214 3.38874
R8380 VSS.n2503 VSS.n2502 3.38874
R8381 VSS.n1819 VSS.n1447 3.38874
R8382 VSS.n4048 VSS.n4047 3.26859
R8383 VSS.n4989 VSS.t774 3.26073
R8384 VSS.n969 VSS.n963 3.21999
R8385 VSS.n2377 VSS.n2322 3.21921
R8386 VSS.n2380 VSS.n2320 3.21921
R8387 VSS.n2897 VSS.n2896 3.21921
R8388 VSS.n2892 VSS.n2891 3.21921
R8389 VSS.n5666 VSS.n53 3.2005
R8390 VSS.n5483 VSS.n131 3.2005
R8391 VSS.n3937 VSS.n3821 3.2005
R8392 VSS.n4084 VSS.n3795 3.2005
R8393 VSS.n3608 VSS.n2962 3.2005
R8394 VSS.n3363 VSS.n3075 3.2005
R8395 VSS.n3301 VSS.n3097 3.2005
R8396 VSS.n2886 VSS.n2885 3.2005
R8397 VSS.n1922 VSS.n1397 3.2005
R8398 VSS.n3894 VSS.n3893 3.13337
R8399 VSS.n5617 VSS.n5616 3.13241
R8400 VSS.n5561 VSS.n5560 3.13241
R8401 VSS.n5526 VSS.n5525 3.13241
R8402 VSS.n5432 VSS.n5431 3.13241
R8403 VSS.n4109 VSS.n4108 3.13241
R8404 VSS.n4225 VSS.n4224 3.13241
R8405 VSS.n4314 VSS.n4313 3.13241
R8406 VSS.n3471 VSS.n3470 3.13241
R8407 VSS.n3454 VSS.n3453 3.13241
R8408 VSS.n3394 VSS.n3393 3.13241
R8409 VSS.n3286 VSS.n3285 3.13241
R8410 VSS.n3279 VSS.n3278 3.13241
R8411 VSS.n2609 VSS.n2608 3.13241
R8412 VSS.n2460 VSS.n2459 3.13241
R8413 VSS.n2717 VSS.n2716 3.13241
R8414 VSS.n2703 VSS.n2675 3.13241
R8415 VSS.n2063 VSS.n2062 3.13241
R8416 VSS.n4874 VSS.n4873 3.13241
R8417 VSS.n5116 VSS.n238 3.13241
R8418 VSS.n230 VSS.n228 3.13241
R8419 VSS.n5203 VSS.n222 3.13241
R8420 VSS.n5221 VSS.n214 3.13241
R8421 VSS.n5238 VSS.n5237 3.13241
R8422 VSS.n456 VSS.n455 3.13241
R8423 VSS.n3295 VSS.n3100 3.11283
R8424 VSS.n2906 VSS.n2903 3.06137
R8425 VSS.n4468 VSS.n4467 3.05276
R8426 VSS.n2900 VSS.n2165 3.04861
R8427 VSS.n5468 VSS.n5467 3.04861
R8428 VSS.n5573 VSS.n5572 3.04861
R8429 VSS.n5689 VSS.n5688 3.04861
R8430 VSS.n5707 VSS.n33 3.04861
R8431 VSS.n5753 VSS.n5752 3.04861
R8432 VSS.n3881 VSS.n3880 3.04861
R8433 VSS.n2126 VSS.n2125 3.04861
R8434 VSS.n3242 VSS.n3241 3.04861
R8435 VSS.n2386 VSS.n2319 3.04861
R8436 VSS.n2630 VSS.n2200 3.04861
R8437 VSS.n1870 VSS.n1422 3.04861
R8438 VSS.n5148 VSS.n5137 3.04861
R8439 VSS.n5160 VSS.n5159 3.04861
R8440 VSS.n5065 VSS.n262 3.04861
R8441 VSS.n5053 VSS.n5052 3.04861
R8442 VSS.n5020 VSS.n283 3.04861
R8443 VSS.n5006 VSS.n291 3.04861
R8444 VSS.n2417 VSS.n2416 3.04386
R8445 VSS.n4329 VSS.n4328 3.01483
R8446 VSS.n1665 VSS.n1664 3.01226
R8447 VSS.n1095 VSS.n1094 3.01194
R8448 VSS.n4047 VSS.n4046 2.99624
R8449 VSS.n2122 VSS.n2071 2.9514
R8450 VSS.n2558 VSS.n2557 2.9514
R8451 VSS.n959 VSS.n324 2.93224
R8452 VSS.n3882 VSS.n3881 2.92166
R8453 VSS.n3891 VSS.n3889 2.88804
R8454 VSS.n1615 VSS.n1614 2.88804
R8455 VSS.n2125 VSS.n2121 2.86855
R8456 VSS.n2387 VSS.n2386 2.86855
R8457 VSS.n3891 VSS.n3890 2.83202
R8458 VSS.n4981 VSS.n4980 2.82936
R8459 VSS.n2889 VSS.n2841 2.76214
R8460 VSS.n2639 VSS.n2194 2.76214
R8461 VSS.n5618 VSS.n5617 2.7239
R8462 VSS.n5562 VSS.n5561 2.7239
R8463 VSS.n5527 VSS.n5526 2.7239
R8464 VSS.n5433 VSS.n5432 2.7239
R8465 VSS.n4108 VSS.n3781 2.7239
R8466 VSS.n4224 VSS.n4223 2.7239
R8467 VSS.n4315 VSS.n4314 2.7239
R8468 VSS.n3472 VSS.n3471 2.7239
R8469 VSS.n3455 VSS.n3454 2.7239
R8470 VSS.n3395 VSS.n3394 2.7239
R8471 VSS.n2608 VSS.n2607 2.7239
R8472 VSS.n2459 VSS.n2284 2.7239
R8473 VSS.n2716 VSS.n2715 2.7239
R8474 VSS.n2677 VSS.n2675 2.7239
R8475 VSS.n2749 VSS.n2748 2.7239
R8476 VSS.n2062 VSS.n1332 2.7239
R8477 VSS.n4873 VSS.n4872 2.7239
R8478 VSS.n240 VSS.n238 2.7239
R8479 VSS.n231 VSS.n230 2.7239
R8480 VSS.n224 VSS.n222 2.7239
R8481 VSS.n216 VSS.n214 2.7239
R8482 VSS.n5237 VSS.n5236 2.7239
R8483 VSS.n455 VSS.n454 2.7239
R8484 VSS.n3971 VSS.n3970 2.63579
R8485 VSS.n4037 VSS.n4036 2.63579
R8486 VSS.n4123 VSS.n4122 2.63579
R8487 VSS.n4390 VSS.n4389 2.63579
R8488 VSS.n3649 VSS.n3648 2.63579
R8489 VSS.n3557 VSS.n3556 2.63579
R8490 VSS.n3534 VSS.n2995 2.63579
R8491 VSS.n3383 VSS.n3065 2.63579
R8492 VSS.n3251 VSS.n3250 2.63579
R8493 VSS.n2615 VSS.n2205 2.63579
R8494 VSS.n2826 VSS.n2825 2.63579
R8495 VSS.n2033 VSS.n2031 2.63579
R8496 VSS.n2019 VSS.n1350 2.63579
R8497 VSS.n2003 VSS.n1358 2.63579
R8498 VSS.n1961 VSS.n1377 2.63579
R8499 VSS.n1767 VSS.n1476 2.63579
R8500 VSS.n1715 VSS.n1712 2.63579
R8501 VSS.n1656 VSS.n1524 2.63579
R8502 VSS.n1144 VSS.n1140 2.63064
R8503 VSS.n5669 VSS.n5668 2.63064
R8504 VSS.n5486 VSS.n5485 2.63064
R8505 VSS.n3940 VSS.n3939 2.63064
R8506 VSS.n4087 VSS.n4086 2.63064
R8507 VSS.n3361 VSS.n3076 2.63064
R8508 VSS.n3304 VSS.n3303 2.63064
R8509 VSS.n2846 VSS.n2842 2.63064
R8510 VSS.n2641 VSS.n2195 2.63064
R8511 VSS.n4663 VSS.n4662 2.63064
R8512 VSS.n2609 VSS.n2606 2.58773
R8513 VSS.n1171 VSS.n1169 2.5605
R8514 VSS.n4801 VSS.n474 2.5605
R8515 VSS.t444 VSS.t445 2.53433
R8516 VSS.t559 VSS.t552 2.53433
R8517 VSS.n2508 VSS.n2253 2.50679
R8518 VSS.n4632 VSS.t89 2.49271
R8519 VSS.n1134 VSS.t260 2.4755
R8520 VSS.n1134 VSS.t250 2.4755
R8521 VSS.n1132 VSS.t258 2.4755
R8522 VSS.n1132 VSS.t252 2.4755
R8523 VSS.n1130 VSS.t254 2.4755
R8524 VSS.n1130 VSS.t256 2.4755
R8525 VSS.n1128 VSS.t248 2.4755
R8526 VSS.n1128 VSS.t308 2.4755
R8527 VSS.n1126 VSS.t314 2.4755
R8528 VSS.n1126 VSS.t310 2.4755
R8529 VSS.n1124 VSS.t312 2.4755
R8530 VSS.n1124 VSS.t453 2.4755
R8531 VSS.n1122 VSS.t451 2.4755
R8532 VSS.n1122 VSS.t2879 2.4755
R8533 VSS.n916 VSS.t3272 2.4755
R8534 VSS.n916 VSS.t3280 2.4755
R8535 VSS.n934 VSS.t3284 2.4755
R8536 VSS.n934 VSS.t3278 2.4755
R8537 VSS.n932 VSS.t3274 2.4755
R8538 VSS.n932 VSS.t3282 2.4755
R8539 VSS.n930 VSS.t367 2.4755
R8540 VSS.n930 VSS.t3276 2.4755
R8541 VSS.n928 VSS.t373 2.4755
R8542 VSS.n928 VSS.t369 2.4755
R8543 VSS.n926 VSS.t2797 2.4755
R8544 VSS.n926 VSS.t371 2.4755
R8545 VSS.n924 VSS.t2826 2.4755
R8546 VSS.n924 VSS.t2795 2.4755
R8547 VSS.n3583 VSS.n2968 2.43528
R8548 VSS.n1158 VSS.n1157 2.40002
R8549 VSS.n4635 VSS.n937 2.39867
R8550 VSS.n4276 VSS.n4275 2.39171
R8551 VSS.n1617 VSS.n1616 2.36572
R8552 VSS.n1097 VSS.n1096 2.341
R8553 VSS.n3907 VSS.n3832 2.33701
R8554 VSS.n3910 VSS.n3832 2.33701
R8555 VSS.n3911 VSS.n3910 2.33701
R8556 VSS.n3912 VSS.n3911 2.33701
R8557 VSS.n4476 VSS.n4429 2.33701
R8558 VSS.n4473 VSS.n4429 2.33701
R8559 VSS.n3183 VSS.n3182 2.33701
R8560 VSS.n3182 VSS.n3181 2.33701
R8561 VSS.n3206 VSS.n3165 2.33701
R8562 VSS.n3203 VSS.n3165 2.33701
R8563 VSS.n2395 VSS.n2316 2.33701
R8564 VSS.n2398 VSS.n2316 2.33701
R8565 VSS.n2402 VSS.n2401 2.33701
R8566 VSS.n2429 VSS.n2428 2.32777
R8567 VSS.n3307 VSS.n3306 2.25932
R8568 VSS.n2501 VSS.n2500 2.25932
R8569 VSS.n3892 VSS.n3837 2.25312
R8570 VSS.n2127 VSS.n2071 2.25312
R8571 VSS.n2557 VSS.n2231 2.25293
R8572 VSS.n314 VSS.n313 2.1939
R8573 VSS.n3893 VSS.n3892 2.13383
R8574 VSS.n3955 VSS.n3954 2.13383
R8575 VSS.n3577 VSS.n2977 2.13383
R8576 VSS.n2748 VSS.n2747 2.11114
R8577 VSS.n1399 VSS.n1395 2.10461
R8578 VSS.n2401 VSS.n2400 2.03225
R8579 VSS.n3584 VSS.n3582 2.01789
R8580 VSS.n2485 VSS.n2484 2.01789
R8581 VSS.n1986 VSS.n1366 2.01789
R8582 VSS.n1615 VSS.n1538 2.01694
R8583 VSS.n3334 VSS.n3333 2.01531
R8584 VSS.n4485 VSS.n4484 1.98299
R8585 VSS.n1609 VSS.n1608 1.98299
R8586 VSS.n1608 VSS.n1539 1.98299
R8587 VSS.n3596 VSS.n3591 1.97497
R8588 VSS.n3449 VSS.n3445 1.97497
R8589 VSS.n2712 VSS.n2668 1.97497
R8590 VSS.n2527 VSS.n2247 1.96973
R8591 VSS.n971 VSS.n969 1.91915
R8592 VSS.n4031 VSS.n4030 1.8968
R8593 VSS.n1639 VSS.n1638 1.8968
R8594 VSS.n4140 VSS.n4139 1.88285
R8595 VSS.n4147 VSS.n4146 1.88285
R8596 VSS.n4232 VSS.n4231 1.88285
R8597 VSS.n4207 VSS.n4182 1.88285
R8598 VSS.n4254 VSS.n3756 1.88285
R8599 VSS.n4405 VSS.n3696 1.88285
R8600 VSS.n3669 VSS.n3668 1.88285
R8601 VSS.n3622 VSS.n3621 1.88285
R8602 VSS.n3525 VSS.n3524 1.88285
R8603 VSS.n3481 VSS.n3480 1.88285
R8604 VSS.n2435 VSS.n2301 1.88285
R8605 VSS.n2730 VSS.n2729 1.88285
R8606 VSS.n2030 VSS.n2029 1.88285
R8607 VSS.n1954 VSS.n1953 1.88285
R8608 VSS.n1774 VSS.n1472 1.88285
R8609 VSS.n1723 VSS.n1722 1.88285
R8610 VSS.n1715 VSS.n1714 1.88285
R8611 VSS.n2906 VSS.n2905 1.87783
R8612 VSS.n4387 VSS.n3705 1.8161
R8613 VSS.n3646 VSS.n2943 1.8161
R8614 VSS.n3554 VSS.n2988 1.8161
R8615 VSS.n3529 VSS.n2997 1.8161
R8616 VSS.n3499 VSS.n3012 1.8161
R8617 VSS.n3491 VSS.n3014 1.8161
R8618 VSS.n701 VSS.n700 1.80797
R8619 VSS.n767 VSS.n766 1.80797
R8620 VSS.n2379 VSS.n2378 1.79699
R8621 VSS.n2895 VSS.n2839 1.79699
R8622 VSS.n4640 VSS.n4639 1.78315
R8623 VSS.n1180 VSS.n1179 1.78315
R8624 VSS.n1153 VSS.n1152 1.77828
R8625 VSS.n948 VSS.n941 1.77828
R8626 VSS.n1912 VSS.n1911 1.77071
R8627 VSS.n1868 VSS.n1425 1.77071
R8628 VSS.n3611 VSS.n3610 1.75392
R8629 VSS.n4484 VSS.n4483 1.72441
R8630 VSS.n4852 VSS.n4851 1.69188
R8631 VSS.n4853 VSS.n4852 1.69188
R8632 VSS.n2040 VSS.n382 1.69188
R8633 VSS.n2025 VSS.n382 1.69188
R8634 VSS.n2939 VSS.n2146 1.69188
R8635 VSS.n2939 VSS.n2938 1.69188
R8636 VSS.n3660 VSS.n3659 1.69188
R8637 VSS.n3659 VSS.n3658 1.69188
R8638 VSS.n4397 VSS.n1 1.69188
R8639 VSS.n4379 VSS.n1 1.69188
R8640 VSS.n5777 VSS.n0 1.69188
R8641 VSS.n5777 VSS.n5776 1.69188
R8642 VSS.n4446 VSS.n4445 1.6821
R8643 VSS.n2091 VSS.n2090 1.6821
R8644 VSS.n2857 VSS.n2856 1.6821
R8645 VSS.n1282 VSS.n1281 1.6821
R8646 VSS.n3855 VSS.n3854 1.6819
R8647 VSS.n3143 VSS.n3142 1.6819
R8648 VSS.n2344 VSS.n2343 1.6819
R8649 VSS.n1564 VSS.n1563 1.6819
R8650 VSS.n2380 VSS.n2379 1.64728
R8651 VSS.n2892 VSS.n2839 1.64728
R8652 VSS.n2422 VSS.n2421 1.61169
R8653 VSS.n4610 VSS.n4609 1.54533
R8654 VSS.n3330 VSS.n3329 1.54124
R8655 VSS.n2566 VSS.n2224 1.52218
R8656 VSS.n3963 VSS.n3962 1.50638
R8657 VSS.n4124 VSS.n4123 1.50638
R8658 VSS.n3152 VSS.n3151 1.50638
R8659 VSS.n2358 VSS.n2331 1.50638
R8660 VSS.n2350 VSS.n2335 1.50638
R8661 VSS.n1706 VSS.n1705 1.50638
R8662 VSS.n1580 VSS.n1579 1.50638
R8663 VSS.n1570 VSS.n1555 1.50638
R8664 VSS.n1297 VSS.n1296 1.50638
R8665 VSS.n3917 VSS.n3916 1.47352
R8666 VSS.n3198 VSS.n3197 1.46433
R8667 VSS.n1097 VSS.n1031 1.43383
R8668 VSS.n3197 VSS.n3196 1.42881
R8669 VSS.n1069 VSS.n308 1.41445
R8670 VSS.n1156 VSS.n1155 1.39283
R8671 VSS.n4666 VSS.n4665 1.39283
R8672 VSS.n2718 VSS.n2667 1.3622
R8673 VSS.n2063 VSS.n2061 1.3622
R8674 VSS.n1672 VSS.n1514 1.3622
R8675 VSS.n348 VSS.n347 1.36141
R8676 VSS.n3175 VSS.n3174 1.3469
R8677 VSS.n4980 VSS.n4979 1.32802
R8678 VSS.n1220 VSS.n978 1.32464
R8679 VSS.n2629 VSS.n2628 1.32281
R8680 VSS.n4449 VSS.n4446 1.30732
R8681 VSS.n2092 VSS.n2091 1.30732
R8682 VSS.n2857 VSS.n2853 1.30732
R8683 VSS.n1285 VSS.n1282 1.30732
R8684 VSS.n3856 VSS.n3855 1.30718
R8685 VSS.n3146 VSS.n3143 1.30718
R8686 VSS.n2345 VSS.n2344 1.30718
R8687 VSS.n1565 VSS.n1564 1.30718
R8688 VSS.n549 VSS.t2341 1.30567
R8689 VSS.n636 VSS.t2430 1.30567
R8690 VSS.n789 VSS.t2547 1.30567
R8691 VSS.n702 VSS.t2377 1.30567
R8692 VSS.n2635 VSS.n2199 1.30065
R8693 VSS.n3944 VSS.n3820 1.27173
R8694 VSS.n4338 VSS.n3721 1.25365
R8695 VSS.n2520 VSS.n2519 1.25365
R8696 VSS.n2921 VSS.n2920 1.25365
R8697 VSS.n2558 VSS.n2228 1.25267
R8698 VSS.n2777 VSS.n2776 1.25267
R8699 VSS.n1891 VSS.n1890 1.25267
R8700 VSS.n3235 VSS.n3131 1.25033
R8701 VSS.n1326 VSS.n1325 1.20723
R8702 VSS.n347 VSS.n338 1.20467
R8703 VSS.n4511 VSS.n4510 1.18311
R8704 VSS.n5740 VSS.n20 1.18311
R8705 VSS.n5589 VSS.n5588 1.18311
R8706 VSS.n5365 VSS.n5364 1.18311
R8707 VSS.n4301 VSS.n4300 1.18311
R8708 VSS.n3589 VSS.n3588 1.18311
R8709 VSS.n3405 VSS.n3055 1.18311
R8710 VSS.n3222 VSS.n3221 1.18311
R8711 VSS.n2487 VSS.n2270 1.18311
R8712 VSS.n2779 VSS.n2778 1.18311
R8713 VSS.n1992 VSS.n1991 1.18311
R8714 VSS.n1893 VSS.n1892 1.18311
R8715 VSS.n1698 VSS.n1503 1.18311
R8716 VSS.n1631 VSS.n1630 1.18311
R8717 VSS.n4823 VSS.n4822 1.18311
R8718 VSS.n5033 VSS.n5032 1.18311
R8719 VSS.n5041 VSS.n5040 1.18311
R8720 VSS.n5277 VSS.n5276 1.18311
R8721 VSS.n5291 VSS.n5290 1.18311
R8722 VSS.n5332 VSS.n5331 1.18311
R8723 VSS.n416 VSS.n415 1.18311
R8724 VSS.n3841 VSS.n3840 1.16896
R8725 VSS.n4627 VSS.t2829 1.16053
R8726 VSS.n3285 VSS.n3284 1.15795
R8727 VSS.n3278 VSS.n3277 1.15795
R8728 VSS.n4319 VSS.n3728 1.15239
R8729 VSS.n5668 VSS.n53 1.14023
R8730 VSS.n5485 VSS.n131 1.14023
R8731 VSS.n3939 VSS.n3821 1.14023
R8732 VSS.n4086 VSS.n3795 1.14023
R8733 VSS.n3610 VSS.n2962 1.14023
R8734 VSS.n3303 VSS.n3097 1.14023
R8735 VSS.n2885 VSS.n2842 1.14023
R8736 VSS.n2642 VSS.n2641 1.14023
R8737 VSS.n1922 VSS.n1921 1.14023
R8738 VSS.n2479 VSS.n2478 1.12991
R8739 VSS.n2656 VSS.n2185 1.12991
R8740 VSS.n549 VSS.t2395 1.1255
R8741 VSS.n550 VSS.t2484 1.1255
R8742 VSS.n551 VSS.t2424 1.1255
R8743 VSS.n552 VSS.t2432 1.1255
R8744 VSS.n553 VSS.t2472 1.1255
R8745 VSS.n554 VSS.t2317 1.1255
R8746 VSS.n555 VSS.t2303 1.1255
R8747 VSS.n556 VSS.t2503 1.1255
R8748 VSS.n557 VSS.t2363 1.1255
R8749 VSS.n558 VSS.t2521 1.1255
R8750 VSS.n559 VSS.t2347 1.1255
R8751 VSS.n560 VSS.t2434 1.1255
R8752 VSS.n561 VSS.t2426 1.1255
R8753 VSS.n562 VSS.t2365 1.1255
R8754 VSS.n563 VSS.t2505 1.1255
R8755 VSS.n564 VSS.t2509 1.1255
R8756 VSS.n565 VSS.t2397 1.1255
R8757 VSS.n566 VSS.t2422 1.1255
R8758 VSS.n567 VSS.t2533 1.1255
R8759 VSS.n568 VSS.t2313 1.1255
R8760 VSS.n569 VSS.t2486 1.1255
R8761 VSS.n570 VSS.t2285 1.1255
R8762 VSS.n571 VSS.t2361 1.1255
R8763 VSS.n572 VSS.t2468 1.1255
R8764 VSS.n573 VSS.t2355 1.1255
R8765 VSS.n574 VSS.t2462 1.1255
R8766 VSS.n575 VSS.t2289 1.1255
R8767 VSS.n576 VSS.t2495 1.1255
R8768 VSS.n577 VSS.t2373 1.1255
R8769 VSS.n578 VSS.t2519 1.1255
R8770 VSS.n579 VSS.t2305 1.1255
R8771 VSS.n580 VSS.t2444 1.1255
R8772 VSS.n581 VSS.t2501 1.1255
R8773 VSS.n582 VSS.t2409 1.1255
R8774 VSS.n583 VSS.t2359 1.1255
R8775 VSS.n584 VSS.t2375 1.1255
R8776 VSS.n585 VSS.t2391 1.1255
R8777 VSS.n586 VSS.t2277 1.1255
R8778 VSS.n587 VSS.t2531 1.1255
R8779 VSS.n588 VSS.t2428 1.1255
R8780 VSS.n589 VSS.t2446 1.1255
R8781 VSS.n590 VSS.t2381 1.1255
R8782 VSS.n591 VSS.t2367 1.1255
R8783 VSS.n592 VSS.t2399 1.1255
R8784 VSS.n593 VSS.t2537 1.1255
R8785 VSS.n594 VSS.t2458 1.1255
R8786 VSS.n595 VSS.t2281 1.1255
R8787 VSS.n596 VSS.t2411 1.1255
R8788 VSS.n597 VSS.t2452 1.1255
R8789 VSS.n598 VSS.t2405 1.1255
R8790 VSS.n599 VSS.t2339 1.1255
R8791 VSS.n600 VSS.t2476 1.1255
R8792 VSS.n601 VSS.t2403 1.1255
R8793 VSS.n602 VSS.t2450 1.1255
R8794 VSS.n603 VSS.t2543 1.1255
R8795 VSS.n604 VSS.t2511 1.1255
R8796 VSS.n605 VSS.t2491 1.1255
R8797 VSS.n606 VSS.t2474 1.1255
R8798 VSS.n607 VSS.t2407 1.1255
R8799 VSS.n608 VSS.t2480 1.1255
R8800 VSS.n609 VSS.t2529 1.1255
R8801 VSS.n610 VSS.t2393 1.1255
R8802 VSS.n611 VSS.t2448 1.1255
R8803 VSS.n612 VSS.t2357 1.1255
R8804 VSS.n613 VSS.t2440 1.1255
R8805 VSS.n636 VSS.t3617 1.1255
R8806 VSS.n637 VSS.t3602 1.1255
R8807 VSS.n638 VSS.t3758 1.1255
R8808 VSS.n639 VSS.t3610 1.1255
R8809 VSS.n640 VSS.t3744 1.1255
R8810 VSS.n641 VSS.t3593 1.1255
R8811 VSS.n642 VSS.t3789 1.1255
R8812 VSS.n643 VSS.t3659 1.1255
R8813 VSS.n644 VSS.t3769 1.1255
R8814 VSS.n645 VSS.t3721 1.1255
R8815 VSS.n646 VSS.t3636 1.1255
R8816 VSS.n647 VSS.t3603 1.1255
R8817 VSS.n648 VSS.t3665 1.1255
R8818 VSS.n649 VSS.t3810 1.1255
R8819 VSS.n650 VSS.t3597 1.1255
R8820 VSS.n651 VSS.t3773 1.1255
R8821 VSS.n652 VSS.t3770 1.1255
R8822 VSS.n653 VSS.t3568 1.1255
R8823 VSS.n654 VSS.t3718 1.1255
R8824 VSS.n655 VSS.t3615 1.1255
R8825 VSS.n656 VSS.t3592 1.1255
R8826 VSS.n657 VSS.t3627 1.1255
R8827 VSS.n658 VSS.t3579 1.1255
R8828 VSS.n659 VSS.t3644 1.1255
R8829 VSS.n660 VSS.t3604 1.1255
R8830 VSS.n661 VSS.t3726 1.1255
R8831 VSS.n662 VSS.t3785 1.1255
R8832 VSS.n663 VSS.t3805 1.1255
R8833 VSS.n664 VSS.t3581 1.1255
R8834 VSS.n665 VSS.t3743 1.1255
R8835 VSS.n666 VSS.t3698 1.1255
R8836 VSS.n667 VSS.t3755 1.1255
R8837 VSS.n668 VSS.t3723 1.1255
R8838 VSS.n669 VSS.t3663 1.1255
R8839 VSS.n670 VSS.t3791 1.1255
R8840 VSS.n671 VSS.t3757 1.1255
R8841 VSS.n672 VSS.t3735 1.1255
R8842 VSS.n673 VSS.t3709 1.1255
R8843 VSS.n674 VSS.t3782 1.1255
R8844 VSS.n675 VSS.t3699 1.1255
R8845 VSS.n676 VSS.t3712 1.1255
R8846 VSS.n677 VSS.t3809 1.1255
R8847 VSS.n678 VSS.t3808 1.1255
R8848 VSS.n679 VSS.t3777 1.1255
R8849 VSS.n680 VSS.t3607 1.1255
R8850 VSS.n681 VSS.t3670 1.1255
R8851 VSS.n682 VSS.t3748 1.1255
R8852 VSS.n683 VSS.t3630 1.1255
R8853 VSS.n684 VSS.t3606 1.1255
R8854 VSS.n685 VSS.t3746 1.1255
R8855 VSS.n686 VSS.t3796 1.1255
R8856 VSS.n687 VSS.t3572 1.1255
R8857 VSS.n688 VSS.t3722 1.1255
R8858 VSS.n689 VSS.t3658 1.1255
R8859 VSS.n690 VSS.t3749 1.1255
R8860 VSS.n691 VSS.t3580 1.1255
R8861 VSS.n692 VSS.t3620 1.1255
R8862 VSS.n693 VSS.t3812 1.1255
R8863 VSS.n694 VSS.t3742 1.1255
R8864 VSS.n695 VSS.t3703 1.1255
R8865 VSS.n696 VSS.t3623 1.1255
R8866 VSS.n697 VSS.t3737 1.1255
R8867 VSS.n698 VSS.t3778 1.1255
R8868 VSS.n699 VSS.t3781 1.1255
R8869 VSS.n700 VSS.t2299 1.1255
R8870 VSS.n789 VSS.t2279 1.1255
R8871 VSS.n790 VSS.t2517 1.1255
R8872 VSS.n791 VSS.t2369 1.1255
R8873 VSS.n792 VSS.t2418 1.1255
R8874 VSS.n793 VSS.t2551 1.1255
R8875 VSS.n794 VSS.t2387 1.1255
R8876 VSS.n795 VSS.t2420 1.1255
R8877 VSS.n796 VSS.t2287 1.1255
R8878 VSS.n797 VSS.t2351 1.1255
R8879 VSS.n798 VSS.t2309 1.1255
R8880 VSS.n799 VSS.t2482 1.1255
R8881 VSS.n800 VSS.t2371 1.1255
R8882 VSS.n801 VSS.t2515 1.1255
R8883 VSS.n802 VSS.t2323 1.1255
R8884 VSS.n803 VSS.t2297 1.1255
R8885 VSS.n804 VSS.t2343 1.1255
R8886 VSS.n805 VSS.t2535 1.1255
R8887 VSS.n806 VSS.t2541 1.1255
R8888 VSS.n807 VSS.t2337 1.1255
R8889 VSS.n808 VSS.t2539 1.1255
R8890 VSS.n809 VSS.t2389 1.1255
R8891 VSS.n810 VSS.t2466 1.1255
R8892 VSS.n811 VSS.t2353 1.1255
R8893 VSS.n812 VSS.t2329 1.1255
R8894 VSS.n813 VSS.t2454 1.1255
R8895 VSS.n814 VSS.t2464 1.1255
R8896 VSS.n815 VSS.t2291 1.1255
R8897 VSS.n816 VSS.t2493 1.1255
R8898 VSS.n817 VSS.t2527 1.1255
R8899 VSS.n818 VSS.t2523 1.1255
R8900 VSS.n819 VSS.t2295 1.1255
R8901 VSS.n820 VSS.t2513 1.1255
R8902 VSS.n821 VSS.t2553 1.1255
R8903 VSS.n822 VSS.t2307 1.1255
R8904 VSS.n823 VSS.t2497 1.1255
R8905 VSS.n824 VSS.t2315 1.1255
R8906 VSS.n825 VSS.t2349 1.1255
R8907 VSS.n826 VSS.t2456 1.1255
R8908 VSS.n827 VSS.t2385 1.1255
R8909 VSS.n828 VSS.t2507 1.1255
R8910 VSS.n829 VSS.t2442 1.1255
R8911 VSS.n830 VSS.t2311 1.1255
R8912 VSS.n831 VSS.t2345 1.1255
R8913 VSS.n832 VSS.t2438 1.1255
R8914 VSS.n833 VSS.t2499 1.1255
R8915 VSS.n834 VSS.t2383 1.1255
R8916 VSS.n835 VSS.t2333 1.1255
R8917 VSS.n836 VSS.t2321 1.1255
R8918 VSS.n837 VSS.t2283 1.1255
R8919 VSS.n838 VSS.t2470 1.1255
R8920 VSS.n839 VSS.t2545 1.1255
R8921 VSS.n840 VSS.t2325 1.1255
R8922 VSS.n841 VSS.t2335 1.1255
R8923 VSS.n842 VSS.t2549 1.1255
R8924 VSS.n843 VSS.t2401 1.1255
R8925 VSS.n844 VSS.t2301 1.1255
R8926 VSS.n845 VSS.t2525 1.1255
R8927 VSS.n846 VSS.t2413 1.1255
R8928 VSS.n847 VSS.t2379 1.1255
R8929 VSS.n848 VSS.t2319 1.1255
R8930 VSS.n849 VSS.t2478 1.1255
R8931 VSS.n850 VSS.t2293 1.1255
R8932 VSS.n851 VSS.t2331 1.1255
R8933 VSS.n852 VSS.t2460 1.1255
R8934 VSS.n853 VSS.t2436 1.1255
R8935 VSS.n702 VSS.t3800 1.1255
R8936 VSS.n703 VSS.t3807 1.1255
R8937 VSS.n704 VSS.t3648 1.1255
R8938 VSS.n705 VSS.t3609 1.1255
R8939 VSS.n706 VSS.t3678 1.1255
R8940 VSS.n707 VSS.t3740 1.1255
R8941 VSS.n708 VSS.t3611 1.1255
R8942 VSS.n709 VSS.t3618 1.1255
R8943 VSS.n710 VSS.t3640 1.1255
R8944 VSS.n711 VSS.t3574 1.1255
R8945 VSS.n712 VSS.t3804 1.1255
R8946 VSS.n713 VSS.t3745 1.1255
R8947 VSS.n714 VSS.t3783 1.1255
R8948 VSS.n715 VSS.t3730 1.1255
R8949 VSS.n716 VSS.t3766 1.1255
R8950 VSS.n717 VSS.t3657 1.1255
R8951 VSS.n718 VSS.t3656 1.1255
R8952 VSS.n719 VSS.t3560 1.1255
R8953 VSS.n720 VSS.t3590 1.1255
R8954 VSS.n721 VSS.t3732 1.1255
R8955 VSS.n722 VSS.t3639 1.1255
R8956 VSS.n723 VSS.t3764 1.1255
R8957 VSS.n724 VSS.t3775 1.1255
R8958 VSS.n725 VSS.t3716 1.1255
R8959 VSS.n726 VSS.t3550 1.1255
R8960 VSS.n727 VSS.t3675 1.1255
R8961 VSS.n728 VSS.t3565 1.1255
R8962 VSS.n729 VSS.t3741 1.1255
R8963 VSS.n730 VSS.t3555 1.1255
R8964 VSS.n731 VSS.t3696 1.1255
R8965 VSS.n732 VSS.t3776 1.1255
R8966 VSS.n733 VSS.t3801 1.1255
R8967 VSS.n734 VSS.t3608 1.1255
R8968 VSS.n735 VSS.t3646 1.1255
R8969 VSS.n736 VSS.t3638 1.1255
R8970 VSS.n737 VSS.t3724 1.1255
R8971 VSS.n738 VSS.t3802 1.1255
R8972 VSS.n739 VSS.t3815 1.1255
R8973 VSS.n740 VSS.t3674 1.1255
R8974 VSS.n741 VSS.t3559 1.1255
R8975 VSS.n742 VSS.t3575 1.1255
R8976 VSS.n743 VSS.t3779 1.1255
R8977 VSS.n744 VSS.t3587 1.1255
R8978 VSS.n745 VSS.t3803 1.1255
R8979 VSS.n746 VSS.t3605 1.1255
R8980 VSS.n747 VSS.t3715 1.1255
R8981 VSS.n748 VSS.t3628 1.1255
R8982 VSS.n749 VSS.t3772 1.1255
R8983 VSS.n750 VSS.t3582 1.1255
R8984 VSS.n751 VSS.t3669 1.1255
R8985 VSS.n752 VSS.t3765 1.1255
R8986 VSS.n753 VSS.t3558 1.1255
R8987 VSS.n754 VSS.t3672 1.1255
R8988 VSS.n755 VSS.t3557 1.1255
R8989 VSS.n756 VSS.t3697 1.1255
R8990 VSS.n757 VSS.t3679 1.1255
R8991 VSS.n758 VSS.t3761 1.1255
R8992 VSS.n759 VSS.t3643 1.1255
R8993 VSS.n760 VSS.t3720 1.1255
R8994 VSS.n761 VSS.t3601 1.1255
R8995 VSS.n762 VSS.t3694 1.1255
R8996 VSS.n763 VSS.t3681 1.1255
R8997 VSS.n764 VSS.t3794 1.1255
R8998 VSS.n765 VSS.t3650 1.1255
R8999 VSS.n766 VSS.t2327 1.1255
R9000 VSS.n3866 VSS.n3865 1.11354
R9001 VSS.n4669 VSS.n325 1.06209
R9002 VSS.n312 VSS.n311 1.04229
R9003 VSS.n2747 VSS.n2746 1.02178
R9004 VSS.n1147 VSS.n1141 1.01637
R9005 VSS.n947 VSS.n946 1.01637
R9006 VSS.n2890 VSS.n2889 1.00931
R9007 VSS.n1136 VSS.n915 0.973907
R9008 VSS.n5751 VSS.n16 0.952566
R9009 VSS.n5706 VSS.n34 0.952566
R9010 VSS.n5687 VSS.n44 0.952566
R9011 VSS.n97 VSS.n96 0.952566
R9012 VSS.n142 VSS.n141 0.952566
R9013 VSS.n3128 VSS.n3127 0.952566
R9014 VSS.n1869 VSS.n1423 0.952566
R9015 VSS.n290 VSS.n289 0.952566
R9016 VSS.n282 VSS.n281 0.952566
R9017 VSS.n5054 VSS.n267 0.952566
R9018 VSS.n261 VSS.n260 0.952566
R9019 VSS.n5158 VSS.n5132 0.952566
R9020 VSS.n5145 VSS.n5144 0.952566
R9021 VSS.n960 VSS.n959 0.951114
R9022 VSS.n634 VSS.n633 0.914923
R9023 VSS.n771 VSS.n769 0.914923
R9024 VSS.n2464 VSS.n2463 0.89958
R9025 VSS.n4598 VSS.n4592 0.883259
R9026 VSS.n987 VSS.n979 0.883259
R9027 VSS.n4762 VSS.n4761 0.881168
R9028 VSS.n528 VSS.n527 0.881168
R9029 VSS.n3612 VSS.n3611 0.877212
R9030 VSS.n3892 VSS.n3891 0.853833
R9031 VSS.n4607 VSS.n4606 0.848387
R9032 VSS.n984 VSS.n980 0.848386
R9033 VSS.n1697 VSS.n1696 0.835283
R9034 VSS.n5666 VSS.n5665 0.833377
R9035 VSS.n5483 VSS.n5482 0.833377
R9036 VSS.n3937 VSS.n3936 0.833377
R9037 VSS.n4084 VSS.n4083 0.833377
R9038 VSS.n3608 VSS.n3607 0.833377
R9039 VSS.n3357 VSS.n3075 0.833377
R9040 VSS.n3362 VSS.n3361 0.833377
R9041 VSS.n3301 VSS.n3300 0.833377
R9042 VSS.n2639 VSS.n2638 0.833377
R9043 VSS.n1917 VSS.n1397 0.833377
R9044 VSS.n340 VSS.n339 0.811095
R9045 VSS.n4730 VSS.n4729 0.769731
R9046 VSS.n4731 VSS.n4730 0.769731
R9047 VSS.n4732 VSS.n4731 0.769731
R9048 VSS.n4733 VSS.n4732 0.769731
R9049 VSS.n4734 VSS.n4733 0.769731
R9050 VSS.n4735 VSS.n4734 0.769731
R9051 VSS.n4736 VSS.n4735 0.769731
R9052 VSS.n4737 VSS.n4736 0.769731
R9053 VSS.n4738 VSS.n4737 0.769731
R9054 VSS.n4739 VSS.n4738 0.769731
R9055 VSS.n4740 VSS.n4739 0.769731
R9056 VSS.n4741 VSS.n4740 0.769731
R9057 VSS.n4742 VSS.n4741 0.769731
R9058 VSS.n4743 VSS.n4742 0.769731
R9059 VSS.n4744 VSS.n4743 0.769731
R9060 VSS.n4694 VSS.n4693 0.769731
R9061 VSS.n4693 VSS.n4692 0.769731
R9062 VSS.n4692 VSS.n4691 0.769731
R9063 VSS.n4691 VSS.n4690 0.769731
R9064 VSS.n4690 VSS.n4689 0.769731
R9065 VSS.n4689 VSS.n4688 0.769731
R9066 VSS.n4688 VSS.n4687 0.769731
R9067 VSS.n4687 VSS.n4686 0.769731
R9068 VSS.n4686 VSS.n4685 0.769731
R9069 VSS.n4685 VSS.n4684 0.769731
R9070 VSS.n4684 VSS.n4683 0.769731
R9071 VSS.n4683 VSS.n4682 0.769731
R9072 VSS.n4682 VSS.n4681 0.769731
R9073 VSS.n4681 VSS.n4680 0.769731
R9074 VSS.n4680 VSS.n4679 0.769731
R9075 VSS.n618 VSS.n547 0.769731
R9076 VSS.n619 VSS.n618 0.769731
R9077 VSS.n620 VSS.n619 0.769731
R9078 VSS.n621 VSS.n620 0.769731
R9079 VSS.n622 VSS.n621 0.769731
R9080 VSS.n623 VSS.n622 0.769731
R9081 VSS.n624 VSS.n623 0.769731
R9082 VSS.n625 VSS.n624 0.769731
R9083 VSS.n626 VSS.n625 0.769731
R9084 VSS.n627 VSS.n626 0.769731
R9085 VSS.n628 VSS.n627 0.769731
R9086 VSS.n629 VSS.n628 0.769731
R9087 VSS.n630 VSS.n629 0.769731
R9088 VSS.n631 VSS.n630 0.769731
R9089 VSS.n632 VSS.n631 0.769731
R9090 VSS.n633 VSS.n632 0.769731
R9091 VSS.n4761 VSS.n4760 0.769731
R9092 VSS.n4760 VSS.n4759 0.769731
R9093 VSS.n4759 VSS.n4758 0.769731
R9094 VSS.n4758 VSS.n4757 0.769731
R9095 VSS.n4757 VSS.n4756 0.769731
R9096 VSS.n4756 VSS.n4755 0.769731
R9097 VSS.n4755 VSS.n4754 0.769731
R9098 VSS.n4754 VSS.n4753 0.769731
R9099 VSS.n4753 VSS.n4752 0.769731
R9100 VSS.n4752 VSS.n4751 0.769731
R9101 VSS.n4751 VSS.n4750 0.769731
R9102 VSS.n4750 VSS.n4749 0.769731
R9103 VSS.n4749 VSS.n4748 0.769731
R9104 VSS.n4748 VSS.n4747 0.769731
R9105 VSS.n4747 VSS.n4746 0.769731
R9106 VSS.n892 VSS.n891 0.769731
R9107 VSS.n893 VSS.n892 0.769731
R9108 VSS.n894 VSS.n893 0.769731
R9109 VSS.n895 VSS.n894 0.769731
R9110 VSS.n896 VSS.n895 0.769731
R9111 VSS.n897 VSS.n896 0.769731
R9112 VSS.n898 VSS.n897 0.769731
R9113 VSS.n899 VSS.n898 0.769731
R9114 VSS.n900 VSS.n899 0.769731
R9115 VSS.n901 VSS.n900 0.769731
R9116 VSS.n902 VSS.n901 0.769731
R9117 VSS.n903 VSS.n902 0.769731
R9118 VSS.n904 VSS.n903 0.769731
R9119 VSS.n905 VSS.n904 0.769731
R9120 VSS.n906 VSS.n905 0.769731
R9121 VSS.n787 VSS.n786 0.769731
R9122 VSS.n786 VSS.n785 0.769731
R9123 VSS.n785 VSS.n784 0.769731
R9124 VSS.n784 VSS.n783 0.769731
R9125 VSS.n783 VSS.n782 0.769731
R9126 VSS.n782 VSS.n781 0.769731
R9127 VSS.n781 VSS.n780 0.769731
R9128 VSS.n780 VSS.n779 0.769731
R9129 VSS.n779 VSS.n778 0.769731
R9130 VSS.n778 VSS.n777 0.769731
R9131 VSS.n777 VSS.n776 0.769731
R9132 VSS.n776 VSS.n775 0.769731
R9133 VSS.n775 VSS.n774 0.769731
R9134 VSS.n774 VSS.n773 0.769731
R9135 VSS.n773 VSS.n772 0.769731
R9136 VSS.n772 VSS.n771 0.769731
R9137 VSS.n480 VSS.n479 0.769731
R9138 VSS.n481 VSS.n480 0.769731
R9139 VSS.n482 VSS.n481 0.769731
R9140 VSS.n483 VSS.n482 0.769731
R9141 VSS.n484 VSS.n483 0.769731
R9142 VSS.n485 VSS.n484 0.769731
R9143 VSS.n486 VSS.n485 0.769731
R9144 VSS.n487 VSS.n486 0.769731
R9145 VSS.n488 VSS.n487 0.769731
R9146 VSS.n489 VSS.n488 0.769731
R9147 VSS.n490 VSS.n489 0.769731
R9148 VSS.n491 VSS.n490 0.769731
R9149 VSS.n492 VSS.n491 0.769731
R9150 VSS.n493 VSS.n492 0.769731
R9151 VSS.n494 VSS.n493 0.769731
R9152 VSS.n543 VSS.n542 0.769731
R9153 VSS.n542 VSS.n541 0.769731
R9154 VSS.n541 VSS.n540 0.769731
R9155 VSS.n540 VSS.n539 0.769731
R9156 VSS.n539 VSS.n538 0.769731
R9157 VSS.n538 VSS.n537 0.769731
R9158 VSS.n537 VSS.n536 0.769731
R9159 VSS.n536 VSS.n535 0.769731
R9160 VSS.n535 VSS.n534 0.769731
R9161 VSS.n534 VSS.n533 0.769731
R9162 VSS.n533 VSS.n532 0.769731
R9163 VSS.n532 VSS.n531 0.769731
R9164 VSS.n531 VSS.n530 0.769731
R9165 VSS.n530 VSS.n529 0.769731
R9166 VSS.n529 VSS.n528 0.769731
R9167 VSS.n4670 VSS.n4669 0.765396
R9168 VSS.n4852 VSS.n325 0.7619
R9169 VSS.n4004 VSS.n3806 0.753441
R9170 VSS.n4099 VSS.n4098 0.753441
R9171 VSS.n4304 VSS.n4303 0.753441
R9172 VSS.n4366 VSS.n4365 0.753441
R9173 VSS.n3580 VSS.n3579 0.753441
R9174 VSS.n3508 VSS.n3008 0.753441
R9175 VSS.n3509 VSS.n3508 0.753441
R9176 VSS.n3487 VSS.n3486 0.753441
R9177 VSS.n3431 VSS.n3040 0.753441
R9178 VSS.n3384 VSS.n3383 0.753441
R9179 VSS.n3151 VSS.n3150 0.753441
R9180 VSS.n2623 VSS.n2622 0.753441
R9181 VSS.n2473 VSS.n2278 0.753441
R9182 VSS.n2358 VSS.n2357 0.753441
R9183 VSS.n2350 VSS.n2349 0.753441
R9184 VSS.n2697 VSS.n2696 0.753441
R9185 VSS.n2790 VSS.n2789 0.753441
R9186 VSS.n2825 VSS.n2824 0.753441
R9187 VSS.n2014 VSS.n2013 0.753441
R9188 VSS.n1999 VSS.n1998 0.753441
R9189 VSS.n1973 VSS.n1972 0.753441
R9190 VSS.n1851 VSS.n1850 0.753441
R9191 VSS.n1811 VSS.n1810 0.753441
R9192 VSS.n1745 VSS.n1486 0.753441
R9193 VSS.n1579 VSS.n1552 0.753441
R9194 VSS.n1570 VSS.n1569 0.753441
R9195 VSS.n1296 VSS.n1295 0.753441
R9196 VSS.n4858 VSS.n4857 0.753441
R9197 VSS.n4977 VSS.n4976 0.752461
R9198 VSS.n1168 VSS.n1166 0.750074
R9199 VSS.n2886 VSS.n2843 0.745706
R9200 VSS.n4328 VSS.n3723 0.743162
R9201 VSS.n473 VSS.n471 0.736693
R9202 VSS.n4695 VSS.n546 0.73175
R9203 VSS.n890 VSS.n856 0.73175
R9204 VSS.n1181 VSS.n1180 0.726407
R9205 VSS.n4641 VSS.n4640 0.726407
R9206 VSS.n4698 VSS.n4697 0.71758
R9207 VSS.n4699 VSS.n4698 0.71758
R9208 VSS.n4700 VSS.n4699 0.71758
R9209 VSS.n4701 VSS.n4700 0.71758
R9210 VSS.n4702 VSS.n4701 0.71758
R9211 VSS.n4703 VSS.n4702 0.71758
R9212 VSS.n4704 VSS.n4703 0.71758
R9213 VSS.n4705 VSS.n4704 0.71758
R9214 VSS.n4706 VSS.n4705 0.71758
R9215 VSS.n4707 VSS.n4706 0.71758
R9216 VSS.n4708 VSS.n4707 0.71758
R9217 VSS.n4709 VSS.n4708 0.71758
R9218 VSS.n4710 VSS.n4709 0.71758
R9219 VSS.n4711 VSS.n4710 0.71758
R9220 VSS.n4712 VSS.n4711 0.71758
R9221 VSS.n4713 VSS.n4712 0.71758
R9222 VSS.n4714 VSS.n4713 0.71758
R9223 VSS.n4715 VSS.n4714 0.71758
R9224 VSS.n4716 VSS.n4715 0.71758
R9225 VSS.n4717 VSS.n4716 0.71758
R9226 VSS.n4718 VSS.n4717 0.71758
R9227 VSS.n4719 VSS.n4718 0.71758
R9228 VSS.n4720 VSS.n4719 0.71758
R9229 VSS.n4721 VSS.n4720 0.71758
R9230 VSS.n4722 VSS.n4721 0.71758
R9231 VSS.n4723 VSS.n4722 0.71758
R9232 VSS.n4724 VSS.n4723 0.71758
R9233 VSS.n4725 VSS.n4724 0.71758
R9234 VSS.n4726 VSS.n4725 0.71758
R9235 VSS.n4727 VSS.n4726 0.71758
R9236 VSS.n4728 VSS.n4727 0.71758
R9237 VSS.n4794 VSS.n4793 0.71758
R9238 VSS.n4793 VSS.n4792 0.71758
R9239 VSS.n4792 VSS.n4791 0.71758
R9240 VSS.n4791 VSS.n4790 0.71758
R9241 VSS.n4790 VSS.n4789 0.71758
R9242 VSS.n4789 VSS.n4788 0.71758
R9243 VSS.n4788 VSS.n4787 0.71758
R9244 VSS.n4787 VSS.n4786 0.71758
R9245 VSS.n4786 VSS.n4785 0.71758
R9246 VSS.n4785 VSS.n4784 0.71758
R9247 VSS.n4784 VSS.n4783 0.71758
R9248 VSS.n4783 VSS.n4782 0.71758
R9249 VSS.n4782 VSS.n4781 0.71758
R9250 VSS.n4781 VSS.n4780 0.71758
R9251 VSS.n4780 VSS.n4779 0.71758
R9252 VSS.n4779 VSS.n4778 0.71758
R9253 VSS.n4778 VSS.n4777 0.71758
R9254 VSS.n4777 VSS.n4776 0.71758
R9255 VSS.n4776 VSS.n4775 0.71758
R9256 VSS.n4775 VSS.n4774 0.71758
R9257 VSS.n4774 VSS.n4773 0.71758
R9258 VSS.n4773 VSS.n4772 0.71758
R9259 VSS.n4772 VSS.n4771 0.71758
R9260 VSS.n4771 VSS.n4770 0.71758
R9261 VSS.n4770 VSS.n4769 0.71758
R9262 VSS.n4769 VSS.n4768 0.71758
R9263 VSS.n4768 VSS.n4767 0.71758
R9264 VSS.n4767 VSS.n4766 0.71758
R9265 VSS.n4766 VSS.n4765 0.71758
R9266 VSS.n4765 VSS.n4764 0.71758
R9267 VSS.n4764 VSS.n4763 0.71758
R9268 VSS.n888 VSS.n887 0.71758
R9269 VSS.n887 VSS.n886 0.71758
R9270 VSS.n886 VSS.n885 0.71758
R9271 VSS.n885 VSS.n884 0.71758
R9272 VSS.n884 VSS.n883 0.71758
R9273 VSS.n883 VSS.n882 0.71758
R9274 VSS.n882 VSS.n881 0.71758
R9275 VSS.n881 VSS.n880 0.71758
R9276 VSS.n880 VSS.n879 0.71758
R9277 VSS.n879 VSS.n878 0.71758
R9278 VSS.n878 VSS.n877 0.71758
R9279 VSS.n877 VSS.n876 0.71758
R9280 VSS.n876 VSS.n875 0.71758
R9281 VSS.n875 VSS.n874 0.71758
R9282 VSS.n874 VSS.n873 0.71758
R9283 VSS.n873 VSS.n872 0.71758
R9284 VSS.n872 VSS.n871 0.71758
R9285 VSS.n871 VSS.n870 0.71758
R9286 VSS.n870 VSS.n869 0.71758
R9287 VSS.n869 VSS.n868 0.71758
R9288 VSS.n868 VSS.n867 0.71758
R9289 VSS.n867 VSS.n866 0.71758
R9290 VSS.n866 VSS.n865 0.71758
R9291 VSS.n865 VSS.n864 0.71758
R9292 VSS.n864 VSS.n863 0.71758
R9293 VSS.n863 VSS.n862 0.71758
R9294 VSS.n862 VSS.n861 0.71758
R9295 VSS.n861 VSS.n860 0.71758
R9296 VSS.n860 VSS.n859 0.71758
R9297 VSS.n859 VSS.n858 0.71758
R9298 VSS.n858 VSS.n857 0.71758
R9299 VSS.n526 VSS.n525 0.71758
R9300 VSS.n525 VSS.n524 0.71758
R9301 VSS.n524 VSS.n523 0.71758
R9302 VSS.n523 VSS.n522 0.71758
R9303 VSS.n522 VSS.n521 0.71758
R9304 VSS.n521 VSS.n520 0.71758
R9305 VSS.n520 VSS.n519 0.71758
R9306 VSS.n519 VSS.n518 0.71758
R9307 VSS.n518 VSS.n517 0.71758
R9308 VSS.n517 VSS.n516 0.71758
R9309 VSS.n516 VSS.n515 0.71758
R9310 VSS.n515 VSS.n514 0.71758
R9311 VSS.n514 VSS.n513 0.71758
R9312 VSS.n513 VSS.n512 0.71758
R9313 VSS.n512 VSS.n511 0.71758
R9314 VSS.n511 VSS.n510 0.71758
R9315 VSS.n510 VSS.n509 0.71758
R9316 VSS.n509 VSS.n508 0.71758
R9317 VSS.n508 VSS.n507 0.71758
R9318 VSS.n507 VSS.n506 0.71758
R9319 VSS.n506 VSS.n505 0.71758
R9320 VSS.n505 VSS.n504 0.71758
R9321 VSS.n504 VSS.n503 0.71758
R9322 VSS.n503 VSS.n502 0.71758
R9323 VSS.n502 VSS.n501 0.71758
R9324 VSS.n501 VSS.n500 0.71758
R9325 VSS.n500 VSS.n499 0.71758
R9326 VSS.n499 VSS.n498 0.71758
R9327 VSS.n498 VSS.n497 0.71758
R9328 VSS.n497 VSS.n496 0.71758
R9329 VSS.n496 VSS.n495 0.71758
R9330 VSS.n3951 VSS.n3816 0.711611
R9331 VSS.n4027 VSS.n4026 0.711611
R9332 VSS.n3574 VSS.n3573 0.711611
R9333 VSS.n1645 VSS.n1642 0.711611
R9334 VSS.n470 VSS.n468 0.6935
R9335 VSS.n1176 VSS.n1160 0.6935
R9336 VSS.n2558 VSS.n2230 0.69032
R9337 VSS.n4257 VSS.n3754 0.681351
R9338 VSS.n4746 VSS.n4745 0.673577
R9339 VSS.n544 VSS.n543 0.673577
R9340 VSS.n4697 VSS.n4696 0.664161
R9341 VSS.n889 VSS.n888 0.664161
R9342 VSS.n527 VSS.n526 0.664161
R9343 VSS.n4763 VSS.n4762 0.664161
R9344 VSS.n1180 VSS.n1158 0.660581
R9345 VSS.n4640 VSS.n4635 0.660581
R9346 VSS.n4638 VSS.n4637 0.627947
R9347 VSS.n1177 VSS.n1159 0.627947
R9348 VSS.n4465 VSS.n4434 0.627073
R9349 VSS.n2576 VSS.n2575 0.627073
R9350 VSS.n2761 VSS.n2760 0.627073
R9351 VSS.n4079 VSS.n4078 0.613266
R9352 VSS.n4107 VSS.n4106 0.613266
R9353 VSS.n3465 VSS.n3464 0.613266
R9354 VSS.n2458 VSS.n2457 0.613266
R9355 VSS.n4637 VSS.n467 0.598603
R9356 VSS.n1161 VSS.n1159 0.598603
R9357 VSS.n4808 VSS.n468 0.596535
R9358 VSS.n1163 VSS.n1160 0.596535
R9359 VSS.n1116 VSS.n1115 0.563
R9360 VSS.n1117 VSS.n1116 0.563
R9361 VSS.n1118 VSS.n1117 0.563
R9362 VSS.n1120 VSS.n1118 0.563
R9363 VSS.n1029 VSS.n1028 0.563
R9364 VSS.n1030 VSS.n1029 0.563
R9365 VSS.n918 VSS.n917 0.563
R9366 VSS.n919 VSS.n918 0.563
R9367 VSS.n920 VSS.n919 0.563
R9368 VSS.n922 VSS.n920 0.563
R9369 VSS.n4806 VSS.n4805 0.561264
R9370 VSS.n1175 VSS.n1165 0.561264
R9371 VSS.n936 VSS.n935 0.559662
R9372 VSS.n4679 VSS.n4678 0.553385
R9373 VSS.n907 VSS.n906 0.553385
R9374 VSS.n4810 VSS.n4809 0.547559
R9375 VSS.n1162 VSS.n1001 0.547559
R9376 VSS.n317 VSS.n316 0.543
R9377 VSS.n4564 VSS.n9 0.537563
R9378 VSS.n4583 VSS.n4558 0.537563
R9379 VSS.n5708 VSS.n32 0.537563
R9380 VSS.n5727 VSS.n5726 0.537563
R9381 VSS.n5620 VSS.n74 0.537563
R9382 VSS.n5639 VSS.n68 0.537563
R9383 VSS.n5530 VSS.n5529 0.537563
R9384 VSS.n5549 VSS.n5548 0.537563
R9385 VSS.n5435 VSS.n153 0.537563
R9386 VSS.n5451 VSS.n147 0.537563
R9387 VSS.n5398 VSS.n5397 0.537563
R9388 VSS.n5417 VSS.n5416 0.537563
R9389 VSS.n4320 VSS.n4319 0.537563
R9390 VSS.n4341 VSS.n4340 0.537563
R9391 VSS.n4461 VSS.n4460 0.537563
R9392 VSS.n2561 VSS.n2226 0.537563
R9393 VSS.n2586 VSS.n2583 0.537563
R9394 VSS.n2532 VSS.n2531 0.537563
R9395 VSS.n2433 VSS.n2303 0.537563
R9396 VSS.n2751 VSS.n2180 0.537563
R9397 VSS.n2926 VSS.n2155 0.537563
R9398 VSS.n1594 VSS.n1593 0.537563
R9399 VSS.n1303 VSS.n1302 0.537563
R9400 VSS.n1133 VSS.n1131 0.53175
R9401 VSS.n935 VSS.n933 0.53175
R9402 VSS.n5662 VSS.n55 0.526527
R9403 VSS.n5478 VSS.n133 0.526527
R9404 VSS.n4080 VSS.n3797 0.526527
R9405 VSS.n3603 VSS.n2964 0.526527
R9406 VSS.n3358 VSS.n3356 0.526527
R9407 VSS.n3296 VSS.n3295 0.526527
R9408 VSS.n1918 VSS.n1916 0.526527
R9409 VSS.n1921 VSS.n1399 0.526527
R9410 VSS.n4808 VSS.n4807 0.52524
R9411 VSS.n1164 VSS.n1163 0.523938
R9412 VSS.n4635 VSS.n467 0.510917
R9413 VSS.n1161 VSS.n1158 0.510917
R9414 VSS.n1121 VSS.n1120 0.507196
R9415 VSS.n923 VSS.n922 0.507196
R9416 VSS.n4695 VSS.n4694 0.505308
R9417 VSS.n891 VSS.n890 0.505308
R9418 VSS.n1125 VSS.n1123 0.5005
R9419 VSS.n1127 VSS.n1125 0.5005
R9420 VSS.n1129 VSS.n1127 0.5005
R9421 VSS.n1131 VSS.n1129 0.5005
R9422 VSS.n927 VSS.n925 0.5005
R9423 VSS.n929 VSS.n927 0.5005
R9424 VSS.n931 VSS.n929 0.5005
R9425 VSS.n933 VSS.n931 0.5005
R9426 VSS.n4605 VSS.n937 0.5005
R9427 VSS.n1157 VSS.n985 0.5005
R9428 VSS.n4807 VSS.n4806 0.496683
R9429 VSS.n1165 VSS.n1164 0.496683
R9430 VSS.n3224 VSS.n3223 0.487457
R9431 VSS.n315 VSS.n314 0.4805
R9432 VSS.n3326 VSS.n3325 0.474574
R9433 VSS.n313 VSS.n312 0.472292
R9434 VSS.n4976 VSS.n4975 0.452653
R9435 VSS.n4978 VSS.n323 0.449932
R9436 VSS.n1135 VSS.n1133 0.444964
R9437 VSS.n4597 VSS.n4596 0.441879
R9438 VSS.n1215 VSS.n1214 0.441879
R9439 VSS.n3931 VSS.n3823 0.438856
R9440 VSS.n2642 VSS.n2194 0.438856
R9441 VSS.n4959 VSS.n362 0.438107
R9442 VSS.n4514 VSS.n4513 0.417891
R9443 VSS.n5739 VSS.n5738 0.417891
R9444 VSS.n5744 VSS.n20 0.417891
R9445 VSS.n5586 VSS.n5585 0.417891
R9446 VSS.n5590 VSS.n5589 0.417891
R9447 VSS.n5369 VSS.n5363 0.417891
R9448 VSS.n3861 VSS.n3846 0.417891
R9449 VSS.n3868 VSS.n3867 0.417891
R9450 VSS.n4296 VSS.n3735 0.417891
R9451 VSS.n4302 VSS.n4301 0.417891
R9452 VSS.n3584 VSS.n3583 0.417891
R9453 VSS.n3590 VSS.n3589 0.417891
R9454 VSS.n3409 VSS.n3055 0.417891
R9455 VSS.n3157 VSS.n3133 0.417891
R9456 VSS.n3221 VSS.n3220 0.417891
R9457 VSS.n2486 VSS.n2485 0.417891
R9458 VSS.n2491 VSS.n2270 0.417891
R9459 VSS.n2780 VSS.n2779 0.417891
R9460 VSS.n1993 VSS.n1992 0.417891
R9461 VSS.n1887 VSS.n1409 0.417891
R9462 VSS.n1894 VSS.n1893 0.417891
R9463 VSS.n1696 VSS.n1695 0.417891
R9464 VSS.n1702 VSS.n1503 0.417891
R9465 VSS.n1629 VSS.n1628 0.417891
R9466 VSS.n1630 VSS.n1530 0.417891
R9467 VSS.n4827 VSS.n390 0.417891
R9468 VSS.n4822 VSS.n4821 0.417891
R9469 VSS.n276 VSS.n273 0.417891
R9470 VSS.n5032 VSS.n5031 0.417891
R9471 VSS.n272 VSS.n270 0.417891
R9472 VSS.n5040 VSS.n5039 0.417891
R9473 VSS.n194 VSS.n192 0.417891
R9474 VSS.n5276 VSS.n5275 0.417891
R9475 VSS.n5294 VSS.n5293 0.417891
R9476 VSS.n5290 VSS.n5289 0.417891
R9477 VSS.n5335 VSS.n5334 0.417891
R9478 VSS.n419 VSS.n418 0.417891
R9479 VSS.n2127 VSS.n2126 0.416381
R9480 VSS.n5746 VSS.n17 0.409011
R9481 VSS.n5701 VSS.n5700 0.409011
R9482 VSS.n5682 VSS.n45 0.409011
R9483 VSS.n5656 VSS.n5655 0.409011
R9484 VSS.n5612 VSS.n5611 0.409011
R9485 VSS.n5619 VSS.n5618 0.409011
R9486 VSS.n5568 VSS.n5567 0.409011
R9487 VSS.n5556 VSS.n101 0.409011
R9488 VSS.n5563 VSS.n5562 0.409011
R9489 VSS.n5521 VSS.n5520 0.409011
R9490 VSS.n5528 VSS.n5527 0.409011
R9491 VSS.n5472 VSS.n5471 0.409011
R9492 VSS.n5463 VSS.n5462 0.409011
R9493 VSS.n5427 VSS.n5426 0.409011
R9494 VSS.n5434 VSS.n5433 0.409011
R9495 VSS.n3923 VSS.n3922 0.409011
R9496 VSS.n4043 VSS.n3983 0.409011
R9497 VSS.n4073 VSS.n4072 0.409011
R9498 VSS.n4105 VSS.n4104 0.409011
R9499 VSS.n4112 VSS.n3781 0.409011
R9500 VSS.n4173 VSS.n4171 0.409011
R9501 VSS.n4256 VSS.n4255 0.409011
R9502 VSS.n4266 VSS.n3750 0.409011
R9503 VSS.n4309 VSS.n3730 0.409011
R9504 VSS.n4316 VSS.n4315 0.409011
R9505 VSS.n3466 VSS.n3465 0.409011
R9506 VSS.n3473 VSS.n3472 0.409011
R9507 VSS.n3457 VSS.n3455 0.409011
R9508 VSS.n3389 VSS.n3062 0.409011
R9509 VSS.n3396 VSS.n3395 0.409011
R9510 VSS.n3350 VSS.n3349 0.409011
R9511 VSS.n3289 VSS.n3103 0.409011
R9512 VSS.n3272 VSS.n3113 0.409011
R9513 VSS.n2604 VSS.n2603 0.409011
R9514 VSS.n2607 VSS.n2208 0.409011
R9515 VSS.n2456 VSS.n2455 0.409011
R9516 VSS.n2463 VSS.n2284 0.409011
R9517 VSS.n2721 VSS.n2665 0.409011
R9518 VSS.n2707 VSS.n2706 0.409011
R9519 VSS.n2700 VSS.n2677 0.409011
R9520 VSS.n2742 VSS.n2741 0.409011
R9521 VSS.n2750 VSS.n2749 0.409011
R9522 VSS.n2059 VSS.n2058 0.409011
R9523 VSS.n2066 VSS.n1332 0.409011
R9524 VSS.n1909 VSS.n1908 0.409011
R9525 VSS.n1864 VSS.n1863 0.409011
R9526 VSS.n1674 VSS.n1673 0.409011
R9527 VSS.n1684 VSS.n1511 0.409011
R9528 VSS.n372 VSS.n370 0.409011
R9529 VSS.n4872 VSS.n4871 0.409011
R9530 VSS.n5011 VSS.n5010 0.409011
R9531 VSS.n5025 VSS.n5024 0.409011
R9532 VSS.n266 VSS.n264 0.409011
R9533 VSS.n5070 VSS.n5069 0.409011
R9534 VSS.n5119 VSS.n5118 0.409011
R9535 VSS.n5113 VSS.n240 0.409011
R9536 VSS.n5153 VSS.n5133 0.409011
R9537 VSS.n5142 VSS.n5141 0.409011
R9538 VSS.n5193 VSS.n5192 0.409011
R9539 VSS.n5187 VSS.n231 0.409011
R9540 VSS.n5206 VSS.n5205 0.409011
R9541 VSS.n5200 VSS.n224 0.409011
R9542 VSS.n5224 VSS.n5223 0.409011
R9543 VSS.n5218 VSS.n216 0.409011
R9544 VSS.n5242 VSS.n208 0.409011
R9545 VSS.n5236 VSS.n5235 0.409011
R9546 VSS.n460 VSS.n395 0.409011
R9547 VSS.n454 VSS.n453 0.409011
R9548 VSS.n4976 VSS.n325 0.406443
R9549 VSS.n3300 VSS.n3100 0.395021
R9550 VSS.n4978 VSS.n4977 0.393625
R9551 VSS.n1144 VSS.n1138 0.388
R9552 VSS.n1147 VSS.n1139 0.388
R9553 VSS.n946 VSS.n945 0.388
R9554 VSS.n4664 VSS.n4663 0.388
R9555 VSS.n4795 VSS.n4794 0.383079
R9556 VSS.n495 VSS.n477 0.383079
R9557 VSS.n4094 VSS.n3789 0.376971
R9558 VSS.n4214 VSS.n4213 0.376971
R9559 VSS.n3626 VSS.n2956 0.376971
R9560 VSS.n3623 VSS.n2956 0.376971
R9561 VSS.n3482 VSS.n3018 0.376971
R9562 VSS.n3271 VSS.n3270 0.376971
R9563 VSS.n2619 VSS.n2618 0.376971
R9564 VSS.n2550 VSS.n2549 0.376971
R9565 VSS.n2471 VSS.n2470 0.376971
R9566 VSS.n2009 VSS.n2008 0.376971
R9567 VSS.n1872 VSS.n1871 0.376971
R9568 VSS.n1856 VSS.n1430 0.376971
R9569 VSS.n1736 VSS.n1735 0.376971
R9570 VSS.n4845 VSS.n4837 0.376971
R9571 VSS.n1092 VSS.n1033 0.376971
R9572 VSS.n4639 VSS.n4636 0.371802
R9573 VSS.n1179 VSS.n1178 0.371802
R9574 VSS.n3161 VSS.n3159 0.358542
R9575 VSS.n3216 VSS.n3215 0.358542
R9576 VSS.n2115 VSS.n2073 0.358542
R9577 VSS.n2109 VSS.n2077 0.358542
R9578 VSS.n2103 VSS.n2080 0.358542
R9579 VSS.n1601 VSS.n1600 0.358542
R9580 VSS.n1312 VSS.n1311 0.358542
R9581 VSS.n1305 VSS.n1304 0.358542
R9582 VSS.n2231 VSS.n2227 0.357692
R9583 VSS.n3334 VSS.n3330 0.356056
R9584 VSS.n4638 VSS.n470 0.343032
R9585 VSS.n1177 VSS.n1176 0.343032
R9586 VSS.n3979 VSS.n3978 0.340926
R9587 VSS.n2715 VSS.n2714 0.340926
R9588 VSS.n4696 VSS.n4695 0.340303
R9589 VSS.n890 VSS.n889 0.340303
R9590 VSS.n1096 VSS.n1095 0.338974
R9591 VSS.n4809 VSS.n467 0.337621
R9592 VSS.n1162 VSS.n1161 0.337621
R9593 VSS.n4795 VSS.n4728 0.335002
R9594 VSS.n857 VSS.n477 0.335002
R9595 VSS.n4636 VSS.n4635 0.333523
R9596 VSS.n1178 VSS.n1158 0.333523
R9597 VSS.n317 VSS.n315 0.333
R9598 VSS.n4980 VSS.n317 0.330857
R9599 VSS.n4809 VSS.n4808 0.328202
R9600 VSS.n1163 VSS.n1162 0.328202
R9601 VSS.n4805 VSS.n470 0.32761
R9602 VSS.n1176 VSS.n1175 0.326799
R9603 VSS.n1155 VSS.n1138 0.326171
R9604 VSS.n4665 VSS.n4664 0.325788
R9605 VSS.n915 VSS.n324 0.324892
R9606 VSS.n4811 VSS.n4810 0.3205
R9607 VSS.n1200 VSS.n1001 0.3205
R9608 VSS.n4639 VSS.n4638 0.318682
R9609 VSS.n1179 VSS.n1177 0.318682
R9610 VSS.n333 VSS.n332 0.311532
R9611 VSS.n4974 VSS.n4973 0.3105
R9612 VSS.n3363 VSS.n3362 0.307349
R9613 VSS.n2637 VSS.n2636 0.307349
R9614 VSS.n3899 VSS.n3898 0.305262
R9615 VSS.n3916 VSS.n3830 0.305262
R9616 VSS.n4428 VSS.n4426 0.305262
R9617 VSS.n4468 VSS.n4431 0.305262
R9618 VSS.n3189 VSS.n3188 0.305262
R9619 VSS.n3176 VSS.n3175 0.305262
R9620 VSS.n3196 VSS.n3195 0.305262
R9621 VSS.n3190 VSS.n3171 0.305262
R9622 VSS.n3164 VSS.n3162 0.305262
R9623 VSS.n3198 VSS.n3167 0.305262
R9624 VSS.n2389 VSS.n2388 0.305262
R9625 VSS.n2400 VSS.n2314 0.305262
R9626 VSS.n3888 VSS.n3837 0.298074
R9627 VSS.n2128 VSS.n2127 0.298074
R9628 VSS.n2555 VSS.n2231 0.29768
R9629 VSS.n321 VSS.n320 0.297375
R9630 VSS.n3896 VSS.n3837 0.297291
R9631 VSS.n4977 VSS.n324 0.288701
R9632 VSS.n3403 VSS.n3057 0.278761
R9633 VSS.n3457 VSS.n3456 0.27331
R9634 VSS.n4222 VSS.n4221 0.27284
R9635 VSS.n3602 VSS.n3601 0.27284
R9636 VSS.n2368 VSS.n2367 0.27284
R9637 VSS.n2510 VSS.n2253 0.269031
R9638 VSS.n2511 VSS.n2510 0.269031
R9639 VSS.n347 VSS.n346 0.267759
R9640 VSS.n5670 VSS.n5669 0.263514
R9641 VSS.n5487 VSS.n5486 0.263514
R9642 VSS.n4088 VSS.n4087 0.263514
R9643 VSS.n3613 VSS.n3612 0.263514
R9644 VSS.n3076 VSS.n3073 0.263514
R9645 VSS.n3305 VSS.n3304 0.263514
R9646 VSS.n2195 VSS.n2191 0.263514
R9647 VSS.n1925 VSS.n1395 0.263514
R9648 VSS.n4327 VSS.n4326 0.262616
R9649 VSS.n4332 VSS.n3723 0.262616
R9650 VSS.n3884 VSS.n3883 0.259086
R9651 VSS.n4425 VSS.n4423 0.259086
R9652 VSS.n4483 VSS.n4482 0.259086
R9653 VSS.n3236 VSS.n3235 0.259086
R9654 VSS.n3239 VSS.n3238 0.259086
R9655 VSS.n1607 VSS.n1606 0.259086
R9656 VSS.n1325 VSS.n1324 0.259086
R9657 VSS.n1318 VSS.n1317 0.259086
R9658 VSS.n1612 VSS.n1537 0.240317
R9659 VSS.n2900 VSS.n2899 0.239726
R9660 VSS.n5467 VSS.n5466 0.239726
R9661 VSS.n5572 VSS.n5571 0.239726
R9662 VSS.n5689 VSS.n43 0.239726
R9663 VSS.n5704 VSS.n33 0.239726
R9664 VSS.n5753 VSS.n15 0.239726
R9665 VSS.n3880 VSS.n3879 0.239726
R9666 VSS.n2126 VSS.n2072 0.239726
R9667 VSS.n3241 VSS.n3240 0.239726
R9668 VSS.n2382 VSS.n2319 0.239726
R9669 VSS.n2626 VSS.n2200 0.239726
R9670 VSS.n1867 VSS.n1422 0.239726
R9671 VSS.n5148 VSS.n5147 0.239726
R9672 VSS.n5160 VSS.n5131 0.239726
R9673 VSS.n5066 VSS.n5065 0.239726
R9674 VSS.n5052 VSS.n265 0.239726
R9675 VSS.n5021 VSS.n5020 0.239726
R9676 VSS.n5007 VSS.n5006 0.239726
R9677 VSS.n5467 VSS.n137 0.239381
R9678 VSS.n5572 VSS.n94 0.239381
R9679 VSS.n5690 VSS.n5689 0.239381
R9680 VSS.n5709 VSS.n33 0.239381
R9681 VSS.n5754 VSS.n5753 0.239381
R9682 VSS.n3880 VSS.n3839 0.239381
R9683 VSS.n3241 VSS.n3126 0.239381
R9684 VSS.n2390 VSS.n2319 0.239381
R9685 VSS.n2633 VSS.n2200 0.239381
R9686 VSS.n2901 VSS.n2900 0.239381
R9687 VSS.n1873 VSS.n1422 0.239381
R9688 VSS.n5149 VSS.n5148 0.239381
R9689 VSS.n5161 VSS.n5160 0.239381
R9690 VSS.n5065 VSS.n5064 0.239381
R9691 VSS.n5052 VSS.n5051 0.239381
R9692 VSS.n5020 VSS.n5019 0.239381
R9693 VSS.n5006 VSS.n5005 0.239381
R9694 VSS.n2374 VSS.n2322 0.225061
R9695 VSS.n2383 VSS.n2320 0.225061
R9696 VSS.n2898 VSS.n2897 0.225061
R9697 VSS.n2891 VSS.n2890 0.225061
R9698 VSS.n2636 VSS.n2635 0.219678
R9699 VSS.n4678 VSS.n547 0.216846
R9700 VSS.n907 VSS.n787 0.216846
R9701 VSS.n4982 VSS.n4981 0.216779
R9702 VSS.n4669 VSS.n4668 0.213625
R9703 VSS.n1988 VSS.n1366 0.209196
R9704 VSS.n1989 VSS.n1988 0.209196
R9705 VSS.n3596 VSS.n3595 0.204755
R9706 VSS.n3595 VSS.n3592 0.204755
R9707 VSS.n3449 VSS.n3448 0.204755
R9708 VSS.n3448 VSS.n3034 0.204755
R9709 VSS.n2741 VSS.n2740 0.204755
R9710 VSS.n1164 VSS.n986 0.203625
R9711 VSS.n4807 VSS.n469 0.202323
R9712 VSS.n1095 VSS.n323 0.190841
R9713 VSS.n550 VSS.n549 0.180667
R9714 VSS.n551 VSS.n550 0.180667
R9715 VSS.n552 VSS.n551 0.180667
R9716 VSS.n553 VSS.n552 0.180667
R9717 VSS.n554 VSS.n553 0.180667
R9718 VSS.n555 VSS.n554 0.180667
R9719 VSS.n556 VSS.n555 0.180667
R9720 VSS.n557 VSS.n556 0.180667
R9721 VSS.n558 VSS.n557 0.180667
R9722 VSS.n559 VSS.n558 0.180667
R9723 VSS.n560 VSS.n559 0.180667
R9724 VSS.n561 VSS.n560 0.180667
R9725 VSS.n562 VSS.n561 0.180667
R9726 VSS.n563 VSS.n562 0.180667
R9727 VSS.n564 VSS.n563 0.180667
R9728 VSS.n565 VSS.n564 0.180667
R9729 VSS.n566 VSS.n565 0.180667
R9730 VSS.n567 VSS.n566 0.180667
R9731 VSS.n568 VSS.n567 0.180667
R9732 VSS.n569 VSS.n568 0.180667
R9733 VSS.n570 VSS.n569 0.180667
R9734 VSS.n571 VSS.n570 0.180667
R9735 VSS.n572 VSS.n571 0.180667
R9736 VSS.n573 VSS.n572 0.180667
R9737 VSS.n574 VSS.n573 0.180667
R9738 VSS.n575 VSS.n574 0.180667
R9739 VSS.n576 VSS.n575 0.180667
R9740 VSS.n577 VSS.n576 0.180667
R9741 VSS.n578 VSS.n577 0.180667
R9742 VSS.n579 VSS.n578 0.180667
R9743 VSS.n580 VSS.n579 0.180667
R9744 VSS.n581 VSS.n580 0.180667
R9745 VSS.n582 VSS.n581 0.180667
R9746 VSS.n583 VSS.n582 0.180667
R9747 VSS.n584 VSS.n583 0.180667
R9748 VSS.n585 VSS.n584 0.180667
R9749 VSS.n586 VSS.n585 0.180667
R9750 VSS.n587 VSS.n586 0.180667
R9751 VSS.n588 VSS.n587 0.180667
R9752 VSS.n589 VSS.n588 0.180667
R9753 VSS.n590 VSS.n589 0.180667
R9754 VSS.n591 VSS.n590 0.180667
R9755 VSS.n592 VSS.n591 0.180667
R9756 VSS.n593 VSS.n592 0.180667
R9757 VSS.n594 VSS.n593 0.180667
R9758 VSS.n595 VSS.n594 0.180667
R9759 VSS.n596 VSS.n595 0.180667
R9760 VSS.n597 VSS.n596 0.180667
R9761 VSS.n598 VSS.n597 0.180667
R9762 VSS.n599 VSS.n598 0.180667
R9763 VSS.n600 VSS.n599 0.180667
R9764 VSS.n601 VSS.n600 0.180667
R9765 VSS.n602 VSS.n601 0.180667
R9766 VSS.n603 VSS.n602 0.180667
R9767 VSS.n604 VSS.n603 0.180667
R9768 VSS.n605 VSS.n604 0.180667
R9769 VSS.n606 VSS.n605 0.180667
R9770 VSS.n607 VSS.n606 0.180667
R9771 VSS.n608 VSS.n607 0.180667
R9772 VSS.n609 VSS.n608 0.180667
R9773 VSS.n610 VSS.n609 0.180667
R9774 VSS.n611 VSS.n610 0.180667
R9775 VSS.n612 VSS.n611 0.180667
R9776 VSS.n613 VSS.n612 0.180667
R9777 VSS.n637 VSS.n636 0.180667
R9778 VSS.n638 VSS.n637 0.180667
R9779 VSS.n639 VSS.n638 0.180667
R9780 VSS.n640 VSS.n639 0.180667
R9781 VSS.n641 VSS.n640 0.180667
R9782 VSS.n642 VSS.n641 0.180667
R9783 VSS.n643 VSS.n642 0.180667
R9784 VSS.n644 VSS.n643 0.180667
R9785 VSS.n645 VSS.n644 0.180667
R9786 VSS.n646 VSS.n645 0.180667
R9787 VSS.n647 VSS.n646 0.180667
R9788 VSS.n648 VSS.n647 0.180667
R9789 VSS.n649 VSS.n648 0.180667
R9790 VSS.n650 VSS.n649 0.180667
R9791 VSS.n651 VSS.n650 0.180667
R9792 VSS.n652 VSS.n651 0.180667
R9793 VSS.n653 VSS.n652 0.180667
R9794 VSS.n654 VSS.n653 0.180667
R9795 VSS.n655 VSS.n654 0.180667
R9796 VSS.n656 VSS.n655 0.180667
R9797 VSS.n657 VSS.n656 0.180667
R9798 VSS.n658 VSS.n657 0.180667
R9799 VSS.n659 VSS.n658 0.180667
R9800 VSS.n660 VSS.n659 0.180667
R9801 VSS.n661 VSS.n660 0.180667
R9802 VSS.n662 VSS.n661 0.180667
R9803 VSS.n663 VSS.n662 0.180667
R9804 VSS.n664 VSS.n663 0.180667
R9805 VSS.n665 VSS.n664 0.180667
R9806 VSS.n666 VSS.n665 0.180667
R9807 VSS.n667 VSS.n666 0.180667
R9808 VSS.n668 VSS.n667 0.180667
R9809 VSS.n669 VSS.n668 0.180667
R9810 VSS.n670 VSS.n669 0.180667
R9811 VSS.n671 VSS.n670 0.180667
R9812 VSS.n672 VSS.n671 0.180667
R9813 VSS.n673 VSS.n672 0.180667
R9814 VSS.n674 VSS.n673 0.180667
R9815 VSS.n675 VSS.n674 0.180667
R9816 VSS.n676 VSS.n675 0.180667
R9817 VSS.n677 VSS.n676 0.180667
R9818 VSS.n678 VSS.n677 0.180667
R9819 VSS.n679 VSS.n678 0.180667
R9820 VSS.n680 VSS.n679 0.180667
R9821 VSS.n681 VSS.n680 0.180667
R9822 VSS.n682 VSS.n681 0.180667
R9823 VSS.n683 VSS.n682 0.180667
R9824 VSS.n684 VSS.n683 0.180667
R9825 VSS.n685 VSS.n684 0.180667
R9826 VSS.n686 VSS.n685 0.180667
R9827 VSS.n687 VSS.n686 0.180667
R9828 VSS.n688 VSS.n687 0.180667
R9829 VSS.n689 VSS.n688 0.180667
R9830 VSS.n690 VSS.n689 0.180667
R9831 VSS.n691 VSS.n690 0.180667
R9832 VSS.n692 VSS.n691 0.180667
R9833 VSS.n693 VSS.n692 0.180667
R9834 VSS.n694 VSS.n693 0.180667
R9835 VSS.n695 VSS.n694 0.180667
R9836 VSS.n696 VSS.n695 0.180667
R9837 VSS.n697 VSS.n696 0.180667
R9838 VSS.n698 VSS.n697 0.180667
R9839 VSS.n699 VSS.n698 0.180667
R9840 VSS.n700 VSS.n699 0.180667
R9841 VSS.n790 VSS.n789 0.180667
R9842 VSS.n791 VSS.n790 0.180667
R9843 VSS.n792 VSS.n791 0.180667
R9844 VSS.n793 VSS.n792 0.180667
R9845 VSS.n794 VSS.n793 0.180667
R9846 VSS.n795 VSS.n794 0.180667
R9847 VSS.n796 VSS.n795 0.180667
R9848 VSS.n797 VSS.n796 0.180667
R9849 VSS.n798 VSS.n797 0.180667
R9850 VSS.n799 VSS.n798 0.180667
R9851 VSS.n800 VSS.n799 0.180667
R9852 VSS.n801 VSS.n800 0.180667
R9853 VSS.n802 VSS.n801 0.180667
R9854 VSS.n803 VSS.n802 0.180667
R9855 VSS.n804 VSS.n803 0.180667
R9856 VSS.n805 VSS.n804 0.180667
R9857 VSS.n806 VSS.n805 0.180667
R9858 VSS.n807 VSS.n806 0.180667
R9859 VSS.n808 VSS.n807 0.180667
R9860 VSS.n809 VSS.n808 0.180667
R9861 VSS.n810 VSS.n809 0.180667
R9862 VSS.n811 VSS.n810 0.180667
R9863 VSS.n812 VSS.n811 0.180667
R9864 VSS.n813 VSS.n812 0.180667
R9865 VSS.n814 VSS.n813 0.180667
R9866 VSS.n815 VSS.n814 0.180667
R9867 VSS.n816 VSS.n815 0.180667
R9868 VSS.n817 VSS.n816 0.180667
R9869 VSS.n818 VSS.n817 0.180667
R9870 VSS.n819 VSS.n818 0.180667
R9871 VSS.n820 VSS.n819 0.180667
R9872 VSS.n821 VSS.n820 0.180667
R9873 VSS.n822 VSS.n821 0.180667
R9874 VSS.n823 VSS.n822 0.180667
R9875 VSS.n824 VSS.n823 0.180667
R9876 VSS.n825 VSS.n824 0.180667
R9877 VSS.n826 VSS.n825 0.180667
R9878 VSS.n827 VSS.n826 0.180667
R9879 VSS.n828 VSS.n827 0.180667
R9880 VSS.n829 VSS.n828 0.180667
R9881 VSS.n830 VSS.n829 0.180667
R9882 VSS.n831 VSS.n830 0.180667
R9883 VSS.n832 VSS.n831 0.180667
R9884 VSS.n833 VSS.n832 0.180667
R9885 VSS.n834 VSS.n833 0.180667
R9886 VSS.n835 VSS.n834 0.180667
R9887 VSS.n836 VSS.n835 0.180667
R9888 VSS.n837 VSS.n836 0.180667
R9889 VSS.n838 VSS.n837 0.180667
R9890 VSS.n839 VSS.n838 0.180667
R9891 VSS.n840 VSS.n839 0.180667
R9892 VSS.n841 VSS.n840 0.180667
R9893 VSS.n842 VSS.n841 0.180667
R9894 VSS.n843 VSS.n842 0.180667
R9895 VSS.n844 VSS.n843 0.180667
R9896 VSS.n845 VSS.n844 0.180667
R9897 VSS.n846 VSS.n845 0.180667
R9898 VSS.n847 VSS.n846 0.180667
R9899 VSS.n848 VSS.n847 0.180667
R9900 VSS.n849 VSS.n848 0.180667
R9901 VSS.n850 VSS.n849 0.180667
R9902 VSS.n851 VSS.n850 0.180667
R9903 VSS.n852 VSS.n851 0.180667
R9904 VSS.n853 VSS.n852 0.180667
R9905 VSS.n703 VSS.n702 0.180667
R9906 VSS.n704 VSS.n703 0.180667
R9907 VSS.n705 VSS.n704 0.180667
R9908 VSS.n706 VSS.n705 0.180667
R9909 VSS.n707 VSS.n706 0.180667
R9910 VSS.n708 VSS.n707 0.180667
R9911 VSS.n709 VSS.n708 0.180667
R9912 VSS.n710 VSS.n709 0.180667
R9913 VSS.n711 VSS.n710 0.180667
R9914 VSS.n712 VSS.n711 0.180667
R9915 VSS.n713 VSS.n712 0.180667
R9916 VSS.n714 VSS.n713 0.180667
R9917 VSS.n715 VSS.n714 0.180667
R9918 VSS.n716 VSS.n715 0.180667
R9919 VSS.n717 VSS.n716 0.180667
R9920 VSS.n718 VSS.n717 0.180667
R9921 VSS.n719 VSS.n718 0.180667
R9922 VSS.n720 VSS.n719 0.180667
R9923 VSS.n721 VSS.n720 0.180667
R9924 VSS.n722 VSS.n721 0.180667
R9925 VSS.n723 VSS.n722 0.180667
R9926 VSS.n724 VSS.n723 0.180667
R9927 VSS.n725 VSS.n724 0.180667
R9928 VSS.n726 VSS.n725 0.180667
R9929 VSS.n727 VSS.n726 0.180667
R9930 VSS.n728 VSS.n727 0.180667
R9931 VSS.n729 VSS.n728 0.180667
R9932 VSS.n730 VSS.n729 0.180667
R9933 VSS.n731 VSS.n730 0.180667
R9934 VSS.n732 VSS.n731 0.180667
R9935 VSS.n733 VSS.n732 0.180667
R9936 VSS.n734 VSS.n733 0.180667
R9937 VSS.n735 VSS.n734 0.180667
R9938 VSS.n736 VSS.n735 0.180667
R9939 VSS.n737 VSS.n736 0.180667
R9940 VSS.n738 VSS.n737 0.180667
R9941 VSS.n739 VSS.n738 0.180667
R9942 VSS.n740 VSS.n739 0.180667
R9943 VSS.n741 VSS.n740 0.180667
R9944 VSS.n742 VSS.n741 0.180667
R9945 VSS.n743 VSS.n742 0.180667
R9946 VSS.n744 VSS.n743 0.180667
R9947 VSS.n745 VSS.n744 0.180667
R9948 VSS.n746 VSS.n745 0.180667
R9949 VSS.n747 VSS.n746 0.180667
R9950 VSS.n748 VSS.n747 0.180667
R9951 VSS.n749 VSS.n748 0.180667
R9952 VSS.n750 VSS.n749 0.180667
R9953 VSS.n751 VSS.n750 0.180667
R9954 VSS.n752 VSS.n751 0.180667
R9955 VSS.n753 VSS.n752 0.180667
R9956 VSS.n754 VSS.n753 0.180667
R9957 VSS.n755 VSS.n754 0.180667
R9958 VSS.n756 VSS.n755 0.180667
R9959 VSS.n757 VSS.n756 0.180667
R9960 VSS.n758 VSS.n757 0.180667
R9961 VSS.n759 VSS.n758 0.180667
R9962 VSS.n760 VSS.n759 0.180667
R9963 VSS.n761 VSS.n760 0.180667
R9964 VSS.n762 VSS.n761 0.180667
R9965 VSS.n763 VSS.n762 0.180667
R9966 VSS.n764 VSS.n763 0.180667
R9967 VSS.n765 VSS.n764 0.180667
R9968 VSS.n766 VSS.n765 0.180667
R9969 VSS.n2163 VSS.n2161 0.180304
R9970 VSS.n2901 VSS.n2163 0.180304
R9971 VSS.n2562 VSS.n2227 0.180304
R9972 VSS.n1613 VSS.n1612 0.180304
R9973 VSS.n1537 VSS.n1536 0.180304
R9974 VSS.n4322 VSS.n3726 0.179521
R9975 VSS.n4460 VSS.n4459 0.179521
R9976 VSS.n3219 VSS.n3159 0.179521
R9977 VSS.n3213 VSS.n3212 0.179521
R9978 VSS.n2120 VSS.n2119 0.179521
R9979 VSS.n2114 VSS.n2113 0.179521
R9980 VSS.n2108 VSS.n2107 0.179521
R9981 VSS.n2080 VSS.n2078 0.179521
R9982 VSS.n2586 VSS.n2585 0.179521
R9983 VSS.n2770 VSS.n2769 0.179521
R9984 VSS.n2911 VSS.n2910 0.179521
R9985 VSS.n1599 VSS.n1598 0.179521
R9986 VSS.n1605 VSS.n1541 0.179521
R9987 VSS.n1316 VSS.n1265 0.179521
R9988 VSS.n1309 VSS.n1267 0.179521
R9989 VSS.n2882 VSS.n2847 0.175842
R9990 VSS.n968 VSS.n967 0.171884
R9991 VSS.n4979 VSS.n322 0.164562
R9992 VSS.n5777 VSS.n1 0.1603
R9993 VSS.n3659 VSS.n1 0.1603
R9994 VSS.n3659 VSS.n2939 0.1603
R9995 VSS.n2939 VSS.n382 0.1603
R9996 VSS.n4852 VSS.n382 0.158581
R9997 VSS.n4673 VSS.n635 0.15675
R9998 VSS.n913 VSS.n768 0.15675
R9999 VSS.n4671 VSS.n914 0.155145
R10000 VSS.n346 VSS.n339 0.145413
R10001 VSS.n4672 VSS.n4671 0.144077
R10002 VSS.n3861 VSS.n3860 0.13963
R10003 VSS.n3404 VSS.n3403 0.13963
R10004 VSS.n4050 VSS.n4049 0.13667
R10005 VSS.n4223 VSS.n4222 0.13667
R10006 VSS.n3349 VSS.n3079 0.13667
R10007 VSS.n3294 VSS.n3293 0.13667
R10008 VSS.n3276 VSS.n3275 0.13667
R10009 VSS.n2367 VSS.n2324 0.13667
R10010 VSS.n2373 VSS.n2372 0.13667
R10011 VSS.n2700 VSS.n2699 0.13667
R10012 VSS.n1680 VSS.n1679 0.13667
R10013 VSS.n3941 VSS.n3940 0.132007
R10014 VSS.n3941 VSS.n3820 0.132007
R10015 VSS.n3174 VSS.n3131 0.126304
R10016 VSS.n4979 VSS.n4978 0.122091
R10017 VSS.n334 VSS.n333 0.120292
R10018 VSS.n334 VSS.n326 0.120292
R10019 VSS.n5368 VSS.n5367 0.120292
R10020 VSS.n5368 VSS.n5362 0.120292
R10021 VSS.n5362 VSS.n5360 0.120292
R10022 VSS.n5373 VSS.n5360 0.120292
R10023 VSS.n5374 VSS.n5373 0.120292
R10024 VSS.n5375 VSS.n5374 0.120292
R10025 VSS.n5375 VSS.n5357 0.120292
R10026 VSS.n5379 VSS.n5357 0.120292
R10027 VSS.n5380 VSS.n5379 0.120292
R10028 VSS.n5381 VSS.n5380 0.120292
R10029 VSS.n5381 VSS.n175 0.120292
R10030 VSS.n5385 VSS.n175 0.120292
R10031 VSS.n5386 VSS.n5385 0.120292
R10032 VSS.n5387 VSS.n5386 0.120292
R10033 VSS.n5387 VSS.n172 0.120292
R10034 VSS.n5391 VSS.n172 0.120292
R10035 VSS.n5392 VSS.n5391 0.120292
R10036 VSS.n5393 VSS.n5392 0.120292
R10037 VSS.n5393 VSS.n169 0.120292
R10038 VSS.n169 VSS.n168 0.120292
R10039 VSS.n5399 VSS.n168 0.120292
R10040 VSS.n5400 VSS.n5399 0.120292
R10041 VSS.n5401 VSS.n5400 0.120292
R10042 VSS.n5401 VSS.n166 0.120292
R10043 VSS.n5405 VSS.n166 0.120292
R10044 VSS.n5406 VSS.n5405 0.120292
R10045 VSS.n5407 VSS.n5406 0.120292
R10046 VSS.n5407 VSS.n164 0.120292
R10047 VSS.n5412 VSS.n164 0.120292
R10048 VSS.n5413 VSS.n5412 0.120292
R10049 VSS.n5414 VSS.n5413 0.120292
R10050 VSS.n5414 VSS.n162 0.120292
R10051 VSS.n5419 VSS.n162 0.120292
R10052 VSS.n5420 VSS.n5419 0.120292
R10053 VSS.n5421 VSS.n5420 0.120292
R10054 VSS.n5421 VSS.n159 0.120292
R10055 VSS.n159 VSS.n157 0.120292
R10056 VSS.n157 VSS.n156 0.120292
R10057 VSS.n5428 VSS.n156 0.120292
R10058 VSS.n5429 VSS.n5428 0.120292
R10059 VSS.n5430 VSS.n5429 0.120292
R10060 VSS.n5430 VSS.n154 0.120292
R10061 VSS.n5436 VSS.n154 0.120292
R10062 VSS.n5437 VSS.n5436 0.120292
R10063 VSS.n5437 VSS.n152 0.120292
R10064 VSS.n5441 VSS.n152 0.120292
R10065 VSS.n5442 VSS.n5441 0.120292
R10066 VSS.n5443 VSS.n5442 0.120292
R10067 VSS.n5443 VSS.n150 0.120292
R10068 VSS.n5447 VSS.n150 0.120292
R10069 VSS.n5448 VSS.n5447 0.120292
R10070 VSS.n5448 VSS.n148 0.120292
R10071 VSS.n5453 VSS.n148 0.120292
R10072 VSS.n5454 VSS.n5453 0.120292
R10073 VSS.n5455 VSS.n5454 0.120292
R10074 VSS.n5455 VSS.n145 0.120292
R10075 VSS.n5459 VSS.n145 0.120292
R10076 VSS.n5460 VSS.n5459 0.120292
R10077 VSS.n5461 VSS.n5460 0.120292
R10078 VSS.n5461 VSS.n143 0.120292
R10079 VSS.n5466 VSS.n143 0.120292
R10080 VSS.n137 VSS.n136 0.120292
R10081 VSS.n5473 VSS.n136 0.120292
R10082 VSS.n5474 VSS.n5473 0.120292
R10083 VSS.n5475 VSS.n5474 0.120292
R10084 VSS.n5475 VSS.n134 0.120292
R10085 VSS.n5479 VSS.n134 0.120292
R10086 VSS.n5481 VSS.n5479 0.120292
R10087 VSS.n5481 VSS.n5480 0.120292
R10088 VSS.n5480 VSS.n130 0.120292
R10089 VSS.n5489 VSS.n130 0.120292
R10090 VSS.n5490 VSS.n5489 0.120292
R10091 VSS.n5491 VSS.n5490 0.120292
R10092 VSS.n5491 VSS.n127 0.120292
R10093 VSS.n5495 VSS.n127 0.120292
R10094 VSS.n5496 VSS.n5495 0.120292
R10095 VSS.n5497 VSS.n5496 0.120292
R10096 VSS.n5497 VSS.n124 0.120292
R10097 VSS.n5501 VSS.n124 0.120292
R10098 VSS.n5502 VSS.n5501 0.120292
R10099 VSS.n5503 VSS.n5502 0.120292
R10100 VSS.n5503 VSS.n121 0.120292
R10101 VSS.n5507 VSS.n121 0.120292
R10102 VSS.n5508 VSS.n5507 0.120292
R10103 VSS.n5509 VSS.n5508 0.120292
R10104 VSS.n5509 VSS.n118 0.120292
R10105 VSS.n118 VSS.n117 0.120292
R10106 VSS.n5514 VSS.n117 0.120292
R10107 VSS.n5515 VSS.n5514 0.120292
R10108 VSS.n5516 VSS.n5515 0.120292
R10109 VSS.n5516 VSS.n114 0.120292
R10110 VSS.n114 VSS.n113 0.120292
R10111 VSS.n5522 VSS.n113 0.120292
R10112 VSS.n5523 VSS.n5522 0.120292
R10113 VSS.n5524 VSS.n5523 0.120292
R10114 VSS.n5524 VSS.n111 0.120292
R10115 VSS.n5531 VSS.n111 0.120292
R10116 VSS.n5532 VSS.n5531 0.120292
R10117 VSS.n5533 VSS.n5532 0.120292
R10118 VSS.n5533 VSS.n109 0.120292
R10119 VSS.n5537 VSS.n109 0.120292
R10120 VSS.n5538 VSS.n5537 0.120292
R10121 VSS.n5539 VSS.n5538 0.120292
R10122 VSS.n5539 VSS.n107 0.120292
R10123 VSS.n5544 VSS.n107 0.120292
R10124 VSS.n5545 VSS.n5544 0.120292
R10125 VSS.n5546 VSS.n5545 0.120292
R10126 VSS.n5546 VSS.n105 0.120292
R10127 VSS.n5551 VSS.n105 0.120292
R10128 VSS.n5552 VSS.n5551 0.120292
R10129 VSS.n5553 VSS.n5552 0.120292
R10130 VSS.n5553 VSS.n102 0.120292
R10131 VSS.n5557 VSS.n102 0.120292
R10132 VSS.n5558 VSS.n5557 0.120292
R10133 VSS.n5558 VSS.n100 0.120292
R10134 VSS.n5564 VSS.n100 0.120292
R10135 VSS.n5565 VSS.n5564 0.120292
R10136 VSS.n5566 VSS.n5565 0.120292
R10137 VSS.n5566 VSS.n98 0.120292
R10138 VSS.n5571 VSS.n98 0.120292
R10139 VSS.n5576 VSS.n94 0.120292
R10140 VSS.n5577 VSS.n5576 0.120292
R10141 VSS.n5578 VSS.n5577 0.120292
R10142 VSS.n5578 VSS.n91 0.120292
R10143 VSS.n5582 VSS.n91 0.120292
R10144 VSS.n5583 VSS.n5582 0.120292
R10145 VSS.n5584 VSS.n5583 0.120292
R10146 VSS.n5584 VSS.n89 0.120292
R10147 VSS.n5591 VSS.n89 0.120292
R10148 VSS.n5592 VSS.n5591 0.120292
R10149 VSS.n5593 VSS.n5592 0.120292
R10150 VSS.n5593 VSS.n86 0.120292
R10151 VSS.n5598 VSS.n86 0.120292
R10152 VSS.n5599 VSS.n5598 0.120292
R10153 VSS.n5600 VSS.n5599 0.120292
R10154 VSS.n5600 VSS.n83 0.120292
R10155 VSS.n5604 VSS.n83 0.120292
R10156 VSS.n5605 VSS.n5604 0.120292
R10157 VSS.n5606 VSS.n5605 0.120292
R10158 VSS.n5606 VSS.n80 0.120292
R10159 VSS.n80 VSS.n78 0.120292
R10160 VSS.n78 VSS.n77 0.120292
R10161 VSS.n5613 VSS.n77 0.120292
R10162 VSS.n5614 VSS.n5613 0.120292
R10163 VSS.n5615 VSS.n5614 0.120292
R10164 VSS.n5615 VSS.n75 0.120292
R10165 VSS.n5621 VSS.n75 0.120292
R10166 VSS.n5622 VSS.n5621 0.120292
R10167 VSS.n5622 VSS.n73 0.120292
R10168 VSS.n5626 VSS.n73 0.120292
R10169 VSS.n5627 VSS.n5626 0.120292
R10170 VSS.n5628 VSS.n5627 0.120292
R10171 VSS.n5628 VSS.n71 0.120292
R10172 VSS.n5632 VSS.n71 0.120292
R10173 VSS.n5633 VSS.n5632 0.120292
R10174 VSS.n5633 VSS.n69 0.120292
R10175 VSS.n5637 VSS.n69 0.120292
R10176 VSS.n5638 VSS.n5637 0.120292
R10177 VSS.n5638 VSS.n67 0.120292
R10178 VSS.n5642 VSS.n67 0.120292
R10179 VSS.n5643 VSS.n5642 0.120292
R10180 VSS.n5644 VSS.n5643 0.120292
R10181 VSS.n5644 VSS.n63 0.120292
R10182 VSS.n63 VSS.n62 0.120292
R10183 VSS.n5649 VSS.n62 0.120292
R10184 VSS.n5650 VSS.n5649 0.120292
R10185 VSS.n5651 VSS.n5650 0.120292
R10186 VSS.n5651 VSS.n60 0.120292
R10187 VSS.n60 VSS.n58 0.120292
R10188 VSS.n5657 VSS.n58 0.120292
R10189 VSS.n5658 VSS.n5657 0.120292
R10190 VSS.n5659 VSS.n5658 0.120292
R10191 VSS.n5659 VSS.n56 0.120292
R10192 VSS.n5663 VSS.n56 0.120292
R10193 VSS.n5664 VSS.n5663 0.120292
R10194 VSS.n5664 VSS.n52 0.120292
R10195 VSS.n5671 VSS.n52 0.120292
R10196 VSS.n5672 VSS.n5671 0.120292
R10197 VSS.n5673 VSS.n5672 0.120292
R10198 VSS.n5673 VSS.n49 0.120292
R10199 VSS.n5677 VSS.n49 0.120292
R10200 VSS.n5678 VSS.n5677 0.120292
R10201 VSS.n5679 VSS.n5678 0.120292
R10202 VSS.n5679 VSS.n46 0.120292
R10203 VSS.n5683 VSS.n46 0.120292
R10204 VSS.n5684 VSS.n5683 0.120292
R10205 VSS.n5684 VSS.n43 0.120292
R10206 VSS.n5691 VSS.n5690 0.120292
R10207 VSS.n5691 VSS.n40 0.120292
R10208 VSS.n5695 VSS.n40 0.120292
R10209 VSS.n5696 VSS.n5695 0.120292
R10210 VSS.n5697 VSS.n5696 0.120292
R10211 VSS.n5697 VSS.n36 0.120292
R10212 VSS.n5702 VSS.n36 0.120292
R10213 VSS.n5703 VSS.n5702 0.120292
R10214 VSS.n5704 VSS.n5703 0.120292
R10215 VSS.n5710 VSS.n5709 0.120292
R10216 VSS.n5710 VSS.n31 0.120292
R10217 VSS.n5714 VSS.n31 0.120292
R10218 VSS.n5715 VSS.n5714 0.120292
R10219 VSS.n5716 VSS.n5715 0.120292
R10220 VSS.n5716 VSS.n29 0.120292
R10221 VSS.n5721 VSS.n29 0.120292
R10222 VSS.n5722 VSS.n5721 0.120292
R10223 VSS.n5723 VSS.n5722 0.120292
R10224 VSS.n5723 VSS.n27 0.120292
R10225 VSS.n5728 VSS.n27 0.120292
R10226 VSS.n5729 VSS.n5728 0.120292
R10227 VSS.n5730 VSS.n5729 0.120292
R10228 VSS.n5730 VSS.n24 0.120292
R10229 VSS.n5734 VSS.n24 0.120292
R10230 VSS.n5735 VSS.n5734 0.120292
R10231 VSS.n5736 VSS.n5735 0.120292
R10232 VSS.n5736 VSS.n21 0.120292
R10233 VSS.n5742 VSS.n21 0.120292
R10234 VSS.n5743 VSS.n5742 0.120292
R10235 VSS.n5743 VSS.n18 0.120292
R10236 VSS.n5747 VSS.n18 0.120292
R10237 VSS.n5748 VSS.n5747 0.120292
R10238 VSS.n5748 VSS.n15 0.120292
R10239 VSS.n5755 VSS.n5754 0.120292
R10240 VSS.n5755 VSS.n13 0.120292
R10241 VSS.n5759 VSS.n13 0.120292
R10242 VSS.n5760 VSS.n5759 0.120292
R10243 VSS.n5761 VSS.n5760 0.120292
R10244 VSS.n4566 VSS.n4565 0.120292
R10245 VSS.n4566 VSS.n4563 0.120292
R10246 VSS.n4570 VSS.n4563 0.120292
R10247 VSS.n4571 VSS.n4570 0.120292
R10248 VSS.n4572 VSS.n4571 0.120292
R10249 VSS.n4572 VSS.n4561 0.120292
R10250 VSS.n4576 VSS.n4561 0.120292
R10251 VSS.n4577 VSS.n4576 0.120292
R10252 VSS.n4577 VSS.n4559 0.120292
R10253 VSS.n4581 VSS.n4559 0.120292
R10254 VSS.n4582 VSS.n4581 0.120292
R10255 VSS.n4582 VSS.n4557 0.120292
R10256 VSS.n4557 VSS.n4556 0.120292
R10257 VSS.n4556 VSS.n4555 0.120292
R10258 VSS.n4555 VSS.n4494 0.120292
R10259 VSS.n4549 VSS.n4494 0.120292
R10260 VSS.n4549 VSS.n4548 0.120292
R10261 VSS.n4548 VSS.n4547 0.120292
R10262 VSS.n4547 VSS.n4496 0.120292
R10263 VSS.n4543 VSS.n4496 0.120292
R10264 VSS.n4543 VSS.n4542 0.120292
R10265 VSS.n4542 VSS.n4541 0.120292
R10266 VSS.n4541 VSS.n4498 0.120292
R10267 VSS.n4536 VSS.n4498 0.120292
R10268 VSS.n4536 VSS.n4535 0.120292
R10269 VSS.n4535 VSS.n4534 0.120292
R10270 VSS.n4534 VSS.n4501 0.120292
R10271 VSS.n4530 VSS.n4501 0.120292
R10272 VSS.n4530 VSS.n4529 0.120292
R10273 VSS.n4529 VSS.n4528 0.120292
R10274 VSS.n4528 VSS.n4504 0.120292
R10275 VSS.n4524 VSS.n4504 0.120292
R10276 VSS.n4524 VSS.n4523 0.120292
R10277 VSS.n4523 VSS.n4522 0.120292
R10278 VSS.n4522 VSS.n4507 0.120292
R10279 VSS.n4517 VSS.n4507 0.120292
R10280 VSS.n4517 VSS.n4516 0.120292
R10281 VSS.n4516 VSS.n4515 0.120292
R10282 VSS.n4515 VSS.n4509 0.120292
R10283 VSS.n3856 VSS.n3849 0.120292
R10284 VSS.n3849 VSS.n3847 0.120292
R10285 VSS.n3862 VSS.n3847 0.120292
R10286 VSS.n3863 VSS.n3862 0.120292
R10287 VSS.n3863 VSS.n3844 0.120292
R10288 VSS.n3871 VSS.n3844 0.120292
R10289 VSS.n3872 VSS.n3871 0.120292
R10290 VSS.n3873 VSS.n3872 0.120292
R10291 VSS.n3873 VSS.n3842 0.120292
R10292 VSS.n3879 VSS.n3842 0.120292
R10293 VSS.n3886 VSS.n3839 0.120292
R10294 VSS.n3887 VSS.n3886 0.120292
R10295 VSS.n3888 VSS.n3887 0.120292
R10296 VSS.n3897 VSS.n3896 0.120292
R10297 VSS.n3897 VSS.n3835 0.120292
R10298 VSS.n3902 VSS.n3835 0.120292
R10299 VSS.n3903 VSS.n3902 0.120292
R10300 VSS.n3904 VSS.n3903 0.120292
R10301 VSS.n3904 VSS.n3833 0.120292
R10302 VSS.n3908 VSS.n3833 0.120292
R10303 VSS.n3909 VSS.n3908 0.120292
R10304 VSS.n3909 VSS.n3831 0.120292
R10305 VSS.n3914 VSS.n3831 0.120292
R10306 VSS.n3915 VSS.n3914 0.120292
R10307 VSS.n3915 VSS.n3829 0.120292
R10308 VSS.n3829 VSS.n3827 0.120292
R10309 VSS.n3924 VSS.n3827 0.120292
R10310 VSS.n3925 VSS.n3924 0.120292
R10311 VSS.n3926 VSS.n3925 0.120292
R10312 VSS.n3926 VSS.n3824 0.120292
R10313 VSS.n3933 VSS.n3824 0.120292
R10314 VSS.n3935 VSS.n3933 0.120292
R10315 VSS.n3935 VSS.n3934 0.120292
R10316 VSS.n3934 VSS.n3819 0.120292
R10317 VSS.n3946 VSS.n3819 0.120292
R10318 VSS.n3947 VSS.n3946 0.120292
R10319 VSS.n3948 VSS.n3947 0.120292
R10320 VSS.n3948 VSS.n3817 0.120292
R10321 VSS.n3956 VSS.n3817 0.120292
R10322 VSS.n3957 VSS.n3956 0.120292
R10323 VSS.n3958 VSS.n3957 0.120292
R10324 VSS.n3958 VSS.n3814 0.120292
R10325 VSS.n3964 VSS.n3814 0.120292
R10326 VSS.n3965 VSS.n3964 0.120292
R10327 VSS.n3966 VSS.n3965 0.120292
R10328 VSS.n3966 VSS.n3811 0.120292
R10329 VSS.n3972 VSS.n3811 0.120292
R10330 VSS.n3973 VSS.n3972 0.120292
R10331 VSS.n3974 VSS.n3973 0.120292
R10332 VSS.n3974 VSS.n3809 0.120292
R10333 VSS.n3980 VSS.n3809 0.120292
R10334 VSS.n3981 VSS.n3980 0.120292
R10335 VSS.n4053 VSS.n3981 0.120292
R10336 VSS.n4053 VSS.n4052 0.120292
R10337 VSS.n4052 VSS.n4051 0.120292
R10338 VSS.n4051 VSS.n3982 0.120292
R10339 VSS.n4045 VSS.n3982 0.120292
R10340 VSS.n4045 VSS.n4044 0.120292
R10341 VSS.n4044 VSS.n3984 0.120292
R10342 VSS.n4040 VSS.n3984 0.120292
R10343 VSS.n4040 VSS.n4039 0.120292
R10344 VSS.n4039 VSS.n4038 0.120292
R10345 VSS.n4038 VSS.n3987 0.120292
R10346 VSS.n4034 VSS.n3987 0.120292
R10347 VSS.n4034 VSS.n4033 0.120292
R10348 VSS.n4033 VSS.n4032 0.120292
R10349 VSS.n4032 VSS.n3992 0.120292
R10350 VSS.n4024 VSS.n3992 0.120292
R10351 VSS.n4024 VSS.n4023 0.120292
R10352 VSS.n4023 VSS.n4022 0.120292
R10353 VSS.n4022 VSS.n3994 0.120292
R10354 VSS.n4018 VSS.n3994 0.120292
R10355 VSS.n4018 VSS.n4017 0.120292
R10356 VSS.n4017 VSS.n4016 0.120292
R10357 VSS.n4016 VSS.n3997 0.120292
R10358 VSS.n4012 VSS.n3997 0.120292
R10359 VSS.n4012 VSS.n4011 0.120292
R10360 VSS.n4011 VSS.n4000 0.120292
R10361 VSS.n4006 VSS.n4000 0.120292
R10362 VSS.n4006 VSS.n4005 0.120292
R10363 VSS.n4005 VSS.n3805 0.120292
R10364 VSS.n4059 VSS.n3805 0.120292
R10365 VSS.n4060 VSS.n4059 0.120292
R10366 VSS.n4061 VSS.n4060 0.120292
R10367 VSS.n4061 VSS.n3803 0.120292
R10368 VSS.n4066 VSS.n3803 0.120292
R10369 VSS.n4067 VSS.n4066 0.120292
R10370 VSS.n4068 VSS.n4067 0.120292
R10371 VSS.n4068 VSS.n3800 0.120292
R10372 VSS.n4074 VSS.n3800 0.120292
R10373 VSS.n4075 VSS.n4074 0.120292
R10374 VSS.n4076 VSS.n4075 0.120292
R10375 VSS.n4076 VSS.n3798 0.120292
R10376 VSS.n4081 VSS.n3798 0.120292
R10377 VSS.n4082 VSS.n4081 0.120292
R10378 VSS.n4082 VSS.n3794 0.120292
R10379 VSS.n4089 VSS.n3794 0.120292
R10380 VSS.n4090 VSS.n4089 0.120292
R10381 VSS.n4091 VSS.n4090 0.120292
R10382 VSS.n4091 VSS.n3790 0.120292
R10383 VSS.n4095 VSS.n3790 0.120292
R10384 VSS.n4096 VSS.n4095 0.120292
R10385 VSS.n4096 VSS.n3786 0.120292
R10386 VSS.n4101 VSS.n3786 0.120292
R10387 VSS.n4102 VSS.n4101 0.120292
R10388 VSS.n4103 VSS.n4102 0.120292
R10389 VSS.n4103 VSS.n3782 0.120292
R10390 VSS.n4110 VSS.n3782 0.120292
R10391 VSS.n4111 VSS.n4110 0.120292
R10392 VSS.n4111 VSS.n3779 0.120292
R10393 VSS.n4117 VSS.n3779 0.120292
R10394 VSS.n4118 VSS.n4117 0.120292
R10395 VSS.n4119 VSS.n4118 0.120292
R10396 VSS.n4119 VSS.n3776 0.120292
R10397 VSS.n4125 VSS.n3776 0.120292
R10398 VSS.n4126 VSS.n4125 0.120292
R10399 VSS.n4127 VSS.n4126 0.120292
R10400 VSS.n4127 VSS.n3772 0.120292
R10401 VSS.n4133 VSS.n3772 0.120292
R10402 VSS.n4134 VSS.n4133 0.120292
R10403 VSS.n4135 VSS.n4134 0.120292
R10404 VSS.n4135 VSS.n3770 0.120292
R10405 VSS.n4141 VSS.n3770 0.120292
R10406 VSS.n4142 VSS.n4141 0.120292
R10407 VSS.n4143 VSS.n4142 0.120292
R10408 VSS.n4143 VSS.n3768 0.120292
R10409 VSS.n4149 VSS.n3768 0.120292
R10410 VSS.n4150 VSS.n4149 0.120292
R10411 VSS.n4151 VSS.n4150 0.120292
R10412 VSS.n4151 VSS.n3765 0.120292
R10413 VSS.n4157 VSS.n3765 0.120292
R10414 VSS.n4158 VSS.n4157 0.120292
R10415 VSS.n4159 VSS.n4158 0.120292
R10416 VSS.n4159 VSS.n3762 0.120292
R10417 VSS.n4164 VSS.n3762 0.120292
R10418 VSS.n4165 VSS.n4164 0.120292
R10419 VSS.n4166 VSS.n4165 0.120292
R10420 VSS.n4237 VSS.n4166 0.120292
R10421 VSS.n4237 VSS.n4236 0.120292
R10422 VSS.n4236 VSS.n4235 0.120292
R10423 VSS.n4235 VSS.n4169 0.120292
R10424 VSS.n4229 VSS.n4169 0.120292
R10425 VSS.n4229 VSS.n4228 0.120292
R10426 VSS.n4228 VSS.n4227 0.120292
R10427 VSS.n4227 VSS.n4172 0.120292
R10428 VSS.n4220 VSS.n4172 0.120292
R10429 VSS.n4220 VSS.n4219 0.120292
R10430 VSS.n4219 VSS.n4218 0.120292
R10431 VSS.n4218 VSS.n4175 0.120292
R10432 VSS.n4212 VSS.n4175 0.120292
R10433 VSS.n4212 VSS.n4211 0.120292
R10434 VSS.n4211 VSS.n4210 0.120292
R10435 VSS.n4210 VSS.n4180 0.120292
R10436 VSS.n4206 VSS.n4180 0.120292
R10437 VSS.n4206 VSS.n4205 0.120292
R10438 VSS.n4205 VSS.n4183 0.120292
R10439 VSS.n4200 VSS.n4183 0.120292
R10440 VSS.n4200 VSS.n4199 0.120292
R10441 VSS.n4199 VSS.n4198 0.120292
R10442 VSS.n4198 VSS.n4186 0.120292
R10443 VSS.n4188 VSS.n4186 0.120292
R10444 VSS.n4193 VSS.n4188 0.120292
R10445 VSS.n4193 VSS.n4192 0.120292
R10446 VSS.n4192 VSS.n4191 0.120292
R10447 VSS.n4191 VSS.n3759 0.120292
R10448 VSS.n4245 VSS.n3759 0.120292
R10449 VSS.n4246 VSS.n4245 0.120292
R10450 VSS.n4247 VSS.n4246 0.120292
R10451 VSS.n4247 VSS.n3757 0.120292
R10452 VSS.n4252 VSS.n3757 0.120292
R10453 VSS.n4253 VSS.n4252 0.120292
R10454 VSS.n4253 VSS.n3755 0.120292
R10455 VSS.n4258 VSS.n3755 0.120292
R10456 VSS.n4259 VSS.n4258 0.120292
R10457 VSS.n4259 VSS.n3751 0.120292
R10458 VSS.n4264 VSS.n3751 0.120292
R10459 VSS.n4265 VSS.n4264 0.120292
R10460 VSS.n4265 VSS.n3749 0.120292
R10461 VSS.n4269 VSS.n3749 0.120292
R10462 VSS.n4270 VSS.n4269 0.120292
R10463 VSS.n4271 VSS.n4270 0.120292
R10464 VSS.n4271 VSS.n3746 0.120292
R10465 VSS.n4277 VSS.n3746 0.120292
R10466 VSS.n4278 VSS.n4277 0.120292
R10467 VSS.n4279 VSS.n4278 0.120292
R10468 VSS.n4279 VSS.n3744 0.120292
R10469 VSS.n4284 VSS.n3744 0.120292
R10470 VSS.n4285 VSS.n4284 0.120292
R10471 VSS.n4285 VSS.n3741 0.120292
R10472 VSS.n4290 VSS.n3741 0.120292
R10473 VSS.n4291 VSS.n4290 0.120292
R10474 VSS.n4292 VSS.n4291 0.120292
R10475 VSS.n4292 VSS.n3736 0.120292
R10476 VSS.n4297 VSS.n3736 0.120292
R10477 VSS.n4298 VSS.n4297 0.120292
R10478 VSS.n4298 VSS.n3734 0.120292
R10479 VSS.n4305 VSS.n3734 0.120292
R10480 VSS.n4306 VSS.n4305 0.120292
R10481 VSS.n4306 VSS.n3731 0.120292
R10482 VSS.n4310 VSS.n3731 0.120292
R10483 VSS.n4311 VSS.n4310 0.120292
R10484 VSS.n4311 VSS.n3729 0.120292
R10485 VSS.n4317 VSS.n3729 0.120292
R10486 VSS.n4318 VSS.n4317 0.120292
R10487 VSS.n4318 VSS.n3727 0.120292
R10488 VSS.n4323 VSS.n3727 0.120292
R10489 VSS.n4324 VSS.n4323 0.120292
R10490 VSS.n4324 VSS.n3724 0.120292
R10491 VSS.n4330 VSS.n3724 0.120292
R10492 VSS.n4331 VSS.n4330 0.120292
R10493 VSS.n4331 VSS.n3722 0.120292
R10494 VSS.n4336 VSS.n3722 0.120292
R10495 VSS.n4337 VSS.n4336 0.120292
R10496 VSS.n4337 VSS.n3719 0.120292
R10497 VSS.n4342 VSS.n3719 0.120292
R10498 VSS.n4343 VSS.n4342 0.120292
R10499 VSS.n4344 VSS.n4343 0.120292
R10500 VSS.n4344 VSS.n3717 0.120292
R10501 VSS.n4350 VSS.n3717 0.120292
R10502 VSS.n4351 VSS.n4350 0.120292
R10503 VSS.n4352 VSS.n4351 0.120292
R10504 VSS.n4352 VSS.n3713 0.120292
R10505 VSS.n4361 VSS.n3713 0.120292
R10506 VSS.n4362 VSS.n4361 0.120292
R10507 VSS.n4363 VSS.n4362 0.120292
R10508 VSS.n4363 VSS.n3710 0.120292
R10509 VSS.n4368 VSS.n3710 0.120292
R10510 VSS.n4369 VSS.n4368 0.120292
R10511 VSS.n4370 VSS.n4369 0.120292
R10512 VSS.n4370 VSS.n3707 0.120292
R10513 VSS.n4375 VSS.n3707 0.120292
R10514 VSS.n4376 VSS.n4375 0.120292
R10515 VSS.n4382 VSS.n4376 0.120292
R10516 VSS.n4401 VSS.n4400 0.120292
R10517 VSS.n4401 VSS.n3697 0.120292
R10518 VSS.n4406 VSS.n3697 0.120292
R10519 VSS.n4407 VSS.n4406 0.120292
R10520 VSS.n4407 VSS.n3694 0.120292
R10521 VSS.n4413 VSS.n3694 0.120292
R10522 VSS.n4414 VSS.n4413 0.120292
R10523 VSS.n4415 VSS.n4414 0.120292
R10524 VSS.n4415 VSS.n3692 0.120292
R10525 VSS.n4419 VSS.n3692 0.120292
R10526 VSS.n4420 VSS.n4419 0.120292
R10527 VSS.n4421 VSS.n4420 0.120292
R10528 VSS.n4489 VSS.n4421 0.120292
R10529 VSS.n4489 VSS.n4488 0.120292
R10530 VSS.n4488 VSS.n4487 0.120292
R10531 VSS.n4487 VSS.n4424 0.120292
R10532 VSS.n4481 VSS.n4424 0.120292
R10533 VSS.n4481 VSS.n4480 0.120292
R10534 VSS.n4480 VSS.n4479 0.120292
R10535 VSS.n4479 VSS.n4427 0.120292
R10536 VSS.n4475 VSS.n4427 0.120292
R10537 VSS.n4475 VSS.n4474 0.120292
R10538 VSS.n4474 VSS.n4430 0.120292
R10539 VSS.n4470 VSS.n4430 0.120292
R10540 VSS.n4470 VSS.n4469 0.120292
R10541 VSS.n4469 VSS.n4432 0.120292
R10542 VSS.n4464 VSS.n4432 0.120292
R10543 VSS.n4464 VSS.n4463 0.120292
R10544 VSS.n4463 VSS.n4435 0.120292
R10545 VSS.n4457 VSS.n4435 0.120292
R10546 VSS.n4457 VSS.n4456 0.120292
R10547 VSS.n4456 VSS.n4455 0.120292
R10548 VSS.n4455 VSS.n4439 0.120292
R10549 VSS.n4451 VSS.n4439 0.120292
R10550 VSS.n4451 VSS.n4450 0.120292
R10551 VSS.n4450 VSS.n4449 0.120292
R10552 VSS.n3147 VSS.n3146 0.120292
R10553 VSS.n3148 VSS.n3147 0.120292
R10554 VSS.n3148 VSS.n3136 0.120292
R10555 VSS.n3154 VSS.n3136 0.120292
R10556 VSS.n3155 VSS.n3154 0.120292
R10557 VSS.n3227 VSS.n3155 0.120292
R10558 VSS.n3227 VSS.n3226 0.120292
R10559 VSS.n3226 VSS.n3225 0.120292
R10560 VSS.n3225 VSS.n3156 0.120292
R10561 VSS.n3218 VSS.n3156 0.120292
R10562 VSS.n3218 VSS.n3217 0.120292
R10563 VSS.n3217 VSS.n3160 0.120292
R10564 VSS.n3211 VSS.n3160 0.120292
R10565 VSS.n3211 VSS.n3210 0.120292
R10566 VSS.n3210 VSS.n3209 0.120292
R10567 VSS.n3209 VSS.n3163 0.120292
R10568 VSS.n3205 VSS.n3163 0.120292
R10569 VSS.n3205 VSS.n3204 0.120292
R10570 VSS.n3204 VSS.n3166 0.120292
R10571 VSS.n3200 VSS.n3166 0.120292
R10572 VSS.n3200 VSS.n3199 0.120292
R10573 VSS.n3199 VSS.n3168 0.120292
R10574 VSS.n3193 VSS.n3168 0.120292
R10575 VSS.n3193 VSS.n3192 0.120292
R10576 VSS.n3192 VSS.n3191 0.120292
R10577 VSS.n3191 VSS.n3170 0.120292
R10578 VSS.n3186 VSS.n3170 0.120292
R10579 VSS.n3186 VSS.n3185 0.120292
R10580 VSS.n3185 VSS.n3184 0.120292
R10581 VSS.n3184 VSS.n3173 0.120292
R10582 VSS.n3179 VSS.n3173 0.120292
R10583 VSS.n3179 VSS.n3178 0.120292
R10584 VSS.n3178 VSS.n3132 0.120292
R10585 VSS.n3233 VSS.n3132 0.120292
R10586 VSS.n3234 VSS.n3233 0.120292
R10587 VSS.n3234 VSS.n3130 0.120292
R10588 VSS.n3240 VSS.n3130 0.120292
R10589 VSS.n3245 VSS.n3126 0.120292
R10590 VSS.n3246 VSS.n3245 0.120292
R10591 VSS.n3247 VSS.n3246 0.120292
R10592 VSS.n3247 VSS.n3123 0.120292
R10593 VSS.n3252 VSS.n3123 0.120292
R10594 VSS.n3253 VSS.n3252 0.120292
R10595 VSS.n3254 VSS.n3253 0.120292
R10596 VSS.n3254 VSS.n3121 0.120292
R10597 VSS.n3121 VSS.n3119 0.120292
R10598 VSS.n3260 VSS.n3119 0.120292
R10599 VSS.n3261 VSS.n3260 0.120292
R10600 VSS.n3261 VSS.n3116 0.120292
R10601 VSS.n3265 VSS.n3116 0.120292
R10602 VSS.n3266 VSS.n3265 0.120292
R10603 VSS.n3267 VSS.n3266 0.120292
R10604 VSS.n3267 VSS.n3114 0.120292
R10605 VSS.n3273 VSS.n3114 0.120292
R10606 VSS.n3274 VSS.n3273 0.120292
R10607 VSS.n3274 VSS.n3108 0.120292
R10608 VSS.n3281 VSS.n3108 0.120292
R10609 VSS.n3282 VSS.n3281 0.120292
R10610 VSS.n3283 VSS.n3282 0.120292
R10611 VSS.n3283 VSS.n3104 0.120292
R10612 VSS.n3290 VSS.n3104 0.120292
R10613 VSS.n3291 VSS.n3290 0.120292
R10614 VSS.n3291 VSS.n3101 0.120292
R10615 VSS.n3297 VSS.n3101 0.120292
R10616 VSS.n3299 VSS.n3297 0.120292
R10617 VSS.n3299 VSS.n3298 0.120292
R10618 VSS.n3298 VSS.n3096 0.120292
R10619 VSS.n3308 VSS.n3096 0.120292
R10620 VSS.n3309 VSS.n3308 0.120292
R10621 VSS.n3309 VSS.n3093 0.120292
R10622 VSS.n3315 VSS.n3093 0.120292
R10623 VSS.n3316 VSS.n3315 0.120292
R10624 VSS.n3317 VSS.n3316 0.120292
R10625 VSS.n3317 VSS.n3089 0.120292
R10626 VSS.n3321 VSS.n3089 0.120292
R10627 VSS.n3322 VSS.n3321 0.120292
R10628 VSS.n3323 VSS.n3322 0.120292
R10629 VSS.n3323 VSS.n3087 0.120292
R10630 VSS.n3335 VSS.n3087 0.120292
R10631 VSS.n3336 VSS.n3335 0.120292
R10632 VSS.n3337 VSS.n3336 0.120292
R10633 VSS.n3337 VSS.n3084 0.120292
R10634 VSS.n3341 VSS.n3084 0.120292
R10635 VSS.n3342 VSS.n3341 0.120292
R10636 VSS.n3343 VSS.n3342 0.120292
R10637 VSS.n3343 VSS.n3080 0.120292
R10638 VSS.n3347 VSS.n3080 0.120292
R10639 VSS.n3348 VSS.n3347 0.120292
R10640 VSS.n3348 VSS.n3078 0.120292
R10641 VSS.n3353 VSS.n3078 0.120292
R10642 VSS.n3354 VSS.n3353 0.120292
R10643 VSS.n3355 VSS.n3354 0.120292
R10644 VSS.n3355 VSS.n3074 0.120292
R10645 VSS.n3364 VSS.n3074 0.120292
R10646 VSS.n3365 VSS.n3364 0.120292
R10647 VSS.n3366 VSS.n3365 0.120292
R10648 VSS.n3366 VSS.n3070 0.120292
R10649 VSS.n3371 VSS.n3070 0.120292
R10650 VSS.n3372 VSS.n3371 0.120292
R10651 VSS.n3373 VSS.n3372 0.120292
R10652 VSS.n3373 VSS.n3068 0.120292
R10653 VSS.n3377 VSS.n3068 0.120292
R10654 VSS.n3378 VSS.n3377 0.120292
R10655 VSS.n3379 VSS.n3378 0.120292
R10656 VSS.n3379 VSS.n3066 0.120292
R10657 VSS.n3385 VSS.n3066 0.120292
R10658 VSS.n3386 VSS.n3385 0.120292
R10659 VSS.n3386 VSS.n3063 0.120292
R10660 VSS.n3390 VSS.n3063 0.120292
R10661 VSS.n3391 VSS.n3390 0.120292
R10662 VSS.n3391 VSS.n3061 0.120292
R10663 VSS.n3397 VSS.n3061 0.120292
R10664 VSS.n3398 VSS.n3397 0.120292
R10665 VSS.n3399 VSS.n3398 0.120292
R10666 VSS.n3399 VSS.n3056 0.120292
R10667 VSS.n3407 VSS.n3056 0.120292
R10668 VSS.n3408 VSS.n3407 0.120292
R10669 VSS.n3408 VSS.n3054 0.120292
R10670 VSS.n3054 VSS.n3052 0.120292
R10671 VSS.n3413 VSS.n3052 0.120292
R10672 VSS.n3414 VSS.n3413 0.120292
R10673 VSS.n3415 VSS.n3414 0.120292
R10674 VSS.n3415 VSS.n3048 0.120292
R10675 VSS.n3419 VSS.n3048 0.120292
R10676 VSS.n3420 VSS.n3419 0.120292
R10677 VSS.n3421 VSS.n3420 0.120292
R10678 VSS.n3421 VSS.n3044 0.120292
R10679 VSS.n3425 VSS.n3044 0.120292
R10680 VSS.n3426 VSS.n3425 0.120292
R10681 VSS.n3427 VSS.n3426 0.120292
R10682 VSS.n3427 VSS.n3041 0.120292
R10683 VSS.n3432 VSS.n3041 0.120292
R10684 VSS.n3433 VSS.n3432 0.120292
R10685 VSS.n3433 VSS.n3038 0.120292
R10686 VSS.n3439 VSS.n3038 0.120292
R10687 VSS.n3440 VSS.n3439 0.120292
R10688 VSS.n3441 VSS.n3440 0.120292
R10689 VSS.n3441 VSS.n3036 0.120292
R10690 VSS.n3036 VSS.n3035 0.120292
R10691 VSS.n3450 VSS.n3035 0.120292
R10692 VSS.n3451 VSS.n3450 0.120292
R10693 VSS.n3451 VSS.n3032 0.120292
R10694 VSS.n3458 VSS.n3032 0.120292
R10695 VSS.n3459 VSS.n3458 0.120292
R10696 VSS.n3460 VSS.n3459 0.120292
R10697 VSS.n3460 VSS.n3028 0.120292
R10698 VSS.n3467 VSS.n3028 0.120292
R10699 VSS.n3468 VSS.n3467 0.120292
R10700 VSS.n3469 VSS.n3468 0.120292
R10701 VSS.n3469 VSS.n3026 0.120292
R10702 VSS.n3475 VSS.n3026 0.120292
R10703 VSS.n3476 VSS.n3475 0.120292
R10704 VSS.n3477 VSS.n3476 0.120292
R10705 VSS.n3477 VSS.n3024 0.120292
R10706 VSS.n3024 VSS.n3021 0.120292
R10707 VSS.n3021 VSS.n3019 0.120292
R10708 VSS.n3483 VSS.n3019 0.120292
R10709 VSS.n3484 VSS.n3483 0.120292
R10710 VSS.n3484 VSS.n3015 0.120292
R10711 VSS.n3492 VSS.n3015 0.120292
R10712 VSS.n3493 VSS.n3492 0.120292
R10713 VSS.n3493 VSS.n3013 0.120292
R10714 VSS.n3500 VSS.n3013 0.120292
R10715 VSS.n3501 VSS.n3500 0.120292
R10716 VSS.n3501 VSS.n3011 0.120292
R10717 VSS.n3011 VSS.n3009 0.120292
R10718 VSS.n3506 VSS.n3009 0.120292
R10719 VSS.n3507 VSS.n3506 0.120292
R10720 VSS.n3507 VSS.n3004 0.120292
R10721 VSS.n3513 VSS.n3004 0.120292
R10722 VSS.n3514 VSS.n3513 0.120292
R10723 VSS.n3515 VSS.n3514 0.120292
R10724 VSS.n3515 VSS.n3001 0.120292
R10725 VSS.n3520 VSS.n3001 0.120292
R10726 VSS.n3521 VSS.n3520 0.120292
R10727 VSS.n3522 VSS.n3521 0.120292
R10728 VSS.n3522 VSS.n2998 0.120292
R10729 VSS.n3530 VSS.n2998 0.120292
R10730 VSS.n3531 VSS.n3530 0.120292
R10731 VSS.n3531 VSS.n2996 0.120292
R10732 VSS.n3535 VSS.n2996 0.120292
R10733 VSS.n3536 VSS.n3535 0.120292
R10734 VSS.n3536 VSS.n2992 0.120292
R10735 VSS.n3540 VSS.n2992 0.120292
R10736 VSS.n3541 VSS.n3540 0.120292
R10737 VSS.n3542 VSS.n3541 0.120292
R10738 VSS.n3542 VSS.n2990 0.120292
R10739 VSS.n3546 VSS.n2990 0.120292
R10740 VSS.n3547 VSS.n3546 0.120292
R10741 VSS.n3549 VSS.n3547 0.120292
R10742 VSS.n3549 VSS.n3548 0.120292
R10743 VSS.n3548 VSS.n2986 0.120292
R10744 VSS.n3558 VSS.n2986 0.120292
R10745 VSS.n3559 VSS.n3558 0.120292
R10746 VSS.n3560 VSS.n3559 0.120292
R10747 VSS.n3560 VSS.n2984 0.120292
R10748 VSS.n2984 VSS.n2980 0.120292
R10749 VSS.n3566 VSS.n2980 0.120292
R10750 VSS.n3567 VSS.n3566 0.120292
R10751 VSS.n3568 VSS.n3567 0.120292
R10752 VSS.n3568 VSS.n2978 0.120292
R10753 VSS.n3575 VSS.n2978 0.120292
R10754 VSS.n3576 VSS.n3575 0.120292
R10755 VSS.n3576 VSS.n2976 0.120292
R10756 VSS.n2976 VSS.n2975 0.120292
R10757 VSS.n2975 VSS.n2973 0.120292
R10758 VSS.n2973 VSS.n2969 0.120292
R10759 VSS.n3585 VSS.n2969 0.120292
R10760 VSS.n3586 VSS.n3585 0.120292
R10761 VSS.n3586 VSS.n2967 0.120292
R10762 VSS.n3597 VSS.n2967 0.120292
R10763 VSS.n3598 VSS.n3597 0.120292
R10764 VSS.n3599 VSS.n3598 0.120292
R10765 VSS.n3599 VSS.n2965 0.120292
R10766 VSS.n3604 VSS.n2965 0.120292
R10767 VSS.n3606 VSS.n3604 0.120292
R10768 VSS.n3606 VSS.n3605 0.120292
R10769 VSS.n3605 VSS.n2960 0.120292
R10770 VSS.n3615 VSS.n2960 0.120292
R10771 VSS.n3616 VSS.n3615 0.120292
R10772 VSS.n3617 VSS.n3616 0.120292
R10773 VSS.n3617 VSS.n2957 0.120292
R10774 VSS.n3624 VSS.n2957 0.120292
R10775 VSS.n3625 VSS.n3624 0.120292
R10776 VSS.n3625 VSS.n2953 0.120292
R10777 VSS.n3629 VSS.n2953 0.120292
R10778 VSS.n3630 VSS.n3629 0.120292
R10779 VSS.n3631 VSS.n3630 0.120292
R10780 VSS.n3631 VSS.n2951 0.120292
R10781 VSS.n2951 VSS.n2949 0.120292
R10782 VSS.n2949 VSS.n2948 0.120292
R10783 VSS.n2948 VSS.n2945 0.120292
R10784 VSS.n3638 VSS.n2945 0.120292
R10785 VSS.n3639 VSS.n3638 0.120292
R10786 VSS.n3641 VSS.n3639 0.120292
R10787 VSS.n3641 VSS.n3640 0.120292
R10788 VSS.n3640 VSS.n2941 0.120292
R10789 VSS.n3650 VSS.n2941 0.120292
R10790 VSS.n3671 VSS.n3670 0.120292
R10791 VSS.n3672 VSS.n3671 0.120292
R10792 VSS.n3672 VSS.n2136 0.120292
R10793 VSS.n3677 VSS.n2136 0.120292
R10794 VSS.n3678 VSS.n3677 0.120292
R10795 VSS.n3679 VSS.n3678 0.120292
R10796 VSS.n3679 VSS.n2134 0.120292
R10797 VSS.n2134 VSS.n2131 0.120292
R10798 VSS.n3685 VSS.n2131 0.120292
R10799 VSS.n3686 VSS.n3685 0.120292
R10800 VSS.n3687 VSS.n3686 0.120292
R10801 VSS.n3687 VSS.n2129 0.120292
R10802 VSS.n2129 VSS.n2128 0.120292
R10803 VSS.n2117 VSS.n2072 0.120292
R10804 VSS.n2117 VSS.n2116 0.120292
R10805 VSS.n2116 VSS.n2074 0.120292
R10806 VSS.n2111 VSS.n2074 0.120292
R10807 VSS.n2111 VSS.n2110 0.120292
R10808 VSS.n2110 VSS.n2076 0.120292
R10809 VSS.n2105 VSS.n2076 0.120292
R10810 VSS.n2105 VSS.n2104 0.120292
R10811 VSS.n2104 VSS.n2079 0.120292
R10812 VSS.n2100 VSS.n2079 0.120292
R10813 VSS.n2100 VSS.n2099 0.120292
R10814 VSS.n2099 VSS.n2098 0.120292
R10815 VSS.n2098 VSS.n2084 0.120292
R10816 VSS.n2093 VSS.n2084 0.120292
R10817 VSS.n2093 VSS.n2092 0.120292
R10818 VSS.n2345 VSS.n2338 0.120292
R10819 VSS.n2338 VSS.n2336 0.120292
R10820 VSS.n2351 VSS.n2336 0.120292
R10821 VSS.n2352 VSS.n2351 0.120292
R10822 VSS.n2352 VSS.n2334 0.120292
R10823 VSS.n2334 VSS.n2332 0.120292
R10824 VSS.n2359 VSS.n2332 0.120292
R10825 VSS.n2360 VSS.n2359 0.120292
R10826 VSS.n2360 VSS.n2329 0.120292
R10827 VSS.n2329 VSS.n2328 0.120292
R10828 VSS.n2328 VSS.n2327 0.120292
R10829 VSS.n2327 VSS.n2326 0.120292
R10830 VSS.n2326 VSS.n2325 0.120292
R10831 VSS.n2369 VSS.n2325 0.120292
R10832 VSS.n2370 VSS.n2369 0.120292
R10833 VSS.n2370 VSS.n2323 0.120292
R10834 VSS.n2375 VSS.n2323 0.120292
R10835 VSS.n2376 VSS.n2375 0.120292
R10836 VSS.n2376 VSS.n2321 0.120292
R10837 VSS.n2381 VSS.n2321 0.120292
R10838 VSS.n2382 VSS.n2381 0.120292
R10839 VSS.n2391 VSS.n2390 0.120292
R10840 VSS.n2392 VSS.n2391 0.120292
R10841 VSS.n2392 VSS.n2317 0.120292
R10842 VSS.n2396 VSS.n2317 0.120292
R10843 VSS.n2397 VSS.n2396 0.120292
R10844 VSS.n2397 VSS.n2315 0.120292
R10845 VSS.n2403 VSS.n2315 0.120292
R10846 VSS.n2404 VSS.n2403 0.120292
R10847 VSS.n2405 VSS.n2404 0.120292
R10848 VSS.n2405 VSS.n2311 0.120292
R10849 VSS.n2410 VSS.n2311 0.120292
R10850 VSS.n2411 VSS.n2410 0.120292
R10851 VSS.n2411 VSS.n2309 0.120292
R10852 VSS.n2418 VSS.n2309 0.120292
R10853 VSS.n2419 VSS.n2418 0.120292
R10854 VSS.n2420 VSS.n2419 0.120292
R10855 VSS.n2420 VSS.n2307 0.120292
R10856 VSS.n2425 VSS.n2307 0.120292
R10857 VSS.n2426 VSS.n2425 0.120292
R10858 VSS.n2426 VSS.n2304 0.120292
R10859 VSS.n2431 VSS.n2304 0.120292
R10860 VSS.n2432 VSS.n2431 0.120292
R10861 VSS.n2432 VSS.n2302 0.120292
R10862 VSS.n2436 VSS.n2302 0.120292
R10863 VSS.n2437 VSS.n2436 0.120292
R10864 VSS.n2437 VSS.n2298 0.120292
R10865 VSS.n2441 VSS.n2298 0.120292
R10866 VSS.n2442 VSS.n2441 0.120292
R10867 VSS.n2443 VSS.n2442 0.120292
R10868 VSS.n2443 VSS.n2296 0.120292
R10869 VSS.n2296 VSS.n2294 0.120292
R10870 VSS.n2294 VSS.n2293 0.120292
R10871 VSS.n2293 VSS.n2291 0.120292
R10872 VSS.n2291 VSS.n2290 0.120292
R10873 VSS.n2290 VSS.n2288 0.120292
R10874 VSS.n2452 VSS.n2288 0.120292
R10875 VSS.n2453 VSS.n2452 0.120292
R10876 VSS.n2454 VSS.n2453 0.120292
R10877 VSS.n2454 VSS.n2285 0.120292
R10878 VSS.n2461 VSS.n2285 0.120292
R10879 VSS.n2462 VSS.n2461 0.120292
R10880 VSS.n2462 VSS.n2282 0.120292
R10881 VSS.n2467 VSS.n2282 0.120292
R10882 VSS.n2468 VSS.n2467 0.120292
R10883 VSS.n2469 VSS.n2468 0.120292
R10884 VSS.n2469 VSS.n2279 0.120292
R10885 VSS.n2474 VSS.n2279 0.120292
R10886 VSS.n2475 VSS.n2474 0.120292
R10887 VSS.n2475 VSS.n2274 0.120292
R10888 VSS.n2480 VSS.n2274 0.120292
R10889 VSS.n2481 VSS.n2480 0.120292
R10890 VSS.n2482 VSS.n2481 0.120292
R10891 VSS.n2482 VSS.n2272 0.120292
R10892 VSS.n2272 VSS.n2271 0.120292
R10893 VSS.n2489 VSS.n2271 0.120292
R10894 VSS.n2490 VSS.n2489 0.120292
R10895 VSS.n2490 VSS.n2269 0.120292
R10896 VSS.n2269 VSS.n2266 0.120292
R10897 VSS.n2495 VSS.n2266 0.120292
R10898 VSS.n2496 VSS.n2495 0.120292
R10899 VSS.n2497 VSS.n2496 0.120292
R10900 VSS.n2497 VSS.n2264 0.120292
R10901 VSS.n2264 VSS.n2261 0.120292
R10902 VSS.n2261 VSS.n2256 0.120292
R10903 VSS.n2504 VSS.n2256 0.120292
R10904 VSS.n2505 VSS.n2504 0.120292
R10905 VSS.n2506 VSS.n2505 0.120292
R10906 VSS.n2506 VSS.n2252 0.120292
R10907 VSS.n2513 VSS.n2252 0.120292
R10908 VSS.n2514 VSS.n2513 0.120292
R10909 VSS.n2515 VSS.n2514 0.120292
R10910 VSS.n2515 VSS.n2250 0.120292
R10911 VSS.n2521 VSS.n2250 0.120292
R10912 VSS.n2522 VSS.n2521 0.120292
R10913 VSS.n2523 VSS.n2522 0.120292
R10914 VSS.n2523 VSS.n2248 0.120292
R10915 VSS.n2528 VSS.n2248 0.120292
R10916 VSS.n2529 VSS.n2528 0.120292
R10917 VSS.n2529 VSS.n2245 0.120292
R10918 VSS.n2534 VSS.n2245 0.120292
R10919 VSS.n2535 VSS.n2534 0.120292
R10920 VSS.n2536 VSS.n2535 0.120292
R10921 VSS.n2536 VSS.n2242 0.120292
R10922 VSS.n2540 VSS.n2242 0.120292
R10923 VSS.n2541 VSS.n2540 0.120292
R10924 VSS.n2542 VSS.n2541 0.120292
R10925 VSS.n2542 VSS.n2238 0.120292
R10926 VSS.n2546 VSS.n2238 0.120292
R10927 VSS.n2547 VSS.n2546 0.120292
R10928 VSS.n2548 VSS.n2547 0.120292
R10929 VSS.n2548 VSS.n2234 0.120292
R10930 VSS.n2553 VSS.n2234 0.120292
R10931 VSS.n2554 VSS.n2553 0.120292
R10932 VSS.n2555 VSS.n2554 0.120292
R10933 VSS.n2563 VSS.n2562 0.120292
R10934 VSS.n2563 VSS.n2225 0.120292
R10935 VSS.n2568 VSS.n2225 0.120292
R10936 VSS.n2569 VSS.n2568 0.120292
R10937 VSS.n2570 VSS.n2569 0.120292
R10938 VSS.n2570 VSS.n2223 0.120292
R10939 VSS.n2577 VSS.n2223 0.120292
R10940 VSS.n2578 VSS.n2577 0.120292
R10941 VSS.n2579 VSS.n2578 0.120292
R10942 VSS.n2579 VSS.n2220 0.120292
R10943 VSS.n2587 VSS.n2220 0.120292
R10944 VSS.n2588 VSS.n2587 0.120292
R10945 VSS.n2589 VSS.n2588 0.120292
R10946 VSS.n2589 VSS.n2217 0.120292
R10947 VSS.n2217 VSS.n2215 0.120292
R10948 VSS.n2595 VSS.n2215 0.120292
R10949 VSS.n2596 VSS.n2595 0.120292
R10950 VSS.n2596 VSS.n2212 0.120292
R10951 VSS.n2600 VSS.n2212 0.120292
R10952 VSS.n2601 VSS.n2600 0.120292
R10953 VSS.n2602 VSS.n2601 0.120292
R10954 VSS.n2602 VSS.n2209 0.120292
R10955 VSS.n2610 VSS.n2209 0.120292
R10956 VSS.n2611 VSS.n2610 0.120292
R10957 VSS.n2612 VSS.n2611 0.120292
R10958 VSS.n2612 VSS.n2206 0.120292
R10959 VSS.n2616 VSS.n2206 0.120292
R10960 VSS.n2617 VSS.n2616 0.120292
R10961 VSS.n2617 VSS.n2202 0.120292
R10962 VSS.n2624 VSS.n2202 0.120292
R10963 VSS.n2625 VSS.n2624 0.120292
R10964 VSS.n2626 VSS.n2625 0.120292
R10965 VSS.n2634 VSS.n2633 0.120292
R10966 VSS.n2634 VSS.n2192 0.120292
R10967 VSS.n2643 VSS.n2192 0.120292
R10968 VSS.n2644 VSS.n2643 0.120292
R10969 VSS.n2645 VSS.n2644 0.120292
R10970 VSS.n2645 VSS.n2190 0.120292
R10971 VSS.n2650 VSS.n2190 0.120292
R10972 VSS.n2651 VSS.n2650 0.120292
R10973 VSS.n2652 VSS.n2651 0.120292
R10974 VSS.n2652 VSS.n2186 0.120292
R10975 VSS.n2657 VSS.n2186 0.120292
R10976 VSS.n2658 VSS.n2657 0.120292
R10977 VSS.n2733 VSS.n2658 0.120292
R10978 VSS.n2733 VSS.n2732 0.120292
R10979 VSS.n2732 VSS.n2731 0.120292
R10980 VSS.n2731 VSS.n2661 0.120292
R10981 VSS.n2726 VSS.n2661 0.120292
R10982 VSS.n2726 VSS.n2725 0.120292
R10983 VSS.n2725 VSS.n2724 0.120292
R10984 VSS.n2724 VSS.n2664 0.120292
R10985 VSS.n2720 VSS.n2664 0.120292
R10986 VSS.n2720 VSS.n2719 0.120292
R10987 VSS.n2719 VSS.n2666 0.120292
R10988 VSS.n2672 VSS.n2666 0.120292
R10989 VSS.n2710 VSS.n2672 0.120292
R10990 VSS.n2710 VSS.n2709 0.120292
R10991 VSS.n2709 VSS.n2708 0.120292
R10992 VSS.n2708 VSS.n2673 0.120292
R10993 VSS.n2702 VSS.n2673 0.120292
R10994 VSS.n2702 VSS.n2701 0.120292
R10995 VSS.n2701 VSS.n2676 0.120292
R10996 VSS.n2695 VSS.n2676 0.120292
R10997 VSS.n2695 VSS.n2694 0.120292
R10998 VSS.n2694 VSS.n2693 0.120292
R10999 VSS.n2693 VSS.n2681 0.120292
R11000 VSS.n2689 VSS.n2681 0.120292
R11001 VSS.n2689 VSS.n2688 0.120292
R11002 VSS.n2688 VSS.n2687 0.120292
R11003 VSS.n2687 VSS.n2685 0.120292
R11004 VSS.n2685 VSS.n2183 0.120292
R11005 VSS.n2743 VSS.n2183 0.120292
R11006 VSS.n2744 VSS.n2743 0.120292
R11007 VSS.n2745 VSS.n2744 0.120292
R11008 VSS.n2745 VSS.n2181 0.120292
R11009 VSS.n2752 VSS.n2181 0.120292
R11010 VSS.n2753 VSS.n2752 0.120292
R11011 VSS.n2753 VSS.n2179 0.120292
R11012 VSS.n2757 VSS.n2179 0.120292
R11013 VSS.n2758 VSS.n2757 0.120292
R11014 VSS.n2759 VSS.n2758 0.120292
R11015 VSS.n2759 VSS.n2176 0.120292
R11016 VSS.n2766 VSS.n2176 0.120292
R11017 VSS.n2767 VSS.n2766 0.120292
R11018 VSS.n2767 VSS.n2173 0.120292
R11019 VSS.n2772 VSS.n2173 0.120292
R11020 VSS.n2773 VSS.n2772 0.120292
R11021 VSS.n2773 VSS.n2171 0.120292
R11022 VSS.n2781 VSS.n2171 0.120292
R11023 VSS.n2782 VSS.n2781 0.120292
R11024 VSS.n2783 VSS.n2782 0.120292
R11025 VSS.n2783 VSS.n2169 0.120292
R11026 VSS.n2791 VSS.n2169 0.120292
R11027 VSS.n2792 VSS.n2791 0.120292
R11028 VSS.n2793 VSS.n2792 0.120292
R11029 VSS.n2793 VSS.n2167 0.120292
R11030 VSS.n2797 VSS.n2167 0.120292
R11031 VSS.n2798 VSS.n2797 0.120292
R11032 VSS.n2799 VSS.n2798 0.120292
R11033 VSS.n2801 VSS.n2799 0.120292
R11034 VSS.n2831 VSS.n2801 0.120292
R11035 VSS.n2831 VSS.n2830 0.120292
R11036 VSS.n2830 VSS.n2829 0.120292
R11037 VSS.n2829 VSS.n2804 0.120292
R11038 VSS.n2823 VSS.n2804 0.120292
R11039 VSS.n2823 VSS.n2822 0.120292
R11040 VSS.n2822 VSS.n2821 0.120292
R11041 VSS.n2821 VSS.n2809 0.120292
R11042 VSS.n2817 VSS.n2809 0.120292
R11043 VSS.n2817 VSS.n2816 0.120292
R11044 VSS.n2816 VSS.n2815 0.120292
R11045 VSS.n2925 VSS.n2924 0.120292
R11046 VSS.n2924 VSS.n2156 0.120292
R11047 VSS.n2919 VSS.n2156 0.120292
R11048 VSS.n2919 VSS.n2918 0.120292
R11049 VSS.n2918 VSS.n2917 0.120292
R11050 VSS.n2917 VSS.n2159 0.120292
R11051 VSS.n2913 VSS.n2159 0.120292
R11052 VSS.n2913 VSS.n2912 0.120292
R11053 VSS.n2912 VSS.n2161 0.120292
R11054 VSS.n2899 VSS.n2837 0.120292
R11055 VSS.n2894 VSS.n2837 0.120292
R11056 VSS.n2894 VSS.n2893 0.120292
R11057 VSS.n2893 VSS.n2840 0.120292
R11058 VSS.n2844 VSS.n2840 0.120292
R11059 VSS.n2884 VSS.n2844 0.120292
R11060 VSS.n2884 VSS.n2883 0.120292
R11061 VSS.n2883 VSS.n2845 0.120292
R11062 VSS.n2879 VSS.n2845 0.120292
R11063 VSS.n2879 VSS.n2878 0.120292
R11064 VSS.n2878 VSS.n2877 0.120292
R11065 VSS.n2877 VSS.n2849 0.120292
R11066 VSS.n2873 VSS.n2849 0.120292
R11067 VSS.n2873 VSS.n2872 0.120292
R11068 VSS.n2872 VSS.n2871 0.120292
R11069 VSS.n2871 VSS.n2851 0.120292
R11070 VSS.n2865 VSS.n2851 0.120292
R11071 VSS.n2865 VSS.n2864 0.120292
R11072 VSS.n2864 VSS.n2863 0.120292
R11073 VSS.n2863 VSS.n2853 0.120292
R11074 VSS.n1565 VSS.n1558 0.120292
R11075 VSS.n1558 VSS.n1556 0.120292
R11076 VSS.n1571 VSS.n1556 0.120292
R11077 VSS.n1572 VSS.n1571 0.120292
R11078 VSS.n1572 VSS.n1553 0.120292
R11079 VSS.n1577 VSS.n1553 0.120292
R11080 VSS.n1578 VSS.n1577 0.120292
R11081 VSS.n1578 VSS.n1550 0.120292
R11082 VSS.n1583 VSS.n1550 0.120292
R11083 VSS.n1584 VSS.n1583 0.120292
R11084 VSS.n1585 VSS.n1584 0.120292
R11085 VSS.n1585 VSS.n1547 0.120292
R11086 VSS.n1547 VSS.n1546 0.120292
R11087 VSS.n1546 VSS.n1545 0.120292
R11088 VSS.n1545 VSS.n1544 0.120292
R11089 VSS.n1595 VSS.n1544 0.120292
R11090 VSS.n1596 VSS.n1595 0.120292
R11091 VSS.n1597 VSS.n1596 0.120292
R11092 VSS.n1597 VSS.n1542 0.120292
R11093 VSS.n1603 VSS.n1542 0.120292
R11094 VSS.n1604 VSS.n1603 0.120292
R11095 VSS.n1604 VSS.n1540 0.120292
R11096 VSS.n1610 VSS.n1540 0.120292
R11097 VSS.n1611 VSS.n1610 0.120292
R11098 VSS.n1613 VSS.n1611 0.120292
R11099 VSS.n1536 VSS.n1533 0.120292
R11100 VSS.n1622 VSS.n1533 0.120292
R11101 VSS.n1623 VSS.n1622 0.120292
R11102 VSS.n1624 VSS.n1623 0.120292
R11103 VSS.n1624 VSS.n1531 0.120292
R11104 VSS.n1633 VSS.n1531 0.120292
R11105 VSS.n1634 VSS.n1633 0.120292
R11106 VSS.n1635 VSS.n1634 0.120292
R11107 VSS.n1635 VSS.n1529 0.120292
R11108 VSS.n1646 VSS.n1529 0.120292
R11109 VSS.n1647 VSS.n1646 0.120292
R11110 VSS.n1648 VSS.n1647 0.120292
R11111 VSS.n1648 VSS.n1526 0.120292
R11112 VSS.n1526 VSS.n1525 0.120292
R11113 VSS.n1654 VSS.n1525 0.120292
R11114 VSS.n1655 VSS.n1654 0.120292
R11115 VSS.n1655 VSS.n1521 0.120292
R11116 VSS.n1659 VSS.n1521 0.120292
R11117 VSS.n1660 VSS.n1659 0.120292
R11118 VSS.n1661 VSS.n1660 0.120292
R11119 VSS.n1661 VSS.n1518 0.120292
R11120 VSS.n1667 VSS.n1518 0.120292
R11121 VSS.n1668 VSS.n1667 0.120292
R11122 VSS.n1669 VSS.n1668 0.120292
R11123 VSS.n1669 VSS.n1515 0.120292
R11124 VSS.n1675 VSS.n1515 0.120292
R11125 VSS.n1676 VSS.n1675 0.120292
R11126 VSS.n1677 VSS.n1676 0.120292
R11127 VSS.n1677 VSS.n1512 0.120292
R11128 VSS.n1682 VSS.n1512 0.120292
R11129 VSS.n1683 VSS.n1682 0.120292
R11130 VSS.n1683 VSS.n1508 0.120292
R11131 VSS.n1689 VSS.n1508 0.120292
R11132 VSS.n1690 VSS.n1689 0.120292
R11133 VSS.n1691 VSS.n1690 0.120292
R11134 VSS.n1691 VSS.n1505 0.120292
R11135 VSS.n1505 VSS.n1504 0.120292
R11136 VSS.n1700 VSS.n1504 0.120292
R11137 VSS.n1701 VSS.n1700 0.120292
R11138 VSS.n1701 VSS.n1501 0.120292
R11139 VSS.n1707 VSS.n1501 0.120292
R11140 VSS.n1708 VSS.n1707 0.120292
R11141 VSS.n1709 VSS.n1708 0.120292
R11142 VSS.n1709 VSS.n1498 0.120292
R11143 VSS.n1716 VSS.n1498 0.120292
R11144 VSS.n1717 VSS.n1716 0.120292
R11145 VSS.n1718 VSS.n1717 0.120292
R11146 VSS.n1718 VSS.n1496 0.120292
R11147 VSS.n1724 VSS.n1496 0.120292
R11148 VSS.n1725 VSS.n1724 0.120292
R11149 VSS.n1726 VSS.n1725 0.120292
R11150 VSS.n1726 VSS.n1494 0.120292
R11151 VSS.n1730 VSS.n1494 0.120292
R11152 VSS.n1731 VSS.n1730 0.120292
R11153 VSS.n1732 VSS.n1731 0.120292
R11154 VSS.n1732 VSS.n1491 0.120292
R11155 VSS.n1738 VSS.n1491 0.120292
R11156 VSS.n1739 VSS.n1738 0.120292
R11157 VSS.n1740 VSS.n1739 0.120292
R11158 VSS.n1740 VSS.n1487 0.120292
R11159 VSS.n1748 VSS.n1487 0.120292
R11160 VSS.n1749 VSS.n1748 0.120292
R11161 VSS.n1750 VSS.n1749 0.120292
R11162 VSS.n1750 VSS.n1485 0.120292
R11163 VSS.n1754 VSS.n1485 0.120292
R11164 VSS.n1755 VSS.n1754 0.120292
R11165 VSS.n1755 VSS.n1482 0.120292
R11166 VSS.n1482 VSS.n1480 0.120292
R11167 VSS.n1761 VSS.n1480 0.120292
R11168 VSS.n1762 VSS.n1761 0.120292
R11169 VSS.n1763 VSS.n1762 0.120292
R11170 VSS.n1763 VSS.n1477 0.120292
R11171 VSS.n1768 VSS.n1477 0.120292
R11172 VSS.n1769 VSS.n1768 0.120292
R11173 VSS.n1769 VSS.n1474 0.120292
R11174 VSS.n1474 VSS.n1473 0.120292
R11175 VSS.n1775 VSS.n1473 0.120292
R11176 VSS.n1776 VSS.n1775 0.120292
R11177 VSS.n1776 VSS.n1469 0.120292
R11178 VSS.n1781 VSS.n1469 0.120292
R11179 VSS.n1782 VSS.n1781 0.120292
R11180 VSS.n1782 VSS.n1467 0.120292
R11181 VSS.n1786 VSS.n1467 0.120292
R11182 VSS.n1787 VSS.n1786 0.120292
R11183 VSS.n1788 VSS.n1787 0.120292
R11184 VSS.n1788 VSS.n1463 0.120292
R11185 VSS.n1463 VSS.n1461 0.120292
R11186 VSS.n1793 VSS.n1461 0.120292
R11187 VSS.n1794 VSS.n1793 0.120292
R11188 VSS.n1794 VSS.n1458 0.120292
R11189 VSS.n1799 VSS.n1458 0.120292
R11190 VSS.n1800 VSS.n1799 0.120292
R11191 VSS.n1800 VSS.n1455 0.120292
R11192 VSS.n1805 VSS.n1455 0.120292
R11193 VSS.n1806 VSS.n1805 0.120292
R11194 VSS.n1807 VSS.n1806 0.120292
R11195 VSS.n1807 VSS.n1451 0.120292
R11196 VSS.n1813 VSS.n1451 0.120292
R11197 VSS.n1814 VSS.n1813 0.120292
R11198 VSS.n1815 VSS.n1814 0.120292
R11199 VSS.n1815 VSS.n1448 0.120292
R11200 VSS.n1820 VSS.n1448 0.120292
R11201 VSS.n1821 VSS.n1820 0.120292
R11202 VSS.n1821 VSS.n1445 0.120292
R11203 VSS.n1825 VSS.n1445 0.120292
R11204 VSS.n1826 VSS.n1825 0.120292
R11205 VSS.n1827 VSS.n1826 0.120292
R11206 VSS.n1827 VSS.n1443 0.120292
R11207 VSS.n1831 VSS.n1443 0.120292
R11208 VSS.n1832 VSS.n1831 0.120292
R11209 VSS.n1833 VSS.n1832 0.120292
R11210 VSS.n1833 VSS.n1440 0.120292
R11211 VSS.n1839 VSS.n1440 0.120292
R11212 VSS.n1840 VSS.n1839 0.120292
R11213 VSS.n1841 VSS.n1840 0.120292
R11214 VSS.n1841 VSS.n1437 0.120292
R11215 VSS.n1437 VSS.n1435 0.120292
R11216 VSS.n1846 VSS.n1435 0.120292
R11217 VSS.n1847 VSS.n1846 0.120292
R11218 VSS.n1848 VSS.n1847 0.120292
R11219 VSS.n1848 VSS.n1431 0.120292
R11220 VSS.n1854 VSS.n1431 0.120292
R11221 VSS.n1855 VSS.n1854 0.120292
R11222 VSS.n1855 VSS.n1428 0.120292
R11223 VSS.n1860 VSS.n1428 0.120292
R11224 VSS.n1861 VSS.n1860 0.120292
R11225 VSS.n1861 VSS.n1426 0.120292
R11226 VSS.n1866 VSS.n1426 0.120292
R11227 VSS.n1867 VSS.n1866 0.120292
R11228 VSS.n1874 VSS.n1873 0.120292
R11229 VSS.n1874 VSS.n1419 0.120292
R11230 VSS.n1419 VSS.n1418 0.120292
R11231 VSS.n1879 VSS.n1418 0.120292
R11232 VSS.n1880 VSS.n1879 0.120292
R11233 VSS.n1881 VSS.n1880 0.120292
R11234 VSS.n1881 VSS.n1416 0.120292
R11235 VSS.n1416 VSS.n1414 0.120292
R11236 VSS.n1414 VSS.n1413 0.120292
R11237 VSS.n1413 VSS.n1410 0.120292
R11238 VSS.n1888 VSS.n1410 0.120292
R11239 VSS.n1889 VSS.n1888 0.120292
R11240 VSS.n1889 VSS.n1408 0.120292
R11241 VSS.n1897 VSS.n1408 0.120292
R11242 VSS.n1898 VSS.n1897 0.120292
R11243 VSS.n1899 VSS.n1898 0.120292
R11244 VSS.n1899 VSS.n1404 0.120292
R11245 VSS.n1905 VSS.n1404 0.120292
R11246 VSS.n1906 VSS.n1905 0.120292
R11247 VSS.n1907 VSS.n1906 0.120292
R11248 VSS.n1907 VSS.n1401 0.120292
R11249 VSS.n1913 VSS.n1401 0.120292
R11250 VSS.n1914 VSS.n1913 0.120292
R11251 VSS.n1915 VSS.n1914 0.120292
R11252 VSS.n1915 VSS.n1396 0.120292
R11253 VSS.n1923 VSS.n1396 0.120292
R11254 VSS.n1924 VSS.n1923 0.120292
R11255 VSS.n1924 VSS.n1394 0.120292
R11256 VSS.n1928 VSS.n1394 0.120292
R11257 VSS.n1929 VSS.n1928 0.120292
R11258 VSS.n1930 VSS.n1929 0.120292
R11259 VSS.n1930 VSS.n1392 0.120292
R11260 VSS.n1935 VSS.n1392 0.120292
R11261 VSS.n1936 VSS.n1935 0.120292
R11262 VSS.n1936 VSS.n1388 0.120292
R11263 VSS.n1940 VSS.n1388 0.120292
R11264 VSS.n1941 VSS.n1940 0.120292
R11265 VSS.n1942 VSS.n1941 0.120292
R11266 VSS.n1942 VSS.n1384 0.120292
R11267 VSS.n1948 VSS.n1384 0.120292
R11268 VSS.n1949 VSS.n1948 0.120292
R11269 VSS.n1950 VSS.n1949 0.120292
R11270 VSS.n1950 VSS.n1380 0.120292
R11271 VSS.n1956 VSS.n1380 0.120292
R11272 VSS.n1957 VSS.n1956 0.120292
R11273 VSS.n1957 VSS.n1378 0.120292
R11274 VSS.n1963 VSS.n1378 0.120292
R11275 VSS.n1964 VSS.n1963 0.120292
R11276 VSS.n1965 VSS.n1964 0.120292
R11277 VSS.n1965 VSS.n1376 0.120292
R11278 VSS.n1376 VSS.n1375 0.120292
R11279 VSS.n1974 VSS.n1375 0.120292
R11280 VSS.n1975 VSS.n1974 0.120292
R11281 VSS.n1976 VSS.n1975 0.120292
R11282 VSS.n1976 VSS.n1372 0.120292
R11283 VSS.n1980 VSS.n1372 0.120292
R11284 VSS.n1981 VSS.n1980 0.120292
R11285 VSS.n1982 VSS.n1981 0.120292
R11286 VSS.n1982 VSS.n1370 0.120292
R11287 VSS.n1370 VSS.n1369 0.120292
R11288 VSS.n1369 VSS.n1368 0.120292
R11289 VSS.n1368 VSS.n1365 0.120292
R11290 VSS.n1994 VSS.n1365 0.120292
R11291 VSS.n1995 VSS.n1994 0.120292
R11292 VSS.n1996 VSS.n1995 0.120292
R11293 VSS.n1996 VSS.n1362 0.120292
R11294 VSS.n1362 VSS.n1360 0.120292
R11295 VSS.n1360 VSS.n1359 0.120292
R11296 VSS.n2004 VSS.n1359 0.120292
R11297 VSS.n2005 VSS.n2004 0.120292
R11298 VSS.n2005 VSS.n1354 0.120292
R11299 VSS.n2011 VSS.n1354 0.120292
R11300 VSS.n2012 VSS.n2011 0.120292
R11301 VSS.n2012 VSS.n1351 0.120292
R11302 VSS.n2017 VSS.n1351 0.120292
R11303 VSS.n2018 VSS.n2017 0.120292
R11304 VSS.n2018 VSS.n1348 0.120292
R11305 VSS.n2022 VSS.n1348 0.120292
R11306 VSS.n2023 VSS.n2022 0.120292
R11307 VSS.n2044 VSS.n2043 0.120292
R11308 VSS.n2044 VSS.n1338 0.120292
R11309 VSS.n2050 VSS.n1338 0.120292
R11310 VSS.n2051 VSS.n2050 0.120292
R11311 VSS.n2051 VSS.n1335 0.120292
R11312 VSS.n2055 VSS.n1335 0.120292
R11313 VSS.n2056 VSS.n2055 0.120292
R11314 VSS.n2057 VSS.n2056 0.120292
R11315 VSS.n2057 VSS.n1333 0.120292
R11316 VSS.n2064 VSS.n1333 0.120292
R11317 VSS.n2065 VSS.n2064 0.120292
R11318 VSS.n2065 VSS.n1330 0.120292
R11319 VSS.n1330 VSS.n1329 0.120292
R11320 VSS.n1329 VSS.n1328 0.120292
R11321 VSS.n1328 VSS.n1262 0.120292
R11322 VSS.n1322 VSS.n1262 0.120292
R11323 VSS.n1322 VSS.n1321 0.120292
R11324 VSS.n1321 VSS.n1320 0.120292
R11325 VSS.n1320 VSS.n1264 0.120292
R11326 VSS.n1315 VSS.n1264 0.120292
R11327 VSS.n1315 VSS.n1314 0.120292
R11328 VSS.n1314 VSS.n1266 0.120292
R11329 VSS.n1308 VSS.n1266 0.120292
R11330 VSS.n1308 VSS.n1307 0.120292
R11331 VSS.n1307 VSS.n1268 0.120292
R11332 VSS.n1301 VSS.n1268 0.120292
R11333 VSS.n1301 VSS.n1300 0.120292
R11334 VSS.n1300 VSS.n1299 0.120292
R11335 VSS.n1299 VSS.n1271 0.120292
R11336 VSS.n1293 VSS.n1271 0.120292
R11337 VSS.n1293 VSS.n1292 0.120292
R11338 VSS.n1292 VSS.n1291 0.120292
R11339 VSS.n1291 VSS.n1275 0.120292
R11340 VSS.n1287 VSS.n1275 0.120292
R11341 VSS.n1287 VSS.n1286 0.120292
R11342 VSS.n1286 VSS.n1285 0.120292
R11343 VSS.n5336 VSS.n5330 0.120292
R11344 VSS.n5337 VSS.n5336 0.120292
R11345 VSS.n5338 VSS.n5337 0.120292
R11346 VSS.n5338 VSS.n5328 0.120292
R11347 VSS.n5328 VSS.n5325 0.120292
R11348 VSS.n5343 VSS.n5325 0.120292
R11349 VSS.n5344 VSS.n5343 0.120292
R11350 VSS.n5345 VSS.n5344 0.120292
R11351 VSS.n5345 VSS.n5323 0.120292
R11352 VSS.n5323 VSS.n5322 0.120292
R11353 VSS.n5322 VSS.n5321 0.120292
R11354 VSS.n5321 VSS.n179 0.120292
R11355 VSS.n5316 VSS.n179 0.120292
R11356 VSS.n5316 VSS.n5315 0.120292
R11357 VSS.n5315 VSS.n5314 0.120292
R11358 VSS.n5314 VSS.n181 0.120292
R11359 VSS.n5309 VSS.n181 0.120292
R11360 VSS.n5309 VSS.n5308 0.120292
R11361 VSS.n5308 VSS.n5307 0.120292
R11362 VSS.n5307 VSS.n183 0.120292
R11363 VSS.n5303 VSS.n183 0.120292
R11364 VSS.n5303 VSS.n5302 0.120292
R11365 VSS.n5302 VSS.n5301 0.120292
R11366 VSS.n5301 VSS.n186 0.120292
R11367 VSS.n5297 VSS.n186 0.120292
R11368 VSS.n5297 VSS.n5296 0.120292
R11369 VSS.n5296 VSS.n5295 0.120292
R11370 VSS.n5295 VSS.n189 0.120292
R11371 VSS.n5288 VSS.n189 0.120292
R11372 VSS.n5288 VSS.n5287 0.120292
R11373 VSS.n5287 VSS.n5286 0.120292
R11374 VSS.n5286 VSS.n191 0.120292
R11375 VSS.n5281 VSS.n191 0.120292
R11376 VSS.n5281 VSS.n5280 0.120292
R11377 VSS.n5280 VSS.n5279 0.120292
R11378 VSS.n5279 VSS.n193 0.120292
R11379 VSS.n5273 VSS.n193 0.120292
R11380 VSS.n5273 VSS.n5272 0.120292
R11381 VSS.n5272 VSS.n5271 0.120292
R11382 VSS.n5271 VSS.n197 0.120292
R11383 VSS.n5267 VSS.n197 0.120292
R11384 VSS.n5267 VSS.n5266 0.120292
R11385 VSS.n5266 VSS.n5265 0.120292
R11386 VSS.n5265 VSS.n200 0.120292
R11387 VSS.n5261 VSS.n200 0.120292
R11388 VSS.n5261 VSS.n5260 0.120292
R11389 VSS.n5260 VSS.n5259 0.120292
R11390 VSS.n5259 VSS.n203 0.120292
R11391 VSS.n5253 VSS.n203 0.120292
R11392 VSS.n5253 VSS.n5252 0.120292
R11393 VSS.n5252 VSS.n5251 0.120292
R11394 VSS.n5251 VSS.n205 0.120292
R11395 VSS.n5247 VSS.n205 0.120292
R11396 VSS.n5247 VSS.n5246 0.120292
R11397 VSS.n5246 VSS.n5245 0.120292
R11398 VSS.n5245 VSS.n207 0.120292
R11399 VSS.n5241 VSS.n207 0.120292
R11400 VSS.n5241 VSS.n5240 0.120292
R11401 VSS.n5240 VSS.n209 0.120292
R11402 VSS.n5234 VSS.n209 0.120292
R11403 VSS.n5234 VSS.n5233 0.120292
R11404 VSS.n5233 VSS.n5232 0.120292
R11405 VSS.n5232 VSS.n211 0.120292
R11406 VSS.n5227 VSS.n211 0.120292
R11407 VSS.n5227 VSS.n5226 0.120292
R11408 VSS.n5226 VSS.n5225 0.120292
R11409 VSS.n5225 VSS.n213 0.120292
R11410 VSS.n5220 VSS.n213 0.120292
R11411 VSS.n5220 VSS.n5219 0.120292
R11412 VSS.n5219 VSS.n215 0.120292
R11413 VSS.n5215 VSS.n215 0.120292
R11414 VSS.n5215 VSS.n5214 0.120292
R11415 VSS.n5214 VSS.n5213 0.120292
R11416 VSS.n5213 VSS.n219 0.120292
R11417 VSS.n5209 VSS.n219 0.120292
R11418 VSS.n5209 VSS.n5208 0.120292
R11419 VSS.n5208 VSS.n5207 0.120292
R11420 VSS.n5207 VSS.n221 0.120292
R11421 VSS.n5202 VSS.n221 0.120292
R11422 VSS.n5202 VSS.n5201 0.120292
R11423 VSS.n5201 VSS.n223 0.120292
R11424 VSS.n5197 VSS.n223 0.120292
R11425 VSS.n5197 VSS.n5196 0.120292
R11426 VSS.n5196 VSS.n5195 0.120292
R11427 VSS.n5195 VSS.n227 0.120292
R11428 VSS.n5190 VSS.n227 0.120292
R11429 VSS.n5190 VSS.n5189 0.120292
R11430 VSS.n5189 VSS.n5188 0.120292
R11431 VSS.n5188 VSS.n229 0.120292
R11432 VSS.n5184 VSS.n229 0.120292
R11433 VSS.n5184 VSS.n5183 0.120292
R11434 VSS.n5183 VSS.n5182 0.120292
R11435 VSS.n5182 VSS.n234 0.120292
R11436 VSS.n5139 VSS.n234 0.120292
R11437 VSS.n5140 VSS.n5139 0.120292
R11438 VSS.n5140 VSS.n5138 0.120292
R11439 VSS.n5147 VSS.n5138 0.120292
R11440 VSS.n5149 VSS.n5136 0.120292
R11441 VSS.n5136 VSS.n5134 0.120292
R11442 VSS.n5154 VSS.n5134 0.120292
R11443 VSS.n5155 VSS.n5154 0.120292
R11444 VSS.n5155 VSS.n5131 0.120292
R11445 VSS.n5162 VSS.n5161 0.120292
R11446 VSS.n5162 VSS.n5128 0.120292
R11447 VSS.n5166 VSS.n5128 0.120292
R11448 VSS.n5167 VSS.n5166 0.120292
R11449 VSS.n5168 VSS.n5167 0.120292
R11450 VSS.n5168 VSS.n5126 0.120292
R11451 VSS.n5126 VSS.n5125 0.120292
R11452 VSS.n5173 VSS.n5125 0.120292
R11453 VSS.n5174 VSS.n5173 0.120292
R11454 VSS.n5175 VSS.n5174 0.120292
R11455 VSS.n5175 VSS.n5122 0.120292
R11456 VSS.n5122 VSS.n5121 0.120292
R11457 VSS.n5121 VSS.n5120 0.120292
R11458 VSS.n5120 VSS.n237 0.120292
R11459 VSS.n5115 VSS.n237 0.120292
R11460 VSS.n5115 VSS.n5114 0.120292
R11461 VSS.n5114 VSS.n239 0.120292
R11462 VSS.n5110 VSS.n239 0.120292
R11463 VSS.n5110 VSS.n5109 0.120292
R11464 VSS.n5109 VSS.n5108 0.120292
R11465 VSS.n5108 VSS.n243 0.120292
R11466 VSS.n5104 VSS.n243 0.120292
R11467 VSS.n5104 VSS.n5103 0.120292
R11468 VSS.n5103 VSS.n5102 0.120292
R11469 VSS.n5102 VSS.n246 0.120292
R11470 VSS.n5098 VSS.n246 0.120292
R11471 VSS.n5098 VSS.n5097 0.120292
R11472 VSS.n5097 VSS.n5096 0.120292
R11473 VSS.n5096 VSS.n248 0.120292
R11474 VSS.n5092 VSS.n248 0.120292
R11475 VSS.n5092 VSS.n5091 0.120292
R11476 VSS.n5091 VSS.n5090 0.120292
R11477 VSS.n5090 VSS.n251 0.120292
R11478 VSS.n5086 VSS.n251 0.120292
R11479 VSS.n5086 VSS.n5085 0.120292
R11480 VSS.n5085 VSS.n5084 0.120292
R11481 VSS.n5084 VSS.n253 0.120292
R11482 VSS.n5080 VSS.n253 0.120292
R11483 VSS.n5080 VSS.n5079 0.120292
R11484 VSS.n5079 VSS.n5078 0.120292
R11485 VSS.n5078 VSS.n255 0.120292
R11486 VSS.n5074 VSS.n255 0.120292
R11487 VSS.n5074 VSS.n5073 0.120292
R11488 VSS.n5073 VSS.n5072 0.120292
R11489 VSS.n5072 VSS.n258 0.120292
R11490 VSS.n5067 VSS.n258 0.120292
R11491 VSS.n5067 VSS.n5066 0.120292
R11492 VSS.n5064 VSS.n263 0.120292
R11493 VSS.n5059 VSS.n263 0.120292
R11494 VSS.n5059 VSS.n5058 0.120292
R11495 VSS.n5058 VSS.n5057 0.120292
R11496 VSS.n5057 VSS.n265 0.120292
R11497 VSS.n5051 VSS.n5050 0.120292
R11498 VSS.n5050 VSS.n269 0.120292
R11499 VSS.n5045 VSS.n269 0.120292
R11500 VSS.n5045 VSS.n5044 0.120292
R11501 VSS.n5044 VSS.n5043 0.120292
R11502 VSS.n5043 VSS.n271 0.120292
R11503 VSS.n5037 VSS.n271 0.120292
R11504 VSS.n5037 VSS.n5036 0.120292
R11505 VSS.n5036 VSS.n5035 0.120292
R11506 VSS.n5035 VSS.n275 0.120292
R11507 VSS.n5029 VSS.n275 0.120292
R11508 VSS.n5029 VSS.n5028 0.120292
R11509 VSS.n5028 VSS.n5027 0.120292
R11510 VSS.n5027 VSS.n279 0.120292
R11511 VSS.n5022 VSS.n279 0.120292
R11512 VSS.n5022 VSS.n5021 0.120292
R11513 VSS.n5019 VSS.n284 0.120292
R11514 VSS.n5015 VSS.n284 0.120292
R11515 VSS.n5015 VSS.n5014 0.120292
R11516 VSS.n5014 VSS.n5013 0.120292
R11517 VSS.n5013 VSS.n287 0.120292
R11518 VSS.n5008 VSS.n287 0.120292
R11519 VSS.n5008 VSS.n5007 0.120292
R11520 VSS.n5005 VSS.n292 0.120292
R11521 VSS.n5000 VSS.n292 0.120292
R11522 VSS.n5000 VSS.n4999 0.120292
R11523 VSS.n4999 VSS.n4998 0.120292
R11524 VSS.n4998 VSS.n294 0.120292
R11525 VSS.n4898 VSS.n294 0.120292
R11526 VSS.n4899 VSS.n4898 0.120292
R11527 VSS.n4900 VSS.n4899 0.120292
R11528 VSS.n4900 VSS.n4894 0.120292
R11529 VSS.n4894 VSS.n4892 0.120292
R11530 VSS.n4905 VSS.n4892 0.120292
R11531 VSS.n4906 VSS.n4905 0.120292
R11532 VSS.n4907 VSS.n4906 0.120292
R11533 VSS.n4907 VSS.n4890 0.120292
R11534 VSS.n4890 VSS.n4889 0.120292
R11535 VSS.n4912 VSS.n4889 0.120292
R11536 VSS.n4913 VSS.n4912 0.120292
R11537 VSS.n4914 VSS.n4913 0.120292
R11538 VSS.n4914 VSS.n4887 0.120292
R11539 VSS.n4887 VSS.n4886 0.120292
R11540 VSS.n4919 VSS.n4886 0.120292
R11541 VSS.n4920 VSS.n4919 0.120292
R11542 VSS.n4921 VSS.n4920 0.120292
R11543 VSS.n4921 VSS.n4883 0.120292
R11544 VSS.n4925 VSS.n4883 0.120292
R11545 VSS.n4926 VSS.n4925 0.120292
R11546 VSS.n4927 VSS.n4926 0.120292
R11547 VSS.n4927 VSS.n4881 0.120292
R11548 VSS.n4931 VSS.n4881 0.120292
R11549 VSS.n4932 VSS.n4931 0.120292
R11550 VSS.n4933 VSS.n4932 0.120292
R11551 VSS.n4933 VSS.n4878 0.120292
R11552 VSS.n4878 VSS.n4877 0.120292
R11553 VSS.n4877 VSS.n4876 0.120292
R11554 VSS.n4876 VSS.n371 0.120292
R11555 VSS.n4870 VSS.n371 0.120292
R11556 VSS.n4870 VSS.n4869 0.120292
R11557 VSS.n4869 VSS.n4868 0.120292
R11558 VSS.n4868 VSS.n374 0.120292
R11559 VSS.n4863 VSS.n374 0.120292
R11560 VSS.n4863 VSS.n4862 0.120292
R11561 VSS.n4862 VSS.n4861 0.120292
R11562 VSS.n4861 VSS.n376 0.120292
R11563 VSS.n4856 VSS.n376 0.120292
R11564 VSS.n4848 VSS.n386 0.120292
R11565 VSS.n4832 VSS.n386 0.120292
R11566 VSS.n4832 VSS.n4831 0.120292
R11567 VSS.n4831 VSS.n4830 0.120292
R11568 VSS.n4830 VSS.n389 0.120292
R11569 VSS.n4826 VSS.n389 0.120292
R11570 VSS.n4826 VSS.n4825 0.120292
R11571 VSS.n4825 VSS.n391 0.120292
R11572 VSS.n4819 VSS.n391 0.120292
R11573 VSS.n4819 VSS.n4818 0.120292
R11574 VSS.n4818 VSS.n4817 0.120292
R11575 VSS.n4817 VSS.n394 0.120292
R11576 VSS.n459 VSS.n394 0.120292
R11577 VSS.n459 VSS.n458 0.120292
R11578 VSS.n458 VSS.n396 0.120292
R11579 VSS.n452 VSS.n396 0.120292
R11580 VSS.n452 VSS.n451 0.120292
R11581 VSS.n451 VSS.n450 0.120292
R11582 VSS.n450 VSS.n398 0.120292
R11583 VSS.n446 VSS.n398 0.120292
R11584 VSS.n446 VSS.n445 0.120292
R11585 VSS.n445 VSS.n444 0.120292
R11586 VSS.n444 VSS.n402 0.120292
R11587 VSS.n440 VSS.n402 0.120292
R11588 VSS.n440 VSS.n439 0.120292
R11589 VSS.n439 VSS.n438 0.120292
R11590 VSS.n438 VSS.n405 0.120292
R11591 VSS.n434 VSS.n405 0.120292
R11592 VSS.n434 VSS.n433 0.120292
R11593 VSS.n433 VSS.n432 0.120292
R11594 VSS.n432 VSS.n408 0.120292
R11595 VSS.n428 VSS.n408 0.120292
R11596 VSS.n428 VSS.n427 0.120292
R11597 VSS.n427 VSS.n426 0.120292
R11598 VSS.n426 VSS.n411 0.120292
R11599 VSS.n422 VSS.n411 0.120292
R11600 VSS.n422 VSS.n421 0.120292
R11601 VSS.n421 VSS.n420 0.120292
R11602 VSS.n420 VSS.n414 0.120292
R11603 VSS.n4600 VSS.n469 0.120292
R11604 VSS.n4601 VSS.n4600 0.120292
R11605 VSS.n4602 VSS.n4601 0.120292
R11606 VSS.n1219 VSS.n1218 0.120292
R11607 VSS.n1218 VSS.n1217 0.120292
R11608 VSS.n1217 VSS.n986 0.120292
R11609 VSS.n1175 VSS.n1174 0.117037
R11610 VSS.n4805 VSS.n4804 0.116225
R11611 VSS.n338 VSS.n326 0.108833
R11612 VSS.n634 VSS.n617 0.104667
R11613 VSS.n4674 VSS.n634 0.104667
R11614 VSS.n548 VSS.n546 0.104667
R11615 VSS.n615 VSS.n546 0.104667
R11616 VSS.n912 VSS.n769 0.104667
R11617 VSS.n910 VSS.n769 0.104667
R11618 VSS.n856 VSS.n788 0.104667
R11619 VSS.n856 VSS.n855 0.104667
R11620 VSS VSS.n5777 0.0972906
R11621 VSS.n4745 VSS.n4744 0.0966538
R11622 VSS.n544 VSS.n494 0.0966538
R11623 VSS.n5775 VSS.n5774 0.0950946
R11624 VSS.n5768 VSS.n7 0.0950946
R11625 VSS.n4380 VSS.n4378 0.0950946
R11626 VSS.n4398 VSS.n3700 0.0950946
R11627 VSS.n3657 VSS.n3656 0.0950946
R11628 VSS.n3662 VSS.n3661 0.0950946
R11629 VSS.n2937 VSS.n2936 0.0950946
R11630 VSS.n2930 VSS.n2152 0.0950946
R11631 VSS.n2026 VSS.n2024 0.0950946
R11632 VSS.n2041 VSS.n1341 0.0950946
R11633 VSS.n4854 VSS.n380 0.0950946
R11634 VSS.n4850 VSS.n384 0.0950946
R11635 VSS.n4565 VSS.n8 0.0916458
R11636 VSS.n4400 VSS.n4399 0.0916458
R11637 VSS.n3670 VSS.n2139 0.0916458
R11638 VSS.n2925 VSS.n2153 0.0916458
R11639 VSS.n2043 VSS.n2042 0.0916458
R11640 VSS.n4849 VSS.n4848 0.0916458
R11641 VSS.n2581 VSS.n2580 0.0900105
R11642 VSS.n2765 VSS.n2764 0.0900105
R11643 VSS.n1593 VSS.n1592 0.0900105
R11644 VSS.n1146 VSS.n1145 0.0882358
R11645 VSS.n1154 VSS.n1153 0.0882358
R11646 VSS.n941 VSS.n938 0.0882358
R11647 VSS.n940 VSS.n939 0.0882358
R11648 VSS.n3932 VSS.n3931 0.0881712
R11649 VSS.n2843 VSS.n2841 0.0881712
R11650 VSS.n2847 VSS.n2846 0.0881712
R11651 VSS.n5773 VSS.n5772 0.0838333
R11652 VSS.n4393 VSS.n3703 0.0838333
R11653 VSS.n3655 VSS.n2143 0.0838333
R11654 VSS.n2935 VSS.n2934 0.0838333
R11655 VSS.n2036 VSS.n1344 0.0838333
R11656 VSS.n4842 VSS.n4838 0.0838333
R11657 VSS.n4607 VSS.n4605 0.0812292
R11658 VSS.n985 VSS.n984 0.0812292
R11659 VSS.n3867 VSS.n3866 0.0700652
R11660 VSS.n3922 VSS.n3921 0.0685851
R11661 VSS.n3928 VSS.n3927 0.0685851
R11662 VSS.n3978 VSS.n3977 0.0685851
R11663 VSS.n4262 VSS.n4261 0.0685851
R11664 VSS.n2714 VSS.n2668 0.0685851
R11665 VSS.n2705 VSS.n2704 0.0685851
R11666 VSS.n5771 VSS.n4 0.0680676
R11667 VSS.n5771 VSS.n5770 0.0680676
R11668 VSS.n4394 VSS.n3702 0.0680676
R11669 VSS.n4395 VSS.n4394 0.0680676
R11670 VSS.n3653 VSS.n3652 0.0680676
R11671 VSS.n3652 VSS.n2144 0.0680676
R11672 VSS.n2933 VSS.n2149 0.0680676
R11673 VSS.n2933 VSS.n2932 0.0680676
R11674 VSS.n2037 VSS.n1343 0.0680676
R11675 VSS.n2038 VSS.n2037 0.0680676
R11676 VSS.n4841 VSS.n4839 0.0680676
R11677 VSS.n4841 VSS.n4840 0.0680676
R11678 VSS.n963 VSS.n958 0.0677515
R11679 VSS.n5 VSS.n3 0.0656042
R11680 VSS.n5767 VSS.n6 0.0656042
R11681 VSS.n4381 VSS.n4377 0.0656042
R11682 VSS.n4392 VSS.n3704 0.0656042
R11683 VSS.n3654 VSS.n3651 0.0656042
R11684 VSS.n3664 VSS.n3663 0.0656042
R11685 VSS.n2150 VSS.n2148 0.0656042
R11686 VSS.n2929 VSS.n2151 0.0656042
R11687 VSS.n2028 VSS.n2027 0.0656042
R11688 VSS.n2035 VSS.n1345 0.0656042
R11689 VSS.n4855 VSS.n379 0.0656042
R11690 VSS.n4844 VSS.n4843 0.0656042
R11691 VSS.n1096 VSS.n1025 0.0620894
R11692 VSS.n5769 VSS.n2 0.0574697
R11693 VSS.n4396 VSS.n3701 0.0574697
R11694 VSS.n2940 VSS.n2145 0.0574697
R11695 VSS.n2931 VSS.n2147 0.0574697
R11696 VSS.n2039 VSS.n1342 0.0574697
R11697 VSS.n383 VSS.n381 0.0574697
R11698 VSS.n5761 VSS.n3 0.0551875
R11699 VSS.n5767 VSS.n5766 0.0551875
R11700 VSS.n4382 VSS.n4381 0.0551875
R11701 VSS.n3704 VSS.n3699 0.0551875
R11702 VSS.n3651 VSS.n3650 0.0551875
R11703 VSS.n3663 VSS.n2140 0.0551875
R11704 VSS.n2815 VSS.n2148 0.0551875
R11705 VSS.n2929 VSS.n2928 0.0551875
R11706 VSS.n2027 VSS.n2023 0.0551875
R11707 VSS.n1345 VSS.n1340 0.0551875
R11708 VSS.n4856 VSS.n4855 0.0551875
R11709 VSS.n4843 VSS.n385 0.0551875
R11710 VSS.n1174 VSS.n1166 0.0550024
R11711 VSS.n4804 VSS.n471 0.0550024
R11712 VSS.n4668 VSS.n936 0.0542119
R11713 VSS.n1136 VSS.n1135 0.0515714
R11714 VSS.n4678 VSS.n4677 0.0513197
R11715 VSS.n908 VSS.n907 0.0513197
R11716 VSS.n4671 VSS.n4670 0.0477304
R11717 VSS.n1031 VSS.n1026 0.0475814
R11718 VSS.n4667 VSS.n4666 0.0469286
R11719 VSS.n1156 VSS.n1137 0.0469286
R11720 VSS.n5774 VSS.n4 0.0410405
R11721 VSS.n5770 VSS.n5768 0.0410405
R11722 VSS.n4378 VSS.n3702 0.0410405
R11723 VSS.n4395 VSS.n3700 0.0410405
R11724 VSS.n3656 VSS.n3653 0.0410405
R11725 VSS.n3662 VSS.n2144 0.0410405
R11726 VSS.n2936 VSS.n2149 0.0410405
R11727 VSS.n2932 VSS.n2930 0.0410405
R11728 VSS.n2024 VSS.n1343 0.0410405
R11729 VSS.n2038 VSS.n1341 0.0410405
R11730 VSS.n4839 VSS.n380 0.0410405
R11731 VSS.n4840 VSS.n384 0.0410405
R11732 VSS.n4605 VSS.n4602 0.0395625
R11733 VSS.n1219 VSS.n985 0.0395625
R11734 VSS.n959 VSS.n958 0.0363187
R11735 VSS.n4853 VSS.n381 0.0292489
R11736 VSS.n4851 VSS.n383 0.0292489
R11737 VSS.n2025 VSS.n1342 0.0292489
R11738 VSS.n2040 VSS.n2039 0.0292489
R11739 VSS.n2938 VSS.n2147 0.0292489
R11740 VSS.n2931 VSS.n2146 0.0292489
R11741 VSS.n3658 VSS.n2940 0.0292489
R11742 VSS.n3660 VSS.n2145 0.0292489
R11743 VSS.n4379 VSS.n3701 0.0292489
R11744 VSS.n4397 VSS.n4396 0.0292489
R11745 VSS.n5776 VSS.n2 0.0292489
R11746 VSS.n5769 VSS.n0 0.0292489
R11747 VSS.n5766 VSS.n8 0.0291458
R11748 VSS.n4399 VSS.n3699 0.0291458
R11749 VSS.n2140 VSS.n2139 0.0291458
R11750 VSS.n2928 VSS.n2153 0.0291458
R11751 VSS.n2042 VSS.n1340 0.0291458
R11752 VSS.n4849 VSS.n385 0.0291458
R11753 VSS.n4974 VSS.n348 0.0258906
R11754 VSS.n5773 VSS.n5 0.0187292
R11755 VSS.n5772 VSS.n6 0.0187292
R11756 VSS.n4377 VSS.n3703 0.0187292
R11757 VSS.n4393 VSS.n4392 0.0187292
R11758 VSS.n3655 VSS.n3654 0.0187292
R11759 VSS.n3664 VSS.n2143 0.0187292
R11760 VSS.n2935 VSS.n2150 0.0187292
R11761 VSS.n2934 VSS.n2151 0.0187292
R11762 VSS.n2028 VSS.n1344 0.0187292
R11763 VSS.n2036 VSS.n2035 0.0187292
R11764 VSS.n4838 VSS.n379 0.0187292
R11765 VSS.n4844 VSS.n4842 0.0187292
R11766 VSS.n1137 VSS.n1136 0.0172857
R11767 VSS.n4668 VSS.n4667 0.0147857
R11768 VSS.n4672 VSS.n701 0.00856395
R11769 VSS.n914 VSS.n767 0.00856395
R11770 VSS.n4975 VSS.n4974 0.00635938
R11771 VSS.n1107 VSS.t3213 0.00492008
R11772 VSS.n4630 VSS.t3469 0.00229169
R11773 VSS.n4670 VSS.n915 0.000960784
R11774 VDAC_N.n0 VDAC_N.t1522 946.489
R11775 VDAC_N.n10 VDAC_N.t1756 946.489
R11776 VDAC_N.n3 VDAC_N.t138 946.489
R11777 VDAC_N.n2 VDAC_N.t1772 945.755
R11778 VDAC_N.n1 VDAC_N.t702 945.755
R11779 VDAC_N.n0 VDAC_N.t1438 945.755
R11780 VDAC_N.n12 VDAC_N.t627 945.755
R11781 VDAC_N.n11 VDAC_N.t1791 945.755
R11782 VDAC_N.n10 VDAC_N.t925 945.755
R11783 VDAC_N.n9 VDAC_N.t284 945.755
R11784 VDAC_N.n8 VDAC_N.t1423 945.755
R11785 VDAC_N.n7 VDAC_N.t1397 945.755
R11786 VDAC_N.n6 VDAC_N.t363 945.755
R11787 VDAC_N.n5 VDAC_N.t955 945.755
R11788 VDAC_N.n4 VDAC_N.t584 945.755
R11789 VDAC_N.n3 VDAC_N.t184 945.755
R11790 VDAC_N.n22 VDAC_N.n14 20.4951
R11791 VDAC_N.n20 VDAC_N.n18 14.894
R11792 VDAC_N.n17 VDAC_N.n15 14.894
R11793 VDAC_N.n17 VDAC_N.n16 14.394
R11794 VDAC_N.n20 VDAC_N.n19 14.394
R11795 VDAC_N.n22 VDAC_N.n21 13.2477
R11796 VDAC_N.n6 VDAC_N.n5 6.84978
R11797 VDAC_N.n14 VDAC_N.n13 3.02654
R11798 VDAC_N.n14 VDAC_N.n2 2.75535
R11799 VDAC_N.n18 VDAC_N.t5 2.4755
R11800 VDAC_N.n18 VDAC_N.t4 2.4755
R11801 VDAC_N.n16 VDAC_N.t6 2.4755
R11802 VDAC_N.n16 VDAC_N.t7 2.4755
R11803 VDAC_N.n15 VDAC_N.t3 2.4755
R11804 VDAC_N.n15 VDAC_N.t2 2.4755
R11805 VDAC_N.n19 VDAC_N.t1 2.4755
R11806 VDAC_N.n19 VDAC_N.t0 2.4755
R11807 VDAC_N VDAC_N.n22 2.17582
R11808 VDAC_N.n116 VDAC_N.t2036 1.1255
R11809 VDAC_N.n117 VDAC_N.t1739 1.1255
R11810 VDAC_N.n118 VDAC_N.t164 1.1255
R11811 VDAC_N.n119 VDAC_N.t829 1.1255
R11812 VDAC_N.n120 VDAC_N.t2091 1.1255
R11813 VDAC_N.n121 VDAC_N.t808 1.1255
R11814 VDAC_N.n122 VDAC_N.t1979 1.1255
R11815 VDAC_N.n123 VDAC_N.t1152 1.1255
R11816 VDAC_N.n124 VDAC_N.t402 1.1255
R11817 VDAC_N.n125 VDAC_N.t1396 1.1255
R11818 VDAC_N.n126 VDAC_N.t1290 1.1255
R11819 VDAC_N.n127 VDAC_N.t2121 1.1255
R11820 VDAC_N.n128 VDAC_N.t552 1.1255
R11821 VDAC_N.n129 VDAC_N.t1022 1.1255
R11822 VDAC_N.n130 VDAC_N.t638 1.1255
R11823 VDAC_N.n131 VDAC_N.t295 1.1255
R11824 VDAC_N.n132 VDAC_N.t1675 1.1255
R11825 VDAC_N.n133 VDAC_N.t1970 1.1255
R11826 VDAC_N.n134 VDAC_N.t1457 1.1255
R11827 VDAC_N.n135 VDAC_N.t1025 1.1255
R11828 VDAC_N.n136 VDAC_N.t111 1.1255
R11829 VDAC_N.n137 VDAC_N.t1809 1.1255
R11830 VDAC_N.n138 VDAC_N.t633 1.1255
R11831 VDAC_N.n139 VDAC_N.t1705 1.1255
R11832 VDAC_N.n140 VDAC_N.t1692 1.1255
R11833 VDAC_N.n141 VDAC_N.t119 1.1255
R11834 VDAC_N.n142 VDAC_N.t2053 1.1255
R11835 VDAC_N.n143 VDAC_N.t1432 1.1255
R11836 VDAC_N.n144 VDAC_N.t1841 1.1255
R11837 VDAC_N.n145 VDAC_N.t1012 1.1255
R11838 VDAC_N.n146 VDAC_N.t241 1.1255
R11839 VDAC_N.n147 VDAC_N.t2012 1.1255
R11840 VDAC_N.n148 VDAC_N.t626 1.1255
R11841 VDAC_N.n149 VDAC_N.t285 1.1255
R11842 VDAC_N.n150 VDAC_N.t1552 1.1255
R11843 VDAC_N.n151 VDAC_N.t134 1.1255
R11844 VDAC_N.n152 VDAC_N.t96 1.1255
R11845 VDAC_N.n153 VDAC_N.t766 1.1255
R11846 VDAC_N.n154 VDAC_N.t1020 1.1255
R11847 VDAC_N.n155 VDAC_N.t654 1.1255
R11848 VDAC_N.n156 VDAC_N.t573 1.1255
R11849 VDAC_N.n157 VDAC_N.t1024 1.1255
R11850 VDAC_N.n158 VDAC_N.t293 1.1255
R11851 VDAC_N.n159 VDAC_N.t793 1.1255
R11852 VDAC_N.n160 VDAC_N.t454 1.1255
R11853 VDAC_N.n161 VDAC_N.t1349 1.1255
R11854 VDAC_N.n162 VDAC_N.t263 1.1255
R11855 VDAC_N.n163 VDAC_N.t329 1.1255
R11856 VDAC_N.n164 VDAC_N.t1701 1.1255
R11857 VDAC_N.n165 VDAC_N.t1125 1.1255
R11858 VDAC_N.n166 VDAC_N.t809 1.1255
R11859 VDAC_N.n167 VDAC_N.t2047 1.1255
R11860 VDAC_N.n168 VDAC_N.t753 1.1255
R11861 VDAC_N.n169 VDAC_N.t1937 1.1255
R11862 VDAC_N.n170 VDAC_N.t1940 1.1255
R11863 VDAC_N.n171 VDAC_N.t877 1.1255
R11864 VDAC_N.n172 VDAC_N.t2060 1.1255
R11865 VDAC_N.n173 VDAC_N.t823 1.1255
R11866 VDAC_N.n174 VDAC_N.t2079 1.1255
R11867 VDAC_N.n175 VDAC_N.t1976 1.1255
R11868 VDAC_N.n176 VDAC_N.t997 1.1255
R11869 VDAC_N.n177 VDAC_N.t1112 1.1255
R11870 VDAC_N.n178 VDAC_N.t1714 1.1255
R11871 VDAC_N.n179 VDAC_N.t1316 1.1255
R11872 VDAC_N.n115 VDAC_N.t835 1.1255
R11873 VDAC_N.n180 VDAC_N.t262 1.1255
R11874 VDAC_N.n181 VDAC_N.t779 1.1255
R11875 VDAC_N.n182 VDAC_N.t1670 1.1255
R11876 VDAC_N.n183 VDAC_N.t351 1.1255
R11877 VDAC_N.n184 VDAC_N.t1775 1.1255
R11878 VDAC_N.n185 VDAC_N.t323 1.1255
R11879 VDAC_N.n186 VDAC_N.t1671 1.1255
R11880 VDAC_N.n187 VDAC_N.t2129 1.1255
R11881 VDAC_N.n188 VDAC_N.t795 1.1255
R11882 VDAC_N.n189 VDAC_N.t1023 1.1255
R11883 VDAC_N.n190 VDAC_N.t359 1.1255
R11884 VDAC_N.n191 VDAC_N.t1911 1.1255
R11885 VDAC_N.n192 VDAC_N.t1732 1.1255
R11886 VDAC_N.n193 VDAC_N.t1720 1.1255
R11887 VDAC_N.n194 VDAC_N.t470 1.1255
R11888 VDAC_N.n195 VDAC_N.t1479 1.1255
R11889 VDAC_N.n196 VDAC_N.t418 1.1255
R11890 VDAC_N.n197 VDAC_N.t337 1.1255
R11891 VDAC_N.n198 VDAC_N.t1835 1.1255
R11892 VDAC_N.n199 VDAC_N.t1159 1.1255
R11893 VDAC_N.n200 VDAC_N.t227 1.1255
R11894 VDAC_N.n201 VDAC_N.t2066 1.1255
R11895 VDAC_N.n202 VDAC_N.t399 1.1255
R11896 VDAC_N.n203 VDAC_N.t1967 1.1255
R11897 VDAC_N.n204 VDAC_N.t1295 1.1255
R11898 VDAC_N.n205 VDAC_N.t1867 1.1255
R11899 VDAC_N.n206 VDAC_N.t676 1.1255
R11900 VDAC_N.n207 VDAC_N.t231 1.1255
R11901 VDAC_N.n208 VDAC_N.t252 1.1255
R11902 VDAC_N.n209 VDAC_N.t785 1.1255
R11903 VDAC_N.n210 VDAC_N.t151 1.1255
R11904 VDAC_N.n211 VDAC_N.t848 1.1255
R11905 VDAC_N.n212 VDAC_N.t961 1.1255
R11906 VDAC_N.n213 VDAC_N.t788 1.1255
R11907 VDAC_N.n214 VDAC_N.t1330 1.1255
R11908 VDAC_N.n215 VDAC_N.t1324 1.1255
R11909 VDAC_N.n216 VDAC_N.t574 1.1255
R11910 VDAC_N.n217 VDAC_N.t2029 1.1255
R11911 VDAC_N.n218 VDAC_N.t248 1.1255
R11912 VDAC_N.n219 VDAC_N.t1830 1.1255
R11913 VDAC_N.n220 VDAC_N.t640 1.1255
R11914 VDAC_N.n221 VDAC_N.t1778 1.1255
R11915 VDAC_N.n222 VDAC_N.t1375 1.1255
R11916 VDAC_N.n223 VDAC_N.t1334 1.1255
R11917 VDAC_N.n224 VDAC_N.t591 1.1255
R11918 VDAC_N.n225 VDAC_N.t1719 1.1255
R11919 VDAC_N.n226 VDAC_N.t1042 1.1255
R11920 VDAC_N.n227 VDAC_N.t1507 1.1255
R11921 VDAC_N.n228 VDAC_N.t934 1.1255
R11922 VDAC_N.n229 VDAC_N.t715 1.1255
R11923 VDAC_N.n230 VDAC_N.t945 1.1255
R11924 VDAC_N.n231 VDAC_N.t1287 1.1255
R11925 VDAC_N.n232 VDAC_N.t891 1.1255
R11926 VDAC_N.n233 VDAC_N.t1660 1.1255
R11927 VDAC_N.n234 VDAC_N.t405 1.1255
R11928 VDAC_N.n235 VDAC_N.t2101 1.1255
R11929 VDAC_N.n236 VDAC_N.t1425 1.1255
R11930 VDAC_N.n237 VDAC_N.t1889 1.1255
R11931 VDAC_N.n238 VDAC_N.t1208 1.1255
R11932 VDAC_N.n239 VDAC_N.t1779 1.1255
R11933 VDAC_N.n240 VDAC_N.t652 1.1255
R11934 VDAC_N.n241 VDAC_N.t350 1.1255
R11935 VDAC_N.n242 VDAC_N.t291 1.1255
R11936 VDAC_N.n114 VDAC_N.t1694 1.1255
R11937 VDAC_N.n243 VDAC_N.t1236 1.1255
R11938 VDAC_N.n244 VDAC_N.t1470 1.1255
R11939 VDAC_N.n245 VDAC_N.t1404 1.1255
R11940 VDAC_N.n246 VDAC_N.t2056 1.1255
R11941 VDAC_N.n247 VDAC_N.t150 1.1255
R11942 VDAC_N.n248 VDAC_N.t1632 1.1255
R11943 VDAC_N.n249 VDAC_N.t1746 1.1255
R11944 VDAC_N.n250 VDAC_N.t361 1.1255
R11945 VDAC_N.n251 VDAC_N.t406 1.1255
R11946 VDAC_N.n252 VDAC_N.t1245 1.1255
R11947 VDAC_N.n253 VDAC_N.t162 1.1255
R11948 VDAC_N.n254 VDAC_N.t1133 1.1255
R11949 VDAC_N.n255 VDAC_N.t421 1.1255
R11950 VDAC_N.n256 VDAC_N.t484 1.1255
R11951 VDAC_N.n257 VDAC_N.t714 1.1255
R11952 VDAC_N.n258 VDAC_N.t343 1.1255
R11953 VDAC_N.n259 VDAC_N.t1190 1.1255
R11954 VDAC_N.n260 VDAC_N.t2110 1.1255
R11955 VDAC_N.n261 VDAC_N.t1647 1.1255
R11956 VDAC_N.n262 VDAC_N.t146 1.1255
R11957 VDAC_N.n263 VDAC_N.t203 1.1255
R11958 VDAC_N.n264 VDAC_N.t1682 1.1255
R11959 VDAC_N.n265 VDAC_N.t109 1.1255
R11960 VDAC_N.n266 VDAC_N.t247 1.1255
R11961 VDAC_N.n267 VDAC_N.t1097 1.1255
R11962 VDAC_N.n268 VDAC_N.t131 1.1255
R11963 VDAC_N.n269 VDAC_N.t2133 1.1255
R11964 VDAC_N.n270 VDAC_N.t1459 1.1255
R11965 VDAC_N.n271 VDAC_N.t2023 1.1255
R11966 VDAC_N.n272 VDAC_N.t1357 1.1255
R11967 VDAC_N.n273 VDAC_N.t919 1.1255
R11968 VDAC_N.n274 VDAC_N.t244 1.1255
R11969 VDAC_N.n275 VDAC_N.t867 1.1255
R11970 VDAC_N.n276 VDAC_N.t412 1.1255
R11971 VDAC_N.n277 VDAC_N.t144 1.1255
R11972 VDAC_N.n278 VDAC_N.t1041 1.1255
R11973 VDAC_N.n279 VDAC_N.t72 1.1255
R11974 VDAC_N.n280 VDAC_N.t935 1.1255
R11975 VDAC_N.n281 VDAC_N.t2004 1.1255
R11976 VDAC_N.n282 VDAC_N.t730 1.1255
R11977 VDAC_N.n283 VDAC_N.t908 1.1255
R11978 VDAC_N.n284 VDAC_N.t1390 1.1255
R11979 VDAC_N.n285 VDAC_N.t601 1.1255
R11980 VDAC_N.n286 VDAC_N.t960 1.1255
R11981 VDAC_N.n287 VDAC_N.t962 1.1255
R11982 VDAC_N.n288 VDAC_N.t1529 1.1255
R11983 VDAC_N.n289 VDAC_N.t1666 1.1255
R11984 VDAC_N.n290 VDAC_N.t1317 1.1255
R11985 VDAC_N.n291 VDAC_N.t382 1.1255
R11986 VDAC_N.n292 VDAC_N.t1205 1.1255
R11987 VDAC_N.n293 VDAC_N.t233 1.1255
R11988 VDAC_N.n294 VDAC_N.t1089 1.1255
R11989 VDAC_N.n295 VDAC_N.t1559 1.1255
R11990 VDAC_N.n296 VDAC_N.t2015 1.1255
R11991 VDAC_N.n297 VDAC_N.t689 1.1255
R11992 VDAC_N.n298 VDAC_N.t1909 1.1255
R11993 VDAC_N.n299 VDAC_N.t1233 1.1255
R11994 VDAC_N.n300 VDAC_N.t1703 1.1255
R11995 VDAC_N.n301 VDAC_N.t812 1.1255
R11996 VDAC_N.n302 VDAC_N.t1591 1.1255
R11997 VDAC_N.n303 VDAC_N.t533 1.1255
R11998 VDAC_N.n304 VDAC_N.t1856 1.1255
R11999 VDAC_N.n305 VDAC_N.t983 1.1255
R12000 VDAC_N.n113 VDAC_N.t1975 1.1255
R12001 VDAC_N.n306 VDAC_N.t1305 1.1255
R12002 VDAC_N.n307 VDAC_N.t489 1.1255
R12003 VDAC_N.n308 VDAC_N.t319 1.1255
R12004 VDAC_N.n309 VDAC_N.t1659 1.1255
R12005 VDAC_N.n310 VDAC_N.t2115 1.1255
R12006 VDAC_N.n311 VDAC_N.t787 1.1255
R12007 VDAC_N.n312 VDAC_N.t1015 1.1255
R12008 VDAC_N.n313 VDAC_N.t1264 1.1255
R12009 VDAC_N.n314 VDAC_N.t1899 1.1255
R12010 VDAC_N.n315 VDAC_N.t420 1.1255
R12011 VDAC_N.n316 VDAC_N.t1693 1.1255
R12012 VDAC_N.n317 VDAC_N.t1420 1.1255
R12013 VDAC_N.n318 VDAC_N.t1134 1.1255
R12014 VDAC_N.n319 VDAC_N.t986 1.1255
R12015 VDAC_N.n320 VDAC_N.t735 1.1255
R12016 VDAC_N.n321 VDAC_N.t275 1.1255
R12017 VDAC_N.n322 VDAC_N.t683 1.1255
R12018 VDAC_N.n323 VDAC_N.t911 1.1255
R12019 VDAC_N.n324 VDAC_N.t1620 1.1255
R12020 VDAC_N.n325 VDAC_N.t861 1.1255
R12021 VDAC_N.n326 VDAC_N.t2118 1.1255
R12022 VDAC_N.n327 VDAC_N.t1577 1.1255
R12023 VDAC_N.n328 VDAC_N.t2039 1.1255
R12024 VDAC_N.n329 VDAC_N.t1368 1.1255
R12025 VDAC_N.n330 VDAC_N.t1823 1.1255
R12026 VDAC_N.n331 VDAC_N.t948 1.1255
R12027 VDAC_N.n332 VDAC_N.t718 1.1255
R12028 VDAC_N.n333 VDAC_N.t290 1.1255
R12029 VDAC_N.n334 VDAC_N.t1194 1.1255
R12030 VDAC_N.n335 VDAC_N.t283 1.1255
R12031 VDAC_N.n336 VDAC_N.t752 1.1255
R12032 VDAC_N.n337 VDAC_N.t974 1.1255
R12033 VDAC_N.n338 VDAC_N.t548 1.1255
R12034 VDAC_N.n339 VDAC_N.t746 1.1255
R12035 VDAC_N.n340 VDAC_N.t1217 1.1255
R12036 VDAC_N.n341 VDAC_N.t1250 1.1255
R12037 VDAC_N.n342 VDAC_N.t565 1.1255
R12038 VDAC_N.n343 VDAC_N.t824 1.1255
R12039 VDAC_N.n344 VDAC_N.t1974 1.1255
R12040 VDAC_N.n345 VDAC_N.t1461 1.1255
R12041 VDAC_N.n346 VDAC_N.t1698 1.1255
R12042 VDAC_N.n347 VDAC_N.t39 1.1255
R12043 VDAC_N.n348 VDAC_N.t1897 1.1255
R12044 VDAC_N.n349 VDAC_N.t177 1.1255
R12045 VDAC_N.n350 VDAC_N.t1685 1.1255
R12046 VDAC_N.n351 VDAC_N.t364 1.1255
R12047 VDAC_N.n352 VDAC_N.t799 1.1255
R12048 VDAC_N.n353 VDAC_N.t2033 1.1255
R12049 VDAC_N.n354 VDAC_N.t1465 1.1255
R12050 VDAC_N.n355 VDAC_N.t1923 1.1255
R12051 VDAC_N.n356 VDAC_N.t84 1.1255
R12052 VDAC_N.n357 VDAC_N.t1815 1.1255
R12053 VDAC_N.n358 VDAC_N.t1836 1.1255
R12054 VDAC_N.n359 VDAC_N.t1182 1.1255
R12055 VDAC_N.n360 VDAC_N.t2061 1.1255
R12056 VDAC_N.n361 VDAC_N.t968 1.1255
R12057 VDAC_N.n362 VDAC_N.t987 1.1255
R12058 VDAC_N.n363 VDAC_N.t36 1.1255
R12059 VDAC_N.n364 VDAC_N.t234 1.1255
R12060 VDAC_N.n365 VDAC_N.t596 1.1255
R12061 VDAC_N.n366 VDAC_N.t1246 1.1255
R12062 VDAC_N.n367 VDAC_N.t619 1.1255
R12063 VDAC_N.n368 VDAC_N.t1032 1.1255
R12064 VDAC_N.n112 VDAC_N.t615 1.1255
R12065 VDAC_N.n369 VDAC_N.t2008 1.1255
R12066 VDAC_N.n370 VDAC_N.t557 1.1255
R12067 VDAC_N.n371 VDAC_N.t40 1.1255
R12068 VDAC_N.n372 VDAC_N.t878 1.1255
R12069 VDAC_N.n373 VDAC_N.t687 1.1255
R12070 VDAC_N.n374 VDAC_N.t770 1.1255
R12071 VDAC_N.n375 VDAC_N.t629 1.1255
R12072 VDAC_N.n376 VDAC_N.t1699 1.1255
R12073 VDAC_N.n377 VDAC_N.t575 1.1255
R12074 VDAC_N.n378 VDAC_N.t807 1.1255
R12075 VDAC_N.n379 VDAC_N.t910 1.1255
R12076 VDAC_N.n380 VDAC_N.t751 1.1255
R12077 VDAC_N.n381 VDAC_N.t1933 1.1255
R12078 VDAC_N.n382 VDAC_N.t790 1.1255
R12079 VDAC_N.n383 VDAC_N.t1249 1.1255
R12080 VDAC_N.n384 VDAC_N.t1817 1.1255
R12081 VDAC_N.n385 VDAC_N.t167 1.1255
R12082 VDAC_N.n386 VDAC_N.t1605 1.1255
R12083 VDAC_N.n387 VDAC_N.t18 1.1255
R12084 VDAC_N.n388 VDAC_N.t1495 1.1255
R12085 VDAC_N.n389 VDAC_N.t1949 1.1255
R12086 VDAC_N.n390 VDAC_N.t1389 1.1255
R12087 VDAC_N.n391 VDAC_N.t1853 1.1255
R12088 VDAC_N.n392 VDAC_N.t1172 1.1255
R12089 VDAC_N.n393 VDAC_N.t831 1.1255
R12090 VDAC_N.n394 VDAC_N.t1212 1.1255
R12091 VDAC_N.n395 VDAC_N.t2040 1.1255
R12092 VDAC_N.n396 VDAC_N.t1005 1.1255
R12093 VDAC_N.n397 VDAC_N.t1600 1.1255
R12094 VDAC_N.n398 VDAC_N.t1883 1.1255
R12095 VDAC_N.n399 VDAC_N.t1428 1.1255
R12096 VDAC_N.n400 VDAC_N.t778 1.1255
R12097 VDAC_N.n401 VDAC_N.t588 1.1255
R12098 VDAC_N.n402 VDAC_N.t1090 1.1255
R12099 VDAC_N.n403 VDAC_N.t1026 1.1255
R12100 VDAC_N.n404 VDAC_N.t1728 1.1255
R12101 VDAC_N.n405 VDAC_N.t1806 1.1255
R12102 VDAC_N.n406 VDAC_N.t436 1.1255
R12103 VDAC_N.n407 VDAC_N.t810 1.1255
R12104 VDAC_N.n408 VDAC_N.t183 1.1255
R12105 VDAC_N.n409 VDAC_N.t666 1.1255
R12106 VDAC_N.n410 VDAC_N.t1243 1.1255
R12107 VDAC_N.n411 VDAC_N.t1707 1.1255
R12108 VDAC_N.n412 VDAC_N.t278 1.1255
R12109 VDAC_N.n413 VDAC_N.t1489 1.1255
R12110 VDAC_N.n414 VDAC_N.t535 1.1255
R12111 VDAC_N.n415 VDAC_N.t1383 1.1255
R12112 VDAC_N.n416 VDAC_N.t937 1.1255
R12113 VDAC_N.n417 VDAC_N.t339 1.1255
R12114 VDAC_N.n418 VDAC_N.t1735 1.1255
R12115 VDAC_N.n419 VDAC_N.t92 1.1255
R12116 VDAC_N.n420 VDAC_N.t1627 1.1255
R12117 VDAC_N.n421 VDAC_N.t543 1.1255
R12118 VDAC_N.n422 VDAC_N.t800 1.1255
R12119 VDAC_N.n423 VDAC_N.t259 1.1255
R12120 VDAC_N.n424 VDAC_N.t1136 1.1255
R12121 VDAC_N.n425 VDAC_N.t895 1.1255
R12122 VDAC_N.n426 VDAC_N.t1100 1.1255
R12123 VDAC_N.n427 VDAC_N.t1286 1.1255
R12124 VDAC_N.n428 VDAC_N.t2117 1.1255
R12125 VDAC_N.n429 VDAC_N.t1712 1.1255
R12126 VDAC_N.n430 VDAC_N.t2010 1.1255
R12127 VDAC_N.n431 VDAC_N.t1272 1.1255
R12128 VDAC_N.n111 VDAC_N.t180 1.1255
R12129 VDAC_N.n432 VDAC_N.t837 1.1255
R12130 VDAC_N.n433 VDAC_N.t1468 1.1255
R12131 VDAC_N.n434 VDAC_N.t781 1.1255
R12132 VDAC_N.n435 VDAC_N.t1991 1.1255
R12133 VDAC_N.n436 VDAC_N.t176 1.1255
R12134 VDAC_N.n437 VDAC_N.t493 1.1255
R12135 VDAC_N.n438 VDAC_N.t1476 1.1255
R12136 VDAC_N.n439 VDAC_N.t1318 1.1255
R12137 VDAC_N.n440 VDAC_N.t1228 1.1255
R12138 VDAC_N.n441 VDAC_N.t566 1.1255
R12139 VDAC_N.n442 VDAC_N.t527 1.1255
R12140 VDAC_N.n443 VDAC_N.t888 1.1255
R12141 VDAC_N.n444 VDAC_N.t922 1.1255
R12142 VDAC_N.n445 VDAC_N.t1511 1.1255
R12143 VDAC_N.n446 VDAC_N.t1963 1.1255
R12144 VDAC_N.n447 VDAC_N.t400 1.1255
R12145 VDAC_N.n448 VDAC_N.t1865 1.1255
R12146 VDAC_N.n449 VDAC_N.t660 1.1255
R12147 VDAC_N.n450 VDAC_N.t1482 1.1255
R12148 VDAC_N.n451 VDAC_N.t892 1.1255
R12149 VDAC_N.n452 VDAC_N.t2080 1.1255
R12150 VDAC_N.n453 VDAC_N.t2103 1.1255
R12151 VDAC_N.n454 VDAC_N.t232 1.1255
R12152 VDAC_N.n455 VDAC_N.t462 1.1255
R12153 VDAC_N.n456 VDAC_N.t404 1.1255
R12154 VDAC_N.n457 VDAC_N.t410 1.1255
R12155 VDAC_N.n458 VDAC_N.t1253 1.1255
R12156 VDAC_N.n459 VDAC_N.t1114 1.1255
R12157 VDAC_N.n460 VDAC_N.t585 1.1255
R12158 VDAC_N.n461 VDAC_N.t1784 1.1255
R12159 VDAC_N.n462 VDAC_N.t1826 1.1255
R12160 VDAC_N.n463 VDAC_N.t1497 1.1255
R12161 VDAC_N.n464 VDAC_N.t822 1.1255
R12162 VDAC_N.n465 VDAC_N.t1281 1.1255
R12163 VDAC_N.n466 VDAC_N.t1747 1.1255
R12164 VDAC_N.n467 VDAC_N.t1171 1.1255
R12165 VDAC_N.n468 VDAC_N.t1639 1.1255
R12166 VDAC_N.n469 VDAC_N.t1890 1.1255
R12167 VDAC_N.n470 VDAC_N.t777 1.1255
R12168 VDAC_N.n471 VDAC_N.t1007 1.1255
R12169 VDAC_N.n472 VDAC_N.t371 1.1255
R12170 VDAC_N.n473 VDAC_N.t1953 1.1255
R12171 VDAC_N.n474 VDAC_N.t1076 1.1255
R12172 VDAC_N.n475 VDAC_N.t1751 1.1255
R12173 VDAC_N.n476 VDAC_N.t1532 1.1255
R12174 VDAC_N.n477 VDAC_N.t642 1.1255
R12175 VDAC_N.n478 VDAC_N.t545 1.1255
R12176 VDAC_N.n479 VDAC_N.t432 1.1255
R12177 VDAC_N.n480 VDAC_N.t1989 1.1255
R12178 VDAC_N.n481 VDAC_N.t320 1.1255
R12179 VDAC_N.n482 VDAC_N.t1546 1.1255
R12180 VDAC_N.n483 VDAC_N.t1460 1.1255
R12181 VDAC_N.n484 VDAC_N.t1310 1.1255
R12182 VDAC_N.n485 VDAC_N.t1137 1.1255
R12183 VDAC_N.n486 VDAC_N.t1760 1.1255
R12184 VDAC_N.n487 VDAC_N.t530 1.1255
R12185 VDAC_N.n488 VDAC_N.t48 1.1255
R12186 VDAC_N.n489 VDAC_N.t1610 1.1255
R12187 VDAC_N.n490 VDAC_N.t113 1.1255
R12188 VDAC_N.n491 VDAC_N.t1366 1.1255
R12189 VDAC_N.n492 VDAC_N.t599 1.1255
R12190 VDAC_N.n493 VDAC_N.t883 1.1255
R12191 VDAC_N.n494 VDAC_N.t2090 1.1255
R12192 VDAC_N.n110 VDAC_N.t407 1.1255
R12193 VDAC_N.n495 VDAC_N.t446 1.1255
R12194 VDAC_N.n496 VDAC_N.t1435 1.1255
R12195 VDAC_N.n497 VDAC_N.t1474 1.1255
R12196 VDAC_N.n498 VDAC_N.t1221 1.1255
R12197 VDAC_N.n499 VDAC_N.t857 1.1255
R12198 VDAC_N.n500 VDAC_N.t1107 1.1255
R12199 VDAC_N.n501 VDAC_N.t1569 1.1255
R12200 VDAC_N.n502 VDAC_N.t2035 1.1255
R12201 VDAC_N.n503 VDAC_N.t387 1.1255
R12202 VDAC_N.n504 VDAC_N.t975 1.1255
R12203 VDAC_N.n505 VDAC_N.t333 1.1255
R12204 VDAC_N.n506 VDAC_N.t475 1.1255
R12205 VDAC_N.n507 VDAC_N.t140 1.1255
R12206 VDAC_N.n508 VDAC_N.t1323 1.1255
R12207 VDAC_N.n509 VDAC_N.t903 1.1255
R12208 VDAC_N.n510 VDAC_N.t388 1.1255
R12209 VDAC_N.n511 VDAC_N.t851 1.1255
R12210 VDAC_N.n512 VDAC_N.t2131 1.1255
R12211 VDAC_N.n513 VDAC_N.t1098 1.1255
R12212 VDAC_N.n514 VDAC_N.t2021 1.1255
R12213 VDAC_N.n515 VDAC_N.t672 1.1255
R12214 VDAC_N.n516 VDAC_N.t1913 1.1255
R12215 VDAC_N.n517 VDAC_N.t1748 1.1255
R12216 VDAC_N.n518 VDAC_N.t1370 1.1255
R12217 VDAC_N.n519 VDAC_N.t924 1.1255
R12218 VDAC_N.n520 VDAC_N.t594 1.1255
R12219 VDAC_N.n521 VDAC_N.t286 1.1255
R12220 VDAC_N.n522 VDAC_N.t1424 1.1255
R12221 VDAC_N.n523 VDAC_N.t1874 1.1255
R12222 VDAC_N.n524 VDAC_N.t1988 1.1255
R12223 VDAC_N.n525 VDAC_N.t378 1.1255
R12224 VDAC_N.n526 VDAC_N.t1309 1.1255
R12225 VDAC_N.n527 VDAC_N.t1222 1.1255
R12226 VDAC_N.n528 VDAC_N.t1083 1.1255
R12227 VDAC_N.n529 VDAC_N.t791 1.1255
R12228 VDAC_N.n530 VDAC_N.t58 1.1255
R12229 VDAC_N.n531 VDAC_N.t1447 1.1255
R12230 VDAC_N.n532 VDAC_N.t74 1.1255
R12231 VDAC_N.n533 VDAC_N.t1341 1.1255
R12232 VDAC_N.n534 VDAC_N.t913 1.1255
R12233 VDAC_N.n535 VDAC_N.t1203 1.1255
R12234 VDAC_N.n536 VDAC_N.t899 1.1255
R12235 VDAC_N.n537 VDAC_N.t172 1.1255
R12236 VDAC_N.n538 VDAC_N.t219 1.1255
R12237 VDAC_N.n539 VDAC_N.t2013 1.1255
R12238 VDAC_N.n540 VDAC_N.t1736 1.1255
R12239 VDAC_N.n541 VDAC_N.t1905 1.1255
R12240 VDAC_N.n542 VDAC_N.t132 1.1255
R12241 VDAC_N.n543 VDAC_N.t915 1.1255
R12242 VDAC_N.n544 VDAC_N.t1580 1.1255
R12243 VDAC_N.n545 VDAC_N.t1150 1.1255
R12244 VDAC_N.n546 VDAC_N.t220 1.1255
R12245 VDAC_N.n547 VDAC_N.t256 1.1255
R12246 VDAC_N.n548 VDAC_N.t946 1.1255
R12247 VDAC_N.n549 VDAC_N.t980 1.1255
R12248 VDAC_N.n550 VDAC_N.t230 1.1255
R12249 VDAC_N.n551 VDAC_N.t1996 1.1255
R12250 VDAC_N.n552 VDAC_N.t1214 1.1255
R12251 VDAC_N.n553 VDAC_N.t1191 1.1255
R12252 VDAC_N.n554 VDAC_N.t512 1.1255
R12253 VDAC_N.n555 VDAC_N.t506 1.1255
R12254 VDAC_N.n556 VDAC_N.t1545 1.1255
R12255 VDAC_N.n557 VDAC_N.t1710 1.1255
R12256 VDAC_N.n109 VDAC_N.t1506 1.1255
R12257 VDAC_N.n558 VDAC_N.t2044 1.1255
R12258 VDAC_N.n559 VDAC_N.t1282 1.1255
R12259 VDAC_N.n560 VDAC_N.t549 1.1255
R12260 VDAC_N.n561 VDAC_N.t80 1.1255
R12261 VDAC_N.n562 VDAC_N.t466 1.1255
R12262 VDAC_N.n563 VDAC_N.t1248 1.1255
R12263 VDAC_N.n564 VDAC_N.t1570 1.1255
R12264 VDAC_N.n565 VDAC_N.t1259 1.1255
R12265 VDAC_N.n566 VDAC_N.t354 1.1255
R12266 VDAC_N.n567 VDAC_N.t589 1.1255
R12267 VDAC_N.n568 VDAC_N.t1808 1.1255
R12268 VDAC_N.n569 VDAC_N.t2050 1.1255
R12269 VDAC_N.n570 VDAC_N.t1503 1.1255
R12270 VDAC_N.n571 VDAC_N.t165 1.1255
R12271 VDAC_N.n572 VDAC_N.t1589 1.1255
R12272 VDAC_N.n573 VDAC_N.t1500 1.1255
R12273 VDAC_N.n574 VDAC_N.t1477 1.1255
R12274 VDAC_N.n575 VDAC_N.t505 1.1255
R12275 VDAC_N.n576 VDAC_N.t1400 1.1255
R12276 VDAC_N.n577 VDAC_N.t931 1.1255
R12277 VDAC_N.n578 VDAC_N.t1036 1.1255
R12278 VDAC_N.n579 VDAC_N.t1723 1.1255
R12279 VDAC_N.n580 VDAC_N.t26 1.1255
R12280 VDAC_N.n581 VDAC_N.t1968 1.1255
R12281 VDAC_N.n582 VDAC_N.t149 1.1255
R12282 VDAC_N.n583 VDAC_N.t1520 1.1255
R12283 VDAC_N.n584 VDAC_N.t870 1.1255
R12284 VDAC_N.n585 VDAC_N.t1300 1.1255
R12285 VDAC_N.n586 VDAC_N.t210 1.1255
R12286 VDAC_N.n587 VDAC_N.t1788 1.1255
R12287 VDAC_N.n588 VDAC_N.t2088 1.1255
R12288 VDAC_N.n589 VDAC_N.t569 1.1255
R12289 VDAC_N.n590 VDAC_N.t1664 1.1255
R12290 VDAC_N.n591 VDAC_N.t1766 1.1255
R12291 VDAC_N.n592 VDAC_N.t1369 1.1255
R12292 VDAC_N.n593 VDAC_N.t1558 1.1255
R12293 VDAC_N.n594 VDAC_N.t641 1.1255
R12294 VDAC_N.n595 VDAC_N.t62 1.1255
R12295 VDAC_N.n596 VDAC_N.t1143 1.1255
R12296 VDAC_N.n597 VDAC_N.t423 1.1255
R12297 VDAC_N.n598 VDAC_N.t2006 1.1255
R12298 VDAC_N.n599 VDAC_N.t417 1.1255
R12299 VDAC_N.n600 VDAC_N.t1035 1.1255
R12300 VDAC_N.n601 VDAC_N.t701 1.1255
R12301 VDAC_N.n602 VDAC_N.t1829 1.1255
R12302 VDAC_N.n603 VDAC_N.t260 1.1255
R12303 VDAC_N.n604 VDAC_N.t1717 1.1255
R12304 VDAC_N.n605 VDAC_N.t24 1.1255
R12305 VDAC_N.n606 VDAC_N.t127 1.1255
R12306 VDAC_N.n607 VDAC_N.t2071 1.1255
R12307 VDAC_N.n608 VDAC_N.t1496 1.1255
R12308 VDAC_N.n609 VDAC_N.t1955 1.1255
R12309 VDAC_N.n610 VDAC_N.t2132 1.1255
R12310 VDAC_N.n611 VDAC_N.t750 1.1255
R12311 VDAC_N.n612 VDAC_N.t1596 1.1255
R12312 VDAC_N.n613 VDAC_N.t1258 1.1255
R12313 VDAC_N.n614 VDAC_N.t287 1.1255
R12314 VDAC_N.n615 VDAC_N.t840 1.1255
R12315 VDAC_N.n616 VDAC_N.t1978 1.1255
R12316 VDAC_N.n617 VDAC_N.t616 1.1255
R12317 VDAC_N.n618 VDAC_N.t1550 1.1255
R12318 VDAC_N.n619 VDAC_N.t1361 1.1255
R12319 VDAC_N.n620 VDAC_N.t1314 1.1255
R12320 VDAC_N.n108 VDAC_N.t57 1.1255
R12321 VDAC_N.n621 VDAC_N.t1207 1.1255
R12322 VDAC_N.n622 VDAC_N.t1771 1.1255
R12323 VDAC_N.n623 VDAC_N.t559 1.1255
R12324 VDAC_N.n624 VDAC_N.t1561 1.1255
R12325 VDAC_N.n625 VDAC_N.t2017 1.1255
R12326 VDAC_N.n626 VDAC_N.t117 1.1255
R12327 VDAC_N.n627 VDAC_N.t969 1.1255
R12328 VDAC_N.n628 VDAC_N.t452 1.1255
R12329 VDAC_N.n629 VDAC_N.t1803 1.1255
R12330 VDAC_N.n630 VDAC_N.t1612 1.1255
R12331 VDAC_N.n631 VDAC_N.t419 1.1255
R12332 VDAC_N.n632 VDAC_N.t732 1.1255
R12333 VDAC_N.n633 VDAC_N.t944 1.1255
R12334 VDAC_N.n634 VDAC_N.t85 1.1255
R12335 VDAC_N.n635 VDAC_N.t308 1.1255
R12336 VDAC_N.n636 VDAC_N.t1446 1.1255
R12337 VDAC_N.n637 VDAC_N.t1148 1.1255
R12338 VDAC_N.n638 VDAC_N.t528 1.1255
R12339 VDAC_N.n639 VDAC_N.t161 1.1255
R12340 VDAC_N.n640 VDAC_N.t1592 1.1255
R12341 VDAC_N.n641 VDAC_N.t1738 1.1255
R12342 VDAC_N.n642 VDAC_N.t592 1.1255
R12343 VDAC_N.n643 VDAC_N.t1526 1.1255
R12344 VDAC_N.n644 VDAC_N.t1235 1.1255
R12345 VDAC_N.n645 VDAC_N.t1082 1.1255
R12346 VDAC_N.n646 VDAC_N.t577 1.1255
R12347 VDAC_N.n647 VDAC_N.t1593 1.1255
R12348 VDAC_N.n648 VDAC_N.t914 1.1255
R12349 VDAC_N.n649 VDAC_N.t391 1.1255
R12350 VDAC_N.n650 VDAC_N.t1590 1.1255
R12351 VDAC_N.n651 VDAC_N.t1265 1.1255
R12352 VDAC_N.n652 VDAC_N.t1837 1.1255
R12353 VDAC_N.n653 VDAC_N.t311 1.1255
R12354 VDAC_N.n654 VDAC_N.t825 1.1255
R12355 VDAC_N.n655 VDAC_N.t1055 1.1255
R12356 VDAC_N.n656 VDAC_N.t1513 1.1255
R12357 VDAC_N.n657 VDAC_N.t1969 1.1255
R12358 VDAC_N.n658 VDAC_N.t663 1.1255
R12359 VDAC_N.n659 VDAC_N.t143 1.1255
R12360 VDAC_N.n660 VDAC_N.t1332 1.1255
R12361 VDAC_N.n661 VDAC_N.t881 1.1255
R12362 VDAC_N.n662 VDAC_N.t1092 1.1255
R12363 VDAC_N.n663 VDAC_N.t1230 1.1255
R12364 VDAC_N.n664 VDAC_N.t1057 1.1255
R12365 VDAC_N.n665 VDAC_N.t1560 1.1255
R12366 VDAC_N.n666 VDAC_N.t990 1.1255
R12367 VDAC_N.n667 VDAC_N.t576 1.1255
R12368 VDAC_N.n668 VDAC_N.t398 1.1255
R12369 VDAC_N.n669 VDAC_N.t1364 1.1255
R12370 VDAC_N.n670 VDAC_N.t342 1.1255
R12371 VDAC_N.n671 VDAC_N.t301 1.1255
R12372 VDAC_N.n672 VDAC_N.t1064 1.1255
R12373 VDAC_N.n673 VDAC_N.t1018 1.1255
R12374 VDAC_N.n674 VDAC_N.t1473 1.1255
R12375 VDAC_N.n675 VDAC_N.t1578 1.1255
R12376 VDAC_N.n676 VDAC_N.t365 1.1255
R12377 VDAC_N.n677 VDAC_N.t682 1.1255
R12378 VDAC_N.n678 VDAC_N.t1155 1.1255
R12379 VDAC_N.n679 VDAC_N.t451 1.1255
R12380 VDAC_N.n680 VDAC_N.t2058 1.1255
R12381 VDAC_N.n681 VDAC_N.t1509 1.1255
R12382 VDAC_N.n682 VDAC_N.t2073 1.1255
R12383 VDAC_N.n683 VDAC_N.t1403 1.1255
R12384 VDAC_N.n107 VDAC_N.t297 1.1255
R12385 VDAC_N.n684 VDAC_N.t128 1.1255
R12386 VDAC_N.n685 VDAC_N.t1002 1.1255
R12387 VDAC_N.n686 VDAC_N.t608 1.1255
R12388 VDAC_N.n687 VDAC_N.t1538 1.1255
R12389 VDAC_N.n688 VDAC_N.t47 1.1255
R12390 VDAC_N.n689 VDAC_N.t1306 1.1255
R12391 VDAC_N.n690 VDAC_N.t97 1.1255
R12392 VDAC_N.n691 VDAC_N.t1599 1.1255
R12393 VDAC_N.n692 VDAC_N.t2030 1.1255
R12394 VDAC_N.n693 VDAC_N.t759 1.1255
R12395 VDAC_N.n694 VDAC_N.t422 1.1255
R12396 VDAC_N.n695 VDAC_N.t1385 1.1255
R12397 VDAC_N.n696 VDAC_N.t483 1.1255
R12398 VDAC_N.n697 VDAC_N.t79 1.1255
R12399 VDAC_N.n698 VDAC_N.t289 1.1255
R12400 VDAC_N.n699 VDAC_N.t2104 1.1255
R12401 VDAC_N.n700 VDAC_N.t2003 1.1255
R12402 VDAC_N.n701 VDAC_N.t648 1.1255
R12403 VDAC_N.n702 VDAC_N.t906 1.1255
R12404 VDAC_N.n703 VDAC_N.t1604 1.1255
R12405 VDAC_N.n704 VDAC_N.t1342 1.1255
R12406 VDAC_N.n705 VDAC_N.t716 1.1255
R12407 VDAC_N.n706 VDAC_N.t166 1.1255
R12408 VDAC_N.n707 VDAC_N.t282 1.1255
R12409 VDAC_N.n708 VDAC_N.t1360 1.1255
R12410 VDAC_N.n709 VDAC_N.t1842 1.1255
R12411 VDAC_N.n710 VDAC_N.t71 1.1255
R12412 VDAC_N.n711 VDAC_N.t114 1.1255
R12413 VDAC_N.n712 VDAC_N.t659 1.1255
R12414 VDAC_N.n713 VDAC_N.t610 1.1255
R12415 VDAC_N.n714 VDAC_N.t10 1.1255
R12416 VDAC_N.n715 VDAC_N.t433 1.1255
R12417 VDAC_N.n716 VDAC_N.t1918 1.1255
R12418 VDAC_N.n717 VDAC_N.t729 1.1255
R12419 VDAC_N.n718 VDAC_N.t1893 1.1255
R12420 VDAC_N.n719 VDAC_N.t677 1.1255
R12421 VDAC_N.n720 VDAC_N.t1783 1.1255
R12422 VDAC_N.n721 VDAC_N.t95 1.1255
R12423 VDAC_N.n722 VDAC_N.t1677 1.1255
R12424 VDAC_N.n723 VDAC_N.t2106 1.1255
R12425 VDAC_N.n724 VDAC_N.t1543 1.1255
R12426 VDAC_N.n725 VDAC_N.t1069 1.1255
R12427 VDAC_N.n726 VDAC_N.t1680 1.1255
R12428 VDAC_N.n727 VDAC_N.t495 1.1255
R12429 VDAC_N.n728 VDAC_N.t52 1.1255
R12430 VDAC_N.n729 VDAC_N.t34 1.1255
R12431 VDAC_N.n730 VDAC_N.t684 1.1255
R12432 VDAC_N.n731 VDAC_N.t302 1.1255
R12433 VDAC_N.n732 VDAC_N.t693 1.1255
R12434 VDAC_N.n733 VDAC_N.t912 1.1255
R12435 VDAC_N.n734 VDAC_N.t1834 1.1255
R12436 VDAC_N.n735 VDAC_N.t1336 1.1255
R12437 VDAC_N.n736 VDAC_N.t1622 1.1255
R12438 VDAC_N.n737 VDAC_N.t185 1.1255
R12439 VDAC_N.n738 VDAC_N.t1178 1.1255
R12440 VDAC_N.n739 VDAC_N.t1177 1.1255
R12441 VDAC_N.n740 VDAC_N.t1896 1.1255
R12442 VDAC_N.n741 VDAC_N.t1902 1.1255
R12443 VDAC_N.n742 VDAC_N.t75 1.1255
R12444 VDAC_N.n743 VDAC_N.t850 1.1255
R12445 VDAC_N.n744 VDAC_N.t1321 1.1255
R12446 VDAC_N.n745 VDAC_N.t957 1.1255
R12447 VDAC_N.n746 VDAC_N.t1209 1.1255
R12448 VDAC_N.n106 VDAC_N.t1006 1.1255
R12449 VDAC_N.n747 VDAC_N.t1216 1.1255
R12450 VDAC_N.n748 VDAC_N.t1750 1.1255
R12451 VDAC_N.n749 VDAC_N.t756 1.1255
R12452 VDAC_N.n750 VDAC_N.t674 1.1255
R12453 VDAC_N.n751 VDAC_N.t1141 1.1255
R12454 VDAC_N.n752 VDAC_N.t1106 1.1255
R12455 VDAC_N.n753 VDAC_N.t2038 1.1255
R12456 VDAC_N.n754 VDAC_N.t395 1.1255
R12457 VDAC_N.n755 VDAC_N.t1818 1.1255
R12458 VDAC_N.n756 VDAC_N.t709 1.1255
R12459 VDAC_N.n757 VDAC_N.t1374 1.1255
R12460 VDAC_N.n758 VDAC_N.t1275 1.1255
R12461 VDAC_N.n759 VDAC_N.t1741 1.1255
R12462 VDAC_N.n760 VDAC_N.t1515 1.1255
R12463 VDAC_N.n761 VDAC_N.t1971 1.1255
R12464 VDAC_N.n762 VDAC_N.t784 1.1255
R12465 VDAC_N.n763 VDAC_N.t949 1.1255
R12466 VDAC_N.n764 VDAC_N.t356 1.1255
R12467 VDAC_N.n765 VDAC_N.t762 1.1255
R12468 VDAC_N.n766 VDAC_N.t508 1.1255
R12469 VDAC_N.n767 VDAC_N.t544 1.1255
R12470 VDAC_N.n768 VDAC_N.t2111 1.1255
R12471 VDAC_N.n769 VDAC_N.t856 1.1255
R12472 VDAC_N.n770 VDAC_N.t246 1.1255
R12473 VDAC_N.n771 VDAC_N.t1572 1.1255
R12474 VDAC_N.n772 VDAC_N.t1566 1.1255
R12475 VDAC_N.n773 VDAC_N.t1257 1.1255
R12476 VDAC_N.n774 VDAC_N.t578 1.1255
R12477 VDAC_N.n775 VDAC_N.t63 1.1255
R12478 VDAC_N.n776 VDAC_N.t1800 1.1255
R12479 VDAC_N.n777 VDAC_N.t1838 1.1255
R12480 VDAC_N.n778 VDAC_N.t765 1.1255
R12481 VDAC_N.n779 VDAC_N.t826 1.1255
R12482 VDAC_N.n780 VDAC_N.t1285 1.1255
R12483 VDAC_N.n781 VDAC_N.t1749 1.1255
R12484 VDAC_N.n782 VDAC_N.t603 1.1255
R12485 VDAC_N.n783 VDAC_N.t129 1.1255
R12486 VDAC_N.n784 VDAC_N.t1906 1.1255
R12487 VDAC_N.n785 VDAC_N.t1533 1.1255
R12488 VDAC_N.n786 VDAC_N.t273 1.1255
R12489 VDAC_N.n787 VDAC_N.t717 1.1255
R12490 VDAC_N.n788 VDAC_N.t511 1.1255
R12491 VDAC_N.n789 VDAC_N.t1096 1.1255
R12492 VDAC_N.n790 VDAC_N.t55 1.1255
R12493 VDAC_N.n791 VDAC_N.t1852 1.1255
R12494 VDAC_N.n792 VDAC_N.t1266 1.1255
R12495 VDAC_N.n793 VDAC_N.t547 1.1255
R12496 VDAC_N.n794 VDAC_N.t1672 1.1255
R12497 VDAC_N.n795 VDAC_N.t1995 1.1255
R12498 VDAC_N.n796 VDAC_N.t328 1.1255
R12499 VDAC_N.n797 VDAC_N.t794 1.1255
R12500 VDAC_N.n798 VDAC_N.t772 1.1255
R12501 VDAC_N.n799 VDAC_N.t190 1.1255
R12502 VDAC_N.n800 VDAC_N.t1145 1.1255
R12503 VDAC_N.n801 VDAC_N.t1792 1.1255
R12504 VDAC_N.n802 VDAC_N.t154 1.1255
R12505 VDAC_N.n803 VDAC_N.t352 1.1255
R12506 VDAC_N.n804 VDAC_N.t1618 1.1255
R12507 VDAC_N.n805 VDAC_N.t711 1.1255
R12508 VDAC_N.n806 VDAC_N.t1382 1.1255
R12509 VDAC_N.n807 VDAC_N.t171 1.1255
R12510 VDAC_N.n808 VDAC_N.t887 1.1255
R12511 VDAC_N.n809 VDAC_N.t2098 1.1255
R12512 VDAC_N.n105 VDAC_N.t804 1.1255
R12513 VDAC_N.n810 VDAC_N.t1689 1.1255
R12514 VDAC_N.n811 VDAC_N.t1388 1.1255
R12515 VDAC_N.n812 VDAC_N.t801 1.1255
R12516 VDAC_N.n813 VDAC_N.t1033 1.1255
R12517 VDAC_N.n814 VDAC_N.t1352 1.1255
R12518 VDAC_N.n815 VDAC_N.t1925 1.1255
R12519 VDAC_N.n816 VDAC_N.t1844 1.1255
R12520 VDAC_N.n817 VDAC_N.t1398 1.1255
R12521 VDAC_N.n818 VDAC_N.t1868 1.1255
R12522 VDAC_N.n819 VDAC_N.t318 1.1255
R12523 VDAC_N.n820 VDAC_N.t537 1.1255
R12524 VDAC_N.n821 VDAC_N.t264 1.1255
R12525 VDAC_N.n822 VDAC_N.t1914 1.1255
R12526 VDAC_N.n823 VDAC_N.t353 1.1255
R12527 VDAC_N.n824 VDAC_N.t1785 1.1255
R12528 VDAC_N.n825 VDAC_N.t1524 1.1255
R12529 VDAC_N.n826 VDAC_N.t441 1.1255
R12530 VDAC_N.n827 VDAC_N.t93 1.1255
R12531 VDAC_N.n828 VDAC_N.t570 1.1255
R12532 VDAC_N.n829 VDAC_N.t153 1.1255
R12533 VDAC_N.n830 VDAC_N.t1328 1.1255
R12534 VDAC_N.n831 VDAC_N.t501 1.1255
R12535 VDAC_N.n832 VDAC_N.t468 1.1255
R12536 VDAC_N.n833 VDAC_N.t706 1.1255
R12537 VDAC_N.n834 VDAC_N.t1180 1.1255
R12538 VDAC_N.n835 VDAC_N.t598 1.1255
R12539 VDAC_N.n836 VDAC_N.t546 1.1255
R12540 VDAC_N.n837 VDAC_N.t384 1.1255
R12541 VDAC_N.n838 VDAC_N.t958 1.1255
R12542 VDAC_N.n839 VDAC_N.t2020 1.1255
R12543 VDAC_N.n840 VDAC_N.t1442 1.1255
R12544 VDAC_N.n841 VDAC_N.t671 1.1255
R12545 VDAC_N.n842 VDAC_N.t630 1.1255
R12546 VDAC_N.n843 VDAC_N.t1087 1.1255
R12547 VDAC_N.n844 VDAC_N.t1555 1.1255
R12548 VDAC_N.n845 VDAC_N.t1954 1.1255
R12549 VDAC_N.n846 VDAC_N.t1451 1.1255
R12550 VDAC_N.n847 VDAC_N.t214 1.1255
R12551 VDAC_N.n848 VDAC_N.t1345 1.1255
R12552 VDAC_N.n849 VDAC_N.t471 1.1255
R12553 VDAC_N.n850 VDAC_N.t1213 1.1255
R12554 VDAC_N.n851 VDAC_N.t465 1.1255
R12555 VDAC_N.n852 VDAC_N.t332 1.1255
R12556 VDAC_N.n853 VDAC_N.t1563 1.1255
R12557 VDAC_N.n854 VDAC_N.t2025 1.1255
R12558 VDAC_N.n855 VDAC_N.t136 1.1255
R12559 VDAC_N.n856 VDAC_N.t971 1.1255
R12560 VDAC_N.n857 VDAC_N.t1764 1.1255
R12561 VDAC_N.n858 VDAC_N.t1807 1.1255
R12562 VDAC_N.n859 VDAC_N.t1676 1.1255
R12563 VDAC_N.n860 VDAC_N.t1162 1.1255
R12564 VDAC_N.n861 VDAC_N.t1116 1.1255
R12565 VDAC_N.n862 VDAC_N.t952 1.1255
R12566 VDAC_N.n863 VDAC_N.t954 1.1255
R12567 VDAC_N.n864 VDAC_N.t276 1.1255
R12568 VDAC_N.n865 VDAC_N.t1654 1.1255
R12569 VDAC_N.n866 VDAC_N.t44 1.1255
R12570 VDAC_N.n867 VDAC_N.t1226 1.1255
R12571 VDAC_N.n868 VDAC_N.t613 1.1255
R12572 VDAC_N.n869 VDAC_N.t1992 1.1255
R12573 VDAC_N.n870 VDAC_N.t1950 1.1255
R12574 VDAC_N.n871 VDAC_N.t409 1.1255
R12575 VDAC_N.n872 VDAC_N.t1718 1.1255
R12576 VDAC_N.n104 VDAC_N.t1585 1.1255
R12577 VDAC_N.n873 VDAC_N.t1782 1.1255
R12578 VDAC_N.n874 VDAC_N.t389 1.1255
R12579 VDAC_N.n875 VDAC_N.t414 1.1255
R12580 VDAC_N.n876 VDAC_N.t105 1.1255
R12581 VDAC_N.n877 VDAC_N.t1721 1.1255
R12582 VDAC_N.n878 VDAC_N.t1153 1.1255
R12583 VDAC_N.n879 VDAC_N.t1613 1.1255
R12584 VDAC_N.n880 VDAC_N.t539 1.1255
R12585 VDAC_N.n881 VDAC_N.t767 1.1255
R12586 VDAC_N.n882 VDAC_N.t993 1.1255
R12587 VDAC_N.n883 VDAC_N.t1289 1.1255
R12588 VDAC_N.n884 VDAC_N.t257 1.1255
R12589 VDAC_N.n885 VDAC_N.t1268 1.1255
R12590 VDAC_N.n886 VDAC_N.t1129 1.1255
R12591 VDAC_N.n887 VDAC_N.t1595 1.1255
R12592 VDAC_N.n888 VDAC_N.t156 1.1255
R12593 VDAC_N.n889 VDAC_N.t1483 1.1255
R12594 VDAC_N.n890 VDAC_N.t1939 1.1255
R12595 VDAC_N.n891 VDAC_N.t376 1.1255
R12596 VDAC_N.n892 VDAC_N.t481 1.1255
R12597 VDAC_N.n893 VDAC_N.t2092 1.1255
R12598 VDAC_N.n894 VDAC_N.t1731 1.1255
R12599 VDAC_N.n895 VDAC_N.t28 1.1255
R12600 VDAC_N.n896 VDAC_N.t520 1.1255
R12601 VDAC_N.n897 VDAC_N.t271 1.1255
R12602 VDAC_N.n898 VDAC_N.t1544 1.1255
R12603 VDAC_N.n899 VDAC_N.t874 1.1255
R12604 VDAC_N.n900 VDAC_N.t1348 1.1255
R12605 VDAC_N.n901 VDAC_N.t1498 1.1255
R12606 VDAC_N.n902 VDAC_N.t1980 1.1255
R12607 VDAC_N.n903 VDAC_N.t2096 1.1255
R12608 VDAC_N.n904 VDAC_N.t45 1.1255
R12609 VDAC_N.n905 VDAC_N.t1688 1.1255
R12610 VDAC_N.n906 VDAC_N.t1774 1.1255
R12611 VDAC_N.n907 VDAC_N.t49 1.1255
R12612 VDAC_N.n908 VDAC_N.t798 1.1255
R12613 VDAC_N.n909 VDAC_N.t643 1.1255
R12614 VDAC_N.n910 VDAC_N.t1130 1.1255
R12615 VDAC_N.n911 VDAC_N.t1149 1.1255
R12616 VDAC_N.n912 VDAC_N.t819 1.1255
R12617 VDAC_N.n913 VDAC_N.t2014 1.1255
R12618 VDAC_N.n914 VDAC_N.t223 1.1255
R12619 VDAC_N.n915 VDAC_N.t2045 1.1255
R12620 VDAC_N.n916 VDAC_N.t1377 1.1255
R12621 VDAC_N.n917 VDAC_N.t141 1.1255
R12622 VDAC_N.n918 VDAC_N.t500 1.1255
R12623 VDAC_N.n919 VDAC_N.t81 1.1255
R12624 VDAC_N.n920 VDAC_N.t988 1.1255
R12625 VDAC_N.n921 VDAC_N.t425 1.1255
R12626 VDAC_N.n922 VDAC_N.t2077 1.1255
R12627 VDAC_N.n923 VDAC_N.t776 1.1255
R12628 VDAC_N.n924 VDAC_N.t995 1.1255
R12629 VDAC_N.n925 VDAC_N.t296 1.1255
R12630 VDAC_N.n926 VDAC_N.t758 1.1255
R12631 VDAC_N.n927 VDAC_N.t956 1.1255
R12632 VDAC_N.n928 VDAC_N.t1270 1.1255
R12633 VDAC_N.n929 VDAC_N.t2105 1.1255
R12634 VDAC_N.n930 VDAC_N.t440 1.1255
R12635 VDAC_N.n931 VDAC_N.t1998 1.1255
R12636 VDAC_N.n932 VDAC_N.t1232 1.1255
R12637 VDAC_N.n933 VDAC_N.t1562 1.1255
R12638 VDAC_N.n934 VDAC_N.t1367 1.1255
R12639 VDAC_N.n935 VDAC_N.t1326 1.1255
R12640 VDAC_N.n103 VDAC_N.t562 1.1255
R12641 VDAC_N.n936 VDAC_N.t2019 1.1255
R12642 VDAC_N.n937 VDAC_N.t456 1.1255
R12643 VDAC_N.n938 VDAC_N.t499 1.1255
R12644 VDAC_N.n939 VDAC_N.t884 1.1255
R12645 VDAC_N.n940 VDAC_N.t1362 1.1255
R12646 VDAC_N.n941 VDAC_N.t1644 1.1255
R12647 VDAC_N.n942 VDAC_N.t310 1.1255
R12648 VDAC_N.n943 VDAC_N.t2086 1.1255
R12649 VDAC_N.n944 VDAC_N.t488 1.1255
R12650 VDAC_N.n945 VDAC_N.t950 1.1255
R12651 VDAC_N.n946 VDAC_N.t516 1.1255
R12652 VDAC_N.n947 VDAC_N.t838 1.1255
R12653 VDAC_N.n948 VDAC_N.t33 1.1255
R12654 VDAC_N.n949 VDAC_N.t1855 1.1255
R12655 VDAC_N.n950 VDAC_N.t1204 1.1255
R12656 VDAC_N.n951 VDAC_N.t386 1.1255
R12657 VDAC_N.n952 VDAC_N.t188 1.1255
R12658 VDAC_N.n953 VDAC_N.t280 1.1255
R12659 VDAC_N.n954 VDAC_N.t1099 1.1255
R12660 VDAC_N.n955 VDAC_N.t1616 1.1255
R12661 VDAC_N.n956 VDAC_N.t1742 1.1255
R12662 VDAC_N.n957 VDAC_N.t1184 1.1255
R12663 VDAC_N.n958 VDAC_N.t1534 1.1255
R12664 VDAC_N.n959 VDAC_N.t331 1.1255
R12665 VDAC_N.n960 VDAC_N.t294 1.1255
R12666 VDAC_N.n961 VDAC_N.t579 1.1255
R12667 VDAC_N.n962 VDAC_N.t1597 1.1255
R12668 VDAC_N.n963 VDAC_N.t474 1.1255
R12669 VDAC_N.n964 VDAC_N.t757 1.1255
R12670 VDAC_N.n965 VDAC_N.t126 1.1255
R12671 VDAC_N.n966 VDAC_N.t1271 1.1255
R12672 VDAC_N.n967 VDAC_N.t255 1.1255
R12673 VDAC_N.n968 VDAC_N.t1163 1.1255
R12674 VDAC_N.n969 VDAC_N.t1625 1.1255
R12675 VDAC_N.n970 VDAC_N.t2085 1.1255
R12676 VDAC_N.n971 VDAC_N.t121 1.1255
R12677 VDAC_N.n972 VDAC_N.t1001 1.1255
R12678 VDAC_N.n973 VDAC_N.t347 1.1255
R12679 VDAC_N.n974 VDAC_N.t1871 1.1255
R12680 VDAC_N.n975 VDAC_N.t692 1.1255
R12681 VDAC_N.n976 VDAC_N.t135 1.1255
R12682 VDAC_N.n977 VDAC_N.t1140 1.1255
R12683 VDAC_N.n978 VDAC_N.t1238 1.1255
R12684 VDAC_N.n979 VDAC_N.t157 1.1255
R12685 VDAC_N.n980 VDAC_N.t816 1.1255
R12686 VDAC_N.n981 VDAC_N.t994 1.1255
R12687 VDAC_N.n982 VDAC_N.t1160 1.1255
R12688 VDAC_N.n983 VDAC_N.t1530 1.1255
R12689 VDAC_N.n984 VDAC_N.t1412 1.1255
R12690 VDAC_N.n985 VDAC_N.t186 1.1255
R12691 VDAC_N.n986 VDAC_N.t1127 1.1255
R12692 VDAC_N.n987 VDAC_N.t2128 1.1255
R12693 VDAC_N.n988 VDAC_N.t2018 1.1255
R12694 VDAC_N.n989 VDAC_N.t755 1.1255
R12695 VDAC_N.n990 VDAC_N.t1594 1.1255
R12696 VDAC_N.n991 VDAC_N.t1379 1.1255
R12697 VDAC_N.n992 VDAC_N.t686 1.1255
R12698 VDAC_N.n993 VDAC_N.t1161 1.1255
R12699 VDAC_N.n994 VDAC_N.t453 1.1255
R12700 VDAC_N.n995 VDAC_N.t2070 1.1255
R12701 VDAC_N.n996 VDAC_N.t771 1.1255
R12702 VDAC_N.n997 VDAC_N.t2081 1.1255
R12703 VDAC_N.n998 VDAC_N.t373 1.1255
R12704 VDAC_N.n102 VDAC_N.t1921 1.1255
R12705 VDAC_N.n999 VDAC_N.t637 1.1255
R12706 VDAC_N.n1000 VDAC_N.t921 1.1255
R12707 VDAC_N.n1001 VDAC_N.t1135 1.1255
R12708 VDAC_N.n1002 VDAC_N.t1601 1.1255
R12709 VDAC_N.n1003 VDAC_N.t1043 1.1255
R12710 VDAC_N.n1004 VDAC_N.t211 1.1255
R12711 VDAC_N.n1005 VDAC_N.t1943 1.1255
R12712 VDAC_N.n1006 VDAC_N.t532 1.1255
R12713 VDAC_N.n1007 VDAC_N.t939 1.1255
R12714 VDAC_N.n1008 VDAC_N.t580 1.1255
R12715 VDAC_N.n1009 VDAC_N.t429 1.1255
R12716 VDAC_N.n1010 VDAC_N.t1084 1.1255
R12717 VDAC_N.n1011 VDAC_N.t2024 1.1255
R12718 VDAC_N.n1012 VDAC_N.t1663 1.1255
R12719 VDAC_N.n1013 VDAC_N.t1075 1.1255
R12720 VDAC_N.n1014 VDAC_N.t1080 1.1255
R12721 VDAC_N.n1015 VDAC_N.t523 1.1255
R12722 VDAC_N.n1016 VDAC_N.t1280 1.1255
R12723 VDAC_N.n1017 VDAC_N.t1798 1.1255
R12724 VDAC_N.n1018 VDAC_N.t1652 1.1255
R12725 VDAC_N.n1019 VDAC_N.t1346 1.1255
R12726 VDAC_N.n1020 VDAC_N.t1548 1.1255
R12727 VDAC_N.n1021 VDAC_N.t586 1.1255
R12728 VDAC_N.n1022 VDAC_N.t1050 1.1255
R12729 VDAC_N.n1023 VDAC_N.t704 1.1255
R12730 VDAC_N.n1024 VDAC_N.t1854 1.1255
R12731 VDAC_N.n1025 VDAC_N.t1409 1.1255
R12732 VDAC_N.n1026 VDAC_N.t374 1.1255
R12733 VDAC_N.n1027 VDAC_N.t1297 1.1255
R12734 VDAC_N.n1028 VDAC_N.t614 1.1255
R12735 VDAC_N.n1029 VDAC_N.t13 1.1255
R12736 VDAC_N.n1030 VDAC_N.t841 1.1255
R12737 VDAC_N.n1031 VDAC_N.t1926 1.1255
R12738 VDAC_N.n1032 VDAC_N.t1433 1.1255
R12739 VDAC_N.n1033 VDAC_N.t1895 1.1255
R12740 VDAC_N.n1034 VDAC_N.t1329 1.1255
R12741 VDAC_N.n1035 VDAC_N.t1787 1.1255
R12742 VDAC_N.n1036 VDAC_N.t567 1.1255
R12743 VDAC_N.n1037 VDAC_N.t855 1.1255
R12744 VDAC_N.n1038 VDAC_N.t1371 1.1255
R12745 VDAC_N.n1039 VDAC_N.t1547 1.1255
R12746 VDAC_N.n1040 VDAC_N.t1071 1.1255
R12747 VDAC_N.n1041 VDAC_N.t864 1.1255
R12748 VDAC_N.n1042 VDAC_N.t145 1.1255
R12749 VDAC_N.n1043 VDAC_N.t228 1.1255
R12750 VDAC_N.n1044 VDAC_N.t802 1.1255
R12751 VDAC_N.n1045 VDAC_N.t1452 1.1255
R12752 VDAC_N.n1046 VDAC_N.t1138 1.1255
R12753 VDAC_N.n1047 VDAC_N.t9 1.1255
R12754 VDAC_N.n1048 VDAC_N.t56 1.1255
R12755 VDAC_N.n1049 VDAC_N.t1846 1.1255
R12756 VDAC_N.n1050 VDAC_N.t360 1.1255
R12757 VDAC_N.n1051 VDAC_N.t1630 1.1255
R12758 VDAC_N.n1052 VDAC_N.t1293 1.1255
R12759 VDAC_N.n1053 VDAC_N.t1198 1.1255
R12760 VDAC_N.n1054 VDAC_N.t605 1.1255
R12761 VDAC_N.n1055 VDAC_N.t1920 1.1255
R12762 VDAC_N.n1056 VDAC_N.t1922 1.1255
R12763 VDAC_N.n1057 VDAC_N.t1539 1.1255
R12764 VDAC_N.n1058 VDAC_N.t1686 1.1255
R12765 VDAC_N.n1059 VDAC_N.t1327 1.1255
R12766 VDAC_N.n1060 VDAC_N.t261 1.1255
R12767 VDAC_N.n1061 VDAC_N.t1215 1.1255
R12768 VDAC_N.n101 VDAC_N.t1786 1.1255
R12769 VDAC_N.n1062 VDAC_N.t820 1.1255
R12770 VDAC_N.n1063 VDAC_N.t1574 1.1255
R12771 VDAC_N.n1064 VDAC_N.t204 1.1255
R12772 VDAC_N.n1065 VDAC_N.t582 1.1255
R12773 VDAC_N.n1066 VDAC_N.t1046 1.1255
R12774 VDAC_N.n1067 VDAC_N.t1816 1.1255
R12775 VDAC_N.n1068 VDAC_N.t482 1.1255
R12776 VDAC_N.n1069 VDAC_N.t1405 1.1255
R12777 VDAC_N.n1070 VDAC_N.t78 1.1255
R12778 VDAC_N.n1071 VDAC_N.t107 1.1255
R12779 VDAC_N.n1072 VDAC_N.t174 1.1255
R12780 VDAC_N.n1073 VDAC_N.t37 1.1255
R12781 VDAC_N.n1074 VDAC_N.t839 1.1255
R12782 VDAC_N.n1075 VDAC_N.t1780 1.1255
R12783 VDAC_N.n1076 VDAC_N.t1378 1.1255
R12784 VDAC_N.n1077 VDAC_N.t653 1.1255
R12785 VDAC_N.n1078 VDAC_N.t1166 1.1255
R12786 VDAC_N.n1079 VDAC_N.t2094 1.1255
R12787 VDAC_N.n1080 VDAC_N.t229 1.1255
R12788 VDAC_N.n1081 VDAC_N.t86 1.1255
R12789 VDAC_N.n1082 VDAC_N.t723 1.1255
R12790 VDAC_N.n1083 VDAC_N.t1662 1.1255
R12791 VDAC_N.n1084 VDAC_N.t349 1.1255
R12792 VDAC_N.n1085 VDAC_N.t1767 1.1255
R12793 VDAC_N.n1086 VDAC_N.t1085 1.1255
R12794 VDAC_N.n1087 VDAC_N.t437 1.1255
R12795 VDAC_N.n1088 VDAC_N.t159 1.1255
R12796 VDAC_N.n1089 VDAC_N.t1449 1.1255
R12797 VDAC_N.n1090 VDAC_N.t1019 1.1255
R12798 VDAC_N.n1091 VDAC_N.t357 1.1255
R12799 VDAC_N.n1092 VDAC_N.t1799 1.1255
R12800 VDAC_N.n1093 VDAC_N.t852 1.1255
R12801 VDAC_N.n1094 VDAC_N.t863 1.1255
R12802 VDAC_N.n1095 VDAC_N.t860 1.1255
R12803 VDAC_N.n1096 VDAC_N.t936 1.1255
R12804 VDAC_N.n1097 VDAC_N.t2043 1.1255
R12805 VDAC_N.n1098 VDAC_N.t368 1.1255
R12806 VDAC_N.n1099 VDAC_N.t929 1.1255
R12807 VDAC_N.n1100 VDAC_N.t1892 1.1255
R12808 VDAC_N.n1101 VDAC_N.t1414 1.1255
R12809 VDAC_N.n1102 VDAC_N.t844 1.1255
R12810 VDAC_N.n1103 VDAC_N.t1358 1.1255
R12811 VDAC_N.n1104 VDAC_N.t597 1.1255
R12812 VDAC_N.n1105 VDAC_N.t1872 1.1255
R12813 VDAC_N.n1106 VDAC_N.t490 1.1255
R12814 VDAC_N.n1107 VDAC_N.t401 1.1255
R12815 VDAC_N.n1108 VDAC_N.t1650 1.1255
R12816 VDAC_N.n1109 VDAC_N.t669 1.1255
R12817 VDAC_N.n1110 VDAC_N.t726 1.1255
R12818 VDAC_N.n1111 VDAC_N.t101 1.1255
R12819 VDAC_N.n1112 VDAC_N.t1661 1.1255
R12820 VDAC_N.n1113 VDAC_N.t25 1.1255
R12821 VDAC_N.n1114 VDAC_N.t789 1.1255
R12822 VDAC_N.n1115 VDAC_N.t1017 1.1255
R12823 VDAC_N.n1116 VDAC_N.t685 1.1255
R12824 VDAC_N.n1117 VDAC_N.t1903 1.1255
R12825 VDAC_N.n1118 VDAC_N.t1227 1.1255
R12826 VDAC_N.n1119 VDAC_N.t445 1.1255
R12827 VDAC_N.n1120 VDAC_N.t1516 1.1255
R12828 VDAC_N.n1121 VDAC_N.t125 1.1255
R12829 VDAC_N.n1122 VDAC_N.t2041 1.1255
R12830 VDAC_N.n1123 VDAC_N.t480 1.1255
R12831 VDAC_N.n1124 VDAC_N.t1929 1.1255
R12832 VDAC_N.n100 VDAC_N.t76 1.1255
R12833 VDAC_N.n1125 VDAC_N.t1587 1.1255
R12834 VDAC_N.n1126 VDAC_N.t1628 1.1255
R12835 VDAC_N.n1127 VDAC_N.t209 1.1255
R12836 VDAC_N.n1128 VDAC_N.t981 1.1255
R12837 VDAC_N.n1129 VDAC_N.t1908 1.1255
R12838 VDAC_N.n1130 VDAC_N.t1833 1.1255
R12839 VDAC_N.n1131 VDAC_N.t1004 1.1255
R12840 VDAC_N.n1132 VDAC_N.t102 1.1255
R12841 VDAC_N.n1133 VDAC_N.t1078 1.1255
R12842 VDAC_N.n1134 VDAC_N.t1960 1.1255
R12843 VDAC_N.n1135 VDAC_N.t1961 1.1255
R12844 VDAC_N.n1136 VDAC_N.t1512 1.1255
R12845 VDAC_N.n1137 VDAC_N.t238 1.1255
R12846 VDAC_N.n1138 VDAC_N.t2130 1.1255
R12847 VDAC_N.n1139 VDAC_N.t1008 1.1255
R12848 VDAC_N.n1140 VDAC_N.t27 1.1255
R12849 VDAC_N.n1141 VDAC_N.t1536 1.1255
R12850 VDAC_N.n1142 VDAC_N.t450 1.1255
R12851 VDAC_N.n1143 VDAC_N.t1445 1.1255
R12852 VDAC_N.n1144 VDAC_N.t1494 1.1255
R12853 VDAC_N.n1145 VDAC_N.t103 1.1255
R12854 VDAC_N.n1146 VDAC_N.t1278 1.1255
R12855 VDAC_N.n1147 VDAC_N.t1115 1.1255
R12856 VDAC_N.n1148 VDAC_N.t1581 1.1255
R12857 VDAC_N.n1149 VDAC_N.t1770 1.1255
R12858 VDAC_N.n1150 VDAC_N.t1469 1.1255
R12859 VDAC_N.n1151 VDAC_N.t979 1.1255
R12860 VDAC_N.n1152 VDAC_N.t335 1.1255
R12861 VDAC_N.n1153 VDAC_N.t1827 1.1255
R12862 VDAC_N.n1154 VDAC_N.t1147 1.1255
R12863 VDAC_N.n1155 VDAC_N.t1609 1.1255
R12864 VDAC_N.n1156 VDAC_N.t2126 1.1255
R12865 VDAC_N.n1157 VDAC_N.t1501 1.1255
R12866 VDAC_N.n1158 VDAC_N.t509 1.1255
R12867 VDAC_N.n1159 VDAC_N.t2116 1.1255
R12868 VDAC_N.n1160 VDAC_N.t485 1.1255
R12869 VDAC_N.n1161 VDAC_N.t628 1.1255
R12870 VDAC_N.n1162 VDAC_N.t1643 1.1255
R12871 VDAC_N.n1163 VDAC_N.t700 1.1255
R12872 VDAC_N.n1164 VDAC_N.t1040 1.1255
R12873 VDAC_N.n1165 VDAC_N.t2135 1.1255
R12874 VDAC_N.n1166 VDAC_N.t1952 1.1255
R12875 VDAC_N.n1167 VDAC_N.t982 1.1255
R12876 VDAC_N.n1168 VDAC_N.t560 1.1255
R12877 VDAC_N.n1169 VDAC_N.t1486 1.1255
R12878 VDAC_N.n1170 VDAC_N.t681 1.1255
R12879 VDAC_N.n1171 VDAC_N.t646 1.1255
R12880 VDAC_N.n1172 VDAC_N.t1111 1.1255
R12881 VDAC_N.n1173 VDAC_N.t2072 1.1255
R12882 VDAC_N.n1174 VDAC_N.t1994 1.1255
R12883 VDAC_N.n1175 VDAC_N.t747 1.1255
R12884 VDAC_N.n1176 VDAC_N.t82 1.1255
R12885 VDAC_N.n1177 VDAC_N.t1365 1.1255
R12886 VDAC_N.n1178 VDAC_N.t1821 1.1255
R12887 VDAC_N.n1179 VDAC_N.t307 1.1255
R12888 VDAC_N.n1180 VDAC_N.t1711 1.1255
R12889 VDAC_N.n1181 VDAC_N.t1034 1.1255
R12890 VDAC_N.n1182 VDAC_N.t763 1.1255
R12891 VDAC_N.n1183 VDAC_N.t1047 1.1255
R12892 VDAC_N.n1184 VDAC_N.t369 1.1255
R12893 VDAC_N.n1185 VDAC_N.t941 1.1255
R12894 VDAC_N.n1186 VDAC_N.t2100 1.1255
R12895 VDAC_N.n1187 VDAC_N.t1743 1.1255
R12896 VDAC_N.n99 VDAC_N.t1487 1.1255
R12897 VDAC_N.n1188 VDAC_N.t1598 1.1255
R12898 VDAC_N.n1189 VDAC_N.t705 1.1255
R12899 VDAC_N.n1190 VDAC_N.t690 1.1255
R12900 VDAC_N.n1191 VDAC_N.t99 1.1255
R12901 VDAC_N.n1192 VDAC_N.t827 1.1255
R12902 VDAC_N.n1193 VDAC_N.t542 1.1255
R12903 VDAC_N.n1194 VDAC_N.t773 1.1255
R12904 VDAC_N.n1195 VDAC_N.t515 1.1255
R12905 VDAC_N.n1196 VDAC_N.t721 1.1255
R12906 VDAC_N.n1197 VDAC_N.t951 1.1255
R12907 VDAC_N.n1198 VDAC_N.t1193 1.1255
R12908 VDAC_N.n1199 VDAC_N.t461 1.1255
R12909 VDAC_N.n1200 VDAC_N.t2108 1.1255
R12910 VDAC_N.n1201 VDAC_N.t1011 1.1255
R12911 VDAC_N.n1202 VDAC_N.t1224 1.1255
R12912 VDAC_N.n1203 VDAC_N.t894 1.1255
R12913 VDAC_N.n1204 VDAC_N.t1508 1.1255
R12914 VDAC_N.n1205 VDAC_N.t1322 1.1255
R12915 VDAC_N.n1206 VDAC_N.t1251 1.1255
R12916 VDAC_N.n1207 VDAC_N.t1110 1.1255
R12917 VDAC_N.n1208 VDAC_N.t2042 1.1255
R12918 VDAC_N.n1209 VDAC_N.t904 1.1255
R12919 VDAC_N.n1210 VDAC_N.t926 1.1255
R12920 VDAC_N.n1211 VDAC_N.t1393 1.1255
R12921 VDAC_N.n1212 VDAC_N.t366 1.1255
R12922 VDAC_N.n1213 VDAC_N.t1279 1.1255
R12923 VDAC_N.n1214 VDAC_N.t457 1.1255
R12924 VDAC_N.n1215 VDAC_N.t1062 1.1255
R12925 VDAC_N.n1216 VDAC_N.t1637 1.1255
R12926 VDAC_N.n1217 VDAC_N.t1886 1.1255
R12927 VDAC_N.n1218 VDAC_N.t1419 1.1255
R12928 VDAC_N.n1219 VDAC_N.t517 1.1255
R12929 VDAC_N.n1220 VDAC_N.t1313 1.1255
R12930 VDAC_N.n1221 VDAC_N.t463 1.1255
R12931 VDAC_N.n1222 VDAC_N.t1164 1.1255
R12932 VDAC_N.n1223 VDAC_N.t1665 1.1255
R12933 VDAC_N.n1224 VDAC_N.t2125 1.1255
R12934 VDAC_N.n1225 VDAC_N.t739 1.1255
R12935 VDAC_N.n1226 VDAC_N.t2011 1.1255
R12936 VDAC_N.n1227 VDAC_N.t1288 1.1255
R12937 VDAC_N.n1228 VDAC_N.t1887 1.1255
R12938 VDAC_N.n1229 VDAC_N.t1192 1.1255
R12939 VDAC_N.n1230 VDAC_N.t1542 1.1255
R12940 VDAC_N.n1231 VDAC_N.t620 1.1255
R12941 VDAC_N.n1232 VDAC_N.t1102 1.1255
R12942 VDAC_N.n1233 VDAC_N.t581 1.1255
R12943 VDAC_N.n1234 VDAC_N.t1744 1.1255
R12944 VDAC_N.n1235 VDAC_N.t1814 1.1255
R12945 VDAC_N.n1236 VDAC_N.t664 1.1255
R12946 VDAC_N.n1237 VDAC_N.t1606 1.1255
R12947 VDAC_N.n1238 VDAC_N.t1273 1.1255
R12948 VDAC_N.n1239 VDAC_N.t694 1.1255
R12949 VDAC_N.n1240 VDAC_N.t1167 1.1255
R12950 VDAC_N.n1241 VDAC_N.t1631 1.1255
R12951 VDAC_N.n1242 VDAC_N.t1878 1.1255
R12952 VDAC_N.n1243 VDAC_N.t1521 1.1255
R12953 VDAC_N.n1244 VDAC_N.t434 1.1255
R12954 VDAC_N.n1245 VDAC_N.t1311 1.1255
R12955 VDAC_N.n1246 VDAC_N.t1879 1.1255
R12956 VDAC_N.n1247 VDAC_N.t1197 1.1255
R12957 VDAC_N.n1248 VDAC_N.t845 1.1255
R12958 VDAC_N.n1249 VDAC_N.t1132 1.1255
R12959 VDAC_N.n1250 VDAC_N.t1551 1.1255
R12960 VDAC_N.n98 VDAC_N.t472 1.1255
R12961 VDAC_N.n1251 VDAC_N.t265 1.1255
R12962 VDAC_N.n1252 VDAC_N.t192 1.1255
R12963 VDAC_N.n1253 VDAC_N.t923 1.1255
R12964 VDAC_N.n1254 VDAC_N.t940 1.1255
R12965 VDAC_N.n1255 VDAC_N.t1186 1.1255
R12966 VDAC_N.n1256 VDAC_N.t16 1.1255
R12967 VDAC_N.n1257 VDAC_N.t1912 1.1255
R12968 VDAC_N.n1258 VDAC_N.t498 1.1255
R12969 VDAC_N.n1259 VDAC_N.t744 1.1255
R12970 VDAC_N.n1260 VDAC_N.t854 1.1255
R12971 VDAC_N.n1261 VDAC_N.t1188 1.1255
R12972 VDAC_N.n1262 VDAC_N.t1450 1.1255
R12973 VDAC_N.n1263 VDAC_N.t65 1.1255
R12974 VDAC_N.n1264 VDAC_N.t1142 1.1255
R12975 VDAC_N.n1265 VDAC_N.t538 1.1255
R12976 VDAC_N.n1266 VDAC_N.t1619 1.1255
R12977 VDAC_N.n1267 VDAC_N.t142 1.1255
R12978 VDAC_N.n1268 VDAC_N.t1407 1.1255
R12979 VDAC_N.n1269 VDAC_N.t513 1.1255
R12980 VDAC_N.n1270 VDAC_N.t345 1.1255
R12981 VDAC_N.n1271 VDAC_N.t1757 1.1255
R12982 VDAC_N.n1272 VDAC_N.t1185 1.1255
R12983 VDAC_N.n1273 VDAC_N.t1653 1.1255
R12984 VDAC_N.n1274 VDAC_N.t2107 1.1255
R12985 VDAC_N.n1275 VDAC_N.t379 1.1255
R12986 VDAC_N.n1276 VDAC_N.t1997 1.1255
R12987 VDAC_N.n1277 VDAC_N.t1240 1.1255
R12988 VDAC_N.n1278 VDAC_N.t907 1.1255
R12989 VDAC_N.n1279 VDAC_N.t1556 1.1255
R12990 VDAC_N.n1280 VDAC_N.t1681 1.1255
R12991 VDAC_N.n1281 VDAC_N.t1417 1.1255
R12992 VDAC_N.n1282 VDAC_N.t1122 1.1255
R12993 VDAC_N.n1283 VDAC_N.t1029 1.1255
R12994 VDAC_N.n1284 VDAC_N.t680 1.1255
R12995 VDAC_N.n1285 VDAC_N.t426 1.1255
R12996 VDAC_N.n1286 VDAC_N.t1796 1.1255
R12997 VDAC_N.n1287 VDAC_N.t198 1.1255
R12998 VDAC_N.n1288 VDAC_N.t796 1.1255
R12999 VDAC_N.n1289 VDAC_N.t1170 1.1255
R13000 VDAC_N.n1290 VDAC_N.t2102 1.1255
R13001 VDAC_N.n1291 VDAC_N.t920 1.1255
R13002 VDAC_N.n1292 VDAC_N.t2054 1.1255
R13003 VDAC_N.n1293 VDAC_N.t213 1.1255
R13004 VDAC_N.n1294 VDAC_N.t1626 1.1255
R13005 VDAC_N.n1295 VDAC_N.t1291 1.1255
R13006 VDAC_N.n1296 VDAC_N.t1861 1.1255
R13007 VDAC_N.n1297 VDAC_N.t1179 1.1255
R13008 VDAC_N.n1298 VDAC_N.t1649 1.1255
R13009 VDAC_N.n1299 VDAC_N.t158 1.1255
R13010 VDAC_N.n1300 VDAC_N.t1537 1.1255
R13011 VDAC_N.n1301 VDAC_N.t519 1.1255
R13012 VDAC_N.n1302 VDAC_N.t727 1.1255
R13013 VDAC_N.n1303 VDAC_N.t959 1.1255
R13014 VDAC_N.n1304 VDAC_N.t212 1.1255
R13015 VDAC_N.n1305 VDAC_N.t853 1.1255
R13016 VDAC_N.n1306 VDAC_N.t1292 1.1255
R13017 VDAC_N.n1307 VDAC_N.t31 1.1255
R13018 VDAC_N.n1308 VDAC_N.t1027 1.1255
R13019 VDAC_N.n1309 VDAC_N.t464 1.1255
R13020 VDAC_N.n1310 VDAC_N.t87 1.1255
R13021 VDAC_N.n1311 VDAC_N.t900 1.1255
R13022 VDAC_N.n1312 VDAC_N.t1614 1.1255
R13023 VDAC_N.n1313 VDAC_N.t1708 1.1255
R13024 VDAC_N.n97 VDAC_N.t253 1.1255
R13025 VDAC_N.n1314 VDAC_N.t1151 1.1255
R13026 VDAC_N.n1315 VDAC_N.t239 1.1255
R13027 VDAC_N.n1316 VDAC_N.t534 1.1255
R13028 VDAC_N.n1317 VDAC_N.t397 1.1255
R13029 VDAC_N.n1318 VDAC_N.t269 1.1255
R13030 VDAC_N.n1319 VDAC_N.t1401 1.1255
R13031 VDAC_N.n1320 VDAC_N.t943 1.1255
R13032 VDAC_N.n1321 VDAC_N.t1252 1.1255
R13033 VDAC_N.n1322 VDAC_N.t459 1.1255
R13034 VDAC_N.n1323 VDAC_N.t124 1.1255
R13035 VDAC_N.n1324 VDAC_N.t1535 1.1255
R13036 VDAC_N.n1325 VDAC_N.t1063 1.1255
R13037 VDAC_N.n1326 VDAC_N.t1648 1.1255
R13038 VDAC_N.n1327 VDAC_N.t1472 1.1255
R13039 VDAC_N.n1328 VDAC_N.t442 1.1255
R13040 VDAC_N.n1329 VDAC_N.t1427 1.1255
R13041 VDAC_N.n1330 VDAC_N.t1458 1.1255
R13042 VDAC_N.n1331 VDAC_N.t621 1.1255
R13043 VDAC_N.n1332 VDAC_N.t1781 1.1255
R13044 VDAC_N.n1333 VDAC_N.t563 1.1255
R13045 VDAC_N.n1334 VDAC_N.t1565 1.1255
R13046 VDAC_N.n1335 VDAC_N.t514 1.1255
R13047 VDAC_N.n1336 VDAC_N.t743 1.1255
R13048 VDAC_N.n1337 VDAC_N.t1917 1.1255
R13049 VDAC_N.n1338 VDAC_N.t1239 1.1255
R13050 VDAC_N.n1339 VDAC_N.t1811 1.1255
R13051 VDAC_N.n1340 VDAC_N.t876 1.1255
R13052 VDAC_N.n1341 VDAC_N.t77 1.1255
R13053 VDAC_N.n1342 VDAC_N.t1436 1.1255
R13054 VDAC_N.n1343 VDAC_N.t1485 1.1255
R13055 VDAC_N.n1344 VDAC_N.t267 1.1255
R13056 VDAC_N.n1345 VDAC_N.t1440 1.1255
R13057 VDAC_N.n1346 VDAC_N.t1843 1.1255
R13058 VDAC_N.n1347 VDAC_N.t2124 1.1255
R13059 VDAC_N.n1348 VDAC_N.t178 1.1255
R13060 VDAC_N.n1349 VDAC_N.t1052 1.1255
R13061 VDAC_N.n1350 VDAC_N.t1016 1.1255
R13062 VDAC_N.n1351 VDAC_N.t1973 1.1255
R13063 VDAC_N.n1352 VDAC_N.t792 1.1255
R13064 VDAC_N.n1353 VDAC_N.t1726 1.1255
R13065 VDAC_N.n1354 VDAC_N.t2052 1.1255
R13066 VDAC_N.n1355 VDAC_N.t438 1.1255
R13067 VDAC_N.n1356 VDAC_N.t673 1.1255
R13068 VDAC_N.n1357 VDAC_N.t1234 1.1255
R13069 VDAC_N.n1358 VDAC_N.t1093 1.1255
R13070 VDAC_N.n1359 VDAC_N.t1669 1.1255
R13071 VDAC_N.n1360 VDAC_N.t510 1.1255
R13072 VDAC_N.n1361 VDAC_N.t1453 1.1255
R13073 VDAC_N.n1362 VDAC_N.t1734 1.1255
R13074 VDAC_N.n1363 VDAC_N.t1351 1.1255
R13075 VDAC_N.n1364 VDAC_N.t139 1.1255
R13076 VDAC_N.n1365 VDAC_N.t631 1.1255
R13077 VDAC_N.n1366 VDAC_N.t865 1.1255
R13078 VDAC_N.n1367 VDAC_N.t1244 1.1255
R13079 VDAC_N.n1368 VDAC_N.t1481 1.1255
R13080 VDAC_N.n1369 VDAC_N.t2049 1.1255
R13081 VDAC_N.n1370 VDAC_N.t703 1.1255
R13082 VDAC_N.n1371 VDAC_N.t933 1.1255
R13083 VDAC_N.n1372 VDAC_N.t1956 1.1255
R13084 VDAC_N.n1373 VDAC_N.t1727 1.1255
R13085 VDAC_N.n1374 VDAC_N.t1564 1.1255
R13086 VDAC_N.n1375 VDAC_N.t1218 1.1255
R13087 VDAC_N.n1376 VDAC_N.t541 1.1255
R13088 VDAC_N.n96 VDAC_N.t814 1.1255
R13089 VDAC_N.n1377 VDAC_N.t428 1.1255
R13090 VDAC_N.n1378 VDAC_N.t194 1.1255
R13091 VDAC_N.n1379 VDAC_N.t348 1.1255
R13092 VDAC_N.n1380 VDAC_N.t1864 1.1255
R13093 VDAC_N.n1381 VDAC_N.t258 1.1255
R13094 VDAC_N.n1382 VDAC_N.t1408 1.1255
R13095 VDAC_N.n1383 VDAC_N.t1646 1.1255
R13096 VDAC_N.n1384 VDAC_N.t667 1.1255
R13097 VDAC_N.n1385 VDAC_N.t1418 1.1255
R13098 VDAC_N.n1386 VDAC_N.t611 1.1255
R13099 VDAC_N.n1387 VDAC_N.t1984 1.1255
R13100 VDAC_N.n1388 VDAC_N.t21 1.1255
R13101 VDAC_N.n1389 VDAC_N.t123 1.1255
R13102 VDAC_N.n1390 VDAC_N.t1113 1.1255
R13103 VDAC_N.n1391 VDAC_N.t803 1.1255
R13104 VDAC_N.n1392 VDAC_N.t550 1.1255
R13105 VDAC_N.n1393 VDAC_N.t73 1.1255
R13106 VDAC_N.n1394 VDAC_N.t1927 1.1255
R13107 VDAC_N.n1395 VDAC_N.t112 1.1255
R13108 VDAC_N.n1396 VDAC_N.t477 1.1255
R13109 VDAC_N.n1397 VDAC_N.t1900 1.1255
R13110 VDAC_N.n1398 VDAC_N.t871 1.1255
R13111 VDAC_N.n1399 VDAC_N.t22 1.1255
R13112 VDAC_N.n1400 VDAC_N.t1928 1.1255
R13113 VDAC_N.n1401 VDAC_N.t1951 1.1255
R13114 VDAC_N.n1402 VDAC_N.t1480 1.1255
R13115 VDAC_N.n1403 VDAC_N.t1690 1.1255
R13116 VDAC_N.n1404 VDAC_N.t324 1.1255
R13117 VDAC_N.n1405 VDAC_N.t1466 1.1255
R13118 VDAC_N.n1406 VDAC_N.t1340 1.1255
R13119 VDAC_N.n1407 VDAC_N.t2048 1.1255
R13120 VDAC_N.n1408 VDAC_N.t1103 1.1255
R13121 VDAC_N.n1409 VDAC_N.t1624 1.1255
R13122 VDAC_N.n1410 VDAC_N.t886 1.1255
R13123 VDAC_N.n1411 VDAC_N.t1359 1.1255
R13124 VDAC_N.n1412 VDAC_N.t782 1.1255
R13125 VDAC_N.n1413 VDAC_N.t635 1.1255
R13126 VDAC_N.n1414 VDAC_N.t1094 1.1255
R13127 VDAC_N.n1415 VDAC_N.t1131 1.1255
R13128 VDAC_N.n1416 VDAC_N.t813 1.1255
R13129 VDAC_N.n1417 VDAC_N.t518 1.1255
R13130 VDAC_N.n1418 VDAC_N.t1571 1.1255
R13131 VDAC_N.n1419 VDAC_N.t1031 1.1255
R13132 VDAC_N.n1420 VDAC_N.t1363 1.1255
R13133 VDAC_N.n1421 VDAC_N.t1819 1.1255
R13134 VDAC_N.n1422 VDAC_N.t1828 1.1255
R13135 VDAC_N.n1423 VDAC_N.t1709 1.1255
R13136 VDAC_N.n1424 VDAC_N.t14 1.1255
R13137 VDAC_N.n1425 VDAC_N.t225 1.1255
R13138 VDAC_N.n1426 VDAC_N.t1045 1.1255
R13139 VDAC_N.n1427 VDAC_N.t1464 1.1255
R13140 VDAC_N.n1428 VDAC_N.t1947 1.1255
R13141 VDAC_N.n1429 VDAC_N.t2084 1.1255
R13142 VDAC_N.n1430 VDAC_N.t1454 1.1255
R13143 VDAC_N.n1431 VDAC_N.t636 1.1255
R13144 VDAC_N.n1432 VDAC_N.t66 1.1255
R13145 VDAC_N.n1433 VDAC_N.t2093 1.1255
R13146 VDAC_N.n1434 VDAC_N.t1608 1.1255
R13147 VDAC_N.n1435 VDAC_N.t998 1.1255
R13148 VDAC_N.n1436 VDAC_N.t600 1.1255
R13149 VDAC_N.n1437 VDAC_N.t122 1.1255
R13150 VDAC_N.n1438 VDAC_N.t1355 1.1255
R13151 VDAC_N.n1439 VDAC_N.t1298 1.1255
R13152 VDAC_N.n95 VDAC_N.t1820 1.1255
R13153 VDAC_N.n1440 VDAC_N.t1491 1.1255
R13154 VDAC_N.n1441 VDAC_N.t2057 1.1255
R13155 VDAC_N.n1442 VDAC_N.t707 1.1255
R13156 VDAC_N.n1443 VDAC_N.t1849 1.1255
R13157 VDAC_N.n1444 VDAC_N.t1124 1.1255
R13158 VDAC_N.n1445 VDAC_N.t1737 1.1255
R13159 VDAC_N.n1446 VDAC_N.t2076 1.1255
R13160 VDAC_N.n1447 VDAC_N.t2016 1.1255
R13161 VDAC_N.n1448 VDAC_N.t1059 1.1255
R13162 VDAC_N.n1449 VDAC_N.t416 1.1255
R13163 VDAC_N.n1450 VDAC_N.t953 1.1255
R13164 VDAC_N.n1451 VDAC_N.t168 1.1255
R13165 VDAC_N.n1452 VDAC_N.t774 1.1255
R13166 VDAC_N.n1453 VDAC_N.t1822 1.1255
R13167 VDAC_N.n1454 VDAC_N.t1391 1.1255
R13168 VDAC_N.n1455 VDAC_N.t43 1.1255
R13169 VDAC_N.n1456 VDAC_N.t1277 1.1255
R13170 VDAC_N.n1457 VDAC_N.t885 1.1255
R13171 VDAC_N.n1458 VDAC_N.t100 1.1255
R13172 VDAC_N.n1459 VDAC_N.t1635 1.1255
R13173 VDAC_N.n1460 VDAC_N.t1061 1.1255
R13174 VDAC_N.n1461 VDAC_N.t1525 1.1255
R13175 VDAC_N.n1462 VDAC_N.t1983 1.1255
R13176 VDAC_N.n1463 VDAC_N.t1176 1.1255
R13177 VDAC_N.n1464 VDAC_N.t897 1.1255
R13178 VDAC_N.n1465 VDAC_N.t116 1.1255
R13179 VDAC_N.n1466 VDAC_N.t346 1.1255
R13180 VDAC_N.n1467 VDAC_N.t2123 1.1255
R13181 VDAC_N.n1468 VDAC_N.t558 1.1255
R13182 VDAC_N.n1469 VDAC_N.t2009 1.1255
R13183 VDAC_N.n1470 VDAC_N.t656 1.1255
R13184 VDAC_N.n1471 VDAC_N.t918 1.1255
R13185 VDAC_N.n1472 VDAC_N.t1668 1.1255
R13186 VDAC_N.n1473 VDAC_N.t1350 1.1255
R13187 VDAC_N.n1474 VDAC_N.t595 1.1255
R13188 VDAC_N.n1475 VDAC_N.t1146 1.1255
R13189 VDAC_N.n1476 VDAC_N.t2078 1.1255
R13190 VDAC_N.n1477 VDAC_N.t1384 1.1255
R13191 VDAC_N.n1478 VDAC_N.t1858 1.1255
R13192 VDAC_N.n1479 VDAC_N.t1411 1.1255
R13193 VDAC_N.n1480 VDAC_N.t1602 1.1255
R13194 VDAC_N.n1481 VDAC_N.t367 1.1255
R13195 VDAC_N.n1482 VDAC_N.t1847 1.1255
R13196 VDAC_N.n1483 VDAC_N.t1165 1.1255
R13197 VDAC_N.n1484 VDAC_N.t1629 1.1255
R13198 VDAC_N.n1485 VDAC_N.t2134 1.1255
R13199 VDAC_N.n1486 VDAC_N.t1519 1.1255
R13200 VDAC_N.n1487 VDAC_N.t1003 1.1255
R13201 VDAC_N.n1488 VDAC_N.t1415 1.1255
R13202 VDAC_N.n1489 VDAC_N.t1877 1.1255
R13203 VDAC_N.n1490 VDAC_N.t708 1.1255
R13204 VDAC_N.n1491 VDAC_N.t1763 1.1255
R13205 VDAC_N.n1492 VDAC_N.t300 1.1255
R13206 VDAC_N.n1493 VDAC_N.t2120 1.1255
R13207 VDAC_N.n1494 VDAC_N.t2005 1.1255
R13208 VDAC_N.n1495 VDAC_N.t872 1.1255
R13209 VDAC_N.n1496 VDAC_N.t1901 1.1255
R13210 VDAC_N.n1497 VDAC_N.t1636 1.1255
R13211 VDAC_N.n1498 VDAC_N.t1586 1.1255
R13212 VDAC_N.n1499 VDAC_N.t1484 1.1255
R13213 VDAC_N.n1500 VDAC_N.t306 1.1255
R13214 VDAC_N.n1501 VDAC_N.t593 1.1255
R13215 VDAC_N.n1502 VDAC_N.t928 1.1255
R13216 VDAC_N.n94 VDAC_N.t713 1.1255
R13217 VDAC_N.n1503 VDAC_N.t710 1.1255
R13218 VDAC_N.n1504 VDAC_N.t1283 1.1255
R13219 VDAC_N.n1505 VDAC_N.t314 1.1255
R13220 VDAC_N.n1506 VDAC_N.t1066 1.1255
R13221 VDAC_N.n1507 VDAC_N.t1531 1.1255
R13222 VDAC_N.n1508 VDAC_N.t1894 1.1255
R13223 VDAC_N.n1509 VDAC_N.t1421 1.1255
R13224 VDAC_N.n1510 VDAC_N.t1885 1.1255
R13225 VDAC_N.n1511 VDAC_N.t189 1.1255
R13226 VDAC_N.n1512 VDAC_N.t1773 1.1255
R13227 VDAC_N.n1513 VDAC_N.t1091 1.1255
R13228 VDAC_N.n1514 VDAC_N.t1667 1.1255
R13229 VDAC_N.n1515 VDAC_N.t2127 1.1255
R13230 VDAC_N.n1516 VDAC_N.t1422 1.1255
R13231 VDAC_N.n1517 VDAC_N.t1195 1.1255
R13232 VDAC_N.n1518 VDAC_N.t245 1.1255
R13233 VDAC_N.n1519 VDAC_N.t23 1.1255
R13234 VDAC_N.n1520 VDAC_N.t1549 1.1255
R13235 VDAC_N.n1521 VDAC_N.t1073 1.1255
R13236 VDAC_N.n1522 VDAC_N.t1443 1.1255
R13237 VDAC_N.n1523 VDAC_N.t965 1.1255
R13238 VDAC_N.n1524 VDAC_N.t1339 1.1255
R13239 VDAC_N.n1525 VDAC_N.t1795 1.1255
R13240 VDAC_N.n1526 VDAC_N.t396 1.1255
R13241 VDAC_N.n1527 VDAC_N.t1579 1.1255
R13242 VDAC_N.n1528 VDAC_N.t1074 1.1255
R13243 VDAC_N.n1529 VDAC_N.t1832 1.1255
R13244 VDAC_N.n1530 VDAC_N.t503 1.1255
R13245 VDAC_N.n1531 VDAC_N.t1376 1.1255
R13246 VDAC_N.n1532 VDAC_N.t1825 1.1255
R13247 VDAC_N.n1533 VDAC_N.t972 1.1255
R13248 VDAC_N.n1534 VDAC_N.t1410 1.1255
R13249 VDAC_N.n1535 VDAC_N.t476 1.1255
R13250 VDAC_N.n1536 VDAC_N.t504 1.1255
R13251 VDAC_N.n1537 VDAC_N.t502 1.1255
R13252 VDAC_N.n1538 VDAC_N.t392 1.1255
R13253 VDAC_N.n1539 VDAC_N.t54 1.1255
R13254 VDAC_N.n1540 VDAC_N.t1220 1.1255
R13255 VDAC_N.n1541 VDAC_N.t118 1.1255
R13256 VDAC_N.n1542 VDAC_N.t623 1.1255
R13257 VDAC_N.n1543 VDAC_N.t618 1.1255
R13258 VDAC_N.n1544 VDAC_N.t1189 1.1255
R13259 VDAC_N.n1545 VDAC_N.t435 1.1255
R13260 VDAC_N.n1546 VDAC_N.t266 1.1255
R13261 VDAC_N.n1547 VDAC_N.t1439 1.1255
R13262 VDAC_N.n1548 VDAC_N.t1999 1.1255
R13263 VDAC_N.n1549 VDAC_N.t191 1.1255
R13264 VDAC_N.n1550 VDAC_N.t909 1.1255
R13265 VDAC_N.n1551 VDAC_N.t1223 1.1255
R13266 VDAC_N.n1552 VDAC_N.t443 1.1255
R13267 VDAC_N.n1553 VDAC_N.t970 1.1255
R13268 VDAC_N.n1554 VDAC_N.t1573 1.1255
R13269 VDAC_N.n1555 VDAC_N.t2037 1.1255
R13270 VDAC_N.n1556 VDAC_N.t688 1.1255
R13271 VDAC_N.n1557 VDAC_N.t35 1.1255
R13272 VDAC_N.n1558 VDAC_N.t932 1.1255
R13273 VDAC_N.n1559 VDAC_N.t869 1.1255
R13274 VDAC_N.n1560 VDAC_N.t12 1.1255
R13275 VDAC_N.n1561 VDAC_N.t606 1.1255
R13276 VDAC_N.n1562 VDAC_N.t2063 1.1255
R13277 VDAC_N.n1563 VDAC_N.t208 1.1255
R13278 VDAC_N.n1564 VDAC_N.t1910 1.1255
R13279 VDAC_N.n1565 VDAC_N.t1060 1.1255
R13280 VDAC_N.n93 VDAC_N.t712 1.1255
R13281 VDAC_N.n1566 VDAC_N.t1831 1.1255
R13282 VDAC_N.n1567 VDAC_N.t964 1.1255
R13283 VDAC_N.n1568 VDAC_N.t875 1.1255
R13284 VDAC_N.n1569 VDAC_N.t540 1.1255
R13285 VDAC_N.n1570 VDAC_N.t992 1.1255
R13286 VDAC_N.n1571 VDAC_N.t2075 1.1255
R13287 VDAC_N.n1572 VDAC_N.t768 1.1255
R13288 VDAC_N.n1573 VDAC_N.t1706 1.1255
R13289 VDAC_N.n1574 VDAC_N.t1088 1.1255
R13290 VDAC_N.n1575 VDAC_N.t754 1.1255
R13291 VDAC_N.n1576 VDAC_N.t1724 1.1255
R13292 VDAC_N.n1577 VDAC_N.t1262 1.1255
R13293 VDAC_N.n1578 VDAC_N.t1109 1.1255
R13294 VDAC_N.n1579 VDAC_N.t385 1.1255
R13295 VDAC_N.n1580 VDAC_N.t1915 1.1255
R13296 VDAC_N.n1581 VDAC_N.t1312 1.1255
R13297 VDAC_N.n1582 VDAC_N.t473 1.1255
R13298 VDAC_N.n1583 VDAC_N.t236 1.1255
R13299 VDAC_N.n1584 VDAC_N.t698 1.1255
R13300 VDAC_N.n1585 VDAC_N.t1948 1.1255
R13301 VDAC_N.n1586 VDAC_N.t1880 1.1255
R13302 VDAC_N.n1587 VDAC_N.t281 1.1255
R13303 VDAC_N.n1588 VDAC_N.t728 1.1255
R13304 VDAC_N.n1589 VDAC_N.t1658 1.1255
R13305 VDAC_N.n1590 VDAC_N.t1068 1.1255
R13306 VDAC_N.n1591 VDAC_N.t1430 1.1255
R13307 VDAC_N.n1592 VDAC_N.t321 1.1255
R13308 VDAC_N.n1593 VDAC_N.t2000 1.1255
R13309 VDAC_N.n1594 VDAC_N.t61 1.1255
R13310 VDAC_N.n1595 VDAC_N.t408 1.1255
R13311 VDAC_N.n1596 VDAC_N.t1722 1.1255
R13312 VDAC_N.n1597 VDAC_N.t383 1.1255
R13313 VDAC_N.n1598 VDAC_N.t1502 1.1255
R13314 VDAC_N.n1599 VDAC_N.t1229 1.1255
R13315 VDAC_N.n1600 VDAC_N.t1697 1.1255
R13316 VDAC_N.n1601 VDAC_N.t1117 1.1255
R13317 VDAC_N.n1602 VDAC_N.t1583 1.1255
R13318 VDAC_N.n1603 VDAC_N.t902 1.1255
R13319 VDAC_N.n1604 VDAC_N.t1471 1.1255
R13320 VDAC_N.n1605 VDAC_N.t1931 1.1255
R13321 VDAC_N.n1606 VDAC_N.t1347 1.1255
R13322 VDAC_N.n1607 VDAC_N.t967 1.1255
R13323 VDAC_N.n1608 VDAC_N.t1700 1.1255
R13324 VDAC_N.n1609 VDAC_N.t237 1.1255
R13325 VDAC_N.n1610 VDAC_N.t1372 1.1255
R13326 VDAC_N.n1611 VDAC_N.t590 1.1255
R13327 VDAC_N.n1612 VDAC_N.t1037 1.1255
R13328 VDAC_N.n1613 VDAC_N.t200 1.1255
R13329 VDAC_N.n1614 VDAC_N.t1935 1.1255
R13330 VDAC_N.n1615 VDAC_N.t1924 1.1255
R13331 VDAC_N.n1616 VDAC_N.t722 1.1255
R13332 VDAC_N.n1617 VDAC_N.t524 1.1255
R13333 VDAC_N.n1618 VDAC_N.t622 1.1255
R13334 VDAC_N.n1619 VDAC_N.t19 1.1255
R13335 VDAC_N.n1620 VDAC_N.t1528 1.1255
R13336 VDAC_N.n1621 VDAC_N.t1942 1.1255
R13337 VDAC_N.n1622 VDAC_N.t1104 1.1255
R13338 VDAC_N.n1623 VDAC_N.t1490 1.1255
R13339 VDAC_N.n1624 VDAC_N.t1337 1.1255
R13340 VDAC_N.n1625 VDAC_N.t650 1.1255
R13341 VDAC_N.n1626 VDAC_N.t299 1.1255
R13342 VDAC_N.n1627 VDAC_N.t41 1.1255
R13343 VDAC_N.n1628 VDAC_N.t1014 1.1255
R13344 VDAC_N.n92 VDAC_N.t1733 1.1255
R13345 VDAC_N.n1629 VDAC_N.t1054 1.1255
R13346 VDAC_N.n1630 VDAC_N.t427 1.1255
R13347 VDAC_N.n1631 VDAC_N.t486 1.1255
R13348 VDAC_N.n1632 VDAC_N.t201 1.1255
R13349 VDAC_N.n1633 VDAC_N.t1873 1.1255
R13350 VDAC_N.n1634 VDAC_N.t665 1.1255
R13351 VDAC_N.n1635 VDAC_N.t1759 1.1255
R13352 VDAC_N.n1636 VDAC_N.t60 1.1255
R13353 VDAC_N.n1637 VDAC_N.t1657 1.1255
R13354 VDAC_N.n1638 VDAC_N.t2113 1.1255
R13355 VDAC_N.n1639 VDAC_N.t381 1.1255
R13356 VDAC_N.n1640 VDAC_N.t521 1.1255
R13357 VDAC_N.n1641 VDAC_N.t1256 1.1255
R13358 VDAC_N.n1642 VDAC_N.t1263 1.1255
R13359 VDAC_N.n1643 VDAC_N.t1725 1.1255
R13360 VDAC_N.n1644 VDAC_N.t2028 1.1255
R13361 VDAC_N.n1645 VDAC_N.t1617 1.1255
R13362 VDAC_N.n1646 VDAC_N.t1053 1.1255
R13363 VDAC_N.n1647 VDAC_N.t1000 1.1255
R13364 VDAC_N.n1648 VDAC_N.t1965 1.1255
R13365 VDAC_N.n1649 VDAC_N.t568 1.1255
R13366 VDAC_N.n1650 VDAC_N.t947 1.1255
R13367 VDAC_N.n1651 VDAC_N.t68 1.1255
R13368 VDAC_N.n1652 VDAC_N.t1274 1.1255
R13369 VDAC_N.n1653 VDAC_N.t1067 1.1255
R13370 VDAC_N.n1654 VDAC_N.t1056 1.1255
R13371 VDAC_N.n1655 VDAC_N.t2002 1.1255
R13372 VDAC_N.n1656 VDAC_N.t632 1.1255
R13373 VDAC_N.n1657 VDAC_N.t898 1.1255
R13374 VDAC_N.n1658 VDAC_N.t1540 1.1255
R13375 VDAC_N.n1659 VDAC_N.t678 1.1255
R13376 VDAC_N.n1660 VDAC_N.t1255 1.1255
R13377 VDAC_N.n1661 VDAC_N.t1118 1.1255
R13378 VDAC_N.n1662 VDAC_N.t1038 1.1255
R13379 VDAC_N.n1663 VDAC_N.t1499 1.1255
R13380 VDAC_N.n1664 VDAC_N.t478 1.1255
R13381 VDAC_N.n1665 VDAC_N.t199 1.1255
R13382 VDAC_N.n1666 VDAC_N.t1386 1.1255
R13383 VDAC_N.n1667 VDAC_N.t655 1.1255
R13384 VDAC_N.n1668 VDAC_N.t243 1.1255
R13385 VDAC_N.n1669 VDAC_N.t309 1.1255
R13386 VDAC_N.n1670 VDAC_N.t873 1.1255
R13387 VDAC_N.n1671 VDAC_N.t1884 1.1255
R13388 VDAC_N.n1672 VDAC_N.t1505 1.1255
R13389 VDAC_N.n1673 VDAC_N.t1957 1.1255
R13390 VDAC_N.n1674 VDAC_N.t120 1.1255
R13391 VDAC_N.n1675 VDAC_N.t1859 1.1255
R13392 VDAC_N.n1676 VDAC_N.t644 1.1255
R13393 VDAC_N.n1677 VDAC_N.t1753 1.1255
R13394 VDAC_N.n1678 VDAC_N.t828 1.1255
R13395 VDAC_N.n1679 VDAC_N.t2064 1.1255
R13396 VDAC_N.n1680 VDAC_N.t2099 1.1255
R13397 VDAC_N.n1681 VDAC_N.t1656 1.1255
R13398 VDAC_N.n1682 VDAC_N.t890 1.1255
R13399 VDAC_N.n1683 VDAC_N.t1492 1.1255
R13400 VDAC_N.n1684 VDAC_N.t218 1.1255
R13401 VDAC_N.n1685 VDAC_N.t1260 1.1255
R13402 VDAC_N.n1686 VDAC_N.t298 1.1255
R13403 VDAC_N.n1687 VDAC_N.t1139 1.1255
R13404 VDAC_N.n1688 VDAC_N.t896 1.1255
R13405 VDAC_N.n1689 VDAC_N.t42 1.1255
R13406 VDAC_N.n1690 VDAC_N.t761 1.1255
R13407 VDAC_N.n1691 VDAC_N.t226 1.1255
R13408 VDAC_N.n91 VDAC_N.t1394 1.1255
R13409 VDAC_N.n1692 VDAC_N.t20 1.1255
R13410 VDAC_N.n1693 VDAC_N.t602 1.1255
R13411 VDAC_N.n1694 VDAC_N.t2059 1.1255
R13412 VDAC_N.n1695 VDAC_N.t1456 1.1255
R13413 VDAC_N.n1696 VDAC_N.t1678 1.1255
R13414 VDAC_N.n1697 VDAC_N.t1044 1.1255
R13415 VDAC_N.n1698 VDAC_N.t738 1.1255
R13416 VDAC_N.n1699 VDAC_N.t1211 1.1255
R13417 VDAC_N.n1700 VDAC_N.t330 1.1255
R13418 VDAC_N.n1701 VDAC_N.t561 1.1255
R13419 VDAC_N.n1702 VDAC_N.t224 1.1255
R13420 VDAC_N.n1703 VDAC_N.t1958 1.1255
R13421 VDAC_N.n1704 VDAC_N.t741 1.1255
R13422 VDAC_N.n1705 VDAC_N.t1981 1.1255
R13423 VDAC_N.n1706 VDAC_N.t312 1.1255
R13424 VDAC_N.n1707 VDAC_N.t882 1.1255
R13425 VDAC_N.n1708 VDAC_N.t724 1.1255
R13426 VDAC_N.n1709 VDAC_N.t1294 1.1255
R13427 VDAC_N.n1710 VDAC_N.t179 1.1255
R13428 VDAC_N.n1711 VDAC_N.t94 1.1255
R13429 VDAC_N.n1712 VDAC_N.t526 1.1255
R13430 VDAC_N.n1713 VDAC_N.t240 1.1255
R13431 VDAC_N.n1714 VDAC_N.t1802 1.1255
R13432 VDAC_N.n1715 VDAC_N.t197 1.1255
R13433 VDAC_N.n1716 VDAC_N.t358 1.1255
R13434 VDAC_N.n1717 VDAC_N.t647 1.1255
R13435 VDAC_N.n1718 VDAC_N.t1729 1.1255
R13436 VDAC_N.n1719 VDAC_N.t2074 1.1255
R13437 VDAC_N.n1720 VDAC_N.t1621 1.1255
R13438 VDAC_N.n1721 VDAC_N.t942 1.1255
R13439 VDAC_N.n1722 VDAC_N.t719 1.1255
R13440 VDAC_N.n1723 VDAC_N.t999 1.1255
R13441 VDAC_N.n1724 VDAC_N.t1299 1.1255
R13442 VDAC_N.n1725 VDAC_N.t893 1.1255
R13443 VDAC_N.n1726 VDAC_N.t1916 1.1255
R13444 VDAC_N.n1727 VDAC_N.t1655 1.1255
R13445 VDAC_N.n1728 VDAC_N.t2109 1.1255
R13446 VDAC_N.n1729 VDAC_N.t731 1.1255
R13447 VDAC_N.n1730 VDAC_N.t1013 1.1255
R13448 VDAC_N.n1731 VDAC_N.t104 1.1255
R13449 VDAC_N.n1732 VDAC_N.t1875 1.1255
R13450 VDAC_N.n1733 VDAC_N.t1128 1.1255
R13451 VDAC_N.n1734 VDAC_N.t1510 1.1255
R13452 VDAC_N.n1735 VDAC_N.t556 1.1255
R13453 VDAC_N.n1736 VDAC_N.t2112 1.1255
R13454 VDAC_N.n1737 VDAC_N.t1121 1.1255
R13455 VDAC_N.n1738 VDAC_N.t1704 1.1255
R13456 VDAC_N.n1739 VDAC_N.t1790 1.1255
R13457 VDAC_N.n1740 VDAC_N.t336 1.1255
R13458 VDAC_N.n1741 VDAC_N.t222 1.1255
R13459 VDAC_N.n1742 VDAC_N.t1261 1.1255
R13460 VDAC_N.n1743 VDAC_N.t1338 1.1255
R13461 VDAC_N.n1744 VDAC_N.t169 1.1255
R13462 VDAC_N.n1745 VDAC_N.t821 1.1255
R13463 VDAC_N.n1746 VDAC_N.t938 1.1255
R13464 VDAC_N.n1747 VDAC_N.t769 1.1255
R13465 VDAC_N.n1748 VDAC_N.t830 1.1255
R13466 VDAC_N.n1749 VDAC_N.t661 1.1255
R13467 VDAC_N.n1750 VDAC_N.t1863 1.1255
R13468 VDAC_N.n1751 VDAC_N.t1183 1.1255
R13469 VDAC_N.n1752 VDAC_N.t1651 1.1255
R13470 VDAC_N.n1753 VDAC_N.t444 1.1255
R13471 VDAC_N.n1754 VDAC_N.t217 1.1255
R13472 VDAC_N.n90 VDAC_N.t1049 1.1255
R13473 VDAC_N.n1755 VDAC_N.t1399 1.1255
R13474 VDAC_N.n1756 VDAC_N.t991 1.1255
R13475 VDAC_N.n1757 VDAC_N.t657 1.1255
R13476 VDAC_N.n1758 VDAC_N.t889 1.1255
R13477 VDAC_N.n1759 VDAC_N.t764 1.1255
R13478 VDAC_N.n1760 VDAC_N.t1645 1.1255
R13479 VDAC_N.n1761 VDAC_N.t2097 1.1255
R13480 VDAC_N.n1762 VDAC_N.t1640 1.1255
R13481 VDAC_N.n1763 VDAC_N.t1009 1.1255
R13482 VDAC_N.n1764 VDAC_N.t1200 1.1255
R13483 VDAC_N.n1765 VDAC_N.t1777 1.1255
R13484 VDAC_N.n1766 VDAC_N.t740 1.1255
R13485 VDAC_N.n1767 VDAC_N.t670 1.1255
R13486 VDAC_N.n1768 VDAC_N.t1793 1.1255
R13487 VDAC_N.n1769 VDAC_N.t748 1.1255
R13488 VDAC_N.n1770 VDAC_N.t110 1.1255
R13489 VDAC_N.n1771 VDAC_N.t2114 1.1255
R13490 VDAC_N.n1772 VDAC_N.t1824 1.1255
R13491 VDAC_N.n1773 VDAC_N.t2062 1.1255
R13492 VDAC_N.n1774 VDAC_N.t696 1.1255
R13493 VDAC_N.n1775 VDAC_N.t1634 1.1255
R13494 VDAC_N.n1776 VDAC_N.t1860 1.1255
R13495 VDAC_N.n1777 VDAC_N.t1406 1.1255
R13496 VDAC_N.n1778 VDAC_N.t317 1.1255
R13497 VDAC_N.n1779 VDAC_N.t976 1.1255
R13498 VDAC_N.n1780 VDAC_N.t11 1.1255
R13499 VDAC_N.n1781 VDAC_N.t1541 1.1255
R13500 VDAC_N.n1782 VDAC_N.t858 1.1255
R13501 VDAC_N.n1783 VDAC_N.t1431 1.1255
R13502 VDAC_N.n1784 VDAC_N.t1462 1.1255
R13503 VDAC_N.n1785 VDAC_N.t325 1.1255
R13504 VDAC_N.n1786 VDAC_N.t467 1.1255
R13505 VDAC_N.n1787 VDAC_N.t1101 1.1255
R13506 VDAC_N.n1788 VDAC_N.t1567 1.1255
R13507 VDAC_N.n1789 VDAC_N.t2027 1.1255
R13508 VDAC_N.n1790 VDAC_N.t207 1.1255
R13509 VDAC_N.n1791 VDAC_N.t1919 1.1255
R13510 VDAC_N.n1792 VDAC_N.t1241 1.1255
R13511 VDAC_N.n1793 VDAC_N.t1813 1.1255
R13512 VDAC_N.n1794 VDAC_N.t460 1.1255
R13513 VDAC_N.n1795 VDAC_N.t235 1.1255
R13514 VDAC_N.n1796 VDAC_N.t1356 1.1255
R13515 VDAC_N.n1797 VDAC_N.t1126 1.1255
R13516 VDAC_N.n1798 VDAC_N.t529 1.1255
R13517 VDAC_N.n1799 VDAC_N.t1344 1.1255
R13518 VDAC_N.n1800 VDAC_N.t254 1.1255
R13519 VDAC_N.n1801 VDAC_N.t1812 1.1255
R13520 VDAC_N.n1802 VDAC_N.t370 1.1255
R13521 VDAC_N.n1803 VDAC_N.t1804 1.1255
R13522 VDAC_N.n1804 VDAC_N.t46 1.1255
R13523 VDAC_N.n1805 VDAC_N.t8 1.1255
R13524 VDAC_N.n1806 VDAC_N.t496 1.1255
R13525 VDAC_N.n1807 VDAC_N.t966 1.1255
R13526 VDAC_N.n1808 VDAC_N.t377 1.1255
R13527 VDAC_N.n1809 VDAC_N.t206 1.1255
R13528 VDAC_N.n1810 VDAC_N.t675 1.1255
R13529 VDAC_N.n1811 VDAC_N.t634 1.1255
R13530 VDAC_N.n1812 VDAC_N.t1095 1.1255
R13531 VDAC_N.n1813 VDAC_N.t1673 1.1255
R13532 VDAC_N.n1814 VDAC_N.t1962 1.1255
R13533 VDAC_N.n1815 VDAC_N.t1455 1.1255
R13534 VDAC_N.n1816 VDAC_N.t277 1.1255
R13535 VDAC_N.n1817 VDAC_N.t1353 1.1255
R13536 VDAC_N.n89 VDAC_N.t187 1.1255
R13537 VDAC_N.n1818 VDAC_N.t1202 1.1255
R13538 VDAC_N.n1819 VDAC_N.t607 1.1255
R13539 VDAC_N.n1820 VDAC_N.t1936 1.1255
R13540 VDAC_N.n1821 VDAC_N.t978 1.1255
R13541 VDAC_N.n1822 VDAC_N.t1437 1.1255
R13542 VDAC_N.n1823 VDAC_N.t862 1.1255
R13543 VDAC_N.n1824 VDAC_N.t679 1.1255
R13544 VDAC_N.n1825 VDAC_N.t83 1.1255
R13545 VDAC_N.n1826 VDAC_N.t1219 1.1255
R13546 VDAC_N.n1827 VDAC_N.t1683 1.1255
R13547 VDAC_N.n1828 VDAC_N.t1982 1.1255
R13548 VDAC_N.n1829 VDAC_N.t413 1.1255
R13549 VDAC_N.n1830 VDAC_N.t2031 1.1255
R13550 VDAC_N.n1831 VDAC_N.t1603 1.1255
R13551 VDAC_N.n1832 VDAC_N.t155 1.1255
R13552 VDAC_N.n1833 VDAC_N.t1904 1.1255
R13553 VDAC_N.n1834 VDAC_N.t1945 1.1255
R13554 VDAC_N.n1835 VDAC_N.t2068 1.1255
R13555 VDAC_N.n1836 VDAC_N.t1674 1.1255
R13556 VDAC_N.n1837 VDAC_N.t1156 1.1255
R13557 VDAC_N.n1838 VDAC_N.t1242 1.1255
R13558 VDAC_N.n1839 VDAC_N.t316 1.1255
R13559 VDAC_N.n1840 VDAC_N.t2032 1.1255
R13560 VDAC_N.n1841 VDAC_N.t270 1.1255
R13561 VDAC_N.n1842 VDAC_N.t1168 1.1255
R13562 VDAC_N.n1843 VDAC_N.t242 1.1255
R13563 VDAC_N.n1844 VDAC_N.t691 1.1255
R13564 VDAC_N.n1845 VDAC_N.t662 1.1255
R13565 VDAC_N.n1846 VDAC_N.t1237 1.1255
R13566 VDAC_N.n1847 VDAC_N.t1086 1.1255
R13567 VDAC_N.n1848 VDAC_N.t2022 1.1255
R13568 VDAC_N.n1849 VDAC_N.t811 1.1255
R13569 VDAC_N.n1850 VDAC_N.t250 1.1255
R13570 VDAC_N.n1851 VDAC_N.t1381 1.1255
R13571 VDAC_N.n1852 VDAC_N.t1839 1.1255
R13572 VDAC_N.n1853 VDAC_N.t1267 1.1255
R13573 VDAC_N.n1854 VDAC_N.t879 1.1255
R13574 VDAC_N.n1855 VDAC_N.t30 1.1255
R13575 VDAC_N.n1856 VDAC_N.t1623 1.1255
R13576 VDAC_N.n1857 VDAC_N.t2083 1.1255
R13577 VDAC_N.n1858 VDAC_N.t393 1.1255
R13578 VDAC_N.n1859 VDAC_N.t2055 1.1255
R13579 VDAC_N.n1860 VDAC_N.t1448 1.1255
R13580 VDAC_N.n1861 VDAC_N.t1845 1.1255
R13581 VDAC_N.n1862 VDAC_N.t1108 1.1255
R13582 VDAC_N.n1863 VDAC_N.t734 1.1255
R13583 VDAC_N.n1864 VDAC_N.t554 1.1255
R13584 VDAC_N.n1865 VDAC_N.t152 1.1255
R13585 VDAC_N.n1866 VDAC_N.t2087 1.1255
R13586 VDAC_N.n1867 VDAC_N.t1568 1.1255
R13587 VDAC_N.n1868 VDAC_N.t1730 1.1255
R13588 VDAC_N.n1869 VDAC_N.t304 1.1255
R13589 VDAC_N.n1870 VDAC_N.t1514 1.1255
R13590 VDAC_N.n1871 VDAC_N.t1231 1.1255
R13591 VDAC_N.n1872 VDAC_N.t1072 1.1255
R13592 VDAC_N.n1873 VDAC_N.t1123 1.1255
R13593 VDAC_N.n1874 VDAC_N.t448 1.1255
R13594 VDAC_N.n1875 VDAC_N.t1794 1.1255
R13595 VDAC_N.n1876 VDAC_N.t1475 1.1255
R13596 VDAC_N.n1877 VDAC_N.t1582 1.1255
R13597 VDAC_N.n1878 VDAC_N.t645 1.1255
R13598 VDAC_N.n1879 VDAC_N.t479 1.1255
R13599 VDAC_N.n1880 VDAC_N.t1157 1.1255
R13600 VDAC_N.n88 VDAC_N.t1028 1.1255
R13601 VDAC_N.n1881 VDAC_N.t455 1.1255
R13602 VDAC_N.n1882 VDAC_N.t564 1.1255
R13603 VDAC_N.n1883 VDAC_N.t53 1.1255
R13604 VDAC_N.n1884 VDAC_N.t2089 1.1255
R13605 VDAC_N.n1885 VDAC_N.t1576 1.1255
R13606 VDAC_N.n1886 VDAC_N.t1977 1.1255
R13607 VDAC_N.n1887 VDAC_N.t1144 1.1255
R13608 VDAC_N.n1888 VDAC_N.t1518 1.1255
R13609 VDAC_N.n1889 VDAC_N.t196 1.1255
R13610 VDAC_N.n1890 VDAC_N.t658 1.1255
R13611 VDAC_N.n1891 VDAC_N.t2119 1.1255
R13612 VDAC_N.n1892 VDAC_N.t288 1.1255
R13613 VDAC_N.n1893 VDAC_N.t90 1.1255
R13614 VDAC_N.n1894 VDAC_N.t1284 1.1255
R13615 VDAC_N.n1895 VDAC_N.t338 1.1255
R13616 VDAC_N.n1896 VDAC_N.t1225 1.1255
R13617 VDAC_N.n1897 VDAC_N.t32 1.1255
R13618 VDAC_N.n1898 VDAC_N.t274 1.1255
R13619 VDAC_N.n1899 VDAC_N.t415 1.1255
R13620 VDAC_N.n1900 VDAC_N.t1762 1.1255
R13621 VDAC_N.n1901 VDAC_N.t697 1.1255
R13622 VDAC_N.n1902 VDAC_N.t1554 1.1255
R13623 VDAC_N.n1903 VDAC_N.t181 1.1255
R13624 VDAC_N.n1904 VDAC_N.t1713 1.1255
R13625 VDAC_N.n1905 VDAC_N.t2046 1.1255
R13626 VDAC_N.n1906 VDAC_N.t1607 1.1255
R13627 VDAC_N.n1907 VDAC_N.t2067 1.1255
R13628 VDAC_N.n1908 VDAC_N.t1395 1.1255
R13629 VDAC_N.n1909 VDAC_N.t989 1.1255
R13630 VDAC_N.n1910 VDAC_N.t341 1.1255
R13631 VDAC_N.n1911 VDAC_N.t1745 1.1255
R13632 VDAC_N.n1912 VDAC_N.t612 1.1255
R13633 VDAC_N.n1913 VDAC_N.t833 1.1255
R13634 VDAC_N.n1914 VDAC_N.t2095 1.1255
R13635 VDAC_N.n1915 VDAC_N.t424 1.1255
R13636 VDAC_N.n1916 VDAC_N.t1985 1.1255
R13637 VDAC_N.n1917 VDAC_N.t64 1.1255
R13638 VDAC_N.n1918 VDAC_N.t1769 1.1255
R13639 VDAC_N.n1919 VDAC_N.t1444 1.1255
R13640 VDAC_N.n1920 VDAC_N.t1302 1.1255
R13641 VDAC_N.n1921 VDAC_N.t380 1.1255
R13642 VDAC_N.n1922 VDAC_N.t1254 1.1255
R13643 VDAC_N.n1923 VDAC_N.t1105 1.1255
R13644 VDAC_N.n1924 VDAC_N.t832 1.1255
R13645 VDAC_N.n1925 VDAC_N.t458 1.1255
R13646 VDAC_N.n1926 VDAC_N.t1463 1.1255
R13647 VDAC_N.n1927 VDAC_N.t786 1.1255
R13648 VDAC_N.n1928 VDAC_N.t1247 1.1255
R13649 VDAC_N.n1929 VDAC_N.t38 1.1255
R13650 VDAC_N.n1930 VDAC_N.t305 1.1255
R13651 VDAC_N.n1931 VDAC_N.t815 1.1255
R13652 VDAC_N.n1932 VDAC_N.t1030 1.1255
R13653 VDAC_N.n1933 VDAC_N.t1493 1.1255
R13654 VDAC_N.n1934 VDAC_N.t507 1.1255
R13655 VDAC_N.n1935 VDAC_N.t651 1.1255
R13656 VDAC_N.n1936 VDAC_N.t1851 1.1255
R13657 VDAC_N.n1937 VDAC_N.t313 1.1255
R13658 VDAC_N.n1938 VDAC_N.t1633 1.1255
R13659 VDAC_N.n1939 VDAC_N.t572 1.1255
R13660 VDAC_N.n1940 VDAC_N.t775 1.1255
R13661 VDAC_N.n1941 VDAC_N.t89 1.1255
R13662 VDAC_N.n1942 VDAC_N.t1584 1.1255
R13663 VDAC_N.n1943 VDAC_N.t491 1.1255
R13664 VDAC_N.n87 VDAC_N.t431 1.1255
R13665 VDAC_N.n86 VDAC_N.t494 1.1255
R13666 VDAC_N.n85 VDAC_N.t403 1.1255
R13667 VDAC_N.n84 VDAC_N.t846 1.1255
R13668 VDAC_N.n83 VDAC_N.t1315 1.1255
R13669 VDAC_N.n82 VDAC_N.t137 1.1255
R13670 VDAC_N.n81 VDAC_N.t175 1.1255
R13671 VDAC_N.n80 VDAC_N.t847 1.1255
R13672 VDAC_N.n79 VDAC_N.t1077 1.1255
R13673 VDAC_N.n78 VDAC_N.t1557 1.1255
R13674 VDAC_N.n77 VDAC_N.t1021 1.1255
R13675 VDAC_N.n76 VDAC_N.t193 1.1255
R13676 VDAC_N.n75 VDAC_N.t1907 1.1255
R13677 VDAC_N.n74 VDAC_N.t868 1.1255
R13678 VDAC_N.n73 VDAC_N.t1079 1.1255
R13679 VDAC_N.n72 VDAC_N.t1752 1.1255
R13680 VDAC_N.n71 VDAC_N.t2034 1.1255
R13681 VDAC_N.n70 VDAC_N.t1304 1.1255
R13682 VDAC_N.n69 VDAC_N.t818 1.1255
R13683 VDAC_N.n68 VDAC_N.t1387 1.1255
R13684 VDAC_N.n67 VDAC_N.t362 1.1255
R13685 VDAC_N.n66 VDAC_N.t1169 1.1255
R13686 VDAC_N.n65 VDAC_N.t1158 1.1255
R13687 VDAC_N.n64 VDAC_N.t1058 1.1255
R13688 VDAC_N.n63 VDAC_N.t1523 1.1255
R13689 VDAC_N.n62 VDAC_N.t842 1.1255
R13690 VDAC_N.n61 VDAC_N.t375 1.1255
R13691 VDAC_N.n60 VDAC_N.t1881 1.1255
R13692 VDAC_N.n59 VDAC_N.t1199 1.1255
R13693 VDAC_N.n58 VDAC_N.t1765 1.1255
R13694 VDAC_N.n57 VDAC_N.t555 1.1255
R13695 VDAC_N.n56 VDAC_N.t1553 1.1255
R13696 VDAC_N.n55 VDAC_N.t551 1.1255
R13697 VDAC_N.n54 VDAC_N.t737 1.1255
R13698 VDAC_N.n53 VDAC_N.t497 1.1255
R13699 VDAC_N.n52 VDAC_N.t836 1.1255
R13700 VDAC_N.n51 VDAC_N.t1797 1.1255
R13701 VDAC_N.n50 VDAC_N.t780 1.1255
R13702 VDAC_N.n49 VDAC_N.t805 1.1255
R13703 VDAC_N.n48 VDAC_N.t2122 1.1255
R13704 VDAC_N.n47 VDAC_N.t1840 1.1255
R13705 VDAC_N.n46 VDAC_N.t59 1.1255
R13706 VDAC_N.n45 VDAC_N.t880 1.1255
R13707 VDAC_N.n44 VDAC_N.t1810 1.1255
R13708 VDAC_N.n43 VDAC_N.t1684 1.1255
R13709 VDAC_N.n42 VDAC_N.t1354 1.1255
R13710 VDAC_N.n41 VDAC_N.t649 1.1255
R13711 VDAC_N.n40 VDAC_N.t98 1.1255
R13712 VDAC_N.n39 VDAC_N.t2082 1.1255
R13713 VDAC_N.n38 VDAC_N.t1848 1.1255
R13714 VDAC_N.n37 VDAC_N.t1862 1.1255
R13715 VDAC_N.n36 VDAC_N.t1413 1.1255
R13716 VDAC_N.n35 VDAC_N.t1642 1.1255
R13717 VDAC_N.n34 VDAC_N.t1303 1.1255
R13718 VDAC_N.n33 VDAC_N.t1761 1.1255
R13719 VDAC_N.n32 VDAC_N.t17 1.1255
R13720 VDAC_N.n31 VDAC_N.t843 1.1255
R13721 VDAC_N.n30 VDAC_N.t1938 1.1255
R13722 VDAC_N.n29 VDAC_N.t1441 1.1255
R13723 VDAC_N.n28 VDAC_N.t2001 1.1255
R13724 VDAC_N.n27 VDAC_N.t1335 1.1255
R13725 VDAC_N.n26 VDAC_N.t469 1.1255
R13726 VDAC_N.n25 VDAC_N.t1588 1.1255
R13727 VDAC_N.n24 VDAC_N.t1691 1.1255
R13728 VDAC_N.n23 VDAC_N.t1380 1.1255
R13729 VDAC_N.n1944 VDAC_N.t372 1.1255
R13730 VDAC_N.n1945 VDAC_N.t1615 1.1255
R13731 VDAC_N.n1946 VDAC_N.t917 1.1255
R13732 VDAC_N.n1947 VDAC_N.t1993 1.1255
R13733 VDAC_N.n1948 VDAC_N.t67 1.1255
R13734 VDAC_N.n1949 VDAC_N.t1467 1.1255
R13735 VDAC_N.n1950 VDAC_N.t742 1.1255
R13736 VDAC_N.n1951 VDAC_N.t1850 1.1255
R13737 VDAC_N.n1952 VDAC_N.t303 1.1255
R13738 VDAC_N.n1953 VDAC_N.t216 1.1255
R13739 VDAC_N.n1954 VDAC_N.t170 1.1255
R13740 VDAC_N.n1955 VDAC_N.t2007 1.1255
R13741 VDAC_N.n1956 VDAC_N.t1276 1.1255
R13742 VDAC_N.n1957 VDAC_N.t1876 1.1255
R13743 VDAC_N.n1958 VDAC_N.t1679 1.1255
R13744 VDAC_N.n1959 VDAC_N.t1869 1.1255
R13745 VDAC_N.n1960 VDAC_N.t587 1.1255
R13746 VDAC_N.n1961 VDAC_N.t1343 1.1255
R13747 VDAC_N.n1962 VDAC_N.t1527 1.1255
R13748 VDAC_N.n1963 VDAC_N.t439 1.1255
R13749 VDAC_N.n1964 VDAC_N.t487 1.1255
R13750 VDAC_N.n1965 VDAC_N.t583 1.1255
R13751 VDAC_N.n1966 VDAC_N.t355 1.1255
R13752 VDAC_N.n1967 VDAC_N.t215 1.1255
R13753 VDAC_N.n1968 VDAC_N.t806 1.1255
R13754 VDAC_N.n1969 VDAC_N.t1966 1.1255
R13755 VDAC_N.n1970 VDAC_N.t148 1.1255
R13756 VDAC_N.n1971 VDAC_N.t1768 1.1255
R13757 VDAC_N.n1972 VDAC_N.t106 1.1255
R13758 VDAC_N.n1973 VDAC_N.t2065 1.1255
R13759 VDAC_N.n1974 VDAC_N.t817 1.1255
R13760 VDAC_N.n1975 VDAC_N.t492 1.1255
R13761 VDAC_N.n1976 VDAC_N.t449 1.1255
R13762 VDAC_N.n1977 VDAC_N.t639 1.1255
R13763 VDAC_N.n1978 VDAC_N.t977 1.1255
R13764 VDAC_N.n1979 VDAC_N.t195 1.1255
R13765 VDAC_N.n1980 VDAC_N.t1758 1.1255
R13766 VDAC_N.n1981 VDAC_N.t1575 1.1255
R13767 VDAC_N.n1982 VDAC_N.t1010 1.1255
R13768 VDAC_N.n1983 VDAC_N.t859 1.1255
R13769 VDAC_N.n1984 VDAC_N.t327 1.1255
R13770 VDAC_N.n1985 VDAC_N.t390 1.1255
R13771 VDAC_N.n1986 VDAC_N.t1333 1.1255
R13772 VDAC_N.n1987 VDAC_N.t866 1.1255
R13773 VDAC_N.n1988 VDAC_N.t1504 1.1255
R13774 VDAC_N.n1989 VDAC_N.t1934 1.1255
R13775 VDAC_N.n1990 VDAC_N.t88 1.1255
R13776 VDAC_N.n1991 VDAC_N.t609 1.1255
R13777 VDAC_N.n1992 VDAC_N.t1210 1.1255
R13778 VDAC_N.n1993 VDAC_N.t1964 1.1255
R13779 VDAC_N.n1994 VDAC_N.t834 1.1255
R13780 VDAC_N.n1995 VDAC_N.t1392 1.1255
R13781 VDAC_N.n1996 VDAC_N.t147 1.1255
R13782 VDAC_N.n1997 VDAC_N.t1488 1.1255
R13783 VDAC_N.n1998 VDAC_N.t2069 1.1255
R13784 VDAC_N.n1999 VDAC_N.t51 1.1255
R13785 VDAC_N.n2000 VDAC_N.t1308 1.1255
R13786 VDAC_N.n2001 VDAC_N.t1715 1.1255
R13787 VDAC_N.n2002 VDAC_N.t1932 1.1255
R13788 VDAC_N.n2003 VDAC_N.t927 1.1255
R13789 VDAC_N.n2004 VDAC_N.t699 1.1255
R13790 VDAC_N.n2005 VDAC_N.t531 1.1255
R13791 VDAC_N.n2006 VDAC_N.t749 1.1255
R13792 VDAC_N.n2007 VDAC_N.t522 1.1255
R13793 VDAC_N.n2008 VDAC_N.t1695 1.1255
R13794 VDAC_N.n2009 VDAC_N.t571 1.1255
R13795 VDAC_N.n2010 VDAC_N.t249 1.1255
R13796 VDAC_N.n2011 VDAC_N.t69 1.1255
R13797 VDAC_N.n2012 VDAC_N.t394 1.1255
R13798 VDAC_N.n2013 VDAC_N.t205 1.1255
R13799 VDAC_N.n2014 VDAC_N.t1946 1.1255
R13800 VDAC_N.n2015 VDAC_N.t272 1.1255
R13801 VDAC_N.n2016 VDAC_N.t29 1.1255
R13802 VDAC_N.n2017 VDAC_N.t326 1.1255
R13803 VDAC_N.n2018 VDAC_N.t1307 1.1255
R13804 VDAC_N.n2019 VDAC_N.t1426 1.1255
R13805 VDAC_N.n2020 VDAC_N.t1972 1.1255
R13806 VDAC_N.n2021 VDAC_N.t1870 1.1255
R13807 VDAC_N.n2022 VDAC_N.t1416 1.1255
R13808 VDAC_N.n2023 VDAC_N.t2051 1.1255
R13809 VDAC_N.n2024 VDAC_N.t279 1.1255
R13810 VDAC_N.n2025 VDAC_N.t221 1.1255
R13811 VDAC_N.n2026 VDAC_N.t1990 1.1255
R13812 VDAC_N.n2027 VDAC_N.t1687 1.1255
R13813 VDAC_N.n2028 VDAC_N.t625 1.1255
R13814 VDAC_N.n2029 VDAC_N.t1789 1.1255
R13815 VDAC_N.n2030 VDAC_N.t1331 1.1255
R13816 VDAC_N.n2031 VDAC_N.t1702 1.1255
R13817 VDAC_N.n2032 VDAC_N.t733 1.1255
R13818 VDAC_N.n2033 VDAC_N.t1930 1.1255
R13819 VDAC_N.n2034 VDAC_N.t1944 1.1255
R13820 VDAC_N.n2035 VDAC_N.t173 1.1255
R13821 VDAC_N.n2036 VDAC_N.t1206 1.1255
R13822 VDAC_N.n2037 VDAC_N.t1301 1.1255
R13823 VDAC_N.n2038 VDAC_N.t1638 1.1255
R13824 VDAC_N.n2039 VDAC_N.t985 1.1255
R13825 VDAC_N.n2040 VDAC_N.t315 1.1255
R13826 VDAC_N.n2041 VDAC_N.t760 1.1255
R13827 VDAC_N.n2042 VDAC_N.t1517 1.1255
R13828 VDAC_N.n2043 VDAC_N.t50 1.1255
R13829 VDAC_N.n2044 VDAC_N.t1857 1.1255
R13830 VDAC_N.n2045 VDAC_N.t15 1.1255
R13831 VDAC_N.n2046 VDAC_N.t1120 1.1255
R13832 VDAC_N.n2047 VDAC_N.t115 1.1255
R13833 VDAC_N.n2048 VDAC_N.t334 1.1255
R13834 VDAC_N.n2049 VDAC_N.t536 1.1255
R13835 VDAC_N.n2050 VDAC_N.t963 1.1255
R13836 VDAC_N.n2051 VDAC_N.t1119 1.1255
R13837 VDAC_N.n2052 VDAC_N.t1196 1.1255
R13838 VDAC_N.n2053 VDAC_N.t745 1.1255
R13839 VDAC_N.n2054 VDAC_N.t1696 1.1255
R13840 VDAC_N.n2055 VDAC_N.t1801 1.1255
R13841 VDAC_N.n2056 VDAC_N.t2026 1.1255
R13842 VDAC_N.n2057 VDAC_N.t1187 1.1255
R13843 VDAC_N.n2058 VDAC_N.t1373 1.1255
R13844 VDAC_N.n2059 VDAC_N.t344 1.1255
R13845 VDAC_N.n2060 VDAC_N.t133 1.1255
R13846 VDAC_N.n2061 VDAC_N.t930 1.1255
R13847 VDAC_N.n2062 VDAC_N.t91 1.1255
R13848 VDAC_N.n2063 VDAC_N.t1269 1.1255
R13849 VDAC_N.n2064 VDAC_N.t916 1.1255
R13850 VDAC_N.n2065 VDAC_N.t1611 1.1255
R13851 VDAC_N.n2066 VDAC_N.t430 1.1255
R13852 VDAC_N.n2067 VDAC_N.t1941 1.1255
R13853 VDAC_N.n2068 VDAC_N.t1173 1.1255
R13854 VDAC_N.n2069 VDAC_N.t268 1.1255
R13855 VDAC_N.n2070 VDAC_N.t322 1.1255
R13856 VDAC_N.n2071 VDAC_N.t1051 1.1255
R13857 VDAC_N.n2072 VDAC_N.t984 1.1255
R13858 VDAC_N.n2073 VDAC_N.t1959 1.1255
R13859 VDAC_N.n2074 VDAC_N.t160 1.1255
R13860 VDAC_N.n2075 VDAC_N.t1478 1.1255
R13861 VDAC_N.n2076 VDAC_N.t340 1.1255
R13862 VDAC_N.n2077 VDAC_N.t182 1.1255
R13863 VDAC_N.n2078 VDAC_N.t163 1.1255
R13864 VDAC_N.n2079 VDAC_N.t1048 1.1255
R13865 VDAC_N.n2080 VDAC_N.t1986 1.1255
R13866 VDAC_N.n2081 VDAC_N.t624 1.1255
R13867 VDAC_N.n2082 VDAC_N.t1754 1.1255
R13868 VDAC_N.n2083 VDAC_N.t695 1.1255
R13869 VDAC_N.n2084 VDAC_N.t1402 1.1255
R13870 VDAC_N.n2085 VDAC_N.t1181 1.1255
R13871 VDAC_N.n2086 VDAC_N.t1755 1.1255
R13872 VDAC_N.n2087 VDAC_N.t1070 1.1255
R13873 VDAC_N.n2088 VDAC_N.t783 1.1255
R13874 VDAC_N.n2089 VDAC_N.t1065 1.1255
R13875 VDAC_N.n2090 VDAC_N.t1429 1.1255
R13876 VDAC_N.n2091 VDAC_N.t1891 1.1255
R13877 VDAC_N.n2092 VDAC_N.t1325 1.1255
R13878 VDAC_N.n2093 VDAC_N.t905 1.1255
R13879 VDAC_N.n2094 VDAC_N.t108 1.1255
R13880 VDAC_N.n2095 VDAC_N.t797 1.1255
R13881 VDAC_N.n2096 VDAC_N.t1081 1.1255
R13882 VDAC_N.n2097 VDAC_N.t1776 1.1255
R13883 VDAC_N.n2098 VDAC_N.t973 1.1255
R13884 VDAC_N.n2099 VDAC_N.t1320 1.1255
R13885 VDAC_N.n2100 VDAC_N.t251 1.1255
R13886 VDAC_N.n2101 VDAC_N.t1740 1.1255
R13887 VDAC_N.n2102 VDAC_N.t70 1.1255
R13888 VDAC_N.n2103 VDAC_N.t668 1.1255
R13889 VDAC_N.n2104 VDAC_N.t1888 1.1255
R13890 VDAC_N.n2105 VDAC_N.t1882 1.1255
R13891 VDAC_N.n2106 VDAC_N.t736 1.1255
R13892 VDAC_N.n2107 VDAC_N.t130 1.1255
R13893 VDAC_N.n2108 VDAC_N.t292 1.1255
R13894 VDAC_N.n2109 VDAC_N.t1434 1.1255
R13895 VDAC_N.n2110 VDAC_N.t1201 1.1255
R13896 VDAC_N.n2111 VDAC_N.t1174 1.1255
R13897 VDAC_N.n2112 VDAC_N.t1175 1.1255
R13898 VDAC_N.n2113 VDAC_N.t1641 1.1255
R13899 VDAC_N.n2114 VDAC_N.t1898 1.1255
R13900 VDAC_N.n2115 VDAC_N.t725 1.1255
R13901 VDAC_N.n2116 VDAC_N.t1987 1.1255
R13902 VDAC_N.n2117 VDAC_N.t1319 1.1255
R13903 VDAC_N.n2118 VDAC_N.t901 1.1255
R13904 VDAC_N.n2119 VDAC_N.t617 1.1255
R13905 VDAC_N.n2120 VDAC_N.t849 1.1255
R13906 VDAC_N.n2121 VDAC_N.t553 1.1255
R13907 VDAC_N.n2122 VDAC_N.t411 1.1255
R13908 VDAC_N.n2123 VDAC_N.t525 1.1255
R13909 VDAC_N.n2124 VDAC_N.t1296 1.1255
R13910 VDAC_N.n2125 VDAC_N.t1805 1.1255
R13911 VDAC_N.n2126 VDAC_N.t1716 1.1255
R13912 VDAC_N.n2127 VDAC_N.t447 1.1255
R13913 VDAC_N.n2128 VDAC_N.t604 1.1255
R13914 VDAC_N.n2129 VDAC_N.t1154 1.1255
R13915 VDAC_N.n2130 VDAC_N.t1039 1.1255
R13916 VDAC_N.n2131 VDAC_N.t720 1.1255
R13917 VDAC_N.n2132 VDAC_N.t1866 1.1255
R13918 VDAC_N.n2133 VDAC_N.t996 1.1255
R13919 VDAC_N.n2134 VDAC_N.t202 1.1255
R13920 VDAC_N.n13 VDAC_N.n9 1.04597
R13921 VDAC_N.n13 VDAC_N.n12 0.929304
R13922 VDAC_N.n1 VDAC_N.n0 0.733109
R13923 VDAC_N.n2 VDAC_N.n1 0.733109
R13924 VDAC_N.n11 VDAC_N.n10 0.733109
R13925 VDAC_N.n12 VDAC_N.n11 0.733109
R13926 VDAC_N.n4 VDAC_N.n3 0.733109
R13927 VDAC_N.n5 VDAC_N.n4 0.733109
R13928 VDAC_N.n7 VDAC_N.n6 0.733109
R13929 VDAC_N.n8 VDAC_N.n7 0.733109
R13930 VDAC_N.n9 VDAC_N.n8 0.733109
R13931 VDAC_N.n21 VDAC_N.n17 0.21925
R13932 VDAC_N.n1944 VDAC_N.n23 0.204167
R13933 VDAC_N.n1945 VDAC_N.n1944 0.204167
R13934 VDAC_N.n1946 VDAC_N.n1945 0.204167
R13935 VDAC_N.n1947 VDAC_N.n1946 0.204167
R13936 VDAC_N.n1948 VDAC_N.n1947 0.204167
R13937 VDAC_N.n1949 VDAC_N.n1948 0.204167
R13938 VDAC_N.n1950 VDAC_N.n1949 0.204167
R13939 VDAC_N.n1951 VDAC_N.n1950 0.204167
R13940 VDAC_N.n1952 VDAC_N.n1951 0.204167
R13941 VDAC_N.n1953 VDAC_N.n1952 0.204167
R13942 VDAC_N.n1954 VDAC_N.n1953 0.204167
R13943 VDAC_N.n1955 VDAC_N.n1954 0.204167
R13944 VDAC_N.n1956 VDAC_N.n1955 0.204167
R13945 VDAC_N.n1957 VDAC_N.n1956 0.204167
R13946 VDAC_N.n1958 VDAC_N.n1957 0.204167
R13947 VDAC_N.n1959 VDAC_N.n1958 0.204167
R13948 VDAC_N.n1960 VDAC_N.n1959 0.204167
R13949 VDAC_N.n1961 VDAC_N.n1960 0.204167
R13950 VDAC_N.n1962 VDAC_N.n1961 0.204167
R13951 VDAC_N.n1963 VDAC_N.n1962 0.204167
R13952 VDAC_N.n1964 VDAC_N.n1963 0.204167
R13953 VDAC_N.n1965 VDAC_N.n1964 0.204167
R13954 VDAC_N.n1966 VDAC_N.n1965 0.204167
R13955 VDAC_N.n1967 VDAC_N.n1966 0.204167
R13956 VDAC_N.n1968 VDAC_N.n1967 0.204167
R13957 VDAC_N.n1969 VDAC_N.n1968 0.204167
R13958 VDAC_N.n1970 VDAC_N.n1969 0.204167
R13959 VDAC_N.n1971 VDAC_N.n1970 0.204167
R13960 VDAC_N.n1972 VDAC_N.n1971 0.204167
R13961 VDAC_N.n2040 VDAC_N.n2039 0.204167
R13962 VDAC_N.n2041 VDAC_N.n2040 0.204167
R13963 VDAC_N.n2042 VDAC_N.n2041 0.204167
R13964 VDAC_N.n2043 VDAC_N.n2042 0.204167
R13965 VDAC_N.n2044 VDAC_N.n2043 0.204167
R13966 VDAC_N.n2045 VDAC_N.n2044 0.204167
R13967 VDAC_N.n2046 VDAC_N.n2045 0.204167
R13968 VDAC_N.n2047 VDAC_N.n2046 0.204167
R13969 VDAC_N.n2048 VDAC_N.n2047 0.204167
R13970 VDAC_N.n2049 VDAC_N.n2048 0.204167
R13971 VDAC_N.n2050 VDAC_N.n2049 0.204167
R13972 VDAC_N.n2051 VDAC_N.n2050 0.204167
R13973 VDAC_N.n2052 VDAC_N.n2051 0.204167
R13974 VDAC_N.n2053 VDAC_N.n2052 0.204167
R13975 VDAC_N.n2054 VDAC_N.n2053 0.204167
R13976 VDAC_N.n2055 VDAC_N.n2054 0.204167
R13977 VDAC_N.n2056 VDAC_N.n2055 0.204167
R13978 VDAC_N.n2057 VDAC_N.n2056 0.204167
R13979 VDAC_N.n2058 VDAC_N.n2057 0.204167
R13980 VDAC_N.n2059 VDAC_N.n2058 0.204167
R13981 VDAC_N.n2060 VDAC_N.n2059 0.204167
R13982 VDAC_N.n2061 VDAC_N.n2060 0.204167
R13983 VDAC_N.n2062 VDAC_N.n2061 0.204167
R13984 VDAC_N.n2063 VDAC_N.n2062 0.204167
R13985 VDAC_N.n2064 VDAC_N.n2063 0.204167
R13986 VDAC_N.n2065 VDAC_N.n2064 0.204167
R13987 VDAC_N.n2066 VDAC_N.n2065 0.204167
R13988 VDAC_N.n2067 VDAC_N.n2066 0.204167
R13989 VDAC_N.n2068 VDAC_N.n2067 0.204167
R13990 VDAC_N.n21 VDAC_N.n20 0.188
R13991 VDAC_N.n117 VDAC_N.n116 0.180667
R13992 VDAC_N.n118 VDAC_N.n117 0.180667
R13993 VDAC_N.n119 VDAC_N.n118 0.180667
R13994 VDAC_N.n120 VDAC_N.n119 0.180667
R13995 VDAC_N.n121 VDAC_N.n120 0.180667
R13996 VDAC_N.n122 VDAC_N.n121 0.180667
R13997 VDAC_N.n123 VDAC_N.n122 0.180667
R13998 VDAC_N.n124 VDAC_N.n123 0.180667
R13999 VDAC_N.n125 VDAC_N.n124 0.180667
R14000 VDAC_N.n126 VDAC_N.n125 0.180667
R14001 VDAC_N.n127 VDAC_N.n126 0.180667
R14002 VDAC_N.n128 VDAC_N.n127 0.180667
R14003 VDAC_N.n129 VDAC_N.n128 0.180667
R14004 VDAC_N.n130 VDAC_N.n129 0.180667
R14005 VDAC_N.n131 VDAC_N.n130 0.180667
R14006 VDAC_N.n132 VDAC_N.n131 0.180667
R14007 VDAC_N.n133 VDAC_N.n132 0.180667
R14008 VDAC_N.n134 VDAC_N.n133 0.180667
R14009 VDAC_N.n135 VDAC_N.n134 0.180667
R14010 VDAC_N.n136 VDAC_N.n135 0.180667
R14011 VDAC_N.n137 VDAC_N.n136 0.180667
R14012 VDAC_N.n138 VDAC_N.n137 0.180667
R14013 VDAC_N.n139 VDAC_N.n138 0.180667
R14014 VDAC_N.n140 VDAC_N.n139 0.180667
R14015 VDAC_N.n141 VDAC_N.n140 0.180667
R14016 VDAC_N.n142 VDAC_N.n141 0.180667
R14017 VDAC_N.n143 VDAC_N.n142 0.180667
R14018 VDAC_N.n144 VDAC_N.n143 0.180667
R14019 VDAC_N.n145 VDAC_N.n144 0.180667
R14020 VDAC_N.n146 VDAC_N.n145 0.180667
R14021 VDAC_N.n147 VDAC_N.n146 0.180667
R14022 VDAC_N.n148 VDAC_N.n147 0.180667
R14023 VDAC_N.n149 VDAC_N.n148 0.180667
R14024 VDAC_N.n150 VDAC_N.n149 0.180667
R14025 VDAC_N.n151 VDAC_N.n150 0.180667
R14026 VDAC_N.n152 VDAC_N.n151 0.180667
R14027 VDAC_N.n153 VDAC_N.n152 0.180667
R14028 VDAC_N.n154 VDAC_N.n153 0.180667
R14029 VDAC_N.n155 VDAC_N.n154 0.180667
R14030 VDAC_N.n156 VDAC_N.n155 0.180667
R14031 VDAC_N.n157 VDAC_N.n156 0.180667
R14032 VDAC_N.n158 VDAC_N.n157 0.180667
R14033 VDAC_N.n159 VDAC_N.n158 0.180667
R14034 VDAC_N.n160 VDAC_N.n159 0.180667
R14035 VDAC_N.n161 VDAC_N.n160 0.180667
R14036 VDAC_N.n162 VDAC_N.n161 0.180667
R14037 VDAC_N.n163 VDAC_N.n162 0.180667
R14038 VDAC_N.n164 VDAC_N.n163 0.180667
R14039 VDAC_N.n165 VDAC_N.n164 0.180667
R14040 VDAC_N.n166 VDAC_N.n165 0.180667
R14041 VDAC_N.n167 VDAC_N.n166 0.180667
R14042 VDAC_N.n168 VDAC_N.n167 0.180667
R14043 VDAC_N.n169 VDAC_N.n168 0.180667
R14044 VDAC_N.n170 VDAC_N.n169 0.180667
R14045 VDAC_N.n171 VDAC_N.n170 0.180667
R14046 VDAC_N.n172 VDAC_N.n171 0.180667
R14047 VDAC_N.n173 VDAC_N.n172 0.180667
R14048 VDAC_N.n174 VDAC_N.n173 0.180667
R14049 VDAC_N.n175 VDAC_N.n174 0.180667
R14050 VDAC_N.n176 VDAC_N.n175 0.180667
R14051 VDAC_N.n177 VDAC_N.n176 0.180667
R14052 VDAC_N.n178 VDAC_N.n177 0.180667
R14053 VDAC_N.n179 VDAC_N.n178 0.180667
R14054 VDAC_N.n180 VDAC_N.n115 0.180667
R14055 VDAC_N.n181 VDAC_N.n180 0.180667
R14056 VDAC_N.n182 VDAC_N.n181 0.180667
R14057 VDAC_N.n183 VDAC_N.n182 0.180667
R14058 VDAC_N.n184 VDAC_N.n183 0.180667
R14059 VDAC_N.n185 VDAC_N.n184 0.180667
R14060 VDAC_N.n186 VDAC_N.n185 0.180667
R14061 VDAC_N.n187 VDAC_N.n186 0.180667
R14062 VDAC_N.n188 VDAC_N.n187 0.180667
R14063 VDAC_N.n189 VDAC_N.n188 0.180667
R14064 VDAC_N.n190 VDAC_N.n189 0.180667
R14065 VDAC_N.n191 VDAC_N.n190 0.180667
R14066 VDAC_N.n192 VDAC_N.n191 0.180667
R14067 VDAC_N.n193 VDAC_N.n192 0.180667
R14068 VDAC_N.n194 VDAC_N.n193 0.180667
R14069 VDAC_N.n195 VDAC_N.n194 0.180667
R14070 VDAC_N.n196 VDAC_N.n195 0.180667
R14071 VDAC_N.n197 VDAC_N.n196 0.180667
R14072 VDAC_N.n198 VDAC_N.n197 0.180667
R14073 VDAC_N.n199 VDAC_N.n198 0.180667
R14074 VDAC_N.n200 VDAC_N.n199 0.180667
R14075 VDAC_N.n201 VDAC_N.n200 0.180667
R14076 VDAC_N.n202 VDAC_N.n201 0.180667
R14077 VDAC_N.n203 VDAC_N.n202 0.180667
R14078 VDAC_N.n204 VDAC_N.n203 0.180667
R14079 VDAC_N.n205 VDAC_N.n204 0.180667
R14080 VDAC_N.n206 VDAC_N.n205 0.180667
R14081 VDAC_N.n207 VDAC_N.n206 0.180667
R14082 VDAC_N.n208 VDAC_N.n207 0.180667
R14083 VDAC_N.n209 VDAC_N.n208 0.180667
R14084 VDAC_N.n210 VDAC_N.n209 0.180667
R14085 VDAC_N.n211 VDAC_N.n210 0.180667
R14086 VDAC_N.n212 VDAC_N.n211 0.180667
R14087 VDAC_N.n213 VDAC_N.n212 0.180667
R14088 VDAC_N.n214 VDAC_N.n213 0.180667
R14089 VDAC_N.n215 VDAC_N.n214 0.180667
R14090 VDAC_N.n216 VDAC_N.n215 0.180667
R14091 VDAC_N.n217 VDAC_N.n216 0.180667
R14092 VDAC_N.n218 VDAC_N.n217 0.180667
R14093 VDAC_N.n219 VDAC_N.n218 0.180667
R14094 VDAC_N.n220 VDAC_N.n219 0.180667
R14095 VDAC_N.n221 VDAC_N.n220 0.180667
R14096 VDAC_N.n222 VDAC_N.n221 0.180667
R14097 VDAC_N.n223 VDAC_N.n222 0.180667
R14098 VDAC_N.n224 VDAC_N.n223 0.180667
R14099 VDAC_N.n225 VDAC_N.n224 0.180667
R14100 VDAC_N.n226 VDAC_N.n225 0.180667
R14101 VDAC_N.n227 VDAC_N.n226 0.180667
R14102 VDAC_N.n228 VDAC_N.n227 0.180667
R14103 VDAC_N.n229 VDAC_N.n228 0.180667
R14104 VDAC_N.n230 VDAC_N.n229 0.180667
R14105 VDAC_N.n231 VDAC_N.n230 0.180667
R14106 VDAC_N.n232 VDAC_N.n231 0.180667
R14107 VDAC_N.n233 VDAC_N.n232 0.180667
R14108 VDAC_N.n234 VDAC_N.n233 0.180667
R14109 VDAC_N.n235 VDAC_N.n234 0.180667
R14110 VDAC_N.n236 VDAC_N.n235 0.180667
R14111 VDAC_N.n237 VDAC_N.n236 0.180667
R14112 VDAC_N.n238 VDAC_N.n237 0.180667
R14113 VDAC_N.n239 VDAC_N.n238 0.180667
R14114 VDAC_N.n240 VDAC_N.n239 0.180667
R14115 VDAC_N.n241 VDAC_N.n240 0.180667
R14116 VDAC_N.n242 VDAC_N.n241 0.180667
R14117 VDAC_N.n243 VDAC_N.n114 0.180667
R14118 VDAC_N.n244 VDAC_N.n243 0.180667
R14119 VDAC_N.n245 VDAC_N.n244 0.180667
R14120 VDAC_N.n246 VDAC_N.n245 0.180667
R14121 VDAC_N.n247 VDAC_N.n246 0.180667
R14122 VDAC_N.n248 VDAC_N.n247 0.180667
R14123 VDAC_N.n249 VDAC_N.n248 0.180667
R14124 VDAC_N.n250 VDAC_N.n249 0.180667
R14125 VDAC_N.n251 VDAC_N.n250 0.180667
R14126 VDAC_N.n252 VDAC_N.n251 0.180667
R14127 VDAC_N.n253 VDAC_N.n252 0.180667
R14128 VDAC_N.n254 VDAC_N.n253 0.180667
R14129 VDAC_N.n255 VDAC_N.n254 0.180667
R14130 VDAC_N.n256 VDAC_N.n255 0.180667
R14131 VDAC_N.n257 VDAC_N.n256 0.180667
R14132 VDAC_N.n258 VDAC_N.n257 0.180667
R14133 VDAC_N.n259 VDAC_N.n258 0.180667
R14134 VDAC_N.n260 VDAC_N.n259 0.180667
R14135 VDAC_N.n261 VDAC_N.n260 0.180667
R14136 VDAC_N.n262 VDAC_N.n261 0.180667
R14137 VDAC_N.n263 VDAC_N.n262 0.180667
R14138 VDAC_N.n264 VDAC_N.n263 0.180667
R14139 VDAC_N.n265 VDAC_N.n264 0.180667
R14140 VDAC_N.n266 VDAC_N.n265 0.180667
R14141 VDAC_N.n267 VDAC_N.n266 0.180667
R14142 VDAC_N.n268 VDAC_N.n267 0.180667
R14143 VDAC_N.n269 VDAC_N.n268 0.180667
R14144 VDAC_N.n270 VDAC_N.n269 0.180667
R14145 VDAC_N.n271 VDAC_N.n270 0.180667
R14146 VDAC_N.n272 VDAC_N.n271 0.180667
R14147 VDAC_N.n273 VDAC_N.n272 0.180667
R14148 VDAC_N.n274 VDAC_N.n273 0.180667
R14149 VDAC_N.n275 VDAC_N.n274 0.180667
R14150 VDAC_N.n276 VDAC_N.n275 0.180667
R14151 VDAC_N.n277 VDAC_N.n276 0.180667
R14152 VDAC_N.n278 VDAC_N.n277 0.180667
R14153 VDAC_N.n279 VDAC_N.n278 0.180667
R14154 VDAC_N.n280 VDAC_N.n279 0.180667
R14155 VDAC_N.n281 VDAC_N.n280 0.180667
R14156 VDAC_N.n282 VDAC_N.n281 0.180667
R14157 VDAC_N.n283 VDAC_N.n282 0.180667
R14158 VDAC_N.n284 VDAC_N.n283 0.180667
R14159 VDAC_N.n285 VDAC_N.n284 0.180667
R14160 VDAC_N.n286 VDAC_N.n285 0.180667
R14161 VDAC_N.n287 VDAC_N.n286 0.180667
R14162 VDAC_N.n288 VDAC_N.n287 0.180667
R14163 VDAC_N.n289 VDAC_N.n288 0.180667
R14164 VDAC_N.n290 VDAC_N.n289 0.180667
R14165 VDAC_N.n291 VDAC_N.n290 0.180667
R14166 VDAC_N.n292 VDAC_N.n291 0.180667
R14167 VDAC_N.n293 VDAC_N.n292 0.180667
R14168 VDAC_N.n294 VDAC_N.n293 0.180667
R14169 VDAC_N.n295 VDAC_N.n294 0.180667
R14170 VDAC_N.n296 VDAC_N.n295 0.180667
R14171 VDAC_N.n297 VDAC_N.n296 0.180667
R14172 VDAC_N.n298 VDAC_N.n297 0.180667
R14173 VDAC_N.n299 VDAC_N.n298 0.180667
R14174 VDAC_N.n300 VDAC_N.n299 0.180667
R14175 VDAC_N.n301 VDAC_N.n300 0.180667
R14176 VDAC_N.n302 VDAC_N.n301 0.180667
R14177 VDAC_N.n303 VDAC_N.n302 0.180667
R14178 VDAC_N.n304 VDAC_N.n303 0.180667
R14179 VDAC_N.n305 VDAC_N.n304 0.180667
R14180 VDAC_N.n306 VDAC_N.n113 0.180667
R14181 VDAC_N.n307 VDAC_N.n306 0.180667
R14182 VDAC_N.n308 VDAC_N.n307 0.180667
R14183 VDAC_N.n309 VDAC_N.n308 0.180667
R14184 VDAC_N.n310 VDAC_N.n309 0.180667
R14185 VDAC_N.n311 VDAC_N.n310 0.180667
R14186 VDAC_N.n312 VDAC_N.n311 0.180667
R14187 VDAC_N.n313 VDAC_N.n312 0.180667
R14188 VDAC_N.n314 VDAC_N.n313 0.180667
R14189 VDAC_N.n315 VDAC_N.n314 0.180667
R14190 VDAC_N.n316 VDAC_N.n315 0.180667
R14191 VDAC_N.n317 VDAC_N.n316 0.180667
R14192 VDAC_N.n318 VDAC_N.n317 0.180667
R14193 VDAC_N.n319 VDAC_N.n318 0.180667
R14194 VDAC_N.n320 VDAC_N.n319 0.180667
R14195 VDAC_N.n321 VDAC_N.n320 0.180667
R14196 VDAC_N.n322 VDAC_N.n321 0.180667
R14197 VDAC_N.n323 VDAC_N.n322 0.180667
R14198 VDAC_N.n324 VDAC_N.n323 0.180667
R14199 VDAC_N.n325 VDAC_N.n324 0.180667
R14200 VDAC_N.n326 VDAC_N.n325 0.180667
R14201 VDAC_N.n327 VDAC_N.n326 0.180667
R14202 VDAC_N.n328 VDAC_N.n327 0.180667
R14203 VDAC_N.n329 VDAC_N.n328 0.180667
R14204 VDAC_N.n330 VDAC_N.n329 0.180667
R14205 VDAC_N.n331 VDAC_N.n330 0.180667
R14206 VDAC_N.n332 VDAC_N.n331 0.180667
R14207 VDAC_N.n333 VDAC_N.n332 0.180667
R14208 VDAC_N.n334 VDAC_N.n333 0.180667
R14209 VDAC_N.n335 VDAC_N.n334 0.180667
R14210 VDAC_N.n336 VDAC_N.n335 0.180667
R14211 VDAC_N.n337 VDAC_N.n336 0.180667
R14212 VDAC_N.n338 VDAC_N.n337 0.180667
R14213 VDAC_N.n339 VDAC_N.n338 0.180667
R14214 VDAC_N.n340 VDAC_N.n339 0.180667
R14215 VDAC_N.n341 VDAC_N.n340 0.180667
R14216 VDAC_N.n342 VDAC_N.n341 0.180667
R14217 VDAC_N.n343 VDAC_N.n342 0.180667
R14218 VDAC_N.n344 VDAC_N.n343 0.180667
R14219 VDAC_N.n345 VDAC_N.n344 0.180667
R14220 VDAC_N.n346 VDAC_N.n345 0.180667
R14221 VDAC_N.n347 VDAC_N.n346 0.180667
R14222 VDAC_N.n348 VDAC_N.n347 0.180667
R14223 VDAC_N.n349 VDAC_N.n348 0.180667
R14224 VDAC_N.n350 VDAC_N.n349 0.180667
R14225 VDAC_N.n351 VDAC_N.n350 0.180667
R14226 VDAC_N.n352 VDAC_N.n351 0.180667
R14227 VDAC_N.n353 VDAC_N.n352 0.180667
R14228 VDAC_N.n354 VDAC_N.n353 0.180667
R14229 VDAC_N.n355 VDAC_N.n354 0.180667
R14230 VDAC_N.n356 VDAC_N.n355 0.180667
R14231 VDAC_N.n357 VDAC_N.n356 0.180667
R14232 VDAC_N.n358 VDAC_N.n357 0.180667
R14233 VDAC_N.n359 VDAC_N.n358 0.180667
R14234 VDAC_N.n360 VDAC_N.n359 0.180667
R14235 VDAC_N.n361 VDAC_N.n360 0.180667
R14236 VDAC_N.n362 VDAC_N.n361 0.180667
R14237 VDAC_N.n363 VDAC_N.n362 0.180667
R14238 VDAC_N.n364 VDAC_N.n363 0.180667
R14239 VDAC_N.n365 VDAC_N.n364 0.180667
R14240 VDAC_N.n366 VDAC_N.n365 0.180667
R14241 VDAC_N.n367 VDAC_N.n366 0.180667
R14242 VDAC_N.n368 VDAC_N.n367 0.180667
R14243 VDAC_N.n369 VDAC_N.n112 0.180667
R14244 VDAC_N.n370 VDAC_N.n369 0.180667
R14245 VDAC_N.n371 VDAC_N.n370 0.180667
R14246 VDAC_N.n372 VDAC_N.n371 0.180667
R14247 VDAC_N.n373 VDAC_N.n372 0.180667
R14248 VDAC_N.n374 VDAC_N.n373 0.180667
R14249 VDAC_N.n375 VDAC_N.n374 0.180667
R14250 VDAC_N.n376 VDAC_N.n375 0.180667
R14251 VDAC_N.n377 VDAC_N.n376 0.180667
R14252 VDAC_N.n378 VDAC_N.n377 0.180667
R14253 VDAC_N.n379 VDAC_N.n378 0.180667
R14254 VDAC_N.n380 VDAC_N.n379 0.180667
R14255 VDAC_N.n381 VDAC_N.n380 0.180667
R14256 VDAC_N.n382 VDAC_N.n381 0.180667
R14257 VDAC_N.n383 VDAC_N.n382 0.180667
R14258 VDAC_N.n384 VDAC_N.n383 0.180667
R14259 VDAC_N.n385 VDAC_N.n384 0.180667
R14260 VDAC_N.n386 VDAC_N.n385 0.180667
R14261 VDAC_N.n387 VDAC_N.n386 0.180667
R14262 VDAC_N.n388 VDAC_N.n387 0.180667
R14263 VDAC_N.n389 VDAC_N.n388 0.180667
R14264 VDAC_N.n390 VDAC_N.n389 0.180667
R14265 VDAC_N.n391 VDAC_N.n390 0.180667
R14266 VDAC_N.n392 VDAC_N.n391 0.180667
R14267 VDAC_N.n393 VDAC_N.n392 0.180667
R14268 VDAC_N.n394 VDAC_N.n393 0.180667
R14269 VDAC_N.n395 VDAC_N.n394 0.180667
R14270 VDAC_N.n396 VDAC_N.n395 0.180667
R14271 VDAC_N.n397 VDAC_N.n396 0.180667
R14272 VDAC_N.n398 VDAC_N.n397 0.180667
R14273 VDAC_N.n399 VDAC_N.n398 0.180667
R14274 VDAC_N.n400 VDAC_N.n399 0.180667
R14275 VDAC_N.n401 VDAC_N.n400 0.180667
R14276 VDAC_N.n402 VDAC_N.n401 0.180667
R14277 VDAC_N.n403 VDAC_N.n402 0.180667
R14278 VDAC_N.n404 VDAC_N.n403 0.180667
R14279 VDAC_N.n405 VDAC_N.n404 0.180667
R14280 VDAC_N.n406 VDAC_N.n405 0.180667
R14281 VDAC_N.n407 VDAC_N.n406 0.180667
R14282 VDAC_N.n408 VDAC_N.n407 0.180667
R14283 VDAC_N.n409 VDAC_N.n408 0.180667
R14284 VDAC_N.n410 VDAC_N.n409 0.180667
R14285 VDAC_N.n411 VDAC_N.n410 0.180667
R14286 VDAC_N.n412 VDAC_N.n411 0.180667
R14287 VDAC_N.n413 VDAC_N.n412 0.180667
R14288 VDAC_N.n414 VDAC_N.n413 0.180667
R14289 VDAC_N.n415 VDAC_N.n414 0.180667
R14290 VDAC_N.n416 VDAC_N.n415 0.180667
R14291 VDAC_N.n417 VDAC_N.n416 0.180667
R14292 VDAC_N.n418 VDAC_N.n417 0.180667
R14293 VDAC_N.n419 VDAC_N.n418 0.180667
R14294 VDAC_N.n420 VDAC_N.n419 0.180667
R14295 VDAC_N.n421 VDAC_N.n420 0.180667
R14296 VDAC_N.n422 VDAC_N.n421 0.180667
R14297 VDAC_N.n423 VDAC_N.n422 0.180667
R14298 VDAC_N.n424 VDAC_N.n423 0.180667
R14299 VDAC_N.n425 VDAC_N.n424 0.180667
R14300 VDAC_N.n426 VDAC_N.n425 0.180667
R14301 VDAC_N.n427 VDAC_N.n426 0.180667
R14302 VDAC_N.n428 VDAC_N.n427 0.180667
R14303 VDAC_N.n429 VDAC_N.n428 0.180667
R14304 VDAC_N.n430 VDAC_N.n429 0.180667
R14305 VDAC_N.n431 VDAC_N.n430 0.180667
R14306 VDAC_N.n432 VDAC_N.n111 0.180667
R14307 VDAC_N.n433 VDAC_N.n432 0.180667
R14308 VDAC_N.n434 VDAC_N.n433 0.180667
R14309 VDAC_N.n435 VDAC_N.n434 0.180667
R14310 VDAC_N.n436 VDAC_N.n435 0.180667
R14311 VDAC_N.n437 VDAC_N.n436 0.180667
R14312 VDAC_N.n438 VDAC_N.n437 0.180667
R14313 VDAC_N.n439 VDAC_N.n438 0.180667
R14314 VDAC_N.n440 VDAC_N.n439 0.180667
R14315 VDAC_N.n441 VDAC_N.n440 0.180667
R14316 VDAC_N.n442 VDAC_N.n441 0.180667
R14317 VDAC_N.n443 VDAC_N.n442 0.180667
R14318 VDAC_N.n444 VDAC_N.n443 0.180667
R14319 VDAC_N.n445 VDAC_N.n444 0.180667
R14320 VDAC_N.n446 VDAC_N.n445 0.180667
R14321 VDAC_N.n447 VDAC_N.n446 0.180667
R14322 VDAC_N.n448 VDAC_N.n447 0.180667
R14323 VDAC_N.n449 VDAC_N.n448 0.180667
R14324 VDAC_N.n450 VDAC_N.n449 0.180667
R14325 VDAC_N.n451 VDAC_N.n450 0.180667
R14326 VDAC_N.n452 VDAC_N.n451 0.180667
R14327 VDAC_N.n453 VDAC_N.n452 0.180667
R14328 VDAC_N.n454 VDAC_N.n453 0.180667
R14329 VDAC_N.n455 VDAC_N.n454 0.180667
R14330 VDAC_N.n456 VDAC_N.n455 0.180667
R14331 VDAC_N.n457 VDAC_N.n456 0.180667
R14332 VDAC_N.n458 VDAC_N.n457 0.180667
R14333 VDAC_N.n459 VDAC_N.n458 0.180667
R14334 VDAC_N.n460 VDAC_N.n459 0.180667
R14335 VDAC_N.n461 VDAC_N.n460 0.180667
R14336 VDAC_N.n462 VDAC_N.n461 0.180667
R14337 VDAC_N.n463 VDAC_N.n462 0.180667
R14338 VDAC_N.n464 VDAC_N.n463 0.180667
R14339 VDAC_N.n465 VDAC_N.n464 0.180667
R14340 VDAC_N.n466 VDAC_N.n465 0.180667
R14341 VDAC_N.n467 VDAC_N.n466 0.180667
R14342 VDAC_N.n468 VDAC_N.n467 0.180667
R14343 VDAC_N.n469 VDAC_N.n468 0.180667
R14344 VDAC_N.n470 VDAC_N.n469 0.180667
R14345 VDAC_N.n471 VDAC_N.n470 0.180667
R14346 VDAC_N.n472 VDAC_N.n471 0.180667
R14347 VDAC_N.n473 VDAC_N.n472 0.180667
R14348 VDAC_N.n474 VDAC_N.n473 0.180667
R14349 VDAC_N.n475 VDAC_N.n474 0.180667
R14350 VDAC_N.n476 VDAC_N.n475 0.180667
R14351 VDAC_N.n477 VDAC_N.n476 0.180667
R14352 VDAC_N.n478 VDAC_N.n477 0.180667
R14353 VDAC_N.n479 VDAC_N.n478 0.180667
R14354 VDAC_N.n480 VDAC_N.n479 0.180667
R14355 VDAC_N.n481 VDAC_N.n480 0.180667
R14356 VDAC_N.n482 VDAC_N.n481 0.180667
R14357 VDAC_N.n483 VDAC_N.n482 0.180667
R14358 VDAC_N.n484 VDAC_N.n483 0.180667
R14359 VDAC_N.n485 VDAC_N.n484 0.180667
R14360 VDAC_N.n486 VDAC_N.n485 0.180667
R14361 VDAC_N.n487 VDAC_N.n486 0.180667
R14362 VDAC_N.n488 VDAC_N.n487 0.180667
R14363 VDAC_N.n489 VDAC_N.n488 0.180667
R14364 VDAC_N.n490 VDAC_N.n489 0.180667
R14365 VDAC_N.n491 VDAC_N.n490 0.180667
R14366 VDAC_N.n492 VDAC_N.n491 0.180667
R14367 VDAC_N.n493 VDAC_N.n492 0.180667
R14368 VDAC_N.n494 VDAC_N.n493 0.180667
R14369 VDAC_N.n495 VDAC_N.n110 0.180667
R14370 VDAC_N.n496 VDAC_N.n495 0.180667
R14371 VDAC_N.n497 VDAC_N.n496 0.180667
R14372 VDAC_N.n498 VDAC_N.n497 0.180667
R14373 VDAC_N.n499 VDAC_N.n498 0.180667
R14374 VDAC_N.n500 VDAC_N.n499 0.180667
R14375 VDAC_N.n501 VDAC_N.n500 0.180667
R14376 VDAC_N.n502 VDAC_N.n501 0.180667
R14377 VDAC_N.n503 VDAC_N.n502 0.180667
R14378 VDAC_N.n504 VDAC_N.n503 0.180667
R14379 VDAC_N.n505 VDAC_N.n504 0.180667
R14380 VDAC_N.n506 VDAC_N.n505 0.180667
R14381 VDAC_N.n507 VDAC_N.n506 0.180667
R14382 VDAC_N.n508 VDAC_N.n507 0.180667
R14383 VDAC_N.n509 VDAC_N.n508 0.180667
R14384 VDAC_N.n510 VDAC_N.n509 0.180667
R14385 VDAC_N.n511 VDAC_N.n510 0.180667
R14386 VDAC_N.n512 VDAC_N.n511 0.180667
R14387 VDAC_N.n513 VDAC_N.n512 0.180667
R14388 VDAC_N.n514 VDAC_N.n513 0.180667
R14389 VDAC_N.n515 VDAC_N.n514 0.180667
R14390 VDAC_N.n516 VDAC_N.n515 0.180667
R14391 VDAC_N.n517 VDAC_N.n516 0.180667
R14392 VDAC_N.n518 VDAC_N.n517 0.180667
R14393 VDAC_N.n519 VDAC_N.n518 0.180667
R14394 VDAC_N.n520 VDAC_N.n519 0.180667
R14395 VDAC_N.n521 VDAC_N.n520 0.180667
R14396 VDAC_N.n522 VDAC_N.n521 0.180667
R14397 VDAC_N.n523 VDAC_N.n522 0.180667
R14398 VDAC_N.n524 VDAC_N.n523 0.180667
R14399 VDAC_N.n525 VDAC_N.n524 0.180667
R14400 VDAC_N.n526 VDAC_N.n525 0.180667
R14401 VDAC_N.n527 VDAC_N.n526 0.180667
R14402 VDAC_N.n528 VDAC_N.n527 0.180667
R14403 VDAC_N.n529 VDAC_N.n528 0.180667
R14404 VDAC_N.n530 VDAC_N.n529 0.180667
R14405 VDAC_N.n531 VDAC_N.n530 0.180667
R14406 VDAC_N.n532 VDAC_N.n531 0.180667
R14407 VDAC_N.n533 VDAC_N.n532 0.180667
R14408 VDAC_N.n534 VDAC_N.n533 0.180667
R14409 VDAC_N.n535 VDAC_N.n534 0.180667
R14410 VDAC_N.n536 VDAC_N.n535 0.180667
R14411 VDAC_N.n537 VDAC_N.n536 0.180667
R14412 VDAC_N.n538 VDAC_N.n537 0.180667
R14413 VDAC_N.n539 VDAC_N.n538 0.180667
R14414 VDAC_N.n540 VDAC_N.n539 0.180667
R14415 VDAC_N.n541 VDAC_N.n540 0.180667
R14416 VDAC_N.n542 VDAC_N.n541 0.180667
R14417 VDAC_N.n543 VDAC_N.n542 0.180667
R14418 VDAC_N.n544 VDAC_N.n543 0.180667
R14419 VDAC_N.n545 VDAC_N.n544 0.180667
R14420 VDAC_N.n546 VDAC_N.n545 0.180667
R14421 VDAC_N.n547 VDAC_N.n546 0.180667
R14422 VDAC_N.n548 VDAC_N.n547 0.180667
R14423 VDAC_N.n549 VDAC_N.n548 0.180667
R14424 VDAC_N.n550 VDAC_N.n549 0.180667
R14425 VDAC_N.n551 VDAC_N.n550 0.180667
R14426 VDAC_N.n552 VDAC_N.n551 0.180667
R14427 VDAC_N.n553 VDAC_N.n552 0.180667
R14428 VDAC_N.n554 VDAC_N.n553 0.180667
R14429 VDAC_N.n555 VDAC_N.n554 0.180667
R14430 VDAC_N.n556 VDAC_N.n555 0.180667
R14431 VDAC_N.n557 VDAC_N.n556 0.180667
R14432 VDAC_N.n558 VDAC_N.n109 0.180667
R14433 VDAC_N.n559 VDAC_N.n558 0.180667
R14434 VDAC_N.n560 VDAC_N.n559 0.180667
R14435 VDAC_N.n561 VDAC_N.n560 0.180667
R14436 VDAC_N.n562 VDAC_N.n561 0.180667
R14437 VDAC_N.n563 VDAC_N.n562 0.180667
R14438 VDAC_N.n564 VDAC_N.n563 0.180667
R14439 VDAC_N.n565 VDAC_N.n564 0.180667
R14440 VDAC_N.n566 VDAC_N.n565 0.180667
R14441 VDAC_N.n567 VDAC_N.n566 0.180667
R14442 VDAC_N.n568 VDAC_N.n567 0.180667
R14443 VDAC_N.n569 VDAC_N.n568 0.180667
R14444 VDAC_N.n570 VDAC_N.n569 0.180667
R14445 VDAC_N.n571 VDAC_N.n570 0.180667
R14446 VDAC_N.n572 VDAC_N.n571 0.180667
R14447 VDAC_N.n573 VDAC_N.n572 0.180667
R14448 VDAC_N.n574 VDAC_N.n573 0.180667
R14449 VDAC_N.n575 VDAC_N.n574 0.180667
R14450 VDAC_N.n576 VDAC_N.n575 0.180667
R14451 VDAC_N.n577 VDAC_N.n576 0.180667
R14452 VDAC_N.n578 VDAC_N.n577 0.180667
R14453 VDAC_N.n579 VDAC_N.n578 0.180667
R14454 VDAC_N.n580 VDAC_N.n579 0.180667
R14455 VDAC_N.n581 VDAC_N.n580 0.180667
R14456 VDAC_N.n582 VDAC_N.n581 0.180667
R14457 VDAC_N.n583 VDAC_N.n582 0.180667
R14458 VDAC_N.n584 VDAC_N.n583 0.180667
R14459 VDAC_N.n585 VDAC_N.n584 0.180667
R14460 VDAC_N.n586 VDAC_N.n585 0.180667
R14461 VDAC_N.n587 VDAC_N.n586 0.180667
R14462 VDAC_N.n588 VDAC_N.n587 0.180667
R14463 VDAC_N.n589 VDAC_N.n588 0.180667
R14464 VDAC_N.n590 VDAC_N.n589 0.180667
R14465 VDAC_N.n591 VDAC_N.n590 0.180667
R14466 VDAC_N.n592 VDAC_N.n591 0.180667
R14467 VDAC_N.n593 VDAC_N.n592 0.180667
R14468 VDAC_N.n594 VDAC_N.n593 0.180667
R14469 VDAC_N.n595 VDAC_N.n594 0.180667
R14470 VDAC_N.n596 VDAC_N.n595 0.180667
R14471 VDAC_N.n597 VDAC_N.n596 0.180667
R14472 VDAC_N.n598 VDAC_N.n597 0.180667
R14473 VDAC_N.n599 VDAC_N.n598 0.180667
R14474 VDAC_N.n600 VDAC_N.n599 0.180667
R14475 VDAC_N.n601 VDAC_N.n600 0.180667
R14476 VDAC_N.n602 VDAC_N.n601 0.180667
R14477 VDAC_N.n603 VDAC_N.n602 0.180667
R14478 VDAC_N.n604 VDAC_N.n603 0.180667
R14479 VDAC_N.n605 VDAC_N.n604 0.180667
R14480 VDAC_N.n606 VDAC_N.n605 0.180667
R14481 VDAC_N.n607 VDAC_N.n606 0.180667
R14482 VDAC_N.n608 VDAC_N.n607 0.180667
R14483 VDAC_N.n609 VDAC_N.n608 0.180667
R14484 VDAC_N.n610 VDAC_N.n609 0.180667
R14485 VDAC_N.n611 VDAC_N.n610 0.180667
R14486 VDAC_N.n612 VDAC_N.n611 0.180667
R14487 VDAC_N.n613 VDAC_N.n612 0.180667
R14488 VDAC_N.n614 VDAC_N.n613 0.180667
R14489 VDAC_N.n615 VDAC_N.n614 0.180667
R14490 VDAC_N.n616 VDAC_N.n615 0.180667
R14491 VDAC_N.n617 VDAC_N.n616 0.180667
R14492 VDAC_N.n618 VDAC_N.n617 0.180667
R14493 VDAC_N.n619 VDAC_N.n618 0.180667
R14494 VDAC_N.n620 VDAC_N.n619 0.180667
R14495 VDAC_N.n621 VDAC_N.n108 0.180667
R14496 VDAC_N.n622 VDAC_N.n621 0.180667
R14497 VDAC_N.n623 VDAC_N.n622 0.180667
R14498 VDAC_N.n624 VDAC_N.n623 0.180667
R14499 VDAC_N.n625 VDAC_N.n624 0.180667
R14500 VDAC_N.n626 VDAC_N.n625 0.180667
R14501 VDAC_N.n627 VDAC_N.n626 0.180667
R14502 VDAC_N.n628 VDAC_N.n627 0.180667
R14503 VDAC_N.n629 VDAC_N.n628 0.180667
R14504 VDAC_N.n630 VDAC_N.n629 0.180667
R14505 VDAC_N.n631 VDAC_N.n630 0.180667
R14506 VDAC_N.n632 VDAC_N.n631 0.180667
R14507 VDAC_N.n633 VDAC_N.n632 0.180667
R14508 VDAC_N.n634 VDAC_N.n633 0.180667
R14509 VDAC_N.n635 VDAC_N.n634 0.180667
R14510 VDAC_N.n636 VDAC_N.n635 0.180667
R14511 VDAC_N.n637 VDAC_N.n636 0.180667
R14512 VDAC_N.n638 VDAC_N.n637 0.180667
R14513 VDAC_N.n639 VDAC_N.n638 0.180667
R14514 VDAC_N.n640 VDAC_N.n639 0.180667
R14515 VDAC_N.n641 VDAC_N.n640 0.180667
R14516 VDAC_N.n642 VDAC_N.n641 0.180667
R14517 VDAC_N.n643 VDAC_N.n642 0.180667
R14518 VDAC_N.n644 VDAC_N.n643 0.180667
R14519 VDAC_N.n645 VDAC_N.n644 0.180667
R14520 VDAC_N.n646 VDAC_N.n645 0.180667
R14521 VDAC_N.n647 VDAC_N.n646 0.180667
R14522 VDAC_N.n648 VDAC_N.n647 0.180667
R14523 VDAC_N.n649 VDAC_N.n648 0.180667
R14524 VDAC_N.n650 VDAC_N.n649 0.180667
R14525 VDAC_N.n651 VDAC_N.n650 0.180667
R14526 VDAC_N.n652 VDAC_N.n651 0.180667
R14527 VDAC_N.n653 VDAC_N.n652 0.180667
R14528 VDAC_N.n654 VDAC_N.n653 0.180667
R14529 VDAC_N.n655 VDAC_N.n654 0.180667
R14530 VDAC_N.n656 VDAC_N.n655 0.180667
R14531 VDAC_N.n657 VDAC_N.n656 0.180667
R14532 VDAC_N.n658 VDAC_N.n657 0.180667
R14533 VDAC_N.n659 VDAC_N.n658 0.180667
R14534 VDAC_N.n660 VDAC_N.n659 0.180667
R14535 VDAC_N.n661 VDAC_N.n660 0.180667
R14536 VDAC_N.n662 VDAC_N.n661 0.180667
R14537 VDAC_N.n663 VDAC_N.n662 0.180667
R14538 VDAC_N.n664 VDAC_N.n663 0.180667
R14539 VDAC_N.n665 VDAC_N.n664 0.180667
R14540 VDAC_N.n666 VDAC_N.n665 0.180667
R14541 VDAC_N.n667 VDAC_N.n666 0.180667
R14542 VDAC_N.n668 VDAC_N.n667 0.180667
R14543 VDAC_N.n669 VDAC_N.n668 0.180667
R14544 VDAC_N.n670 VDAC_N.n669 0.180667
R14545 VDAC_N.n671 VDAC_N.n670 0.180667
R14546 VDAC_N.n672 VDAC_N.n671 0.180667
R14547 VDAC_N.n673 VDAC_N.n672 0.180667
R14548 VDAC_N.n674 VDAC_N.n673 0.180667
R14549 VDAC_N.n675 VDAC_N.n674 0.180667
R14550 VDAC_N.n676 VDAC_N.n675 0.180667
R14551 VDAC_N.n677 VDAC_N.n676 0.180667
R14552 VDAC_N.n678 VDAC_N.n677 0.180667
R14553 VDAC_N.n679 VDAC_N.n678 0.180667
R14554 VDAC_N.n680 VDAC_N.n679 0.180667
R14555 VDAC_N.n681 VDAC_N.n680 0.180667
R14556 VDAC_N.n682 VDAC_N.n681 0.180667
R14557 VDAC_N.n683 VDAC_N.n682 0.180667
R14558 VDAC_N.n684 VDAC_N.n107 0.180667
R14559 VDAC_N.n685 VDAC_N.n684 0.180667
R14560 VDAC_N.n686 VDAC_N.n685 0.180667
R14561 VDAC_N.n687 VDAC_N.n686 0.180667
R14562 VDAC_N.n688 VDAC_N.n687 0.180667
R14563 VDAC_N.n689 VDAC_N.n688 0.180667
R14564 VDAC_N.n690 VDAC_N.n689 0.180667
R14565 VDAC_N.n691 VDAC_N.n690 0.180667
R14566 VDAC_N.n692 VDAC_N.n691 0.180667
R14567 VDAC_N.n693 VDAC_N.n692 0.180667
R14568 VDAC_N.n694 VDAC_N.n693 0.180667
R14569 VDAC_N.n695 VDAC_N.n694 0.180667
R14570 VDAC_N.n696 VDAC_N.n695 0.180667
R14571 VDAC_N.n697 VDAC_N.n696 0.180667
R14572 VDAC_N.n698 VDAC_N.n697 0.180667
R14573 VDAC_N.n699 VDAC_N.n698 0.180667
R14574 VDAC_N.n700 VDAC_N.n699 0.180667
R14575 VDAC_N.n701 VDAC_N.n700 0.180667
R14576 VDAC_N.n702 VDAC_N.n701 0.180667
R14577 VDAC_N.n703 VDAC_N.n702 0.180667
R14578 VDAC_N.n704 VDAC_N.n703 0.180667
R14579 VDAC_N.n705 VDAC_N.n704 0.180667
R14580 VDAC_N.n706 VDAC_N.n705 0.180667
R14581 VDAC_N.n707 VDAC_N.n706 0.180667
R14582 VDAC_N.n708 VDAC_N.n707 0.180667
R14583 VDAC_N.n709 VDAC_N.n708 0.180667
R14584 VDAC_N.n710 VDAC_N.n709 0.180667
R14585 VDAC_N.n711 VDAC_N.n710 0.180667
R14586 VDAC_N.n712 VDAC_N.n711 0.180667
R14587 VDAC_N.n713 VDAC_N.n712 0.180667
R14588 VDAC_N.n714 VDAC_N.n713 0.180667
R14589 VDAC_N.n715 VDAC_N.n714 0.180667
R14590 VDAC_N.n716 VDAC_N.n715 0.180667
R14591 VDAC_N.n717 VDAC_N.n716 0.180667
R14592 VDAC_N.n718 VDAC_N.n717 0.180667
R14593 VDAC_N.n719 VDAC_N.n718 0.180667
R14594 VDAC_N.n720 VDAC_N.n719 0.180667
R14595 VDAC_N.n721 VDAC_N.n720 0.180667
R14596 VDAC_N.n722 VDAC_N.n721 0.180667
R14597 VDAC_N.n723 VDAC_N.n722 0.180667
R14598 VDAC_N.n724 VDAC_N.n723 0.180667
R14599 VDAC_N.n725 VDAC_N.n724 0.180667
R14600 VDAC_N.n726 VDAC_N.n725 0.180667
R14601 VDAC_N.n727 VDAC_N.n726 0.180667
R14602 VDAC_N.n728 VDAC_N.n727 0.180667
R14603 VDAC_N.n729 VDAC_N.n728 0.180667
R14604 VDAC_N.n730 VDAC_N.n729 0.180667
R14605 VDAC_N.n731 VDAC_N.n730 0.180667
R14606 VDAC_N.n732 VDAC_N.n731 0.180667
R14607 VDAC_N.n733 VDAC_N.n732 0.180667
R14608 VDAC_N.n734 VDAC_N.n733 0.180667
R14609 VDAC_N.n735 VDAC_N.n734 0.180667
R14610 VDAC_N.n736 VDAC_N.n735 0.180667
R14611 VDAC_N.n737 VDAC_N.n736 0.180667
R14612 VDAC_N.n738 VDAC_N.n737 0.180667
R14613 VDAC_N.n739 VDAC_N.n738 0.180667
R14614 VDAC_N.n740 VDAC_N.n739 0.180667
R14615 VDAC_N.n741 VDAC_N.n740 0.180667
R14616 VDAC_N.n742 VDAC_N.n741 0.180667
R14617 VDAC_N.n743 VDAC_N.n742 0.180667
R14618 VDAC_N.n744 VDAC_N.n743 0.180667
R14619 VDAC_N.n745 VDAC_N.n744 0.180667
R14620 VDAC_N.n746 VDAC_N.n745 0.180667
R14621 VDAC_N.n747 VDAC_N.n106 0.180667
R14622 VDAC_N.n748 VDAC_N.n747 0.180667
R14623 VDAC_N.n749 VDAC_N.n748 0.180667
R14624 VDAC_N.n750 VDAC_N.n749 0.180667
R14625 VDAC_N.n751 VDAC_N.n750 0.180667
R14626 VDAC_N.n752 VDAC_N.n751 0.180667
R14627 VDAC_N.n753 VDAC_N.n752 0.180667
R14628 VDAC_N.n754 VDAC_N.n753 0.180667
R14629 VDAC_N.n755 VDAC_N.n754 0.180667
R14630 VDAC_N.n756 VDAC_N.n755 0.180667
R14631 VDAC_N.n757 VDAC_N.n756 0.180667
R14632 VDAC_N.n758 VDAC_N.n757 0.180667
R14633 VDAC_N.n759 VDAC_N.n758 0.180667
R14634 VDAC_N.n760 VDAC_N.n759 0.180667
R14635 VDAC_N.n761 VDAC_N.n760 0.180667
R14636 VDAC_N.n762 VDAC_N.n761 0.180667
R14637 VDAC_N.n763 VDAC_N.n762 0.180667
R14638 VDAC_N.n764 VDAC_N.n763 0.180667
R14639 VDAC_N.n765 VDAC_N.n764 0.180667
R14640 VDAC_N.n766 VDAC_N.n765 0.180667
R14641 VDAC_N.n767 VDAC_N.n766 0.180667
R14642 VDAC_N.n768 VDAC_N.n767 0.180667
R14643 VDAC_N.n769 VDAC_N.n768 0.180667
R14644 VDAC_N.n770 VDAC_N.n769 0.180667
R14645 VDAC_N.n771 VDAC_N.n770 0.180667
R14646 VDAC_N.n772 VDAC_N.n771 0.180667
R14647 VDAC_N.n773 VDAC_N.n772 0.180667
R14648 VDAC_N.n774 VDAC_N.n773 0.180667
R14649 VDAC_N.n775 VDAC_N.n774 0.180667
R14650 VDAC_N.n776 VDAC_N.n775 0.180667
R14651 VDAC_N.n777 VDAC_N.n776 0.180667
R14652 VDAC_N.n778 VDAC_N.n777 0.180667
R14653 VDAC_N.n779 VDAC_N.n778 0.180667
R14654 VDAC_N.n780 VDAC_N.n779 0.180667
R14655 VDAC_N.n781 VDAC_N.n780 0.180667
R14656 VDAC_N.n782 VDAC_N.n781 0.180667
R14657 VDAC_N.n783 VDAC_N.n782 0.180667
R14658 VDAC_N.n784 VDAC_N.n783 0.180667
R14659 VDAC_N.n785 VDAC_N.n784 0.180667
R14660 VDAC_N.n786 VDAC_N.n785 0.180667
R14661 VDAC_N.n787 VDAC_N.n786 0.180667
R14662 VDAC_N.n788 VDAC_N.n787 0.180667
R14663 VDAC_N.n789 VDAC_N.n788 0.180667
R14664 VDAC_N.n790 VDAC_N.n789 0.180667
R14665 VDAC_N.n791 VDAC_N.n790 0.180667
R14666 VDAC_N.n792 VDAC_N.n791 0.180667
R14667 VDAC_N.n793 VDAC_N.n792 0.180667
R14668 VDAC_N.n794 VDAC_N.n793 0.180667
R14669 VDAC_N.n795 VDAC_N.n794 0.180667
R14670 VDAC_N.n796 VDAC_N.n795 0.180667
R14671 VDAC_N.n797 VDAC_N.n796 0.180667
R14672 VDAC_N.n798 VDAC_N.n797 0.180667
R14673 VDAC_N.n799 VDAC_N.n798 0.180667
R14674 VDAC_N.n800 VDAC_N.n799 0.180667
R14675 VDAC_N.n801 VDAC_N.n800 0.180667
R14676 VDAC_N.n802 VDAC_N.n801 0.180667
R14677 VDAC_N.n803 VDAC_N.n802 0.180667
R14678 VDAC_N.n804 VDAC_N.n803 0.180667
R14679 VDAC_N.n805 VDAC_N.n804 0.180667
R14680 VDAC_N.n806 VDAC_N.n805 0.180667
R14681 VDAC_N.n807 VDAC_N.n806 0.180667
R14682 VDAC_N.n808 VDAC_N.n807 0.180667
R14683 VDAC_N.n809 VDAC_N.n808 0.180667
R14684 VDAC_N.n810 VDAC_N.n105 0.180667
R14685 VDAC_N.n811 VDAC_N.n810 0.180667
R14686 VDAC_N.n812 VDAC_N.n811 0.180667
R14687 VDAC_N.n813 VDAC_N.n812 0.180667
R14688 VDAC_N.n814 VDAC_N.n813 0.180667
R14689 VDAC_N.n815 VDAC_N.n814 0.180667
R14690 VDAC_N.n816 VDAC_N.n815 0.180667
R14691 VDAC_N.n817 VDAC_N.n816 0.180667
R14692 VDAC_N.n818 VDAC_N.n817 0.180667
R14693 VDAC_N.n819 VDAC_N.n818 0.180667
R14694 VDAC_N.n820 VDAC_N.n819 0.180667
R14695 VDAC_N.n821 VDAC_N.n820 0.180667
R14696 VDAC_N.n822 VDAC_N.n821 0.180667
R14697 VDAC_N.n823 VDAC_N.n822 0.180667
R14698 VDAC_N.n824 VDAC_N.n823 0.180667
R14699 VDAC_N.n825 VDAC_N.n824 0.180667
R14700 VDAC_N.n826 VDAC_N.n825 0.180667
R14701 VDAC_N.n827 VDAC_N.n826 0.180667
R14702 VDAC_N.n828 VDAC_N.n827 0.180667
R14703 VDAC_N.n829 VDAC_N.n828 0.180667
R14704 VDAC_N.n830 VDAC_N.n829 0.180667
R14705 VDAC_N.n831 VDAC_N.n830 0.180667
R14706 VDAC_N.n832 VDAC_N.n831 0.180667
R14707 VDAC_N.n833 VDAC_N.n832 0.180667
R14708 VDAC_N.n834 VDAC_N.n833 0.180667
R14709 VDAC_N.n835 VDAC_N.n834 0.180667
R14710 VDAC_N.n836 VDAC_N.n835 0.180667
R14711 VDAC_N.n837 VDAC_N.n836 0.180667
R14712 VDAC_N.n838 VDAC_N.n837 0.180667
R14713 VDAC_N.n839 VDAC_N.n838 0.180667
R14714 VDAC_N.n840 VDAC_N.n839 0.180667
R14715 VDAC_N.n841 VDAC_N.n840 0.180667
R14716 VDAC_N.n842 VDAC_N.n841 0.180667
R14717 VDAC_N.n843 VDAC_N.n842 0.180667
R14718 VDAC_N.n844 VDAC_N.n843 0.180667
R14719 VDAC_N.n845 VDAC_N.n844 0.180667
R14720 VDAC_N.n846 VDAC_N.n845 0.180667
R14721 VDAC_N.n847 VDAC_N.n846 0.180667
R14722 VDAC_N.n848 VDAC_N.n847 0.180667
R14723 VDAC_N.n849 VDAC_N.n848 0.180667
R14724 VDAC_N.n850 VDAC_N.n849 0.180667
R14725 VDAC_N.n851 VDAC_N.n850 0.180667
R14726 VDAC_N.n852 VDAC_N.n851 0.180667
R14727 VDAC_N.n853 VDAC_N.n852 0.180667
R14728 VDAC_N.n854 VDAC_N.n853 0.180667
R14729 VDAC_N.n855 VDAC_N.n854 0.180667
R14730 VDAC_N.n856 VDAC_N.n855 0.180667
R14731 VDAC_N.n857 VDAC_N.n856 0.180667
R14732 VDAC_N.n858 VDAC_N.n857 0.180667
R14733 VDAC_N.n859 VDAC_N.n858 0.180667
R14734 VDAC_N.n860 VDAC_N.n859 0.180667
R14735 VDAC_N.n861 VDAC_N.n860 0.180667
R14736 VDAC_N.n862 VDAC_N.n861 0.180667
R14737 VDAC_N.n863 VDAC_N.n862 0.180667
R14738 VDAC_N.n864 VDAC_N.n863 0.180667
R14739 VDAC_N.n865 VDAC_N.n864 0.180667
R14740 VDAC_N.n866 VDAC_N.n865 0.180667
R14741 VDAC_N.n867 VDAC_N.n866 0.180667
R14742 VDAC_N.n868 VDAC_N.n867 0.180667
R14743 VDAC_N.n869 VDAC_N.n868 0.180667
R14744 VDAC_N.n870 VDAC_N.n869 0.180667
R14745 VDAC_N.n871 VDAC_N.n870 0.180667
R14746 VDAC_N.n872 VDAC_N.n871 0.180667
R14747 VDAC_N.n873 VDAC_N.n104 0.180667
R14748 VDAC_N.n874 VDAC_N.n873 0.180667
R14749 VDAC_N.n875 VDAC_N.n874 0.180667
R14750 VDAC_N.n876 VDAC_N.n875 0.180667
R14751 VDAC_N.n877 VDAC_N.n876 0.180667
R14752 VDAC_N.n878 VDAC_N.n877 0.180667
R14753 VDAC_N.n879 VDAC_N.n878 0.180667
R14754 VDAC_N.n880 VDAC_N.n879 0.180667
R14755 VDAC_N.n881 VDAC_N.n880 0.180667
R14756 VDAC_N.n882 VDAC_N.n881 0.180667
R14757 VDAC_N.n883 VDAC_N.n882 0.180667
R14758 VDAC_N.n884 VDAC_N.n883 0.180667
R14759 VDAC_N.n885 VDAC_N.n884 0.180667
R14760 VDAC_N.n886 VDAC_N.n885 0.180667
R14761 VDAC_N.n887 VDAC_N.n886 0.180667
R14762 VDAC_N.n888 VDAC_N.n887 0.180667
R14763 VDAC_N.n889 VDAC_N.n888 0.180667
R14764 VDAC_N.n890 VDAC_N.n889 0.180667
R14765 VDAC_N.n891 VDAC_N.n890 0.180667
R14766 VDAC_N.n892 VDAC_N.n891 0.180667
R14767 VDAC_N.n893 VDAC_N.n892 0.180667
R14768 VDAC_N.n894 VDAC_N.n893 0.180667
R14769 VDAC_N.n895 VDAC_N.n894 0.180667
R14770 VDAC_N.n896 VDAC_N.n895 0.180667
R14771 VDAC_N.n897 VDAC_N.n896 0.180667
R14772 VDAC_N.n898 VDAC_N.n897 0.180667
R14773 VDAC_N.n899 VDAC_N.n898 0.180667
R14774 VDAC_N.n900 VDAC_N.n899 0.180667
R14775 VDAC_N.n901 VDAC_N.n900 0.180667
R14776 VDAC_N.n902 VDAC_N.n901 0.180667
R14777 VDAC_N.n903 VDAC_N.n902 0.180667
R14778 VDAC_N.n904 VDAC_N.n903 0.180667
R14779 VDAC_N.n905 VDAC_N.n904 0.180667
R14780 VDAC_N.n906 VDAC_N.n905 0.180667
R14781 VDAC_N.n907 VDAC_N.n906 0.180667
R14782 VDAC_N.n908 VDAC_N.n907 0.180667
R14783 VDAC_N.n909 VDAC_N.n908 0.180667
R14784 VDAC_N.n910 VDAC_N.n909 0.180667
R14785 VDAC_N.n911 VDAC_N.n910 0.180667
R14786 VDAC_N.n912 VDAC_N.n911 0.180667
R14787 VDAC_N.n913 VDAC_N.n912 0.180667
R14788 VDAC_N.n914 VDAC_N.n913 0.180667
R14789 VDAC_N.n915 VDAC_N.n914 0.180667
R14790 VDAC_N.n916 VDAC_N.n915 0.180667
R14791 VDAC_N.n917 VDAC_N.n916 0.180667
R14792 VDAC_N.n918 VDAC_N.n917 0.180667
R14793 VDAC_N.n919 VDAC_N.n918 0.180667
R14794 VDAC_N.n920 VDAC_N.n919 0.180667
R14795 VDAC_N.n921 VDAC_N.n920 0.180667
R14796 VDAC_N.n922 VDAC_N.n921 0.180667
R14797 VDAC_N.n923 VDAC_N.n922 0.180667
R14798 VDAC_N.n924 VDAC_N.n923 0.180667
R14799 VDAC_N.n925 VDAC_N.n924 0.180667
R14800 VDAC_N.n926 VDAC_N.n925 0.180667
R14801 VDAC_N.n927 VDAC_N.n926 0.180667
R14802 VDAC_N.n928 VDAC_N.n927 0.180667
R14803 VDAC_N.n929 VDAC_N.n928 0.180667
R14804 VDAC_N.n930 VDAC_N.n929 0.180667
R14805 VDAC_N.n931 VDAC_N.n930 0.180667
R14806 VDAC_N.n932 VDAC_N.n931 0.180667
R14807 VDAC_N.n933 VDAC_N.n932 0.180667
R14808 VDAC_N.n934 VDAC_N.n933 0.180667
R14809 VDAC_N.n935 VDAC_N.n934 0.180667
R14810 VDAC_N.n936 VDAC_N.n103 0.180667
R14811 VDAC_N.n937 VDAC_N.n936 0.180667
R14812 VDAC_N.n938 VDAC_N.n937 0.180667
R14813 VDAC_N.n939 VDAC_N.n938 0.180667
R14814 VDAC_N.n940 VDAC_N.n939 0.180667
R14815 VDAC_N.n941 VDAC_N.n940 0.180667
R14816 VDAC_N.n942 VDAC_N.n941 0.180667
R14817 VDAC_N.n943 VDAC_N.n942 0.180667
R14818 VDAC_N.n944 VDAC_N.n943 0.180667
R14819 VDAC_N.n945 VDAC_N.n944 0.180667
R14820 VDAC_N.n946 VDAC_N.n945 0.180667
R14821 VDAC_N.n947 VDAC_N.n946 0.180667
R14822 VDAC_N.n948 VDAC_N.n947 0.180667
R14823 VDAC_N.n949 VDAC_N.n948 0.180667
R14824 VDAC_N.n950 VDAC_N.n949 0.180667
R14825 VDAC_N.n951 VDAC_N.n950 0.180667
R14826 VDAC_N.n952 VDAC_N.n951 0.180667
R14827 VDAC_N.n953 VDAC_N.n952 0.180667
R14828 VDAC_N.n954 VDAC_N.n953 0.180667
R14829 VDAC_N.n955 VDAC_N.n954 0.180667
R14830 VDAC_N.n956 VDAC_N.n955 0.180667
R14831 VDAC_N.n957 VDAC_N.n956 0.180667
R14832 VDAC_N.n958 VDAC_N.n957 0.180667
R14833 VDAC_N.n959 VDAC_N.n958 0.180667
R14834 VDAC_N.n960 VDAC_N.n959 0.180667
R14835 VDAC_N.n961 VDAC_N.n960 0.180667
R14836 VDAC_N.n962 VDAC_N.n961 0.180667
R14837 VDAC_N.n963 VDAC_N.n962 0.180667
R14838 VDAC_N.n964 VDAC_N.n963 0.180667
R14839 VDAC_N.n965 VDAC_N.n964 0.180667
R14840 VDAC_N.n966 VDAC_N.n965 0.180667
R14841 VDAC_N.n967 VDAC_N.n966 0.180667
R14842 VDAC_N.n968 VDAC_N.n967 0.180667
R14843 VDAC_N.n969 VDAC_N.n968 0.180667
R14844 VDAC_N.n970 VDAC_N.n969 0.180667
R14845 VDAC_N.n971 VDAC_N.n970 0.180667
R14846 VDAC_N.n972 VDAC_N.n971 0.180667
R14847 VDAC_N.n973 VDAC_N.n972 0.180667
R14848 VDAC_N.n974 VDAC_N.n973 0.180667
R14849 VDAC_N.n975 VDAC_N.n974 0.180667
R14850 VDAC_N.n976 VDAC_N.n975 0.180667
R14851 VDAC_N.n977 VDAC_N.n976 0.180667
R14852 VDAC_N.n978 VDAC_N.n977 0.180667
R14853 VDAC_N.n979 VDAC_N.n978 0.180667
R14854 VDAC_N.n980 VDAC_N.n979 0.180667
R14855 VDAC_N.n981 VDAC_N.n980 0.180667
R14856 VDAC_N.n982 VDAC_N.n981 0.180667
R14857 VDAC_N.n983 VDAC_N.n982 0.180667
R14858 VDAC_N.n984 VDAC_N.n983 0.180667
R14859 VDAC_N.n985 VDAC_N.n984 0.180667
R14860 VDAC_N.n986 VDAC_N.n985 0.180667
R14861 VDAC_N.n987 VDAC_N.n986 0.180667
R14862 VDAC_N.n988 VDAC_N.n987 0.180667
R14863 VDAC_N.n989 VDAC_N.n988 0.180667
R14864 VDAC_N.n990 VDAC_N.n989 0.180667
R14865 VDAC_N.n991 VDAC_N.n990 0.180667
R14866 VDAC_N.n992 VDAC_N.n991 0.180667
R14867 VDAC_N.n993 VDAC_N.n992 0.180667
R14868 VDAC_N.n994 VDAC_N.n993 0.180667
R14869 VDAC_N.n995 VDAC_N.n994 0.180667
R14870 VDAC_N.n996 VDAC_N.n995 0.180667
R14871 VDAC_N.n997 VDAC_N.n996 0.180667
R14872 VDAC_N.n998 VDAC_N.n997 0.180667
R14873 VDAC_N.n999 VDAC_N.n102 0.180667
R14874 VDAC_N.n1000 VDAC_N.n999 0.180667
R14875 VDAC_N.n1001 VDAC_N.n1000 0.180667
R14876 VDAC_N.n1002 VDAC_N.n1001 0.180667
R14877 VDAC_N.n1003 VDAC_N.n1002 0.180667
R14878 VDAC_N.n1004 VDAC_N.n1003 0.180667
R14879 VDAC_N.n1005 VDAC_N.n1004 0.180667
R14880 VDAC_N.n1006 VDAC_N.n1005 0.180667
R14881 VDAC_N.n1007 VDAC_N.n1006 0.180667
R14882 VDAC_N.n1008 VDAC_N.n1007 0.180667
R14883 VDAC_N.n1009 VDAC_N.n1008 0.180667
R14884 VDAC_N.n1010 VDAC_N.n1009 0.180667
R14885 VDAC_N.n1011 VDAC_N.n1010 0.180667
R14886 VDAC_N.n1012 VDAC_N.n1011 0.180667
R14887 VDAC_N.n1013 VDAC_N.n1012 0.180667
R14888 VDAC_N.n1014 VDAC_N.n1013 0.180667
R14889 VDAC_N.n1015 VDAC_N.n1014 0.180667
R14890 VDAC_N.n1016 VDAC_N.n1015 0.180667
R14891 VDAC_N.n1017 VDAC_N.n1016 0.180667
R14892 VDAC_N.n1018 VDAC_N.n1017 0.180667
R14893 VDAC_N.n1019 VDAC_N.n1018 0.180667
R14894 VDAC_N.n1020 VDAC_N.n1019 0.180667
R14895 VDAC_N.n1021 VDAC_N.n1020 0.180667
R14896 VDAC_N.n1022 VDAC_N.n1021 0.180667
R14897 VDAC_N.n1023 VDAC_N.n1022 0.180667
R14898 VDAC_N.n1024 VDAC_N.n1023 0.180667
R14899 VDAC_N.n1025 VDAC_N.n1024 0.180667
R14900 VDAC_N.n1026 VDAC_N.n1025 0.180667
R14901 VDAC_N.n1027 VDAC_N.n1026 0.180667
R14902 VDAC_N.n1028 VDAC_N.n1027 0.180667
R14903 VDAC_N.n1029 VDAC_N.n1028 0.180667
R14904 VDAC_N.n1030 VDAC_N.n1029 0.180667
R14905 VDAC_N.n1031 VDAC_N.n1030 0.180667
R14906 VDAC_N.n1032 VDAC_N.n1031 0.180667
R14907 VDAC_N.n1033 VDAC_N.n1032 0.180667
R14908 VDAC_N.n1034 VDAC_N.n1033 0.180667
R14909 VDAC_N.n1035 VDAC_N.n1034 0.180667
R14910 VDAC_N.n1036 VDAC_N.n1035 0.180667
R14911 VDAC_N.n1037 VDAC_N.n1036 0.180667
R14912 VDAC_N.n1038 VDAC_N.n1037 0.180667
R14913 VDAC_N.n1039 VDAC_N.n1038 0.180667
R14914 VDAC_N.n1040 VDAC_N.n1039 0.180667
R14915 VDAC_N.n1041 VDAC_N.n1040 0.180667
R14916 VDAC_N.n1042 VDAC_N.n1041 0.180667
R14917 VDAC_N.n1043 VDAC_N.n1042 0.180667
R14918 VDAC_N.n1044 VDAC_N.n1043 0.180667
R14919 VDAC_N.n1045 VDAC_N.n1044 0.180667
R14920 VDAC_N.n1046 VDAC_N.n1045 0.180667
R14921 VDAC_N.n1047 VDAC_N.n1046 0.180667
R14922 VDAC_N.n1048 VDAC_N.n1047 0.180667
R14923 VDAC_N.n1049 VDAC_N.n1048 0.180667
R14924 VDAC_N.n1050 VDAC_N.n1049 0.180667
R14925 VDAC_N.n1051 VDAC_N.n1050 0.180667
R14926 VDAC_N.n1052 VDAC_N.n1051 0.180667
R14927 VDAC_N.n1053 VDAC_N.n1052 0.180667
R14928 VDAC_N.n1054 VDAC_N.n1053 0.180667
R14929 VDAC_N.n1055 VDAC_N.n1054 0.180667
R14930 VDAC_N.n1056 VDAC_N.n1055 0.180667
R14931 VDAC_N.n1057 VDAC_N.n1056 0.180667
R14932 VDAC_N.n1058 VDAC_N.n1057 0.180667
R14933 VDAC_N.n1059 VDAC_N.n1058 0.180667
R14934 VDAC_N.n1060 VDAC_N.n1059 0.180667
R14935 VDAC_N.n1061 VDAC_N.n1060 0.180667
R14936 VDAC_N.n1062 VDAC_N.n101 0.180667
R14937 VDAC_N.n1063 VDAC_N.n1062 0.180667
R14938 VDAC_N.n1064 VDAC_N.n1063 0.180667
R14939 VDAC_N.n1065 VDAC_N.n1064 0.180667
R14940 VDAC_N.n1066 VDAC_N.n1065 0.180667
R14941 VDAC_N.n1067 VDAC_N.n1066 0.180667
R14942 VDAC_N.n1068 VDAC_N.n1067 0.180667
R14943 VDAC_N.n1069 VDAC_N.n1068 0.180667
R14944 VDAC_N.n1070 VDAC_N.n1069 0.180667
R14945 VDAC_N.n1071 VDAC_N.n1070 0.180667
R14946 VDAC_N.n1072 VDAC_N.n1071 0.180667
R14947 VDAC_N.n1073 VDAC_N.n1072 0.180667
R14948 VDAC_N.n1074 VDAC_N.n1073 0.180667
R14949 VDAC_N.n1075 VDAC_N.n1074 0.180667
R14950 VDAC_N.n1076 VDAC_N.n1075 0.180667
R14951 VDAC_N.n1077 VDAC_N.n1076 0.180667
R14952 VDAC_N.n1078 VDAC_N.n1077 0.180667
R14953 VDAC_N.n1079 VDAC_N.n1078 0.180667
R14954 VDAC_N.n1080 VDAC_N.n1079 0.180667
R14955 VDAC_N.n1081 VDAC_N.n1080 0.180667
R14956 VDAC_N.n1082 VDAC_N.n1081 0.180667
R14957 VDAC_N.n1083 VDAC_N.n1082 0.180667
R14958 VDAC_N.n1084 VDAC_N.n1083 0.180667
R14959 VDAC_N.n1085 VDAC_N.n1084 0.180667
R14960 VDAC_N.n1086 VDAC_N.n1085 0.180667
R14961 VDAC_N.n1087 VDAC_N.n1086 0.180667
R14962 VDAC_N.n1088 VDAC_N.n1087 0.180667
R14963 VDAC_N.n1089 VDAC_N.n1088 0.180667
R14964 VDAC_N.n1090 VDAC_N.n1089 0.180667
R14965 VDAC_N.n1091 VDAC_N.n1090 0.180667
R14966 VDAC_N.n1092 VDAC_N.n1091 0.180667
R14967 VDAC_N.n1093 VDAC_N.n1092 0.180667
R14968 VDAC_N.n1094 VDAC_N.n1093 0.180667
R14969 VDAC_N.n1095 VDAC_N.n1094 0.180667
R14970 VDAC_N.n1096 VDAC_N.n1095 0.180667
R14971 VDAC_N.n1097 VDAC_N.n1096 0.180667
R14972 VDAC_N.n1098 VDAC_N.n1097 0.180667
R14973 VDAC_N.n1099 VDAC_N.n1098 0.180667
R14974 VDAC_N.n1100 VDAC_N.n1099 0.180667
R14975 VDAC_N.n1101 VDAC_N.n1100 0.180667
R14976 VDAC_N.n1102 VDAC_N.n1101 0.180667
R14977 VDAC_N.n1103 VDAC_N.n1102 0.180667
R14978 VDAC_N.n1104 VDAC_N.n1103 0.180667
R14979 VDAC_N.n1105 VDAC_N.n1104 0.180667
R14980 VDAC_N.n1106 VDAC_N.n1105 0.180667
R14981 VDAC_N.n1107 VDAC_N.n1106 0.180667
R14982 VDAC_N.n1108 VDAC_N.n1107 0.180667
R14983 VDAC_N.n1109 VDAC_N.n1108 0.180667
R14984 VDAC_N.n1110 VDAC_N.n1109 0.180667
R14985 VDAC_N.n1111 VDAC_N.n1110 0.180667
R14986 VDAC_N.n1112 VDAC_N.n1111 0.180667
R14987 VDAC_N.n1113 VDAC_N.n1112 0.180667
R14988 VDAC_N.n1114 VDAC_N.n1113 0.180667
R14989 VDAC_N.n1115 VDAC_N.n1114 0.180667
R14990 VDAC_N.n1116 VDAC_N.n1115 0.180667
R14991 VDAC_N.n1117 VDAC_N.n1116 0.180667
R14992 VDAC_N.n1118 VDAC_N.n1117 0.180667
R14993 VDAC_N.n1119 VDAC_N.n1118 0.180667
R14994 VDAC_N.n1120 VDAC_N.n1119 0.180667
R14995 VDAC_N.n1121 VDAC_N.n1120 0.180667
R14996 VDAC_N.n1122 VDAC_N.n1121 0.180667
R14997 VDAC_N.n1123 VDAC_N.n1122 0.180667
R14998 VDAC_N.n1124 VDAC_N.n1123 0.180667
R14999 VDAC_N.n1125 VDAC_N.n100 0.180667
R15000 VDAC_N.n1126 VDAC_N.n1125 0.180667
R15001 VDAC_N.n1127 VDAC_N.n1126 0.180667
R15002 VDAC_N.n1128 VDAC_N.n1127 0.180667
R15003 VDAC_N.n1129 VDAC_N.n1128 0.180667
R15004 VDAC_N.n1130 VDAC_N.n1129 0.180667
R15005 VDAC_N.n1131 VDAC_N.n1130 0.180667
R15006 VDAC_N.n1132 VDAC_N.n1131 0.180667
R15007 VDAC_N.n1133 VDAC_N.n1132 0.180667
R15008 VDAC_N.n1134 VDAC_N.n1133 0.180667
R15009 VDAC_N.n1135 VDAC_N.n1134 0.180667
R15010 VDAC_N.n1136 VDAC_N.n1135 0.180667
R15011 VDAC_N.n1137 VDAC_N.n1136 0.180667
R15012 VDAC_N.n1138 VDAC_N.n1137 0.180667
R15013 VDAC_N.n1139 VDAC_N.n1138 0.180667
R15014 VDAC_N.n1140 VDAC_N.n1139 0.180667
R15015 VDAC_N.n1141 VDAC_N.n1140 0.180667
R15016 VDAC_N.n1142 VDAC_N.n1141 0.180667
R15017 VDAC_N.n1143 VDAC_N.n1142 0.180667
R15018 VDAC_N.n1144 VDAC_N.n1143 0.180667
R15019 VDAC_N.n1145 VDAC_N.n1144 0.180667
R15020 VDAC_N.n1146 VDAC_N.n1145 0.180667
R15021 VDAC_N.n1147 VDAC_N.n1146 0.180667
R15022 VDAC_N.n1148 VDAC_N.n1147 0.180667
R15023 VDAC_N.n1149 VDAC_N.n1148 0.180667
R15024 VDAC_N.n1150 VDAC_N.n1149 0.180667
R15025 VDAC_N.n1151 VDAC_N.n1150 0.180667
R15026 VDAC_N.n1152 VDAC_N.n1151 0.180667
R15027 VDAC_N.n1153 VDAC_N.n1152 0.180667
R15028 VDAC_N.n1154 VDAC_N.n1153 0.180667
R15029 VDAC_N.n1155 VDAC_N.n1154 0.180667
R15030 VDAC_N.n1156 VDAC_N.n1155 0.180667
R15031 VDAC_N.n1157 VDAC_N.n1156 0.180667
R15032 VDAC_N.n1158 VDAC_N.n1157 0.180667
R15033 VDAC_N.n1159 VDAC_N.n1158 0.180667
R15034 VDAC_N.n1160 VDAC_N.n1159 0.180667
R15035 VDAC_N.n1161 VDAC_N.n1160 0.180667
R15036 VDAC_N.n1162 VDAC_N.n1161 0.180667
R15037 VDAC_N.n1163 VDAC_N.n1162 0.180667
R15038 VDAC_N.n1164 VDAC_N.n1163 0.180667
R15039 VDAC_N.n1165 VDAC_N.n1164 0.180667
R15040 VDAC_N.n1166 VDAC_N.n1165 0.180667
R15041 VDAC_N.n1167 VDAC_N.n1166 0.180667
R15042 VDAC_N.n1168 VDAC_N.n1167 0.180667
R15043 VDAC_N.n1169 VDAC_N.n1168 0.180667
R15044 VDAC_N.n1170 VDAC_N.n1169 0.180667
R15045 VDAC_N.n1171 VDAC_N.n1170 0.180667
R15046 VDAC_N.n1172 VDAC_N.n1171 0.180667
R15047 VDAC_N.n1173 VDAC_N.n1172 0.180667
R15048 VDAC_N.n1174 VDAC_N.n1173 0.180667
R15049 VDAC_N.n1175 VDAC_N.n1174 0.180667
R15050 VDAC_N.n1176 VDAC_N.n1175 0.180667
R15051 VDAC_N.n1177 VDAC_N.n1176 0.180667
R15052 VDAC_N.n1178 VDAC_N.n1177 0.180667
R15053 VDAC_N.n1179 VDAC_N.n1178 0.180667
R15054 VDAC_N.n1180 VDAC_N.n1179 0.180667
R15055 VDAC_N.n1181 VDAC_N.n1180 0.180667
R15056 VDAC_N.n1182 VDAC_N.n1181 0.180667
R15057 VDAC_N.n1183 VDAC_N.n1182 0.180667
R15058 VDAC_N.n1184 VDAC_N.n1183 0.180667
R15059 VDAC_N.n1185 VDAC_N.n1184 0.180667
R15060 VDAC_N.n1186 VDAC_N.n1185 0.180667
R15061 VDAC_N.n1187 VDAC_N.n1186 0.180667
R15062 VDAC_N.n1188 VDAC_N.n99 0.180667
R15063 VDAC_N.n1189 VDAC_N.n1188 0.180667
R15064 VDAC_N.n1190 VDAC_N.n1189 0.180667
R15065 VDAC_N.n1191 VDAC_N.n1190 0.180667
R15066 VDAC_N.n1192 VDAC_N.n1191 0.180667
R15067 VDAC_N.n1193 VDAC_N.n1192 0.180667
R15068 VDAC_N.n1194 VDAC_N.n1193 0.180667
R15069 VDAC_N.n1195 VDAC_N.n1194 0.180667
R15070 VDAC_N.n1196 VDAC_N.n1195 0.180667
R15071 VDAC_N.n1197 VDAC_N.n1196 0.180667
R15072 VDAC_N.n1198 VDAC_N.n1197 0.180667
R15073 VDAC_N.n1199 VDAC_N.n1198 0.180667
R15074 VDAC_N.n1200 VDAC_N.n1199 0.180667
R15075 VDAC_N.n1201 VDAC_N.n1200 0.180667
R15076 VDAC_N.n1202 VDAC_N.n1201 0.180667
R15077 VDAC_N.n1203 VDAC_N.n1202 0.180667
R15078 VDAC_N.n1204 VDAC_N.n1203 0.180667
R15079 VDAC_N.n1205 VDAC_N.n1204 0.180667
R15080 VDAC_N.n1206 VDAC_N.n1205 0.180667
R15081 VDAC_N.n1207 VDAC_N.n1206 0.180667
R15082 VDAC_N.n1208 VDAC_N.n1207 0.180667
R15083 VDAC_N.n1209 VDAC_N.n1208 0.180667
R15084 VDAC_N.n1210 VDAC_N.n1209 0.180667
R15085 VDAC_N.n1211 VDAC_N.n1210 0.180667
R15086 VDAC_N.n1212 VDAC_N.n1211 0.180667
R15087 VDAC_N.n1213 VDAC_N.n1212 0.180667
R15088 VDAC_N.n1214 VDAC_N.n1213 0.180667
R15089 VDAC_N.n1215 VDAC_N.n1214 0.180667
R15090 VDAC_N.n1216 VDAC_N.n1215 0.180667
R15091 VDAC_N.n1217 VDAC_N.n1216 0.180667
R15092 VDAC_N.n1218 VDAC_N.n1217 0.180667
R15093 VDAC_N.n1219 VDAC_N.n1218 0.180667
R15094 VDAC_N.n1220 VDAC_N.n1219 0.180667
R15095 VDAC_N.n1221 VDAC_N.n1220 0.180667
R15096 VDAC_N.n1222 VDAC_N.n1221 0.180667
R15097 VDAC_N.n1223 VDAC_N.n1222 0.180667
R15098 VDAC_N.n1224 VDAC_N.n1223 0.180667
R15099 VDAC_N.n1225 VDAC_N.n1224 0.180667
R15100 VDAC_N.n1226 VDAC_N.n1225 0.180667
R15101 VDAC_N.n1227 VDAC_N.n1226 0.180667
R15102 VDAC_N.n1228 VDAC_N.n1227 0.180667
R15103 VDAC_N.n1229 VDAC_N.n1228 0.180667
R15104 VDAC_N.n1230 VDAC_N.n1229 0.180667
R15105 VDAC_N.n1231 VDAC_N.n1230 0.180667
R15106 VDAC_N.n1232 VDAC_N.n1231 0.180667
R15107 VDAC_N.n1233 VDAC_N.n1232 0.180667
R15108 VDAC_N.n1234 VDAC_N.n1233 0.180667
R15109 VDAC_N.n1235 VDAC_N.n1234 0.180667
R15110 VDAC_N.n1236 VDAC_N.n1235 0.180667
R15111 VDAC_N.n1237 VDAC_N.n1236 0.180667
R15112 VDAC_N.n1238 VDAC_N.n1237 0.180667
R15113 VDAC_N.n1239 VDAC_N.n1238 0.180667
R15114 VDAC_N.n1240 VDAC_N.n1239 0.180667
R15115 VDAC_N.n1241 VDAC_N.n1240 0.180667
R15116 VDAC_N.n1242 VDAC_N.n1241 0.180667
R15117 VDAC_N.n1243 VDAC_N.n1242 0.180667
R15118 VDAC_N.n1244 VDAC_N.n1243 0.180667
R15119 VDAC_N.n1245 VDAC_N.n1244 0.180667
R15120 VDAC_N.n1246 VDAC_N.n1245 0.180667
R15121 VDAC_N.n1247 VDAC_N.n1246 0.180667
R15122 VDAC_N.n1248 VDAC_N.n1247 0.180667
R15123 VDAC_N.n1249 VDAC_N.n1248 0.180667
R15124 VDAC_N.n1250 VDAC_N.n1249 0.180667
R15125 VDAC_N.n1251 VDAC_N.n98 0.180667
R15126 VDAC_N.n1252 VDAC_N.n1251 0.180667
R15127 VDAC_N.n1253 VDAC_N.n1252 0.180667
R15128 VDAC_N.n1254 VDAC_N.n1253 0.180667
R15129 VDAC_N.n1255 VDAC_N.n1254 0.180667
R15130 VDAC_N.n1256 VDAC_N.n1255 0.180667
R15131 VDAC_N.n1257 VDAC_N.n1256 0.180667
R15132 VDAC_N.n1258 VDAC_N.n1257 0.180667
R15133 VDAC_N.n1259 VDAC_N.n1258 0.180667
R15134 VDAC_N.n1260 VDAC_N.n1259 0.180667
R15135 VDAC_N.n1261 VDAC_N.n1260 0.180667
R15136 VDAC_N.n1262 VDAC_N.n1261 0.180667
R15137 VDAC_N.n1263 VDAC_N.n1262 0.180667
R15138 VDAC_N.n1264 VDAC_N.n1263 0.180667
R15139 VDAC_N.n1265 VDAC_N.n1264 0.180667
R15140 VDAC_N.n1266 VDAC_N.n1265 0.180667
R15141 VDAC_N.n1267 VDAC_N.n1266 0.180667
R15142 VDAC_N.n1268 VDAC_N.n1267 0.180667
R15143 VDAC_N.n1269 VDAC_N.n1268 0.180667
R15144 VDAC_N.n1270 VDAC_N.n1269 0.180667
R15145 VDAC_N.n1271 VDAC_N.n1270 0.180667
R15146 VDAC_N.n1272 VDAC_N.n1271 0.180667
R15147 VDAC_N.n1273 VDAC_N.n1272 0.180667
R15148 VDAC_N.n1274 VDAC_N.n1273 0.180667
R15149 VDAC_N.n1275 VDAC_N.n1274 0.180667
R15150 VDAC_N.n1276 VDAC_N.n1275 0.180667
R15151 VDAC_N.n1277 VDAC_N.n1276 0.180667
R15152 VDAC_N.n1278 VDAC_N.n1277 0.180667
R15153 VDAC_N.n1279 VDAC_N.n1278 0.180667
R15154 VDAC_N.n1280 VDAC_N.n1279 0.180667
R15155 VDAC_N.n1281 VDAC_N.n1280 0.180667
R15156 VDAC_N.n1282 VDAC_N.n1281 0.180667
R15157 VDAC_N.n1283 VDAC_N.n1282 0.180667
R15158 VDAC_N.n1284 VDAC_N.n1283 0.180667
R15159 VDAC_N.n1285 VDAC_N.n1284 0.180667
R15160 VDAC_N.n1286 VDAC_N.n1285 0.180667
R15161 VDAC_N.n1287 VDAC_N.n1286 0.180667
R15162 VDAC_N.n1288 VDAC_N.n1287 0.180667
R15163 VDAC_N.n1289 VDAC_N.n1288 0.180667
R15164 VDAC_N.n1290 VDAC_N.n1289 0.180667
R15165 VDAC_N.n1291 VDAC_N.n1290 0.180667
R15166 VDAC_N.n1292 VDAC_N.n1291 0.180667
R15167 VDAC_N.n1293 VDAC_N.n1292 0.180667
R15168 VDAC_N.n1294 VDAC_N.n1293 0.180667
R15169 VDAC_N.n1295 VDAC_N.n1294 0.180667
R15170 VDAC_N.n1296 VDAC_N.n1295 0.180667
R15171 VDAC_N.n1297 VDAC_N.n1296 0.180667
R15172 VDAC_N.n1298 VDAC_N.n1297 0.180667
R15173 VDAC_N.n1299 VDAC_N.n1298 0.180667
R15174 VDAC_N.n1300 VDAC_N.n1299 0.180667
R15175 VDAC_N.n1301 VDAC_N.n1300 0.180667
R15176 VDAC_N.n1302 VDAC_N.n1301 0.180667
R15177 VDAC_N.n1303 VDAC_N.n1302 0.180667
R15178 VDAC_N.n1304 VDAC_N.n1303 0.180667
R15179 VDAC_N.n1305 VDAC_N.n1304 0.180667
R15180 VDAC_N.n1306 VDAC_N.n1305 0.180667
R15181 VDAC_N.n1307 VDAC_N.n1306 0.180667
R15182 VDAC_N.n1308 VDAC_N.n1307 0.180667
R15183 VDAC_N.n1309 VDAC_N.n1308 0.180667
R15184 VDAC_N.n1310 VDAC_N.n1309 0.180667
R15185 VDAC_N.n1311 VDAC_N.n1310 0.180667
R15186 VDAC_N.n1312 VDAC_N.n1311 0.180667
R15187 VDAC_N.n1313 VDAC_N.n1312 0.180667
R15188 VDAC_N.n1314 VDAC_N.n97 0.180667
R15189 VDAC_N.n1315 VDAC_N.n1314 0.180667
R15190 VDAC_N.n1316 VDAC_N.n1315 0.180667
R15191 VDAC_N.n1317 VDAC_N.n1316 0.180667
R15192 VDAC_N.n1318 VDAC_N.n1317 0.180667
R15193 VDAC_N.n1319 VDAC_N.n1318 0.180667
R15194 VDAC_N.n1320 VDAC_N.n1319 0.180667
R15195 VDAC_N.n1321 VDAC_N.n1320 0.180667
R15196 VDAC_N.n1322 VDAC_N.n1321 0.180667
R15197 VDAC_N.n1323 VDAC_N.n1322 0.180667
R15198 VDAC_N.n1324 VDAC_N.n1323 0.180667
R15199 VDAC_N.n1325 VDAC_N.n1324 0.180667
R15200 VDAC_N.n1326 VDAC_N.n1325 0.180667
R15201 VDAC_N.n1327 VDAC_N.n1326 0.180667
R15202 VDAC_N.n1328 VDAC_N.n1327 0.180667
R15203 VDAC_N.n1329 VDAC_N.n1328 0.180667
R15204 VDAC_N.n1330 VDAC_N.n1329 0.180667
R15205 VDAC_N.n1331 VDAC_N.n1330 0.180667
R15206 VDAC_N.n1332 VDAC_N.n1331 0.180667
R15207 VDAC_N.n1333 VDAC_N.n1332 0.180667
R15208 VDAC_N.n1334 VDAC_N.n1333 0.180667
R15209 VDAC_N.n1335 VDAC_N.n1334 0.180667
R15210 VDAC_N.n1336 VDAC_N.n1335 0.180667
R15211 VDAC_N.n1337 VDAC_N.n1336 0.180667
R15212 VDAC_N.n1338 VDAC_N.n1337 0.180667
R15213 VDAC_N.n1339 VDAC_N.n1338 0.180667
R15214 VDAC_N.n1340 VDAC_N.n1339 0.180667
R15215 VDAC_N.n1341 VDAC_N.n1340 0.180667
R15216 VDAC_N.n1342 VDAC_N.n1341 0.180667
R15217 VDAC_N.n1343 VDAC_N.n1342 0.180667
R15218 VDAC_N.n1344 VDAC_N.n1343 0.180667
R15219 VDAC_N.n1345 VDAC_N.n1344 0.180667
R15220 VDAC_N.n1346 VDAC_N.n1345 0.180667
R15221 VDAC_N.n1347 VDAC_N.n1346 0.180667
R15222 VDAC_N.n1348 VDAC_N.n1347 0.180667
R15223 VDAC_N.n1349 VDAC_N.n1348 0.180667
R15224 VDAC_N.n1350 VDAC_N.n1349 0.180667
R15225 VDAC_N.n1351 VDAC_N.n1350 0.180667
R15226 VDAC_N.n1352 VDAC_N.n1351 0.180667
R15227 VDAC_N.n1353 VDAC_N.n1352 0.180667
R15228 VDAC_N.n1354 VDAC_N.n1353 0.180667
R15229 VDAC_N.n1355 VDAC_N.n1354 0.180667
R15230 VDAC_N.n1356 VDAC_N.n1355 0.180667
R15231 VDAC_N.n1357 VDAC_N.n1356 0.180667
R15232 VDAC_N.n1358 VDAC_N.n1357 0.180667
R15233 VDAC_N.n1359 VDAC_N.n1358 0.180667
R15234 VDAC_N.n1360 VDAC_N.n1359 0.180667
R15235 VDAC_N.n1361 VDAC_N.n1360 0.180667
R15236 VDAC_N.n1362 VDAC_N.n1361 0.180667
R15237 VDAC_N.n1363 VDAC_N.n1362 0.180667
R15238 VDAC_N.n1364 VDAC_N.n1363 0.180667
R15239 VDAC_N.n1365 VDAC_N.n1364 0.180667
R15240 VDAC_N.n1366 VDAC_N.n1365 0.180667
R15241 VDAC_N.n1367 VDAC_N.n1366 0.180667
R15242 VDAC_N.n1368 VDAC_N.n1367 0.180667
R15243 VDAC_N.n1369 VDAC_N.n1368 0.180667
R15244 VDAC_N.n1370 VDAC_N.n1369 0.180667
R15245 VDAC_N.n1371 VDAC_N.n1370 0.180667
R15246 VDAC_N.n1372 VDAC_N.n1371 0.180667
R15247 VDAC_N.n1373 VDAC_N.n1372 0.180667
R15248 VDAC_N.n1374 VDAC_N.n1373 0.180667
R15249 VDAC_N.n1375 VDAC_N.n1374 0.180667
R15250 VDAC_N.n1376 VDAC_N.n1375 0.180667
R15251 VDAC_N.n1377 VDAC_N.n96 0.180667
R15252 VDAC_N.n1378 VDAC_N.n1377 0.180667
R15253 VDAC_N.n1379 VDAC_N.n1378 0.180667
R15254 VDAC_N.n1380 VDAC_N.n1379 0.180667
R15255 VDAC_N.n1381 VDAC_N.n1380 0.180667
R15256 VDAC_N.n1382 VDAC_N.n1381 0.180667
R15257 VDAC_N.n1383 VDAC_N.n1382 0.180667
R15258 VDAC_N.n1384 VDAC_N.n1383 0.180667
R15259 VDAC_N.n1385 VDAC_N.n1384 0.180667
R15260 VDAC_N.n1386 VDAC_N.n1385 0.180667
R15261 VDAC_N.n1387 VDAC_N.n1386 0.180667
R15262 VDAC_N.n1388 VDAC_N.n1387 0.180667
R15263 VDAC_N.n1389 VDAC_N.n1388 0.180667
R15264 VDAC_N.n1390 VDAC_N.n1389 0.180667
R15265 VDAC_N.n1391 VDAC_N.n1390 0.180667
R15266 VDAC_N.n1392 VDAC_N.n1391 0.180667
R15267 VDAC_N.n1393 VDAC_N.n1392 0.180667
R15268 VDAC_N.n1394 VDAC_N.n1393 0.180667
R15269 VDAC_N.n1395 VDAC_N.n1394 0.180667
R15270 VDAC_N.n1396 VDAC_N.n1395 0.180667
R15271 VDAC_N.n1397 VDAC_N.n1396 0.180667
R15272 VDAC_N.n1398 VDAC_N.n1397 0.180667
R15273 VDAC_N.n1399 VDAC_N.n1398 0.180667
R15274 VDAC_N.n1400 VDAC_N.n1399 0.180667
R15275 VDAC_N.n1401 VDAC_N.n1400 0.180667
R15276 VDAC_N.n1402 VDAC_N.n1401 0.180667
R15277 VDAC_N.n1403 VDAC_N.n1402 0.180667
R15278 VDAC_N.n1404 VDAC_N.n1403 0.180667
R15279 VDAC_N.n1405 VDAC_N.n1404 0.180667
R15280 VDAC_N.n1406 VDAC_N.n1405 0.180667
R15281 VDAC_N.n1407 VDAC_N.n1406 0.180667
R15282 VDAC_N.n1408 VDAC_N.n1407 0.180667
R15283 VDAC_N.n1409 VDAC_N.n1408 0.180667
R15284 VDAC_N.n1410 VDAC_N.n1409 0.180667
R15285 VDAC_N.n1411 VDAC_N.n1410 0.180667
R15286 VDAC_N.n1412 VDAC_N.n1411 0.180667
R15287 VDAC_N.n1413 VDAC_N.n1412 0.180667
R15288 VDAC_N.n1414 VDAC_N.n1413 0.180667
R15289 VDAC_N.n1415 VDAC_N.n1414 0.180667
R15290 VDAC_N.n1416 VDAC_N.n1415 0.180667
R15291 VDAC_N.n1417 VDAC_N.n1416 0.180667
R15292 VDAC_N.n1418 VDAC_N.n1417 0.180667
R15293 VDAC_N.n1419 VDAC_N.n1418 0.180667
R15294 VDAC_N.n1420 VDAC_N.n1419 0.180667
R15295 VDAC_N.n1421 VDAC_N.n1420 0.180667
R15296 VDAC_N.n1422 VDAC_N.n1421 0.180667
R15297 VDAC_N.n1423 VDAC_N.n1422 0.180667
R15298 VDAC_N.n1424 VDAC_N.n1423 0.180667
R15299 VDAC_N.n1425 VDAC_N.n1424 0.180667
R15300 VDAC_N.n1426 VDAC_N.n1425 0.180667
R15301 VDAC_N.n1427 VDAC_N.n1426 0.180667
R15302 VDAC_N.n1428 VDAC_N.n1427 0.180667
R15303 VDAC_N.n1429 VDAC_N.n1428 0.180667
R15304 VDAC_N.n1430 VDAC_N.n1429 0.180667
R15305 VDAC_N.n1431 VDAC_N.n1430 0.180667
R15306 VDAC_N.n1432 VDAC_N.n1431 0.180667
R15307 VDAC_N.n1433 VDAC_N.n1432 0.180667
R15308 VDAC_N.n1434 VDAC_N.n1433 0.180667
R15309 VDAC_N.n1435 VDAC_N.n1434 0.180667
R15310 VDAC_N.n1436 VDAC_N.n1435 0.180667
R15311 VDAC_N.n1437 VDAC_N.n1436 0.180667
R15312 VDAC_N.n1438 VDAC_N.n1437 0.180667
R15313 VDAC_N.n1439 VDAC_N.n1438 0.180667
R15314 VDAC_N.n1440 VDAC_N.n95 0.180667
R15315 VDAC_N.n1441 VDAC_N.n1440 0.180667
R15316 VDAC_N.n1442 VDAC_N.n1441 0.180667
R15317 VDAC_N.n1443 VDAC_N.n1442 0.180667
R15318 VDAC_N.n1444 VDAC_N.n1443 0.180667
R15319 VDAC_N.n1445 VDAC_N.n1444 0.180667
R15320 VDAC_N.n1446 VDAC_N.n1445 0.180667
R15321 VDAC_N.n1447 VDAC_N.n1446 0.180667
R15322 VDAC_N.n1448 VDAC_N.n1447 0.180667
R15323 VDAC_N.n1449 VDAC_N.n1448 0.180667
R15324 VDAC_N.n1450 VDAC_N.n1449 0.180667
R15325 VDAC_N.n1451 VDAC_N.n1450 0.180667
R15326 VDAC_N.n1452 VDAC_N.n1451 0.180667
R15327 VDAC_N.n1453 VDAC_N.n1452 0.180667
R15328 VDAC_N.n1454 VDAC_N.n1453 0.180667
R15329 VDAC_N.n1455 VDAC_N.n1454 0.180667
R15330 VDAC_N.n1456 VDAC_N.n1455 0.180667
R15331 VDAC_N.n1457 VDAC_N.n1456 0.180667
R15332 VDAC_N.n1458 VDAC_N.n1457 0.180667
R15333 VDAC_N.n1459 VDAC_N.n1458 0.180667
R15334 VDAC_N.n1460 VDAC_N.n1459 0.180667
R15335 VDAC_N.n1461 VDAC_N.n1460 0.180667
R15336 VDAC_N.n1462 VDAC_N.n1461 0.180667
R15337 VDAC_N.n1463 VDAC_N.n1462 0.180667
R15338 VDAC_N.n1464 VDAC_N.n1463 0.180667
R15339 VDAC_N.n1465 VDAC_N.n1464 0.180667
R15340 VDAC_N.n1466 VDAC_N.n1465 0.180667
R15341 VDAC_N.n1467 VDAC_N.n1466 0.180667
R15342 VDAC_N.n1468 VDAC_N.n1467 0.180667
R15343 VDAC_N.n1469 VDAC_N.n1468 0.180667
R15344 VDAC_N.n1470 VDAC_N.n1469 0.180667
R15345 VDAC_N.n1471 VDAC_N.n1470 0.180667
R15346 VDAC_N.n1472 VDAC_N.n1471 0.180667
R15347 VDAC_N.n1473 VDAC_N.n1472 0.180667
R15348 VDAC_N.n1474 VDAC_N.n1473 0.180667
R15349 VDAC_N.n1475 VDAC_N.n1474 0.180667
R15350 VDAC_N.n1476 VDAC_N.n1475 0.180667
R15351 VDAC_N.n1477 VDAC_N.n1476 0.180667
R15352 VDAC_N.n1478 VDAC_N.n1477 0.180667
R15353 VDAC_N.n1479 VDAC_N.n1478 0.180667
R15354 VDAC_N.n1480 VDAC_N.n1479 0.180667
R15355 VDAC_N.n1481 VDAC_N.n1480 0.180667
R15356 VDAC_N.n1482 VDAC_N.n1481 0.180667
R15357 VDAC_N.n1483 VDAC_N.n1482 0.180667
R15358 VDAC_N.n1484 VDAC_N.n1483 0.180667
R15359 VDAC_N.n1485 VDAC_N.n1484 0.180667
R15360 VDAC_N.n1486 VDAC_N.n1485 0.180667
R15361 VDAC_N.n1487 VDAC_N.n1486 0.180667
R15362 VDAC_N.n1488 VDAC_N.n1487 0.180667
R15363 VDAC_N.n1489 VDAC_N.n1488 0.180667
R15364 VDAC_N.n1490 VDAC_N.n1489 0.180667
R15365 VDAC_N.n1491 VDAC_N.n1490 0.180667
R15366 VDAC_N.n1492 VDAC_N.n1491 0.180667
R15367 VDAC_N.n1493 VDAC_N.n1492 0.180667
R15368 VDAC_N.n1494 VDAC_N.n1493 0.180667
R15369 VDAC_N.n1495 VDAC_N.n1494 0.180667
R15370 VDAC_N.n1496 VDAC_N.n1495 0.180667
R15371 VDAC_N.n1497 VDAC_N.n1496 0.180667
R15372 VDAC_N.n1498 VDAC_N.n1497 0.180667
R15373 VDAC_N.n1499 VDAC_N.n1498 0.180667
R15374 VDAC_N.n1500 VDAC_N.n1499 0.180667
R15375 VDAC_N.n1501 VDAC_N.n1500 0.180667
R15376 VDAC_N.n1502 VDAC_N.n1501 0.180667
R15377 VDAC_N.n1503 VDAC_N.n94 0.180667
R15378 VDAC_N.n1504 VDAC_N.n1503 0.180667
R15379 VDAC_N.n1505 VDAC_N.n1504 0.180667
R15380 VDAC_N.n1506 VDAC_N.n1505 0.180667
R15381 VDAC_N.n1507 VDAC_N.n1506 0.180667
R15382 VDAC_N.n1508 VDAC_N.n1507 0.180667
R15383 VDAC_N.n1509 VDAC_N.n1508 0.180667
R15384 VDAC_N.n1510 VDAC_N.n1509 0.180667
R15385 VDAC_N.n1511 VDAC_N.n1510 0.180667
R15386 VDAC_N.n1512 VDAC_N.n1511 0.180667
R15387 VDAC_N.n1513 VDAC_N.n1512 0.180667
R15388 VDAC_N.n1514 VDAC_N.n1513 0.180667
R15389 VDAC_N.n1515 VDAC_N.n1514 0.180667
R15390 VDAC_N.n1516 VDAC_N.n1515 0.180667
R15391 VDAC_N.n1517 VDAC_N.n1516 0.180667
R15392 VDAC_N.n1518 VDAC_N.n1517 0.180667
R15393 VDAC_N.n1519 VDAC_N.n1518 0.180667
R15394 VDAC_N.n1520 VDAC_N.n1519 0.180667
R15395 VDAC_N.n1521 VDAC_N.n1520 0.180667
R15396 VDAC_N.n1522 VDAC_N.n1521 0.180667
R15397 VDAC_N.n1523 VDAC_N.n1522 0.180667
R15398 VDAC_N.n1524 VDAC_N.n1523 0.180667
R15399 VDAC_N.n1525 VDAC_N.n1524 0.180667
R15400 VDAC_N.n1526 VDAC_N.n1525 0.180667
R15401 VDAC_N.n1527 VDAC_N.n1526 0.180667
R15402 VDAC_N.n1528 VDAC_N.n1527 0.180667
R15403 VDAC_N.n1529 VDAC_N.n1528 0.180667
R15404 VDAC_N.n1530 VDAC_N.n1529 0.180667
R15405 VDAC_N.n1531 VDAC_N.n1530 0.180667
R15406 VDAC_N.n1532 VDAC_N.n1531 0.180667
R15407 VDAC_N.n1533 VDAC_N.n1532 0.180667
R15408 VDAC_N.n1534 VDAC_N.n1533 0.180667
R15409 VDAC_N.n1535 VDAC_N.n1534 0.180667
R15410 VDAC_N.n1536 VDAC_N.n1535 0.180667
R15411 VDAC_N.n1537 VDAC_N.n1536 0.180667
R15412 VDAC_N.n1538 VDAC_N.n1537 0.180667
R15413 VDAC_N.n1539 VDAC_N.n1538 0.180667
R15414 VDAC_N.n1540 VDAC_N.n1539 0.180667
R15415 VDAC_N.n1541 VDAC_N.n1540 0.180667
R15416 VDAC_N.n1542 VDAC_N.n1541 0.180667
R15417 VDAC_N.n1543 VDAC_N.n1542 0.180667
R15418 VDAC_N.n1544 VDAC_N.n1543 0.180667
R15419 VDAC_N.n1545 VDAC_N.n1544 0.180667
R15420 VDAC_N.n1546 VDAC_N.n1545 0.180667
R15421 VDAC_N.n1547 VDAC_N.n1546 0.180667
R15422 VDAC_N.n1548 VDAC_N.n1547 0.180667
R15423 VDAC_N.n1549 VDAC_N.n1548 0.180667
R15424 VDAC_N.n1550 VDAC_N.n1549 0.180667
R15425 VDAC_N.n1551 VDAC_N.n1550 0.180667
R15426 VDAC_N.n1552 VDAC_N.n1551 0.180667
R15427 VDAC_N.n1553 VDAC_N.n1552 0.180667
R15428 VDAC_N.n1554 VDAC_N.n1553 0.180667
R15429 VDAC_N.n1555 VDAC_N.n1554 0.180667
R15430 VDAC_N.n1556 VDAC_N.n1555 0.180667
R15431 VDAC_N.n1557 VDAC_N.n1556 0.180667
R15432 VDAC_N.n1558 VDAC_N.n1557 0.180667
R15433 VDAC_N.n1559 VDAC_N.n1558 0.180667
R15434 VDAC_N.n1560 VDAC_N.n1559 0.180667
R15435 VDAC_N.n1561 VDAC_N.n1560 0.180667
R15436 VDAC_N.n1562 VDAC_N.n1561 0.180667
R15437 VDAC_N.n1563 VDAC_N.n1562 0.180667
R15438 VDAC_N.n1564 VDAC_N.n1563 0.180667
R15439 VDAC_N.n1565 VDAC_N.n1564 0.180667
R15440 VDAC_N.n1566 VDAC_N.n93 0.180667
R15441 VDAC_N.n1567 VDAC_N.n1566 0.180667
R15442 VDAC_N.n1568 VDAC_N.n1567 0.180667
R15443 VDAC_N.n1569 VDAC_N.n1568 0.180667
R15444 VDAC_N.n1570 VDAC_N.n1569 0.180667
R15445 VDAC_N.n1571 VDAC_N.n1570 0.180667
R15446 VDAC_N.n1572 VDAC_N.n1571 0.180667
R15447 VDAC_N.n1573 VDAC_N.n1572 0.180667
R15448 VDAC_N.n1574 VDAC_N.n1573 0.180667
R15449 VDAC_N.n1575 VDAC_N.n1574 0.180667
R15450 VDAC_N.n1576 VDAC_N.n1575 0.180667
R15451 VDAC_N.n1577 VDAC_N.n1576 0.180667
R15452 VDAC_N.n1578 VDAC_N.n1577 0.180667
R15453 VDAC_N.n1579 VDAC_N.n1578 0.180667
R15454 VDAC_N.n1580 VDAC_N.n1579 0.180667
R15455 VDAC_N.n1581 VDAC_N.n1580 0.180667
R15456 VDAC_N.n1582 VDAC_N.n1581 0.180667
R15457 VDAC_N.n1583 VDAC_N.n1582 0.180667
R15458 VDAC_N.n1584 VDAC_N.n1583 0.180667
R15459 VDAC_N.n1585 VDAC_N.n1584 0.180667
R15460 VDAC_N.n1586 VDAC_N.n1585 0.180667
R15461 VDAC_N.n1587 VDAC_N.n1586 0.180667
R15462 VDAC_N.n1588 VDAC_N.n1587 0.180667
R15463 VDAC_N.n1589 VDAC_N.n1588 0.180667
R15464 VDAC_N.n1590 VDAC_N.n1589 0.180667
R15465 VDAC_N.n1591 VDAC_N.n1590 0.180667
R15466 VDAC_N.n1592 VDAC_N.n1591 0.180667
R15467 VDAC_N.n1593 VDAC_N.n1592 0.180667
R15468 VDAC_N.n1594 VDAC_N.n1593 0.180667
R15469 VDAC_N.n1595 VDAC_N.n1594 0.180667
R15470 VDAC_N.n1596 VDAC_N.n1595 0.180667
R15471 VDAC_N.n1597 VDAC_N.n1596 0.180667
R15472 VDAC_N.n1598 VDAC_N.n1597 0.180667
R15473 VDAC_N.n1599 VDAC_N.n1598 0.180667
R15474 VDAC_N.n1600 VDAC_N.n1599 0.180667
R15475 VDAC_N.n1601 VDAC_N.n1600 0.180667
R15476 VDAC_N.n1602 VDAC_N.n1601 0.180667
R15477 VDAC_N.n1603 VDAC_N.n1602 0.180667
R15478 VDAC_N.n1604 VDAC_N.n1603 0.180667
R15479 VDAC_N.n1605 VDAC_N.n1604 0.180667
R15480 VDAC_N.n1606 VDAC_N.n1605 0.180667
R15481 VDAC_N.n1607 VDAC_N.n1606 0.180667
R15482 VDAC_N.n1608 VDAC_N.n1607 0.180667
R15483 VDAC_N.n1609 VDAC_N.n1608 0.180667
R15484 VDAC_N.n1610 VDAC_N.n1609 0.180667
R15485 VDAC_N.n1611 VDAC_N.n1610 0.180667
R15486 VDAC_N.n1612 VDAC_N.n1611 0.180667
R15487 VDAC_N.n1613 VDAC_N.n1612 0.180667
R15488 VDAC_N.n1614 VDAC_N.n1613 0.180667
R15489 VDAC_N.n1615 VDAC_N.n1614 0.180667
R15490 VDAC_N.n1616 VDAC_N.n1615 0.180667
R15491 VDAC_N.n1617 VDAC_N.n1616 0.180667
R15492 VDAC_N.n1618 VDAC_N.n1617 0.180667
R15493 VDAC_N.n1619 VDAC_N.n1618 0.180667
R15494 VDAC_N.n1620 VDAC_N.n1619 0.180667
R15495 VDAC_N.n1621 VDAC_N.n1620 0.180667
R15496 VDAC_N.n1622 VDAC_N.n1621 0.180667
R15497 VDAC_N.n1623 VDAC_N.n1622 0.180667
R15498 VDAC_N.n1624 VDAC_N.n1623 0.180667
R15499 VDAC_N.n1625 VDAC_N.n1624 0.180667
R15500 VDAC_N.n1626 VDAC_N.n1625 0.180667
R15501 VDAC_N.n1627 VDAC_N.n1626 0.180667
R15502 VDAC_N.n1628 VDAC_N.n1627 0.180667
R15503 VDAC_N.n1629 VDAC_N.n92 0.180667
R15504 VDAC_N.n1630 VDAC_N.n1629 0.180667
R15505 VDAC_N.n1631 VDAC_N.n1630 0.180667
R15506 VDAC_N.n1632 VDAC_N.n1631 0.180667
R15507 VDAC_N.n1633 VDAC_N.n1632 0.180667
R15508 VDAC_N.n1634 VDAC_N.n1633 0.180667
R15509 VDAC_N.n1635 VDAC_N.n1634 0.180667
R15510 VDAC_N.n1636 VDAC_N.n1635 0.180667
R15511 VDAC_N.n1637 VDAC_N.n1636 0.180667
R15512 VDAC_N.n1638 VDAC_N.n1637 0.180667
R15513 VDAC_N.n1639 VDAC_N.n1638 0.180667
R15514 VDAC_N.n1640 VDAC_N.n1639 0.180667
R15515 VDAC_N.n1641 VDAC_N.n1640 0.180667
R15516 VDAC_N.n1642 VDAC_N.n1641 0.180667
R15517 VDAC_N.n1643 VDAC_N.n1642 0.180667
R15518 VDAC_N.n1644 VDAC_N.n1643 0.180667
R15519 VDAC_N.n1645 VDAC_N.n1644 0.180667
R15520 VDAC_N.n1646 VDAC_N.n1645 0.180667
R15521 VDAC_N.n1647 VDAC_N.n1646 0.180667
R15522 VDAC_N.n1648 VDAC_N.n1647 0.180667
R15523 VDAC_N.n1649 VDAC_N.n1648 0.180667
R15524 VDAC_N.n1650 VDAC_N.n1649 0.180667
R15525 VDAC_N.n1651 VDAC_N.n1650 0.180667
R15526 VDAC_N.n1652 VDAC_N.n1651 0.180667
R15527 VDAC_N.n1653 VDAC_N.n1652 0.180667
R15528 VDAC_N.n1654 VDAC_N.n1653 0.180667
R15529 VDAC_N.n1655 VDAC_N.n1654 0.180667
R15530 VDAC_N.n1656 VDAC_N.n1655 0.180667
R15531 VDAC_N.n1657 VDAC_N.n1656 0.180667
R15532 VDAC_N.n1658 VDAC_N.n1657 0.180667
R15533 VDAC_N.n1659 VDAC_N.n1658 0.180667
R15534 VDAC_N.n1660 VDAC_N.n1659 0.180667
R15535 VDAC_N.n1661 VDAC_N.n1660 0.180667
R15536 VDAC_N.n1662 VDAC_N.n1661 0.180667
R15537 VDAC_N.n1663 VDAC_N.n1662 0.180667
R15538 VDAC_N.n1664 VDAC_N.n1663 0.180667
R15539 VDAC_N.n1665 VDAC_N.n1664 0.180667
R15540 VDAC_N.n1666 VDAC_N.n1665 0.180667
R15541 VDAC_N.n1667 VDAC_N.n1666 0.180667
R15542 VDAC_N.n1668 VDAC_N.n1667 0.180667
R15543 VDAC_N.n1669 VDAC_N.n1668 0.180667
R15544 VDAC_N.n1670 VDAC_N.n1669 0.180667
R15545 VDAC_N.n1671 VDAC_N.n1670 0.180667
R15546 VDAC_N.n1672 VDAC_N.n1671 0.180667
R15547 VDAC_N.n1673 VDAC_N.n1672 0.180667
R15548 VDAC_N.n1674 VDAC_N.n1673 0.180667
R15549 VDAC_N.n1675 VDAC_N.n1674 0.180667
R15550 VDAC_N.n1676 VDAC_N.n1675 0.180667
R15551 VDAC_N.n1677 VDAC_N.n1676 0.180667
R15552 VDAC_N.n1678 VDAC_N.n1677 0.180667
R15553 VDAC_N.n1679 VDAC_N.n1678 0.180667
R15554 VDAC_N.n1680 VDAC_N.n1679 0.180667
R15555 VDAC_N.n1681 VDAC_N.n1680 0.180667
R15556 VDAC_N.n1682 VDAC_N.n1681 0.180667
R15557 VDAC_N.n1683 VDAC_N.n1682 0.180667
R15558 VDAC_N.n1684 VDAC_N.n1683 0.180667
R15559 VDAC_N.n1685 VDAC_N.n1684 0.180667
R15560 VDAC_N.n1686 VDAC_N.n1685 0.180667
R15561 VDAC_N.n1687 VDAC_N.n1686 0.180667
R15562 VDAC_N.n1688 VDAC_N.n1687 0.180667
R15563 VDAC_N.n1689 VDAC_N.n1688 0.180667
R15564 VDAC_N.n1690 VDAC_N.n1689 0.180667
R15565 VDAC_N.n1691 VDAC_N.n1690 0.180667
R15566 VDAC_N.n1692 VDAC_N.n91 0.180667
R15567 VDAC_N.n1693 VDAC_N.n1692 0.180667
R15568 VDAC_N.n1694 VDAC_N.n1693 0.180667
R15569 VDAC_N.n1695 VDAC_N.n1694 0.180667
R15570 VDAC_N.n1696 VDAC_N.n1695 0.180667
R15571 VDAC_N.n1697 VDAC_N.n1696 0.180667
R15572 VDAC_N.n1698 VDAC_N.n1697 0.180667
R15573 VDAC_N.n1699 VDAC_N.n1698 0.180667
R15574 VDAC_N.n1700 VDAC_N.n1699 0.180667
R15575 VDAC_N.n1701 VDAC_N.n1700 0.180667
R15576 VDAC_N.n1702 VDAC_N.n1701 0.180667
R15577 VDAC_N.n1703 VDAC_N.n1702 0.180667
R15578 VDAC_N.n1704 VDAC_N.n1703 0.180667
R15579 VDAC_N.n1705 VDAC_N.n1704 0.180667
R15580 VDAC_N.n1706 VDAC_N.n1705 0.180667
R15581 VDAC_N.n1707 VDAC_N.n1706 0.180667
R15582 VDAC_N.n1708 VDAC_N.n1707 0.180667
R15583 VDAC_N.n1709 VDAC_N.n1708 0.180667
R15584 VDAC_N.n1710 VDAC_N.n1709 0.180667
R15585 VDAC_N.n1711 VDAC_N.n1710 0.180667
R15586 VDAC_N.n1712 VDAC_N.n1711 0.180667
R15587 VDAC_N.n1713 VDAC_N.n1712 0.180667
R15588 VDAC_N.n1714 VDAC_N.n1713 0.180667
R15589 VDAC_N.n1715 VDAC_N.n1714 0.180667
R15590 VDAC_N.n1716 VDAC_N.n1715 0.180667
R15591 VDAC_N.n1717 VDAC_N.n1716 0.180667
R15592 VDAC_N.n1718 VDAC_N.n1717 0.180667
R15593 VDAC_N.n1719 VDAC_N.n1718 0.180667
R15594 VDAC_N.n1720 VDAC_N.n1719 0.180667
R15595 VDAC_N.n1721 VDAC_N.n1720 0.180667
R15596 VDAC_N.n1722 VDAC_N.n1721 0.180667
R15597 VDAC_N.n1723 VDAC_N.n1722 0.180667
R15598 VDAC_N.n1724 VDAC_N.n1723 0.180667
R15599 VDAC_N.n1725 VDAC_N.n1724 0.180667
R15600 VDAC_N.n1726 VDAC_N.n1725 0.180667
R15601 VDAC_N.n1727 VDAC_N.n1726 0.180667
R15602 VDAC_N.n1728 VDAC_N.n1727 0.180667
R15603 VDAC_N.n1729 VDAC_N.n1728 0.180667
R15604 VDAC_N.n1730 VDAC_N.n1729 0.180667
R15605 VDAC_N.n1731 VDAC_N.n1730 0.180667
R15606 VDAC_N.n1732 VDAC_N.n1731 0.180667
R15607 VDAC_N.n1733 VDAC_N.n1732 0.180667
R15608 VDAC_N.n1734 VDAC_N.n1733 0.180667
R15609 VDAC_N.n1735 VDAC_N.n1734 0.180667
R15610 VDAC_N.n1736 VDAC_N.n1735 0.180667
R15611 VDAC_N.n1737 VDAC_N.n1736 0.180667
R15612 VDAC_N.n1738 VDAC_N.n1737 0.180667
R15613 VDAC_N.n1739 VDAC_N.n1738 0.180667
R15614 VDAC_N.n1740 VDAC_N.n1739 0.180667
R15615 VDAC_N.n1741 VDAC_N.n1740 0.180667
R15616 VDAC_N.n1742 VDAC_N.n1741 0.180667
R15617 VDAC_N.n1743 VDAC_N.n1742 0.180667
R15618 VDAC_N.n1744 VDAC_N.n1743 0.180667
R15619 VDAC_N.n1745 VDAC_N.n1744 0.180667
R15620 VDAC_N.n1746 VDAC_N.n1745 0.180667
R15621 VDAC_N.n1747 VDAC_N.n1746 0.180667
R15622 VDAC_N.n1748 VDAC_N.n1747 0.180667
R15623 VDAC_N.n1749 VDAC_N.n1748 0.180667
R15624 VDAC_N.n1750 VDAC_N.n1749 0.180667
R15625 VDAC_N.n1751 VDAC_N.n1750 0.180667
R15626 VDAC_N.n1752 VDAC_N.n1751 0.180667
R15627 VDAC_N.n1753 VDAC_N.n1752 0.180667
R15628 VDAC_N.n1754 VDAC_N.n1753 0.180667
R15629 VDAC_N.n1755 VDAC_N.n90 0.180667
R15630 VDAC_N.n1756 VDAC_N.n1755 0.180667
R15631 VDAC_N.n1757 VDAC_N.n1756 0.180667
R15632 VDAC_N.n1758 VDAC_N.n1757 0.180667
R15633 VDAC_N.n1759 VDAC_N.n1758 0.180667
R15634 VDAC_N.n1760 VDAC_N.n1759 0.180667
R15635 VDAC_N.n1761 VDAC_N.n1760 0.180667
R15636 VDAC_N.n1762 VDAC_N.n1761 0.180667
R15637 VDAC_N.n1763 VDAC_N.n1762 0.180667
R15638 VDAC_N.n1764 VDAC_N.n1763 0.180667
R15639 VDAC_N.n1765 VDAC_N.n1764 0.180667
R15640 VDAC_N.n1766 VDAC_N.n1765 0.180667
R15641 VDAC_N.n1767 VDAC_N.n1766 0.180667
R15642 VDAC_N.n1768 VDAC_N.n1767 0.180667
R15643 VDAC_N.n1769 VDAC_N.n1768 0.180667
R15644 VDAC_N.n1770 VDAC_N.n1769 0.180667
R15645 VDAC_N.n1771 VDAC_N.n1770 0.180667
R15646 VDAC_N.n1772 VDAC_N.n1771 0.180667
R15647 VDAC_N.n1773 VDAC_N.n1772 0.180667
R15648 VDAC_N.n1774 VDAC_N.n1773 0.180667
R15649 VDAC_N.n1775 VDAC_N.n1774 0.180667
R15650 VDAC_N.n1776 VDAC_N.n1775 0.180667
R15651 VDAC_N.n1777 VDAC_N.n1776 0.180667
R15652 VDAC_N.n1778 VDAC_N.n1777 0.180667
R15653 VDAC_N.n1779 VDAC_N.n1778 0.180667
R15654 VDAC_N.n1780 VDAC_N.n1779 0.180667
R15655 VDAC_N.n1781 VDAC_N.n1780 0.180667
R15656 VDAC_N.n1782 VDAC_N.n1781 0.180667
R15657 VDAC_N.n1783 VDAC_N.n1782 0.180667
R15658 VDAC_N.n1784 VDAC_N.n1783 0.180667
R15659 VDAC_N.n1785 VDAC_N.n1784 0.180667
R15660 VDAC_N.n1786 VDAC_N.n1785 0.180667
R15661 VDAC_N.n1787 VDAC_N.n1786 0.180667
R15662 VDAC_N.n1788 VDAC_N.n1787 0.180667
R15663 VDAC_N.n1789 VDAC_N.n1788 0.180667
R15664 VDAC_N.n1790 VDAC_N.n1789 0.180667
R15665 VDAC_N.n1791 VDAC_N.n1790 0.180667
R15666 VDAC_N.n1792 VDAC_N.n1791 0.180667
R15667 VDAC_N.n1793 VDAC_N.n1792 0.180667
R15668 VDAC_N.n1794 VDAC_N.n1793 0.180667
R15669 VDAC_N.n1795 VDAC_N.n1794 0.180667
R15670 VDAC_N.n1796 VDAC_N.n1795 0.180667
R15671 VDAC_N.n1797 VDAC_N.n1796 0.180667
R15672 VDAC_N.n1798 VDAC_N.n1797 0.180667
R15673 VDAC_N.n1799 VDAC_N.n1798 0.180667
R15674 VDAC_N.n1800 VDAC_N.n1799 0.180667
R15675 VDAC_N.n1801 VDAC_N.n1800 0.180667
R15676 VDAC_N.n1802 VDAC_N.n1801 0.180667
R15677 VDAC_N.n1803 VDAC_N.n1802 0.180667
R15678 VDAC_N.n1804 VDAC_N.n1803 0.180667
R15679 VDAC_N.n1805 VDAC_N.n1804 0.180667
R15680 VDAC_N.n1806 VDAC_N.n1805 0.180667
R15681 VDAC_N.n1807 VDAC_N.n1806 0.180667
R15682 VDAC_N.n1808 VDAC_N.n1807 0.180667
R15683 VDAC_N.n1809 VDAC_N.n1808 0.180667
R15684 VDAC_N.n1810 VDAC_N.n1809 0.180667
R15685 VDAC_N.n1811 VDAC_N.n1810 0.180667
R15686 VDAC_N.n1812 VDAC_N.n1811 0.180667
R15687 VDAC_N.n1813 VDAC_N.n1812 0.180667
R15688 VDAC_N.n1814 VDAC_N.n1813 0.180667
R15689 VDAC_N.n1815 VDAC_N.n1814 0.180667
R15690 VDAC_N.n1816 VDAC_N.n1815 0.180667
R15691 VDAC_N.n1817 VDAC_N.n1816 0.180667
R15692 VDAC_N.n1818 VDAC_N.n89 0.180667
R15693 VDAC_N.n1819 VDAC_N.n1818 0.180667
R15694 VDAC_N.n1820 VDAC_N.n1819 0.180667
R15695 VDAC_N.n1821 VDAC_N.n1820 0.180667
R15696 VDAC_N.n1822 VDAC_N.n1821 0.180667
R15697 VDAC_N.n1823 VDAC_N.n1822 0.180667
R15698 VDAC_N.n1824 VDAC_N.n1823 0.180667
R15699 VDAC_N.n1825 VDAC_N.n1824 0.180667
R15700 VDAC_N.n1826 VDAC_N.n1825 0.180667
R15701 VDAC_N.n1827 VDAC_N.n1826 0.180667
R15702 VDAC_N.n1828 VDAC_N.n1827 0.180667
R15703 VDAC_N.n1829 VDAC_N.n1828 0.180667
R15704 VDAC_N.n1830 VDAC_N.n1829 0.180667
R15705 VDAC_N.n1831 VDAC_N.n1830 0.180667
R15706 VDAC_N.n1832 VDAC_N.n1831 0.180667
R15707 VDAC_N.n1833 VDAC_N.n1832 0.180667
R15708 VDAC_N.n1834 VDAC_N.n1833 0.180667
R15709 VDAC_N.n1835 VDAC_N.n1834 0.180667
R15710 VDAC_N.n1836 VDAC_N.n1835 0.180667
R15711 VDAC_N.n1837 VDAC_N.n1836 0.180667
R15712 VDAC_N.n1838 VDAC_N.n1837 0.180667
R15713 VDAC_N.n1839 VDAC_N.n1838 0.180667
R15714 VDAC_N.n1840 VDAC_N.n1839 0.180667
R15715 VDAC_N.n1841 VDAC_N.n1840 0.180667
R15716 VDAC_N.n1842 VDAC_N.n1841 0.180667
R15717 VDAC_N.n1843 VDAC_N.n1842 0.180667
R15718 VDAC_N.n1844 VDAC_N.n1843 0.180667
R15719 VDAC_N.n1845 VDAC_N.n1844 0.180667
R15720 VDAC_N.n1846 VDAC_N.n1845 0.180667
R15721 VDAC_N.n1847 VDAC_N.n1846 0.180667
R15722 VDAC_N.n1848 VDAC_N.n1847 0.180667
R15723 VDAC_N.n1849 VDAC_N.n1848 0.180667
R15724 VDAC_N.n1850 VDAC_N.n1849 0.180667
R15725 VDAC_N.n1851 VDAC_N.n1850 0.180667
R15726 VDAC_N.n1852 VDAC_N.n1851 0.180667
R15727 VDAC_N.n1853 VDAC_N.n1852 0.180667
R15728 VDAC_N.n1854 VDAC_N.n1853 0.180667
R15729 VDAC_N.n1855 VDAC_N.n1854 0.180667
R15730 VDAC_N.n1856 VDAC_N.n1855 0.180667
R15731 VDAC_N.n1857 VDAC_N.n1856 0.180667
R15732 VDAC_N.n1858 VDAC_N.n1857 0.180667
R15733 VDAC_N.n1859 VDAC_N.n1858 0.180667
R15734 VDAC_N.n1860 VDAC_N.n1859 0.180667
R15735 VDAC_N.n1861 VDAC_N.n1860 0.180667
R15736 VDAC_N.n1862 VDAC_N.n1861 0.180667
R15737 VDAC_N.n1863 VDAC_N.n1862 0.180667
R15738 VDAC_N.n1864 VDAC_N.n1863 0.180667
R15739 VDAC_N.n1865 VDAC_N.n1864 0.180667
R15740 VDAC_N.n1866 VDAC_N.n1865 0.180667
R15741 VDAC_N.n1867 VDAC_N.n1866 0.180667
R15742 VDAC_N.n1868 VDAC_N.n1867 0.180667
R15743 VDAC_N.n1869 VDAC_N.n1868 0.180667
R15744 VDAC_N.n1870 VDAC_N.n1869 0.180667
R15745 VDAC_N.n1871 VDAC_N.n1870 0.180667
R15746 VDAC_N.n1872 VDAC_N.n1871 0.180667
R15747 VDAC_N.n1873 VDAC_N.n1872 0.180667
R15748 VDAC_N.n1874 VDAC_N.n1873 0.180667
R15749 VDAC_N.n1875 VDAC_N.n1874 0.180667
R15750 VDAC_N.n1876 VDAC_N.n1875 0.180667
R15751 VDAC_N.n1877 VDAC_N.n1876 0.180667
R15752 VDAC_N.n1878 VDAC_N.n1877 0.180667
R15753 VDAC_N.n1879 VDAC_N.n1878 0.180667
R15754 VDAC_N.n1880 VDAC_N.n1879 0.180667
R15755 VDAC_N.n1881 VDAC_N.n88 0.180667
R15756 VDAC_N.n1882 VDAC_N.n1881 0.180667
R15757 VDAC_N.n1883 VDAC_N.n1882 0.180667
R15758 VDAC_N.n1884 VDAC_N.n1883 0.180667
R15759 VDAC_N.n1885 VDAC_N.n1884 0.180667
R15760 VDAC_N.n1886 VDAC_N.n1885 0.180667
R15761 VDAC_N.n1887 VDAC_N.n1886 0.180667
R15762 VDAC_N.n1888 VDAC_N.n1887 0.180667
R15763 VDAC_N.n1889 VDAC_N.n1888 0.180667
R15764 VDAC_N.n1890 VDAC_N.n1889 0.180667
R15765 VDAC_N.n1891 VDAC_N.n1890 0.180667
R15766 VDAC_N.n1892 VDAC_N.n1891 0.180667
R15767 VDAC_N.n1893 VDAC_N.n1892 0.180667
R15768 VDAC_N.n1894 VDAC_N.n1893 0.180667
R15769 VDAC_N.n1895 VDAC_N.n1894 0.180667
R15770 VDAC_N.n1896 VDAC_N.n1895 0.180667
R15771 VDAC_N.n1897 VDAC_N.n1896 0.180667
R15772 VDAC_N.n1898 VDAC_N.n1897 0.180667
R15773 VDAC_N.n1899 VDAC_N.n1898 0.180667
R15774 VDAC_N.n1900 VDAC_N.n1899 0.180667
R15775 VDAC_N.n1901 VDAC_N.n1900 0.180667
R15776 VDAC_N.n1902 VDAC_N.n1901 0.180667
R15777 VDAC_N.n1903 VDAC_N.n1902 0.180667
R15778 VDAC_N.n1904 VDAC_N.n1903 0.180667
R15779 VDAC_N.n1905 VDAC_N.n1904 0.180667
R15780 VDAC_N.n1906 VDAC_N.n1905 0.180667
R15781 VDAC_N.n1907 VDAC_N.n1906 0.180667
R15782 VDAC_N.n1908 VDAC_N.n1907 0.180667
R15783 VDAC_N.n1909 VDAC_N.n1908 0.180667
R15784 VDAC_N.n1910 VDAC_N.n1909 0.180667
R15785 VDAC_N.n1911 VDAC_N.n1910 0.180667
R15786 VDAC_N.n1912 VDAC_N.n1911 0.180667
R15787 VDAC_N.n1913 VDAC_N.n1912 0.180667
R15788 VDAC_N.n1914 VDAC_N.n1913 0.180667
R15789 VDAC_N.n1915 VDAC_N.n1914 0.180667
R15790 VDAC_N.n1916 VDAC_N.n1915 0.180667
R15791 VDAC_N.n1917 VDAC_N.n1916 0.180667
R15792 VDAC_N.n1918 VDAC_N.n1917 0.180667
R15793 VDAC_N.n1919 VDAC_N.n1918 0.180667
R15794 VDAC_N.n1920 VDAC_N.n1919 0.180667
R15795 VDAC_N.n1921 VDAC_N.n1920 0.180667
R15796 VDAC_N.n1922 VDAC_N.n1921 0.180667
R15797 VDAC_N.n1923 VDAC_N.n1922 0.180667
R15798 VDAC_N.n1924 VDAC_N.n1923 0.180667
R15799 VDAC_N.n1925 VDAC_N.n1924 0.180667
R15800 VDAC_N.n1926 VDAC_N.n1925 0.180667
R15801 VDAC_N.n1927 VDAC_N.n1926 0.180667
R15802 VDAC_N.n1928 VDAC_N.n1927 0.180667
R15803 VDAC_N.n1929 VDAC_N.n1928 0.180667
R15804 VDAC_N.n1930 VDAC_N.n1929 0.180667
R15805 VDAC_N.n1931 VDAC_N.n1930 0.180667
R15806 VDAC_N.n1932 VDAC_N.n1931 0.180667
R15807 VDAC_N.n1933 VDAC_N.n1932 0.180667
R15808 VDAC_N.n1934 VDAC_N.n1933 0.180667
R15809 VDAC_N.n1935 VDAC_N.n1934 0.180667
R15810 VDAC_N.n1936 VDAC_N.n1935 0.180667
R15811 VDAC_N.n1937 VDAC_N.n1936 0.180667
R15812 VDAC_N.n1938 VDAC_N.n1937 0.180667
R15813 VDAC_N.n1939 VDAC_N.n1938 0.180667
R15814 VDAC_N.n1940 VDAC_N.n1939 0.180667
R15815 VDAC_N.n1941 VDAC_N.n1940 0.180667
R15816 VDAC_N.n1942 VDAC_N.n1941 0.180667
R15817 VDAC_N.n1943 VDAC_N.n1942 0.180667
R15818 VDAC_N.n87 VDAC_N.n86 0.180667
R15819 VDAC_N.n86 VDAC_N.n85 0.180667
R15820 VDAC_N.n85 VDAC_N.n84 0.180667
R15821 VDAC_N.n84 VDAC_N.n83 0.180667
R15822 VDAC_N.n83 VDAC_N.n82 0.180667
R15823 VDAC_N.n82 VDAC_N.n81 0.180667
R15824 VDAC_N.n81 VDAC_N.n80 0.180667
R15825 VDAC_N.n80 VDAC_N.n79 0.180667
R15826 VDAC_N.n79 VDAC_N.n78 0.180667
R15827 VDAC_N.n78 VDAC_N.n77 0.180667
R15828 VDAC_N.n77 VDAC_N.n76 0.180667
R15829 VDAC_N.n76 VDAC_N.n75 0.180667
R15830 VDAC_N.n75 VDAC_N.n74 0.180667
R15831 VDAC_N.n74 VDAC_N.n73 0.180667
R15832 VDAC_N.n73 VDAC_N.n72 0.180667
R15833 VDAC_N.n72 VDAC_N.n71 0.180667
R15834 VDAC_N.n71 VDAC_N.n70 0.180667
R15835 VDAC_N.n70 VDAC_N.n69 0.180667
R15836 VDAC_N.n69 VDAC_N.n68 0.180667
R15837 VDAC_N.n68 VDAC_N.n67 0.180667
R15838 VDAC_N.n67 VDAC_N.n66 0.180667
R15839 VDAC_N.n66 VDAC_N.n65 0.180667
R15840 VDAC_N.n65 VDAC_N.n64 0.180667
R15841 VDAC_N.n64 VDAC_N.n63 0.180667
R15842 VDAC_N.n63 VDAC_N.n62 0.180667
R15843 VDAC_N.n62 VDAC_N.n61 0.180667
R15844 VDAC_N.n61 VDAC_N.n60 0.180667
R15845 VDAC_N.n60 VDAC_N.n59 0.180667
R15846 VDAC_N.n59 VDAC_N.n58 0.180667
R15847 VDAC_N.n58 VDAC_N.n57 0.180667
R15848 VDAC_N.n57 VDAC_N.n56 0.180667
R15849 VDAC_N.n56 VDAC_N.n55 0.180667
R15850 VDAC_N.n55 VDAC_N.n54 0.180667
R15851 VDAC_N.n54 VDAC_N.n53 0.180667
R15852 VDAC_N.n53 VDAC_N.n52 0.180667
R15853 VDAC_N.n52 VDAC_N.n51 0.180667
R15854 VDAC_N.n51 VDAC_N.n50 0.180667
R15855 VDAC_N.n50 VDAC_N.n49 0.180667
R15856 VDAC_N.n49 VDAC_N.n48 0.180667
R15857 VDAC_N.n48 VDAC_N.n47 0.180667
R15858 VDAC_N.n47 VDAC_N.n46 0.180667
R15859 VDAC_N.n46 VDAC_N.n45 0.180667
R15860 VDAC_N.n45 VDAC_N.n44 0.180667
R15861 VDAC_N.n44 VDAC_N.n43 0.180667
R15862 VDAC_N.n43 VDAC_N.n42 0.180667
R15863 VDAC_N.n42 VDAC_N.n41 0.180667
R15864 VDAC_N.n41 VDAC_N.n40 0.180667
R15865 VDAC_N.n40 VDAC_N.n39 0.180667
R15866 VDAC_N.n39 VDAC_N.n38 0.180667
R15867 VDAC_N.n38 VDAC_N.n37 0.180667
R15868 VDAC_N.n37 VDAC_N.n36 0.180667
R15869 VDAC_N.n36 VDAC_N.n35 0.180667
R15870 VDAC_N.n35 VDAC_N.n34 0.180667
R15871 VDAC_N.n34 VDAC_N.n33 0.180667
R15872 VDAC_N.n33 VDAC_N.n32 0.180667
R15873 VDAC_N.n32 VDAC_N.n31 0.180667
R15874 VDAC_N.n31 VDAC_N.n30 0.180667
R15875 VDAC_N.n30 VDAC_N.n29 0.180667
R15876 VDAC_N.n29 VDAC_N.n28 0.180667
R15877 VDAC_N.n28 VDAC_N.n27 0.180667
R15878 VDAC_N.n27 VDAC_N.n26 0.180667
R15879 VDAC_N.n26 VDAC_N.n25 0.180667
R15880 VDAC_N.n25 VDAC_N.n24 0.180667
R15881 VDAC_N.n2134 VDAC_N.n23 0.180667
R15882 VDAC_N.n1973 VDAC_N.n1972 0.180667
R15883 VDAC_N.n1974 VDAC_N.n1973 0.180667
R15884 VDAC_N.n1975 VDAC_N.n1974 0.180667
R15885 VDAC_N.n1976 VDAC_N.n1975 0.180667
R15886 VDAC_N.n1977 VDAC_N.n1976 0.180667
R15887 VDAC_N.n1978 VDAC_N.n1977 0.180667
R15888 VDAC_N.n1979 VDAC_N.n1978 0.180667
R15889 VDAC_N.n1980 VDAC_N.n1979 0.180667
R15890 VDAC_N.n1981 VDAC_N.n1980 0.180667
R15891 VDAC_N.n1982 VDAC_N.n1981 0.180667
R15892 VDAC_N.n1983 VDAC_N.n1982 0.180667
R15893 VDAC_N.n1984 VDAC_N.n1983 0.180667
R15894 VDAC_N.n1985 VDAC_N.n1984 0.180667
R15895 VDAC_N.n1986 VDAC_N.n1985 0.180667
R15896 VDAC_N.n1987 VDAC_N.n1986 0.180667
R15897 VDAC_N.n1988 VDAC_N.n1987 0.180667
R15898 VDAC_N.n1989 VDAC_N.n1988 0.180667
R15899 VDAC_N.n1990 VDAC_N.n1989 0.180667
R15900 VDAC_N.n1991 VDAC_N.n1990 0.180667
R15901 VDAC_N.n1992 VDAC_N.n1991 0.180667
R15902 VDAC_N.n1993 VDAC_N.n1992 0.180667
R15903 VDAC_N.n1994 VDAC_N.n1993 0.180667
R15904 VDAC_N.n1995 VDAC_N.n1994 0.180667
R15905 VDAC_N.n1996 VDAC_N.n1995 0.180667
R15906 VDAC_N.n1997 VDAC_N.n1996 0.180667
R15907 VDAC_N.n1998 VDAC_N.n1997 0.180667
R15908 VDAC_N.n1999 VDAC_N.n1998 0.180667
R15909 VDAC_N.n2000 VDAC_N.n1999 0.180667
R15910 VDAC_N.n2001 VDAC_N.n2000 0.180667
R15911 VDAC_N.n2002 VDAC_N.n2001 0.180667
R15912 VDAC_N.n2003 VDAC_N.n2002 0.180667
R15913 VDAC_N.n2004 VDAC_N.n2003 0.180667
R15914 VDAC_N.n2005 VDAC_N.n2004 0.180667
R15915 VDAC_N.n2006 VDAC_N.n2005 0.180667
R15916 VDAC_N.n2007 VDAC_N.n2006 0.180667
R15917 VDAC_N.n2008 VDAC_N.n2007 0.180667
R15918 VDAC_N.n2009 VDAC_N.n2008 0.180667
R15919 VDAC_N.n2010 VDAC_N.n2009 0.180667
R15920 VDAC_N.n2011 VDAC_N.n2010 0.180667
R15921 VDAC_N.n2012 VDAC_N.n2011 0.180667
R15922 VDAC_N.n2013 VDAC_N.n2012 0.180667
R15923 VDAC_N.n2014 VDAC_N.n2013 0.180667
R15924 VDAC_N.n2015 VDAC_N.n2014 0.180667
R15925 VDAC_N.n2016 VDAC_N.n2015 0.180667
R15926 VDAC_N.n2017 VDAC_N.n2016 0.180667
R15927 VDAC_N.n2018 VDAC_N.n2017 0.180667
R15928 VDAC_N.n2019 VDAC_N.n2018 0.180667
R15929 VDAC_N.n2020 VDAC_N.n2019 0.180667
R15930 VDAC_N.n2021 VDAC_N.n2020 0.180667
R15931 VDAC_N.n2022 VDAC_N.n2021 0.180667
R15932 VDAC_N.n2023 VDAC_N.n2022 0.180667
R15933 VDAC_N.n2024 VDAC_N.n2023 0.180667
R15934 VDAC_N.n2025 VDAC_N.n2024 0.180667
R15935 VDAC_N.n2026 VDAC_N.n2025 0.180667
R15936 VDAC_N.n2027 VDAC_N.n2026 0.180667
R15937 VDAC_N.n2028 VDAC_N.n2027 0.180667
R15938 VDAC_N.n2029 VDAC_N.n2028 0.180667
R15939 VDAC_N.n2030 VDAC_N.n2029 0.180667
R15940 VDAC_N.n2031 VDAC_N.n2030 0.180667
R15941 VDAC_N.n2032 VDAC_N.n2031 0.180667
R15942 VDAC_N.n2033 VDAC_N.n2032 0.180667
R15943 VDAC_N.n2034 VDAC_N.n2033 0.180667
R15944 VDAC_N.n2035 VDAC_N.n2034 0.180667
R15945 VDAC_N.n2036 VDAC_N.n2035 0.180667
R15946 VDAC_N.n2037 VDAC_N.n2036 0.180667
R15947 VDAC_N.n2038 VDAC_N.n2037 0.180667
R15948 VDAC_N.n2039 VDAC_N.n2038 0.180667
R15949 VDAC_N.n2069 VDAC_N.n2068 0.180667
R15950 VDAC_N.n2070 VDAC_N.n2069 0.180667
R15951 VDAC_N.n2071 VDAC_N.n2070 0.180667
R15952 VDAC_N.n2072 VDAC_N.n2071 0.180667
R15953 VDAC_N.n2073 VDAC_N.n2072 0.180667
R15954 VDAC_N.n2074 VDAC_N.n2073 0.180667
R15955 VDAC_N.n2075 VDAC_N.n2074 0.180667
R15956 VDAC_N.n2076 VDAC_N.n2075 0.180667
R15957 VDAC_N.n2077 VDAC_N.n2076 0.180667
R15958 VDAC_N.n2078 VDAC_N.n2077 0.180667
R15959 VDAC_N.n2079 VDAC_N.n2078 0.180667
R15960 VDAC_N.n2080 VDAC_N.n2079 0.180667
R15961 VDAC_N.n2081 VDAC_N.n2080 0.180667
R15962 VDAC_N.n2082 VDAC_N.n2081 0.180667
R15963 VDAC_N.n2083 VDAC_N.n2082 0.180667
R15964 VDAC_N.n2084 VDAC_N.n2083 0.180667
R15965 VDAC_N.n2085 VDAC_N.n2084 0.180667
R15966 VDAC_N.n2086 VDAC_N.n2085 0.180667
R15967 VDAC_N.n2087 VDAC_N.n2086 0.180667
R15968 VDAC_N.n2088 VDAC_N.n2087 0.180667
R15969 VDAC_N.n2089 VDAC_N.n2088 0.180667
R15970 VDAC_N.n2090 VDAC_N.n2089 0.180667
R15971 VDAC_N.n2091 VDAC_N.n2090 0.180667
R15972 VDAC_N.n2092 VDAC_N.n2091 0.180667
R15973 VDAC_N.n2093 VDAC_N.n2092 0.180667
R15974 VDAC_N.n2094 VDAC_N.n2093 0.180667
R15975 VDAC_N.n2095 VDAC_N.n2094 0.180667
R15976 VDAC_N.n2096 VDAC_N.n2095 0.180667
R15977 VDAC_N.n2097 VDAC_N.n2096 0.180667
R15978 VDAC_N.n2098 VDAC_N.n2097 0.180667
R15979 VDAC_N.n2099 VDAC_N.n2098 0.180667
R15980 VDAC_N.n2100 VDAC_N.n2099 0.180667
R15981 VDAC_N.n2101 VDAC_N.n2100 0.180667
R15982 VDAC_N.n2102 VDAC_N.n2101 0.180667
R15983 VDAC_N.n2103 VDAC_N.n2102 0.180667
R15984 VDAC_N.n2104 VDAC_N.n2103 0.180667
R15985 VDAC_N.n2105 VDAC_N.n2104 0.180667
R15986 VDAC_N.n2106 VDAC_N.n2105 0.180667
R15987 VDAC_N.n2107 VDAC_N.n2106 0.180667
R15988 VDAC_N.n2108 VDAC_N.n2107 0.180667
R15989 VDAC_N.n2109 VDAC_N.n2108 0.180667
R15990 VDAC_N.n2110 VDAC_N.n2109 0.180667
R15991 VDAC_N.n2111 VDAC_N.n2110 0.180667
R15992 VDAC_N.n2112 VDAC_N.n2111 0.180667
R15993 VDAC_N.n2113 VDAC_N.n2112 0.180667
R15994 VDAC_N.n2114 VDAC_N.n2113 0.180667
R15995 VDAC_N.n2115 VDAC_N.n2114 0.180667
R15996 VDAC_N.n2116 VDAC_N.n2115 0.180667
R15997 VDAC_N.n2117 VDAC_N.n2116 0.180667
R15998 VDAC_N.n2118 VDAC_N.n2117 0.180667
R15999 VDAC_N.n2119 VDAC_N.n2118 0.180667
R16000 VDAC_N.n2120 VDAC_N.n2119 0.180667
R16001 VDAC_N.n2121 VDAC_N.n2120 0.180667
R16002 VDAC_N.n2122 VDAC_N.n2121 0.180667
R16003 VDAC_N.n2123 VDAC_N.n2122 0.180667
R16004 VDAC_N.n2124 VDAC_N.n2123 0.180667
R16005 VDAC_N.n2125 VDAC_N.n2124 0.180667
R16006 VDAC_N.n2126 VDAC_N.n2125 0.180667
R16007 VDAC_N.n2127 VDAC_N.n2126 0.180667
R16008 VDAC_N.n2128 VDAC_N.n2127 0.180667
R16009 VDAC_N.n2129 VDAC_N.n2128 0.180667
R16010 VDAC_N.n2130 VDAC_N.n2129 0.180667
R16011 VDAC_N.n2131 VDAC_N.n2130 0.180667
R16012 VDAC_N.n2132 VDAC_N.n2131 0.180667
R16013 VDAC_N.n2133 VDAC_N.n2132 0.180667
R16014 VDAC_N.n2134 VDAC_N.n2133 0.180667
R16015 VDAC_N.n2039 VDAC_N.n116 0.157167
R16016 VDAC_N.n1972 VDAC_N.n179 0.157167
R16017 VDAC_N.n2040 VDAC_N.n115 0.157167
R16018 VDAC_N.n1971 VDAC_N.n242 0.157167
R16019 VDAC_N.n2041 VDAC_N.n114 0.157167
R16020 VDAC_N.n1970 VDAC_N.n305 0.157167
R16021 VDAC_N.n2042 VDAC_N.n113 0.157167
R16022 VDAC_N.n1969 VDAC_N.n368 0.157167
R16023 VDAC_N.n2043 VDAC_N.n112 0.157167
R16024 VDAC_N.n1968 VDAC_N.n431 0.157167
R16025 VDAC_N.n2044 VDAC_N.n111 0.157167
R16026 VDAC_N.n1967 VDAC_N.n494 0.157167
R16027 VDAC_N.n2045 VDAC_N.n110 0.157167
R16028 VDAC_N.n1966 VDAC_N.n557 0.157167
R16029 VDAC_N.n2046 VDAC_N.n109 0.157167
R16030 VDAC_N.n1965 VDAC_N.n620 0.157167
R16031 VDAC_N.n2047 VDAC_N.n108 0.157167
R16032 VDAC_N.n1964 VDAC_N.n683 0.157167
R16033 VDAC_N.n2048 VDAC_N.n107 0.157167
R16034 VDAC_N.n1963 VDAC_N.n746 0.157167
R16035 VDAC_N.n2049 VDAC_N.n106 0.157167
R16036 VDAC_N.n1962 VDAC_N.n809 0.157167
R16037 VDAC_N.n2050 VDAC_N.n105 0.157167
R16038 VDAC_N.n1961 VDAC_N.n872 0.157167
R16039 VDAC_N.n2051 VDAC_N.n104 0.157167
R16040 VDAC_N.n1960 VDAC_N.n935 0.157167
R16041 VDAC_N.n2052 VDAC_N.n103 0.157167
R16042 VDAC_N.n1959 VDAC_N.n998 0.157167
R16043 VDAC_N.n2053 VDAC_N.n102 0.157167
R16044 VDAC_N.n1958 VDAC_N.n1061 0.157167
R16045 VDAC_N.n2054 VDAC_N.n101 0.157167
R16046 VDAC_N.n1957 VDAC_N.n1124 0.157167
R16047 VDAC_N.n2055 VDAC_N.n100 0.157167
R16048 VDAC_N.n1956 VDAC_N.n1187 0.157167
R16049 VDAC_N.n2056 VDAC_N.n99 0.157167
R16050 VDAC_N.n1955 VDAC_N.n1250 0.157167
R16051 VDAC_N.n2057 VDAC_N.n98 0.157167
R16052 VDAC_N.n1954 VDAC_N.n1313 0.157167
R16053 VDAC_N.n2058 VDAC_N.n97 0.157167
R16054 VDAC_N.n1953 VDAC_N.n1376 0.157167
R16055 VDAC_N.n2059 VDAC_N.n96 0.157167
R16056 VDAC_N.n1952 VDAC_N.n1439 0.157167
R16057 VDAC_N.n2060 VDAC_N.n95 0.157167
R16058 VDAC_N.n1951 VDAC_N.n1502 0.157167
R16059 VDAC_N.n2061 VDAC_N.n94 0.157167
R16060 VDAC_N.n1950 VDAC_N.n1565 0.157167
R16061 VDAC_N.n2062 VDAC_N.n93 0.157167
R16062 VDAC_N.n1949 VDAC_N.n1628 0.157167
R16063 VDAC_N.n2063 VDAC_N.n92 0.157167
R16064 VDAC_N.n1948 VDAC_N.n1691 0.157167
R16065 VDAC_N.n2064 VDAC_N.n91 0.157167
R16066 VDAC_N.n1947 VDAC_N.n1754 0.157167
R16067 VDAC_N.n2065 VDAC_N.n90 0.157167
R16068 VDAC_N.n1946 VDAC_N.n1817 0.157167
R16069 VDAC_N.n2066 VDAC_N.n89 0.157167
R16070 VDAC_N.n1945 VDAC_N.n1880 0.157167
R16071 VDAC_N.n2067 VDAC_N.n88 0.157167
R16072 VDAC_N.n1944 VDAC_N.n1943 0.157167
R16073 VDAC_N.n2068 VDAC_N.n87 0.157167
R16074 VDAC_N.n24 VDAC_N.n23 0.157167
R16075 VDAC_N VDAC_N.n2134 0.071
R16076 C6_N_btm.n4 C6_N_btm.t0 97.811
R16077 C6_N_btm.n3 C6_N_btm.t1 68.0518
R16078 C6_N_btm C6_N_btm.n4 59.5317
R16079 C6_N_btm.n2 C6_N_btm.n0 45.0311
R16080 C6_N_btm.n2 C6_N_btm.n1 37.4635
R16081 C6_N_btm.n1 C6_N_btm.t73 9.9005
R16082 C6_N_btm.n1 C6_N_btm.t72 9.9005
R16083 C6_N_btm.n0 C6_N_btm.t71 9.9005
R16084 C6_N_btm.n0 C6_N_btm.t70 9.9005
R16085 C6_N_btm.n4 C6_N_btm.n3 8.0005
R16086 C6_N_btm C6_N_btm.n187 7.24425
R16087 C6_N_btm.n3 C6_N_btm.n2 6.58904
R16088 C6_N_btm.n39 C6_N_btm.t66 5.03712
R16089 C6_N_btm.n36 C6_N_btm.t67 5.03712
R16090 C6_N_btm.n183 C6_N_btm.t68 5.03712
R16091 C6_N_btm.n163 C6_N_btm.n162 4.60698
R16092 C6_N_btm.n162 C6_N_btm.n161 4.60698
R16093 C6_N_btm.n143 C6_N_btm.n142 4.60698
R16094 C6_N_btm.n144 C6_N_btm.n143 4.60698
R16095 C6_N_btm.n146 C6_N_btm.n145 4.60698
R16096 C6_N_btm.n147 C6_N_btm.n146 4.60698
R16097 C6_N_btm.n149 C6_N_btm.n148 4.60698
R16098 C6_N_btm.n150 C6_N_btm.n149 4.60698
R16099 C6_N_btm.n152 C6_N_btm.n151 4.60698
R16100 C6_N_btm.n151 C6_N_btm.n13 4.60698
R16101 C6_N_btm.n157 C6_N_btm.n156 4.60698
R16102 C6_N_btm.n156 C6_N_btm.n155 4.60698
R16103 C6_N_btm.n160 C6_N_btm.n159 4.60698
R16104 C6_N_btm.n159 C6_N_btm.n158 4.60698
R16105 C6_N_btm.n76 C6_N_btm.n75 4.60698
R16106 C6_N_btm.n77 C6_N_btm.n76 4.60698
R16107 C6_N_btm.n79 C6_N_btm.n78 4.60698
R16108 C6_N_btm.n80 C6_N_btm.n79 4.60698
R16109 C6_N_btm.n82 C6_N_btm.n81 4.60698
R16110 C6_N_btm.n83 C6_N_btm.n82 4.60698
R16111 C6_N_btm.n85 C6_N_btm.n84 4.60698
R16112 C6_N_btm.n86 C6_N_btm.n85 4.60698
R16113 C6_N_btm.n88 C6_N_btm.n87 4.60698
R16114 C6_N_btm.n89 C6_N_btm.n88 4.60698
R16115 C6_N_btm.n91 C6_N_btm.n90 4.60698
R16116 C6_N_btm.n92 C6_N_btm.n91 4.60698
R16117 C6_N_btm.n94 C6_N_btm.n93 4.60698
R16118 C6_N_btm.n95 C6_N_btm.n94 4.60698
R16119 C6_N_btm.n97 C6_N_btm.n96 4.60698
R16120 C6_N_btm.n98 C6_N_btm.n97 4.60698
R16121 C6_N_btm.n103 C6_N_btm.n102 4.60698
R16122 C6_N_btm.n104 C6_N_btm.n103 4.60698
R16123 C6_N_btm.n106 C6_N_btm.n105 4.60698
R16124 C6_N_btm.n107 C6_N_btm.n106 4.60698
R16125 C6_N_btm.n109 C6_N_btm.n108 4.60698
R16126 C6_N_btm.n110 C6_N_btm.n109 4.60698
R16127 C6_N_btm.n112 C6_N_btm.n111 4.60698
R16128 C6_N_btm.n113 C6_N_btm.n112 4.60698
R16129 C6_N_btm.n115 C6_N_btm.n114 4.60698
R16130 C6_N_btm.n116 C6_N_btm.n115 4.60698
R16131 C6_N_btm.n118 C6_N_btm.n117 4.60698
R16132 C6_N_btm.n119 C6_N_btm.n118 4.60698
R16133 C6_N_btm.n122 C6_N_btm.n121 4.60698
R16134 C6_N_btm.n121 C6_N_btm.n120 4.60698
R16135 C6_N_btm.n124 C6_N_btm.n123 4.60698
R16136 C6_N_btm.n125 C6_N_btm.n124 4.60698
R16137 C6_N_btm.n127 C6_N_btm.n126 4.60698
R16138 C6_N_btm.n128 C6_N_btm.n127 4.60698
R16139 C6_N_btm.n130 C6_N_btm.n129 4.60698
R16140 C6_N_btm.n131 C6_N_btm.n130 4.60698
R16141 C6_N_btm.n133 C6_N_btm.n132 4.60698
R16142 C6_N_btm.n134 C6_N_btm.n133 4.60698
R16143 C6_N_btm.n137 C6_N_btm.n135 4.60698
R16144 C6_N_btm.n138 C6_N_btm.n137 4.60698
R16145 C6_N_btm.n62 C6_N_btm.n61 4.60698
R16146 C6_N_btm.n61 C6_N_btm.n60 4.60698
R16147 C6_N_btm.n65 C6_N_btm.n64 4.60698
R16148 C6_N_btm.n64 C6_N_btm.n63 4.60698
R16149 C6_N_btm.n68 C6_N_btm.n67 4.60698
R16150 C6_N_btm.n67 C6_N_btm.n66 4.60698
R16151 C6_N_btm.n187 C6_N_btm.t69 4.03712
R16152 C6_N_btm.n185 C6_N_btm.t21 3.98193
R16153 C6_N_btm.n180 C6_N_btm.t47 3.98193
R16154 C6_N_btm.n177 C6_N_btm.t59 3.98193
R16155 C6_N_btm.n174 C6_N_btm.t63 3.98193
R16156 C6_N_btm.n171 C6_N_btm.t38 3.98193
R16157 C6_N_btm.n166 C6_N_btm.t44 3.98193
R16158 C6_N_btm.n154 C6_N_btm.t64 3.98193
R16159 C6_N_btm.n99 C6_N_btm.t30 3.98193
R16160 C6_N_btm.n101 C6_N_btm.t9 3.98193
R16161 C6_N_btm.n20 C6_N_btm.t12 3.98193
R16162 C6_N_btm.n21 C6_N_btm.t31 3.98193
R16163 C6_N_btm.n136 C6_N_btm.t2 3.98193
R16164 C6_N_btm.n59 C6_N_btm.t54 3.98193
R16165 C6_N_btm.n55 C6_N_btm.t48 3.98193
R16166 C6_N_btm.n52 C6_N_btm.t65 3.98193
R16167 C6_N_btm.n49 C6_N_btm.t37 3.98193
R16168 C6_N_btm.n44 C6_N_btm.t29 3.98193
R16169 C6_N_btm.n41 C6_N_btm.t57 3.98193
R16170 C6_N_btm.n38 C6_N_btm.t8 3.98193
R16171 C6_N_btm.n37 C6_N_btm.t50 3.98193
R16172 C6_N_btm.n42 C6_N_btm.t5 3.98193
R16173 C6_N_btm.n45 C6_N_btm.t26 3.98193
R16174 C6_N_btm.n48 C6_N_btm.t61 3.98193
R16175 C6_N_btm.n51 C6_N_btm.t53 3.98193
R16176 C6_N_btm.n56 C6_N_btm.t22 3.98193
R16177 C6_N_btm.n69 C6_N_btm.t36 3.98193
R16178 C6_N_btm.n141 C6_N_btm.t7 3.98193
R16179 C6_N_btm.n164 C6_N_btm.t60 3.98193
R16180 C6_N_btm.n167 C6_N_btm.t23 3.98193
R16181 C6_N_btm.n170 C6_N_btm.t17 3.98193
R16182 C6_N_btm.n173 C6_N_btm.t10 3.98193
R16183 C6_N_btm.n178 C6_N_btm.t35 3.98193
R16184 C6_N_btm.n181 C6_N_btm.t58 3.98193
R16185 C6_N_btm.n184 C6_N_btm.t55 3.98193
R16186 C6_N_btm.n162 C6_N_btm.t20 1.67819
R16187 C6_N_btm.n143 C6_N_btm.t56 1.67819
R16188 C6_N_btm.n146 C6_N_btm.t41 1.67819
R16189 C6_N_btm.n149 C6_N_btm.t19 1.67819
R16190 C6_N_btm.n151 C6_N_btm.t39 1.67819
R16191 C6_N_btm.n156 C6_N_btm.t51 1.67819
R16192 C6_N_btm.n159 C6_N_btm.t34 1.67819
R16193 C6_N_btm.n76 C6_N_btm.t15 1.67819
R16194 C6_N_btm.n79 C6_N_btm.t62 1.67819
R16195 C6_N_btm.n82 C6_N_btm.t4 1.67819
R16196 C6_N_btm.n85 C6_N_btm.t49 1.67819
R16197 C6_N_btm.n88 C6_N_btm.t42 1.67819
R16198 C6_N_btm.n91 C6_N_btm.t11 1.67819
R16199 C6_N_btm.n94 C6_N_btm.t40 1.67819
R16200 C6_N_btm.n97 C6_N_btm.t3 1.67819
R16201 C6_N_btm.n103 C6_N_btm.t27 1.67819
R16202 C6_N_btm.n106 C6_N_btm.t14 1.67819
R16203 C6_N_btm.n109 C6_N_btm.t33 1.67819
R16204 C6_N_btm.n112 C6_N_btm.t18 1.67819
R16205 C6_N_btm.n115 C6_N_btm.t52 1.67819
R16206 C6_N_btm.n118 C6_N_btm.t25 1.67819
R16207 C6_N_btm.n121 C6_N_btm.t6 1.67819
R16208 C6_N_btm.n124 C6_N_btm.t28 1.67819
R16209 C6_N_btm.n127 C6_N_btm.t13 1.67819
R16210 C6_N_btm.n130 C6_N_btm.t45 1.67819
R16211 C6_N_btm.n133 C6_N_btm.t16 1.67819
R16212 C6_N_btm.n137 C6_N_btm.t43 1.67819
R16213 C6_N_btm.n61 C6_N_btm.t46 1.67819
R16214 C6_N_btm.n64 C6_N_btm.t32 1.67819
R16215 C6_N_btm.n67 C6_N_btm.t24 1.67819
R16216 C6_N_btm.n154 C6_N_btm.n153 1.05569
R16217 C6_N_btm.n22 C6_N_btm.n21 1.05569
R16218 C6_N_btm.n20 C6_N_btm.n19 1.05569
R16219 C6_N_btm.n136 C6_N_btm.n8 1.05569
R16220 C6_N_btm.n101 C6_N_btm.n100 1.05569
R16221 C6_N_btm.n70 C6_N_btm.n69 1.05569
R16222 C6_N_btm.n140 C6_N_btm.n9 1.0005
R16223 C6_N_btm.n14 C6_N_btm.n11 1.0005
R16224 C6_N_btm.n15 C6_N_btm.n10 1.0005
R16225 C6_N_btm.n29 C6_N_btm.n27 1.0005
R16226 C6_N_btm.n30 C6_N_btm.n26 1.0005
R16227 C6_N_btm.n31 C6_N_btm.n25 1.0005
R16228 C6_N_btm.n70 C6_N_btm.n24 1.0005
R16229 C6_N_btm.n71 C6_N_btm.n23 1.0005
R16230 C6_N_btm.n72 C6_N_btm.n22 1.0005
R16231 C6_N_btm.n73 C6_N_btm.n19 1.0005
R16232 C6_N_btm.n74 C6_N_btm.n18 1.0005
R16233 C6_N_btm.n153 C6_N_btm.n12 1.0005
R16234 C6_N_btm.n17 C6_N_btm.n14 1.0005
R16235 C6_N_btm.n16 C6_N_btm.n15 1.0005
R16236 C6_N_btm.n140 C6_N_btm.n139 1.0005
R16237 C6_N_btm.n43 C6_N_btm.n36 1.0005
R16238 C6_N_btm.n40 C6_N_btm.n39 1.0005
R16239 C6_N_btm.n40 C6_N_btm.n35 1.0005
R16240 C6_N_btm.n46 C6_N_btm.n43 1.0005
R16241 C6_N_btm.n47 C6_N_btm.n46 1.0005
R16242 C6_N_btm.n50 C6_N_btm.n35 1.0005
R16243 C6_N_btm.n53 C6_N_btm.n50 1.0005
R16244 C6_N_btm.n47 C6_N_btm.n34 1.0005
R16245 C6_N_btm.n57 C6_N_btm.n34 1.0005
R16246 C6_N_btm.n54 C6_N_btm.n53 1.0005
R16247 C6_N_btm.n54 C6_N_btm.n28 1.0005
R16248 C6_N_btm.n58 C6_N_btm.n57 1.0005
R16249 C6_N_btm.n58 C6_N_btm.n29 1.0005
R16250 C6_N_btm.n33 C6_N_btm.n30 1.0005
R16251 C6_N_btm.n32 C6_N_btm.n31 1.0005
R16252 C6_N_btm.n100 C6_N_btm.n28 1.0005
R16253 C6_N_btm.n168 C6_N_btm.n165 1.0005
R16254 C6_N_btm.n165 C6_N_btm.n8 1.0005
R16255 C6_N_btm.n172 C6_N_btm.n7 1.0005
R16256 C6_N_btm.n9 C6_N_btm.n7 1.0005
R16257 C6_N_btm.n169 C6_N_btm.n6 1.0005
R16258 C6_N_btm.n169 C6_N_btm.n168 1.0005
R16259 C6_N_btm.n176 C6_N_btm.n175 1.0005
R16260 C6_N_btm.n175 C6_N_btm.n172 1.0005
R16261 C6_N_btm.n182 C6_N_btm.n179 1.0005
R16262 C6_N_btm.n179 C6_N_btm.n6 1.0005
R16263 C6_N_btm.n186 C6_N_btm.n5 1.0005
R16264 C6_N_btm.n176 C6_N_btm.n5 1.0005
R16265 C6_N_btm.n183 C6_N_btm.n182 1.0005
R16266 C6_N_btm.n187 C6_N_btm.n186 1.0005
R16267 C6_N_btm.n21 C6_N_btm.n20 0.733338
R16268 C6_N_btm.n38 C6_N_btm.n37 0.733338
R16269 C6_N_btm.n42 C6_N_btm.n41 0.733338
R16270 C6_N_btm.n45 C6_N_btm.n44 0.733338
R16271 C6_N_btm.n49 C6_N_btm.n48 0.733338
R16272 C6_N_btm.n52 C6_N_btm.n51 0.733338
R16273 C6_N_btm.n56 C6_N_btm.n55 0.733338
R16274 C6_N_btm.n167 C6_N_btm.n166 0.733338
R16275 C6_N_btm.n171 C6_N_btm.n170 0.733338
R16276 C6_N_btm.n174 C6_N_btm.n173 0.733338
R16277 C6_N_btm.n178 C6_N_btm.n177 0.733338
R16278 C6_N_btm.n181 C6_N_btm.n180 0.733338
R16279 C6_N_btm.n185 C6_N_btm.n184 0.733338
R16280 C6_N_btm.n155 C6_N_btm.n154 0.679419
R16281 C6_N_btm.n138 C6_N_btm.n136 0.679419
R16282 C6_N_btm.n102 C6_N_btm.n101 0.679419
R16283 C6_N_btm.n69 C6_N_btm.n68 0.679419
R16284 C6_N_btm.n60 C6_N_btm.n59 0.679419
R16285 C6_N_btm.n99 C6_N_btm.n98 0.679419
R16286 C6_N_btm.n142 C6_N_btm.n141 0.679419
R16287 C6_N_btm.n164 C6_N_btm.n163 0.679419
R16288 C6_N_btm.n161 C6_N_btm.n160 0.6255
R16289 C6_N_btm.n158 C6_N_btm.n157 0.6255
R16290 C6_N_btm.n135 C6_N_btm.n134 0.6255
R16291 C6_N_btm.n132 C6_N_btm.n131 0.6255
R16292 C6_N_btm.n129 C6_N_btm.n128 0.6255
R16293 C6_N_btm.n126 C6_N_btm.n125 0.6255
R16294 C6_N_btm.n123 C6_N_btm.n122 0.6255
R16295 C6_N_btm.n120 C6_N_btm.n119 0.6255
R16296 C6_N_btm.n117 C6_N_btm.n116 0.6255
R16297 C6_N_btm.n114 C6_N_btm.n113 0.6255
R16298 C6_N_btm.n111 C6_N_btm.n110 0.6255
R16299 C6_N_btm.n108 C6_N_btm.n107 0.6255
R16300 C6_N_btm.n105 C6_N_btm.n104 0.6255
R16301 C6_N_btm.n66 C6_N_btm.n65 0.6255
R16302 C6_N_btm.n63 C6_N_btm.n62 0.6255
R16303 C6_N_btm.n96 C6_N_btm.n95 0.6255
R16304 C6_N_btm.n93 C6_N_btm.n92 0.6255
R16305 C6_N_btm.n90 C6_N_btm.n89 0.6255
R16306 C6_N_btm.n87 C6_N_btm.n86 0.6255
R16307 C6_N_btm.n84 C6_N_btm.n83 0.6255
R16308 C6_N_btm.n81 C6_N_btm.n80 0.6255
R16309 C6_N_btm.n78 C6_N_btm.n77 0.6255
R16310 C6_N_btm.n75 C6_N_btm.n13 0.6255
R16311 C6_N_btm.n152 C6_N_btm.n150 0.6255
R16312 C6_N_btm.n148 C6_N_btm.n147 0.6255
R16313 C6_N_btm.n145 C6_N_btm.n144 0.6255
R16314 C6_N_btm.n158 C6_N_btm.n10 0.109875
R16315 C6_N_btm.n160 C6_N_btm.n10 0.109875
R16316 C6_N_btm.n155 C6_N_btm.n11 0.109875
R16317 C6_N_btm.n157 C6_N_btm.n11 0.109875
R16318 C6_N_btm.n139 C6_N_btm.n135 0.109875
R16319 C6_N_btm.n139 C6_N_btm.n138 0.109875
R16320 C6_N_btm.n132 C6_N_btm.n16 0.109875
R16321 C6_N_btm.n134 C6_N_btm.n16 0.109875
R16322 C6_N_btm.n129 C6_N_btm.n17 0.109875
R16323 C6_N_btm.n131 C6_N_btm.n17 0.109875
R16324 C6_N_btm.n126 C6_N_btm.n12 0.109875
R16325 C6_N_btm.n128 C6_N_btm.n12 0.109875
R16326 C6_N_btm.n123 C6_N_btm.n18 0.109875
R16327 C6_N_btm.n125 C6_N_btm.n18 0.109875
R16328 C6_N_btm.n120 C6_N_btm.n19 0.109875
R16329 C6_N_btm.n122 C6_N_btm.n19 0.109875
R16330 C6_N_btm.n117 C6_N_btm.n22 0.109875
R16331 C6_N_btm.n119 C6_N_btm.n22 0.109875
R16332 C6_N_btm.n114 C6_N_btm.n23 0.109875
R16333 C6_N_btm.n116 C6_N_btm.n23 0.109875
R16334 C6_N_btm.n111 C6_N_btm.n24 0.109875
R16335 C6_N_btm.n113 C6_N_btm.n24 0.109875
R16336 C6_N_btm.n108 C6_N_btm.n25 0.109875
R16337 C6_N_btm.n110 C6_N_btm.n25 0.109875
R16338 C6_N_btm.n105 C6_N_btm.n26 0.109875
R16339 C6_N_btm.n107 C6_N_btm.n26 0.109875
R16340 C6_N_btm.n102 C6_N_btm.n27 0.109875
R16341 C6_N_btm.n104 C6_N_btm.n27 0.109875
R16342 C6_N_btm.n66 C6_N_btm.n32 0.109875
R16343 C6_N_btm.n68 C6_N_btm.n32 0.109875
R16344 C6_N_btm.n63 C6_N_btm.n33 0.109875
R16345 C6_N_btm.n65 C6_N_btm.n33 0.109875
R16346 C6_N_btm.n60 C6_N_btm.n58 0.109875
R16347 C6_N_btm.n62 C6_N_btm.n58 0.109875
R16348 C6_N_btm.n98 C6_N_btm.n29 0.109875
R16349 C6_N_btm.n96 C6_N_btm.n29 0.109875
R16350 C6_N_btm.n95 C6_N_btm.n30 0.109875
R16351 C6_N_btm.n93 C6_N_btm.n30 0.109875
R16352 C6_N_btm.n92 C6_N_btm.n31 0.109875
R16353 C6_N_btm.n90 C6_N_btm.n31 0.109875
R16354 C6_N_btm.n89 C6_N_btm.n70 0.109875
R16355 C6_N_btm.n87 C6_N_btm.n70 0.109875
R16356 C6_N_btm.n86 C6_N_btm.n71 0.109875
R16357 C6_N_btm.n84 C6_N_btm.n71 0.109875
R16358 C6_N_btm.n83 C6_N_btm.n72 0.109875
R16359 C6_N_btm.n81 C6_N_btm.n72 0.109875
R16360 C6_N_btm.n80 C6_N_btm.n73 0.109875
R16361 C6_N_btm.n78 C6_N_btm.n73 0.109875
R16362 C6_N_btm.n77 C6_N_btm.n74 0.109875
R16363 C6_N_btm.n75 C6_N_btm.n74 0.109875
R16364 C6_N_btm.n153 C6_N_btm.n13 0.109875
R16365 C6_N_btm.n153 C6_N_btm.n152 0.109875
R16366 C6_N_btm.n150 C6_N_btm.n14 0.109875
R16367 C6_N_btm.n148 C6_N_btm.n14 0.109875
R16368 C6_N_btm.n147 C6_N_btm.n15 0.109875
R16369 C6_N_btm.n145 C6_N_btm.n15 0.109875
R16370 C6_N_btm.n144 C6_N_btm.n140 0.109875
R16371 C6_N_btm.n142 C6_N_btm.n140 0.109875
R16372 C6_N_btm.n161 C6_N_btm.n9 0.109875
R16373 C6_N_btm.n163 C6_N_btm.n9 0.109875
R16374 C6_N_btm.n37 C6_N_btm.n36 0.0556875
R16375 C6_N_btm.n39 C6_N_btm.n38 0.0556875
R16376 C6_N_btm.n41 C6_N_btm.n40 0.0556875
R16377 C6_N_btm.n43 C6_N_btm.n42 0.0556875
R16378 C6_N_btm.n46 C6_N_btm.n45 0.0556875
R16379 C6_N_btm.n44 C6_N_btm.n35 0.0556875
R16380 C6_N_btm.n50 C6_N_btm.n49 0.0556875
R16381 C6_N_btm.n48 C6_N_btm.n47 0.0556875
R16382 C6_N_btm.n51 C6_N_btm.n34 0.0556875
R16383 C6_N_btm.n53 C6_N_btm.n52 0.0556875
R16384 C6_N_btm.n55 C6_N_btm.n54 0.0556875
R16385 C6_N_btm.n57 C6_N_btm.n56 0.0556875
R16386 C6_N_btm.n59 C6_N_btm.n28 0.0556875
R16387 C6_N_btm.n100 C6_N_btm.n99 0.0556875
R16388 C6_N_btm.n141 C6_N_btm.n8 0.0556875
R16389 C6_N_btm.n165 C6_N_btm.n164 0.0556875
R16390 C6_N_btm.n166 C6_N_btm.n7 0.0556875
R16391 C6_N_btm.n168 C6_N_btm.n167 0.0556875
R16392 C6_N_btm.n170 C6_N_btm.n169 0.0556875
R16393 C6_N_btm.n172 C6_N_btm.n171 0.0556875
R16394 C6_N_btm.n175 C6_N_btm.n174 0.0556875
R16395 C6_N_btm.n173 C6_N_btm.n6 0.0556875
R16396 C6_N_btm.n179 C6_N_btm.n178 0.0556875
R16397 C6_N_btm.n177 C6_N_btm.n176 0.0556875
R16398 C6_N_btm.n180 C6_N_btm.n5 0.0556875
R16399 C6_N_btm.n182 C6_N_btm.n181 0.0556875
R16400 C6_N_btm.n184 C6_N_btm.n183 0.0556875
R16401 C6_N_btm.n186 C6_N_btm.n185 0.0556875
R16402 VDAC_P.n3 VDAC_P.t320 946.489
R16403 VDAC_P.n0 VDAC_P.t1085 946.489
R16404 VDAC_P.n7 VDAC_P.t602 946.345
R16405 VDAC_P.n13 VDAC_P.t941 945.764
R16406 VDAC_P.n12 VDAC_P.t165 945.755
R16407 VDAC_P.n11 VDAC_P.t1087 945.755
R16408 VDAC_P.n10 VDAC_P.t2078 945.755
R16409 VDAC_P.n9 VDAC_P.t221 945.755
R16410 VDAC_P.n8 VDAC_P.t1081 945.755
R16411 VDAC_P.n7 VDAC_P.t668 945.755
R16412 VDAC_P.n5 VDAC_P.t1537 945.755
R16413 VDAC_P.n4 VDAC_P.t2091 945.755
R16414 VDAC_P.n3 VDAC_P.t2131 945.755
R16415 VDAC_P.n2 VDAC_P.t456 945.755
R16416 VDAC_P.n1 VDAC_P.t90 945.755
R16417 VDAC_P.n0 VDAC_P.t1050 945.755
R16418 VDAC_P.n20 VDAC_P.n18 14.894
R16419 VDAC_P.n17 VDAC_P.n15 14.894
R16420 VDAC_P.n17 VDAC_P.n16 14.394
R16421 VDAC_P.n20 VDAC_P.n19 14.394
R16422 VDAC_P.n22 VDAC_P.n14 13.701
R16423 VDAC_P.n22 VDAC_P.n21 13.3496
R16424 VDAC_P.n10 VDAC_P.n9 6.67373
R16425 VDAC_P.n6 VDAC_P.n2 6.20847
R16426 VDAC_P.n14 VDAC_P.n6 5.45883
R16427 VDAC_P.n14 VDAC_P.n13 4.5005
R16428 VDAC_P.n16 VDAC_P.t3 2.4755
R16429 VDAC_P.n16 VDAC_P.t2 2.4755
R16430 VDAC_P.n19 VDAC_P.t4 2.4755
R16431 VDAC_P.n19 VDAC_P.t6 2.4755
R16432 VDAC_P.n18 VDAC_P.t7 2.4755
R16433 VDAC_P.n18 VDAC_P.t5 2.4755
R16434 VDAC_P.n15 VDAC_P.t1 2.4755
R16435 VDAC_P.n15 VDAC_P.t0 2.4755
R16436 VDAC_P VDAC_P.n22 2.28
R16437 VDAC_P.n116 VDAC_P.t87 1.1255
R16438 VDAC_P.n117 VDAC_P.t1251 1.1255
R16439 VDAC_P.n118 VDAC_P.t919 1.1255
R16440 VDAC_P.n119 VDAC_P.t1147 1.1255
R16441 VDAC_P.n120 VDAC_P.t421 1.1255
R16442 VDAC_P.n121 VDAC_P.t1041 1.1255
R16443 VDAC_P.n122 VDAC_P.t761 1.1255
R16444 VDAC_P.n123 VDAC_P.t43 1.1255
R16445 VDAC_P.n124 VDAC_P.t2020 1.1255
R16446 VDAC_P.n125 VDAC_P.t933 1.1255
R16447 VDAC_P.n126 VDAC_P.t164 1.1255
R16448 VDAC_P.n127 VDAC_P.t1631 1.1255
R16449 VDAC_P.n128 VDAC_P.t2134 1.1255
R16450 VDAC_P.n129 VDAC_P.t152 1.1255
R16451 VDAC_P.n130 VDAC_P.t1074 1.1255
R16452 VDAC_P.n131 VDAC_P.t480 1.1255
R16453 VDAC_P.n132 VDAC_P.t1046 1.1255
R16454 VDAC_P.n133 VDAC_P.t704 1.1255
R16455 VDAC_P.n134 VDAC_P.t430 1.1255
R16456 VDAC_P.n135 VDAC_P.t713 1.1255
R16457 VDAC_P.n136 VDAC_P.t202 1.1255
R16458 VDAC_P.n137 VDAC_P.t1191 1.1255
R16459 VDAC_P.n138 VDAC_P.t614 1.1255
R16460 VDAC_P.n139 VDAC_P.t19 1.1255
R16461 VDAC_P.n140 VDAC_P.t785 1.1255
R16462 VDAC_P.n141 VDAC_P.t862 1.1255
R16463 VDAC_P.n142 VDAC_P.t1429 1.1255
R16464 VDAC_P.n143 VDAC_P.t1889 1.1255
R16465 VDAC_P.n144 VDAC_P.t103 1.1255
R16466 VDAC_P.n145 VDAC_P.t467 1.1255
R16467 VDAC_P.n146 VDAC_P.t571 1.1255
R16468 VDAC_P.n147 VDAC_P.t1573 1.1255
R16469 VDAC_P.n148 VDAC_P.t2115 1.1255
R16470 VDAC_P.n149 VDAC_P.t747 1.1255
R16471 VDAC_P.n150 VDAC_P.t1917 1.1255
R16472 VDAC_P.n151 VDAC_P.t1828 1.1255
R16473 VDAC_P.n152 VDAC_P.t1811 1.1255
R16474 VDAC_P.n153 VDAC_P.t908 1.1255
R16475 VDAC_P.n154 VDAC_P.t1601 1.1255
R16476 VDAC_P.n155 VDAC_P.t1436 1.1255
R16477 VDAC_P.n156 VDAC_P.t1904 1.1255
R16478 VDAC_P.n157 VDAC_P.t279 1.1255
R16479 VDAC_P.n158 VDAC_P.t1808 1.1255
R16480 VDAC_P.n159 VDAC_P.t1850 1.1255
R16481 VDAC_P.n160 VDAC_P.t1860 1.1255
R16482 VDAC_P.n161 VDAC_P.t1410 1.1255
R16483 VDAC_P.n162 VDAC_P.t107 1.1255
R16484 VDAC_P.n163 VDAC_P.t174 1.1255
R16485 VDAC_P.n164 VDAC_P.t11 1.1255
R16486 VDAC_P.n165 VDAC_P.t1920 1.1255
R16487 VDAC_P.n166 VDAC_P.t970 1.1255
R16488 VDAC_P.n167 VDAC_P.t727 1.1255
R16489 VDAC_P.n168 VDAC_P.t1682 1.1255
R16490 VDAC_P.n169 VDAC_P.t353 1.1255
R16491 VDAC_P.n170 VDAC_P.t903 1.1255
R16492 VDAC_P.n171 VDAC_P.t569 1.1255
R16493 VDAC_P.n172 VDAC_P.t1679 1.1255
R16494 VDAC_P.n173 VDAC_P.t998 1.1255
R16495 VDAC_P.n174 VDAC_P.t1463 1.1255
R16496 VDAC_P.n175 VDAC_P.t2025 1.1255
R16497 VDAC_P.n176 VDAC_P.t1357 1.1255
R16498 VDAC_P.n177 VDAC_P.t473 1.1255
R16499 VDAC_P.n178 VDAC_P.t1764 1.1255
R16500 VDAC_P.n179 VDAC_P.t447 1.1255
R16501 VDAC_P.n115 VDAC_P.t591 1.1255
R16502 VDAC_P.n180 VDAC_P.t1800 1.1255
R16503 VDAC_P.n181 VDAC_P.t1038 1.1255
R16504 VDAC_P.n182 VDAC_P.t1344 1.1255
R16505 VDAC_P.n183 VDAC_P.t1622 1.1255
R16506 VDAC_P.n184 VDAC_P.t657 1.1255
R16507 VDAC_P.n185 VDAC_P.t1398 1.1255
R16508 VDAC_P.n186 VDAC_P.t317 1.1255
R16509 VDAC_P.n187 VDAC_P.t1639 1.1255
R16510 VDAC_P.n188 VDAC_P.t158 1.1255
R16511 VDAC_P.n189 VDAC_P.t1529 1.1255
R16512 VDAC_P.n190 VDAC_P.t234 1.1255
R16513 VDAC_P.n191 VDAC_P.t1419 1.1255
R16514 VDAC_P.n192 VDAC_P.t1873 1.1255
R16515 VDAC_P.n193 VDAC_P.t1953 1.1255
R16516 VDAC_P.n194 VDAC_P.t1060 1.1255
R16517 VDAC_P.n195 VDAC_P.t442 1.1255
R16518 VDAC_P.n196 VDAC_P.t1188 1.1255
R16519 VDAC_P.n197 VDAC_P.t1258 1.1255
R16520 VDAC_P.n198 VDAC_P.t625 1.1255
R16521 VDAC_P.n199 VDAC_P.t1040 1.1255
R16522 VDAC_P.n200 VDAC_P.t1970 1.1255
R16523 VDAC_P.n201 VDAC_P.t1624 1.1255
R16524 VDAC_P.n202 VDAC_P.t1750 1.1255
R16525 VDAC_P.n203 VDAC_P.t693 1.1255
R16526 VDAC_P.n204 VDAC_P.t1318 1.1255
R16527 VDAC_P.n205 VDAC_P.t333 1.1255
R16528 VDAC_P.n206 VDAC_P.t1705 1.1255
R16529 VDAC_P.n207 VDAC_P.t2034 1.1255
R16530 VDAC_P.n208 VDAC_P.t77 1.1255
R16531 VDAC_P.n209 VDAC_P.t1810 1.1255
R16532 VDAC_P.n210 VDAC_P.t197 1.1255
R16533 VDAC_P.n211 VDAC_P.t985 1.1255
R16534 VDAC_P.n212 VDAC_P.t339 1.1255
R16535 VDAC_P.n213 VDAC_P.t1729 1.1255
R16536 VDAC_P.n214 VDAC_P.t92 1.1255
R16537 VDAC_P.n215 VDAC_P.t1623 1.1255
R16538 VDAC_P.n216 VDAC_P.t2081 1.1255
R16539 VDAC_P.n217 VDAC_P.t1405 1.1255
R16540 VDAC_P.n218 VDAC_P.t1001 1.1255
R16541 VDAC_P.n219 VDAC_P.t1128 1.1255
R16542 VDAC_P.n220 VDAC_P.t1841 1.1255
R16543 VDAC_P.n221 VDAC_P.t1028 1.1255
R16544 VDAC_P.n222 VDAC_P.t390 1.1255
R16545 VDAC_P.n223 VDAC_P.t316 1.1255
R16546 VDAC_P.n224 VDAC_P.t1032 1.1255
R16547 VDAC_P.n225 VDAC_P.t1101 1.1255
R16548 VDAC_P.n226 VDAC_P.t424 1.1255
R16549 VDAC_P.n227 VDAC_P.t886 1.1255
R16550 VDAC_P.n228 VDAC_P.t584 1.1255
R16551 VDAC_P.n229 VDAC_P.t1538 1.1255
R16552 VDAC_P.n230 VDAC_P.t637 1.1255
R16553 VDAC_P.n231 VDAC_P.t346 1.1255
R16554 VDAC_P.n232 VDAC_P.t1139 1.1255
R16555 VDAC_P.n233 VDAC_P.t1591 1.1255
R16556 VDAC_P.n234 VDAC_P.t1802 1.1255
R16557 VDAC_P.n235 VDAC_P.t757 1.1255
R16558 VDAC_P.n236 VDAC_P.t222 1.1255
R16559 VDAC_P.n237 VDAC_P.t1269 1.1255
R16560 VDAC_P.n238 VDAC_P.t253 1.1255
R16561 VDAC_P.n239 VDAC_P.t1167 1.1255
R16562 VDAC_P.n240 VDAC_P.t1621 1.1255
R16563 VDAC_P.n241 VDAC_P.t540 1.1255
R16564 VDAC_P.n242 VDAC_P.t771 1.1255
R16565 VDAC_P.n114 VDAC_P.t1376 1.1255
R16566 VDAC_P.n243 VDAC_P.t35 1.1255
R16567 VDAC_P.n244 VDAC_P.t948 1.1255
R16568 VDAC_P.n245 VDAC_P.t1713 1.1255
R16569 VDAC_P.n246 VDAC_P.t22 1.1255
R16570 VDAC_P.n247 VDAC_P.t1936 1.1255
R16571 VDAC_P.n248 VDAC_P.t1045 1.1255
R16572 VDAC_P.n249 VDAC_P.t400 1.1255
R16573 VDAC_P.n250 VDAC_P.t1694 1.1255
R16574 VDAC_P.n251 VDAC_P.t2116 1.1255
R16575 VDAC_P.n252 VDAC_P.t1490 1.1255
R16576 VDAC_P.n253 VDAC_P.t1340 1.1255
R16577 VDAC_P.n254 VDAC_P.t1262 1.1255
R16578 VDAC_P.n255 VDAC_P.t1113 1.1255
R16579 VDAC_P.n256 VDAC_P.t1763 1.1255
R16580 VDAC_P.n257 VDAC_P.t2108 1.1255
R16581 VDAC_P.n258 VDAC_P.t1302 1.1255
R16582 VDAC_P.n259 VDAC_P.t2113 1.1255
R16583 VDAC_P.n260 VDAC_P.t1736 1.1255
R16584 VDAC_P.n261 VDAC_P.t2010 1.1255
R16585 VDAC_P.n262 VDAC_P.t1256 1.1255
R16586 VDAC_P.n263 VDAC_P.t1582 1.1255
R16587 VDAC_P.n264 VDAC_P.t1636 1.1255
R16588 VDAC_P.n265 VDAC_P.t1354 1.1255
R16589 VDAC_P.n266 VDAC_P.t313 1.1255
R16590 VDAC_P.n267 VDAC_P.t1840 1.1255
R16591 VDAC_P.n268 VDAC_P.t2066 1.1255
R16592 VDAC_P.n269 VDAC_P.t1515 1.1255
R16593 VDAC_P.n270 VDAC_P.t1638 1.1255
R16594 VDAC_P.n271 VDAC_P.t1399 1.1255
R16595 VDAC_P.n272 VDAC_P.t1422 1.1255
R16596 VDAC_P.n273 VDAC_P.t319 1.1255
R16597 VDAC_P.n274 VDAC_P.t889 1.1255
R16598 VDAC_P.n275 VDAC_P.t21 1.1255
R16599 VDAC_P.n276 VDAC_P.t1543 1.1255
R16600 VDAC_P.n277 VDAC_P.t521 1.1255
R16601 VDAC_P.n278 VDAC_P.t729 1.1255
R16602 VDAC_P.n279 VDAC_P.t959 1.1255
R16603 VDAC_P.n280 VDAC_P.t1229 1.1255
R16604 VDAC_P.n281 VDAC_P.t1785 1.1255
R16605 VDAC_P.n282 VDAC_P.t1292 1.1255
R16606 VDAC_P.n283 VDAC_P.t841 1.1255
R16607 VDAC_P.n284 VDAC_P.t1852 1.1255
R16608 VDAC_P.n285 VDAC_P.t1080 1.1255
R16609 VDAC_P.n286 VDAC_P.t2005 1.1255
R16610 VDAC_P.n287 VDAC_P.t632 1.1255
R16611 VDAC_P.n288 VDAC_P.t1786 1.1255
R16612 VDAC_P.n289 VDAC_P.t1588 1.1255
R16613 VDAC_P.n290 VDAC_P.t1350 1.1255
R16614 VDAC_P.n291 VDAC_P.t364 1.1255
R16615 VDAC_P.n292 VDAC_P.t582 1.1255
R16616 VDAC_P.n293 VDAC_P.t282 1.1255
R16617 VDAC_P.n294 VDAC_P.t920 1.1255
R16618 VDAC_P.n295 VDAC_P.t142 1.1255
R16619 VDAC_P.n296 VDAC_P.t1395 1.1255
R16620 VDAC_P.n297 VDAC_P.t374 1.1255
R16621 VDAC_P.n298 VDAC_P.t661 1.1255
R16622 VDAC_P.n299 VDAC_P.t1198 1.1255
R16623 VDAC_P.n300 VDAC_P.t13 1.1255
R16624 VDAC_P.n301 VDAC_P.t129 1.1255
R16625 VDAC_P.n302 VDAC_P.t1914 1.1255
R16626 VDAC_P.n303 VDAC_P.t1427 1.1255
R16627 VDAC_P.n304 VDAC_P.t519 1.1255
R16628 VDAC_P.n305 VDAC_P.t1329 1.1255
R16629 VDAC_P.n113 VDAC_P.t211 1.1255
R16630 VDAC_P.n306 VDAC_P.t1590 1.1255
R16631 VDAC_P.n307 VDAC_P.t1379 1.1255
R16632 VDAC_P.n308 VDAC_P.t1370 1.1255
R16633 VDAC_P.n309 VDAC_P.t1171 1.1255
R16634 VDAC_P.n310 VDAC_P.t827 1.1255
R16635 VDAC_P.n311 VDAC_P.t30 1.1255
R16636 VDAC_P.n312 VDAC_P.t401 1.1255
R16637 VDAC_P.n313 VDAC_P.t1977 1.1255
R16638 VDAC_P.n314 VDAC_P.t71 1.1255
R16639 VDAC_P.n315 VDAC_P.t1861 1.1255
R16640 VDAC_P.n316 VDAC_P.t613 1.1255
R16641 VDAC_P.n317 VDAC_P.t1757 1.1255
R16642 VDAC_P.n318 VDAC_P.t252 1.1255
R16643 VDAC_P.n319 VDAC_P.t672 1.1255
R16644 VDAC_P.n320 VDAC_P.t1610 1.1255
R16645 VDAC_P.n321 VDAC_P.t367 1.1255
R16646 VDAC_P.n322 VDAC_P.t706 1.1255
R16647 VDAC_P.n323 VDAC_P.t1179 1.1255
R16648 VDAC_P.n324 VDAC_P.t1735 1.1255
R16649 VDAC_P.n325 VDAC_P.t1062 1.1255
R16650 VDAC_P.n326 VDAC_P.t777 1.1255
R16651 VDAC_P.n327 VDAC_P.t86 1.1255
R16652 VDAC_P.n328 VDAC_P.t201 1.1255
R16653 VDAC_P.n329 VDAC_P.t949 1.1255
R16654 VDAC_P.n330 VDAC_P.t1209 1.1255
R16655 VDAC_P.n331 VDAC_P.t245 1.1255
R16656 VDAC_P.n332 VDAC_P.t556 1.1255
R16657 VDAC_P.n333 VDAC_P.t1561 1.1255
R16658 VDAC_P.n334 VDAC_P.t289 1.1255
R16659 VDAC_P.n335 VDAC_P.t383 1.1255
R16660 VDAC_P.n336 VDAC_P.t965 1.1255
R16661 VDAC_P.n337 VDAC_P.t336 1.1255
R16662 VDAC_P.n338 VDAC_P.t1797 1.1255
R16663 VDAC_P.n339 VDAC_P.t1484 1.1255
R16664 VDAC_P.n340 VDAC_P.t1158 1.1255
R16665 VDAC_P.n341 VDAC_P.t2122 1.1255
R16666 VDAC_P.n342 VDAC_P.t1848 1.1255
R16667 VDAC_P.n343 VDAC_P.t1929 1.1255
R16668 VDAC_P.n344 VDAC_P.t368 1.1255
R16669 VDAC_P.n345 VDAC_P.t834 1.1255
R16670 VDAC_P.n346 VDAC_P.t868 1.1255
R16671 VDAC_P.n347 VDAC_P.t1594 1.1255
R16672 VDAC_P.n348 VDAC_P.t1277 1.1255
R16673 VDAC_P.n349 VDAC_P.t170 1.1255
R16674 VDAC_P.n350 VDAC_P.t2082 1.1255
R16675 VDAC_P.n351 VDAC_P.t1629 1.1255
R16676 VDAC_P.n352 VDAC_P.t490 1.1255
R16677 VDAC_P.n353 VDAC_P.t1407 1.1255
R16678 VDAC_P.n354 VDAC_P.t1650 1.1255
R16679 VDAC_P.n355 VDAC_P.t1309 1.1255
R16680 VDAC_P.n356 VDAC_P.t1761 1.1255
R16681 VDAC_P.n357 VDAC_P.t1201 1.1255
R16682 VDAC_P.n358 VDAC_P.t843 1.1255
R16683 VDAC_P.n359 VDAC_P.t2111 1.1255
R16684 VDAC_P.n360 VDAC_P.t735 1.1255
R16685 VDAC_P.n361 VDAC_P.t523 1.1255
R16686 VDAC_P.n362 VDAC_P.t1339 1.1255
R16687 VDAC_P.n363 VDAC_P.t911 1.1255
R16688 VDAC_P.n364 VDAC_P.t1620 1.1255
R16689 VDAC_P.n365 VDAC_P.t859 1.1255
R16690 VDAC_P.n366 VDAC_P.t550 1.1255
R16691 VDAC_P.n367 VDAC_P.t1142 1.1255
R16692 VDAC_P.n368 VDAC_P.t2037 1.1255
R16693 VDAC_P.n112 VDAC_P.t198 1.1255
R16694 VDAC_P.n369 VDAC_P.t412 1.1255
R16695 VDAC_P.n370 VDAC_P.t1174 1.1255
R16696 VDAC_P.n371 VDAC_P.t2051 1.1255
R16697 VDAC_P.n372 VDAC_P.t744 1.1255
R16698 VDAC_P.n373 VDAC_P.t1666 1.1255
R16699 VDAC_P.n374 VDAC_P.t276 1.1255
R16700 VDAC_P.n375 VDAC_P.t1462 1.1255
R16701 VDAC_P.n376 VDAC_P.t1211 1.1255
R16702 VDAC_P.n377 VDAC_P.t634 1.1255
R16703 VDAC_P.n378 VDAC_P.t1095 1.1255
R16704 VDAC_P.n379 VDAC_P.t1584 1.1255
R16705 VDAC_P.n380 VDAC_P.t58 1.1255
R16706 VDAC_P.n381 VDAC_P.t739 1.1255
R16707 VDAC_P.n382 VDAC_P.t1036 1.1255
R16708 VDAC_P.n383 VDAC_P.t626 1.1255
R16709 VDAC_P.n384 VDAC_P.t615 1.1255
R16710 VDAC_P.n385 VDAC_P.t1984 1.1255
R16711 VDAC_P.n386 VDAC_P.t982 1.1255
R16712 VDAC_P.n387 VDAC_P.t1553 1.1255
R16713 VDAC_P.n388 VDAC_P.t1714 1.1255
R16714 VDAC_P.n389 VDAC_P.t69 1.1255
R16715 VDAC_P.n390 VDAC_P.t398 1.1255
R16716 VDAC_P.n391 VDAC_P.t631 1.1255
R16717 VDAC_P.n392 VDAC_P.t1691 1.1255
R16718 VDAC_P.n393 VDAC_P.t1010 1.1255
R16719 VDAC_P.n394 VDAC_P.t803 1.1255
R16720 VDAC_P.n395 VDAC_P.t1033 1.1255
R16721 VDAC_P.n396 VDAC_P.t363 1.1255
R16722 VDAC_P.n397 VDAC_P.t265 1.1255
R16723 VDAC_P.n398 VDAC_P.t105 1.1255
R16724 VDAC_P.n399 VDAC_P.t449 1.1255
R16725 VDAC_P.n400 VDAC_P.t1868 1.1255
R16726 VDAC_P.n401 VDAC_P.t1609 1.1255
R16727 VDAC_P.n402 VDAC_P.t2061 1.1255
R16728 VDAC_P.n403 VDAC_P.t768 1.1255
R16729 VDAC_P.n404 VDAC_P.t991 1.1255
R16730 VDAC_P.n405 VDAC_P.t548 1.1255
R16731 VDAC_P.n406 VDAC_P.t1743 1.1255
R16732 VDAC_P.n407 VDAC_P.t612 1.1255
R16733 VDAC_P.n408 VDAC_P.t182 1.1255
R16734 VDAC_P.n409 VDAC_P.t1308 1.1255
R16735 VDAC_P.n410 VDAC_P.t618 1.1255
R16736 VDAC_P.n411 VDAC_P.t1083 1.1255
R16737 VDAC_P.n412 VDAC_P.t1528 1.1255
R16738 VDAC_P.n413 VDAC_P.t1698 1.1255
R16739 VDAC_P.n414 VDAC_P.t731 1.1255
R16740 VDAC_P.n415 VDAC_P.t762 1.1255
R16741 VDAC_P.n416 VDAC_P.t629 1.1255
R16742 VDAC_P.n417 VDAC_P.t338 1.1255
R16743 VDAC_P.n418 VDAC_P.t45 1.1255
R16744 VDAC_P.n419 VDAC_P.t1575 1.1255
R16745 VDAC_P.n420 VDAC_P.t1974 1.1255
R16746 VDAC_P.n421 VDAC_P.t1469 1.1255
R16747 VDAC_P.n422 VDAC_P.t1921 1.1255
R16748 VDAC_P.n423 VDAC_P.t1255 1.1255
R16749 VDAC_P.n424 VDAC_P.t921 1.1255
R16750 VDAC_P.n425 VDAC_P.t309 1.1255
R16751 VDAC_P.n426 VDAC_P.t817 1.1255
R16752 VDAC_P.n427 VDAC_P.t1820 1.1255
R16753 VDAC_P.n428 VDAC_P.t51 1.1255
R16754 VDAC_P.n429 VDAC_P.t509 1.1255
R16755 VDAC_P.n430 VDAC_P.t1480 1.1255
R16756 VDAC_P.n431 VDAC_P.t1843 1.1255
R16757 VDAC_P.n111 VDAC_P.t925 1.1255
R16758 VDAC_P.n432 VDAC_P.t1157 1.1255
R16759 VDAC_P.n433 VDAC_P.t871 1.1255
R16760 VDAC_P.n434 VDAC_P.t534 1.1255
R16761 VDAC_P.n435 VDAC_P.t1507 1.1255
R16762 VDAC_P.n436 VDAC_P.t993 1.1255
R16763 VDAC_P.n437 VDAC_P.t1389 1.1255
R16764 VDAC_P.n438 VDAC_P.t1849 1.1255
R16765 VDAC_P.n439 VDAC_P.t1220 1.1255
R16766 VDAC_P.n440 VDAC_P.t457 1.1255
R16767 VDAC_P.n441 VDAC_P.t700 1.1255
R16768 VDAC_P.n442 VDAC_P.t1531 1.1255
R16769 VDAC_P.n443 VDAC_P.t1059 1.1255
R16770 VDAC_P.n444 VDAC_P.t1648 1.1255
R16771 VDAC_P.n445 VDAC_P.t458 1.1255
R16772 VDAC_P.n446 VDAC_P.t1353 1.1255
R16773 VDAC_P.n447 VDAC_P.t1911 1.1255
R16774 VDAC_P.n448 VDAC_P.t1247 1.1255
R16775 VDAC_P.n449 VDAC_P.t1701 1.1255
R16776 VDAC_P.n450 VDAC_P.t1612 1.1255
R16777 VDAC_P.n451 VDAC_P.t1593 1.1255
R16778 VDAC_P.n452 VDAC_P.t2047 1.1255
R16779 VDAC_P.n453 VDAC_P.t393 1.1255
R16780 VDAC_P.n454 VDAC_P.t267 1.1255
R16781 VDAC_P.n455 VDAC_P.t516 1.1255
R16782 VDAC_P.n456 VDAC_P.t453 1.1255
R16783 VDAC_P.n457 VDAC_P.t44 1.1255
R16784 VDAC_P.n458 VDAC_P.t1230 1.1255
R16785 VDAC_P.n459 VDAC_P.t1053 1.1255
R16786 VDAC_P.n460 VDAC_P.t1008 1.1255
R16787 VDAC_P.n461 VDAC_P.t1973 1.1255
R16788 VDAC_P.n462 VDAC_P.t576 1.1255
R16789 VDAC_P.n463 VDAC_P.t1718 1.1255
R16790 VDAC_P.n464 VDAC_P.t356 1.1255
R16791 VDAC_P.n465 VDAC_P.t1290 1.1255
R16792 VDAC_P.n466 VDAC_P.t1129 1.1255
R16793 VDAC_P.n467 VDAC_P.t2112 1.1255
R16794 VDAC_P.n468 VDAC_P.t1014 1.1255
R16795 VDAC_P.n469 VDAC_P.t1224 1.1255
R16796 VDAC_P.n470 VDAC_P.t1774 1.1255
R16797 VDAC_P.n471 VDAC_P.t699 1.1255
R16798 VDAC_P.n472 VDAC_P.t782 1.1255
R16799 VDAC_P.n473 VDAC_P.t1345 1.1255
R16800 VDAC_P.n474 VDAC_P.t1801 1.1255
R16801 VDAC_P.n475 VDAC_P.t583 1.1255
R16802 VDAC_P.n476 VDAC_P.t1587 1.1255
R16803 VDAC_P.n477 VDAC_P.t1500 1.1255
R16804 VDAC_P.n478 VDAC_P.t755 1.1255
R16805 VDAC_P.n479 VDAC_P.t505 1.1255
R16806 VDAC_P.n480 VDAC_P.t49 1.1255
R16807 VDAC_P.n481 VDAC_P.t1825 1.1255
R16808 VDAC_P.n482 VDAC_P.t1996 1.1255
R16809 VDAC_P.n483 VDAC_P.t873 1.1255
R16810 VDAC_P.n484 VDAC_P.t24 1.1255
R16811 VDAC_P.n485 VDAC_P.t1968 1.1255
R16812 VDAC_P.n486 VDAC_P.t1967 1.1255
R16813 VDAC_P.n487 VDAC_P.t216 1.1255
R16814 VDAC_P.n488 VDAC_P.t1855 1.1255
R16815 VDAC_P.n489 VDAC_P.t1300 1.1255
R16816 VDAC_P.n490 VDAC_P.t74 1.1255
R16817 VDAC_P.n491 VDAC_P.t828 1.1255
R16818 VDAC_P.n492 VDAC_P.t2096 1.1255
R16819 VDAC_P.n493 VDAC_P.t573 1.1255
R16820 VDAC_P.n494 VDAC_P.t440 1.1255
R16821 VDAC_P.n110 VDAC_P.t538 1.1255
R16822 VDAC_P.n495 VDAC_P.t1384 1.1255
R16823 VDAC_P.n496 VDAC_P.t1858 1.1255
R16824 VDAC_P.n497 VDAC_P.t1892 1.1255
R16825 VDAC_P.n498 VDAC_P.t726 1.1255
R16826 VDAC_P.n499 VDAC_P.t1193 1.1255
R16827 VDAC_P.n500 VDAC_P.t322 1.1255
R16828 VDAC_P.n501 VDAC_P.t23 1.1255
R16829 VDAC_P.n502 VDAC_P.t1545 1.1255
R16830 VDAC_P.n503 VDAC_P.t974 1.1255
R16831 VDAC_P.n504 VDAC_P.t1431 1.1255
R16832 VDAC_P.n505 VDAC_P.t394 1.1255
R16833 VDAC_P.n506 VDAC_P.t191 1.1255
R16834 VDAC_P.n507 VDAC_P.t907 1.1255
R16835 VDAC_P.n508 VDAC_P.t690 1.1255
R16836 VDAC_P.n509 VDAC_P.t1165 1.1255
R16837 VDAC_P.n510 VDAC_P.t1719 1.1255
R16838 VDAC_P.n511 VDAC_P.t2062 1.1255
R16839 VDAC_P.n512 VDAC_P.t1513 1.1255
R16840 VDAC_P.n513 VDAC_P.t1047 1.1255
R16841 VDAC_P.n514 VDAC_P.t1397 1.1255
R16842 VDAC_P.n515 VDAC_P.t485 1.1255
R16843 VDAC_P.n516 VDAC_P.t1297 1.1255
R16844 VDAC_P.n517 VDAC_P.t1749 1.1255
R16845 VDAC_P.n518 VDAC_P.t1660 1.1255
R16846 VDAC_P.n519 VDAC_P.t1541 1.1255
R16847 VDAC_P.n520 VDAC_P.t545 1.1255
R16848 VDAC_P.n521 VDAC_P.t1680 1.1255
R16849 VDAC_P.n522 VDAC_P.t493 1.1255
R16850 VDAC_P.n523 VDAC_P.t1200 1.1255
R16851 VDAC_P.n524 VDAC_P.t1783 1.1255
R16852 VDAC_P.n525 VDAC_P.t652 1.1255
R16853 VDAC_P.n526 VDAC_P.t354 1.1255
R16854 VDAC_P.n527 VDAC_P.t2106 1.1255
R16855 VDAC_P.n528 VDAC_P.t1792 1.1255
R16856 VDAC_P.n529 VDAC_P.t1834 1.1255
R16857 VDAC_P.n530 VDAC_P.t352 1.1255
R16858 VDAC_P.n531 VDAC_P.t1618 1.1255
R16859 VDAC_P.n532 VDAC_P.t1772 1.1255
R16860 VDAC_P.n533 VDAC_P.t1390 1.1255
R16861 VDAC_P.n534 VDAC_P.t605 1.1255
R16862 VDAC_P.n535 VDAC_P.t166 1.1255
R16863 VDAC_P.n536 VDAC_P.t1159 1.1255
R16864 VDAC_P.n537 VDAC_P.t821 1.1255
R16865 VDAC_P.n538 VDAC_P.t938 1.1255
R16866 VDAC_P.n539 VDAC_P.t369 1.1255
R16867 VDAC_P.n540 VDAC_P.t1959 1.1255
R16868 VDAC_P.n541 VDAC_P.t1291 1.1255
R16869 VDAC_P.n542 VDAC_P.t1747 1.1255
R16870 VDAC_P.n543 VDAC_P.t607 1.1255
R16871 VDAC_P.n544 VDAC_P.t1643 1.1255
R16872 VDAC_P.n545 VDAC_P.t1061 1.1255
R16873 VDAC_P.n546 VDAC_P.t75 1.1255
R16874 VDAC_P.n547 VDAC_P.t1991 1.1255
R16875 VDAC_P.n548 VDAC_P.t64 1.1255
R16876 VDAC_P.n549 VDAC_P.t465 1.1255
R16877 VDAC_P.n550 VDAC_P.t1476 1.1255
R16878 VDAC_P.n551 VDAC_P.t1677 1.1255
R16879 VDAC_P.n552 VDAC_P.t1079 1.1255
R16880 VDAC_P.n553 VDAC_P.t566 1.1255
R16881 VDAC_P.n554 VDAC_P.t2023 1.1255
R16882 VDAC_P.n555 VDAC_P.t1312 1.1255
R16883 VDAC_P.n556 VDAC_P.t1814 1.1255
R16884 VDAC_P.n557 VDAC_P.t1748 1.1255
R16885 VDAC_P.n109 VDAC_P.t1972 1.1255
R16886 VDAC_P.n558 VDAC_P.t1727 1.1255
R16887 VDAC_P.n559 VDAC_P.t2060 1.1255
R16888 VDAC_P.n560 VDAC_P.t825 1.1255
R16889 VDAC_P.n561 VDAC_P.t2077 1.1255
R16890 VDAC_P.n562 VDAC_P.t40 1.1255
R16891 VDAC_P.n563 VDAC_P.t271 1.1255
R16892 VDAC_P.n564 VDAC_P.t96 1.1255
R16893 VDAC_P.n565 VDAC_P.t1518 1.1255
R16894 VDAC_P.n566 VDAC_P.t1332 1.1255
R16895 VDAC_P.n567 VDAC_P.t1286 1.1255
R16896 VDAC_P.n568 VDAC_P.t2103 1.1255
R16897 VDAC_P.n569 VDAC_P.t288 1.1255
R16898 VDAC_P.n570 VDAC_P.t274 1.1255
R16899 VDAC_P.n571 VDAC_P.t264 1.1255
R16900 VDAC_P.n572 VDAC_P.t1910 1.1255
R16901 VDAC_P.n573 VDAC_P.t1533 1.1255
R16902 VDAC_P.n574 VDAC_P.t854 1.1255
R16903 VDAC_P.n575 VDAC_P.t1327 1.1255
R16904 VDAC_P.n576 VDAC_P.t259 1.1255
R16905 VDAC_P.n577 VDAC_P.t1221 1.1255
R16906 VDAC_P.n578 VDAC_P.t853 1.1255
R16907 VDAC_P.n579 VDAC_P.t297 1.1255
R16908 VDAC_P.n580 VDAC_P.t797 1.1255
R16909 VDAC_P.n581 VDAC_P.t527 1.1255
R16910 VDAC_P.n582 VDAC_P.t1355 1.1255
R16911 VDAC_P.n583 VDAC_P.t499 1.1255
R16912 VDAC_P.n584 VDAC_P.t244 1.1255
R16913 VDAC_P.n585 VDAC_P.t1703 1.1255
R16914 VDAC_P.n586 VDAC_P.t428 1.1255
R16915 VDAC_P.n587 VDAC_P.t1595 1.1255
R16916 VDAC_P.n588 VDAC_P.t2049 1.1255
R16917 VDAC_P.n589 VDAC_P.t488 1.1255
R16918 VDAC_P.n590 VDAC_P.t1941 1.1255
R16919 VDAC_P.n591 VDAC_P.t1012 1.1255
R16920 VDAC_P.n592 VDAC_P.t1454 1.1255
R16921 VDAC_P.n593 VDAC_P.t2092 1.1255
R16922 VDAC_P.n594 VDAC_P.t1234 1.1255
R16923 VDAC_P.n595 VDAC_P.t541 1.1255
R16924 VDAC_P.n596 VDAC_P.t1992 1.1255
R16925 VDAC_P.n597 VDAC_P.t1942 1.1255
R16926 VDAC_P.n598 VDAC_P.t752 1.1255
R16927 VDAC_P.n599 VDAC_P.t962 1.1255
R16928 VDAC_P.n600 VDAC_P.t115 1.1255
R16929 VDAC_P.n601 VDAC_P.t1474 1.1255
R16930 VDAC_P.n602 VDAC_P.t1217 1.1255
R16931 VDAC_P.n603 VDAC_P.t463 1.1255
R16932 VDAC_P.n604 VDAC_P.t1099 1.1255
R16933 VDAC_P.n605 VDAC_P.t1563 1.1255
R16934 VDAC_P.n606 VDAC_P.t510 1.1255
R16935 VDAC_P.n607 VDAC_P.t1455 1.1255
R16936 VDAC_P.n608 VDAC_P.t1907 1.1255
R16937 VDAC_P.n609 VDAC_P.t687 1.1255
R16938 VDAC_P.n610 VDAC_P.t915 1.1255
R16939 VDAC_P.n611 VDAC_P.t76 1.1255
R16940 VDAC_P.n612 VDAC_P.t223 1.1255
R16941 VDAC_P.n613 VDAC_P.t732 1.1255
R16942 VDAC_P.n614 VDAC_P.t1485 1.1255
R16943 VDAC_P.n615 VDAC_P.t1937 1.1255
R16944 VDAC_P.n616 VDAC_P.t200 1.1255
R16945 VDAC_P.n617 VDAC_P.t1827 1.1255
R16946 VDAC_P.n618 VDAC_P.t2028 1.1255
R16947 VDAC_P.n619 VDAC_P.t50 1.1255
R16948 VDAC_P.n620 VDAC_P.t1884 1.1255
R16949 VDAC_P.n108 VDAC_P.t1581 1.1255
R16950 VDAC_P.n621 VDAC_P.t906 1.1255
R16951 VDAC_P.n622 VDAC_P.t1477 1.1255
R16952 VDAC_P.n623 VDAC_P.t1570 1.1255
R16953 VDAC_P.n624 VDAC_P.t337 1.1255
R16954 VDAC_P.n625 VDAC_P.t239 1.1255
R16955 VDAC_P.n626 VDAC_P.t311 1.1255
R16956 VDAC_P.n627 VDAC_P.t1615 1.1255
R16957 VDAC_P.n628 VDAC_P.t537 1.1255
R16958 VDAC_P.n629 VDAC_P.t213 1.1255
R16959 VDAC_P.n630 VDAC_P.t511 1.1255
R16960 VDAC_P.n631 VDAC_P.t1293 1.1255
R16961 VDAC_P.n632 VDAC_P.t939 1.1255
R16962 VDAC_P.n633 VDAC_P.t628 1.1255
R16963 VDAC_P.n634 VDAC_P.t609 1.1255
R16964 VDAC_P.n635 VDAC_P.t839 1.1255
R16965 VDAC_P.n636 VDAC_P.t1596 1.1255
R16966 VDAC_P.n637 VDAC_P.t217 1.1255
R16967 VDAC_P.n638 VDAC_P.t1013 1.1255
R16968 VDAC_P.n639 VDAC_P.t1672 1.1255
R16969 VDAC_P.n640 VDAC_P.t1887 1.1255
R16970 VDAC_P.n641 VDAC_P.t404 1.1255
R16971 VDAC_P.n642 VDAC_P.t905 1.1255
R16972 VDAC_P.n643 VDAC_P.t1260 1.1255
R16973 VDAC_P.n644 VDAC_P.t1122 1.1255
R16974 VDAC_P.n645 VDAC_P.t1029 1.1255
R16975 VDAC_P.n646 VDAC_P.t248 1.1255
R16976 VDAC_P.n647 VDAC_P.t930 1.1255
R16977 VDAC_P.n648 VDAC_P.t84 1.1255
R16978 VDAC_P.n649 VDAC_P.t822 1.1255
R16979 VDAC_P.n650 VDAC_P.t460 1.1255
R16980 VDAC_P.n651 VDAC_P.t1182 1.1255
R16981 VDAC_P.n652 VDAC_P.t1181 1.1255
R16982 VDAC_P.n653 VDAC_P.t496 1.1255
R16983 VDAC_P.n654 VDAC_P.t1894 1.1255
R16984 VDAC_P.n655 VDAC_P.t723 1.1255
R16985 VDAC_P.n656 VDAC_P.t438 1.1255
R16986 VDAC_P.n657 VDAC_P.t1319 1.1255
R16987 VDAC_P.n658 VDAC_P.t66 1.1255
R16988 VDAC_P.n659 VDAC_P.t1213 1.1255
R16989 VDAC_P.n660 VDAC_P.t233 1.1255
R16990 VDAC_P.n661 VDAC_P.t10 1.1255
R16991 VDAC_P.n662 VDAC_P.t835 1.1255
R16992 VDAC_P.n663 VDAC_P.t2093 1.1255
R16993 VDAC_P.n664 VDAC_P.t377 1.1255
R16994 VDAC_P.n665 VDAC_P.t491 1.1255
R16995 VDAC_P.n666 VDAC_P.t600 1.1255
R16996 VDAC_P.n667 VDAC_P.t901 1.1255
R16997 VDAC_P.n668 VDAC_P.t1164 1.1255
R16998 VDAC_P.n669 VDAC_P.t131 1.1255
R16999 VDAC_P.n670 VDAC_P.t553 1.1255
R17000 VDAC_P.n671 VDAC_P.t464 1.1255
R17001 VDAC_P.n672 VDAC_P.t277 1.1255
R17002 VDAC_P.n673 VDAC_P.t1304 1.1255
R17003 VDAC_P.n674 VDAC_P.t1606 1.1255
R17004 VDAC_P.n675 VDAC_P.t1676 1.1255
R17005 VDAC_P.n676 VDAC_P.t1378 1.1255
R17006 VDAC_P.n677 VDAC_P.t1116 1.1255
R17007 VDAC_P.n678 VDAC_P.t144 1.1255
R17008 VDAC_P.n679 VDAC_P.t286 1.1255
R17009 VDAC_P.n680 VDAC_P.t72 1.1255
R17010 VDAC_P.n681 VDAC_P.t130 1.1255
R17011 VDAC_P.n682 VDAC_P.t719 1.1255
R17012 VDAC_P.n683 VDAC_P.t738 1.1255
R17013 VDAC_P.n107 VDAC_P.t418 1.1255
R17014 VDAC_P.n684 VDAC_P.t1516 1.1255
R17015 VDAC_P.n685 VDAC_P.t1366 1.1255
R17016 VDAC_P.n686 VDAC_P.t1628 1.1255
R17017 VDAC_P.n687 VDAC_P.t1856 1.1255
R17018 VDAC_P.n688 VDAC_P.t258 1.1255
R17019 VDAC_P.n689 VDAC_P.t1400 1.1255
R17020 VDAC_P.n690 VDAC_P.t230 1.1255
R17021 VDAC_P.n691 VDAC_P.t1303 1.1255
R17022 VDAC_P.n692 VDAC_P.t1434 1.1255
R17023 VDAC_P.n693 VDAC_P.t101 1.1255
R17024 VDAC_P.n694 VDAC_P.t88 1.1255
R17025 VDAC_P.n695 VDAC_P.t555 1.1255
R17026 VDAC_P.n696 VDAC_P.t1547 1.1255
R17027 VDAC_P.n697 VDAC_P.t270 1.1255
R17028 VDAC_P.n698 VDAC_P.t207 1.1255
R17029 VDAC_P.n699 VDAC_P.t1025 1.1255
R17030 VDAC_P.n700 VDAC_P.t691 1.1255
R17031 VDAC_P.n701 VDAC_P.t1805 1.1255
R17032 VDAC_P.n702 VDAC_P.t884 1.1255
R17033 VDAC_P.n703 VDAC_P.t865 1.1255
R17034 VDAC_P.n704 VDAC_P.t156 1.1255
R17035 VDAC_P.n705 VDAC_P.t811 1.1255
R17036 VDAC_P.n706 VDAC_P.t533 1.1255
R17037 VDAC_P.n707 VDAC_P.t736 1.1255
R17038 VDAC_P.n708 VDAC_P.t931 1.1255
R17039 VDAC_P.n709 VDAC_P.t1988 1.1255
R17040 VDAC_P.n710 VDAC_P.t206 1.1255
R17041 VDAC_P.n711 VDAC_P.t2012 1.1255
R17042 VDAC_P.n712 VDAC_P.t630 1.1255
R17043 VDAC_P.n713 VDAC_P.t2079 1.1255
R17044 VDAC_P.n714 VDAC_P.t1568 1.1255
R17045 VDAC_P.n715 VDAC_P.t506 1.1255
R17046 VDAC_P.n716 VDAC_P.t1120 1.1255
R17047 VDAC_P.n717 VDAC_P.t774 1.1255
R17048 VDAC_P.n718 VDAC_P.t1239 1.1255
R17049 VDAC_P.n719 VDAC_P.t658 1.1255
R17050 VDAC_P.n720 VDAC_P.t303 1.1255
R17051 VDAC_P.n721 VDAC_P.t448 1.1255
R17052 VDAC_P.n722 VDAC_P.t1998 1.1255
R17053 VDAC_P.n723 VDAC_P.t209 1.1255
R17054 VDAC_P.n724 VDAC_P.t242 1.1255
R17055 VDAC_P.n725 VDAC_P.t741 1.1255
R17056 VDAC_P.n726 VDAC_P.t967 1.1255
R17057 VDAC_P.n727 VDAC_P.t47 1.1255
R17058 VDAC_P.n728 VDAC_P.t1697 1.1255
R17059 VDAC_P.n729 VDAC_P.t1548 1.1255
R17060 VDAC_P.n730 VDAC_P.t807 1.1255
R17061 VDAC_P.n731 VDAC_P.t91 1.1255
R17062 VDAC_P.n732 VDAC_P.t119 1.1255
R17063 VDAC_P.n733 VDAC_P.t1935 1.1255
R17064 VDAC_P.n734 VDAC_P.t148 1.1255
R17065 VDAC_P.n735 VDAC_P.t927 1.1255
R17066 VDAC_P.n736 VDAC_P.t524 1.1255
R17067 VDAC_P.n737 VDAC_P.t326 1.1255
R17068 VDAC_P.n738 VDAC_P.t539 1.1255
R17069 VDAC_P.n739 VDAC_P.t1000 1.1255
R17070 VDAC_P.n740 VDAC_P.t513 1.1255
R17071 VDAC_P.n741 VDAC_P.t296 1.1255
R17072 VDAC_P.n742 VDAC_P.t1710 1.1255
R17073 VDAC_P.n743 VDAC_P.t68 1.1255
R17074 VDAC_P.n744 VDAC_P.t1282 1.1255
R17075 VDAC_P.n745 VDAC_P.t1233 1.1255
R17076 VDAC_P.n746 VDAC_P.t544 1.1255
R17077 VDAC_P.n106 VDAC_P.t1670 1.1255
R17078 VDAC_P.n747 VDAC_P.t1124 1.1255
R17079 VDAC_P.n748 VDAC_P.t1466 1.1255
R17080 VDAC_P.n749 VDAC_P.t2076 1.1255
R17081 VDAC_P.n750 VDAC_P.t2016 1.1255
R17082 VDAC_P.n751 VDAC_P.t1958 1.1255
R17083 VDAC_P.n752 VDAC_P.t808 1.1255
R17084 VDAC_P.n753 VDAC_P.t1734 1.1255
R17085 VDAC_P.n754 VDAC_P.t1347 1.1255
R17086 VDAC_P.n755 VDAC_P.t778 1.1255
R17087 VDAC_P.n756 VDAC_P.t1241 1.1255
R17088 VDAC_P.n757 VDAC_P.t1082 1.1255
R17089 VDAC_P.n758 VDAC_P.t581 1.1255
R17090 VDAC_P.n759 VDAC_P.t1583 1.1255
R17091 VDAC_P.n760 VDAC_P.t1273 1.1255
R17092 VDAC_P.n761 VDAC_P.t879 1.1255
R17093 VDAC_P.n762 VDAC_P.t292 1.1255
R17094 VDAC_P.n763 VDAC_P.t427 1.1255
R17095 VDAC_P.n764 VDAC_P.t1055 1.1255
R17096 VDAC_P.n765 VDAC_P.t1016 1.1255
R17097 VDAC_P.n766 VDAC_P.t1975 1.1255
R17098 VDAC_P.n767 VDAC_P.t1136 1.1255
R17099 VDAC_P.n768 VDAC_P.t1859 1.1255
R17100 VDAC_P.n769 VDAC_P.t692 1.1255
R17101 VDAC_P.n770 VDAC_P.t1294 1.1255
R17102 VDAC_P.n771 VDAC_P.t2105 1.1255
R17103 VDAC_P.n772 VDAC_P.t552 1.1255
R17104 VDAC_P.n773 VDAC_P.t522 1.1255
R17105 VDAC_P.n774 VDAC_P.t1232 1.1255
R17106 VDAC_P.n775 VDAC_P.t466 1.1255
R17107 VDAC_P.n776 VDAC_P.t804 1.1255
R17108 VDAC_P.n777 VDAC_P.t358 1.1255
R17109 VDAC_P.n778 VDAC_P.t1263 1.1255
R17110 VDAC_P.n779 VDAC_P.t1134 1.1255
R17111 VDAC_P.n780 VDAC_P.t1042 1.1255
R17112 VDAC_P.n781 VDAC_P.t769 1.1255
R17113 VDAC_P.n782 VDAC_P.t1846 1.1255
R17114 VDAC_P.n783 VDAC_P.t1393 1.1255
R17115 VDAC_P.n784 VDAC_P.t1406 1.1255
R17116 VDAC_P.n785 VDAC_P.t659 1.1255
R17117 VDAC_P.n786 VDAC_P.t887 1.1255
R17118 VDAC_P.n787 VDAC_P.t1169 1.1255
R17119 VDAC_P.n788 VDAC_P.t1723 1.1255
R17120 VDAC_P.n789 VDAC_P.t988 1.1255
R17121 VDAC_P.n790 VDAC_P.t121 1.1255
R17122 VDAC_P.n791 VDAC_P.t1971 1.1255
R17123 VDAC_P.n792 VDAC_P.t408 1.1255
R17124 VDAC_P.n793 VDAC_P.t1857 1.1255
R17125 VDAC_P.n794 VDAC_P.t676 1.1255
R17126 VDAC_P.n795 VDAC_P.t459 1.1255
R17127 VDAC_P.n796 VDAC_P.t1724 1.1255
R17128 VDAC_P.n797 VDAC_P.t2104 1.1255
R17129 VDAC_P.n798 VDAC_P.t287 1.1255
R17130 VDAC_P.n799 VDAC_P.t80 1.1255
R17131 VDAC_P.n800 VDAC_P.t246 1.1255
R17132 VDAC_P.n801 VDAC_P.t1556 1.1255
R17133 VDAC_P.n802 VDAC_P.t34 1.1255
R17134 VDAC_P.n803 VDAC_P.t1324 1.1255
R17135 VDAC_P.n804 VDAC_P.t578 1.1255
R17136 VDAC_P.n805 VDAC_P.t1155 1.1255
R17137 VDAC_P.n806 VDAC_P.t472 1.1255
R17138 VDAC_P.n807 VDAC_P.t1838 1.1255
R17139 VDAC_P.n808 VDAC_P.t1503 1.1255
R17140 VDAC_P.n809 VDAC_P.t826 1.1255
R17141 VDAC_P.n105 VDAC_P.t53 1.1255
R17142 VDAC_P.n810 VDAC_P.t1874 1.1255
R17143 VDAC_P.n811 VDAC_P.t1521 1.1255
R17144 VDAC_P.n812 VDAC_P.t838 1.1255
R17145 VDAC_P.n813 VDAC_P.t1307 1.1255
R17146 VDAC_P.n814 VDAC_P.t461 1.1255
R17147 VDAC_P.n815 VDAC_P.t1199 1.1255
R17148 VDAC_P.n816 VDAC_P.t435 1.1255
R17149 VDAC_P.n817 VDAC_P.t93 1.1255
R17150 VDAC_P.n818 VDAC_P.t1551 1.1255
R17151 VDAC_P.n819 VDAC_P.t1017 1.1255
R17152 VDAC_P.n820 VDAC_P.t683 1.1255
R17153 VDAC_P.n821 VDAC_P.t1893 1.1255
R17154 VDAC_P.n822 VDAC_P.t1604 1.1255
R17155 VDAC_P.n823 VDAC_P.t1467 1.1255
R17156 VDAC_P.n824 VDAC_P.t973 1.1255
R17157 VDAC_P.n825 VDAC_P.t192 1.1255
R17158 VDAC_P.n826 VDAC_P.t1813 1.1255
R17159 VDAC_P.n827 VDAC_P.t1804 1.1255
R17160 VDAC_P.n828 VDAC_P.t370 1.1255
R17161 VDAC_P.n829 VDAC_P.t284 1.1255
R17162 VDAC_P.n830 VDAC_P.t1912 1.1255
R17163 VDAC_P.n831 VDAC_P.t2053 1.1255
R17164 VDAC_P.n832 VDAC_P.t1472 1.1255
R17165 VDAC_P.n833 VDAC_P.t1674 1.1255
R17166 VDAC_P.n834 VDAC_P.t1140 1.1255
R17167 VDAC_P.n835 VDAC_P.t750 1.1255
R17168 VDAC_P.n836 VDAC_P.t325 1.1255
R17169 VDAC_P.n837 VDAC_P.t528 1.1255
R17170 VDAC_P.n838 VDAC_P.t563 1.1255
R17171 VDAC_P.n839 VDAC_P.t1600 1.1255
R17172 VDAC_P.n840 VDAC_P.t1738 1.1255
R17173 VDAC_P.n841 VDAC_P.t1453 1.1255
R17174 VDAC_P.n842 VDAC_P.t122 1.1255
R17175 VDAC_P.n843 VDAC_P.t1243 1.1255
R17176 VDAC_P.n844 VDAC_P.t445 1.1255
R17177 VDAC_P.n845 VDAC_P.t1137 1.1255
R17178 VDAC_P.n846 VDAC_P.t1585 1.1255
R17179 VDAC_P.n847 VDAC_P.t910 1.1255
R17180 VDAC_P.n848 VDAC_P.t1483 1.1255
R17181 VDAC_P.n849 VDAC_P.t981 1.1255
R17182 VDAC_P.n850 VDAC_P.t1359 1.1255
R17183 VDAC_P.n851 VDAC_P.t971 1.1255
R17184 VDAC_P.n852 VDAC_P.t468 1.1255
R17185 VDAC_P.n853 VDAC_P.t867 1.1255
R17186 VDAC_P.n854 VDAC_P.t1692 1.1255
R17187 VDAC_P.n855 VDAC_P.t314 1.1255
R17188 VDAC_P.n856 VDAC_P.t1039 1.1255
R17189 VDAC_P.n857 VDAC_P.t384 1.1255
R17190 VDAC_P.n858 VDAC_P.t507 1.1255
R17191 VDAC_P.n859 VDAC_P.t2004 1.1255
R17192 VDAC_P.n860 VDAC_P.t1458 1.1255
R17193 VDAC_P.n861 VDAC_P.t2124 1.1255
R17194 VDAC_P.n862 VDAC_P.t1238 1.1255
R17195 VDAC_P.n863 VDAC_P.t1093 1.1255
R17196 VDAC_P.n864 VDAC_P.t416 1.1255
R17197 VDAC_P.n865 VDAC_P.t1946 1.1255
R17198 VDAC_P.n866 VDAC_P.t304 1.1255
R17199 VDAC_P.n867 VDAC_P.t402 1.1255
R17200 VDAC_P.n868 VDAC_P.t685 1.1255
R17201 VDAC_P.n869 VDAC_P.t186 1.1255
R17202 VDAC_P.n870 VDAC_P.t1131 1.1255
R17203 VDAC_P.n871 VDAC_P.t1693 1.1255
R17204 VDAC_P.n872 VDAC_P.t2002 1.1255
R17205 VDAC_P.n104 VDAC_P.t500 1.1255
R17206 VDAC_P.n873 VDAC_P.t451 1.1255
R17207 VDAC_P.n874 VDAC_P.t1964 1.1255
R17208 VDAC_P.n875 VDAC_P.t823 1.1255
R17209 VDAC_P.n876 VDAC_P.t2067 1.1255
R17210 VDAC_P.n877 VDAC_P.t1536 1.1255
R17211 VDAC_P.n878 VDAC_P.t1963 1.1255
R17212 VDAC_P.n879 VDAC_P.t2132 1.1255
R17213 VDAC_P.n880 VDAC_P.t1502 1.1255
R17214 VDAC_P.n881 VDAC_P.t644 1.1255
R17215 VDAC_P.n882 VDAC_P.t650 1.1255
R17216 VDAC_P.n883 VDAC_P.t2097 1.1255
R17217 VDAC_P.n884 VDAC_P.t32 1.1255
R17218 VDAC_P.n885 VDAC_P.t1982 1.1255
R17219 VDAC_P.n886 VDAC_P.t1653 1.1255
R17220 VDAC_P.n887 VDAC_P.t547 1.1255
R17221 VDAC_P.n888 VDAC_P.t2120 1.1255
R17222 VDAC_P.n889 VDAC_P.t2003 1.1255
R17223 VDAC_P.n890 VDAC_P.t328 1.1255
R17224 VDAC_P.n891 VDAC_P.t1778 1.1255
R17225 VDAC_P.n892 VDAC_P.t1572 1.1255
R17226 VDAC_P.n893 VDAC_P.t1346 1.1255
R17227 VDAC_P.n894 VDAC_P.t1356 1.1255
R17228 VDAC_P.n895 VDAC_P.t1130 1.1255
R17229 VDAC_P.n896 VDAC_P.t2054 1.1255
R17230 VDAC_P.n897 VDAC_P.t360 1.1255
R17231 VDAC_P.n898 VDAC_P.t482 1.1255
R17232 VDAC_P.n899 VDAC_P.t1391 1.1255
R17233 VDAC_P.n900 VDAC_P.t1402 1.1255
R17234 VDAC_P.n901 VDAC_P.t1289 1.1255
R17235 VDAC_P.n902 VDAC_P.t610 1.1255
R17236 VDAC_P.n903 VDAC_P.t1070 1.1255
R17237 VDAC_P.n904 VDAC_P.t1641 1.1255
R17238 VDAC_P.n905 VDAC_P.t498 1.1255
R17239 VDAC_P.n906 VDAC_P.t1423 1.1255
R17240 VDAC_P.n907 VDAC_P.t1879 1.1255
R17241 VDAC_P.n908 VDAC_P.t677 1.1255
R17242 VDAC_P.n909 VDAC_P.t1773 1.1255
R17243 VDAC_P.n910 VDAC_P.t1107 1.1255
R17244 VDAC_P.n911 VDAC_P.t1675 1.1255
R17245 VDAC_P.n912 VDAC_P.t2127 1.1255
R17246 VDAC_P.n913 VDAC_P.t407 1.1255
R17247 VDAC_P.n914 VDAC_P.t2099 1.1255
R17248 VDAC_P.n915 VDAC_P.t1688 1.1255
R17249 VDAC_P.n916 VDAC_P.t1891 1.1255
R17250 VDAC_P.n917 VDAC_P.t788 1.1255
R17251 VDAC_P.n918 VDAC_P.t1562 1.1255
R17252 VDAC_P.n919 VDAC_P.t108 1.1255
R17253 VDAC_P.n920 VDAC_P.t1126 1.1255
R17254 VDAC_P.n921 VDAC_P.t65 1.1255
R17255 VDAC_P.n922 VDAC_P.t912 1.1255
R17256 VDAC_P.n923 VDAC_P.t254 1.1255
R17257 VDAC_P.n924 VDAC_P.t680 1.1255
R17258 VDAC_P.n925 VDAC_P.t426 1.1255
R17259 VDAC_P.n926 VDAC_P.t1285 1.1255
R17260 VDAC_P.n927 VDAC_P.t606 1.1255
R17261 VDAC_P.n928 VDAC_P.t1183 1.1255
R17262 VDAC_P.n929 VDAC_P.t968 1.1255
R17263 VDAC_P.n930 VDAC_P.t1898 1.1255
R17264 VDAC_P.n931 VDAC_P.t403 1.1255
R17265 VDAC_P.n932 VDAC_P.t850 1.1255
R17266 VDAC_P.n933 VDAC_P.t351 1.1255
R17267 VDAC_P.n934 VDAC_P.t1871 1.1255
R17268 VDAC_P.n935 VDAC_P.t1215 1.1255
R17269 VDAC_P.n103 VDAC_P.t117 1.1255
R17270 VDAC_P.n936 VDAC_P.t1526 1.1255
R17271 VDAC_P.n937 VDAC_P.t357 1.1255
R17272 VDAC_P.n938 VDAC_P.t1298 1.1255
R17273 VDAC_P.n939 VDAC_P.t1133 1.1255
R17274 VDAC_P.n940 VDAC_P.t805 1.1255
R17275 VDAC_P.n941 VDAC_P.t1018 1.1255
R17276 VDAC_P.n942 VDAC_P.t391 1.1255
R17277 VDAC_P.n943 VDAC_P.t1931 1.1255
R17278 VDAC_P.n944 VDAC_P.t1371 1.1255
R17279 VDAC_P.n945 VDAC_P.t477 1.1255
R17280 VDAC_P.n946 VDAC_P.t1163 1.1255
R17281 VDAC_P.n947 VDAC_P.t1717 1.1255
R17282 VDAC_P.n948 VDAC_P.t2126 1.1255
R17283 VDAC_P.n949 VDAC_P.t1425 1.1255
R17284 VDAC_P.n950 VDAC_P.t955 1.1255
R17285 VDAC_P.n951 VDAC_P.t1176 1.1255
R17286 VDAC_P.n952 VDAC_P.t1775 1.1255
R17287 VDAC_P.n953 VDAC_P.t1196 1.1255
R17288 VDAC_P.n954 VDAC_P.t190 1.1255
R17289 VDAC_P.n955 VDAC_P.t2129 1.1255
R17290 VDAC_P.n956 VDAC_P.t904 1.1255
R17291 VDAC_P.n957 VDAC_P.t2021 1.1255
R17292 VDAC_P.n958 VDAC_P.t48 1.1255
R17293 VDAC_P.n959 VDAC_P.t818 1.1255
R17294 VDAC_P.n960 VDAC_P.t236 1.1255
R17295 VDAC_P.n961 VDAC_P.t366 1.1255
R17296 VDAC_P.n962 VDAC_P.t603 1.1255
R17297 VDAC_P.n963 VDAC_P.t1888 1.1255
R17298 VDAC_P.n964 VDAC_P.t2094 1.1255
R17299 VDAC_P.n965 VDAC_P.t1440 1.1255
R17300 VDAC_P.n966 VDAC_P.t1662 1.1255
R17301 VDAC_P.n967 VDAC_P.t1411 1.1255
R17302 VDAC_P.n968 VDAC_P.t1450 1.1255
R17303 VDAC_P.n969 VDAC_P.t323 1.1255
R17304 VDAC_P.n970 VDAC_P.t1663 1.1255
R17305 VDAC_P.n971 VDAC_P.t161 1.1255
R17306 VDAC_P.n972 VDAC_P.t1559 1.1255
R17307 VDAC_P.n973 VDAC_P.t878 1.1255
R17308 VDAC_P.n974 VDAC_P.t1447 1.1255
R17309 VDAC_P.n975 VDAC_P.t1901 1.1255
R17310 VDAC_P.n976 VDAC_P.t1321 1.1255
R17311 VDAC_P.n977 VDAC_P.t489 1.1255
R17312 VDAC_P.n978 VDAC_P.t1444 1.1255
R17313 VDAC_P.n979 VDAC_P.t849 1.1255
R17314 VDAC_P.n980 VDAC_P.t2121 1.1255
R17315 VDAC_P.n981 VDAC_P.t1098 1.1255
R17316 VDAC_P.n982 VDAC_P.t2015 1.1255
R17317 VDAC_P.n983 VDAC_P.t1296 1.1255
R17318 VDAC_P.n984 VDAC_P.t1905 1.1255
R17319 VDAC_P.n985 VDAC_P.t1700 1.1255
R17320 VDAC_P.n986 VDAC_P.t70 1.1255
R17321 VDAC_P.n987 VDAC_P.t780 1.1255
R17322 VDAC_P.n988 VDAC_P.t594 1.1255
R17323 VDAC_P.n989 VDAC_P.t1054 1.1255
R17324 VDAC_P.n990 VDAC_P.t720 1.1255
R17325 VDAC_P.n991 VDAC_P.t950 1.1255
R17326 VDAC_P.n992 VDAC_P.t1940 1.1255
R17327 VDAC_P.n993 VDAC_P.t734 1.1255
R17328 VDAC_P.n994 VDAC_P.t667 1.1255
R17329 VDAC_P.n995 VDAC_P.t1218 1.1255
R17330 VDAC_P.n996 VDAC_P.t293 1.1255
R17331 VDAC_P.n997 VDAC_P.t1655 1.1255
R17332 VDAC_P.n998 VDAC_P.t266 1.1255
R17333 VDAC_P.n102 VDAC_P.t956 1.1255
R17334 VDAC_P.n999 VDAC_P.t789 1.1255
R17335 VDAC_P.n1000 VDAC_P.t1067 1.1255
R17336 VDAC_P.n1001 VDAC_P.t733 1.1255
R17337 VDAC_P.n1002 VDAC_P.t261 1.1255
R17338 VDAC_P.n1003 VDAC_P.t420 1.1255
R17339 VDAC_P.n1004 VDAC_P.t1791 1.1255
R17340 VDAC_P.n1005 VDAC_P.t1388 1.1255
R17341 VDAC_P.n1006 VDAC_P.t1138 1.1255
R17342 VDAC_P.n1007 VDAC_P.t388 1.1255
R17343 VDAC_P.n1008 VDAC_P.t1816 1.1255
R17344 VDAC_P.n1009 VDAC_P.t1923 1.1255
R17345 VDAC_P.n1010 VDAC_P.t1360 1.1255
R17346 VDAC_P.n1011 VDAC_P.t1626 1.1255
R17347 VDAC_P.n1012 VDAC_P.t1619 1.1255
R17348 VDAC_P.n1013 VDAC_P.t2071 1.1255
R17349 VDAC_P.n1014 VDAC_P.t512 1.1255
R17350 VDAC_P.n1015 VDAC_P.t997 1.1255
R17351 VDAC_P.n1016 VDAC_P.t1096 1.1255
R17352 VDAC_P.n1017 VDAC_P.t238 1.1255
R17353 VDAC_P.n1018 VDAC_P.t660 1.1255
R17354 VDAC_P.n1019 VDAC_P.t654 1.1255
R17355 VDAC_P.n1020 VDAC_P.t124 1.1255
R17356 VDAC_P.n1021 VDAC_P.t2088 1.1255
R17357 VDAC_P.n1022 VDAC_P.t518 1.1255
R17358 VDAC_P.n1023 VDAC_P.t1216 1.1255
R17359 VDAC_P.n1024 VDAC_P.t898 1.1255
R17360 VDAC_P.n1025 VDAC_P.t697 1.1255
R17361 VDAC_P.n1026 VDAC_P.t110 1.1255
R17362 VDAC_P.n1027 VDAC_P.t1259 1.1255
R17363 VDAC_P.n1028 VDAC_P.t574 1.1255
R17364 VDAC_P.n1029 VDAC_P.t2046 1.1255
R17365 VDAC_P.n1030 VDAC_P.t423 1.1255
R17366 VDAC_P.n1031 VDAC_P.t1830 1.1255
R17367 VDAC_P.n1032 VDAC_P.t113 1.1255
R17368 VDAC_P.n1033 VDAC_P.t937 1.1255
R17369 VDAC_P.n1034 VDAC_P.t185 1.1255
R17370 VDAC_P.n1035 VDAC_P.t1741 1.1255
R17371 VDAC_P.n1036 VDAC_P.t8 1.1255
R17372 VDAC_P.n1037 VDAC_P.t833 1.1255
R17373 VDAC_P.n1038 VDAC_P.t2089 1.1255
R17374 VDAC_P.n1039 VDAC_P.t1509 1.1255
R17375 VDAC_P.n1040 VDAC_P.t2063 1.1255
R17376 VDAC_P.n1041 VDAC_P.t1520 1.1255
R17377 VDAC_P.n1042 VDAC_P.t85 1.1255
R17378 VDAC_P.n1043 VDAC_P.t180 1.1255
R17379 VDAC_P.n1044 VDAC_P.t1494 1.1255
R17380 VDAC_P.n1045 VDAC_P.t380 1.1255
R17381 VDAC_P.n1046 VDAC_P.t2072 1.1255
R17382 VDAC_P.n1047 VDAC_P.t157 1.1255
R17383 VDAC_P.n1048 VDAC_P.t232 1.1255
R17384 VDAC_P.n1049 VDAC_P.t894 1.1255
R17385 VDAC_P.n1050 VDAC_P.t1168 1.1255
R17386 VDAC_P.n1051 VDAC_P.t410 1.1255
R17387 VDAC_P.n1052 VDAC_P.t1253 1.1255
R17388 VDAC_P.n1053 VDAC_P.t298 1.1255
R17389 VDAC_P.n1054 VDAC_P.t1151 1.1255
R17390 VDAC_P.n1055 VDAC_P.t1768 1.1255
R17391 VDAC_P.n1056 VDAC_P.t42 1.1255
R17392 VDAC_P.n1057 VDAC_P.t763 1.1255
R17393 VDAC_P.n1058 VDAC_P.t422 1.1255
R17394 VDAC_P.n1059 VDAC_P.t341 1.1255
R17395 VDAC_P.n1060 VDAC_P.t935 1.1255
R17396 VDAC_P.n1061 VDAC_P.t1177 1.1255
R17397 VDAC_P.n101 VDAC_P.t1115 1.1255
R17398 VDAC_P.n1062 VDAC_P.t840 1.1255
R17399 VDAC_P.n1063 VDAC_P.t514 1.1255
R17400 VDAC_P.n1064 VDAC_P.t312 1.1255
R17401 VDAC_P.n1065 VDAC_P.t1554 1.1255
R17402 VDAC_P.n1066 VDAC_P.t181 1.1255
R17403 VDAC_P.n1067 VDAC_P.t1322 1.1255
R17404 VDAC_P.n1068 VDAC_P.t589 1.1255
R17405 VDAC_P.n1069 VDAC_P.t1603 1.1255
R17406 VDAC_P.n1070 VDAC_P.t530 1.1255
R17407 VDAC_P.n1071 VDAC_P.t1497 1.1255
R17408 VDAC_P.n1072 VDAC_P.t1598 1.1255
R17409 VDAC_P.n1073 VDAC_P.t1383 1.1255
R17410 VDAC_P.n1074 VDAC_P.t481 1.1255
R17411 VDAC_P.n1075 VDAC_P.t1762 1.1255
R17412 VDAC_P.n1076 VDAC_P.t1361 1.1255
R17413 VDAC_P.n1077 VDAC_P.t501 1.1255
R17414 VDAC_P.n1078 VDAC_P.t641 1.1255
R17415 VDAC_P.n1079 VDAC_P.t133 1.1255
R17416 VDAC_P.n1080 VDAC_P.t1836 1.1255
R17417 VDAC_P.n1081 VDAC_P.t1605 1.1255
R17418 VDAC_P.n1082 VDAC_P.t1043 1.1255
R17419 VDAC_P.n1083 VDAC_P.t1499 1.1255
R17420 VDAC_P.n1084 VDAC_P.t1951 1.1255
R17421 VDAC_P.n1085 VDAC_P.t2068 1.1255
R17422 VDAC_P.n1086 VDAC_P.t883 1.1255
R17423 VDAC_P.n1087 VDAC_P.t1172 1.1255
R17424 VDAC_P.n1088 VDAC_P.t334 1.1255
R17425 VDAC_P.n1089 VDAC_P.t1057 1.1255
R17426 VDAC_P.n1090 VDAC_P.t2048 1.1255
R17427 VDAC_P.n1091 VDAC_P.t1987 1.1255
R17428 VDAC_P.n1092 VDAC_P.t1160 1.1255
R17429 VDAC_P.n1093 VDAC_P.t1746 1.1255
R17430 VDAC_P.n1094 VDAC_P.t1428 1.1255
R17431 VDAC_P.n1095 VDAC_P.t350 1.1255
R17432 VDAC_P.n1096 VDAC_P.t585 1.1255
R17433 VDAC_P.n1097 VDAC_P.t562 1.1255
R17434 VDAC_P.n1098 VDAC_P.t278 1.1255
R17435 VDAC_P.n1099 VDAC_P.t1288 1.1255
R17436 VDAC_P.n1100 VDAC_P.t918 1.1255
R17437 VDAC_P.n1101 VDAC_P.t703 1.1255
R17438 VDAC_P.n1102 VDAC_P.t790 1.1255
R17439 VDAC_P.n1103 VDAC_P.t361 1.1255
R17440 VDAC_P.n1104 VDAC_P.t251 1.1255
R17441 VDAC_P.n1105 VDAC_P.t63 1.1255
R17442 VDAC_P.n1106 VDAC_P.t815 1.1255
R17443 VDAC_P.n1107 VDAC_P.t1180 1.1255
R17444 VDAC_P.n1108 VDAC_P.t1495 1.1255
R17445 VDAC_P.n1109 VDAC_P.t1949 1.1255
R17446 VDAC_P.n1110 VDAC_P.t705 1.1255
R17447 VDAC_P.n1111 VDAC_P.t1839 1.1255
R17448 VDAC_P.n1112 VDAC_P.t580 1.1255
R17449 VDAC_P.n1113 VDAC_P.t1733 1.1255
R17450 VDAC_P.n1114 VDAC_P.t572 1.1255
R17451 VDAC_P.n1115 VDAC_P.t2024 1.1255
R17452 VDAC_P.n1116 VDAC_P.t89 1.1255
R17453 VDAC_P.n1117 VDAC_P.t816 1.1255
R17454 VDAC_P.n1118 VDAC_P.t947 1.1255
R17455 VDAC_P.n1119 VDAC_P.t708 1.1255
R17456 VDAC_P.n1120 VDAC_P.t1534 1.1255
R17457 VDAC_P.n1121 VDAC_P.t1020 1.1255
R17458 VDAC_P.n1122 VDAC_P.t1086 1.1255
R17459 VDAC_P.n1123 VDAC_P.t305 1.1255
R17460 VDAC_P.n1124 VDAC_P.t240 1.1255
R17461 VDAC_P.n100 VDAC_P.t951 1.1255
R17462 VDAC_P.n1125 VDAC_P.t1219 1.1255
R17463 VDAC_P.n1126 VDAC_P.t1769 1.1255
R17464 VDAC_P.n1127 VDAC_P.t565 1.1255
R17465 VDAC_P.n1128 VDAC_P.t31 1.1255
R17466 VDAC_P.n1129 VDAC_P.t2017 1.1255
R17467 VDAC_P.n1130 VDAC_P.t385 1.1255
R17468 VDAC_P.n1131 VDAC_P.t263 1.1255
R17469 VDAC_P.n1132 VDAC_P.t1716 1.1255
R17470 VDAC_P.n1133 VDAC_P.t1803 1.1255
R17471 VDAC_P.n1134 VDAC_P.t1580 1.1255
R17472 VDAC_P.n1135 VDAC_P.t419 1.1255
R17473 VDAC_P.n1136 VDAC_P.t1372 1.1255
R17474 VDAC_P.n1137 VDAC_P.t1864 1.1255
R17475 VDAC_P.n1138 VDAC_P.t1089 1.1255
R17476 VDAC_P.n1139 VDAC_P.t1555 1.1255
R17477 VDAC_P.n1140 VDAC_P.t1069 1.1255
R17478 VDAC_P.n1141 VDAC_P.t1441 1.1255
R17479 VDAC_P.n1142 VDAC_P.t1897 1.1255
R17480 VDAC_P.n1143 VDAC_P.t1248 1.1255
R17481 VDAC_P.n1144 VDAC_P.t1793 1.1255
R17482 VDAC_P.n1145 VDAC_P.t748 1.1255
R17483 VDAC_P.n1146 VDAC_P.t443 1.1255
R17484 VDAC_P.n1147 VDAC_P.t2114 1.1255
R17485 VDAC_P.n1148 VDAC_P.t1832 1.1255
R17486 VDAC_P.n1149 VDAC_P.t977 1.1255
R17487 VDAC_P.n1150 VDAC_P.t1368 1.1255
R17488 VDAC_P.n1151 VDAC_P.t1634 1.1255
R17489 VDAC_P.n1152 VDAC_P.t972 1.1255
R17490 VDAC_P.n1153 VDAC_P.t1418 1.1255
R17491 VDAC_P.n1154 VDAC_P.t9 1.1255
R17492 VDAC_P.n1155 VDAC_P.t504 1.1255
R17493 VDAC_P.n1156 VDAC_P.t17 1.1255
R17494 VDAC_P.n1157 VDAC_P.t1504 1.1255
R17495 VDAC_P.n1158 VDAC_P.t54 1.1255
R17496 VDAC_P.n1159 VDAC_P.t1331 1.1255
R17497 VDAC_P.n1160 VDAC_P.t758 1.1255
R17498 VDAC_P.n1161 VDAC_P.t1227 1.1255
R17499 VDAC_P.n1162 VDAC_P.t2064 1.1255
R17500 VDAC_P.n1163 VDAC_P.t299 1.1255
R17501 VDAC_P.n1164 VDAC_P.t1571 1.1255
R17502 VDAC_P.n1165 VDAC_P.t1926 1.1255
R17503 VDAC_P.n1166 VDAC_P.t123 1.1255
R17504 VDAC_P.n1167 VDAC_P.t1015 1.1255
R17505 VDAC_P.n1168 VDAC_P.t681 1.1255
R17506 VDAC_P.n1169 VDAC_P.t83 1.1255
R17507 VDAC_P.n1170 VDAC_P.t52 1.1255
R17508 VDAC_P.n1171 VDAC_P.t1683 1.1255
R17509 VDAC_P.n1172 VDAC_P.t864 1.1255
R17510 VDAC_P.n1173 VDAC_P.t801 1.1255
R17511 VDAC_P.n1174 VDAC_P.t529 1.1255
R17512 VDAC_P.n1175 VDAC_P.t1352 1.1255
R17513 VDAC_P.n1176 VDAC_P.t1919 1.1255
R17514 VDAC_P.n1177 VDAC_P.t932 1.1255
R17515 VDAC_P.n1178 VDAC_P.t114 1.1255
R17516 VDAC_P.n1179 VDAC_P.t796 1.1255
R17517 VDAC_P.n1180 VDAC_P.t1190 1.1255
R17518 VDAC_P.n1181 VDAC_P.t2057 1.1255
R17519 VDAC_P.n1182 VDAC_P.t1488 1.1255
R17520 VDAC_P.n1183 VDAC_P.t1906 1.1255
R17521 VDAC_P.n1184 VDAC_P.t1044 1.1255
R17522 VDAC_P.n1185 VDAC_P.t754 1.1255
R17523 VDAC_P.n1186 VDAC_P.t1325 1.1255
R17524 VDAC_P.n1187 VDAC_P.t1250 1.1255
R17525 VDAC_P.n99 VDAC_P.t2032 1.1255
R17526 VDAC_P.n1188 VDAC_P.t1981 1.1255
R17527 VDAC_P.n1189 VDAC_P.t1608 1.1255
R17528 VDAC_P.n1190 VDAC_P.t143 1.1255
R17529 VDAC_P.n1191 VDAC_P.t1396 1.1255
R17530 VDAC_P.n1192 VDAC_P.t1306 1.1255
R17531 VDAC_P.n1193 VDAC_P.t60 1.1255
R17532 VDAC_P.n1194 VDAC_P.t558 1.1255
R17533 VDAC_P.n1195 VDAC_P.t1022 1.1255
R17534 VDAC_P.n1196 VDAC_P.t1728 1.1255
R17535 VDAC_P.n1197 VDAC_P.t1798 1.1255
R17536 VDAC_P.n1198 VDAC_P.t436 1.1255
R17537 VDAC_P.n1199 VDAC_P.t1578 1.1255
R17538 VDAC_P.n1200 VDAC_P.t1267 1.1255
R17539 VDAC_P.n1201 VDAC_P.t1281 1.1255
R17540 VDAC_P.n1202 VDAC_P.t1737 1.1255
R17541 VDAC_P.n1203 VDAC_P.t596 1.1255
R17542 VDAC_P.n1204 VDAC_P.t229 1.1255
R17543 VDAC_P.n1205 VDAC_P.t2085 1.1255
R17544 VDAC_P.n1206 VDAC_P.t280 1.1255
R17545 VDAC_P.n1207 VDAC_P.t1007 1.1255
R17546 VDAC_P.n1208 VDAC_P.t592 1.1255
R17547 VDAC_P.n1209 VDAC_P.t1869 1.1255
R17548 VDAC_P.n1210 VDAC_P.t724 1.1255
R17549 VDAC_P.n1211 VDAC_P.t1314 1.1255
R17550 VDAC_P.n1212 VDAC_P.t2119 1.1255
R17551 VDAC_P.n1213 VDAC_P.t1094 1.1255
R17552 VDAC_P.n1214 VDAC_P.t2026 1.1255
R17553 VDAC_P.n1215 VDAC_P.t1280 1.1255
R17554 VDAC_P.n1216 VDAC_P.t1806 1.1255
R17555 VDAC_P.n1217 VDAC_P.t1684 1.1255
R17556 VDAC_P.n1218 VDAC_P.t362 1.1255
R17557 VDAC_P.n1219 VDAC_P.t1271 1.1255
R17558 VDAC_P.n1220 VDAC_P.t310 1.1255
R17559 VDAC_P.n1221 VDAC_P.t2074 1.1255
R17560 VDAC_P.n1222 VDAC_P.t773 1.1255
R17561 VDAC_P.n1223 VDAC_P.t946 1.1255
R17562 VDAC_P.n1224 VDAC_P.t1403 1.1255
R17563 VDAC_P.n1225 VDAC_P.t730 1.1255
R17564 VDAC_P.n1226 VDAC_P.t1301 1.1255
R17565 VDAC_P.n1227 VDAC_P.t55 1.1255
R17566 VDAC_P.n1228 VDAC_P.t601 1.1255
R17567 VDAC_P.n1229 VDAC_P.t1731 1.1255
R17568 VDAC_P.n1230 VDAC_P.t1084 1.1255
R17569 VDAC_P.n1231 VDAC_P.t1523 1.1255
R17570 VDAC_P.n1232 VDAC_P.t1979 1.1255
R17571 VDAC_P.n1233 VDAC_P.t1592 1.1255
R17572 VDAC_P.n1234 VDAC_P.t487 1.1255
R17573 VDAC_P.n1235 VDAC_P.t1380 1.1255
R17574 VDAC_P.n1236 VDAC_P.t1759 1.1255
R17575 VDAC_P.n1237 VDAC_P.t508 1.1255
R17576 VDAC_P.n1238 VDAC_P.t94 1.1255
R17577 VDAC_P.n1239 VDAC_P.t2107 1.1255
R17578 VDAC_P.n1240 VDAC_P.t1720 1.1255
R17579 VDAC_P.n1241 VDAC_P.t138 1.1255
R17580 VDAC_P.n1242 VDAC_P.t836 1.1255
R17581 VDAC_P.n1243 VDAC_P.t802 1.1255
R17582 VDAC_P.n1244 VDAC_P.t1452 1.1255
R17583 VDAC_P.n1245 VDAC_P.t98 1.1255
R17584 VDAC_P.n1246 VDAC_P.t99 1.1255
R17585 VDAC_P.n1247 VDAC_P.t928 1.1255
R17586 VDAC_P.n1248 VDAC_P.t942 1.1255
R17587 VDAC_P.n1249 VDAC_P.t399 1.1255
R17588 VDAC_P.n1250 VDAC_P.t830 1.1255
R17589 VDAC_P.n98 VDAC_P.t1549 1.1255
R17590 VDAC_P.n1251 VDAC_P.t1702 1.1255
R17591 VDAC_P.n1252 VDAC_P.t1435 1.1255
R17592 VDAC_P.n1253 VDAC_P.t1498 1.1255
R17593 VDAC_P.n1254 VDAC_P.t1231 1.1255
R17594 VDAC_P.n1255 VDAC_P.t1685 1.1255
R17595 VDAC_P.n1256 VDAC_P.t1117 1.1255
R17596 VDAC_P.n1257 VDAC_P.t415 1.1255
R17597 VDAC_P.n1258 VDAC_P.t2033 1.1255
R17598 VDAC_P.n1259 VDAC_P.t749 1.1255
R17599 VDAC_P.n1260 VDAC_P.t975 1.1255
R17600 VDAC_P.n1261 VDAC_P.t335 1.1255
R17601 VDAC_P.n1262 VDAC_P.t1815 1.1255
R17602 VDAC_P.n1263 VDAC_P.t940 1.1255
R17603 VDAC_P.n1264 VDAC_P.t294 1.1255
R17604 VDAC_P.n1265 VDAC_P.t526 1.1255
R17605 VDAC_P.n1266 VDAC_P.t809 1.1255
R17606 VDAC_P.n1267 VDAC_P.t914 1.1255
R17607 VDAC_P.n1268 VDAC_P.t1375 1.1255
R17608 VDAC_P.n1269 VDAC_P.t983 1.1255
R17609 VDAC_P.n1270 VDAC_P.t183 1.1255
R17610 VDAC_P.n1271 VDAC_P.t877 1.1255
R17611 VDAC_P.n1272 VDAC_P.t597 1.1255
R17612 VDAC_P.n1273 VDAC_P.t227 1.1255
R17613 VDAC_P.n1274 VDAC_P.t2075 1.1255
R17614 VDAC_P.n1275 VDAC_P.t1401 1.1255
R17615 VDAC_P.n1276 VDAC_P.t1969 1.1255
R17616 VDAC_P.n1277 VDAC_P.t1112 1.1255
R17617 VDAC_P.n1278 VDAC_P.t891 1.1255
R17618 VDAC_P.n1279 VDAC_P.t1316 1.1255
R17619 VDAC_P.n1280 VDAC_P.t1651 1.1255
R17620 VDAC_P.n1281 VDAC_P.t1065 1.1255
R17621 VDAC_P.n1282 VDAC_P.t1064 1.1255
R17622 VDAC_P.n1283 VDAC_P.t1999 1.1255
R17623 VDAC_P.n1284 VDAC_P.t624 1.1255
R17624 VDAC_P.n1285 VDAC_P.t1566 1.1255
R17625 VDAC_P.n1286 VDAC_P.t1540 1.1255
R17626 VDAC_P.n1287 VDAC_P.t686 1.1255
R17627 VDAC_P.n1288 VDAC_P.t95 1.1255
R17628 VDAC_P.n1289 VDAC_P.t302 1.1255
R17629 VDAC_P.n1290 VDAC_P.t2050 1.1255
R17630 VDAC_P.n1291 VDAC_P.t872 1.1255
R17631 VDAC_P.n1292 VDAC_P.t2006 1.1255
R17632 VDAC_P.n1293 VDAC_P.t1479 1.1255
R17633 VDAC_P.n1294 VDAC_P.t414 1.1255
R17634 VDAC_P.n1295 VDAC_P.t1265 1.1255
R17635 VDAC_P.n1296 VDAC_P.t1823 1.1255
R17636 VDAC_P.n1297 VDAC_P.t1161 1.1255
R17637 VDAC_P.n1298 VDAC_P.t1617 1.1255
R17638 VDAC_P.n1299 VDAC_P.t2058 1.1255
R17639 VDAC_P.n1300 VDAC_P.t1511 1.1255
R17640 VDAC_P.n1301 VDAC_P.t995 1.1255
R17641 VDAC_P.n1302 VDAC_P.t711 1.1255
R17642 VDAC_P.n1303 VDAC_P.t1853 1.1255
R17643 VDAC_P.n1304 VDAC_P.t1252 1.1255
R17644 VDAC_P.n1305 VDAC_P.t1647 1.1255
R17645 VDAC_P.n1306 VDAC_P.t764 1.1255
R17646 VDAC_P.n1307 VDAC_P.t783 1.1255
R17647 VDAC_P.n1308 VDAC_P.t151 1.1255
R17648 VDAC_P.n1309 VDAC_P.t1664 1.1255
R17649 VDAC_P.n1310 VDAC_P.t1883 1.1255
R17650 VDAC_P.n1311 VDAC_P.t1508 1.1255
R17651 VDAC_P.n1312 VDAC_P.t1558 1.1255
R17652 VDAC_P.n1313 VDAC_P.t620 1.1255
R17653 VDAC_P.n97 VDAC_P.t1236 1.1255
R17654 VDAC_P.n1314 VDAC_P.t1645 1.1255
R17655 VDAC_P.n1315 VDAC_P.t1468 1.1255
R17656 VDAC_P.n1316 VDAC_P.t405 1.1255
R17657 VDAC_P.n1317 VDAC_P.t1011 1.1255
R17658 VDAC_P.n1318 VDAC_P.t1184 1.1255
R17659 VDAC_P.n1319 VDAC_P.t1881 1.1255
R17660 VDAC_P.n1320 VDAC_P.t1492 1.1255
R17661 VDAC_P.n1321 VDAC_P.t1326 1.1255
R17662 VDAC_P.n1322 VDAC_P.t172 1.1255
R17663 VDAC_P.n1323 VDAC_P.t1110 1.1255
R17664 VDAC_P.n1324 VDAC_P.t1027 1.1255
R17665 VDAC_P.n1325 VDAC_P.t1776 1.1255
R17666 VDAC_P.n1326 VDAC_P.t1822 1.1255
R17667 VDAC_P.n1327 VDAC_P.t210 1.1255
R17668 VDAC_P.n1328 VDAC_P.t327 1.1255
R17669 VDAC_P.n1329 VDAC_P.t1777 1.1255
R17670 VDAC_P.n1330 VDAC_P.t1109 1.1255
R17671 VDAC_P.n1331 VDAC_P.t413 1.1255
R17672 VDAC_P.n1332 VDAC_P.t291 1.1255
R17673 VDAC_P.n1333 VDAC_P.t745 1.1255
R17674 VDAC_P.n1334 VDAC_P.t1915 1.1255
R17675 VDAC_P.n1335 VDAC_P.t111 1.1255
R17676 VDAC_P.n1336 VDAC_P.t1807 1.1255
R17677 VDAC_P.n1337 VDAC_P.t1708 1.1255
R17678 VDAC_P.n1338 VDAC_P.t813 1.1255
R17679 VDAC_P.n1339 VDAC_P.t1948 1.1255
R17680 VDAC_P.n1340 VDAC_P.t960 1.1255
R17681 VDAC_P.n1341 VDAC_P.t987 1.1255
R17682 VDAC_P.n1342 VDAC_P.t1448 1.1255
R17683 VDAC_P.n1343 VDAC_P.t141 1.1255
R17684 VDAC_P.n1344 VDAC_P.t564 1.1255
R17685 VDAC_P.n1345 VDAC_P.t742 1.1255
R17686 VDAC_P.n1346 VDAC_P.t554 1.1255
R17687 VDAC_P.n1347 VDAC_P.t2008 1.1255
R17688 VDAC_P.n1348 VDAC_P.t1950 1.1255
R17689 VDAC_P.n1349 VDAC_P.t1576 1.1255
R17690 VDAC_P.n1350 VDAC_P.t1730 1.1255
R17691 VDAC_P.n1351 VDAC_P.t196 1.1255
R17692 VDAC_P.n1352 VDAC_P.t1522 1.1255
R17693 VDAC_P.n1353 VDAC_P.t331 1.1255
R17694 VDAC_P.n1354 VDAC_P.t1246 1.1255
R17695 VDAC_P.n1355 VDAC_P.t623 1.1255
R17696 VDAC_P.n1356 VDAC_P.t1671 1.1255
R17697 VDAC_P.n1357 VDAC_P.t994 1.1255
R17698 VDAC_P.n1358 VDAC_P.t1457 1.1255
R17699 VDAC_P.n1359 VDAC_P.t525 1.1255
R17700 VDAC_P.n1360 VDAC_P.t689 1.1255
R17701 VDAC_P.n1361 VDAC_P.t139 1.1255
R17702 VDAC_P.n1362 VDAC_P.t1245 1.1255
R17703 VDAC_P.n1363 VDAC_P.t1699 1.1255
R17704 VDAC_P.n1364 VDAC_P.t348 1.1255
R17705 VDAC_P.n1365 VDAC_P.t1589 1.1255
R17706 VDAC_P.n1366 VDAC_P.t2045 1.1255
R17707 VDAC_P.n1367 VDAC_P.t1416 1.1255
R17708 VDAC_P.n1368 VDAC_P.t1831 1.1255
R17709 VDAC_P.n1369 VDAC_P.t1956 1.1255
R17710 VDAC_P.n1370 VDAC_P.t1725 1.1255
R17711 VDAC_P.n1371 VDAC_P.t2130 1.1255
R17712 VDAC_P.n1372 VDAC_P.t1222 1.1255
R17713 VDAC_P.n1373 VDAC_P.t1051 1.1255
R17714 VDAC_P.n1374 VDAC_P.t1552 1.1255
R17715 VDAC_P.n1375 VDAC_P.t1934 1.1255
R17716 VDAC_P.n1376 VDAC_P.t568 1.1255
R17717 VDAC_P.n96 VDAC_P.t621 1.1255
R17718 VDAC_P.n1377 VDAC_P.t1024 1.1255
R17719 VDAC_P.n1378 VDAC_P.t1097 1.1255
R17720 VDAC_P.n1379 VDAC_P.t224 1.1255
R17721 VDAC_P.n1380 VDAC_P.t882 1.1255
R17722 VDAC_P.n1381 VDAC_P.t193 1.1255
R17723 VDAC_P.n1382 VDAC_P.t1530 1.1255
R17724 VDAC_P.n1383 VDAC_P.t635 1.1255
R17725 VDAC_P.n1384 VDAC_P.t1695 1.1255
R17726 VDAC_P.n1385 VDAC_P.t1135 1.1255
R17727 VDAC_P.n1386 VDAC_P.t417 1.1255
R17728 VDAC_P.n1387 VDAC_P.t1790 1.1255
R17729 VDAC_P.n1388 VDAC_P.t1481 1.1255
R17730 VDAC_P.n1389 VDAC_P.t1933 1.1255
R17731 VDAC_P.n1390 VDAC_P.t1244 1.1255
R17732 VDAC_P.n1391 VDAC_P.t1872 1.1255
R17733 VDAC_P.n1392 VDAC_P.t1058 1.1255
R17734 VDAC_P.n1393 VDAC_P.t376 1.1255
R17735 VDAC_P.n1394 VDAC_P.t1654 1.1255
R17736 VDAC_P.n1395 VDAC_P.t1409 1.1255
R17737 VDAC_P.n1396 VDAC_P.t1442 1.1255
R17738 VDAC_P.n1397 VDAC_P.t1205 1.1255
R17739 VDAC_P.n1398 VDAC_P.t178 1.1255
R17740 VDAC_P.n1399 VDAC_P.t559 1.1255
R17741 VDAC_P.n1400 VDAC_P.t1557 1.1255
R17742 VDAC_P.n1401 VDAC_P.t1722 1.1255
R17743 VDAC_P.n1402 VDAC_P.t1445 1.1255
R17744 VDAC_P.n1403 VDAC_P.t1899 1.1255
R17745 VDAC_P.n1404 VDAC_P.t179 1.1255
R17746 VDAC_P.n1405 VDAC_P.t249 1.1255
R17747 VDAC_P.n1406 VDAC_P.t577 1.1255
R17748 VDAC_P.n1407 VDAC_P.t125 1.1255
R17749 VDAC_P.n1408 VDAC_P.t2118 1.1255
R17750 VDAC_P.n1409 VDAC_P.t751 1.1255
R17751 VDAC_P.n1410 VDAC_P.t503 1.1255
R17752 VDAC_P.n1411 VDAC_P.t260 1.1255
R17753 VDAC_P.n1412 VDAC_P.t1821 1.1255
R17754 VDAC_P.n1413 VDAC_P.t268 1.1255
R17755 VDAC_P.n1414 VDAC_P.t127 1.1255
R17756 VDAC_P.n1415 VDAC_P.t476 1.1255
R17757 VDAC_P.n1416 VDAC_P.t984 1.1255
R17758 VDAC_P.n1417 VDAC_P.t1035 1.1255
R17759 VDAC_P.n1418 VDAC_P.t944 1.1255
R17760 VDAC_P.n1419 VDAC_P.t1870 1.1255
R17761 VDAC_P.n1420 VDAC_P.t1908 1.1255
R17762 VDAC_P.n1421 VDAC_P.t1438 1.1255
R17763 VDAC_P.n1422 VDAC_P.t1305 1.1255
R17764 VDAC_P.n1423 VDAC_P.t102 1.1255
R17765 VDAC_P.n1424 VDAC_P.t557 1.1255
R17766 VDAC_P.n1425 VDAC_P.t992 1.1255
R17767 VDAC_P.n1426 VDAC_P.t1930 1.1255
R17768 VDAC_P.n1427 VDAC_P.t1437 1.1255
R17769 VDAC_P.n1428 VDAC_P.t1706 1.1255
R17770 VDAC_P.n1429 VDAC_P.t1337 1.1255
R17771 VDAC_P.n1430 VDAC_P.t909 1.1255
R17772 VDAC_P.n1431 VDAC_P.t301 1.1255
R17773 VDAC_P.n1432 VDAC_P.t1687 1.1255
R17774 VDAC_P.n1433 VDAC_P.t150 1.1255
R17775 VDAC_P.n1434 VDAC_P.t389 1.1255
R17776 VDAC_P.n1435 VDAC_P.t2035 1.1255
R17777 VDAC_P.n1436 VDAC_P.t1363 1.1255
R17778 VDAC_P.n1437 VDAC_P.t1817 1.1255
R17779 VDAC_P.n1438 VDAC_P.t484 1.1255
R17780 VDAC_P.n1439 VDAC_P.t869 1.1255
R17781 VDAC_P.n95 VDAC_P.t1003 1.1255
R17782 VDAC_P.n1440 VDAC_P.t33 1.1255
R17783 VDAC_P.n1441 VDAC_P.t945 1.1255
R17784 VDAC_P.n1442 VDAC_P.t321 1.1255
R17785 VDAC_P.n1443 VDAC_P.t1657 1.1255
R17786 VDAC_P.n1444 VDAC_P.t2109 1.1255
R17787 VDAC_P.n1445 VDAC_P.t409 1.1255
R17788 VDAC_P.n1446 VDAC_P.t2007 1.1255
R17789 VDAC_P.n1447 VDAC_P.t104 1.1255
R17790 VDAC_P.n1448 VDAC_P.t961 1.1255
R17791 VDAC_P.n1449 VDAC_P.t820 1.1255
R17792 VDAC_P.n1450 VDAC_P.t1689 1.1255
R17793 VDAC_P.n1451 VDAC_P.t716 1.1255
R17794 VDAC_P.n1452 VDAC_P.t306 1.1255
R17795 VDAC_P.n1453 VDAC_P.t772 1.1255
R17796 VDAC_P.n1454 VDAC_P.t1334 1.1255
R17797 VDAC_P.n1455 VDAC_P.t643 1.1255
R17798 VDAC_P.n1456 VDAC_P.t1114 1.1255
R17799 VDAC_P.n1457 VDAC_P.t1034 1.1255
R17800 VDAC_P.n1458 VDAC_P.t1607 1.1255
R17801 VDAC_P.n1459 VDAC_P.t926 1.1255
R17802 VDAC_P.n1460 VDAC_P.t1387 1.1255
R17803 VDAC_P.n1461 VDAC_P.t226 1.1255
R17804 VDAC_P.n1462 VDAC_P.t655 1.1255
R17805 VDAC_P.n1463 VDAC_P.t135 1.1255
R17806 VDAC_P.n1464 VDAC_P.t546 1.1255
R17807 VDAC_P.n1465 VDAC_P.t1637 1.1255
R17808 VDAC_P.n1466 VDAC_P.t543 1.1255
R17809 VDAC_P.n1467 VDAC_P.t1415 1.1255
R17810 VDAC_P.n1468 VDAC_P.t273 1.1255
R17811 VDAC_P.n1469 VDAC_P.t189 1.1255
R17812 VDAC_P.n1470 VDAC_P.t897 1.1255
R17813 VDAC_P.n1471 VDAC_P.t116 1.1255
R17814 VDAC_P.n1472 VDAC_P.t1665 1.1255
R17815 VDAC_P.n1473 VDAC_P.t551 1.1255
R17816 VDAC_P.n1474 VDAC_P.t888 1.1255
R17817 VDAC_P.n1475 VDAC_P.t1021 1.1255
R17818 VDAC_P.n1476 VDAC_P.t344 1.1255
R17819 VDAC_P.n1477 VDAC_P.t1799 1.1255
R17820 VDAC_P.n1478 VDAC_P.t132 1.1255
R17821 VDAC_P.n1479 VDAC_P.t698 1.1255
R17822 VDAC_P.n1480 VDAC_P.t1132 1.1255
R17823 VDAC_P.n1481 VDAC_P.t674 1.1255
R17824 VDAC_P.n1482 VDAC_P.t1149 1.1255
R17825 VDAC_P.n1483 VDAC_P.t136 1.1255
R17826 VDAC_P.n1484 VDAC_P.t922 1.1255
R17827 VDAC_P.n1485 VDAC_P.t395 1.1255
R17828 VDAC_P.n1486 VDAC_P.t126 1.1255
R17829 VDAC_P.n1487 VDAC_P.t1279 1.1255
R17830 VDAC_P.n1488 VDAC_P.t1374 1.1255
R17831 VDAC_P.n1489 VDAC_P.t1175 1.1255
R17832 VDAC_P.n1490 VDAC_P.t429 1.1255
R17833 VDAC_P.n1491 VDAC_P.t2086 1.1255
R17834 VDAC_P.n1492 VDAC_P.t215 1.1255
R17835 VDAC_P.n1493 VDAC_P.t1005 1.1255
R17836 VDAC_P.n1494 VDAC_P.t349 1.1255
R17837 VDAC_P.n1495 VDAC_P.t1867 1.1255
R17838 VDAC_P.n1496 VDAC_P.t175 1.1255
R17839 VDAC_P.n1497 VDAC_P.t845 1.1255
R17840 VDAC_P.n1498 VDAC_P.t2044 1.1255
R17841 VDAC_P.n1499 VDAC_P.t219 1.1255
R17842 VDAC_P.n1500 VDAC_P.t2011 1.1255
R17843 VDAC_P.n1501 VDAC_P.t880 1.1255
R17844 VDAC_P.n1502 VDAC_P.t963 1.1255
R17845 VDAC_P.n94 VDAC_P.t1214 1.1255
R17846 VDAC_P.n1503 VDAC_P.t283 1.1255
R17847 VDAC_P.n1504 VDAC_P.t1960 1.1255
R17848 VDAC_P.n1505 VDAC_P.t1965 1.1255
R17849 VDAC_P.n1506 VDAC_P.t1088 1.1255
R17850 VDAC_P.n1507 VDAC_P.t766 1.1255
R17851 VDAC_P.n1508 VDAC_P.t340 1.1255
R17852 VDAC_P.n1509 VDAC_P.t106 1.1255
R17853 VDAC_P.n1510 VDAC_P.t575 1.1255
R17854 VDAC_P.n1511 VDAC_P.t2080 1.1255
R17855 VDAC_P.n1512 VDAC_P.t1986 1.1255
R17856 VDAC_P.n1513 VDAC_P.t1208 1.1255
R17857 VDAC_P.n1514 VDAC_P.t1766 1.1255
R17858 VDAC_P.n1515 VDAC_P.t1365 1.1255
R17859 VDAC_P.n1516 VDAC_P.t792 1.1255
R17860 VDAC_P.n1517 VDAC_P.t874 1.1255
R17861 VDAC_P.n1518 VDAC_P.t205 1.1255
R17862 VDAC_P.n1519 VDAC_P.t1514 1.1255
R17863 VDAC_P.n1520 VDAC_P.t1235 1.1255
R17864 VDAC_P.n1521 VDAC_P.t1795 1.1255
R17865 VDAC_P.n1522 VDAC_P.t1125 1.1255
R17866 VDAC_P.n1523 VDAC_P.t1579 1.1255
R17867 VDAC_P.n1524 VDAC_P.t1994 1.1255
R17868 VDAC_P.n1525 VDAC_P.t1473 1.1255
R17869 VDAC_P.n1526 VDAC_P.t1927 1.1255
R17870 VDAC_P.n1527 VDAC_P.t1261 1.1255
R17871 VDAC_P.n1528 VDAC_P.t1819 1.1255
R17872 VDAC_P.n1529 VDAC_P.t1932 1.1255
R17873 VDAC_P.n1530 VDAC_P.t1611 1.1255
R17874 VDAC_P.n1531 VDAC_P.t290 1.1255
R17875 VDAC_P.n1532 VDAC_P.t1505 1.1255
R17876 VDAC_P.n1533 VDAC_P.t269 1.1255
R17877 VDAC_P.n1534 VDAC_P.t1512 1.1255
R17878 VDAC_P.n1535 VDAC_P.t483 1.1255
R17879 VDAC_P.n1536 VDAC_P.t324 1.1255
R17880 VDAC_P.n1537 VDAC_P.t646 1.1255
R17881 VDAC_P.n1538 VDAC_P.t188 1.1255
R17882 VDAC_P.n1539 VDAC_P.t1048 1.1255
R17883 VDAC_P.n1540 VDAC_P.t1009 1.1255
R17884 VDAC_P.n1541 VDAC_P.t432 1.1255
R17885 VDAC_P.n1542 VDAC_P.t1758 1.1255
R17886 VDAC_P.n1543 VDAC_P.t1076 1.1255
R17887 VDAC_P.n1544 VDAC_P.t446 1.1255
R17888 VDAC_P.n1545 VDAC_P.t1335 1.1255
R17889 VDAC_P.n1546 VDAC_P.t1270 1.1255
R17890 VDAC_P.n1547 VDAC_P.t1119 1.1255
R17891 VDAC_P.n1548 VDAC_P.t235 1.1255
R17892 VDAC_P.n1549 VDAC_P.t1002 1.1255
R17893 VDAC_P.n1550 VDAC_P.t1471 1.1255
R17894 VDAC_P.n1551 VDAC_P.t462 1.1255
R17895 VDAC_P.n1552 VDAC_P.t695 1.1255
R17896 VDAC_P.n1553 VDAC_P.t475 1.1255
R17897 VDAC_P.n1554 VDAC_P.t1257 1.1255
R17898 VDAC_P.n1555 VDAC_P.t1709 1.1255
R17899 VDAC_P.n1556 VDAC_P.t20 1.1255
R17900 VDAC_P.n1557 VDAC_P.t1501 1.1255
R17901 VDAC_P.n1558 VDAC_P.t155 1.1255
R17902 VDAC_P.n1559 VDAC_P.t707 1.1255
R17903 VDAC_P.n1560 VDAC_P.t1845 1.1255
R17904 VDAC_P.n1561 VDAC_P.t2084 1.1255
R17905 VDAC_P.n1562 VDAC_P.t1739 1.1255
R17906 VDAC_P.n1563 VDAC_P.t636 1.1255
R17907 VDAC_P.n1564 VDAC_P.t642 1.1255
R17908 VDAC_P.n1565 VDAC_P.t2087 1.1255
R17909 VDAC_P.n93 VDAC_P.t431 1.1255
R17910 VDAC_P.n1566 VDAC_P.t1902 1.1255
R17911 VDAC_P.n1567 VDAC_P.t779 1.1255
R17912 VDAC_P.n1568 VDAC_P.t1678 1.1255
R17913 VDAC_P.n1569 VDAC_P.t1323 1.1255
R17914 VDAC_P.n1570 VDAC_P.t899 1.1255
R17915 VDAC_P.n1571 VDAC_P.t177 1.1255
R17916 VDAC_P.n1572 VDAC_P.t1673 1.1255
R17917 VDAC_P.n1573 VDAC_P.t159 1.1255
R17918 VDAC_P.n1574 VDAC_P.t1565 1.1255
R17919 VDAC_P.n1575 VDAC_P.t2019 1.1255
R17920 VDAC_P.n1576 VDAC_P.t359 1.1255
R17921 VDAC_P.n1577 VDAC_P.t969 1.1255
R17922 VDAC_P.n1578 VDAC_P.t1732 1.1255
R17923 VDAC_P.n1579 VDAC_P.t923 1.1255
R17924 VDAC_P.n1580 VDAC_P.t492 1.1255
R17925 VDAC_P.n1581 VDAC_P.t722 1.1255
R17926 VDAC_P.n1582 VDAC_P.t14 1.1255
R17927 VDAC_P.n1583 VDAC_P.t976 1.1255
R17928 VDAC_P.n1584 VDAC_P.t15 1.1255
R17929 VDAC_P.n1585 VDAC_P.t1496 1.1255
R17930 VDAC_P.n1586 VDAC_P.t1690 1.1255
R17931 VDAC_P.n1587 VDAC_P.t2100 1.1255
R17932 VDAC_P.n1588 VDAC_P.t1486 1.1255
R17933 VDAC_P.n1589 VDAC_P.t627 1.1255
R17934 VDAC_P.n1590 VDAC_P.t2056 1.1255
R17935 VDAC_P.n1591 VDAC_P.t1111 1.1255
R17936 VDAC_P.n1592 VDAC_P.t799 1.1255
R17937 VDAC_P.n1593 VDAC_P.t1754 1.1255
R17938 VDAC_P.n1594 VDAC_P.t387 1.1255
R17939 VDAC_P.n1595 VDAC_P.t218 1.1255
R17940 VDAC_P.n1596 VDAC_P.t639 1.1255
R17941 VDAC_P.n1597 VDAC_P.t1809 1.1255
R17942 VDAC_P.n1598 VDAC_P.t307 1.1255
R17943 VDAC_P.n1599 VDAC_P.t1599 1.1255
R17944 VDAC_P.n1600 VDAC_P.t281 1.1255
R17945 VDAC_P.n1601 VDAC_P.t1493 1.1255
R17946 VDAC_P.n1602 VDAC_P.t1947 1.1255
R17947 VDAC_P.n1603 VDAC_P.t1275 1.1255
R17948 VDAC_P.n1604 VDAC_P.t1837 1.1255
R17949 VDAC_P.n1605 VDAC_P.t1108 1.1255
R17950 VDAC_P.n1606 VDAC_P.t1707 1.1255
R17951 VDAC_P.n1607 VDAC_P.t140 1.1255
R17952 VDAC_P.n1608 VDAC_P.t1186 1.1255
R17953 VDAC_P.n1609 VDAC_P.t2055 1.1255
R17954 VDAC_P.n1610 VDAC_P.t392 1.1255
R17955 VDAC_P.n1611 VDAC_P.t262 1.1255
R17956 VDAC_P.n1612 VDAC_P.t532 1.1255
R17957 VDAC_P.n1613 VDAC_P.t1478 1.1255
R17958 VDAC_P.n1614 VDAC_P.t1156 1.1255
R17959 VDAC_P.n1615 VDAC_P.t638 1.1255
R17960 VDAC_P.n1616 VDAC_P.t1103 1.1255
R17961 VDAC_P.n1617 VDAC_P.t2040 1.1255
R17962 VDAC_P.n1618 VDAC_P.t1962 1.1255
R17963 VDAC_P.n1619 VDAC_P.t743 1.1255
R17964 VDAC_P.n1620 VDAC_P.t1542 1.1255
R17965 VDAC_P.n1621 VDAC_P.t1351 1.1255
R17966 VDAC_P.n1622 VDAC_P.t1310 1.1255
R17967 VDAC_P.n1623 VDAC_P.t1141 1.1255
R17968 VDAC_P.n1624 VDAC_P.t237 1.1255
R17969 VDAC_P.n1625 VDAC_P.t2022 1.1255
R17970 VDAC_P.n1626 VDAC_P.t1489 1.1255
R17971 VDAC_P.n1627 VDAC_P.t1037 1.1255
R17972 VDAC_P.n1628 VDAC_P.t365 1.1255
R17973 VDAC_P.n92 VDAC_P.t2036 1.1255
R17974 VDAC_P.n1629 VDAC_P.t881 1.1255
R17975 VDAC_P.n1630 VDAC_P.t308 1.1255
R17976 VDAC_P.n1631 VDAC_P.t1633 1.1255
R17977 VDAC_P.n1632 VDAC_P.t2083 1.1255
R17978 VDAC_P.n1633 VDAC_P.t1616 1.1255
R17979 VDAC_P.n1634 VDAC_P.t1983 1.1255
R17980 VDAC_P.n1635 VDAC_P.t168 1.1255
R17981 VDAC_P.n1636 VDAC_P.t406 1.1255
R17982 VDAC_P.n1637 VDAC_P.t372 1.1255
R17983 VDAC_P.n1638 VDAC_P.t38 1.1255
R17984 VDAC_P.n1639 VDAC_P.t1071 1.1255
R17985 VDAC_P.n1640 VDAC_P.t1090 1.1255
R17986 VDAC_P.n1641 VDAC_P.t2018 1.1255
R17987 VDAC_P.n1642 VDAC_P.t59 1.1255
R17988 VDAC_P.n1643 VDAC_P.t648 1.1255
R17989 VDAC_P.n1644 VDAC_P.t250 1.1255
R17990 VDAC_P.n1645 VDAC_P.t1668 1.1255
R17991 VDAC_P.n1646 VDAC_P.t1358 1.1255
R17992 VDAC_P.n1647 VDAC_P.t649 1.1255
R17993 VDAC_P.n1648 VDAC_P.t590 1.1255
R17994 VDAC_P.n1649 VDAC_P.t2070 1.1255
R17995 VDAC_P.n1650 VDAC_P.t936 1.1255
R17996 VDAC_P.n1651 VDAC_P.t486 1.1255
R17997 VDAC_P.n1652 VDAC_P.t715 1.1255
R17998 VDAC_P.n1653 VDAC_P.t1426 1.1255
R17999 VDAC_P.n1654 VDAC_P.t187 1.1255
R18000 VDAC_P.n1655 VDAC_P.t1755 1.1255
R18001 VDAC_P.n1656 VDAC_P.t25 1.1255
R18002 VDAC_P.n1657 VDAC_P.t231 1.1255
R18003 VDAC_P.n1658 VDAC_P.t1922 1.1255
R18004 VDAC_P.n1659 VDAC_P.t379 1.1255
R18005 VDAC_P.n1660 VDAC_P.t2001 1.1255
R18006 VDAC_P.n1661 VDAC_P.t1333 1.1255
R18007 VDAC_P.n1662 VDAC_P.t1787 1.1255
R18008 VDAC_P.n1663 VDAC_P.t684 1.1255
R18009 VDAC_P.n1664 VDAC_P.t855 1.1255
R18010 VDAC_P.n1665 VDAC_P.t450 1.1255
R18011 VDAC_P.n1666 VDAC_P.t73 1.1255
R18012 VDAC_P.n1667 VDAC_P.t2031 1.1255
R18013 VDAC_P.n1668 VDAC_P.t688 1.1255
R18014 VDAC_P.n1669 VDAC_P.t1895 1.1255
R18015 VDAC_P.n1670 VDAC_P.t1240 1.1255
R18016 VDAC_P.n1671 VDAC_P.t1574 1.1255
R18017 VDAC_P.n1672 VDAC_P.t1420 1.1255
R18018 VDAC_P.n1673 VDAC_P.t586 1.1255
R18019 VDAC_P.n1674 VDAC_P.t595 1.1255
R18020 VDAC_P.n1675 VDAC_P.t56 1.1255
R18021 VDAC_P.n1676 VDAC_P.t1854 1.1255
R18022 VDAC_P.n1677 VDAC_P.t696 1.1255
R18023 VDAC_P.n1678 VDAC_P.t78 1.1255
R18024 VDAC_P.n1679 VDAC_P.t345 1.1255
R18025 VDAC_P.n1680 VDAC_P.t1414 1.1255
R18026 VDAC_P.n1681 VDAC_P.t173 1.1255
R18027 VDAC_P.n1682 VDAC_P.t433 1.1255
R18028 VDAC_P.n1683 VDAC_P.t146 1.1255
R18029 VDAC_P.n1684 VDAC_P.t1539 1.1255
R18030 VDAC_P.n1685 VDAC_P.t858 1.1255
R18031 VDAC_P.n1686 VDAC_P.t679 1.1255
R18032 VDAC_P.n1687 VDAC_P.t57 1.1255
R18033 VDAC_P.n1688 VDAC_P.t1225 1.1255
R18034 VDAC_P.n1689 VDAC_P.t441 1.1255
R18035 VDAC_P.n1690 VDAC_P.t1228 1.1255
R18036 VDAC_P.n1691 VDAC_P.t1569 1.1255
R18037 VDAC_P.n91 VDAC_P.t347 1.1255
R18038 VDAC_P.n1692 VDAC_P.t1210 1.1255
R18039 VDAC_P.n1693 VDAC_P.t1197 1.1255
R18040 VDAC_P.n1694 VDAC_P.t1952 1.1255
R18041 VDAC_P.n1695 VDAC_P.t978 1.1255
R18042 VDAC_P.n1696 VDAC_P.t39 1.1255
R18043 VDAC_P.n1697 VDAC_P.t866 1.1255
R18044 VDAC_P.n1698 VDAC_P.t355 1.1255
R18045 VDAC_P.n1699 VDAC_P.t1789 1.1255
R18046 VDAC_P.n1700 VDAC_P.t329 1.1255
R18047 VDAC_P.n1701 VDAC_P.t857 1.1255
R18048 VDAC_P.n1702 VDAC_P.t1978 1.1255
R18049 VDAC_P.n1703 VDAC_P.t1577 1.1255
R18050 VDAC_P.n1704 VDAC_P.t1031 1.1255
R18051 VDAC_P.n1705 VDAC_P.t1299 1.1255
R18052 VDAC_P.n1706 VDAC_P.t1751 1.1255
R18053 VDAC_P.n1707 VDAC_P.t1284 1.1255
R18054 VDAC_P.n1708 VDAC_P.t1649 1.1255
R18055 VDAC_P.n1709 VDAC_P.t1063 1.1255
R18056 VDAC_P.n1710 VDAC_P.t1056 1.1255
R18057 VDAC_P.n1711 VDAC_P.t1997 1.1255
R18058 VDAC_P.n1712 VDAC_P.t176 1.1255
R18059 VDAC_P.n1713 VDAC_P.t957 1.1255
R18060 VDAC_P.n1714 VDAC_P.t1524 1.1255
R18061 VDAC_P.n1715 VDAC_P.t1338 1.1255
R18062 VDAC_P.n1716 VDAC_P.t587 1.1255
R18063 VDAC_P.n1717 VDAC_P.t1118 1.1255
R18064 VDAC_P.n1718 VDAC_P.t154 1.1255
R18065 VDAC_P.n1719 VDAC_P.t1336 1.1255
R18066 VDAC_P.n1720 VDAC_P.t478 1.1255
R18067 VDAC_P.n1721 VDAC_P.t1812 1.1255
R18068 VDAC_P.n1722 VDAC_P.t1394 1.1255
R18069 VDAC_P.n1723 VDAC_P.t1283 1.1255
R18070 VDAC_P.n1724 VDAC_P.t46 1.1255
R18071 VDAC_P.n1725 VDAC_P.t1066 1.1255
R18072 VDAC_P.n1726 VDAC_P.t1527 1.1255
R18073 VDAC_P.n1727 VDAC_P.t494 1.1255
R18074 VDAC_P.n1728 VDAC_P.t1417 1.1255
R18075 VDAC_P.n1729 VDAC_P.t118 1.1255
R18076 VDAC_P.n1730 VDAC_P.t673 1.1255
R18077 VDAC_P.n1731 VDAC_P.t1767 1.1255
R18078 VDAC_P.n1732 VDAC_P.t1187 1.1255
R18079 VDAC_P.n1733 VDAC_P.t1745 1.1255
R18080 VDAC_P.n1734 VDAC_P.t1404 1.1255
R18081 VDAC_P.n1735 VDAC_P.t1535 1.1255
R18082 VDAC_P.n1736 VDAC_P.t1993 1.1255
R18083 VDAC_P.n1737 VDAC_P.t1656 1.1255
R18084 VDAC_P.n1738 VDAC_P.t953 1.1255
R18085 VDAC_P.n1739 VDAC_P.t756 1.1255
R18086 VDAC_P.n1740 VDAC_P.t137 1.1255
R18087 VDAC_P.n1741 VDAC_P.t588 1.1255
R18088 VDAC_P.n1742 VDAC_P.t1106 1.1255
R18089 VDAC_P.n1743 VDAC_P.t1077 1.1255
R18090 VDAC_P.n1744 VDAC_P.t896 1.1255
R18091 VDAC_P.n1745 VDAC_P.t1818 1.1255
R18092 VDAC_P.n1746 VDAC_P.t1780 1.1255
R18093 VDAC_P.n1747 VDAC_P.t1602 1.1255
R18094 VDAC_P.n1748 VDAC_P.t844 1.1255
R18095 VDAC_P.n1749 VDAC_P.t1170 1.1255
R18096 VDAC_P.n1750 VDAC_P.t315 1.1255
R18097 VDAC_P.n1751 VDAC_P.t1880 1.1255
R18098 VDAC_P.n1752 VDAC_P.t1886 1.1255
R18099 VDAC_P.n1753 VDAC_P.t1525 1.1255
R18100 VDAC_P.n1754 VDAC_P.t1658 1.1255
R18101 VDAC_P.n90 VDAC_P.t2065 1.1255
R18102 VDAC_P.n1755 VDAC_P.t199 1.1255
R18103 VDAC_P.n1756 VDAC_P.t1961 1.1255
R18104 VDAC_P.n1757 VDAC_P.t1295 1.1255
R18105 VDAC_P.n1758 VDAC_P.t243 1.1255
R18106 VDAC_P.n1759 VDAC_P.t1532 1.1255
R18107 VDAC_P.n1760 VDAC_P.t837 1.1255
R18108 VDAC_P.n1761 VDAC_P.t2095 1.1255
R18109 VDAC_P.n1762 VDAC_P.t848 1.1255
R18110 VDAC_P.n1763 VDAC_P.t1995 1.1255
R18111 VDAC_P.n1764 VDAC_P.t608 1.1255
R18112 VDAC_P.n1765 VDAC_P.t247 1.1255
R18113 VDAC_P.n1766 VDAC_P.t212 1.1255
R18114 VDAC_P.n1767 VDAC_P.t678 1.1255
R18115 VDAC_P.n1768 VDAC_P.t759 1.1255
R18116 VDAC_P.n1769 VDAC_P.t1943 1.1255
R18117 VDAC_P.n1770 VDAC_P.t1432 1.1255
R18118 VDAC_P.n1771 VDAC_P.t1833 1.1255
R18119 VDAC_P.n1772 VDAC_P.t1068 1.1255
R18120 VDAC_P.n1773 VDAC_P.t1446 1.1255
R18121 VDAC_P.n1774 VDAC_P.t28 1.1255
R18122 VDAC_P.n1775 VDAC_P.t2000 1.1255
R18123 VDAC_P.n1776 VDAC_P.t2135 1.1255
R18124 VDAC_P.n1777 VDAC_P.t1560 1.1255
R18125 VDAC_P.n1778 VDAC_P.t1726 1.1255
R18126 VDAC_P.n1779 VDAC_P.t1348 1.1255
R18127 VDAC_P.n1780 VDAC_P.t214 1.1255
R18128 VDAC_P.n1781 VDAC_P.t633 1.1255
R18129 VDAC_P.n1782 VDAC_P.t1072 1.1255
R18130 VDAC_P.n1783 VDAC_P.t1127 1.1255
R18131 VDAC_P.n1784 VDAC_P.t1704 1.1255
R18132 VDAC_P.n1785 VDAC_P.t902 1.1255
R18133 VDAC_P.n1786 VDAC_P.t1475 1.1255
R18134 VDAC_P.n1787 VDAC_P.t798 1.1255
R18135 VDAC_P.n1788 VDAC_P.t645 1.1255
R18136 VDAC_P.n1789 VDAC_P.t1715 1.1255
R18137 VDAC_P.n1790 VDAC_P.t593 1.1255
R18138 VDAC_P.n1791 VDAC_P.t1613 1.1255
R18139 VDAC_P.n1792 VDAC_P.t934 1.1255
R18140 VDAC_P.n1793 VDAC_P.t767 1.1255
R18141 VDAC_P.n1794 VDAC_P.t1957 1.1255
R18142 VDAC_P.n1795 VDAC_P.t1373 1.1255
R18143 VDAC_P.n1796 VDAC_P.t147 1.1255
R18144 VDAC_P.n1797 VDAC_P.t1924 1.1255
R18145 VDAC_P.n1798 VDAC_P.t1721 1.1255
R18146 VDAC_P.n1799 VDAC_P.t1078 1.1255
R18147 VDAC_P.n1800 VDAC_P.t622 1.1255
R18148 VDAC_P.n1801 VDAC_P.t2069 1.1255
R18149 VDAC_P.n1802 VDAC_P.t784 1.1255
R18150 VDAC_P.n1803 VDAC_P.t149 1.1255
R18151 VDAC_P.n1804 VDAC_P.t160 1.1255
R18152 VDAC_P.n1805 VDAC_P.t1506 1.1255
R18153 VDAC_P.n1806 VDAC_P.t1268 1.1255
R18154 VDAC_P.n1807 VDAC_P.t1274 1.1255
R18155 VDAC_P.n1808 VDAC_P.t1121 1.1255
R18156 VDAC_P.n1809 VDAC_P.t856 1.1255
R18157 VDAC_P.n1810 VDAC_P.t1006 1.1255
R18158 VDAC_P.n1811 VDAC_P.t616 1.1255
R18159 VDAC_P.n1812 VDAC_P.t794 1.1255
R18160 VDAC_P.n1813 VDAC_P.t195 1.1255
R18161 VDAC_P.n1814 VDAC_P.t682 1.1255
R18162 VDAC_P.n1815 VDAC_P.t1153 1.1255
R18163 VDAC_P.n1816 VDAC_P.t1711 1.1255
R18164 VDAC_P.n1817 VDAC_P.t2042 1.1255
R18165 VDAC_P.n89 VDAC_P.t718 1.1255
R18166 VDAC_P.n1818 VDAC_P.t18 1.1255
R18167 VDAC_P.n1819 VDAC_P.t1194 1.1255
R18168 VDAC_P.n1820 VDAC_P.t2059 1.1255
R18169 VDAC_P.n1821 VDAC_P.t760 1.1255
R18170 VDAC_P.n1822 VDAC_P.t1686 1.1255
R18171 VDAC_P.n1823 VDAC_P.t36 1.1255
R18172 VDAC_P.n1824 VDAC_P.t1482 1.1255
R18173 VDAC_P.n1825 VDAC_P.t1223 1.1255
R18174 VDAC_P.n1826 VDAC_P.t1254 1.1255
R18175 VDAC_P.n1827 VDAC_P.t163 1.1255
R18176 VDAC_P.n1828 VDAC_P.t128 1.1255
R18177 VDAC_P.n1829 VDAC_P.t1966 1.1255
R18178 VDAC_P.n1830 VDAC_P.t1459 1.1255
R18179 VDAC_P.n1831 VDAC_P.t1681 1.1255
R18180 VDAC_P.n1832 VDAC_P.t1367 1.1255
R18181 VDAC_P.n1833 VDAC_P.t62 1.1255
R18182 VDAC_P.n1834 VDAC_P.t2029 1.1255
R18183 VDAC_P.n1835 VDAC_P.t1328 1.1255
R18184 VDAC_P.n1836 VDAC_P.t1826 1.1255
R18185 VDAC_P.n1837 VDAC_P.t916 1.1255
R18186 VDAC_P.n1838 VDAC_P.t710 1.1255
R18187 VDAC_P.n1839 VDAC_P.t1740 1.1255
R18188 VDAC_P.n1840 VDAC_P.t1178 1.1255
R18189 VDAC_P.n1841 VDAC_P.t2102 1.1255
R18190 VDAC_P.n1842 VDAC_P.t1464 1.1255
R18191 VDAC_P.n1843 VDAC_P.t1890 1.1255
R18192 VDAC_P.n1844 VDAC_P.t375 1.1255
R18193 VDAC_P.n1845 VDAC_P.t746 1.1255
R18194 VDAC_P.n1846 VDAC_P.t1317 1.1255
R18195 VDAC_P.n1847 VDAC_P.t1242 1.1255
R18196 VDAC_P.n1848 VDAC_P.t295 1.1255
R18197 VDAC_P.n1849 VDAC_P.t1667 1.1255
R18198 VDAC_P.n1850 VDAC_P.t990 1.1255
R18199 VDAC_P.n1851 VDAC_P.t1451 1.1255
R18200 VDAC_P.n1852 VDAC_P.t497 1.1255
R18201 VDAC_P.n1853 VDAC_P.t1343 1.1255
R18202 VDAC_P.n1854 VDAC_P.t471 1.1255
R18203 VDAC_P.n1855 VDAC_P.t97 1.1255
R18204 VDAC_P.n1856 VDAC_P.t861 1.1255
R18205 VDAC_P.n1857 VDAC_P.t220 1.1255
R18206 VDAC_P.n1858 VDAC_P.t1567 1.1255
R18207 VDAC_P.n1859 VDAC_P.t2123 1.1255
R18208 VDAC_P.n1860 VDAC_P.t1760 1.1255
R18209 VDAC_P.n1861 VDAC_P.t1913 1.1255
R18210 VDAC_P.n1862 VDAC_P.t900 1.1255
R18211 VDAC_P.n1863 VDAC_P.t814 1.1255
R18212 VDAC_P.n1864 VDAC_P.t1644 1.1255
R18213 VDAC_P.n1865 VDAC_P.t598 1.1255
R18214 VDAC_P.n1866 VDAC_P.t604 1.1255
R18215 VDAC_P.n1867 VDAC_P.t952 1.1255
R18216 VDAC_P.n1868 VDAC_P.t1882 1.1255
R18217 VDAC_P.n1869 VDAC_P.t728 1.1255
R18218 VDAC_P.n1870 VDAC_P.t842 1.1255
R18219 VDAC_P.n1871 VDAC_P.t1313 1.1255
R18220 VDAC_P.n1872 VDAC_P.t330 1.1255
R18221 VDAC_P.n1873 VDAC_P.t617 1.1255
R18222 VDAC_P.n1874 VDAC_P.t520 1.1255
R18223 VDAC_P.n1875 VDAC_P.t986 1.1255
R18224 VDAC_P.n1876 VDAC_P.t793 1.1255
R18225 VDAC_P.n1877 VDAC_P.t134 1.1255
R18226 VDAC_P.n1878 VDAC_P.t1341 1.1255
R18227 VDAC_P.n1879 VDAC_P.t145 1.1255
R18228 VDAC_P.n1880 VDAC_P.t1237 1.1255
R18229 VDAC_P.n88 VDAC_P.t241 1.1255
R18230 VDAC_P.n1881 VDAC_P.t542 1.1255
R18231 VDAC_P.n1882 VDAC_P.t829 1.1255
R18232 VDAC_P.n1883 VDAC_P.t1878 1.1255
R18233 VDAC_P.n1884 VDAC_P.t373 1.1255
R18234 VDAC_P.n1885 VDAC_P.t1865 1.1255
R18235 VDAC_P.n1886 VDAC_P.t669 1.1255
R18236 VDAC_P.n1887 VDAC_P.t895 1.1255
R18237 VDAC_P.n1888 VDAC_P.t1980 1.1255
R18238 VDAC_P.n1889 VDAC_P.t1659 1.1255
R18239 VDAC_P.n1890 VDAC_P.t549 1.1255
R18240 VDAC_P.n1891 VDAC_P.t1443 1.1255
R18241 VDAC_P.n1892 VDAC_P.t2009 1.1255
R18242 VDAC_P.n1893 VDAC_P.t640 1.1255
R18243 VDAC_P.n1894 VDAC_P.t958 1.1255
R18244 VDAC_P.n1895 VDAC_P.t721 1.1255
R18245 VDAC_P.n1896 VDAC_P.t1985 1.1255
R18246 VDAC_P.n1897 VDAC_P.t1315 1.1255
R18247 VDAC_P.n1898 VDAC_P.t1765 1.1255
R18248 VDAC_P.n1899 VDAC_P.t1412 1.1255
R18249 VDAC_P.n1900 VDAC_P.t437 1.1255
R18250 VDAC_P.n1901 VDAC_P.t1073 1.1255
R18251 VDAC_P.n1902 VDAC_P.t411 1.1255
R18252 VDAC_P.n1903 VDAC_P.t2013 1.1255
R18253 VDAC_P.n1904 VDAC_P.t184 1.1255
R18254 VDAC_P.n1905 VDAC_P.t913 1.1255
R18255 VDAC_P.n1906 VDAC_P.t852 1.1255
R18256 VDAC_P.n1907 VDAC_P.t1362 1.1255
R18257 VDAC_P.n1908 VDAC_P.t860 1.1255
R18258 VDAC_P.n1909 VDAC_P.t1154 1.1255
R18259 VDAC_P.n1910 VDAC_P.t2041 1.1255
R18260 VDAC_P.n1911 VDAC_P.t712 1.1255
R18261 VDAC_P.n1912 VDAC_P.t1862 1.1255
R18262 VDAC_P.n1913 VDAC_P.t964 1.1255
R18263 VDAC_P.n1914 VDAC_P.t1430 1.1255
R18264 VDAC_P.n1915 VDAC_P.t1195 1.1255
R18265 VDAC_P.n1916 VDAC_P.t1206 1.1255
R18266 VDAC_P.n1917 VDAC_P.t29 1.1255
R18267 VDAC_P.n1918 VDAC_P.t776 1.1255
R18268 VDAC_P.n1919 VDAC_P.t502 1.1255
R18269 VDAC_P.n1920 VDAC_P.t1433 1.1255
R18270 VDAC_P.n1921 VDAC_P.t434 1.1255
R18271 VDAC_P.n1922 VDAC_P.t717 1.1255
R18272 VDAC_P.n1923 VDAC_P.t1863 1.1255
R18273 VDAC_P.n1924 VDAC_P.t1203 1.1255
R18274 VDAC_P.n1925 VDAC_P.t1661 1.1255
R18275 VDAC_P.n1926 VDAC_P.t1916 1.1255
R18276 VDAC_P.n1927 VDAC_P.t791 1.1255
R18277 VDAC_P.n1928 VDAC_P.t1019 1.1255
R18278 VDAC_P.n1929 VDAC_P.t381 1.1255
R18279 VDAC_P.n1930 VDAC_P.t495 1.1255
R18280 VDAC_P.n1931 VDAC_P.t228 1.1255
R18281 VDAC_P.n1932 VDAC_P.t469 1.1255
R18282 VDAC_P.n1933 VDAC_P.t204 1.1255
R18283 VDAC_P.n1934 VDAC_P.t1146 1.1255
R18284 VDAC_P.n1935 VDAC_P.t531 1.1255
R18285 VDAC_P.n1936 VDAC_P.t1824 1.1255
R18286 VDAC_P.n1937 VDAC_P.t1925 1.1255
R18287 VDAC_P.n1938 VDAC_P.t1876 1.1255
R18288 VDAC_P.n1939 VDAC_P.t1630 1.1255
R18289 VDAC_P.n1940 VDAC_P.t1900 1.1255
R18290 VDAC_P.n1941 VDAC_P.t1202 1.1255
R18291 VDAC_P.n1942 VDAC_P.t1189 1.1255
R18292 VDAC_P.n1943 VDAC_P.t1928 1.1255
R18293 VDAC_P.n87 VDAC_P.t1408 1.1255
R18294 VDAC_P.n86 VDAC_P.t1829 1.1255
R18295 VDAC_P.n85 VDAC_P.t980 1.1255
R18296 VDAC_P.n84 VDAC_P.t875 1.1255
R18297 VDAC_P.n83 VDAC_P.t26 1.1255
R18298 VDAC_P.n82 VDAC_P.t272 1.1255
R18299 VDAC_P.n81 VDAC_P.t1049 1.1255
R18300 VDAC_P.n80 VDAC_P.t1544 1.1255
R18301 VDAC_P.n79 VDAC_P.t870 1.1255
R18302 VDAC_P.n78 VDAC_P.t560 1.1255
R18303 VDAC_P.n77 VDAC_P.t1510 1.1255
R18304 VDAC_P.n76 VDAC_P.t444 1.1255
R18305 VDAC_P.n75 VDAC_P.t1278 1.1255
R18306 VDAC_P.n74 VDAC_P.t1123 1.1255
R18307 VDAC_P.n73 VDAC_P.t169 1.1255
R18308 VDAC_P.n72 VDAC_P.t819 1.1255
R18309 VDAC_P.n71 VDAC_P.t12 1.1255
R18310 VDAC_P.n70 VDAC_P.t397 1.1255
R18311 VDAC_P.n69 VDAC_P.t1955 1.1255
R18312 VDAC_P.n68 VDAC_P.t120 1.1255
R18313 VDAC_P.n67 VDAC_P.t1847 1.1255
R18314 VDAC_P.n66 VDAC_P.t1204 1.1255
R18315 VDAC_P.n65 VDAC_P.t885 1.1255
R18316 VDAC_P.n64 VDAC_P.t1276 1.1255
R18317 VDAC_P.n63 VDAC_P.t536 1.1255
R18318 VDAC_P.n62 VDAC_P.t1989 1.1255
R18319 VDAC_P.n61 VDAC_P.t1640 1.1255
R18320 VDAC_P.n60 VDAC_P.t82 1.1255
R18321 VDAC_P.n59 VDAC_P.t740 1.1255
R18322 VDAC_P.n58 VDAC_P.t1550 1.1255
R18323 VDAC_P.n57 VDAC_P.t300 1.1255
R18324 VDAC_P.n56 VDAC_P.t162 1.1255
R18325 VDAC_P.n55 VDAC_P.t1145 1.1255
R18326 VDAC_P.n54 VDAC_P.t1752 1.1255
R18327 VDAC_P.n53 VDAC_P.t474 1.1255
R18328 VDAC_P.n52 VDAC_P.t1381 1.1255
R18329 VDAC_P.n51 VDAC_P.t810 1.1255
R18330 VDAC_P.n50 VDAC_P.t67 1.1255
R18331 VDAC_P.n49 VDAC_P.t1162 1.1255
R18332 VDAC_P.n48 VDAC_P.t171 1.1255
R18333 VDAC_P.n47 VDAC_P.t1627 1.1255
R18334 VDAC_P.n46 VDAC_P.t2038 1.1255
R18335 VDAC_P.n45 VDAC_P.t225 1.1255
R18336 VDAC_P.n44 VDAC_P.t535 1.1255
R18337 VDAC_P.n43 VDAC_P.t1385 1.1255
R18338 VDAC_P.n42 VDAC_P.t255 1.1255
R18339 VDAC_P.n41 VDAC_P.t2052 1.1255
R18340 VDAC_P.n40 VDAC_P.t455 1.1255
R18341 VDAC_P.n39 VDAC_P.t1212 1.1255
R18342 VDAC_P.n38 VDAC_P.t1635 1.1255
R18343 VDAC_P.n37 VDAC_P.t285 1.1255
R18344 VDAC_P.n36 VDAC_P.t824 1.1255
R18345 VDAC_P.n35 VDAC_P.t517 1.1255
R18346 VDAC_P.n34 VDAC_P.t1152 1.1255
R18347 VDAC_P.n33 VDAC_P.t786 1.1255
R18348 VDAC_P.n32 VDAC_P.t1100 1.1255
R18349 VDAC_P.n31 VDAC_P.t670 1.1255
R18350 VDAC_P.n30 VDAC_P.t2117 1.1255
R18351 VDAC_P.n29 VDAC_P.t1744 1.1255
R18352 VDAC_P.n28 VDAC_P.t1026 1.1255
R18353 VDAC_P.n27 VDAC_P.t1272 1.1255
R18354 VDAC_P.n26 VDAC_P.t1586 1.1255
R18355 VDAC_P.n25 VDAC_P.t1377 1.1255
R18356 VDAC_P.n24 VDAC_P.t694 1.1255
R18357 VDAC_P.n23 VDAC_P.t599 1.1255
R18358 VDAC_P.n1944 VDAC_P.t1918 1.1255
R18359 VDAC_P.n1945 VDAC_P.t41 1.1255
R18360 VDAC_P.n1946 VDAC_P.t765 1.1255
R18361 VDAC_P.n1947 VDAC_P.t671 1.1255
R18362 VDAC_P.n1948 VDAC_P.t153 1.1255
R18363 VDAC_P.n1949 VDAC_P.t479 1.1255
R18364 VDAC_P.n1950 VDAC_P.t1632 1.1255
R18365 VDAC_P.n1951 VDAC_P.t1652 1.1255
R18366 VDAC_P.n1952 VDAC_P.t16 1.1255
R18367 VDAC_P.n1953 VDAC_P.t770 1.1255
R18368 VDAC_P.n1954 VDAC_P.t570 1.1255
R18369 VDAC_P.n1955 VDAC_P.t663 1.1255
R18370 VDAC_P.n1956 VDAC_P.t567 1.1255
R18371 VDAC_P.n1957 VDAC_P.t1794 1.1255
R18372 VDAC_P.n1958 VDAC_P.t831 1.1255
R18373 VDAC_P.n1959 VDAC_P.t1439 1.1255
R18374 VDAC_P.n1960 VDAC_P.t1669 1.1255
R18375 VDAC_P.n1961 VDAC_P.t753 1.1255
R18376 VDAC_P.n1962 VDAC_P.t1287 1.1255
R18377 VDAC_P.n1963 VDAC_P.t1990 1.1255
R18378 VDAC_P.n1964 VDAC_P.t1207 1.1255
R18379 VDAC_P.n1965 VDAC_P.t1976 1.1255
R18380 VDAC_P.n1966 VDAC_P.t1382 1.1255
R18381 VDAC_P.n1967 VDAC_P.t1770 1.1255
R18382 VDAC_P.n1968 VDAC_P.t100 1.1255
R18383 VDAC_P.n1969 VDAC_P.t112 1.1255
R18384 VDAC_P.n1970 VDAC_P.t1779 1.1255
R18385 VDAC_P.n1971 VDAC_P.t999 1.1255
R18386 VDAC_P.n1972 VDAC_P.t924 1.1255
R18387 VDAC_P.n1973 VDAC_P.t737 1.1255
R18388 VDAC_P.n1974 VDAC_P.t1938 1.1255
R18389 VDAC_P.n1975 VDAC_P.t79 1.1255
R18390 VDAC_P.n1976 VDAC_P.t1091 1.1255
R18391 VDAC_P.n1977 VDAC_P.t1226 1.1255
R18392 VDAC_P.n1978 VDAC_P.t1311 1.1255
R18393 VDAC_P.n1979 VDAC_P.t382 1.1255
R18394 VDAC_P.n1980 VDAC_P.t996 1.1255
R18395 VDAC_P.n1981 VDAC_P.t954 1.1255
R18396 VDAC_P.n1982 VDAC_P.t1424 1.1255
R18397 VDAC_P.n1983 VDAC_P.t2090 1.1255
R18398 VDAC_P.n1984 VDAC_P.t1166 1.1255
R18399 VDAC_P.n1985 VDAC_P.t812 1.1255
R18400 VDAC_P.n1986 VDAC_P.t702 1.1255
R18401 VDAC_P.n1987 VDAC_P.t452 1.1255
R18402 VDAC_P.n1988 VDAC_P.t1909 1.1255
R18403 VDAC_P.n1989 VDAC_P.t664 1.1255
R18404 VDAC_P.n1990 VDAC_P.t1023 1.1255
R18405 VDAC_P.n1991 VDAC_P.t1102 1.1255
R18406 VDAC_P.n1992 VDAC_P.t1075 1.1255
R18407 VDAC_P.n1993 VDAC_P.t439 1.1255
R18408 VDAC_P.n1994 VDAC_P.t1460 1.1255
R18409 VDAC_P.n1995 VDAC_P.t1875 1.1255
R18410 VDAC_P.n1996 VDAC_P.t675 1.1255
R18411 VDAC_P.n1997 VDAC_P.t1903 1.1255
R18412 VDAC_P.n1998 VDAC_P.t1449 1.1255
R18413 VDAC_P.n1999 VDAC_P.t454 1.1255
R18414 VDAC_P.n2000 VDAC_P.t795 1.1255
R18415 VDAC_P.n2001 VDAC_P.t561 1.1255
R18416 VDAC_P.n2002 VDAC_P.t847 1.1255
R18417 VDAC_P.n2003 VDAC_P.t619 1.1255
R18418 VDAC_P.n2004 VDAC_P.t386 1.1255
R18419 VDAC_P.n2005 VDAC_P.t1413 1.1255
R18420 VDAC_P.n2006 VDAC_P.t846 1.1255
R18421 VDAC_P.n2007 VDAC_P.t1456 1.1255
R18422 VDAC_P.n2008 VDAC_P.t2098 1.1255
R18423 VDAC_P.n2009 VDAC_P.t1896 1.1255
R18424 VDAC_P.n2010 VDAC_P.t37 1.1255
R18425 VDAC_P.n2011 VDAC_P.t1386 1.1255
R18426 VDAC_P.n2012 VDAC_P.t876 1.1255
R18427 VDAC_P.n2013 VDAC_P.t1614 1.1255
R18428 VDAC_P.n2014 VDAC_P.t1320 1.1255
R18429 VDAC_P.n2015 VDAC_P.t2027 1.1255
R18430 VDAC_P.n2016 VDAC_P.t1784 1.1255
R18431 VDAC_P.n2017 VDAC_P.t2133 1.1255
R18432 VDAC_P.n2018 VDAC_P.t1330 1.1255
R18433 VDAC_P.n2019 VDAC_P.t332 1.1255
R18434 VDAC_P.n2020 VDAC_P.t1781 1.1255
R18435 VDAC_P.n2021 VDAC_P.t1192 1.1255
R18436 VDAC_P.n2022 VDAC_P.t1885 1.1255
R18437 VDAC_P.n2023 VDAC_P.t203 1.1255
R18438 VDAC_P.n2024 VDAC_P.t787 1.1255
R18439 VDAC_P.n2025 VDAC_P.t27 1.1255
R18440 VDAC_P.n2026 VDAC_P.t1944 1.1255
R18441 VDAC_P.n2027 VDAC_P.t611 1.1255
R18442 VDAC_P.n2028 VDAC_P.t378 1.1255
R18443 VDAC_P.n2029 VDAC_P.t665 1.1255
R18444 VDAC_P.n2030 VDAC_P.t1642 1.1255
R18445 VDAC_P.n2031 VDAC_P.t1392 1.1255
R18446 VDAC_P.n2032 VDAC_P.t1866 1.1255
R18447 VDAC_P.n2033 VDAC_P.t256 1.1255
R18448 VDAC_P.n2034 VDAC_P.t1756 1.1255
R18449 VDAC_P.n2035 VDAC_P.t194 1.1255
R18450 VDAC_P.n2036 VDAC_P.t396 1.1255
R18451 VDAC_P.n2037 VDAC_P.t806 1.1255
R18452 VDAC_P.n2038 VDAC_P.t1264 1.1255
R18453 VDAC_P.n2039 VDAC_P.t1465 1.1255
R18454 VDAC_P.n2040 VDAC_P.t1342 1.1255
R18455 VDAC_P.n2041 VDAC_P.t2039 1.1255
R18456 VDAC_P.n2042 VDAC_P.t1030 1.1255
R18457 VDAC_P.n2043 VDAC_P.t1796 1.1255
R18458 VDAC_P.n2044 VDAC_P.t1369 1.1255
R18459 VDAC_P.n2045 VDAC_P.t1150 1.1255
R18460 VDAC_P.n2046 VDAC_P.t1939 1.1255
R18461 VDAC_P.n2047 VDAC_P.t579 1.1255
R18462 VDAC_P.n2048 VDAC_P.t656 1.1255
R18463 VDAC_P.n2049 VDAC_P.t208 1.1255
R18464 VDAC_P.n2050 VDAC_P.t1173 1.1255
R18465 VDAC_P.n2051 VDAC_P.t979 1.1255
R18466 VDAC_P.n2052 VDAC_P.t1954 1.1255
R18467 VDAC_P.n2053 VDAC_P.t893 1.1255
R18468 VDAC_P.n2054 VDAC_P.t1266 1.1255
R18469 VDAC_P.n2055 VDAC_P.t1421 1.1255
R18470 VDAC_P.n2056 VDAC_P.t1148 1.1255
R18471 VDAC_P.n2057 VDAC_P.t61 1.1255
R18472 VDAC_P.n2058 VDAC_P.t1851 1.1255
R18473 VDAC_P.n2059 VDAC_P.t1470 1.1255
R18474 VDAC_P.n2060 VDAC_P.t775 1.1255
R18475 VDAC_P.n2061 VDAC_P.t1004 1.1255
R18476 VDAC_P.n2062 VDAC_P.t1185 1.1255
R18477 VDAC_P.n2063 VDAC_P.t989 1.1255
R18478 VDAC_P.n2064 VDAC_P.t1646 1.1255
R18479 VDAC_P.n2065 VDAC_P.t425 1.1255
R18480 VDAC_P.n2066 VDAC_P.t1844 1.1255
R18481 VDAC_P.n2067 VDAC_P.t653 1.1255
R18482 VDAC_P.n2068 VDAC_P.t2043 1.1255
R18483 VDAC_P.n2069 VDAC_P.t1842 1.1255
R18484 VDAC_P.n2070 VDAC_P.t709 1.1255
R18485 VDAC_P.n2071 VDAC_P.t714 1.1255
R18486 VDAC_P.n2072 VDAC_P.t343 1.1255
R18487 VDAC_P.n2073 VDAC_P.t318 1.1255
R18488 VDAC_P.n2074 VDAC_P.t2110 1.1255
R18489 VDAC_P.n2075 VDAC_P.t781 1.1255
R18490 VDAC_P.n2076 VDAC_P.t966 1.1255
R18491 VDAC_P.n2077 VDAC_P.t725 1.1255
R18492 VDAC_P.n2078 VDAC_P.t1877 1.1255
R18493 VDAC_P.n2079 VDAC_P.t109 1.1255
R18494 VDAC_P.n2080 VDAC_P.t1771 1.1255
R18495 VDAC_P.n2081 VDAC_P.t1105 1.1255
R18496 VDAC_P.n2082 VDAC_P.t851 1.1255
R18497 VDAC_P.n2083 VDAC_P.t2125 1.1255
R18498 VDAC_P.n2084 VDAC_P.t832 1.1255
R18499 VDAC_P.n2085 VDAC_P.t890 1.1255
R18500 VDAC_P.n2086 VDAC_P.t1461 1.1255
R18501 VDAC_P.n2087 VDAC_P.t1546 1.1255
R18502 VDAC_P.n2088 VDAC_P.t1249 1.1255
R18503 VDAC_P.n2089 VDAC_P.t917 1.1255
R18504 VDAC_P.n2090 VDAC_P.t1143 1.1255
R18505 VDAC_P.n2091 VDAC_P.t1597 1.1255
R18506 VDAC_P.n2092 VDAC_P.t2030 1.1255
R18507 VDAC_P.n2093 VDAC_P.t1491 1.1255
R18508 VDAC_P.n2094 VDAC_P.t1945 1.1255
R18509 VDAC_P.n2095 VDAC_P.t651 1.1255
R18510 VDAC_P.n2096 VDAC_P.t1835 1.1255
R18511 VDAC_P.n2097 VDAC_P.t1092 1.1255
R18512 VDAC_P.n2098 VDAC_P.t1625 1.1255
R18513 VDAC_P.n2099 VDAC_P.t1052 1.1255
R18514 VDAC_P.n2100 VDAC_P.t1519 1.1255
R18515 VDAC_P.n2101 VDAC_P.t515 1.1255
R18516 VDAC_P.n2102 VDAC_P.t800 1.1255
R18517 VDAC_P.n2103 VDAC_P.t257 1.1255
R18518 VDAC_P.n2104 VDAC_P.t1364 1.1255
R18519 VDAC_P.n2105 VDAC_P.t662 1.1255
R18520 VDAC_P.n2106 VDAC_P.t1788 1.1255
R18521 VDAC_P.n2107 VDAC_P.t2128 1.1255
R18522 VDAC_P.n2108 VDAC_P.t275 1.1255
R18523 VDAC_P.n2109 VDAC_P.t1712 1.1255
R18524 VDAC_P.n2110 VDAC_P.t1782 1.1255
R18525 VDAC_P.n2111 VDAC_P.t1144 1.1255
R18526 VDAC_P.n2112 VDAC_P.t1742 1.1255
R18527 VDAC_P.n2113 VDAC_P.t1349 1.1255
R18528 VDAC_P.n2114 VDAC_P.t666 1.1255
R18529 VDAC_P.n2115 VDAC_P.t167 1.1255
R18530 VDAC_P.n2116 VDAC_P.t863 1.1255
R18531 VDAC_P.n2117 VDAC_P.t2014 1.1255
R18532 VDAC_P.n2118 VDAC_P.t1487 1.1255
R18533 VDAC_P.n2119 VDAC_P.t470 1.1255
R18534 VDAC_P.n2120 VDAC_P.t701 1.1255
R18535 VDAC_P.n2121 VDAC_P.t929 1.1255
R18536 VDAC_P.n2122 VDAC_P.t647 1.1255
R18537 VDAC_P.n2123 VDAC_P.t81 1.1255
R18538 VDAC_P.n2124 VDAC_P.t1564 1.1255
R18539 VDAC_P.n2125 VDAC_P.t1517 1.1255
R18540 VDAC_P.n2126 VDAC_P.t2073 1.1255
R18541 VDAC_P.n2127 VDAC_P.t371 1.1255
R18542 VDAC_P.n2128 VDAC_P.t943 1.1255
R18543 VDAC_P.n2129 VDAC_P.t1104 1.1255
R18544 VDAC_P.n2130 VDAC_P.t1753 1.1255
R18545 VDAC_P.n2131 VDAC_P.t892 1.1255
R18546 VDAC_P.n2132 VDAC_P.t342 1.1255
R18547 VDAC_P.n2133 VDAC_P.t2101 1.1255
R18548 VDAC_P.n2134 VDAC_P.t1696 1.1255
R18549 VDAC_P.n11 VDAC_P.n10 0.733109
R18550 VDAC_P.n12 VDAC_P.n11 0.733109
R18551 VDAC_P.n4 VDAC_P.n3 0.733109
R18552 VDAC_P.n5 VDAC_P.n4 0.733109
R18553 VDAC_P.n1 VDAC_P.n0 0.733109
R18554 VDAC_P.n2 VDAC_P.n1 0.733109
R18555 VDAC_P.n13 VDAC_P.n12 0.675138
R18556 VDAC_P.n8 VDAC_P.n7 0.589359
R18557 VDAC_P.n9 VDAC_P.n8 0.589359
R18558 VDAC_P.n6 VDAC_P.n5 0.491804
R18559 VDAC_P.n21 VDAC_P.n20 0.21925
R18560 VDAC_P.n1944 VDAC_P.n23 0.204167
R18561 VDAC_P.n1945 VDAC_P.n1944 0.204167
R18562 VDAC_P.n1946 VDAC_P.n1945 0.204167
R18563 VDAC_P.n1947 VDAC_P.n1946 0.204167
R18564 VDAC_P.n1948 VDAC_P.n1947 0.204167
R18565 VDAC_P.n1949 VDAC_P.n1948 0.204167
R18566 VDAC_P.n1950 VDAC_P.n1949 0.204167
R18567 VDAC_P.n1951 VDAC_P.n1950 0.204167
R18568 VDAC_P.n1952 VDAC_P.n1951 0.204167
R18569 VDAC_P.n1953 VDAC_P.n1952 0.204167
R18570 VDAC_P.n1954 VDAC_P.n1953 0.204167
R18571 VDAC_P.n1955 VDAC_P.n1954 0.204167
R18572 VDAC_P.n1956 VDAC_P.n1955 0.204167
R18573 VDAC_P.n1957 VDAC_P.n1956 0.204167
R18574 VDAC_P.n1958 VDAC_P.n1957 0.204167
R18575 VDAC_P.n1959 VDAC_P.n1958 0.204167
R18576 VDAC_P.n1960 VDAC_P.n1959 0.204167
R18577 VDAC_P.n1961 VDAC_P.n1960 0.204167
R18578 VDAC_P.n1962 VDAC_P.n1961 0.204167
R18579 VDAC_P.n1963 VDAC_P.n1962 0.204167
R18580 VDAC_P.n1964 VDAC_P.n1963 0.204167
R18581 VDAC_P.n1965 VDAC_P.n1964 0.204167
R18582 VDAC_P.n1966 VDAC_P.n1965 0.204167
R18583 VDAC_P.n1967 VDAC_P.n1966 0.204167
R18584 VDAC_P.n1968 VDAC_P.n1967 0.204167
R18585 VDAC_P.n1969 VDAC_P.n1968 0.204167
R18586 VDAC_P.n1970 VDAC_P.n1969 0.204167
R18587 VDAC_P.n1971 VDAC_P.n1970 0.204167
R18588 VDAC_P.n1972 VDAC_P.n1971 0.204167
R18589 VDAC_P.n2040 VDAC_P.n2039 0.204167
R18590 VDAC_P.n2041 VDAC_P.n2040 0.204167
R18591 VDAC_P.n2042 VDAC_P.n2041 0.204167
R18592 VDAC_P.n2043 VDAC_P.n2042 0.204167
R18593 VDAC_P.n2044 VDAC_P.n2043 0.204167
R18594 VDAC_P.n2045 VDAC_P.n2044 0.204167
R18595 VDAC_P.n2046 VDAC_P.n2045 0.204167
R18596 VDAC_P.n2047 VDAC_P.n2046 0.204167
R18597 VDAC_P.n2048 VDAC_P.n2047 0.204167
R18598 VDAC_P.n2049 VDAC_P.n2048 0.204167
R18599 VDAC_P.n2050 VDAC_P.n2049 0.204167
R18600 VDAC_P.n2051 VDAC_P.n2050 0.204167
R18601 VDAC_P.n2052 VDAC_P.n2051 0.204167
R18602 VDAC_P.n2053 VDAC_P.n2052 0.204167
R18603 VDAC_P.n2054 VDAC_P.n2053 0.204167
R18604 VDAC_P.n2055 VDAC_P.n2054 0.204167
R18605 VDAC_P.n2056 VDAC_P.n2055 0.204167
R18606 VDAC_P.n2057 VDAC_P.n2056 0.204167
R18607 VDAC_P.n2058 VDAC_P.n2057 0.204167
R18608 VDAC_P.n2059 VDAC_P.n2058 0.204167
R18609 VDAC_P.n2060 VDAC_P.n2059 0.204167
R18610 VDAC_P.n2061 VDAC_P.n2060 0.204167
R18611 VDAC_P.n2062 VDAC_P.n2061 0.204167
R18612 VDAC_P.n2063 VDAC_P.n2062 0.204167
R18613 VDAC_P.n2064 VDAC_P.n2063 0.204167
R18614 VDAC_P.n2065 VDAC_P.n2064 0.204167
R18615 VDAC_P.n2066 VDAC_P.n2065 0.204167
R18616 VDAC_P.n2067 VDAC_P.n2066 0.204167
R18617 VDAC_P.n2068 VDAC_P.n2067 0.204167
R18618 VDAC_P.n21 VDAC_P.n17 0.188
R18619 VDAC_P.n117 VDAC_P.n116 0.180667
R18620 VDAC_P.n118 VDAC_P.n117 0.180667
R18621 VDAC_P.n119 VDAC_P.n118 0.180667
R18622 VDAC_P.n120 VDAC_P.n119 0.180667
R18623 VDAC_P.n121 VDAC_P.n120 0.180667
R18624 VDAC_P.n122 VDAC_P.n121 0.180667
R18625 VDAC_P.n123 VDAC_P.n122 0.180667
R18626 VDAC_P.n124 VDAC_P.n123 0.180667
R18627 VDAC_P.n125 VDAC_P.n124 0.180667
R18628 VDAC_P.n126 VDAC_P.n125 0.180667
R18629 VDAC_P.n127 VDAC_P.n126 0.180667
R18630 VDAC_P.n128 VDAC_P.n127 0.180667
R18631 VDAC_P.n129 VDAC_P.n128 0.180667
R18632 VDAC_P.n130 VDAC_P.n129 0.180667
R18633 VDAC_P.n131 VDAC_P.n130 0.180667
R18634 VDAC_P.n132 VDAC_P.n131 0.180667
R18635 VDAC_P.n133 VDAC_P.n132 0.180667
R18636 VDAC_P.n134 VDAC_P.n133 0.180667
R18637 VDAC_P.n135 VDAC_P.n134 0.180667
R18638 VDAC_P.n136 VDAC_P.n135 0.180667
R18639 VDAC_P.n137 VDAC_P.n136 0.180667
R18640 VDAC_P.n138 VDAC_P.n137 0.180667
R18641 VDAC_P.n139 VDAC_P.n138 0.180667
R18642 VDAC_P.n140 VDAC_P.n139 0.180667
R18643 VDAC_P.n141 VDAC_P.n140 0.180667
R18644 VDAC_P.n142 VDAC_P.n141 0.180667
R18645 VDAC_P.n143 VDAC_P.n142 0.180667
R18646 VDAC_P.n144 VDAC_P.n143 0.180667
R18647 VDAC_P.n145 VDAC_P.n144 0.180667
R18648 VDAC_P.n146 VDAC_P.n145 0.180667
R18649 VDAC_P.n147 VDAC_P.n146 0.180667
R18650 VDAC_P.n148 VDAC_P.n147 0.180667
R18651 VDAC_P.n149 VDAC_P.n148 0.180667
R18652 VDAC_P.n150 VDAC_P.n149 0.180667
R18653 VDAC_P.n151 VDAC_P.n150 0.180667
R18654 VDAC_P.n152 VDAC_P.n151 0.180667
R18655 VDAC_P.n153 VDAC_P.n152 0.180667
R18656 VDAC_P.n154 VDAC_P.n153 0.180667
R18657 VDAC_P.n155 VDAC_P.n154 0.180667
R18658 VDAC_P.n156 VDAC_P.n155 0.180667
R18659 VDAC_P.n157 VDAC_P.n156 0.180667
R18660 VDAC_P.n158 VDAC_P.n157 0.180667
R18661 VDAC_P.n159 VDAC_P.n158 0.180667
R18662 VDAC_P.n160 VDAC_P.n159 0.180667
R18663 VDAC_P.n161 VDAC_P.n160 0.180667
R18664 VDAC_P.n162 VDAC_P.n161 0.180667
R18665 VDAC_P.n163 VDAC_P.n162 0.180667
R18666 VDAC_P.n164 VDAC_P.n163 0.180667
R18667 VDAC_P.n165 VDAC_P.n164 0.180667
R18668 VDAC_P.n166 VDAC_P.n165 0.180667
R18669 VDAC_P.n167 VDAC_P.n166 0.180667
R18670 VDAC_P.n168 VDAC_P.n167 0.180667
R18671 VDAC_P.n169 VDAC_P.n168 0.180667
R18672 VDAC_P.n170 VDAC_P.n169 0.180667
R18673 VDAC_P.n171 VDAC_P.n170 0.180667
R18674 VDAC_P.n172 VDAC_P.n171 0.180667
R18675 VDAC_P.n173 VDAC_P.n172 0.180667
R18676 VDAC_P.n174 VDAC_P.n173 0.180667
R18677 VDAC_P.n175 VDAC_P.n174 0.180667
R18678 VDAC_P.n176 VDAC_P.n175 0.180667
R18679 VDAC_P.n177 VDAC_P.n176 0.180667
R18680 VDAC_P.n178 VDAC_P.n177 0.180667
R18681 VDAC_P.n179 VDAC_P.n178 0.180667
R18682 VDAC_P.n180 VDAC_P.n115 0.180667
R18683 VDAC_P.n181 VDAC_P.n180 0.180667
R18684 VDAC_P.n182 VDAC_P.n181 0.180667
R18685 VDAC_P.n183 VDAC_P.n182 0.180667
R18686 VDAC_P.n184 VDAC_P.n183 0.180667
R18687 VDAC_P.n185 VDAC_P.n184 0.180667
R18688 VDAC_P.n186 VDAC_P.n185 0.180667
R18689 VDAC_P.n187 VDAC_P.n186 0.180667
R18690 VDAC_P.n188 VDAC_P.n187 0.180667
R18691 VDAC_P.n189 VDAC_P.n188 0.180667
R18692 VDAC_P.n190 VDAC_P.n189 0.180667
R18693 VDAC_P.n191 VDAC_P.n190 0.180667
R18694 VDAC_P.n192 VDAC_P.n191 0.180667
R18695 VDAC_P.n193 VDAC_P.n192 0.180667
R18696 VDAC_P.n194 VDAC_P.n193 0.180667
R18697 VDAC_P.n195 VDAC_P.n194 0.180667
R18698 VDAC_P.n196 VDAC_P.n195 0.180667
R18699 VDAC_P.n197 VDAC_P.n196 0.180667
R18700 VDAC_P.n198 VDAC_P.n197 0.180667
R18701 VDAC_P.n199 VDAC_P.n198 0.180667
R18702 VDAC_P.n200 VDAC_P.n199 0.180667
R18703 VDAC_P.n201 VDAC_P.n200 0.180667
R18704 VDAC_P.n202 VDAC_P.n201 0.180667
R18705 VDAC_P.n203 VDAC_P.n202 0.180667
R18706 VDAC_P.n204 VDAC_P.n203 0.180667
R18707 VDAC_P.n205 VDAC_P.n204 0.180667
R18708 VDAC_P.n206 VDAC_P.n205 0.180667
R18709 VDAC_P.n207 VDAC_P.n206 0.180667
R18710 VDAC_P.n208 VDAC_P.n207 0.180667
R18711 VDAC_P.n209 VDAC_P.n208 0.180667
R18712 VDAC_P.n210 VDAC_P.n209 0.180667
R18713 VDAC_P.n211 VDAC_P.n210 0.180667
R18714 VDAC_P.n212 VDAC_P.n211 0.180667
R18715 VDAC_P.n213 VDAC_P.n212 0.180667
R18716 VDAC_P.n214 VDAC_P.n213 0.180667
R18717 VDAC_P.n215 VDAC_P.n214 0.180667
R18718 VDAC_P.n216 VDAC_P.n215 0.180667
R18719 VDAC_P.n217 VDAC_P.n216 0.180667
R18720 VDAC_P.n218 VDAC_P.n217 0.180667
R18721 VDAC_P.n219 VDAC_P.n218 0.180667
R18722 VDAC_P.n220 VDAC_P.n219 0.180667
R18723 VDAC_P.n221 VDAC_P.n220 0.180667
R18724 VDAC_P.n222 VDAC_P.n221 0.180667
R18725 VDAC_P.n223 VDAC_P.n222 0.180667
R18726 VDAC_P.n224 VDAC_P.n223 0.180667
R18727 VDAC_P.n225 VDAC_P.n224 0.180667
R18728 VDAC_P.n226 VDAC_P.n225 0.180667
R18729 VDAC_P.n227 VDAC_P.n226 0.180667
R18730 VDAC_P.n228 VDAC_P.n227 0.180667
R18731 VDAC_P.n229 VDAC_P.n228 0.180667
R18732 VDAC_P.n230 VDAC_P.n229 0.180667
R18733 VDAC_P.n231 VDAC_P.n230 0.180667
R18734 VDAC_P.n232 VDAC_P.n231 0.180667
R18735 VDAC_P.n233 VDAC_P.n232 0.180667
R18736 VDAC_P.n234 VDAC_P.n233 0.180667
R18737 VDAC_P.n235 VDAC_P.n234 0.180667
R18738 VDAC_P.n236 VDAC_P.n235 0.180667
R18739 VDAC_P.n237 VDAC_P.n236 0.180667
R18740 VDAC_P.n238 VDAC_P.n237 0.180667
R18741 VDAC_P.n239 VDAC_P.n238 0.180667
R18742 VDAC_P.n240 VDAC_P.n239 0.180667
R18743 VDAC_P.n241 VDAC_P.n240 0.180667
R18744 VDAC_P.n242 VDAC_P.n241 0.180667
R18745 VDAC_P.n243 VDAC_P.n114 0.180667
R18746 VDAC_P.n244 VDAC_P.n243 0.180667
R18747 VDAC_P.n245 VDAC_P.n244 0.180667
R18748 VDAC_P.n246 VDAC_P.n245 0.180667
R18749 VDAC_P.n247 VDAC_P.n246 0.180667
R18750 VDAC_P.n248 VDAC_P.n247 0.180667
R18751 VDAC_P.n249 VDAC_P.n248 0.180667
R18752 VDAC_P.n250 VDAC_P.n249 0.180667
R18753 VDAC_P.n251 VDAC_P.n250 0.180667
R18754 VDAC_P.n252 VDAC_P.n251 0.180667
R18755 VDAC_P.n253 VDAC_P.n252 0.180667
R18756 VDAC_P.n254 VDAC_P.n253 0.180667
R18757 VDAC_P.n255 VDAC_P.n254 0.180667
R18758 VDAC_P.n256 VDAC_P.n255 0.180667
R18759 VDAC_P.n257 VDAC_P.n256 0.180667
R18760 VDAC_P.n258 VDAC_P.n257 0.180667
R18761 VDAC_P.n259 VDAC_P.n258 0.180667
R18762 VDAC_P.n260 VDAC_P.n259 0.180667
R18763 VDAC_P.n261 VDAC_P.n260 0.180667
R18764 VDAC_P.n262 VDAC_P.n261 0.180667
R18765 VDAC_P.n263 VDAC_P.n262 0.180667
R18766 VDAC_P.n264 VDAC_P.n263 0.180667
R18767 VDAC_P.n265 VDAC_P.n264 0.180667
R18768 VDAC_P.n266 VDAC_P.n265 0.180667
R18769 VDAC_P.n267 VDAC_P.n266 0.180667
R18770 VDAC_P.n268 VDAC_P.n267 0.180667
R18771 VDAC_P.n269 VDAC_P.n268 0.180667
R18772 VDAC_P.n270 VDAC_P.n269 0.180667
R18773 VDAC_P.n271 VDAC_P.n270 0.180667
R18774 VDAC_P.n272 VDAC_P.n271 0.180667
R18775 VDAC_P.n273 VDAC_P.n272 0.180667
R18776 VDAC_P.n274 VDAC_P.n273 0.180667
R18777 VDAC_P.n275 VDAC_P.n274 0.180667
R18778 VDAC_P.n276 VDAC_P.n275 0.180667
R18779 VDAC_P.n277 VDAC_P.n276 0.180667
R18780 VDAC_P.n278 VDAC_P.n277 0.180667
R18781 VDAC_P.n279 VDAC_P.n278 0.180667
R18782 VDAC_P.n280 VDAC_P.n279 0.180667
R18783 VDAC_P.n281 VDAC_P.n280 0.180667
R18784 VDAC_P.n282 VDAC_P.n281 0.180667
R18785 VDAC_P.n283 VDAC_P.n282 0.180667
R18786 VDAC_P.n284 VDAC_P.n283 0.180667
R18787 VDAC_P.n285 VDAC_P.n284 0.180667
R18788 VDAC_P.n286 VDAC_P.n285 0.180667
R18789 VDAC_P.n287 VDAC_P.n286 0.180667
R18790 VDAC_P.n288 VDAC_P.n287 0.180667
R18791 VDAC_P.n289 VDAC_P.n288 0.180667
R18792 VDAC_P.n290 VDAC_P.n289 0.180667
R18793 VDAC_P.n291 VDAC_P.n290 0.180667
R18794 VDAC_P.n292 VDAC_P.n291 0.180667
R18795 VDAC_P.n293 VDAC_P.n292 0.180667
R18796 VDAC_P.n294 VDAC_P.n293 0.180667
R18797 VDAC_P.n295 VDAC_P.n294 0.180667
R18798 VDAC_P.n296 VDAC_P.n295 0.180667
R18799 VDAC_P.n297 VDAC_P.n296 0.180667
R18800 VDAC_P.n298 VDAC_P.n297 0.180667
R18801 VDAC_P.n299 VDAC_P.n298 0.180667
R18802 VDAC_P.n300 VDAC_P.n299 0.180667
R18803 VDAC_P.n301 VDAC_P.n300 0.180667
R18804 VDAC_P.n302 VDAC_P.n301 0.180667
R18805 VDAC_P.n303 VDAC_P.n302 0.180667
R18806 VDAC_P.n304 VDAC_P.n303 0.180667
R18807 VDAC_P.n305 VDAC_P.n304 0.180667
R18808 VDAC_P.n306 VDAC_P.n113 0.180667
R18809 VDAC_P.n307 VDAC_P.n306 0.180667
R18810 VDAC_P.n308 VDAC_P.n307 0.180667
R18811 VDAC_P.n309 VDAC_P.n308 0.180667
R18812 VDAC_P.n310 VDAC_P.n309 0.180667
R18813 VDAC_P.n311 VDAC_P.n310 0.180667
R18814 VDAC_P.n312 VDAC_P.n311 0.180667
R18815 VDAC_P.n313 VDAC_P.n312 0.180667
R18816 VDAC_P.n314 VDAC_P.n313 0.180667
R18817 VDAC_P.n315 VDAC_P.n314 0.180667
R18818 VDAC_P.n316 VDAC_P.n315 0.180667
R18819 VDAC_P.n317 VDAC_P.n316 0.180667
R18820 VDAC_P.n318 VDAC_P.n317 0.180667
R18821 VDAC_P.n319 VDAC_P.n318 0.180667
R18822 VDAC_P.n320 VDAC_P.n319 0.180667
R18823 VDAC_P.n321 VDAC_P.n320 0.180667
R18824 VDAC_P.n322 VDAC_P.n321 0.180667
R18825 VDAC_P.n323 VDAC_P.n322 0.180667
R18826 VDAC_P.n324 VDAC_P.n323 0.180667
R18827 VDAC_P.n325 VDAC_P.n324 0.180667
R18828 VDAC_P.n326 VDAC_P.n325 0.180667
R18829 VDAC_P.n327 VDAC_P.n326 0.180667
R18830 VDAC_P.n328 VDAC_P.n327 0.180667
R18831 VDAC_P.n329 VDAC_P.n328 0.180667
R18832 VDAC_P.n330 VDAC_P.n329 0.180667
R18833 VDAC_P.n331 VDAC_P.n330 0.180667
R18834 VDAC_P.n332 VDAC_P.n331 0.180667
R18835 VDAC_P.n333 VDAC_P.n332 0.180667
R18836 VDAC_P.n334 VDAC_P.n333 0.180667
R18837 VDAC_P.n335 VDAC_P.n334 0.180667
R18838 VDAC_P.n336 VDAC_P.n335 0.180667
R18839 VDAC_P.n337 VDAC_P.n336 0.180667
R18840 VDAC_P.n338 VDAC_P.n337 0.180667
R18841 VDAC_P.n339 VDAC_P.n338 0.180667
R18842 VDAC_P.n340 VDAC_P.n339 0.180667
R18843 VDAC_P.n341 VDAC_P.n340 0.180667
R18844 VDAC_P.n342 VDAC_P.n341 0.180667
R18845 VDAC_P.n343 VDAC_P.n342 0.180667
R18846 VDAC_P.n344 VDAC_P.n343 0.180667
R18847 VDAC_P.n345 VDAC_P.n344 0.180667
R18848 VDAC_P.n346 VDAC_P.n345 0.180667
R18849 VDAC_P.n347 VDAC_P.n346 0.180667
R18850 VDAC_P.n348 VDAC_P.n347 0.180667
R18851 VDAC_P.n349 VDAC_P.n348 0.180667
R18852 VDAC_P.n350 VDAC_P.n349 0.180667
R18853 VDAC_P.n351 VDAC_P.n350 0.180667
R18854 VDAC_P.n352 VDAC_P.n351 0.180667
R18855 VDAC_P.n353 VDAC_P.n352 0.180667
R18856 VDAC_P.n354 VDAC_P.n353 0.180667
R18857 VDAC_P.n355 VDAC_P.n354 0.180667
R18858 VDAC_P.n356 VDAC_P.n355 0.180667
R18859 VDAC_P.n357 VDAC_P.n356 0.180667
R18860 VDAC_P.n358 VDAC_P.n357 0.180667
R18861 VDAC_P.n359 VDAC_P.n358 0.180667
R18862 VDAC_P.n360 VDAC_P.n359 0.180667
R18863 VDAC_P.n361 VDAC_P.n360 0.180667
R18864 VDAC_P.n362 VDAC_P.n361 0.180667
R18865 VDAC_P.n363 VDAC_P.n362 0.180667
R18866 VDAC_P.n364 VDAC_P.n363 0.180667
R18867 VDAC_P.n365 VDAC_P.n364 0.180667
R18868 VDAC_P.n366 VDAC_P.n365 0.180667
R18869 VDAC_P.n367 VDAC_P.n366 0.180667
R18870 VDAC_P.n368 VDAC_P.n367 0.180667
R18871 VDAC_P.n369 VDAC_P.n112 0.180667
R18872 VDAC_P.n370 VDAC_P.n369 0.180667
R18873 VDAC_P.n371 VDAC_P.n370 0.180667
R18874 VDAC_P.n372 VDAC_P.n371 0.180667
R18875 VDAC_P.n373 VDAC_P.n372 0.180667
R18876 VDAC_P.n374 VDAC_P.n373 0.180667
R18877 VDAC_P.n375 VDAC_P.n374 0.180667
R18878 VDAC_P.n376 VDAC_P.n375 0.180667
R18879 VDAC_P.n377 VDAC_P.n376 0.180667
R18880 VDAC_P.n378 VDAC_P.n377 0.180667
R18881 VDAC_P.n379 VDAC_P.n378 0.180667
R18882 VDAC_P.n380 VDAC_P.n379 0.180667
R18883 VDAC_P.n381 VDAC_P.n380 0.180667
R18884 VDAC_P.n382 VDAC_P.n381 0.180667
R18885 VDAC_P.n383 VDAC_P.n382 0.180667
R18886 VDAC_P.n384 VDAC_P.n383 0.180667
R18887 VDAC_P.n385 VDAC_P.n384 0.180667
R18888 VDAC_P.n386 VDAC_P.n385 0.180667
R18889 VDAC_P.n387 VDAC_P.n386 0.180667
R18890 VDAC_P.n388 VDAC_P.n387 0.180667
R18891 VDAC_P.n389 VDAC_P.n388 0.180667
R18892 VDAC_P.n390 VDAC_P.n389 0.180667
R18893 VDAC_P.n391 VDAC_P.n390 0.180667
R18894 VDAC_P.n392 VDAC_P.n391 0.180667
R18895 VDAC_P.n393 VDAC_P.n392 0.180667
R18896 VDAC_P.n394 VDAC_P.n393 0.180667
R18897 VDAC_P.n395 VDAC_P.n394 0.180667
R18898 VDAC_P.n396 VDAC_P.n395 0.180667
R18899 VDAC_P.n397 VDAC_P.n396 0.180667
R18900 VDAC_P.n398 VDAC_P.n397 0.180667
R18901 VDAC_P.n399 VDAC_P.n398 0.180667
R18902 VDAC_P.n400 VDAC_P.n399 0.180667
R18903 VDAC_P.n401 VDAC_P.n400 0.180667
R18904 VDAC_P.n402 VDAC_P.n401 0.180667
R18905 VDAC_P.n403 VDAC_P.n402 0.180667
R18906 VDAC_P.n404 VDAC_P.n403 0.180667
R18907 VDAC_P.n405 VDAC_P.n404 0.180667
R18908 VDAC_P.n406 VDAC_P.n405 0.180667
R18909 VDAC_P.n407 VDAC_P.n406 0.180667
R18910 VDAC_P.n408 VDAC_P.n407 0.180667
R18911 VDAC_P.n409 VDAC_P.n408 0.180667
R18912 VDAC_P.n410 VDAC_P.n409 0.180667
R18913 VDAC_P.n411 VDAC_P.n410 0.180667
R18914 VDAC_P.n412 VDAC_P.n411 0.180667
R18915 VDAC_P.n413 VDAC_P.n412 0.180667
R18916 VDAC_P.n414 VDAC_P.n413 0.180667
R18917 VDAC_P.n415 VDAC_P.n414 0.180667
R18918 VDAC_P.n416 VDAC_P.n415 0.180667
R18919 VDAC_P.n417 VDAC_P.n416 0.180667
R18920 VDAC_P.n418 VDAC_P.n417 0.180667
R18921 VDAC_P.n419 VDAC_P.n418 0.180667
R18922 VDAC_P.n420 VDAC_P.n419 0.180667
R18923 VDAC_P.n421 VDAC_P.n420 0.180667
R18924 VDAC_P.n422 VDAC_P.n421 0.180667
R18925 VDAC_P.n423 VDAC_P.n422 0.180667
R18926 VDAC_P.n424 VDAC_P.n423 0.180667
R18927 VDAC_P.n425 VDAC_P.n424 0.180667
R18928 VDAC_P.n426 VDAC_P.n425 0.180667
R18929 VDAC_P.n427 VDAC_P.n426 0.180667
R18930 VDAC_P.n428 VDAC_P.n427 0.180667
R18931 VDAC_P.n429 VDAC_P.n428 0.180667
R18932 VDAC_P.n430 VDAC_P.n429 0.180667
R18933 VDAC_P.n431 VDAC_P.n430 0.180667
R18934 VDAC_P.n432 VDAC_P.n111 0.180667
R18935 VDAC_P.n433 VDAC_P.n432 0.180667
R18936 VDAC_P.n434 VDAC_P.n433 0.180667
R18937 VDAC_P.n435 VDAC_P.n434 0.180667
R18938 VDAC_P.n436 VDAC_P.n435 0.180667
R18939 VDAC_P.n437 VDAC_P.n436 0.180667
R18940 VDAC_P.n438 VDAC_P.n437 0.180667
R18941 VDAC_P.n439 VDAC_P.n438 0.180667
R18942 VDAC_P.n440 VDAC_P.n439 0.180667
R18943 VDAC_P.n441 VDAC_P.n440 0.180667
R18944 VDAC_P.n442 VDAC_P.n441 0.180667
R18945 VDAC_P.n443 VDAC_P.n442 0.180667
R18946 VDAC_P.n444 VDAC_P.n443 0.180667
R18947 VDAC_P.n445 VDAC_P.n444 0.180667
R18948 VDAC_P.n446 VDAC_P.n445 0.180667
R18949 VDAC_P.n447 VDAC_P.n446 0.180667
R18950 VDAC_P.n448 VDAC_P.n447 0.180667
R18951 VDAC_P.n449 VDAC_P.n448 0.180667
R18952 VDAC_P.n450 VDAC_P.n449 0.180667
R18953 VDAC_P.n451 VDAC_P.n450 0.180667
R18954 VDAC_P.n452 VDAC_P.n451 0.180667
R18955 VDAC_P.n453 VDAC_P.n452 0.180667
R18956 VDAC_P.n454 VDAC_P.n453 0.180667
R18957 VDAC_P.n455 VDAC_P.n454 0.180667
R18958 VDAC_P.n456 VDAC_P.n455 0.180667
R18959 VDAC_P.n457 VDAC_P.n456 0.180667
R18960 VDAC_P.n458 VDAC_P.n457 0.180667
R18961 VDAC_P.n459 VDAC_P.n458 0.180667
R18962 VDAC_P.n460 VDAC_P.n459 0.180667
R18963 VDAC_P.n461 VDAC_P.n460 0.180667
R18964 VDAC_P.n462 VDAC_P.n461 0.180667
R18965 VDAC_P.n463 VDAC_P.n462 0.180667
R18966 VDAC_P.n464 VDAC_P.n463 0.180667
R18967 VDAC_P.n465 VDAC_P.n464 0.180667
R18968 VDAC_P.n466 VDAC_P.n465 0.180667
R18969 VDAC_P.n467 VDAC_P.n466 0.180667
R18970 VDAC_P.n468 VDAC_P.n467 0.180667
R18971 VDAC_P.n469 VDAC_P.n468 0.180667
R18972 VDAC_P.n470 VDAC_P.n469 0.180667
R18973 VDAC_P.n471 VDAC_P.n470 0.180667
R18974 VDAC_P.n472 VDAC_P.n471 0.180667
R18975 VDAC_P.n473 VDAC_P.n472 0.180667
R18976 VDAC_P.n474 VDAC_P.n473 0.180667
R18977 VDAC_P.n475 VDAC_P.n474 0.180667
R18978 VDAC_P.n476 VDAC_P.n475 0.180667
R18979 VDAC_P.n477 VDAC_P.n476 0.180667
R18980 VDAC_P.n478 VDAC_P.n477 0.180667
R18981 VDAC_P.n479 VDAC_P.n478 0.180667
R18982 VDAC_P.n480 VDAC_P.n479 0.180667
R18983 VDAC_P.n481 VDAC_P.n480 0.180667
R18984 VDAC_P.n482 VDAC_P.n481 0.180667
R18985 VDAC_P.n483 VDAC_P.n482 0.180667
R18986 VDAC_P.n484 VDAC_P.n483 0.180667
R18987 VDAC_P.n485 VDAC_P.n484 0.180667
R18988 VDAC_P.n486 VDAC_P.n485 0.180667
R18989 VDAC_P.n487 VDAC_P.n486 0.180667
R18990 VDAC_P.n488 VDAC_P.n487 0.180667
R18991 VDAC_P.n489 VDAC_P.n488 0.180667
R18992 VDAC_P.n490 VDAC_P.n489 0.180667
R18993 VDAC_P.n491 VDAC_P.n490 0.180667
R18994 VDAC_P.n492 VDAC_P.n491 0.180667
R18995 VDAC_P.n493 VDAC_P.n492 0.180667
R18996 VDAC_P.n494 VDAC_P.n493 0.180667
R18997 VDAC_P.n495 VDAC_P.n110 0.180667
R18998 VDAC_P.n496 VDAC_P.n495 0.180667
R18999 VDAC_P.n497 VDAC_P.n496 0.180667
R19000 VDAC_P.n498 VDAC_P.n497 0.180667
R19001 VDAC_P.n499 VDAC_P.n498 0.180667
R19002 VDAC_P.n500 VDAC_P.n499 0.180667
R19003 VDAC_P.n501 VDAC_P.n500 0.180667
R19004 VDAC_P.n502 VDAC_P.n501 0.180667
R19005 VDAC_P.n503 VDAC_P.n502 0.180667
R19006 VDAC_P.n504 VDAC_P.n503 0.180667
R19007 VDAC_P.n505 VDAC_P.n504 0.180667
R19008 VDAC_P.n506 VDAC_P.n505 0.180667
R19009 VDAC_P.n507 VDAC_P.n506 0.180667
R19010 VDAC_P.n508 VDAC_P.n507 0.180667
R19011 VDAC_P.n509 VDAC_P.n508 0.180667
R19012 VDAC_P.n510 VDAC_P.n509 0.180667
R19013 VDAC_P.n511 VDAC_P.n510 0.180667
R19014 VDAC_P.n512 VDAC_P.n511 0.180667
R19015 VDAC_P.n513 VDAC_P.n512 0.180667
R19016 VDAC_P.n514 VDAC_P.n513 0.180667
R19017 VDAC_P.n515 VDAC_P.n514 0.180667
R19018 VDAC_P.n516 VDAC_P.n515 0.180667
R19019 VDAC_P.n517 VDAC_P.n516 0.180667
R19020 VDAC_P.n518 VDAC_P.n517 0.180667
R19021 VDAC_P.n519 VDAC_P.n518 0.180667
R19022 VDAC_P.n520 VDAC_P.n519 0.180667
R19023 VDAC_P.n521 VDAC_P.n520 0.180667
R19024 VDAC_P.n522 VDAC_P.n521 0.180667
R19025 VDAC_P.n523 VDAC_P.n522 0.180667
R19026 VDAC_P.n524 VDAC_P.n523 0.180667
R19027 VDAC_P.n525 VDAC_P.n524 0.180667
R19028 VDAC_P.n526 VDAC_P.n525 0.180667
R19029 VDAC_P.n527 VDAC_P.n526 0.180667
R19030 VDAC_P.n528 VDAC_P.n527 0.180667
R19031 VDAC_P.n529 VDAC_P.n528 0.180667
R19032 VDAC_P.n530 VDAC_P.n529 0.180667
R19033 VDAC_P.n531 VDAC_P.n530 0.180667
R19034 VDAC_P.n532 VDAC_P.n531 0.180667
R19035 VDAC_P.n533 VDAC_P.n532 0.180667
R19036 VDAC_P.n534 VDAC_P.n533 0.180667
R19037 VDAC_P.n535 VDAC_P.n534 0.180667
R19038 VDAC_P.n536 VDAC_P.n535 0.180667
R19039 VDAC_P.n537 VDAC_P.n536 0.180667
R19040 VDAC_P.n538 VDAC_P.n537 0.180667
R19041 VDAC_P.n539 VDAC_P.n538 0.180667
R19042 VDAC_P.n540 VDAC_P.n539 0.180667
R19043 VDAC_P.n541 VDAC_P.n540 0.180667
R19044 VDAC_P.n542 VDAC_P.n541 0.180667
R19045 VDAC_P.n543 VDAC_P.n542 0.180667
R19046 VDAC_P.n544 VDAC_P.n543 0.180667
R19047 VDAC_P.n545 VDAC_P.n544 0.180667
R19048 VDAC_P.n546 VDAC_P.n545 0.180667
R19049 VDAC_P.n547 VDAC_P.n546 0.180667
R19050 VDAC_P.n548 VDAC_P.n547 0.180667
R19051 VDAC_P.n549 VDAC_P.n548 0.180667
R19052 VDAC_P.n550 VDAC_P.n549 0.180667
R19053 VDAC_P.n551 VDAC_P.n550 0.180667
R19054 VDAC_P.n552 VDAC_P.n551 0.180667
R19055 VDAC_P.n553 VDAC_P.n552 0.180667
R19056 VDAC_P.n554 VDAC_P.n553 0.180667
R19057 VDAC_P.n555 VDAC_P.n554 0.180667
R19058 VDAC_P.n556 VDAC_P.n555 0.180667
R19059 VDAC_P.n557 VDAC_P.n556 0.180667
R19060 VDAC_P.n558 VDAC_P.n109 0.180667
R19061 VDAC_P.n559 VDAC_P.n558 0.180667
R19062 VDAC_P.n560 VDAC_P.n559 0.180667
R19063 VDAC_P.n561 VDAC_P.n560 0.180667
R19064 VDAC_P.n562 VDAC_P.n561 0.180667
R19065 VDAC_P.n563 VDAC_P.n562 0.180667
R19066 VDAC_P.n564 VDAC_P.n563 0.180667
R19067 VDAC_P.n565 VDAC_P.n564 0.180667
R19068 VDAC_P.n566 VDAC_P.n565 0.180667
R19069 VDAC_P.n567 VDAC_P.n566 0.180667
R19070 VDAC_P.n568 VDAC_P.n567 0.180667
R19071 VDAC_P.n569 VDAC_P.n568 0.180667
R19072 VDAC_P.n570 VDAC_P.n569 0.180667
R19073 VDAC_P.n571 VDAC_P.n570 0.180667
R19074 VDAC_P.n572 VDAC_P.n571 0.180667
R19075 VDAC_P.n573 VDAC_P.n572 0.180667
R19076 VDAC_P.n574 VDAC_P.n573 0.180667
R19077 VDAC_P.n575 VDAC_P.n574 0.180667
R19078 VDAC_P.n576 VDAC_P.n575 0.180667
R19079 VDAC_P.n577 VDAC_P.n576 0.180667
R19080 VDAC_P.n578 VDAC_P.n577 0.180667
R19081 VDAC_P.n579 VDAC_P.n578 0.180667
R19082 VDAC_P.n580 VDAC_P.n579 0.180667
R19083 VDAC_P.n581 VDAC_P.n580 0.180667
R19084 VDAC_P.n582 VDAC_P.n581 0.180667
R19085 VDAC_P.n583 VDAC_P.n582 0.180667
R19086 VDAC_P.n584 VDAC_P.n583 0.180667
R19087 VDAC_P.n585 VDAC_P.n584 0.180667
R19088 VDAC_P.n586 VDAC_P.n585 0.180667
R19089 VDAC_P.n587 VDAC_P.n586 0.180667
R19090 VDAC_P.n588 VDAC_P.n587 0.180667
R19091 VDAC_P.n589 VDAC_P.n588 0.180667
R19092 VDAC_P.n590 VDAC_P.n589 0.180667
R19093 VDAC_P.n591 VDAC_P.n590 0.180667
R19094 VDAC_P.n592 VDAC_P.n591 0.180667
R19095 VDAC_P.n593 VDAC_P.n592 0.180667
R19096 VDAC_P.n594 VDAC_P.n593 0.180667
R19097 VDAC_P.n595 VDAC_P.n594 0.180667
R19098 VDAC_P.n596 VDAC_P.n595 0.180667
R19099 VDAC_P.n597 VDAC_P.n596 0.180667
R19100 VDAC_P.n598 VDAC_P.n597 0.180667
R19101 VDAC_P.n599 VDAC_P.n598 0.180667
R19102 VDAC_P.n600 VDAC_P.n599 0.180667
R19103 VDAC_P.n601 VDAC_P.n600 0.180667
R19104 VDAC_P.n602 VDAC_P.n601 0.180667
R19105 VDAC_P.n603 VDAC_P.n602 0.180667
R19106 VDAC_P.n604 VDAC_P.n603 0.180667
R19107 VDAC_P.n605 VDAC_P.n604 0.180667
R19108 VDAC_P.n606 VDAC_P.n605 0.180667
R19109 VDAC_P.n607 VDAC_P.n606 0.180667
R19110 VDAC_P.n608 VDAC_P.n607 0.180667
R19111 VDAC_P.n609 VDAC_P.n608 0.180667
R19112 VDAC_P.n610 VDAC_P.n609 0.180667
R19113 VDAC_P.n611 VDAC_P.n610 0.180667
R19114 VDAC_P.n612 VDAC_P.n611 0.180667
R19115 VDAC_P.n613 VDAC_P.n612 0.180667
R19116 VDAC_P.n614 VDAC_P.n613 0.180667
R19117 VDAC_P.n615 VDAC_P.n614 0.180667
R19118 VDAC_P.n616 VDAC_P.n615 0.180667
R19119 VDAC_P.n617 VDAC_P.n616 0.180667
R19120 VDAC_P.n618 VDAC_P.n617 0.180667
R19121 VDAC_P.n619 VDAC_P.n618 0.180667
R19122 VDAC_P.n620 VDAC_P.n619 0.180667
R19123 VDAC_P.n621 VDAC_P.n108 0.180667
R19124 VDAC_P.n622 VDAC_P.n621 0.180667
R19125 VDAC_P.n623 VDAC_P.n622 0.180667
R19126 VDAC_P.n624 VDAC_P.n623 0.180667
R19127 VDAC_P.n625 VDAC_P.n624 0.180667
R19128 VDAC_P.n626 VDAC_P.n625 0.180667
R19129 VDAC_P.n627 VDAC_P.n626 0.180667
R19130 VDAC_P.n628 VDAC_P.n627 0.180667
R19131 VDAC_P.n629 VDAC_P.n628 0.180667
R19132 VDAC_P.n630 VDAC_P.n629 0.180667
R19133 VDAC_P.n631 VDAC_P.n630 0.180667
R19134 VDAC_P.n632 VDAC_P.n631 0.180667
R19135 VDAC_P.n633 VDAC_P.n632 0.180667
R19136 VDAC_P.n634 VDAC_P.n633 0.180667
R19137 VDAC_P.n635 VDAC_P.n634 0.180667
R19138 VDAC_P.n636 VDAC_P.n635 0.180667
R19139 VDAC_P.n637 VDAC_P.n636 0.180667
R19140 VDAC_P.n638 VDAC_P.n637 0.180667
R19141 VDAC_P.n639 VDAC_P.n638 0.180667
R19142 VDAC_P.n640 VDAC_P.n639 0.180667
R19143 VDAC_P.n641 VDAC_P.n640 0.180667
R19144 VDAC_P.n642 VDAC_P.n641 0.180667
R19145 VDAC_P.n643 VDAC_P.n642 0.180667
R19146 VDAC_P.n644 VDAC_P.n643 0.180667
R19147 VDAC_P.n645 VDAC_P.n644 0.180667
R19148 VDAC_P.n646 VDAC_P.n645 0.180667
R19149 VDAC_P.n647 VDAC_P.n646 0.180667
R19150 VDAC_P.n648 VDAC_P.n647 0.180667
R19151 VDAC_P.n649 VDAC_P.n648 0.180667
R19152 VDAC_P.n650 VDAC_P.n649 0.180667
R19153 VDAC_P.n651 VDAC_P.n650 0.180667
R19154 VDAC_P.n652 VDAC_P.n651 0.180667
R19155 VDAC_P.n653 VDAC_P.n652 0.180667
R19156 VDAC_P.n654 VDAC_P.n653 0.180667
R19157 VDAC_P.n655 VDAC_P.n654 0.180667
R19158 VDAC_P.n656 VDAC_P.n655 0.180667
R19159 VDAC_P.n657 VDAC_P.n656 0.180667
R19160 VDAC_P.n658 VDAC_P.n657 0.180667
R19161 VDAC_P.n659 VDAC_P.n658 0.180667
R19162 VDAC_P.n660 VDAC_P.n659 0.180667
R19163 VDAC_P.n661 VDAC_P.n660 0.180667
R19164 VDAC_P.n662 VDAC_P.n661 0.180667
R19165 VDAC_P.n663 VDAC_P.n662 0.180667
R19166 VDAC_P.n664 VDAC_P.n663 0.180667
R19167 VDAC_P.n665 VDAC_P.n664 0.180667
R19168 VDAC_P.n666 VDAC_P.n665 0.180667
R19169 VDAC_P.n667 VDAC_P.n666 0.180667
R19170 VDAC_P.n668 VDAC_P.n667 0.180667
R19171 VDAC_P.n669 VDAC_P.n668 0.180667
R19172 VDAC_P.n670 VDAC_P.n669 0.180667
R19173 VDAC_P.n671 VDAC_P.n670 0.180667
R19174 VDAC_P.n672 VDAC_P.n671 0.180667
R19175 VDAC_P.n673 VDAC_P.n672 0.180667
R19176 VDAC_P.n674 VDAC_P.n673 0.180667
R19177 VDAC_P.n675 VDAC_P.n674 0.180667
R19178 VDAC_P.n676 VDAC_P.n675 0.180667
R19179 VDAC_P.n677 VDAC_P.n676 0.180667
R19180 VDAC_P.n678 VDAC_P.n677 0.180667
R19181 VDAC_P.n679 VDAC_P.n678 0.180667
R19182 VDAC_P.n680 VDAC_P.n679 0.180667
R19183 VDAC_P.n681 VDAC_P.n680 0.180667
R19184 VDAC_P.n682 VDAC_P.n681 0.180667
R19185 VDAC_P.n683 VDAC_P.n682 0.180667
R19186 VDAC_P.n684 VDAC_P.n107 0.180667
R19187 VDAC_P.n685 VDAC_P.n684 0.180667
R19188 VDAC_P.n686 VDAC_P.n685 0.180667
R19189 VDAC_P.n687 VDAC_P.n686 0.180667
R19190 VDAC_P.n688 VDAC_P.n687 0.180667
R19191 VDAC_P.n689 VDAC_P.n688 0.180667
R19192 VDAC_P.n690 VDAC_P.n689 0.180667
R19193 VDAC_P.n691 VDAC_P.n690 0.180667
R19194 VDAC_P.n692 VDAC_P.n691 0.180667
R19195 VDAC_P.n693 VDAC_P.n692 0.180667
R19196 VDAC_P.n694 VDAC_P.n693 0.180667
R19197 VDAC_P.n695 VDAC_P.n694 0.180667
R19198 VDAC_P.n696 VDAC_P.n695 0.180667
R19199 VDAC_P.n697 VDAC_P.n696 0.180667
R19200 VDAC_P.n698 VDAC_P.n697 0.180667
R19201 VDAC_P.n699 VDAC_P.n698 0.180667
R19202 VDAC_P.n700 VDAC_P.n699 0.180667
R19203 VDAC_P.n701 VDAC_P.n700 0.180667
R19204 VDAC_P.n702 VDAC_P.n701 0.180667
R19205 VDAC_P.n703 VDAC_P.n702 0.180667
R19206 VDAC_P.n704 VDAC_P.n703 0.180667
R19207 VDAC_P.n705 VDAC_P.n704 0.180667
R19208 VDAC_P.n706 VDAC_P.n705 0.180667
R19209 VDAC_P.n707 VDAC_P.n706 0.180667
R19210 VDAC_P.n708 VDAC_P.n707 0.180667
R19211 VDAC_P.n709 VDAC_P.n708 0.180667
R19212 VDAC_P.n710 VDAC_P.n709 0.180667
R19213 VDAC_P.n711 VDAC_P.n710 0.180667
R19214 VDAC_P.n712 VDAC_P.n711 0.180667
R19215 VDAC_P.n713 VDAC_P.n712 0.180667
R19216 VDAC_P.n714 VDAC_P.n713 0.180667
R19217 VDAC_P.n715 VDAC_P.n714 0.180667
R19218 VDAC_P.n716 VDAC_P.n715 0.180667
R19219 VDAC_P.n717 VDAC_P.n716 0.180667
R19220 VDAC_P.n718 VDAC_P.n717 0.180667
R19221 VDAC_P.n719 VDAC_P.n718 0.180667
R19222 VDAC_P.n720 VDAC_P.n719 0.180667
R19223 VDAC_P.n721 VDAC_P.n720 0.180667
R19224 VDAC_P.n722 VDAC_P.n721 0.180667
R19225 VDAC_P.n723 VDAC_P.n722 0.180667
R19226 VDAC_P.n724 VDAC_P.n723 0.180667
R19227 VDAC_P.n725 VDAC_P.n724 0.180667
R19228 VDAC_P.n726 VDAC_P.n725 0.180667
R19229 VDAC_P.n727 VDAC_P.n726 0.180667
R19230 VDAC_P.n728 VDAC_P.n727 0.180667
R19231 VDAC_P.n729 VDAC_P.n728 0.180667
R19232 VDAC_P.n730 VDAC_P.n729 0.180667
R19233 VDAC_P.n731 VDAC_P.n730 0.180667
R19234 VDAC_P.n732 VDAC_P.n731 0.180667
R19235 VDAC_P.n733 VDAC_P.n732 0.180667
R19236 VDAC_P.n734 VDAC_P.n733 0.180667
R19237 VDAC_P.n735 VDAC_P.n734 0.180667
R19238 VDAC_P.n736 VDAC_P.n735 0.180667
R19239 VDAC_P.n737 VDAC_P.n736 0.180667
R19240 VDAC_P.n738 VDAC_P.n737 0.180667
R19241 VDAC_P.n739 VDAC_P.n738 0.180667
R19242 VDAC_P.n740 VDAC_P.n739 0.180667
R19243 VDAC_P.n741 VDAC_P.n740 0.180667
R19244 VDAC_P.n742 VDAC_P.n741 0.180667
R19245 VDAC_P.n743 VDAC_P.n742 0.180667
R19246 VDAC_P.n744 VDAC_P.n743 0.180667
R19247 VDAC_P.n745 VDAC_P.n744 0.180667
R19248 VDAC_P.n746 VDAC_P.n745 0.180667
R19249 VDAC_P.n747 VDAC_P.n106 0.180667
R19250 VDAC_P.n748 VDAC_P.n747 0.180667
R19251 VDAC_P.n749 VDAC_P.n748 0.180667
R19252 VDAC_P.n750 VDAC_P.n749 0.180667
R19253 VDAC_P.n751 VDAC_P.n750 0.180667
R19254 VDAC_P.n752 VDAC_P.n751 0.180667
R19255 VDAC_P.n753 VDAC_P.n752 0.180667
R19256 VDAC_P.n754 VDAC_P.n753 0.180667
R19257 VDAC_P.n755 VDAC_P.n754 0.180667
R19258 VDAC_P.n756 VDAC_P.n755 0.180667
R19259 VDAC_P.n757 VDAC_P.n756 0.180667
R19260 VDAC_P.n758 VDAC_P.n757 0.180667
R19261 VDAC_P.n759 VDAC_P.n758 0.180667
R19262 VDAC_P.n760 VDAC_P.n759 0.180667
R19263 VDAC_P.n761 VDAC_P.n760 0.180667
R19264 VDAC_P.n762 VDAC_P.n761 0.180667
R19265 VDAC_P.n763 VDAC_P.n762 0.180667
R19266 VDAC_P.n764 VDAC_P.n763 0.180667
R19267 VDAC_P.n765 VDAC_P.n764 0.180667
R19268 VDAC_P.n766 VDAC_P.n765 0.180667
R19269 VDAC_P.n767 VDAC_P.n766 0.180667
R19270 VDAC_P.n768 VDAC_P.n767 0.180667
R19271 VDAC_P.n769 VDAC_P.n768 0.180667
R19272 VDAC_P.n770 VDAC_P.n769 0.180667
R19273 VDAC_P.n771 VDAC_P.n770 0.180667
R19274 VDAC_P.n772 VDAC_P.n771 0.180667
R19275 VDAC_P.n773 VDAC_P.n772 0.180667
R19276 VDAC_P.n774 VDAC_P.n773 0.180667
R19277 VDAC_P.n775 VDAC_P.n774 0.180667
R19278 VDAC_P.n776 VDAC_P.n775 0.180667
R19279 VDAC_P.n777 VDAC_P.n776 0.180667
R19280 VDAC_P.n778 VDAC_P.n777 0.180667
R19281 VDAC_P.n779 VDAC_P.n778 0.180667
R19282 VDAC_P.n780 VDAC_P.n779 0.180667
R19283 VDAC_P.n781 VDAC_P.n780 0.180667
R19284 VDAC_P.n782 VDAC_P.n781 0.180667
R19285 VDAC_P.n783 VDAC_P.n782 0.180667
R19286 VDAC_P.n784 VDAC_P.n783 0.180667
R19287 VDAC_P.n785 VDAC_P.n784 0.180667
R19288 VDAC_P.n786 VDAC_P.n785 0.180667
R19289 VDAC_P.n787 VDAC_P.n786 0.180667
R19290 VDAC_P.n788 VDAC_P.n787 0.180667
R19291 VDAC_P.n789 VDAC_P.n788 0.180667
R19292 VDAC_P.n790 VDAC_P.n789 0.180667
R19293 VDAC_P.n791 VDAC_P.n790 0.180667
R19294 VDAC_P.n792 VDAC_P.n791 0.180667
R19295 VDAC_P.n793 VDAC_P.n792 0.180667
R19296 VDAC_P.n794 VDAC_P.n793 0.180667
R19297 VDAC_P.n795 VDAC_P.n794 0.180667
R19298 VDAC_P.n796 VDAC_P.n795 0.180667
R19299 VDAC_P.n797 VDAC_P.n796 0.180667
R19300 VDAC_P.n798 VDAC_P.n797 0.180667
R19301 VDAC_P.n799 VDAC_P.n798 0.180667
R19302 VDAC_P.n800 VDAC_P.n799 0.180667
R19303 VDAC_P.n801 VDAC_P.n800 0.180667
R19304 VDAC_P.n802 VDAC_P.n801 0.180667
R19305 VDAC_P.n803 VDAC_P.n802 0.180667
R19306 VDAC_P.n804 VDAC_P.n803 0.180667
R19307 VDAC_P.n805 VDAC_P.n804 0.180667
R19308 VDAC_P.n806 VDAC_P.n805 0.180667
R19309 VDAC_P.n807 VDAC_P.n806 0.180667
R19310 VDAC_P.n808 VDAC_P.n807 0.180667
R19311 VDAC_P.n809 VDAC_P.n808 0.180667
R19312 VDAC_P.n810 VDAC_P.n105 0.180667
R19313 VDAC_P.n811 VDAC_P.n810 0.180667
R19314 VDAC_P.n812 VDAC_P.n811 0.180667
R19315 VDAC_P.n813 VDAC_P.n812 0.180667
R19316 VDAC_P.n814 VDAC_P.n813 0.180667
R19317 VDAC_P.n815 VDAC_P.n814 0.180667
R19318 VDAC_P.n816 VDAC_P.n815 0.180667
R19319 VDAC_P.n817 VDAC_P.n816 0.180667
R19320 VDAC_P.n818 VDAC_P.n817 0.180667
R19321 VDAC_P.n819 VDAC_P.n818 0.180667
R19322 VDAC_P.n820 VDAC_P.n819 0.180667
R19323 VDAC_P.n821 VDAC_P.n820 0.180667
R19324 VDAC_P.n822 VDAC_P.n821 0.180667
R19325 VDAC_P.n823 VDAC_P.n822 0.180667
R19326 VDAC_P.n824 VDAC_P.n823 0.180667
R19327 VDAC_P.n825 VDAC_P.n824 0.180667
R19328 VDAC_P.n826 VDAC_P.n825 0.180667
R19329 VDAC_P.n827 VDAC_P.n826 0.180667
R19330 VDAC_P.n828 VDAC_P.n827 0.180667
R19331 VDAC_P.n829 VDAC_P.n828 0.180667
R19332 VDAC_P.n830 VDAC_P.n829 0.180667
R19333 VDAC_P.n831 VDAC_P.n830 0.180667
R19334 VDAC_P.n832 VDAC_P.n831 0.180667
R19335 VDAC_P.n833 VDAC_P.n832 0.180667
R19336 VDAC_P.n834 VDAC_P.n833 0.180667
R19337 VDAC_P.n835 VDAC_P.n834 0.180667
R19338 VDAC_P.n836 VDAC_P.n835 0.180667
R19339 VDAC_P.n837 VDAC_P.n836 0.180667
R19340 VDAC_P.n838 VDAC_P.n837 0.180667
R19341 VDAC_P.n839 VDAC_P.n838 0.180667
R19342 VDAC_P.n840 VDAC_P.n839 0.180667
R19343 VDAC_P.n841 VDAC_P.n840 0.180667
R19344 VDAC_P.n842 VDAC_P.n841 0.180667
R19345 VDAC_P.n843 VDAC_P.n842 0.180667
R19346 VDAC_P.n844 VDAC_P.n843 0.180667
R19347 VDAC_P.n845 VDAC_P.n844 0.180667
R19348 VDAC_P.n846 VDAC_P.n845 0.180667
R19349 VDAC_P.n847 VDAC_P.n846 0.180667
R19350 VDAC_P.n848 VDAC_P.n847 0.180667
R19351 VDAC_P.n849 VDAC_P.n848 0.180667
R19352 VDAC_P.n850 VDAC_P.n849 0.180667
R19353 VDAC_P.n851 VDAC_P.n850 0.180667
R19354 VDAC_P.n852 VDAC_P.n851 0.180667
R19355 VDAC_P.n853 VDAC_P.n852 0.180667
R19356 VDAC_P.n854 VDAC_P.n853 0.180667
R19357 VDAC_P.n855 VDAC_P.n854 0.180667
R19358 VDAC_P.n856 VDAC_P.n855 0.180667
R19359 VDAC_P.n857 VDAC_P.n856 0.180667
R19360 VDAC_P.n858 VDAC_P.n857 0.180667
R19361 VDAC_P.n859 VDAC_P.n858 0.180667
R19362 VDAC_P.n860 VDAC_P.n859 0.180667
R19363 VDAC_P.n861 VDAC_P.n860 0.180667
R19364 VDAC_P.n862 VDAC_P.n861 0.180667
R19365 VDAC_P.n863 VDAC_P.n862 0.180667
R19366 VDAC_P.n864 VDAC_P.n863 0.180667
R19367 VDAC_P.n865 VDAC_P.n864 0.180667
R19368 VDAC_P.n866 VDAC_P.n865 0.180667
R19369 VDAC_P.n867 VDAC_P.n866 0.180667
R19370 VDAC_P.n868 VDAC_P.n867 0.180667
R19371 VDAC_P.n869 VDAC_P.n868 0.180667
R19372 VDAC_P.n870 VDAC_P.n869 0.180667
R19373 VDAC_P.n871 VDAC_P.n870 0.180667
R19374 VDAC_P.n872 VDAC_P.n871 0.180667
R19375 VDAC_P.n873 VDAC_P.n104 0.180667
R19376 VDAC_P.n874 VDAC_P.n873 0.180667
R19377 VDAC_P.n875 VDAC_P.n874 0.180667
R19378 VDAC_P.n876 VDAC_P.n875 0.180667
R19379 VDAC_P.n877 VDAC_P.n876 0.180667
R19380 VDAC_P.n878 VDAC_P.n877 0.180667
R19381 VDAC_P.n879 VDAC_P.n878 0.180667
R19382 VDAC_P.n880 VDAC_P.n879 0.180667
R19383 VDAC_P.n881 VDAC_P.n880 0.180667
R19384 VDAC_P.n882 VDAC_P.n881 0.180667
R19385 VDAC_P.n883 VDAC_P.n882 0.180667
R19386 VDAC_P.n884 VDAC_P.n883 0.180667
R19387 VDAC_P.n885 VDAC_P.n884 0.180667
R19388 VDAC_P.n886 VDAC_P.n885 0.180667
R19389 VDAC_P.n887 VDAC_P.n886 0.180667
R19390 VDAC_P.n888 VDAC_P.n887 0.180667
R19391 VDAC_P.n889 VDAC_P.n888 0.180667
R19392 VDAC_P.n890 VDAC_P.n889 0.180667
R19393 VDAC_P.n891 VDAC_P.n890 0.180667
R19394 VDAC_P.n892 VDAC_P.n891 0.180667
R19395 VDAC_P.n893 VDAC_P.n892 0.180667
R19396 VDAC_P.n894 VDAC_P.n893 0.180667
R19397 VDAC_P.n895 VDAC_P.n894 0.180667
R19398 VDAC_P.n896 VDAC_P.n895 0.180667
R19399 VDAC_P.n897 VDAC_P.n896 0.180667
R19400 VDAC_P.n898 VDAC_P.n897 0.180667
R19401 VDAC_P.n899 VDAC_P.n898 0.180667
R19402 VDAC_P.n900 VDAC_P.n899 0.180667
R19403 VDAC_P.n901 VDAC_P.n900 0.180667
R19404 VDAC_P.n902 VDAC_P.n901 0.180667
R19405 VDAC_P.n903 VDAC_P.n902 0.180667
R19406 VDAC_P.n904 VDAC_P.n903 0.180667
R19407 VDAC_P.n905 VDAC_P.n904 0.180667
R19408 VDAC_P.n906 VDAC_P.n905 0.180667
R19409 VDAC_P.n907 VDAC_P.n906 0.180667
R19410 VDAC_P.n908 VDAC_P.n907 0.180667
R19411 VDAC_P.n909 VDAC_P.n908 0.180667
R19412 VDAC_P.n910 VDAC_P.n909 0.180667
R19413 VDAC_P.n911 VDAC_P.n910 0.180667
R19414 VDAC_P.n912 VDAC_P.n911 0.180667
R19415 VDAC_P.n913 VDAC_P.n912 0.180667
R19416 VDAC_P.n914 VDAC_P.n913 0.180667
R19417 VDAC_P.n915 VDAC_P.n914 0.180667
R19418 VDAC_P.n916 VDAC_P.n915 0.180667
R19419 VDAC_P.n917 VDAC_P.n916 0.180667
R19420 VDAC_P.n918 VDAC_P.n917 0.180667
R19421 VDAC_P.n919 VDAC_P.n918 0.180667
R19422 VDAC_P.n920 VDAC_P.n919 0.180667
R19423 VDAC_P.n921 VDAC_P.n920 0.180667
R19424 VDAC_P.n922 VDAC_P.n921 0.180667
R19425 VDAC_P.n923 VDAC_P.n922 0.180667
R19426 VDAC_P.n924 VDAC_P.n923 0.180667
R19427 VDAC_P.n925 VDAC_P.n924 0.180667
R19428 VDAC_P.n926 VDAC_P.n925 0.180667
R19429 VDAC_P.n927 VDAC_P.n926 0.180667
R19430 VDAC_P.n928 VDAC_P.n927 0.180667
R19431 VDAC_P.n929 VDAC_P.n928 0.180667
R19432 VDAC_P.n930 VDAC_P.n929 0.180667
R19433 VDAC_P.n931 VDAC_P.n930 0.180667
R19434 VDAC_P.n932 VDAC_P.n931 0.180667
R19435 VDAC_P.n933 VDAC_P.n932 0.180667
R19436 VDAC_P.n934 VDAC_P.n933 0.180667
R19437 VDAC_P.n935 VDAC_P.n934 0.180667
R19438 VDAC_P.n936 VDAC_P.n103 0.180667
R19439 VDAC_P.n937 VDAC_P.n936 0.180667
R19440 VDAC_P.n938 VDAC_P.n937 0.180667
R19441 VDAC_P.n939 VDAC_P.n938 0.180667
R19442 VDAC_P.n940 VDAC_P.n939 0.180667
R19443 VDAC_P.n941 VDAC_P.n940 0.180667
R19444 VDAC_P.n942 VDAC_P.n941 0.180667
R19445 VDAC_P.n943 VDAC_P.n942 0.180667
R19446 VDAC_P.n944 VDAC_P.n943 0.180667
R19447 VDAC_P.n945 VDAC_P.n944 0.180667
R19448 VDAC_P.n946 VDAC_P.n945 0.180667
R19449 VDAC_P.n947 VDAC_P.n946 0.180667
R19450 VDAC_P.n948 VDAC_P.n947 0.180667
R19451 VDAC_P.n949 VDAC_P.n948 0.180667
R19452 VDAC_P.n950 VDAC_P.n949 0.180667
R19453 VDAC_P.n951 VDAC_P.n950 0.180667
R19454 VDAC_P.n952 VDAC_P.n951 0.180667
R19455 VDAC_P.n953 VDAC_P.n952 0.180667
R19456 VDAC_P.n954 VDAC_P.n953 0.180667
R19457 VDAC_P.n955 VDAC_P.n954 0.180667
R19458 VDAC_P.n956 VDAC_P.n955 0.180667
R19459 VDAC_P.n957 VDAC_P.n956 0.180667
R19460 VDAC_P.n958 VDAC_P.n957 0.180667
R19461 VDAC_P.n959 VDAC_P.n958 0.180667
R19462 VDAC_P.n960 VDAC_P.n959 0.180667
R19463 VDAC_P.n961 VDAC_P.n960 0.180667
R19464 VDAC_P.n962 VDAC_P.n961 0.180667
R19465 VDAC_P.n963 VDAC_P.n962 0.180667
R19466 VDAC_P.n964 VDAC_P.n963 0.180667
R19467 VDAC_P.n965 VDAC_P.n964 0.180667
R19468 VDAC_P.n966 VDAC_P.n965 0.180667
R19469 VDAC_P.n967 VDAC_P.n966 0.180667
R19470 VDAC_P.n968 VDAC_P.n967 0.180667
R19471 VDAC_P.n969 VDAC_P.n968 0.180667
R19472 VDAC_P.n970 VDAC_P.n969 0.180667
R19473 VDAC_P.n971 VDAC_P.n970 0.180667
R19474 VDAC_P.n972 VDAC_P.n971 0.180667
R19475 VDAC_P.n973 VDAC_P.n972 0.180667
R19476 VDAC_P.n974 VDAC_P.n973 0.180667
R19477 VDAC_P.n975 VDAC_P.n974 0.180667
R19478 VDAC_P.n976 VDAC_P.n975 0.180667
R19479 VDAC_P.n977 VDAC_P.n976 0.180667
R19480 VDAC_P.n978 VDAC_P.n977 0.180667
R19481 VDAC_P.n979 VDAC_P.n978 0.180667
R19482 VDAC_P.n980 VDAC_P.n979 0.180667
R19483 VDAC_P.n981 VDAC_P.n980 0.180667
R19484 VDAC_P.n982 VDAC_P.n981 0.180667
R19485 VDAC_P.n983 VDAC_P.n982 0.180667
R19486 VDAC_P.n984 VDAC_P.n983 0.180667
R19487 VDAC_P.n985 VDAC_P.n984 0.180667
R19488 VDAC_P.n986 VDAC_P.n985 0.180667
R19489 VDAC_P.n987 VDAC_P.n986 0.180667
R19490 VDAC_P.n988 VDAC_P.n987 0.180667
R19491 VDAC_P.n989 VDAC_P.n988 0.180667
R19492 VDAC_P.n990 VDAC_P.n989 0.180667
R19493 VDAC_P.n991 VDAC_P.n990 0.180667
R19494 VDAC_P.n992 VDAC_P.n991 0.180667
R19495 VDAC_P.n993 VDAC_P.n992 0.180667
R19496 VDAC_P.n994 VDAC_P.n993 0.180667
R19497 VDAC_P.n995 VDAC_P.n994 0.180667
R19498 VDAC_P.n996 VDAC_P.n995 0.180667
R19499 VDAC_P.n997 VDAC_P.n996 0.180667
R19500 VDAC_P.n998 VDAC_P.n997 0.180667
R19501 VDAC_P.n999 VDAC_P.n102 0.180667
R19502 VDAC_P.n1000 VDAC_P.n999 0.180667
R19503 VDAC_P.n1001 VDAC_P.n1000 0.180667
R19504 VDAC_P.n1002 VDAC_P.n1001 0.180667
R19505 VDAC_P.n1003 VDAC_P.n1002 0.180667
R19506 VDAC_P.n1004 VDAC_P.n1003 0.180667
R19507 VDAC_P.n1005 VDAC_P.n1004 0.180667
R19508 VDAC_P.n1006 VDAC_P.n1005 0.180667
R19509 VDAC_P.n1007 VDAC_P.n1006 0.180667
R19510 VDAC_P.n1008 VDAC_P.n1007 0.180667
R19511 VDAC_P.n1009 VDAC_P.n1008 0.180667
R19512 VDAC_P.n1010 VDAC_P.n1009 0.180667
R19513 VDAC_P.n1011 VDAC_P.n1010 0.180667
R19514 VDAC_P.n1012 VDAC_P.n1011 0.180667
R19515 VDAC_P.n1013 VDAC_P.n1012 0.180667
R19516 VDAC_P.n1014 VDAC_P.n1013 0.180667
R19517 VDAC_P.n1015 VDAC_P.n1014 0.180667
R19518 VDAC_P.n1016 VDAC_P.n1015 0.180667
R19519 VDAC_P.n1017 VDAC_P.n1016 0.180667
R19520 VDAC_P.n1018 VDAC_P.n1017 0.180667
R19521 VDAC_P.n1019 VDAC_P.n1018 0.180667
R19522 VDAC_P.n1020 VDAC_P.n1019 0.180667
R19523 VDAC_P.n1021 VDAC_P.n1020 0.180667
R19524 VDAC_P.n1022 VDAC_P.n1021 0.180667
R19525 VDAC_P.n1023 VDAC_P.n1022 0.180667
R19526 VDAC_P.n1024 VDAC_P.n1023 0.180667
R19527 VDAC_P.n1025 VDAC_P.n1024 0.180667
R19528 VDAC_P.n1026 VDAC_P.n1025 0.180667
R19529 VDAC_P.n1027 VDAC_P.n1026 0.180667
R19530 VDAC_P.n1028 VDAC_P.n1027 0.180667
R19531 VDAC_P.n1029 VDAC_P.n1028 0.180667
R19532 VDAC_P.n1030 VDAC_P.n1029 0.180667
R19533 VDAC_P.n1031 VDAC_P.n1030 0.180667
R19534 VDAC_P.n1032 VDAC_P.n1031 0.180667
R19535 VDAC_P.n1033 VDAC_P.n1032 0.180667
R19536 VDAC_P.n1034 VDAC_P.n1033 0.180667
R19537 VDAC_P.n1035 VDAC_P.n1034 0.180667
R19538 VDAC_P.n1036 VDAC_P.n1035 0.180667
R19539 VDAC_P.n1037 VDAC_P.n1036 0.180667
R19540 VDAC_P.n1038 VDAC_P.n1037 0.180667
R19541 VDAC_P.n1039 VDAC_P.n1038 0.180667
R19542 VDAC_P.n1040 VDAC_P.n1039 0.180667
R19543 VDAC_P.n1041 VDAC_P.n1040 0.180667
R19544 VDAC_P.n1042 VDAC_P.n1041 0.180667
R19545 VDAC_P.n1043 VDAC_P.n1042 0.180667
R19546 VDAC_P.n1044 VDAC_P.n1043 0.180667
R19547 VDAC_P.n1045 VDAC_P.n1044 0.180667
R19548 VDAC_P.n1046 VDAC_P.n1045 0.180667
R19549 VDAC_P.n1047 VDAC_P.n1046 0.180667
R19550 VDAC_P.n1048 VDAC_P.n1047 0.180667
R19551 VDAC_P.n1049 VDAC_P.n1048 0.180667
R19552 VDAC_P.n1050 VDAC_P.n1049 0.180667
R19553 VDAC_P.n1051 VDAC_P.n1050 0.180667
R19554 VDAC_P.n1052 VDAC_P.n1051 0.180667
R19555 VDAC_P.n1053 VDAC_P.n1052 0.180667
R19556 VDAC_P.n1054 VDAC_P.n1053 0.180667
R19557 VDAC_P.n1055 VDAC_P.n1054 0.180667
R19558 VDAC_P.n1056 VDAC_P.n1055 0.180667
R19559 VDAC_P.n1057 VDAC_P.n1056 0.180667
R19560 VDAC_P.n1058 VDAC_P.n1057 0.180667
R19561 VDAC_P.n1059 VDAC_P.n1058 0.180667
R19562 VDAC_P.n1060 VDAC_P.n1059 0.180667
R19563 VDAC_P.n1061 VDAC_P.n1060 0.180667
R19564 VDAC_P.n1062 VDAC_P.n101 0.180667
R19565 VDAC_P.n1063 VDAC_P.n1062 0.180667
R19566 VDAC_P.n1064 VDAC_P.n1063 0.180667
R19567 VDAC_P.n1065 VDAC_P.n1064 0.180667
R19568 VDAC_P.n1066 VDAC_P.n1065 0.180667
R19569 VDAC_P.n1067 VDAC_P.n1066 0.180667
R19570 VDAC_P.n1068 VDAC_P.n1067 0.180667
R19571 VDAC_P.n1069 VDAC_P.n1068 0.180667
R19572 VDAC_P.n1070 VDAC_P.n1069 0.180667
R19573 VDAC_P.n1071 VDAC_P.n1070 0.180667
R19574 VDAC_P.n1072 VDAC_P.n1071 0.180667
R19575 VDAC_P.n1073 VDAC_P.n1072 0.180667
R19576 VDAC_P.n1074 VDAC_P.n1073 0.180667
R19577 VDAC_P.n1075 VDAC_P.n1074 0.180667
R19578 VDAC_P.n1076 VDAC_P.n1075 0.180667
R19579 VDAC_P.n1077 VDAC_P.n1076 0.180667
R19580 VDAC_P.n1078 VDAC_P.n1077 0.180667
R19581 VDAC_P.n1079 VDAC_P.n1078 0.180667
R19582 VDAC_P.n1080 VDAC_P.n1079 0.180667
R19583 VDAC_P.n1081 VDAC_P.n1080 0.180667
R19584 VDAC_P.n1082 VDAC_P.n1081 0.180667
R19585 VDAC_P.n1083 VDAC_P.n1082 0.180667
R19586 VDAC_P.n1084 VDAC_P.n1083 0.180667
R19587 VDAC_P.n1085 VDAC_P.n1084 0.180667
R19588 VDAC_P.n1086 VDAC_P.n1085 0.180667
R19589 VDAC_P.n1087 VDAC_P.n1086 0.180667
R19590 VDAC_P.n1088 VDAC_P.n1087 0.180667
R19591 VDAC_P.n1089 VDAC_P.n1088 0.180667
R19592 VDAC_P.n1090 VDAC_P.n1089 0.180667
R19593 VDAC_P.n1091 VDAC_P.n1090 0.180667
R19594 VDAC_P.n1092 VDAC_P.n1091 0.180667
R19595 VDAC_P.n1093 VDAC_P.n1092 0.180667
R19596 VDAC_P.n1094 VDAC_P.n1093 0.180667
R19597 VDAC_P.n1095 VDAC_P.n1094 0.180667
R19598 VDAC_P.n1096 VDAC_P.n1095 0.180667
R19599 VDAC_P.n1097 VDAC_P.n1096 0.180667
R19600 VDAC_P.n1098 VDAC_P.n1097 0.180667
R19601 VDAC_P.n1099 VDAC_P.n1098 0.180667
R19602 VDAC_P.n1100 VDAC_P.n1099 0.180667
R19603 VDAC_P.n1101 VDAC_P.n1100 0.180667
R19604 VDAC_P.n1102 VDAC_P.n1101 0.180667
R19605 VDAC_P.n1103 VDAC_P.n1102 0.180667
R19606 VDAC_P.n1104 VDAC_P.n1103 0.180667
R19607 VDAC_P.n1105 VDAC_P.n1104 0.180667
R19608 VDAC_P.n1106 VDAC_P.n1105 0.180667
R19609 VDAC_P.n1107 VDAC_P.n1106 0.180667
R19610 VDAC_P.n1108 VDAC_P.n1107 0.180667
R19611 VDAC_P.n1109 VDAC_P.n1108 0.180667
R19612 VDAC_P.n1110 VDAC_P.n1109 0.180667
R19613 VDAC_P.n1111 VDAC_P.n1110 0.180667
R19614 VDAC_P.n1112 VDAC_P.n1111 0.180667
R19615 VDAC_P.n1113 VDAC_P.n1112 0.180667
R19616 VDAC_P.n1114 VDAC_P.n1113 0.180667
R19617 VDAC_P.n1115 VDAC_P.n1114 0.180667
R19618 VDAC_P.n1116 VDAC_P.n1115 0.180667
R19619 VDAC_P.n1117 VDAC_P.n1116 0.180667
R19620 VDAC_P.n1118 VDAC_P.n1117 0.180667
R19621 VDAC_P.n1119 VDAC_P.n1118 0.180667
R19622 VDAC_P.n1120 VDAC_P.n1119 0.180667
R19623 VDAC_P.n1121 VDAC_P.n1120 0.180667
R19624 VDAC_P.n1122 VDAC_P.n1121 0.180667
R19625 VDAC_P.n1123 VDAC_P.n1122 0.180667
R19626 VDAC_P.n1124 VDAC_P.n1123 0.180667
R19627 VDAC_P.n1125 VDAC_P.n100 0.180667
R19628 VDAC_P.n1126 VDAC_P.n1125 0.180667
R19629 VDAC_P.n1127 VDAC_P.n1126 0.180667
R19630 VDAC_P.n1128 VDAC_P.n1127 0.180667
R19631 VDAC_P.n1129 VDAC_P.n1128 0.180667
R19632 VDAC_P.n1130 VDAC_P.n1129 0.180667
R19633 VDAC_P.n1131 VDAC_P.n1130 0.180667
R19634 VDAC_P.n1132 VDAC_P.n1131 0.180667
R19635 VDAC_P.n1133 VDAC_P.n1132 0.180667
R19636 VDAC_P.n1134 VDAC_P.n1133 0.180667
R19637 VDAC_P.n1135 VDAC_P.n1134 0.180667
R19638 VDAC_P.n1136 VDAC_P.n1135 0.180667
R19639 VDAC_P.n1137 VDAC_P.n1136 0.180667
R19640 VDAC_P.n1138 VDAC_P.n1137 0.180667
R19641 VDAC_P.n1139 VDAC_P.n1138 0.180667
R19642 VDAC_P.n1140 VDAC_P.n1139 0.180667
R19643 VDAC_P.n1141 VDAC_P.n1140 0.180667
R19644 VDAC_P.n1142 VDAC_P.n1141 0.180667
R19645 VDAC_P.n1143 VDAC_P.n1142 0.180667
R19646 VDAC_P.n1144 VDAC_P.n1143 0.180667
R19647 VDAC_P.n1145 VDAC_P.n1144 0.180667
R19648 VDAC_P.n1146 VDAC_P.n1145 0.180667
R19649 VDAC_P.n1147 VDAC_P.n1146 0.180667
R19650 VDAC_P.n1148 VDAC_P.n1147 0.180667
R19651 VDAC_P.n1149 VDAC_P.n1148 0.180667
R19652 VDAC_P.n1150 VDAC_P.n1149 0.180667
R19653 VDAC_P.n1151 VDAC_P.n1150 0.180667
R19654 VDAC_P.n1152 VDAC_P.n1151 0.180667
R19655 VDAC_P.n1153 VDAC_P.n1152 0.180667
R19656 VDAC_P.n1154 VDAC_P.n1153 0.180667
R19657 VDAC_P.n1155 VDAC_P.n1154 0.180667
R19658 VDAC_P.n1156 VDAC_P.n1155 0.180667
R19659 VDAC_P.n1157 VDAC_P.n1156 0.180667
R19660 VDAC_P.n1158 VDAC_P.n1157 0.180667
R19661 VDAC_P.n1159 VDAC_P.n1158 0.180667
R19662 VDAC_P.n1160 VDAC_P.n1159 0.180667
R19663 VDAC_P.n1161 VDAC_P.n1160 0.180667
R19664 VDAC_P.n1162 VDAC_P.n1161 0.180667
R19665 VDAC_P.n1163 VDAC_P.n1162 0.180667
R19666 VDAC_P.n1164 VDAC_P.n1163 0.180667
R19667 VDAC_P.n1165 VDAC_P.n1164 0.180667
R19668 VDAC_P.n1166 VDAC_P.n1165 0.180667
R19669 VDAC_P.n1167 VDAC_P.n1166 0.180667
R19670 VDAC_P.n1168 VDAC_P.n1167 0.180667
R19671 VDAC_P.n1169 VDAC_P.n1168 0.180667
R19672 VDAC_P.n1170 VDAC_P.n1169 0.180667
R19673 VDAC_P.n1171 VDAC_P.n1170 0.180667
R19674 VDAC_P.n1172 VDAC_P.n1171 0.180667
R19675 VDAC_P.n1173 VDAC_P.n1172 0.180667
R19676 VDAC_P.n1174 VDAC_P.n1173 0.180667
R19677 VDAC_P.n1175 VDAC_P.n1174 0.180667
R19678 VDAC_P.n1176 VDAC_P.n1175 0.180667
R19679 VDAC_P.n1177 VDAC_P.n1176 0.180667
R19680 VDAC_P.n1178 VDAC_P.n1177 0.180667
R19681 VDAC_P.n1179 VDAC_P.n1178 0.180667
R19682 VDAC_P.n1180 VDAC_P.n1179 0.180667
R19683 VDAC_P.n1181 VDAC_P.n1180 0.180667
R19684 VDAC_P.n1182 VDAC_P.n1181 0.180667
R19685 VDAC_P.n1183 VDAC_P.n1182 0.180667
R19686 VDAC_P.n1184 VDAC_P.n1183 0.180667
R19687 VDAC_P.n1185 VDAC_P.n1184 0.180667
R19688 VDAC_P.n1186 VDAC_P.n1185 0.180667
R19689 VDAC_P.n1187 VDAC_P.n1186 0.180667
R19690 VDAC_P.n1188 VDAC_P.n99 0.180667
R19691 VDAC_P.n1189 VDAC_P.n1188 0.180667
R19692 VDAC_P.n1190 VDAC_P.n1189 0.180667
R19693 VDAC_P.n1191 VDAC_P.n1190 0.180667
R19694 VDAC_P.n1192 VDAC_P.n1191 0.180667
R19695 VDAC_P.n1193 VDAC_P.n1192 0.180667
R19696 VDAC_P.n1194 VDAC_P.n1193 0.180667
R19697 VDAC_P.n1195 VDAC_P.n1194 0.180667
R19698 VDAC_P.n1196 VDAC_P.n1195 0.180667
R19699 VDAC_P.n1197 VDAC_P.n1196 0.180667
R19700 VDAC_P.n1198 VDAC_P.n1197 0.180667
R19701 VDAC_P.n1199 VDAC_P.n1198 0.180667
R19702 VDAC_P.n1200 VDAC_P.n1199 0.180667
R19703 VDAC_P.n1201 VDAC_P.n1200 0.180667
R19704 VDAC_P.n1202 VDAC_P.n1201 0.180667
R19705 VDAC_P.n1203 VDAC_P.n1202 0.180667
R19706 VDAC_P.n1204 VDAC_P.n1203 0.180667
R19707 VDAC_P.n1205 VDAC_P.n1204 0.180667
R19708 VDAC_P.n1206 VDAC_P.n1205 0.180667
R19709 VDAC_P.n1207 VDAC_P.n1206 0.180667
R19710 VDAC_P.n1208 VDAC_P.n1207 0.180667
R19711 VDAC_P.n1209 VDAC_P.n1208 0.180667
R19712 VDAC_P.n1210 VDAC_P.n1209 0.180667
R19713 VDAC_P.n1211 VDAC_P.n1210 0.180667
R19714 VDAC_P.n1212 VDAC_P.n1211 0.180667
R19715 VDAC_P.n1213 VDAC_P.n1212 0.180667
R19716 VDAC_P.n1214 VDAC_P.n1213 0.180667
R19717 VDAC_P.n1215 VDAC_P.n1214 0.180667
R19718 VDAC_P.n1216 VDAC_P.n1215 0.180667
R19719 VDAC_P.n1217 VDAC_P.n1216 0.180667
R19720 VDAC_P.n1218 VDAC_P.n1217 0.180667
R19721 VDAC_P.n1219 VDAC_P.n1218 0.180667
R19722 VDAC_P.n1220 VDAC_P.n1219 0.180667
R19723 VDAC_P.n1221 VDAC_P.n1220 0.180667
R19724 VDAC_P.n1222 VDAC_P.n1221 0.180667
R19725 VDAC_P.n1223 VDAC_P.n1222 0.180667
R19726 VDAC_P.n1224 VDAC_P.n1223 0.180667
R19727 VDAC_P.n1225 VDAC_P.n1224 0.180667
R19728 VDAC_P.n1226 VDAC_P.n1225 0.180667
R19729 VDAC_P.n1227 VDAC_P.n1226 0.180667
R19730 VDAC_P.n1228 VDAC_P.n1227 0.180667
R19731 VDAC_P.n1229 VDAC_P.n1228 0.180667
R19732 VDAC_P.n1230 VDAC_P.n1229 0.180667
R19733 VDAC_P.n1231 VDAC_P.n1230 0.180667
R19734 VDAC_P.n1232 VDAC_P.n1231 0.180667
R19735 VDAC_P.n1233 VDAC_P.n1232 0.180667
R19736 VDAC_P.n1234 VDAC_P.n1233 0.180667
R19737 VDAC_P.n1235 VDAC_P.n1234 0.180667
R19738 VDAC_P.n1236 VDAC_P.n1235 0.180667
R19739 VDAC_P.n1237 VDAC_P.n1236 0.180667
R19740 VDAC_P.n1238 VDAC_P.n1237 0.180667
R19741 VDAC_P.n1239 VDAC_P.n1238 0.180667
R19742 VDAC_P.n1240 VDAC_P.n1239 0.180667
R19743 VDAC_P.n1241 VDAC_P.n1240 0.180667
R19744 VDAC_P.n1242 VDAC_P.n1241 0.180667
R19745 VDAC_P.n1243 VDAC_P.n1242 0.180667
R19746 VDAC_P.n1244 VDAC_P.n1243 0.180667
R19747 VDAC_P.n1245 VDAC_P.n1244 0.180667
R19748 VDAC_P.n1246 VDAC_P.n1245 0.180667
R19749 VDAC_P.n1247 VDAC_P.n1246 0.180667
R19750 VDAC_P.n1248 VDAC_P.n1247 0.180667
R19751 VDAC_P.n1249 VDAC_P.n1248 0.180667
R19752 VDAC_P.n1250 VDAC_P.n1249 0.180667
R19753 VDAC_P.n1251 VDAC_P.n98 0.180667
R19754 VDAC_P.n1252 VDAC_P.n1251 0.180667
R19755 VDAC_P.n1253 VDAC_P.n1252 0.180667
R19756 VDAC_P.n1254 VDAC_P.n1253 0.180667
R19757 VDAC_P.n1255 VDAC_P.n1254 0.180667
R19758 VDAC_P.n1256 VDAC_P.n1255 0.180667
R19759 VDAC_P.n1257 VDAC_P.n1256 0.180667
R19760 VDAC_P.n1258 VDAC_P.n1257 0.180667
R19761 VDAC_P.n1259 VDAC_P.n1258 0.180667
R19762 VDAC_P.n1260 VDAC_P.n1259 0.180667
R19763 VDAC_P.n1261 VDAC_P.n1260 0.180667
R19764 VDAC_P.n1262 VDAC_P.n1261 0.180667
R19765 VDAC_P.n1263 VDAC_P.n1262 0.180667
R19766 VDAC_P.n1264 VDAC_P.n1263 0.180667
R19767 VDAC_P.n1265 VDAC_P.n1264 0.180667
R19768 VDAC_P.n1266 VDAC_P.n1265 0.180667
R19769 VDAC_P.n1267 VDAC_P.n1266 0.180667
R19770 VDAC_P.n1268 VDAC_P.n1267 0.180667
R19771 VDAC_P.n1269 VDAC_P.n1268 0.180667
R19772 VDAC_P.n1270 VDAC_P.n1269 0.180667
R19773 VDAC_P.n1271 VDAC_P.n1270 0.180667
R19774 VDAC_P.n1272 VDAC_P.n1271 0.180667
R19775 VDAC_P.n1273 VDAC_P.n1272 0.180667
R19776 VDAC_P.n1274 VDAC_P.n1273 0.180667
R19777 VDAC_P.n1275 VDAC_P.n1274 0.180667
R19778 VDAC_P.n1276 VDAC_P.n1275 0.180667
R19779 VDAC_P.n1277 VDAC_P.n1276 0.180667
R19780 VDAC_P.n1278 VDAC_P.n1277 0.180667
R19781 VDAC_P.n1279 VDAC_P.n1278 0.180667
R19782 VDAC_P.n1280 VDAC_P.n1279 0.180667
R19783 VDAC_P.n1281 VDAC_P.n1280 0.180667
R19784 VDAC_P.n1282 VDAC_P.n1281 0.180667
R19785 VDAC_P.n1283 VDAC_P.n1282 0.180667
R19786 VDAC_P.n1284 VDAC_P.n1283 0.180667
R19787 VDAC_P.n1285 VDAC_P.n1284 0.180667
R19788 VDAC_P.n1286 VDAC_P.n1285 0.180667
R19789 VDAC_P.n1287 VDAC_P.n1286 0.180667
R19790 VDAC_P.n1288 VDAC_P.n1287 0.180667
R19791 VDAC_P.n1289 VDAC_P.n1288 0.180667
R19792 VDAC_P.n1290 VDAC_P.n1289 0.180667
R19793 VDAC_P.n1291 VDAC_P.n1290 0.180667
R19794 VDAC_P.n1292 VDAC_P.n1291 0.180667
R19795 VDAC_P.n1293 VDAC_P.n1292 0.180667
R19796 VDAC_P.n1294 VDAC_P.n1293 0.180667
R19797 VDAC_P.n1295 VDAC_P.n1294 0.180667
R19798 VDAC_P.n1296 VDAC_P.n1295 0.180667
R19799 VDAC_P.n1297 VDAC_P.n1296 0.180667
R19800 VDAC_P.n1298 VDAC_P.n1297 0.180667
R19801 VDAC_P.n1299 VDAC_P.n1298 0.180667
R19802 VDAC_P.n1300 VDAC_P.n1299 0.180667
R19803 VDAC_P.n1301 VDAC_P.n1300 0.180667
R19804 VDAC_P.n1302 VDAC_P.n1301 0.180667
R19805 VDAC_P.n1303 VDAC_P.n1302 0.180667
R19806 VDAC_P.n1304 VDAC_P.n1303 0.180667
R19807 VDAC_P.n1305 VDAC_P.n1304 0.180667
R19808 VDAC_P.n1306 VDAC_P.n1305 0.180667
R19809 VDAC_P.n1307 VDAC_P.n1306 0.180667
R19810 VDAC_P.n1308 VDAC_P.n1307 0.180667
R19811 VDAC_P.n1309 VDAC_P.n1308 0.180667
R19812 VDAC_P.n1310 VDAC_P.n1309 0.180667
R19813 VDAC_P.n1311 VDAC_P.n1310 0.180667
R19814 VDAC_P.n1312 VDAC_P.n1311 0.180667
R19815 VDAC_P.n1313 VDAC_P.n1312 0.180667
R19816 VDAC_P.n1314 VDAC_P.n97 0.180667
R19817 VDAC_P.n1315 VDAC_P.n1314 0.180667
R19818 VDAC_P.n1316 VDAC_P.n1315 0.180667
R19819 VDAC_P.n1317 VDAC_P.n1316 0.180667
R19820 VDAC_P.n1318 VDAC_P.n1317 0.180667
R19821 VDAC_P.n1319 VDAC_P.n1318 0.180667
R19822 VDAC_P.n1320 VDAC_P.n1319 0.180667
R19823 VDAC_P.n1321 VDAC_P.n1320 0.180667
R19824 VDAC_P.n1322 VDAC_P.n1321 0.180667
R19825 VDAC_P.n1323 VDAC_P.n1322 0.180667
R19826 VDAC_P.n1324 VDAC_P.n1323 0.180667
R19827 VDAC_P.n1325 VDAC_P.n1324 0.180667
R19828 VDAC_P.n1326 VDAC_P.n1325 0.180667
R19829 VDAC_P.n1327 VDAC_P.n1326 0.180667
R19830 VDAC_P.n1328 VDAC_P.n1327 0.180667
R19831 VDAC_P.n1329 VDAC_P.n1328 0.180667
R19832 VDAC_P.n1330 VDAC_P.n1329 0.180667
R19833 VDAC_P.n1331 VDAC_P.n1330 0.180667
R19834 VDAC_P.n1332 VDAC_P.n1331 0.180667
R19835 VDAC_P.n1333 VDAC_P.n1332 0.180667
R19836 VDAC_P.n1334 VDAC_P.n1333 0.180667
R19837 VDAC_P.n1335 VDAC_P.n1334 0.180667
R19838 VDAC_P.n1336 VDAC_P.n1335 0.180667
R19839 VDAC_P.n1337 VDAC_P.n1336 0.180667
R19840 VDAC_P.n1338 VDAC_P.n1337 0.180667
R19841 VDAC_P.n1339 VDAC_P.n1338 0.180667
R19842 VDAC_P.n1340 VDAC_P.n1339 0.180667
R19843 VDAC_P.n1341 VDAC_P.n1340 0.180667
R19844 VDAC_P.n1342 VDAC_P.n1341 0.180667
R19845 VDAC_P.n1343 VDAC_P.n1342 0.180667
R19846 VDAC_P.n1344 VDAC_P.n1343 0.180667
R19847 VDAC_P.n1345 VDAC_P.n1344 0.180667
R19848 VDAC_P.n1346 VDAC_P.n1345 0.180667
R19849 VDAC_P.n1347 VDAC_P.n1346 0.180667
R19850 VDAC_P.n1348 VDAC_P.n1347 0.180667
R19851 VDAC_P.n1349 VDAC_P.n1348 0.180667
R19852 VDAC_P.n1350 VDAC_P.n1349 0.180667
R19853 VDAC_P.n1351 VDAC_P.n1350 0.180667
R19854 VDAC_P.n1352 VDAC_P.n1351 0.180667
R19855 VDAC_P.n1353 VDAC_P.n1352 0.180667
R19856 VDAC_P.n1354 VDAC_P.n1353 0.180667
R19857 VDAC_P.n1355 VDAC_P.n1354 0.180667
R19858 VDAC_P.n1356 VDAC_P.n1355 0.180667
R19859 VDAC_P.n1357 VDAC_P.n1356 0.180667
R19860 VDAC_P.n1358 VDAC_P.n1357 0.180667
R19861 VDAC_P.n1359 VDAC_P.n1358 0.180667
R19862 VDAC_P.n1360 VDAC_P.n1359 0.180667
R19863 VDAC_P.n1361 VDAC_P.n1360 0.180667
R19864 VDAC_P.n1362 VDAC_P.n1361 0.180667
R19865 VDAC_P.n1363 VDAC_P.n1362 0.180667
R19866 VDAC_P.n1364 VDAC_P.n1363 0.180667
R19867 VDAC_P.n1365 VDAC_P.n1364 0.180667
R19868 VDAC_P.n1366 VDAC_P.n1365 0.180667
R19869 VDAC_P.n1367 VDAC_P.n1366 0.180667
R19870 VDAC_P.n1368 VDAC_P.n1367 0.180667
R19871 VDAC_P.n1369 VDAC_P.n1368 0.180667
R19872 VDAC_P.n1370 VDAC_P.n1369 0.180667
R19873 VDAC_P.n1371 VDAC_P.n1370 0.180667
R19874 VDAC_P.n1372 VDAC_P.n1371 0.180667
R19875 VDAC_P.n1373 VDAC_P.n1372 0.180667
R19876 VDAC_P.n1374 VDAC_P.n1373 0.180667
R19877 VDAC_P.n1375 VDAC_P.n1374 0.180667
R19878 VDAC_P.n1376 VDAC_P.n1375 0.180667
R19879 VDAC_P.n1377 VDAC_P.n96 0.180667
R19880 VDAC_P.n1378 VDAC_P.n1377 0.180667
R19881 VDAC_P.n1379 VDAC_P.n1378 0.180667
R19882 VDAC_P.n1380 VDAC_P.n1379 0.180667
R19883 VDAC_P.n1381 VDAC_P.n1380 0.180667
R19884 VDAC_P.n1382 VDAC_P.n1381 0.180667
R19885 VDAC_P.n1383 VDAC_P.n1382 0.180667
R19886 VDAC_P.n1384 VDAC_P.n1383 0.180667
R19887 VDAC_P.n1385 VDAC_P.n1384 0.180667
R19888 VDAC_P.n1386 VDAC_P.n1385 0.180667
R19889 VDAC_P.n1387 VDAC_P.n1386 0.180667
R19890 VDAC_P.n1388 VDAC_P.n1387 0.180667
R19891 VDAC_P.n1389 VDAC_P.n1388 0.180667
R19892 VDAC_P.n1390 VDAC_P.n1389 0.180667
R19893 VDAC_P.n1391 VDAC_P.n1390 0.180667
R19894 VDAC_P.n1392 VDAC_P.n1391 0.180667
R19895 VDAC_P.n1393 VDAC_P.n1392 0.180667
R19896 VDAC_P.n1394 VDAC_P.n1393 0.180667
R19897 VDAC_P.n1395 VDAC_P.n1394 0.180667
R19898 VDAC_P.n1396 VDAC_P.n1395 0.180667
R19899 VDAC_P.n1397 VDAC_P.n1396 0.180667
R19900 VDAC_P.n1398 VDAC_P.n1397 0.180667
R19901 VDAC_P.n1399 VDAC_P.n1398 0.180667
R19902 VDAC_P.n1400 VDAC_P.n1399 0.180667
R19903 VDAC_P.n1401 VDAC_P.n1400 0.180667
R19904 VDAC_P.n1402 VDAC_P.n1401 0.180667
R19905 VDAC_P.n1403 VDAC_P.n1402 0.180667
R19906 VDAC_P.n1404 VDAC_P.n1403 0.180667
R19907 VDAC_P.n1405 VDAC_P.n1404 0.180667
R19908 VDAC_P.n1406 VDAC_P.n1405 0.180667
R19909 VDAC_P.n1407 VDAC_P.n1406 0.180667
R19910 VDAC_P.n1408 VDAC_P.n1407 0.180667
R19911 VDAC_P.n1409 VDAC_P.n1408 0.180667
R19912 VDAC_P.n1410 VDAC_P.n1409 0.180667
R19913 VDAC_P.n1411 VDAC_P.n1410 0.180667
R19914 VDAC_P.n1412 VDAC_P.n1411 0.180667
R19915 VDAC_P.n1413 VDAC_P.n1412 0.180667
R19916 VDAC_P.n1414 VDAC_P.n1413 0.180667
R19917 VDAC_P.n1415 VDAC_P.n1414 0.180667
R19918 VDAC_P.n1416 VDAC_P.n1415 0.180667
R19919 VDAC_P.n1417 VDAC_P.n1416 0.180667
R19920 VDAC_P.n1418 VDAC_P.n1417 0.180667
R19921 VDAC_P.n1419 VDAC_P.n1418 0.180667
R19922 VDAC_P.n1420 VDAC_P.n1419 0.180667
R19923 VDAC_P.n1421 VDAC_P.n1420 0.180667
R19924 VDAC_P.n1422 VDAC_P.n1421 0.180667
R19925 VDAC_P.n1423 VDAC_P.n1422 0.180667
R19926 VDAC_P.n1424 VDAC_P.n1423 0.180667
R19927 VDAC_P.n1425 VDAC_P.n1424 0.180667
R19928 VDAC_P.n1426 VDAC_P.n1425 0.180667
R19929 VDAC_P.n1427 VDAC_P.n1426 0.180667
R19930 VDAC_P.n1428 VDAC_P.n1427 0.180667
R19931 VDAC_P.n1429 VDAC_P.n1428 0.180667
R19932 VDAC_P.n1430 VDAC_P.n1429 0.180667
R19933 VDAC_P.n1431 VDAC_P.n1430 0.180667
R19934 VDAC_P.n1432 VDAC_P.n1431 0.180667
R19935 VDAC_P.n1433 VDAC_P.n1432 0.180667
R19936 VDAC_P.n1434 VDAC_P.n1433 0.180667
R19937 VDAC_P.n1435 VDAC_P.n1434 0.180667
R19938 VDAC_P.n1436 VDAC_P.n1435 0.180667
R19939 VDAC_P.n1437 VDAC_P.n1436 0.180667
R19940 VDAC_P.n1438 VDAC_P.n1437 0.180667
R19941 VDAC_P.n1439 VDAC_P.n1438 0.180667
R19942 VDAC_P.n1440 VDAC_P.n95 0.180667
R19943 VDAC_P.n1441 VDAC_P.n1440 0.180667
R19944 VDAC_P.n1442 VDAC_P.n1441 0.180667
R19945 VDAC_P.n1443 VDAC_P.n1442 0.180667
R19946 VDAC_P.n1444 VDAC_P.n1443 0.180667
R19947 VDAC_P.n1445 VDAC_P.n1444 0.180667
R19948 VDAC_P.n1446 VDAC_P.n1445 0.180667
R19949 VDAC_P.n1447 VDAC_P.n1446 0.180667
R19950 VDAC_P.n1448 VDAC_P.n1447 0.180667
R19951 VDAC_P.n1449 VDAC_P.n1448 0.180667
R19952 VDAC_P.n1450 VDAC_P.n1449 0.180667
R19953 VDAC_P.n1451 VDAC_P.n1450 0.180667
R19954 VDAC_P.n1452 VDAC_P.n1451 0.180667
R19955 VDAC_P.n1453 VDAC_P.n1452 0.180667
R19956 VDAC_P.n1454 VDAC_P.n1453 0.180667
R19957 VDAC_P.n1455 VDAC_P.n1454 0.180667
R19958 VDAC_P.n1456 VDAC_P.n1455 0.180667
R19959 VDAC_P.n1457 VDAC_P.n1456 0.180667
R19960 VDAC_P.n1458 VDAC_P.n1457 0.180667
R19961 VDAC_P.n1459 VDAC_P.n1458 0.180667
R19962 VDAC_P.n1460 VDAC_P.n1459 0.180667
R19963 VDAC_P.n1461 VDAC_P.n1460 0.180667
R19964 VDAC_P.n1462 VDAC_P.n1461 0.180667
R19965 VDAC_P.n1463 VDAC_P.n1462 0.180667
R19966 VDAC_P.n1464 VDAC_P.n1463 0.180667
R19967 VDAC_P.n1465 VDAC_P.n1464 0.180667
R19968 VDAC_P.n1466 VDAC_P.n1465 0.180667
R19969 VDAC_P.n1467 VDAC_P.n1466 0.180667
R19970 VDAC_P.n1468 VDAC_P.n1467 0.180667
R19971 VDAC_P.n1469 VDAC_P.n1468 0.180667
R19972 VDAC_P.n1470 VDAC_P.n1469 0.180667
R19973 VDAC_P.n1471 VDAC_P.n1470 0.180667
R19974 VDAC_P.n1472 VDAC_P.n1471 0.180667
R19975 VDAC_P.n1473 VDAC_P.n1472 0.180667
R19976 VDAC_P.n1474 VDAC_P.n1473 0.180667
R19977 VDAC_P.n1475 VDAC_P.n1474 0.180667
R19978 VDAC_P.n1476 VDAC_P.n1475 0.180667
R19979 VDAC_P.n1477 VDAC_P.n1476 0.180667
R19980 VDAC_P.n1478 VDAC_P.n1477 0.180667
R19981 VDAC_P.n1479 VDAC_P.n1478 0.180667
R19982 VDAC_P.n1480 VDAC_P.n1479 0.180667
R19983 VDAC_P.n1481 VDAC_P.n1480 0.180667
R19984 VDAC_P.n1482 VDAC_P.n1481 0.180667
R19985 VDAC_P.n1483 VDAC_P.n1482 0.180667
R19986 VDAC_P.n1484 VDAC_P.n1483 0.180667
R19987 VDAC_P.n1485 VDAC_P.n1484 0.180667
R19988 VDAC_P.n1486 VDAC_P.n1485 0.180667
R19989 VDAC_P.n1487 VDAC_P.n1486 0.180667
R19990 VDAC_P.n1488 VDAC_P.n1487 0.180667
R19991 VDAC_P.n1489 VDAC_P.n1488 0.180667
R19992 VDAC_P.n1490 VDAC_P.n1489 0.180667
R19993 VDAC_P.n1491 VDAC_P.n1490 0.180667
R19994 VDAC_P.n1492 VDAC_P.n1491 0.180667
R19995 VDAC_P.n1493 VDAC_P.n1492 0.180667
R19996 VDAC_P.n1494 VDAC_P.n1493 0.180667
R19997 VDAC_P.n1495 VDAC_P.n1494 0.180667
R19998 VDAC_P.n1496 VDAC_P.n1495 0.180667
R19999 VDAC_P.n1497 VDAC_P.n1496 0.180667
R20000 VDAC_P.n1498 VDAC_P.n1497 0.180667
R20001 VDAC_P.n1499 VDAC_P.n1498 0.180667
R20002 VDAC_P.n1500 VDAC_P.n1499 0.180667
R20003 VDAC_P.n1501 VDAC_P.n1500 0.180667
R20004 VDAC_P.n1502 VDAC_P.n1501 0.180667
R20005 VDAC_P.n1503 VDAC_P.n94 0.180667
R20006 VDAC_P.n1504 VDAC_P.n1503 0.180667
R20007 VDAC_P.n1505 VDAC_P.n1504 0.180667
R20008 VDAC_P.n1506 VDAC_P.n1505 0.180667
R20009 VDAC_P.n1507 VDAC_P.n1506 0.180667
R20010 VDAC_P.n1508 VDAC_P.n1507 0.180667
R20011 VDAC_P.n1509 VDAC_P.n1508 0.180667
R20012 VDAC_P.n1510 VDAC_P.n1509 0.180667
R20013 VDAC_P.n1511 VDAC_P.n1510 0.180667
R20014 VDAC_P.n1512 VDAC_P.n1511 0.180667
R20015 VDAC_P.n1513 VDAC_P.n1512 0.180667
R20016 VDAC_P.n1514 VDAC_P.n1513 0.180667
R20017 VDAC_P.n1515 VDAC_P.n1514 0.180667
R20018 VDAC_P.n1516 VDAC_P.n1515 0.180667
R20019 VDAC_P.n1517 VDAC_P.n1516 0.180667
R20020 VDAC_P.n1518 VDAC_P.n1517 0.180667
R20021 VDAC_P.n1519 VDAC_P.n1518 0.180667
R20022 VDAC_P.n1520 VDAC_P.n1519 0.180667
R20023 VDAC_P.n1521 VDAC_P.n1520 0.180667
R20024 VDAC_P.n1522 VDAC_P.n1521 0.180667
R20025 VDAC_P.n1523 VDAC_P.n1522 0.180667
R20026 VDAC_P.n1524 VDAC_P.n1523 0.180667
R20027 VDAC_P.n1525 VDAC_P.n1524 0.180667
R20028 VDAC_P.n1526 VDAC_P.n1525 0.180667
R20029 VDAC_P.n1527 VDAC_P.n1526 0.180667
R20030 VDAC_P.n1528 VDAC_P.n1527 0.180667
R20031 VDAC_P.n1529 VDAC_P.n1528 0.180667
R20032 VDAC_P.n1530 VDAC_P.n1529 0.180667
R20033 VDAC_P.n1531 VDAC_P.n1530 0.180667
R20034 VDAC_P.n1532 VDAC_P.n1531 0.180667
R20035 VDAC_P.n1533 VDAC_P.n1532 0.180667
R20036 VDAC_P.n1534 VDAC_P.n1533 0.180667
R20037 VDAC_P.n1535 VDAC_P.n1534 0.180667
R20038 VDAC_P.n1536 VDAC_P.n1535 0.180667
R20039 VDAC_P.n1537 VDAC_P.n1536 0.180667
R20040 VDAC_P.n1538 VDAC_P.n1537 0.180667
R20041 VDAC_P.n1539 VDAC_P.n1538 0.180667
R20042 VDAC_P.n1540 VDAC_P.n1539 0.180667
R20043 VDAC_P.n1541 VDAC_P.n1540 0.180667
R20044 VDAC_P.n1542 VDAC_P.n1541 0.180667
R20045 VDAC_P.n1543 VDAC_P.n1542 0.180667
R20046 VDAC_P.n1544 VDAC_P.n1543 0.180667
R20047 VDAC_P.n1545 VDAC_P.n1544 0.180667
R20048 VDAC_P.n1546 VDAC_P.n1545 0.180667
R20049 VDAC_P.n1547 VDAC_P.n1546 0.180667
R20050 VDAC_P.n1548 VDAC_P.n1547 0.180667
R20051 VDAC_P.n1549 VDAC_P.n1548 0.180667
R20052 VDAC_P.n1550 VDAC_P.n1549 0.180667
R20053 VDAC_P.n1551 VDAC_P.n1550 0.180667
R20054 VDAC_P.n1552 VDAC_P.n1551 0.180667
R20055 VDAC_P.n1553 VDAC_P.n1552 0.180667
R20056 VDAC_P.n1554 VDAC_P.n1553 0.180667
R20057 VDAC_P.n1555 VDAC_P.n1554 0.180667
R20058 VDAC_P.n1556 VDAC_P.n1555 0.180667
R20059 VDAC_P.n1557 VDAC_P.n1556 0.180667
R20060 VDAC_P.n1558 VDAC_P.n1557 0.180667
R20061 VDAC_P.n1559 VDAC_P.n1558 0.180667
R20062 VDAC_P.n1560 VDAC_P.n1559 0.180667
R20063 VDAC_P.n1561 VDAC_P.n1560 0.180667
R20064 VDAC_P.n1562 VDAC_P.n1561 0.180667
R20065 VDAC_P.n1563 VDAC_P.n1562 0.180667
R20066 VDAC_P.n1564 VDAC_P.n1563 0.180667
R20067 VDAC_P.n1565 VDAC_P.n1564 0.180667
R20068 VDAC_P.n1566 VDAC_P.n93 0.180667
R20069 VDAC_P.n1567 VDAC_P.n1566 0.180667
R20070 VDAC_P.n1568 VDAC_P.n1567 0.180667
R20071 VDAC_P.n1569 VDAC_P.n1568 0.180667
R20072 VDAC_P.n1570 VDAC_P.n1569 0.180667
R20073 VDAC_P.n1571 VDAC_P.n1570 0.180667
R20074 VDAC_P.n1572 VDAC_P.n1571 0.180667
R20075 VDAC_P.n1573 VDAC_P.n1572 0.180667
R20076 VDAC_P.n1574 VDAC_P.n1573 0.180667
R20077 VDAC_P.n1575 VDAC_P.n1574 0.180667
R20078 VDAC_P.n1576 VDAC_P.n1575 0.180667
R20079 VDAC_P.n1577 VDAC_P.n1576 0.180667
R20080 VDAC_P.n1578 VDAC_P.n1577 0.180667
R20081 VDAC_P.n1579 VDAC_P.n1578 0.180667
R20082 VDAC_P.n1580 VDAC_P.n1579 0.180667
R20083 VDAC_P.n1581 VDAC_P.n1580 0.180667
R20084 VDAC_P.n1582 VDAC_P.n1581 0.180667
R20085 VDAC_P.n1583 VDAC_P.n1582 0.180667
R20086 VDAC_P.n1584 VDAC_P.n1583 0.180667
R20087 VDAC_P.n1585 VDAC_P.n1584 0.180667
R20088 VDAC_P.n1586 VDAC_P.n1585 0.180667
R20089 VDAC_P.n1587 VDAC_P.n1586 0.180667
R20090 VDAC_P.n1588 VDAC_P.n1587 0.180667
R20091 VDAC_P.n1589 VDAC_P.n1588 0.180667
R20092 VDAC_P.n1590 VDAC_P.n1589 0.180667
R20093 VDAC_P.n1591 VDAC_P.n1590 0.180667
R20094 VDAC_P.n1592 VDAC_P.n1591 0.180667
R20095 VDAC_P.n1593 VDAC_P.n1592 0.180667
R20096 VDAC_P.n1594 VDAC_P.n1593 0.180667
R20097 VDAC_P.n1595 VDAC_P.n1594 0.180667
R20098 VDAC_P.n1596 VDAC_P.n1595 0.180667
R20099 VDAC_P.n1597 VDAC_P.n1596 0.180667
R20100 VDAC_P.n1598 VDAC_P.n1597 0.180667
R20101 VDAC_P.n1599 VDAC_P.n1598 0.180667
R20102 VDAC_P.n1600 VDAC_P.n1599 0.180667
R20103 VDAC_P.n1601 VDAC_P.n1600 0.180667
R20104 VDAC_P.n1602 VDAC_P.n1601 0.180667
R20105 VDAC_P.n1603 VDAC_P.n1602 0.180667
R20106 VDAC_P.n1604 VDAC_P.n1603 0.180667
R20107 VDAC_P.n1605 VDAC_P.n1604 0.180667
R20108 VDAC_P.n1606 VDAC_P.n1605 0.180667
R20109 VDAC_P.n1607 VDAC_P.n1606 0.180667
R20110 VDAC_P.n1608 VDAC_P.n1607 0.180667
R20111 VDAC_P.n1609 VDAC_P.n1608 0.180667
R20112 VDAC_P.n1610 VDAC_P.n1609 0.180667
R20113 VDAC_P.n1611 VDAC_P.n1610 0.180667
R20114 VDAC_P.n1612 VDAC_P.n1611 0.180667
R20115 VDAC_P.n1613 VDAC_P.n1612 0.180667
R20116 VDAC_P.n1614 VDAC_P.n1613 0.180667
R20117 VDAC_P.n1615 VDAC_P.n1614 0.180667
R20118 VDAC_P.n1616 VDAC_P.n1615 0.180667
R20119 VDAC_P.n1617 VDAC_P.n1616 0.180667
R20120 VDAC_P.n1618 VDAC_P.n1617 0.180667
R20121 VDAC_P.n1619 VDAC_P.n1618 0.180667
R20122 VDAC_P.n1620 VDAC_P.n1619 0.180667
R20123 VDAC_P.n1621 VDAC_P.n1620 0.180667
R20124 VDAC_P.n1622 VDAC_P.n1621 0.180667
R20125 VDAC_P.n1623 VDAC_P.n1622 0.180667
R20126 VDAC_P.n1624 VDAC_P.n1623 0.180667
R20127 VDAC_P.n1625 VDAC_P.n1624 0.180667
R20128 VDAC_P.n1626 VDAC_P.n1625 0.180667
R20129 VDAC_P.n1627 VDAC_P.n1626 0.180667
R20130 VDAC_P.n1628 VDAC_P.n1627 0.180667
R20131 VDAC_P.n1629 VDAC_P.n92 0.180667
R20132 VDAC_P.n1630 VDAC_P.n1629 0.180667
R20133 VDAC_P.n1631 VDAC_P.n1630 0.180667
R20134 VDAC_P.n1632 VDAC_P.n1631 0.180667
R20135 VDAC_P.n1633 VDAC_P.n1632 0.180667
R20136 VDAC_P.n1634 VDAC_P.n1633 0.180667
R20137 VDAC_P.n1635 VDAC_P.n1634 0.180667
R20138 VDAC_P.n1636 VDAC_P.n1635 0.180667
R20139 VDAC_P.n1637 VDAC_P.n1636 0.180667
R20140 VDAC_P.n1638 VDAC_P.n1637 0.180667
R20141 VDAC_P.n1639 VDAC_P.n1638 0.180667
R20142 VDAC_P.n1640 VDAC_P.n1639 0.180667
R20143 VDAC_P.n1641 VDAC_P.n1640 0.180667
R20144 VDAC_P.n1642 VDAC_P.n1641 0.180667
R20145 VDAC_P.n1643 VDAC_P.n1642 0.180667
R20146 VDAC_P.n1644 VDAC_P.n1643 0.180667
R20147 VDAC_P.n1645 VDAC_P.n1644 0.180667
R20148 VDAC_P.n1646 VDAC_P.n1645 0.180667
R20149 VDAC_P.n1647 VDAC_P.n1646 0.180667
R20150 VDAC_P.n1648 VDAC_P.n1647 0.180667
R20151 VDAC_P.n1649 VDAC_P.n1648 0.180667
R20152 VDAC_P.n1650 VDAC_P.n1649 0.180667
R20153 VDAC_P.n1651 VDAC_P.n1650 0.180667
R20154 VDAC_P.n1652 VDAC_P.n1651 0.180667
R20155 VDAC_P.n1653 VDAC_P.n1652 0.180667
R20156 VDAC_P.n1654 VDAC_P.n1653 0.180667
R20157 VDAC_P.n1655 VDAC_P.n1654 0.180667
R20158 VDAC_P.n1656 VDAC_P.n1655 0.180667
R20159 VDAC_P.n1657 VDAC_P.n1656 0.180667
R20160 VDAC_P.n1658 VDAC_P.n1657 0.180667
R20161 VDAC_P.n1659 VDAC_P.n1658 0.180667
R20162 VDAC_P.n1660 VDAC_P.n1659 0.180667
R20163 VDAC_P.n1661 VDAC_P.n1660 0.180667
R20164 VDAC_P.n1662 VDAC_P.n1661 0.180667
R20165 VDAC_P.n1663 VDAC_P.n1662 0.180667
R20166 VDAC_P.n1664 VDAC_P.n1663 0.180667
R20167 VDAC_P.n1665 VDAC_P.n1664 0.180667
R20168 VDAC_P.n1666 VDAC_P.n1665 0.180667
R20169 VDAC_P.n1667 VDAC_P.n1666 0.180667
R20170 VDAC_P.n1668 VDAC_P.n1667 0.180667
R20171 VDAC_P.n1669 VDAC_P.n1668 0.180667
R20172 VDAC_P.n1670 VDAC_P.n1669 0.180667
R20173 VDAC_P.n1671 VDAC_P.n1670 0.180667
R20174 VDAC_P.n1672 VDAC_P.n1671 0.180667
R20175 VDAC_P.n1673 VDAC_P.n1672 0.180667
R20176 VDAC_P.n1674 VDAC_P.n1673 0.180667
R20177 VDAC_P.n1675 VDAC_P.n1674 0.180667
R20178 VDAC_P.n1676 VDAC_P.n1675 0.180667
R20179 VDAC_P.n1677 VDAC_P.n1676 0.180667
R20180 VDAC_P.n1678 VDAC_P.n1677 0.180667
R20181 VDAC_P.n1679 VDAC_P.n1678 0.180667
R20182 VDAC_P.n1680 VDAC_P.n1679 0.180667
R20183 VDAC_P.n1681 VDAC_P.n1680 0.180667
R20184 VDAC_P.n1682 VDAC_P.n1681 0.180667
R20185 VDAC_P.n1683 VDAC_P.n1682 0.180667
R20186 VDAC_P.n1684 VDAC_P.n1683 0.180667
R20187 VDAC_P.n1685 VDAC_P.n1684 0.180667
R20188 VDAC_P.n1686 VDAC_P.n1685 0.180667
R20189 VDAC_P.n1687 VDAC_P.n1686 0.180667
R20190 VDAC_P.n1688 VDAC_P.n1687 0.180667
R20191 VDAC_P.n1689 VDAC_P.n1688 0.180667
R20192 VDAC_P.n1690 VDAC_P.n1689 0.180667
R20193 VDAC_P.n1691 VDAC_P.n1690 0.180667
R20194 VDAC_P.n1692 VDAC_P.n91 0.180667
R20195 VDAC_P.n1693 VDAC_P.n1692 0.180667
R20196 VDAC_P.n1694 VDAC_P.n1693 0.180667
R20197 VDAC_P.n1695 VDAC_P.n1694 0.180667
R20198 VDAC_P.n1696 VDAC_P.n1695 0.180667
R20199 VDAC_P.n1697 VDAC_P.n1696 0.180667
R20200 VDAC_P.n1698 VDAC_P.n1697 0.180667
R20201 VDAC_P.n1699 VDAC_P.n1698 0.180667
R20202 VDAC_P.n1700 VDAC_P.n1699 0.180667
R20203 VDAC_P.n1701 VDAC_P.n1700 0.180667
R20204 VDAC_P.n1702 VDAC_P.n1701 0.180667
R20205 VDAC_P.n1703 VDAC_P.n1702 0.180667
R20206 VDAC_P.n1704 VDAC_P.n1703 0.180667
R20207 VDAC_P.n1705 VDAC_P.n1704 0.180667
R20208 VDAC_P.n1706 VDAC_P.n1705 0.180667
R20209 VDAC_P.n1707 VDAC_P.n1706 0.180667
R20210 VDAC_P.n1708 VDAC_P.n1707 0.180667
R20211 VDAC_P.n1709 VDAC_P.n1708 0.180667
R20212 VDAC_P.n1710 VDAC_P.n1709 0.180667
R20213 VDAC_P.n1711 VDAC_P.n1710 0.180667
R20214 VDAC_P.n1712 VDAC_P.n1711 0.180667
R20215 VDAC_P.n1713 VDAC_P.n1712 0.180667
R20216 VDAC_P.n1714 VDAC_P.n1713 0.180667
R20217 VDAC_P.n1715 VDAC_P.n1714 0.180667
R20218 VDAC_P.n1716 VDAC_P.n1715 0.180667
R20219 VDAC_P.n1717 VDAC_P.n1716 0.180667
R20220 VDAC_P.n1718 VDAC_P.n1717 0.180667
R20221 VDAC_P.n1719 VDAC_P.n1718 0.180667
R20222 VDAC_P.n1720 VDAC_P.n1719 0.180667
R20223 VDAC_P.n1721 VDAC_P.n1720 0.180667
R20224 VDAC_P.n1722 VDAC_P.n1721 0.180667
R20225 VDAC_P.n1723 VDAC_P.n1722 0.180667
R20226 VDAC_P.n1724 VDAC_P.n1723 0.180667
R20227 VDAC_P.n1725 VDAC_P.n1724 0.180667
R20228 VDAC_P.n1726 VDAC_P.n1725 0.180667
R20229 VDAC_P.n1727 VDAC_P.n1726 0.180667
R20230 VDAC_P.n1728 VDAC_P.n1727 0.180667
R20231 VDAC_P.n1729 VDAC_P.n1728 0.180667
R20232 VDAC_P.n1730 VDAC_P.n1729 0.180667
R20233 VDAC_P.n1731 VDAC_P.n1730 0.180667
R20234 VDAC_P.n1732 VDAC_P.n1731 0.180667
R20235 VDAC_P.n1733 VDAC_P.n1732 0.180667
R20236 VDAC_P.n1734 VDAC_P.n1733 0.180667
R20237 VDAC_P.n1735 VDAC_P.n1734 0.180667
R20238 VDAC_P.n1736 VDAC_P.n1735 0.180667
R20239 VDAC_P.n1737 VDAC_P.n1736 0.180667
R20240 VDAC_P.n1738 VDAC_P.n1737 0.180667
R20241 VDAC_P.n1739 VDAC_P.n1738 0.180667
R20242 VDAC_P.n1740 VDAC_P.n1739 0.180667
R20243 VDAC_P.n1741 VDAC_P.n1740 0.180667
R20244 VDAC_P.n1742 VDAC_P.n1741 0.180667
R20245 VDAC_P.n1743 VDAC_P.n1742 0.180667
R20246 VDAC_P.n1744 VDAC_P.n1743 0.180667
R20247 VDAC_P.n1745 VDAC_P.n1744 0.180667
R20248 VDAC_P.n1746 VDAC_P.n1745 0.180667
R20249 VDAC_P.n1747 VDAC_P.n1746 0.180667
R20250 VDAC_P.n1748 VDAC_P.n1747 0.180667
R20251 VDAC_P.n1749 VDAC_P.n1748 0.180667
R20252 VDAC_P.n1750 VDAC_P.n1749 0.180667
R20253 VDAC_P.n1751 VDAC_P.n1750 0.180667
R20254 VDAC_P.n1752 VDAC_P.n1751 0.180667
R20255 VDAC_P.n1753 VDAC_P.n1752 0.180667
R20256 VDAC_P.n1754 VDAC_P.n1753 0.180667
R20257 VDAC_P.n1755 VDAC_P.n90 0.180667
R20258 VDAC_P.n1756 VDAC_P.n1755 0.180667
R20259 VDAC_P.n1757 VDAC_P.n1756 0.180667
R20260 VDAC_P.n1758 VDAC_P.n1757 0.180667
R20261 VDAC_P.n1759 VDAC_P.n1758 0.180667
R20262 VDAC_P.n1760 VDAC_P.n1759 0.180667
R20263 VDAC_P.n1761 VDAC_P.n1760 0.180667
R20264 VDAC_P.n1762 VDAC_P.n1761 0.180667
R20265 VDAC_P.n1763 VDAC_P.n1762 0.180667
R20266 VDAC_P.n1764 VDAC_P.n1763 0.180667
R20267 VDAC_P.n1765 VDAC_P.n1764 0.180667
R20268 VDAC_P.n1766 VDAC_P.n1765 0.180667
R20269 VDAC_P.n1767 VDAC_P.n1766 0.180667
R20270 VDAC_P.n1768 VDAC_P.n1767 0.180667
R20271 VDAC_P.n1769 VDAC_P.n1768 0.180667
R20272 VDAC_P.n1770 VDAC_P.n1769 0.180667
R20273 VDAC_P.n1771 VDAC_P.n1770 0.180667
R20274 VDAC_P.n1772 VDAC_P.n1771 0.180667
R20275 VDAC_P.n1773 VDAC_P.n1772 0.180667
R20276 VDAC_P.n1774 VDAC_P.n1773 0.180667
R20277 VDAC_P.n1775 VDAC_P.n1774 0.180667
R20278 VDAC_P.n1776 VDAC_P.n1775 0.180667
R20279 VDAC_P.n1777 VDAC_P.n1776 0.180667
R20280 VDAC_P.n1778 VDAC_P.n1777 0.180667
R20281 VDAC_P.n1779 VDAC_P.n1778 0.180667
R20282 VDAC_P.n1780 VDAC_P.n1779 0.180667
R20283 VDAC_P.n1781 VDAC_P.n1780 0.180667
R20284 VDAC_P.n1782 VDAC_P.n1781 0.180667
R20285 VDAC_P.n1783 VDAC_P.n1782 0.180667
R20286 VDAC_P.n1784 VDAC_P.n1783 0.180667
R20287 VDAC_P.n1785 VDAC_P.n1784 0.180667
R20288 VDAC_P.n1786 VDAC_P.n1785 0.180667
R20289 VDAC_P.n1787 VDAC_P.n1786 0.180667
R20290 VDAC_P.n1788 VDAC_P.n1787 0.180667
R20291 VDAC_P.n1789 VDAC_P.n1788 0.180667
R20292 VDAC_P.n1790 VDAC_P.n1789 0.180667
R20293 VDAC_P.n1791 VDAC_P.n1790 0.180667
R20294 VDAC_P.n1792 VDAC_P.n1791 0.180667
R20295 VDAC_P.n1793 VDAC_P.n1792 0.180667
R20296 VDAC_P.n1794 VDAC_P.n1793 0.180667
R20297 VDAC_P.n1795 VDAC_P.n1794 0.180667
R20298 VDAC_P.n1796 VDAC_P.n1795 0.180667
R20299 VDAC_P.n1797 VDAC_P.n1796 0.180667
R20300 VDAC_P.n1798 VDAC_P.n1797 0.180667
R20301 VDAC_P.n1799 VDAC_P.n1798 0.180667
R20302 VDAC_P.n1800 VDAC_P.n1799 0.180667
R20303 VDAC_P.n1801 VDAC_P.n1800 0.180667
R20304 VDAC_P.n1802 VDAC_P.n1801 0.180667
R20305 VDAC_P.n1803 VDAC_P.n1802 0.180667
R20306 VDAC_P.n1804 VDAC_P.n1803 0.180667
R20307 VDAC_P.n1805 VDAC_P.n1804 0.180667
R20308 VDAC_P.n1806 VDAC_P.n1805 0.180667
R20309 VDAC_P.n1807 VDAC_P.n1806 0.180667
R20310 VDAC_P.n1808 VDAC_P.n1807 0.180667
R20311 VDAC_P.n1809 VDAC_P.n1808 0.180667
R20312 VDAC_P.n1810 VDAC_P.n1809 0.180667
R20313 VDAC_P.n1811 VDAC_P.n1810 0.180667
R20314 VDAC_P.n1812 VDAC_P.n1811 0.180667
R20315 VDAC_P.n1813 VDAC_P.n1812 0.180667
R20316 VDAC_P.n1814 VDAC_P.n1813 0.180667
R20317 VDAC_P.n1815 VDAC_P.n1814 0.180667
R20318 VDAC_P.n1816 VDAC_P.n1815 0.180667
R20319 VDAC_P.n1817 VDAC_P.n1816 0.180667
R20320 VDAC_P.n1818 VDAC_P.n89 0.180667
R20321 VDAC_P.n1819 VDAC_P.n1818 0.180667
R20322 VDAC_P.n1820 VDAC_P.n1819 0.180667
R20323 VDAC_P.n1821 VDAC_P.n1820 0.180667
R20324 VDAC_P.n1822 VDAC_P.n1821 0.180667
R20325 VDAC_P.n1823 VDAC_P.n1822 0.180667
R20326 VDAC_P.n1824 VDAC_P.n1823 0.180667
R20327 VDAC_P.n1825 VDAC_P.n1824 0.180667
R20328 VDAC_P.n1826 VDAC_P.n1825 0.180667
R20329 VDAC_P.n1827 VDAC_P.n1826 0.180667
R20330 VDAC_P.n1828 VDAC_P.n1827 0.180667
R20331 VDAC_P.n1829 VDAC_P.n1828 0.180667
R20332 VDAC_P.n1830 VDAC_P.n1829 0.180667
R20333 VDAC_P.n1831 VDAC_P.n1830 0.180667
R20334 VDAC_P.n1832 VDAC_P.n1831 0.180667
R20335 VDAC_P.n1833 VDAC_P.n1832 0.180667
R20336 VDAC_P.n1834 VDAC_P.n1833 0.180667
R20337 VDAC_P.n1835 VDAC_P.n1834 0.180667
R20338 VDAC_P.n1836 VDAC_P.n1835 0.180667
R20339 VDAC_P.n1837 VDAC_P.n1836 0.180667
R20340 VDAC_P.n1838 VDAC_P.n1837 0.180667
R20341 VDAC_P.n1839 VDAC_P.n1838 0.180667
R20342 VDAC_P.n1840 VDAC_P.n1839 0.180667
R20343 VDAC_P.n1841 VDAC_P.n1840 0.180667
R20344 VDAC_P.n1842 VDAC_P.n1841 0.180667
R20345 VDAC_P.n1843 VDAC_P.n1842 0.180667
R20346 VDAC_P.n1844 VDAC_P.n1843 0.180667
R20347 VDAC_P.n1845 VDAC_P.n1844 0.180667
R20348 VDAC_P.n1846 VDAC_P.n1845 0.180667
R20349 VDAC_P.n1847 VDAC_P.n1846 0.180667
R20350 VDAC_P.n1848 VDAC_P.n1847 0.180667
R20351 VDAC_P.n1849 VDAC_P.n1848 0.180667
R20352 VDAC_P.n1850 VDAC_P.n1849 0.180667
R20353 VDAC_P.n1851 VDAC_P.n1850 0.180667
R20354 VDAC_P.n1852 VDAC_P.n1851 0.180667
R20355 VDAC_P.n1853 VDAC_P.n1852 0.180667
R20356 VDAC_P.n1854 VDAC_P.n1853 0.180667
R20357 VDAC_P.n1855 VDAC_P.n1854 0.180667
R20358 VDAC_P.n1856 VDAC_P.n1855 0.180667
R20359 VDAC_P.n1857 VDAC_P.n1856 0.180667
R20360 VDAC_P.n1858 VDAC_P.n1857 0.180667
R20361 VDAC_P.n1859 VDAC_P.n1858 0.180667
R20362 VDAC_P.n1860 VDAC_P.n1859 0.180667
R20363 VDAC_P.n1861 VDAC_P.n1860 0.180667
R20364 VDAC_P.n1862 VDAC_P.n1861 0.180667
R20365 VDAC_P.n1863 VDAC_P.n1862 0.180667
R20366 VDAC_P.n1864 VDAC_P.n1863 0.180667
R20367 VDAC_P.n1865 VDAC_P.n1864 0.180667
R20368 VDAC_P.n1866 VDAC_P.n1865 0.180667
R20369 VDAC_P.n1867 VDAC_P.n1866 0.180667
R20370 VDAC_P.n1868 VDAC_P.n1867 0.180667
R20371 VDAC_P.n1869 VDAC_P.n1868 0.180667
R20372 VDAC_P.n1870 VDAC_P.n1869 0.180667
R20373 VDAC_P.n1871 VDAC_P.n1870 0.180667
R20374 VDAC_P.n1872 VDAC_P.n1871 0.180667
R20375 VDAC_P.n1873 VDAC_P.n1872 0.180667
R20376 VDAC_P.n1874 VDAC_P.n1873 0.180667
R20377 VDAC_P.n1875 VDAC_P.n1874 0.180667
R20378 VDAC_P.n1876 VDAC_P.n1875 0.180667
R20379 VDAC_P.n1877 VDAC_P.n1876 0.180667
R20380 VDAC_P.n1878 VDAC_P.n1877 0.180667
R20381 VDAC_P.n1879 VDAC_P.n1878 0.180667
R20382 VDAC_P.n1880 VDAC_P.n1879 0.180667
R20383 VDAC_P.n1881 VDAC_P.n88 0.180667
R20384 VDAC_P.n1882 VDAC_P.n1881 0.180667
R20385 VDAC_P.n1883 VDAC_P.n1882 0.180667
R20386 VDAC_P.n1884 VDAC_P.n1883 0.180667
R20387 VDAC_P.n1885 VDAC_P.n1884 0.180667
R20388 VDAC_P.n1886 VDAC_P.n1885 0.180667
R20389 VDAC_P.n1887 VDAC_P.n1886 0.180667
R20390 VDAC_P.n1888 VDAC_P.n1887 0.180667
R20391 VDAC_P.n1889 VDAC_P.n1888 0.180667
R20392 VDAC_P.n1890 VDAC_P.n1889 0.180667
R20393 VDAC_P.n1891 VDAC_P.n1890 0.180667
R20394 VDAC_P.n1892 VDAC_P.n1891 0.180667
R20395 VDAC_P.n1893 VDAC_P.n1892 0.180667
R20396 VDAC_P.n1894 VDAC_P.n1893 0.180667
R20397 VDAC_P.n1895 VDAC_P.n1894 0.180667
R20398 VDAC_P.n1896 VDAC_P.n1895 0.180667
R20399 VDAC_P.n1897 VDAC_P.n1896 0.180667
R20400 VDAC_P.n1898 VDAC_P.n1897 0.180667
R20401 VDAC_P.n1899 VDAC_P.n1898 0.180667
R20402 VDAC_P.n1900 VDAC_P.n1899 0.180667
R20403 VDAC_P.n1901 VDAC_P.n1900 0.180667
R20404 VDAC_P.n1902 VDAC_P.n1901 0.180667
R20405 VDAC_P.n1903 VDAC_P.n1902 0.180667
R20406 VDAC_P.n1904 VDAC_P.n1903 0.180667
R20407 VDAC_P.n1905 VDAC_P.n1904 0.180667
R20408 VDAC_P.n1906 VDAC_P.n1905 0.180667
R20409 VDAC_P.n1907 VDAC_P.n1906 0.180667
R20410 VDAC_P.n1908 VDAC_P.n1907 0.180667
R20411 VDAC_P.n1909 VDAC_P.n1908 0.180667
R20412 VDAC_P.n1910 VDAC_P.n1909 0.180667
R20413 VDAC_P.n1911 VDAC_P.n1910 0.180667
R20414 VDAC_P.n1912 VDAC_P.n1911 0.180667
R20415 VDAC_P.n1913 VDAC_P.n1912 0.180667
R20416 VDAC_P.n1914 VDAC_P.n1913 0.180667
R20417 VDAC_P.n1915 VDAC_P.n1914 0.180667
R20418 VDAC_P.n1916 VDAC_P.n1915 0.180667
R20419 VDAC_P.n1917 VDAC_P.n1916 0.180667
R20420 VDAC_P.n1918 VDAC_P.n1917 0.180667
R20421 VDAC_P.n1919 VDAC_P.n1918 0.180667
R20422 VDAC_P.n1920 VDAC_P.n1919 0.180667
R20423 VDAC_P.n1921 VDAC_P.n1920 0.180667
R20424 VDAC_P.n1922 VDAC_P.n1921 0.180667
R20425 VDAC_P.n1923 VDAC_P.n1922 0.180667
R20426 VDAC_P.n1924 VDAC_P.n1923 0.180667
R20427 VDAC_P.n1925 VDAC_P.n1924 0.180667
R20428 VDAC_P.n1926 VDAC_P.n1925 0.180667
R20429 VDAC_P.n1927 VDAC_P.n1926 0.180667
R20430 VDAC_P.n1928 VDAC_P.n1927 0.180667
R20431 VDAC_P.n1929 VDAC_P.n1928 0.180667
R20432 VDAC_P.n1930 VDAC_P.n1929 0.180667
R20433 VDAC_P.n1931 VDAC_P.n1930 0.180667
R20434 VDAC_P.n1932 VDAC_P.n1931 0.180667
R20435 VDAC_P.n1933 VDAC_P.n1932 0.180667
R20436 VDAC_P.n1934 VDAC_P.n1933 0.180667
R20437 VDAC_P.n1935 VDAC_P.n1934 0.180667
R20438 VDAC_P.n1936 VDAC_P.n1935 0.180667
R20439 VDAC_P.n1937 VDAC_P.n1936 0.180667
R20440 VDAC_P.n1938 VDAC_P.n1937 0.180667
R20441 VDAC_P.n1939 VDAC_P.n1938 0.180667
R20442 VDAC_P.n1940 VDAC_P.n1939 0.180667
R20443 VDAC_P.n1941 VDAC_P.n1940 0.180667
R20444 VDAC_P.n1942 VDAC_P.n1941 0.180667
R20445 VDAC_P.n1943 VDAC_P.n1942 0.180667
R20446 VDAC_P.n87 VDAC_P.n86 0.180667
R20447 VDAC_P.n86 VDAC_P.n85 0.180667
R20448 VDAC_P.n85 VDAC_P.n84 0.180667
R20449 VDAC_P.n84 VDAC_P.n83 0.180667
R20450 VDAC_P.n83 VDAC_P.n82 0.180667
R20451 VDAC_P.n82 VDAC_P.n81 0.180667
R20452 VDAC_P.n81 VDAC_P.n80 0.180667
R20453 VDAC_P.n80 VDAC_P.n79 0.180667
R20454 VDAC_P.n79 VDAC_P.n78 0.180667
R20455 VDAC_P.n78 VDAC_P.n77 0.180667
R20456 VDAC_P.n77 VDAC_P.n76 0.180667
R20457 VDAC_P.n76 VDAC_P.n75 0.180667
R20458 VDAC_P.n75 VDAC_P.n74 0.180667
R20459 VDAC_P.n74 VDAC_P.n73 0.180667
R20460 VDAC_P.n73 VDAC_P.n72 0.180667
R20461 VDAC_P.n72 VDAC_P.n71 0.180667
R20462 VDAC_P.n71 VDAC_P.n70 0.180667
R20463 VDAC_P.n70 VDAC_P.n69 0.180667
R20464 VDAC_P.n69 VDAC_P.n68 0.180667
R20465 VDAC_P.n68 VDAC_P.n67 0.180667
R20466 VDAC_P.n67 VDAC_P.n66 0.180667
R20467 VDAC_P.n66 VDAC_P.n65 0.180667
R20468 VDAC_P.n65 VDAC_P.n64 0.180667
R20469 VDAC_P.n64 VDAC_P.n63 0.180667
R20470 VDAC_P.n63 VDAC_P.n62 0.180667
R20471 VDAC_P.n62 VDAC_P.n61 0.180667
R20472 VDAC_P.n61 VDAC_P.n60 0.180667
R20473 VDAC_P.n60 VDAC_P.n59 0.180667
R20474 VDAC_P.n59 VDAC_P.n58 0.180667
R20475 VDAC_P.n58 VDAC_P.n57 0.180667
R20476 VDAC_P.n57 VDAC_P.n56 0.180667
R20477 VDAC_P.n56 VDAC_P.n55 0.180667
R20478 VDAC_P.n55 VDAC_P.n54 0.180667
R20479 VDAC_P.n54 VDAC_P.n53 0.180667
R20480 VDAC_P.n53 VDAC_P.n52 0.180667
R20481 VDAC_P.n52 VDAC_P.n51 0.180667
R20482 VDAC_P.n51 VDAC_P.n50 0.180667
R20483 VDAC_P.n50 VDAC_P.n49 0.180667
R20484 VDAC_P.n49 VDAC_P.n48 0.180667
R20485 VDAC_P.n48 VDAC_P.n47 0.180667
R20486 VDAC_P.n47 VDAC_P.n46 0.180667
R20487 VDAC_P.n46 VDAC_P.n45 0.180667
R20488 VDAC_P.n45 VDAC_P.n44 0.180667
R20489 VDAC_P.n44 VDAC_P.n43 0.180667
R20490 VDAC_P.n43 VDAC_P.n42 0.180667
R20491 VDAC_P.n42 VDAC_P.n41 0.180667
R20492 VDAC_P.n41 VDAC_P.n40 0.180667
R20493 VDAC_P.n40 VDAC_P.n39 0.180667
R20494 VDAC_P.n39 VDAC_P.n38 0.180667
R20495 VDAC_P.n38 VDAC_P.n37 0.180667
R20496 VDAC_P.n37 VDAC_P.n36 0.180667
R20497 VDAC_P.n36 VDAC_P.n35 0.180667
R20498 VDAC_P.n35 VDAC_P.n34 0.180667
R20499 VDAC_P.n34 VDAC_P.n33 0.180667
R20500 VDAC_P.n33 VDAC_P.n32 0.180667
R20501 VDAC_P.n32 VDAC_P.n31 0.180667
R20502 VDAC_P.n31 VDAC_P.n30 0.180667
R20503 VDAC_P.n30 VDAC_P.n29 0.180667
R20504 VDAC_P.n29 VDAC_P.n28 0.180667
R20505 VDAC_P.n28 VDAC_P.n27 0.180667
R20506 VDAC_P.n27 VDAC_P.n26 0.180667
R20507 VDAC_P.n26 VDAC_P.n25 0.180667
R20508 VDAC_P.n25 VDAC_P.n24 0.180667
R20509 VDAC_P.n2134 VDAC_P.n23 0.180667
R20510 VDAC_P.n1973 VDAC_P.n1972 0.180667
R20511 VDAC_P.n1974 VDAC_P.n1973 0.180667
R20512 VDAC_P.n1975 VDAC_P.n1974 0.180667
R20513 VDAC_P.n1976 VDAC_P.n1975 0.180667
R20514 VDAC_P.n1977 VDAC_P.n1976 0.180667
R20515 VDAC_P.n1978 VDAC_P.n1977 0.180667
R20516 VDAC_P.n1979 VDAC_P.n1978 0.180667
R20517 VDAC_P.n1980 VDAC_P.n1979 0.180667
R20518 VDAC_P.n1981 VDAC_P.n1980 0.180667
R20519 VDAC_P.n1982 VDAC_P.n1981 0.180667
R20520 VDAC_P.n1983 VDAC_P.n1982 0.180667
R20521 VDAC_P.n1984 VDAC_P.n1983 0.180667
R20522 VDAC_P.n1985 VDAC_P.n1984 0.180667
R20523 VDAC_P.n1986 VDAC_P.n1985 0.180667
R20524 VDAC_P.n1987 VDAC_P.n1986 0.180667
R20525 VDAC_P.n1988 VDAC_P.n1987 0.180667
R20526 VDAC_P.n1989 VDAC_P.n1988 0.180667
R20527 VDAC_P.n1990 VDAC_P.n1989 0.180667
R20528 VDAC_P.n1991 VDAC_P.n1990 0.180667
R20529 VDAC_P.n1992 VDAC_P.n1991 0.180667
R20530 VDAC_P.n1993 VDAC_P.n1992 0.180667
R20531 VDAC_P.n1994 VDAC_P.n1993 0.180667
R20532 VDAC_P.n1995 VDAC_P.n1994 0.180667
R20533 VDAC_P.n1996 VDAC_P.n1995 0.180667
R20534 VDAC_P.n1997 VDAC_P.n1996 0.180667
R20535 VDAC_P.n1998 VDAC_P.n1997 0.180667
R20536 VDAC_P.n1999 VDAC_P.n1998 0.180667
R20537 VDAC_P.n2000 VDAC_P.n1999 0.180667
R20538 VDAC_P.n2001 VDAC_P.n2000 0.180667
R20539 VDAC_P.n2002 VDAC_P.n2001 0.180667
R20540 VDAC_P.n2003 VDAC_P.n2002 0.180667
R20541 VDAC_P.n2004 VDAC_P.n2003 0.180667
R20542 VDAC_P.n2005 VDAC_P.n2004 0.180667
R20543 VDAC_P.n2006 VDAC_P.n2005 0.180667
R20544 VDAC_P.n2007 VDAC_P.n2006 0.180667
R20545 VDAC_P.n2008 VDAC_P.n2007 0.180667
R20546 VDAC_P.n2009 VDAC_P.n2008 0.180667
R20547 VDAC_P.n2010 VDAC_P.n2009 0.180667
R20548 VDAC_P.n2011 VDAC_P.n2010 0.180667
R20549 VDAC_P.n2012 VDAC_P.n2011 0.180667
R20550 VDAC_P.n2013 VDAC_P.n2012 0.180667
R20551 VDAC_P.n2014 VDAC_P.n2013 0.180667
R20552 VDAC_P.n2015 VDAC_P.n2014 0.180667
R20553 VDAC_P.n2016 VDAC_P.n2015 0.180667
R20554 VDAC_P.n2017 VDAC_P.n2016 0.180667
R20555 VDAC_P.n2018 VDAC_P.n2017 0.180667
R20556 VDAC_P.n2019 VDAC_P.n2018 0.180667
R20557 VDAC_P.n2020 VDAC_P.n2019 0.180667
R20558 VDAC_P.n2021 VDAC_P.n2020 0.180667
R20559 VDAC_P.n2022 VDAC_P.n2021 0.180667
R20560 VDAC_P.n2023 VDAC_P.n2022 0.180667
R20561 VDAC_P.n2024 VDAC_P.n2023 0.180667
R20562 VDAC_P.n2025 VDAC_P.n2024 0.180667
R20563 VDAC_P.n2026 VDAC_P.n2025 0.180667
R20564 VDAC_P.n2027 VDAC_P.n2026 0.180667
R20565 VDAC_P.n2028 VDAC_P.n2027 0.180667
R20566 VDAC_P.n2029 VDAC_P.n2028 0.180667
R20567 VDAC_P.n2030 VDAC_P.n2029 0.180667
R20568 VDAC_P.n2031 VDAC_P.n2030 0.180667
R20569 VDAC_P.n2032 VDAC_P.n2031 0.180667
R20570 VDAC_P.n2033 VDAC_P.n2032 0.180667
R20571 VDAC_P.n2034 VDAC_P.n2033 0.180667
R20572 VDAC_P.n2035 VDAC_P.n2034 0.180667
R20573 VDAC_P.n2036 VDAC_P.n2035 0.180667
R20574 VDAC_P.n2037 VDAC_P.n2036 0.180667
R20575 VDAC_P.n2038 VDAC_P.n2037 0.180667
R20576 VDAC_P.n2039 VDAC_P.n2038 0.180667
R20577 VDAC_P.n2069 VDAC_P.n2068 0.180667
R20578 VDAC_P.n2070 VDAC_P.n2069 0.180667
R20579 VDAC_P.n2071 VDAC_P.n2070 0.180667
R20580 VDAC_P.n2072 VDAC_P.n2071 0.180667
R20581 VDAC_P.n2073 VDAC_P.n2072 0.180667
R20582 VDAC_P.n2074 VDAC_P.n2073 0.180667
R20583 VDAC_P.n2075 VDAC_P.n2074 0.180667
R20584 VDAC_P.n2076 VDAC_P.n2075 0.180667
R20585 VDAC_P.n2077 VDAC_P.n2076 0.180667
R20586 VDAC_P.n2078 VDAC_P.n2077 0.180667
R20587 VDAC_P.n2079 VDAC_P.n2078 0.180667
R20588 VDAC_P.n2080 VDAC_P.n2079 0.180667
R20589 VDAC_P.n2081 VDAC_P.n2080 0.180667
R20590 VDAC_P.n2082 VDAC_P.n2081 0.180667
R20591 VDAC_P.n2083 VDAC_P.n2082 0.180667
R20592 VDAC_P.n2084 VDAC_P.n2083 0.180667
R20593 VDAC_P.n2085 VDAC_P.n2084 0.180667
R20594 VDAC_P.n2086 VDAC_P.n2085 0.180667
R20595 VDAC_P.n2087 VDAC_P.n2086 0.180667
R20596 VDAC_P.n2088 VDAC_P.n2087 0.180667
R20597 VDAC_P.n2089 VDAC_P.n2088 0.180667
R20598 VDAC_P.n2090 VDAC_P.n2089 0.180667
R20599 VDAC_P.n2091 VDAC_P.n2090 0.180667
R20600 VDAC_P.n2092 VDAC_P.n2091 0.180667
R20601 VDAC_P.n2093 VDAC_P.n2092 0.180667
R20602 VDAC_P.n2094 VDAC_P.n2093 0.180667
R20603 VDAC_P.n2095 VDAC_P.n2094 0.180667
R20604 VDAC_P.n2096 VDAC_P.n2095 0.180667
R20605 VDAC_P.n2097 VDAC_P.n2096 0.180667
R20606 VDAC_P.n2098 VDAC_P.n2097 0.180667
R20607 VDAC_P.n2099 VDAC_P.n2098 0.180667
R20608 VDAC_P.n2100 VDAC_P.n2099 0.180667
R20609 VDAC_P.n2101 VDAC_P.n2100 0.180667
R20610 VDAC_P.n2102 VDAC_P.n2101 0.180667
R20611 VDAC_P.n2103 VDAC_P.n2102 0.180667
R20612 VDAC_P.n2104 VDAC_P.n2103 0.180667
R20613 VDAC_P.n2105 VDAC_P.n2104 0.180667
R20614 VDAC_P.n2106 VDAC_P.n2105 0.180667
R20615 VDAC_P.n2107 VDAC_P.n2106 0.180667
R20616 VDAC_P.n2108 VDAC_P.n2107 0.180667
R20617 VDAC_P.n2109 VDAC_P.n2108 0.180667
R20618 VDAC_P.n2110 VDAC_P.n2109 0.180667
R20619 VDAC_P.n2111 VDAC_P.n2110 0.180667
R20620 VDAC_P.n2112 VDAC_P.n2111 0.180667
R20621 VDAC_P.n2113 VDAC_P.n2112 0.180667
R20622 VDAC_P.n2114 VDAC_P.n2113 0.180667
R20623 VDAC_P.n2115 VDAC_P.n2114 0.180667
R20624 VDAC_P.n2116 VDAC_P.n2115 0.180667
R20625 VDAC_P.n2117 VDAC_P.n2116 0.180667
R20626 VDAC_P.n2118 VDAC_P.n2117 0.180667
R20627 VDAC_P.n2119 VDAC_P.n2118 0.180667
R20628 VDAC_P.n2120 VDAC_P.n2119 0.180667
R20629 VDAC_P.n2121 VDAC_P.n2120 0.180667
R20630 VDAC_P.n2122 VDAC_P.n2121 0.180667
R20631 VDAC_P.n2123 VDAC_P.n2122 0.180667
R20632 VDAC_P.n2124 VDAC_P.n2123 0.180667
R20633 VDAC_P.n2125 VDAC_P.n2124 0.180667
R20634 VDAC_P.n2126 VDAC_P.n2125 0.180667
R20635 VDAC_P.n2127 VDAC_P.n2126 0.180667
R20636 VDAC_P.n2128 VDAC_P.n2127 0.180667
R20637 VDAC_P.n2129 VDAC_P.n2128 0.180667
R20638 VDAC_P.n2130 VDAC_P.n2129 0.180667
R20639 VDAC_P.n2131 VDAC_P.n2130 0.180667
R20640 VDAC_P.n2132 VDAC_P.n2131 0.180667
R20641 VDAC_P.n2133 VDAC_P.n2132 0.180667
R20642 VDAC_P.n2134 VDAC_P.n2133 0.180667
R20643 VDAC_P.n2039 VDAC_P.n116 0.157167
R20644 VDAC_P.n1972 VDAC_P.n179 0.157167
R20645 VDAC_P.n2040 VDAC_P.n115 0.157167
R20646 VDAC_P.n1971 VDAC_P.n242 0.157167
R20647 VDAC_P.n2041 VDAC_P.n114 0.157167
R20648 VDAC_P.n1970 VDAC_P.n305 0.157167
R20649 VDAC_P.n2042 VDAC_P.n113 0.157167
R20650 VDAC_P.n1969 VDAC_P.n368 0.157167
R20651 VDAC_P.n2043 VDAC_P.n112 0.157167
R20652 VDAC_P.n1968 VDAC_P.n431 0.157167
R20653 VDAC_P.n2044 VDAC_P.n111 0.157167
R20654 VDAC_P.n1967 VDAC_P.n494 0.157167
R20655 VDAC_P.n2045 VDAC_P.n110 0.157167
R20656 VDAC_P.n1966 VDAC_P.n557 0.157167
R20657 VDAC_P.n2046 VDAC_P.n109 0.157167
R20658 VDAC_P.n1965 VDAC_P.n620 0.157167
R20659 VDAC_P.n2047 VDAC_P.n108 0.157167
R20660 VDAC_P.n1964 VDAC_P.n683 0.157167
R20661 VDAC_P.n2048 VDAC_P.n107 0.157167
R20662 VDAC_P.n1963 VDAC_P.n746 0.157167
R20663 VDAC_P.n2049 VDAC_P.n106 0.157167
R20664 VDAC_P.n1962 VDAC_P.n809 0.157167
R20665 VDAC_P.n2050 VDAC_P.n105 0.157167
R20666 VDAC_P.n1961 VDAC_P.n872 0.157167
R20667 VDAC_P.n2051 VDAC_P.n104 0.157167
R20668 VDAC_P.n1960 VDAC_P.n935 0.157167
R20669 VDAC_P.n2052 VDAC_P.n103 0.157167
R20670 VDAC_P.n1959 VDAC_P.n998 0.157167
R20671 VDAC_P.n2053 VDAC_P.n102 0.157167
R20672 VDAC_P.n1958 VDAC_P.n1061 0.157167
R20673 VDAC_P.n2054 VDAC_P.n101 0.157167
R20674 VDAC_P.n1957 VDAC_P.n1124 0.157167
R20675 VDAC_P.n2055 VDAC_P.n100 0.157167
R20676 VDAC_P.n1956 VDAC_P.n1187 0.157167
R20677 VDAC_P.n2056 VDAC_P.n99 0.157167
R20678 VDAC_P.n1955 VDAC_P.n1250 0.157167
R20679 VDAC_P.n2057 VDAC_P.n98 0.157167
R20680 VDAC_P.n1954 VDAC_P.n1313 0.157167
R20681 VDAC_P.n2058 VDAC_P.n97 0.157167
R20682 VDAC_P.n1953 VDAC_P.n1376 0.157167
R20683 VDAC_P.n2059 VDAC_P.n96 0.157167
R20684 VDAC_P.n1952 VDAC_P.n1439 0.157167
R20685 VDAC_P.n2060 VDAC_P.n95 0.157167
R20686 VDAC_P.n1951 VDAC_P.n1502 0.157167
R20687 VDAC_P.n2061 VDAC_P.n94 0.157167
R20688 VDAC_P.n1950 VDAC_P.n1565 0.157167
R20689 VDAC_P.n2062 VDAC_P.n93 0.157167
R20690 VDAC_P.n1949 VDAC_P.n1628 0.157167
R20691 VDAC_P.n2063 VDAC_P.n92 0.157167
R20692 VDAC_P.n1948 VDAC_P.n1691 0.157167
R20693 VDAC_P.n2064 VDAC_P.n91 0.157167
R20694 VDAC_P.n1947 VDAC_P.n1754 0.157167
R20695 VDAC_P.n2065 VDAC_P.n90 0.157167
R20696 VDAC_P.n1946 VDAC_P.n1817 0.157167
R20697 VDAC_P.n2066 VDAC_P.n89 0.157167
R20698 VDAC_P.n1945 VDAC_P.n1880 0.157167
R20699 VDAC_P.n2067 VDAC_P.n88 0.157167
R20700 VDAC_P.n1944 VDAC_P.n1943 0.157167
R20701 VDAC_P.n2068 VDAC_P.n87 0.157167
R20702 VDAC_P.n24 VDAC_P.n23 0.157167
R20703 VDAC_P VDAC_P.n2134 0.071
R20704 a_5088_37509.n16 a_5088_37509.t1 120.862
R20705 a_5088_37509.n15 a_5088_37509.t3 120.564
R20706 a_5088_37509.n17 a_5088_37509.n16 104.312
R20707 a_5088_37509.n2 a_5088_37509.n0 40.84
R20708 a_5088_37509.n6 a_5088_37509.n5 40.5431
R20709 a_5088_37509.n4 a_5088_37509.n3 40.5431
R20710 a_5088_37509.n2 a_5088_37509.n1 40.5431
R20711 a_5088_37509.n9 a_5088_37509.n7 40.4813
R20712 a_5088_37509.n13 a_5088_37509.n12 40.1844
R20713 a_5088_37509.n11 a_5088_37509.n10 40.1844
R20714 a_5088_37509.n9 a_5088_37509.n8 40.1844
R20715 a_5088_37509.n15 a_5088_37509.n14 24.9745
R20716 a_5088_37509.n17 a_5088_37509.t2 16.253
R20717 a_5088_37509.t0 a_5088_37509.n17 16.253
R20718 a_5088_37509.n14 a_5088_37509.n13 13.188
R20719 a_5088_37509.n12 a_5088_37509.t14 4.76133
R20720 a_5088_37509.n12 a_5088_37509.t6 4.76133
R20721 a_5088_37509.n10 a_5088_37509.t13 4.76133
R20722 a_5088_37509.n10 a_5088_37509.t5 4.76133
R20723 a_5088_37509.n8 a_5088_37509.t9 4.76133
R20724 a_5088_37509.n8 a_5088_37509.t15 4.76133
R20725 a_5088_37509.n7 a_5088_37509.t11 4.76133
R20726 a_5088_37509.n7 a_5088_37509.t19 4.76133
R20727 a_5088_37509.n5 a_5088_37509.t17 4.76133
R20728 a_5088_37509.n5 a_5088_37509.t7 4.76133
R20729 a_5088_37509.n3 a_5088_37509.t18 4.76133
R20730 a_5088_37509.n3 a_5088_37509.t12 4.76133
R20731 a_5088_37509.n1 a_5088_37509.t8 4.76133
R20732 a_5088_37509.n1 a_5088_37509.t4 4.76133
R20733 a_5088_37509.n0 a_5088_37509.t16 4.76133
R20734 a_5088_37509.n0 a_5088_37509.t10 4.76133
R20735 a_5088_37509.n11 a_5088_37509.n9 0.313
R20736 a_5088_37509.n13 a_5088_37509.n11 0.313
R20737 a_5088_37509.n4 a_5088_37509.n2 0.313
R20738 a_5088_37509.n6 a_5088_37509.n4 0.313
R20739 a_5088_37509.n14 a_5088_37509.n6 0.297375
R20740 a_5088_37509.n16 a_5088_37509.n15 0.297375
R20741 a_8912_37509.n1 a_8912_37509.t25 45.8845
R20742 a_8912_37509.n30 a_8912_37509.t16 45.6616
R20743 a_8912_37509.n6 a_8912_37509.t34 45.6572
R20744 a_8912_37509.n7 a_8912_37509.t7 45.6572
R20745 a_8912_37509.n14 a_8912_37509.t11 45.6572
R20746 a_8912_37509.n35 a_8912_37509.t8 45.4344
R20747 a_8912_37509.n36 a_8912_37509.t24 45.4344
R20748 a_8912_37509.n43 a_8912_37509.t29 45.4344
R20749 a_8912_37509.n1 a_8912_37509.n0 40.8964
R20750 a_8912_37509.n3 a_8912_37509.n2 40.8964
R20751 a_8912_37509.n5 a_8912_37509.n4 40.8964
R20752 a_8912_37509.n9 a_8912_37509.n8 40.8964
R20753 a_8912_37509.n11 a_8912_37509.n10 40.8964
R20754 a_8912_37509.n13 a_8912_37509.n12 40.8964
R20755 a_8912_37509.n30 a_8912_37509.n29 40.6735
R20756 a_8912_37509.n32 a_8912_37509.n31 40.6735
R20757 a_8912_37509.n34 a_8912_37509.n33 40.6735
R20758 a_8912_37509.n38 a_8912_37509.n37 40.6735
R20759 a_8912_37509.n40 a_8912_37509.n39 40.6735
R20760 a_8912_37509.n42 a_8912_37509.n41 40.6735
R20761 a_8912_37509.n27 a_8912_37509.t4 30.0869
R20762 a_8912_37509.n24 a_8912_37509.t2 30.0869
R20763 a_8912_37509.n22 a_8912_37509.t3 30.0869
R20764 a_8912_37509.n19 a_8912_37509.t5 30.0869
R20765 a_8912_37509.n18 a_8912_37509.t1 30.0869
R20766 a_8912_37509.t0 a_8912_37509.n45 30.0869
R20767 a_8912_37509.n18 a_8912_37509.n17 5.95542
R20768 a_8912_37509.n27 a_8912_37509.n26 5.6486
R20769 a_8912_37509.n25 a_8912_37509.n24 5.6486
R20770 a_8912_37509.n23 a_8912_37509.n22 5.6486
R20771 a_8912_37509.n19 a_8912_37509.n17 5.6486
R20772 a_8912_37509.n45 a_8912_37509.n15 5.6486
R20773 a_8912_37509.n20 a_8912_37509.n18 4.80732
R20774 a_8912_37509.n29 a_8912_37509.t6 4.76133
R20775 a_8912_37509.n29 a_8912_37509.t14 4.76133
R20776 a_8912_37509.n31 a_8912_37509.t13 4.76133
R20777 a_8912_37509.n31 a_8912_37509.t20 4.76133
R20778 a_8912_37509.n33 a_8912_37509.t21 4.76133
R20779 a_8912_37509.n33 a_8912_37509.t12 4.76133
R20780 a_8912_37509.n37 a_8912_37509.t23 4.76133
R20781 a_8912_37509.n37 a_8912_37509.t32 4.76133
R20782 a_8912_37509.n39 a_8912_37509.t33 4.76133
R20783 a_8912_37509.n39 a_8912_37509.t31 4.76133
R20784 a_8912_37509.n41 a_8912_37509.t37 4.76133
R20785 a_8912_37509.n41 a_8912_37509.t27 4.76133
R20786 a_8912_37509.n0 a_8912_37509.t30 4.76133
R20787 a_8912_37509.n0 a_8912_37509.t35 4.76133
R20788 a_8912_37509.n2 a_8912_37509.t22 4.76133
R20789 a_8912_37509.n2 a_8912_37509.t36 4.76133
R20790 a_8912_37509.n4 a_8912_37509.t28 4.76133
R20791 a_8912_37509.n4 a_8912_37509.t26 4.76133
R20792 a_8912_37509.n8 a_8912_37509.t19 4.76133
R20793 a_8912_37509.n8 a_8912_37509.t15 4.76133
R20794 a_8912_37509.n10 a_8912_37509.t18 4.76133
R20795 a_8912_37509.n10 a_8912_37509.t10 4.76133
R20796 a_8912_37509.n12 a_8912_37509.t17 4.76133
R20797 a_8912_37509.n12 a_8912_37509.t9 4.76133
R20798 a_8912_37509.n20 a_8912_37509.n19 4.5005
R20799 a_8912_37509.n22 a_8912_37509.n21 4.5005
R20800 a_8912_37509.n24 a_8912_37509.n16 4.5005
R20801 a_8912_37509.n28 a_8912_37509.n27 4.5005
R20802 a_8912_37509.n45 a_8912_37509.n44 4.5005
R20803 a_8912_37509.n15 a_8912_37509.n14 1.19141
R20804 a_8912_37509.n44 a_8912_37509.n43 1.18686
R20805 a_8912_37509.n21 a_8912_37509.n16 0.614136
R20806 a_8912_37509.n25 a_8912_37509.n23 0.614136
R20807 a_8912_37509.n28 a_8912_37509.n16 0.318682
R20808 a_8912_37509.n26 a_8912_37509.n25 0.318682
R20809 a_8912_37509.n21 a_8912_37509.n20 0.307318
R20810 a_8912_37509.n44 a_8912_37509.n28 0.307318
R20811 a_8912_37509.n23 a_8912_37509.n17 0.307318
R20812 a_8912_37509.n26 a_8912_37509.n15 0.307318
R20813 a_8912_37509.n36 a_8912_37509.n35 0.261864
R20814 a_8912_37509.n7 a_8912_37509.n6 0.261864
R20815 a_8912_37509.n42 a_8912_37509.n40 0.227773
R20816 a_8912_37509.n40 a_8912_37509.n38 0.227773
R20817 a_8912_37509.n35 a_8912_37509.n34 0.227773
R20818 a_8912_37509.n34 a_8912_37509.n32 0.227773
R20819 a_8912_37509.n14 a_8912_37509.n13 0.227773
R20820 a_8912_37509.n11 a_8912_37509.n9 0.227773
R20821 a_8912_37509.n6 a_8912_37509.n5 0.227773
R20822 a_8912_37509.n5 a_8912_37509.n3 0.227773
R20823 a_8912_37509.n43 a_8912_37509.n42 0.216409
R20824 a_8912_37509.n38 a_8912_37509.n36 0.216409
R20825 a_8912_37509.n32 a_8912_37509.n30 0.216409
R20826 a_8912_37509.n13 a_8912_37509.n11 0.216409
R20827 a_8912_37509.n9 a_8912_37509.n7 0.216409
R20828 a_8912_37509.n3 a_8912_37509.n1 0.216409
R20829 VDD.n219 VDD.t2917 187509
R20830 VDD.n321 VDD.n219 135375
R20831 VDD.n321 VDD.t2253 115781
R20832 VDD.n147 VDD.n107 15352.9
R20833 VDD.n147 VDD.n108 15352.9
R20834 VDD.n146 VDD.n134 15352.9
R20835 VDD.n146 VDD.n137 15352.9
R20836 VDD.n75 VDD.n67 13260
R20837 VDD.n72 VDD.n68 13260
R20838 VDD.n38 VDD.n31 13260
R20839 VDD.n35 VDD.n32 13260
R20840 VDD.n72 VDD.n67 13154.1
R20841 VDD.n75 VDD.n68 13154.1
R20842 VDD.n35 VDD.n31 13154.1
R20843 VDD.n38 VDD.n32 13154.1
R20844 VDD.n110 VDD.n109 11297.6
R20845 VDD.n135 VDD.n109 11297.6
R20846 VDD.n320 VDD.n319 9790.59
R20847 VDD.n319 VDD.n221 8022.35
R20848 VDD.n215 VDD.n192 6963.53
R20849 VDD.n215 VDD.n194 6963.53
R20850 VDD.n320 VDD.n185 6374.12
R20851 VDD.n226 VDD.n186 5516.47
R20852 VDD.n140 VDD.n105 5440
R20853 VDD.n210 VDD.n186 5379.02
R20854 VDD.n191 VDD.n189 5177.65
R20855 VDD.n209 VDD.n189 5177.65
R20856 VDD.n134 VDD.n110 4055.29
R20857 VDD.n137 VDD.n135 4055.29
R20858 VDD.n135 VDD.n108 4055.29
R20859 VDD.n323 VDD.n185 3220
R20860 VDD.n323 VDD.n186 3220
R20861 VDD.n127 VDD.n126 2771.2
R20862 VDD.n128 VDD.n127 2662.4
R20863 VDD.n259 VDD.n256 2311.76
R20864 VDD.n261 VDD.n256 2311.76
R20865 VDD.n267 VDD.n253 2311.76
R20866 VDD.n265 VDD.n253 2311.76
R20867 VDD.n2456 VDD.n2406 2296.22
R20868 VDD.n229 VDD.n228 2068.24
R20869 VDD.n228 VDD.n227 2068.24
R20870 VDD.n4139 VDD.n3720 2060.8
R20871 VDD.n4269 VDD.n4266 2060.8
R20872 VDD.n344 VDD.n336 1937.65
R20873 VDD.n345 VDD.n344 1937.65
R20874 VDD.n191 VDD.n188 1785.88
R20875 VDD.n192 VDD.n191 1785.88
R20876 VDD.n210 VDD.n209 1785.88
R20877 VDD.n209 VDD.n194 1785.88
R20878 VDD.n221 VDD.n220 1768.24
R20879 VDD.n347 VDD.n343 1757.65
R20880 VDD.n389 VDD.n340 1757.65
R20881 VDD.n364 VDD.n347 1757.65
R20882 VDD.n124 VDD.n112 1754.12
R20883 VDD.n130 VDD.n113 1754.12
R20884 VDD.n389 VDD.n337 1750.59
R20885 VDD.n188 VDD.n185 1718.82
R20886 VDD.t2274 VDD.t2526 1698.59
R20887 VDD.n4139 VDD.n4138 1612.8
R20888 VDD.n4270 VDD.n4269 1612.8
R20889 VDD.n376 VDD.n374 1436.47
R20890 VDD.n384 VDD.n378 1436.47
R20891 VDD.n2457 VDD.n2456 1411.01
R20892 VDD.n116 VDD.n115 1348.24
R20893 VDD.n115 VDD.n114 1348.24
R20894 VDD.n202 VDD.n197 1312.94
R20895 VDD.n200 VDD.n197 1312.94
R20896 VDD.n200 VDD.n198 1312.94
R20897 VDD.t2333 VDD.t2283 1235.34
R20898 VDD.t2566 VDD.t2363 1235.34
R20899 VDD.n257 VDD.n252 1231.76
R20900 VDD.n257 VDD.n254 1231.76
R20901 VDD.n141 VDD.n140 1195.67
R20902 VDD.n142 VDD.n141 1187.39
R20903 VDD.n128 VDD.n119 1113.6
R20904 VDD.t137 VDD.t2506 1099.38
R20905 VDD.t2283 VDD.t113 1084.28
R20906 VDD.n259 VDD.n252 1080
R20907 VDD.n267 VDD.n252 1080
R20908 VDD.n261 VDD.n254 1080
R20909 VDD.n265 VDD.n254 1080
R20910 VDD.n114 VDD.n112 1080
R20911 VDD.n130 VDD.n116 1080
R20912 VDD.n122 VDD.n111 1080
R20913 VDD.n115 VDD.n111 1080
R20914 VDD.n412 VDD.t1718 1001.47
R20915 VDD.t587 VDD.t2277 929.86
R20916 VDD.t2628 VDD.t264 929.86
R20917 VDD.t2487 VDD.t2443 926.503
R20918 VDD.n425 VDD.t1728 879.831
R20919 VDD.n384 VDD.n377 878.823
R20920 VDD.n352 VDD.n351 878.823
R20921 VDD.n353 VDD.n352 878.823
R20922 VDD.n50 VDD.t2763 877.016
R20923 VDD.n12 VDD.t2721 877.016
R20924 VDD.n2714 VDD.t159 873.438
R20925 VDD.n2634 VDD.t2950 873.438
R20926 VDD.n2620 VDD.t1746 873.438
R20927 VDD.n1876 VDD.t514 873.438
R20928 VDD.n1877 VDD.t2668 872.107
R20929 VDD.n55 VDD.t3053 871.962
R20930 VDD.n15 VDD.t3057 871.962
R20931 VDD.n377 VDD.n376 871.765
R20932 VDD.n2359 VDD.t1838 871.529
R20933 VDD.n2383 VDD.t1712 871.529
R20934 VDD.n2626 VDD.t914 870.754
R20935 VDD.n1364 VDD.t1592 870.754
R20936 VDD.n1879 VDD.t2666 870.754
R20937 VDD.n2720 VDD.t660 870.024
R20938 VDD.n2640 VDD.t747 870.024
R20939 VDD.n2715 VDD.t658 869.086
R20940 VDD.n2635 VDD.t749 869.086
R20941 VDD.n2621 VDD.t916 869.086
R20942 VDD.n2391 VDD.t2705 869.086
R20943 VDD.n2514 VDD.t1976 869.086
R20944 VDD.n1378 VDD.t1594 869.086
R20945 VDD.n1362 VDD.t757 869.086
R20946 VDD.n1406 VDD.t1630 869.086
R20947 VDD.n2049 VDD.t1737 869.086
R20948 VDD.n2009 VDD.t1993 869.086
R20949 VDD.n2006 VDD.t1393 869.086
R20950 VDD.n1745 VDD.t1203 869.086
R20951 VDD.n1745 VDD.t3101 869.086
R20952 VDD.n3290 VDD.t1219 868.721
R20953 VDD.n2995 VDD.t1852 868.721
R20954 VDD.n2389 VDD.t1978 867.003
R20955 VDD.n1404 VDD.t1739 867.003
R20956 VDD.n2014 VDD.t1991 867.003
R20957 VDD.n1750 VDD.t1201 867.003
R20958 VDD.n71 VDD.n69 861.352
R20959 VDD.n34 VDD.n29 861.268
R20960 VDD.n226 VDD.n220 857.648
R20961 VDD.n71 VDD.n70 857.359
R20962 VDD.n34 VDD.n33 857.183
R20963 VDD.n3134 VDD.t2622 849.293
R20964 VDD.t2643 VDD.t2601 849.293
R20965 VDD.n149 VDD.n105 845.83
R20966 VDD.n3227 VDD.t1435 838.817
R20967 VDD.n4094 VDD.t1377 836.124
R20968 VDD.n4343 VDD.t1087 836.124
R20969 VDD.n3953 VDD.t1113 836.124
R20970 VDD.n2966 VDD.t1464 836.124
R20971 VDD.n2987 VDD.t2156 836.124
R20972 VDD.n2380 VDD.t1290 836.124
R20973 VDD.n4244 VDD.t2111 832.876
R20974 VDD.n4131 VDD.t1188 832.876
R20975 VDD.n3908 VDD.t1035 832.876
R20976 VDD.n1894 VDD.t2182 832.876
R20977 VDD.n3107 VDD.t2528 812.141
R20978 VDD.n3105 VDD.t2275 811.918
R20979 VDD.n3039 VDD.t2624 809.322
R20980 VDD.n1584 VDD.t2507 809.232
R20981 VDD.n2396 VDD.t2270 807.567
R20982 VDD.n1574 VDD.t2399 807.548
R20983 VDD.n2500 VDD.t2588 807.481
R20984 VDD.n2917 VDD.t3090 806.511
R20985 VDD.n3481 VDD.t2107 806.511
R20986 VDD.n3392 VDD.t1229 806.511
R20987 VDD.n2976 VDD.t1490 806.511
R20988 VDD.n3320 VDD.t2119 806.511
R20989 VDD.n3545 VDD.t623 806.511
R20990 VDD.n3540 VDD.t1259 806.511
R20991 VDD.n3166 VDD.t1425 806.511
R20992 VDD.n3174 VDD.t627 806.511
R20993 VDD.n2238 VDD.t1915 806.511
R20994 VDD.n1971 VDD.t857 806.511
R20995 VDD.n1709 VDD.t921 806.511
R20996 VDD.n1563 VDD.t1888 806.511
R20997 VDD.n1543 VDD.t1417 806.511
R20998 VDD.n1072 VDD.t2113 806.511
R20999 VDD.n2838 VDD.t2466 805.957
R21000 VDD.n3693 VDD.t2583 804.731
R21001 VDD.n4182 VDD.t2407 804.731
R21002 VDD.n4240 VDD.t2632 804.731
R21003 VDD.n3712 VDD.t2469 804.731
R21004 VDD.n3721 VDD.t2468 804.731
R21005 VDD.n3739 VDD.t2433 804.731
R21006 VDD.t2488 VDD.n3876 804.731
R21007 VDD.n3879 VDD.t2444 804.731
R21008 VDD.n3900 VDD.t2445 804.731
R21009 VDD.n3821 VDD.t2462 804.731
R21010 VDD.n3907 VDD.t2463 804.731
R21011 VDD.n3830 VDD.t2448 804.731
R21012 VDD.n3850 VDD.t2289 804.731
R21013 VDD.n3853 VDD.t2513 804.731
R21014 VDD.n4376 VDD.t2442 804.731
R21015 VDD.n4368 VDD.t2441 804.731
R21016 VDD.n3670 VDD.t2618 804.731
R21017 VDD.n4323 VDD.t2617 804.731
R21018 VDD.n3679 VDD.t2436 804.731
R21019 VDD.n4289 VDD.t2516 804.731
R21020 VDD.n3685 VDD.t2435 804.731
R21021 VDD.n4272 VDD.t2515 804.731
R21022 VDD.n3675 VDD.t2347 804.731
R21023 VDD.n4063 VDD.t2380 804.731
R21024 VDD.n4045 VDD.t2457 804.731
R21025 VDD.n4025 VDD.t2456 804.731
R21026 VDD.n3792 VDD.t2426 804.731
R21027 VDD.n3799 VDD.t2504 804.731
R21028 VDD.n3942 VDD.t2627 804.731
R21029 VDD.n3920 VDD.t2626 804.731
R21030 VDD.t2361 VDD.n3917 804.731
R21031 VDD.n4392 VDD.t2499 804.731
R21032 VDD.n4395 VDD.t2344 804.731
R21033 VDD.n2924 VDD.t2497 804.731
R21034 VDD.n3589 VDD.t2560 804.731
R21035 VDD.n3583 VDD.t2559 804.731
R21036 VDD.n3589 VDD.t2285 804.731
R21037 VDD.n3583 VDD.t2284 804.731
R21038 VDD.n3079 VDD.t2623 804.731
R21039 VDD.n3087 VDD.t2276 804.731
R21040 VDD.n3125 VDD.t2527 804.731
R21041 VDD.n3077 VDD.t2630 804.731
R21042 VDD.n3071 VDD.t2629 804.731
R21043 VDD.n3050 VDD.t2413 804.731
R21044 VDD.n3053 VDD.t2322 804.731
R21045 VDD.n3042 VDD.t2405 804.731
R21046 VDD.n3070 VDD.t2586 804.731
R21047 VDD.n3579 VDD.t2335 804.731
R21048 VDD.n3582 VDD.t2454 804.731
R21049 VDD.n3601 VDD.t2301 804.731
R21050 VDD.n3604 VDD.t2421 804.731
R21051 VDD.n2520 VDD.t2589 804.731
R21052 VDD.n2375 VDD.t2591 804.731
R21053 VDD.t2592 VDD.n2370 804.731
R21054 VDD.n2557 VDD.t2410 804.731
R21055 VDD.t2389 VDD.n2596 804.731
R21056 VDD.n2339 VDD.t2477 804.731
R21057 VDD.n2329 VDD.t2478 804.731
R21058 VDD.t2614 VDD.n2643 804.731
R21059 VDD.n2647 VDD.t2615 804.731
R21060 VDD.n2680 VDD.t2460 804.731
R21061 VDD.n2660 VDD.t2459 804.731
R21062 VDD.n2824 VDD.t2465 804.731
R21063 VDD.n2840 VDD.t2602 804.731
R21064 VDD.n2099 VDD.t2598 804.731
R21065 VDD.n2177 VDD.t2597 804.731
R21066 VDD.n2229 VDD.t2645 804.731
R21067 VDD.n2358 VDD.t2549 804.731
R21068 VDD.n2431 VDD.t2269 804.731
R21069 VDD.n2418 VDD.t2568 804.731
R21070 VDD.n2415 VDD.t2365 804.731
R21071 VDD.n2439 VDD.t2567 804.731
R21072 VDD.n2407 VDD.t2364 804.731
R21073 VDD.n2476 VDD.t2292 804.731
R21074 VDD.n2479 VDD.t2486 804.731
R21075 VDD.n2109 VDD.t2359 804.731
R21076 VDD.t2423 VDD.n2112 804.731
R21077 VDD.t2358 VDD.n2101 804.731
R21078 VDD.n2104 VDD.t2338 804.731
R21079 VDD.n2129 VDD.t2368 804.731
R21080 VDD.n2132 VDD.t2562 804.731
R21081 VDD.n1344 VDD.t2620 804.731
R21082 VDD.n1454 VDD.t2266 804.731
R21083 VDD.n1748 VDD.t2313 804.731
R21084 VDD.t2524 VDD.n1681 804.731
R21085 VDD.n1612 VDD.t2398 804.731
R21086 VDD.n1591 VDD.t2508 804.731
R21087 VDD.n1658 VDD.t2332 804.731
R21088 VDD.n1661 VDD.t2298 804.731
R21089 VDD.n1318 VDD.t2430 804.731
R21090 VDD.n1338 VDD.t2429 804.731
R21091 VDD.t2573 VDD.n1271 804.731
R21092 VDD.n1295 VDD.t2419 804.731
R21093 VDD.n1298 VDD.t2600 804.731
R21094 VDD.n797 VDD.t2636 804.731
R21095 VDD.t2415 VDD.n908 804.731
R21096 VDD.t2530 VDD.n1120 804.731
R21097 VDD.n661 VDD.t2608 804.731
R21098 VDD.n637 VDD.t2383 804.731
R21099 VDD.n629 VDD.t2474 804.731
R21100 VDD.t2384 VDD.n633 804.731
R21101 VDD.n593 VDD.t2350 804.731
R21102 VDD.n650 VDD.t2396 804.731
R21103 VDD.n773 VDD.t2537 804.731
R21104 VDD.n854 VDD.t2327 804.731
R21105 VDD.n857 VDD.t2260 804.731
R21106 VDD.n462 VDD.t2471 804.731
R21107 VDD.n458 VDD.t2511 804.731
R21108 VDD.t2510 VDD.n453 804.731
R21109 VDD.n485 VDD.t2519 804.731
R21110 VDD.n488 VDD.t2579 804.731
R21111 VDD.n1025 VDD.t1504 804.095
R21112 VDD.n4100 VDD.t1566 803.572
R21113 VDD.n3439 VDD.t2078 803.572
R21114 VDD.n2761 VDD.t872 803.572
R21115 VDD.n1360 VDD.t886 803.572
R21116 VDD.n2024 VDD.t1153 803.572
R21117 VDD.n1464 VDD.t955 803.572
R21118 VDD.n1900 VDD.t1582 803.572
R21119 VDD.n1509 VDD.t723 803.572
R21120 VDD.n555 VDD.t719 803.572
R21121 VDD.n1194 VDD.t721 803.572
R21122 VDD.n951 VDD.t1647 803.572
R21123 VDD.t2360 VDD.t1809 802.298
R21124 VDD.n139 VDD.n138 799.532
R21125 VDD.n1432 VDD.t1791 789.686
R21126 VDD.n1862 VDD.t2814 789.686
R21127 VDD.n1511 VDD.t2962 789.686
R21128 VDD.n1151 VDD.t3013 789.686
R21129 VDD.n1140 VDD.t210 789.686
R21130 VDD.n681 VDD.t1 789.686
R21131 VDD.n140 VDD.n103 787.201
R21132 VDD.n1773 VDD.t599 786.62
R21133 VDD.n1216 VDD.t2890 786.62
R21134 VDD.n1217 VDD.t341 786.62
R21135 VDD.n2223 VDD.t100 780.119
R21136 VDD.t2550 VDD.t3063 778.799
R21137 VDD.t2556 VDD.t2650 778.799
R21138 VDD.t2877 VDD.t2388 775.442
R21139 VDD.n229 VDD.n226 755.294
R21140 VDD.n227 VDD.n221 755.294
R21141 VDD.t2504 VDD.n3798 752.703
R21142 VDD.t2407 VDD.n4181 751.692
R21143 VDD.t2632 VDD.n4239 751.692
R21144 VDD.n3877 VDD.t2488 751.692
R21145 VDD.t2380 VDD.n4062 751.692
R21146 VDD.t2426 VDD.n3791 751.692
R21147 VDD.n3918 VDD.t2361 751.692
R21148 VDD.t2335 VDD.n3578 751.692
R21149 VDD.t2454 VDD.n3581 751.692
R21150 VDD.t2591 VDD.n2374 751.692
R21151 VDD.n2372 VDD.t2592 751.692
R21152 VDD.t2410 VDD.n2369 751.692
R21153 VDD.n2597 VDD.t2389 751.692
R21154 VDD.t2602 VDD.n2226 751.692
R21155 VDD.t2359 VDD.n2108 751.692
R21156 VDD.n2113 VDD.t2423 751.692
R21157 VDD.n2106 VDD.t2358 751.692
R21158 VDD.n1274 VDD.t2573 751.692
R21159 VDD.n909 VDD.t2415 751.692
R21160 VDD.n1121 VDD.t2530 751.692
R21161 VDD.t2608 VDD.n660 751.692
R21162 VDD.t2383 VDD.n636 751.692
R21163 VDD.t2474 VDD.n628 751.692
R21164 VDD.n634 VDD.t2384 751.692
R21165 VDD.t2471 VDD.n461 751.692
R21166 VDD.t2511 VDD.n457 751.692
R21167 VDD.n455 VDD.t2510 751.692
R21168 VDD.n214 VDD.n213 742.777
R21169 VDD.n148 VDD.n106 728.284
R21170 VDD.t2583 VDD.n3692 725.173
R21171 VDD.t2433 VDD.n3738 725.173
R21172 VDD.t2448 VDD.n3829 725.173
R21173 VDD.t2289 VDD.n3849 725.173
R21174 VDD.t2513 VDD.n3852 725.173
R21175 VDD.t2347 VDD.n3674 725.173
R21176 VDD.t2499 VDD.n4391 725.173
R21177 VDD.t2344 VDD.n4394 725.173
R21178 VDD.t2497 VDD.n2923 725.173
R21179 VDD.t2413 VDD.n3049 725.173
R21180 VDD.t2322 VDD.n3052 725.173
R21181 VDD.t2405 VDD.n3041 725.173
R21182 VDD.t2586 VDD.n3069 725.173
R21183 VDD.t2301 VDD.n3600 725.173
R21184 VDD.t2421 VDD.n3603 725.173
R21185 VDD.n2644 VDD.t2614 725.173
R21186 VDD.t2615 VDD.n2646 725.173
R21187 VDD.t2645 VDD.n2228 725.173
R21188 VDD.t2549 VDD.n2357 725.173
R21189 VDD.t2292 VDD.n2475 725.173
R21190 VDD.t2486 VDD.n2478 725.173
R21191 VDD.t2338 VDD.n2103 725.173
R21192 VDD.t2368 VDD.n2128 725.173
R21193 VDD.t2562 VDD.n2131 725.173
R21194 VDD.t2620 VDD.n1343 725.173
R21195 VDD.t2266 VDD.n1453 725.173
R21196 VDD.t2313 VDD.n1747 725.173
R21197 VDD.n1682 VDD.t2524 725.173
R21198 VDD.t2332 VDD.n1657 725.173
R21199 VDD.t2298 VDD.n1660 725.173
R21200 VDD.t2419 VDD.n1294 725.173
R21201 VDD.t2600 VDD.n1297 725.173
R21202 VDD.t2636 VDD.n796 725.173
R21203 VDD.t2350 VDD.n592 725.173
R21204 VDD.t2396 VDD.n649 725.173
R21205 VDD.t2537 VDD.n772 725.173
R21206 VDD.t2327 VDD.n853 725.173
R21207 VDD.t2260 VDD.n856 725.173
R21208 VDD.t2519 VDD.n484 725.173
R21209 VDD.t2579 VDD.n487 725.173
R21210 VDD.t3033 VDD.t1719 725.078
R21211 VDD.n2349 VDD.n2348 721.278
R21212 VDD.n3769 VDD.n3768 713.668
R21213 VDD.n3243 VDD.t2968 700.506
R21214 VDD.n2165 VDD.t2888 700.506
R21215 VDD.n2294 VDD.t18 700.506
R21216 VDD.n1347 VDD.t343 700.506
R21217 VDD.n1944 VDD.t3022 700.506
R21218 VDD.n3354 VDD.t220 699.889
R21219 VDD.n2494 VDD.t981 698.234
R21220 VDD.n2858 VDD.t106 696.322
R21221 VDD.n2650 VDD.t2825 696.322
R21222 VDD.n1779 VDD.t593 696.322
R21223 VDD.n2059 VDD.t2572 694.876
R21224 VDD.n4163 VDD.t163 677.308
R21225 VDD.n2291 VDD.t1748 675.293
R21226 VDD.n1884 VDD.t510 675.293
R21227 VDD.n768 VDD.t1696 675.293
R21228 VDD.n1757 VDD.t1678 674.705
R21229 VDD.n124 VDD.n122 674.119
R21230 VDD.n122 VDD.n113 674.119
R21231 VDD.n157 VDD.t643 672.854
R21232 VDD.n157 VDD.t728 672.77
R21233 VDD.n159 VDD.t2793 671.86
R21234 VDD.n156 VDD.t2796 671.86
R21235 VDD.n4099 VDD.t2946 671.408
R21236 VDD.n3669 VDD.t976 671.408
R21237 VDD.n2093 VDD.t1627 671.408
R21238 VDD.n2873 VDD.t268 671.408
R21239 VDD.n2258 VDD.t2692 671.408
R21240 VDD.n2048 VDD.t761 671.408
R21241 VDD.n724 VDD.t3096 671.408
R21242 VDD.n896 VDD.t2910 671.408
R21243 VDD.n2594 VDD.t2878 669.491
R21244 VDD.n2926 VDD.t2684 668.702
R21245 VDD.n3493 VDD.t1512 667.778
R21246 VDD.n2973 VDD.t1040 667.778
R21247 VDD.n3651 VDD.t1938 667.778
R21248 VDD.n3161 VDD.t1215 667.778
R21249 VDD.n3179 VDD.t1894 667.778
R21250 VDD.n2775 VDD.t1974 667.778
R21251 VDD.n1368 VDD.t1450 667.778
R21252 VDD.n2038 VDD.t1343 667.778
R21253 VDD.n1984 VDD.t2013 667.778
R21254 VDD.n1938 VDD.t1931 667.778
R21255 VDD.n1886 VDD.t829 667.778
R21256 VDD.n1857 VDD.t944 667.778
R21257 VDD.n1724 VDD.t1922 667.778
R21258 VDD.n1725 VDD.t1217 667.778
R21259 VDD.n1237 VDD.t1848 667.778
R21260 VDD.n603 VDD.t1269 667.778
R21261 VDD.n1084 VDD.t1042 667.778
R21262 VDD.n730 VDD.t711 667.778
R21263 VDD.n3472 VDD.t1018 667.751
R21264 VDD.n3449 VDD.t938 667.751
R21265 VDD.n3401 VDD.t838 667.751
R21266 VDD.n2981 VDD.t790 667.751
R21267 VDD.n2984 VDD.t1901 667.751
R21268 VDD.n3527 VDD.t2154 667.751
R21269 VDD.n3530 VDD.t855 667.751
R21270 VDD.n2747 VDD.t715 667.751
R21271 VDD.n1701 VDD.t1073 667.751
R21272 VDD.n1757 VDD.t1496 667.751
R21273 VDD.n1446 VDD.t1164 667.721
R21274 VDD.n1013 VDD.t782 667.721
R21275 VDD.n3270 VDD.t392 665.163
R21276 VDD.n3275 VDD.t545 665.163
R21277 VDD.n4112 VDD.t686 664.455
R21278 VDD.n3154 VDD.t743 664.455
R21279 VDD.n3022 VDD.t1514 664.455
R21280 VDD.n2798 VDD.t1271 664.455
R21281 VDD.n1392 VDD.t797 664.455
R21282 VDD.n1423 VDD.t616 664.455
R21283 VDD.n1469 VDD.t1536 664.455
R21284 VDD.n1912 VDD.t2739 664.455
R21285 VDD.n1832 VDD.t1617 664.455
R21286 VDD.n1699 VDD.t2783 664.455
R21287 VDD.n545 VDD.t2082 664.455
R21288 VDD.n616 VDD.t2184 664.455
R21289 VDD.n1064 VDD.t1850 664.455
R21290 VDD.n938 VDD.t1325 664.455
R21291 VDD.n3744 VDD.t1929 663.426
R21292 VDD.n3425 VDD.t1946 663.426
R21293 VDD.n3377 VDD.t1283 663.426
R21294 VDD.n2971 VDD.t809 663.426
R21295 VDD.n3567 VDD.t2779 663.426
R21296 VDD.n3644 VDD.t1235 663.426
R21297 VDD.n2233 VDD.t1193 663.426
R21298 VDD.n1780 VDD.t1121 663.426
R21299 VDD.n706 VDD.t1486 663.426
R21300 VDD.n2629 VDD.t1782 662.841
R21301 VDD.n3780 VDD.t641 662.22
R21302 VDD.n3281 VDD.t536 662.22
R21303 VDD.n3234 VDD.t405 662.22
R21304 VDD.n759 VDD.t1298 662.22
R21305 VDD.n1955 VDD.t3015 659.593
R21306 VDD.n1827 VDD.t2957 659.593
R21307 VDD.n77 VDD.n65 657.715
R21308 VDD.n41 VDD.n40 657.715
R21309 VDD.n4053 VDD.n4052 656.938
R21310 VDD.n2272 VDD.n2271 656.938
R21311 VDD.n2720 VDD.n2277 656.938
R21312 VDD.n2640 VDD.n2314 656.938
R21313 VDD.n2567 VDD.n2365 656.938
R21314 VDD.n1979 VDD.n1438 656.938
R21315 VDD.n1877 VDD.n1491 656.938
R21316 VDD.n3146 VDD.n3144 653.917
R21317 VDD.n1417 VDD.n1416 653.917
R21318 VDD.n544 VDD.n543 653.917
R21319 VDD.n577 VDD.n537 653.917
R21320 VDD.n76 VDD.n66 647.111
R21321 VDD.n39 VDD.n30 647.111
R21322 VDD.t2455 VDD.t717 636.131
R21323 VDD.n991 VDD.n990 634.25
R21324 VDD.n3704 VDD.n3703 629.801
R21325 VDD.n4319 VDD.n4318 629.801
R21326 VDD.n2920 VDD.n2919 629.801
R21327 VDD.n3460 VDD.n3458 629.801
R21328 VDD.n3362 VDD.n3361 629.801
R21329 VDD.n3414 VDD.n3349 629.801
R21330 VDD.n2991 VDD.n2990 629.801
R21331 VDD.n3566 VDD.n3521 629.801
R21332 VDD.n2172 VDD.n2171 629.801
R21333 VDD.n2197 VDD.n2173 629.801
R21334 VDD.n2256 VDD.n2255 629.801
R21335 VDD.n2740 VDD.n2739 629.801
R21336 VDD.n2300 VDD.n2299 629.801
R21337 VDD.n1369 VDD.n1366 629.801
R21338 VDD.n1804 VDD.n1803 629.801
R21339 VDD.n1097 VDD.n677 629.801
R21340 VDD.t2593 VDD.t2020 624.383
R21341 VDD.t683 VDD.t2400 621.025
R21342 VDD.t2631 VDD.t2110 621.025
R21343 VDD.t2369 VDD.t1150 621.025
R21344 VDD.t2443 VDD.t2461 617.668
R21345 VDD.t2503 VDD.t2425 617.668
R21346 VDD.t2323 VDD.t2479 617.668
R21347 VDD.t2351 VDD.t2514 617.668
R21348 VDD.t2514 VDD.t2434 617.668
R21349 VDD.t2268 VDD.t2566 617.668
R21350 VDD.t2572 VDD.t2428 617.668
R21351 VDD.t2529 VDD.t2607 617.668
R21352 VDD.n2592 VDD.n2346 615.659
R21353 VDD.n2043 VDD.n1408 610.51
R21354 VDD.n4019 VDD.n4018 609.38
R21355 VDD.n2282 VDD.n2281 607.212
R21356 VDD.n2319 VDD.n2318 607.212
R21357 VDD.n2615 VDD.n2614 607.212
R21358 VDD.n2509 VDD.n2393 607.212
R21359 VDD.n1383 VDD.n1359 607.212
R21360 VDD.n2001 VDD.n2000 607.212
R21361 VDD.n1874 VDD.n1496 607.212
R21362 VDD.n1744 VDD.n1550 607.212
R21363 VDD.n4048 VDD.n4047 604.881
R21364 VDD.n1875 VDD.n1494 604.881
R21365 VDD.n4109 VDD.n3734 604.457
R21366 VDD.n2933 VDD.n2932 604.457
R21367 VDD.n3475 VDD.n2942 604.457
R21368 VDD.n3447 VDD.n2956 604.457
R21369 VDD.n3399 VDD.n3357 604.457
R21370 VDD.n3319 VDD.n2980 604.457
R21371 VDD.n3546 VDD.n3532 604.457
R21372 VDD.n3160 VDD.n3159 604.457
R21373 VDD.n3181 VDD.n3180 604.457
R21374 VDD.n2801 VDD.n2244 604.457
R21375 VDD.n1390 VDD.n1389 604.457
R21376 VDD.n1918 VDD.n1468 604.457
R21377 VDD.n1909 VDD.n1471 604.457
R21378 VDD.n1835 VDD.n1513 604.457
R21379 VDD.n1703 VDD.n1702 604.457
R21380 VDD.n1566 VDD.n1565 604.457
R21381 VDD.n1187 VDD.n614 604.457
R21382 VDD.n1066 VDD.n693 604.457
R21383 VDD.n943 VDD.n737 604.457
R21384 VDD.n2929 VDD.n2927 604.394
R21385 VDD.n3344 VDD.n2970 604.394
R21386 VDD.n3523 VDD.n3522 604.394
R21387 VDD.n3575 VDD.n2911 604.394
R21388 VDD.n2252 VDD.n2251 604.394
R21389 VDD.n2080 VDD.n2079 604.394
R21390 VDD.n2043 VDD.n1409 604.394
R21391 VDD.n1943 VDD.n1457 604.394
R21392 VDD.n1489 VDD.n1488 604.394
R21393 VDD.n1729 VDD.n1559 604.394
R21394 VDD.n1731 VDD.n1730 604.394
R21395 VDD.n1787 VDD.n1786 604.394
R21396 VDD.n1232 VDD.n529 604.394
R21397 VDD.n1209 VDD.n600 604.394
R21398 VDD.n1432 VDD.n1431 604.163
R21399 VDD.n1862 VDD.n1502 604.163
R21400 VDD.n681 VDD.n680 604.163
R21401 VDD.n4337 VDD.n4336 604.076
R21402 VDD.n886 VDD.n762 603.619
R21403 VDD.n3226 VDD.n3000 603.231
R21404 VDD.n1810 VDD.n1526 603.231
R21405 VDD.n2732 VDD.n2731 602.457
R21406 VDD.n535 VDD.n534 602.457
R21407 VDD.n2363 VDD.n2362 602.456
R21408 VDD.n2387 VDD.n2386 602.456
R21409 VDD.n3780 VDD.n3779 602.266
R21410 VDD.n2929 VDD.n2928 602.213
R21411 VDD.n1847 VDD.n1846 602.009
R21412 VDD.n3387 VDD.n3386 601.679
R21413 VDD.n3330 VDD.n2975 601.679
R21414 VDD.n3323 VDD.n3322 601.679
R21415 VDD.n3537 VDD.n3536 601.679
R21416 VDD.n2899 VDD.n2898 601.679
R21417 VDD.n3203 VDD.n3015 601.679
R21418 VDD.n3169 VDD.n3168 601.679
R21419 VDD.n3027 VDD.n3026 601.679
R21420 VDD.n1715 VDD.n1714 601.679
R21421 VDD.n1718 VDD.n1717 601.679
R21422 VDD.n1077 VDD.n687 601.679
R21423 VDD.n3143 VDD.n3036 601.585
R21424 VDD.n2279 VDD.n2278 601.585
R21425 VDD.n2316 VDD.n2315 601.585
R21426 VDD.n2564 VDD.n2366 601.585
R21427 VDD.n2023 VDD.n1419 601.585
R21428 VDD.n1976 VDD.n1440 601.585
R21429 VDD.n3748 VDD.n3747 601.097
R21430 VDD.n3371 VDD.n3370 601.097
R21431 VDD.n3369 VDD.n3368 601.097
R21432 VDD.n3338 VDD.n3337 601.097
R21433 VDD.n3645 VDD.n2910 601.097
R21434 VDD.n3153 VDD.n3033 601.097
R21435 VDD.n3186 VDD.n3021 601.097
R21436 VDD.n2831 VDD.n2830 601.097
R21437 VDD.n703 VDD.n702 601.097
R21438 VDD.n973 VDD.n971 601.097
R21439 VDD.n992 VDD.n988 600.304
R21440 VDD.n3503 VDD.n3502 600.105
R21441 VDD.n3314 VDD.n2983 600.105
R21442 VDD.n3551 VDD.n3529 600.105
R21443 VDD.n2754 VDD.n2264 600.105
R21444 VDD.n2016 VDD.n1422 600.105
R21445 VDD.n1965 VDD.n1445 600.105
R21446 VDD.n1760 VDD.n1759 600.105
R21447 VDD.n1017 VDD.n1016 600.105
R21448 VDD.n562 VDD.n547 600.105
R21449 VDD.n4198 VDD.n4197 599.933
R21450 VDD.n564 VDD.n546 599.886
R21451 VDD.n4207 VDD.n4200 599.808
R21452 VDD.n4231 VDD.n4188 599.808
R21453 VDD.n3708 VDD.n3707 599.808
R21454 VDD.n4151 VDD.n4150 599.808
R21455 VDD.n3730 VDD.n3729 599.808
R21456 VDD.n4075 VDD.n4074 599.808
R21457 VDD.n4298 VDD.n4297 599.808
R21458 VDD.n4436 VDD.n4369 599.808
R21459 VDD.n4404 VDD.n4387 599.808
R21460 VDD.n1596 VDD.n1595 599.808
R21461 VDD.n866 VDD.n849 599.808
R21462 VDD.n497 VDD.n480 599.808
R21463 VDD.n3262 VDD.n3261 599.74
R21464 VDD.n3241 VDD.n3240 599.74
R21465 VDD.n3277 VDD.n3276 599.74
R21466 VDD.n3283 VDD.n3282 599.74
R21467 VDD.n2627 VDD.n2324 599.74
R21468 VDD.n1951 VDD.n1451 599.74
R21469 VDD.n1824 VDD.n1518 599.74
R21470 VDD.n3741 VDD.n3740 599.282
R21471 VDD.n3516 VDD.n2915 598.383
R21472 VDD.n3486 VDD.n2935 598.383
R21473 VDD.n3433 VDD.n3432 598.383
R21474 VDD.n2765 VDD.n2764 598.383
R21475 VDD.n1376 VDD.n1363 598.383
R21476 VDD.n2029 VDD.n1415 598.383
R21477 VDD.n1977 VDD.n1439 598.383
R21478 VDD.n1930 VDD.n1463 598.383
R21479 VDD.n1893 VDD.n1892 598.383
R21480 VDD.n1772 VDD.n1542 598.383
R21481 VDD.n445 VDD.n444 598.383
R21482 VDD.n608 VDD.n607 598.383
R21483 VDD.n1031 VDD.n711 598.383
R21484 VDD.n956 VDD.n954 598.383
R21485 VDD.n2814 VDD.n2813 598.274
R21486 VDD.n2583 VDD.n2354 596.567
R21487 VDD.n3983 VDD.n3783 591.962
R21488 VDD.n231 VDD.n184 588.424
R21489 VDD.n3988 VDD.n3987 585
R21490 VDD.n3986 VDD.n3985 585
R21491 VDD.n2577 VDD.n2576 585
R21492 VDD.n2575 VDD.n2574 585
R21493 VDD.n2533 VDD.n2532 585
R21494 VDD.n2531 VDD.n2530 585
R21495 VDD.n211 VDD.n184 573.763
R21496 VDD.n3946 VDD.n3945 564.811
R21497 VDD.n356 VDD.n343 557.648
R21498 VDD.n366 VDD.n343 557.648
R21499 VDD.n366 VDD.n345 557.648
R21500 VDD.n345 VDD.n338 557.648
R21501 VDD.n340 VDD.n338 557.648
R21502 VDD.n378 VDD.n340 557.648
R21503 VDD.n364 VDD.n363 557.648
R21504 VDD.n365 VDD.n364 557.648
R21505 VDD.n365 VDD.n336 557.648
R21506 VDD.n391 VDD.n336 557.648
R21507 VDD.n391 VDD.n337 557.648
R21508 VDD.n374 VDD.n337 557.648
R21509 VDD.n145 VDD.n144 557.184
R21510 VDD.n375 VDD.t3033 556.386
R21511 VDD.n208 VDD.n207 552.283
R21512 VDD.n212 VDD.n208 552.283
R21513 VDD.n214 VDD.n205 552.283
R21514 VDD.n227 VDD.t2941 545.926
R21515 VDD.n229 VDD.t145 545.926
R21516 VDD.t1148 VDD.t162 545.495
R21517 VDD.n3841 VDD.t2500 540.46
R21518 VDD.t2400 VDD.n3840 540.46
R21519 VDD.n114 VDD.n107 504.707
R21520 VDD.n119 VDD.n118 497.493
R21521 VDD.n116 VDD.n110 494.118
R21522 VDD.t2434 VDD.t2001 481.714
R21523 VDD.t1019 VDD.t2828 469.966
R21524 VDD.t1517 VDD.t2351 469.966
R21525 VDD.t2461 VDD.t155 468.286
R21526 VDD.t2479 VDD.t84 468.286
R21527 VDD.n375 VDD.t58 467.601
R21528 VDD.t2811 VDD.t2302 466.608
R21529 VDD.t366 VDD.t2333 466.608
R21530 VDD.t1971 VDD.t2382 466.608
R21531 VDD.t2590 VDD.t2409 463.252
R21532 VDD.t2388 VDD.t2476 463.252
R21533 VDD.t2357 VDD.t2422 463.252
R21534 VDD.t2414 VDD.t2261 463.252
R21535 VDD.t2382 VDD.t2473 463.252
R21536 VDD.n383 VDD.t462 461.5
R21537 VDD.t2241 VDD.n193 451.502
R21538 VDD.n2867 VDD.t267 449.824
R21539 VDD.t1192 VDD.t2114 448.146
R21540 VDD.t1485 VDD.t3067 441.432
R21541 VDD.t710 VDD.t2563 438.075
R21542 VDD.t406 VDD.t2030 436.397
R21543 VDD.t1603 VDD.t323 433.039
R21544 VDD.n410 VDD.t3034 431.428
R21545 VDD.t462 VDD.t2768 419.767
R21546 VDD.t151 VDD.t146 409.875
R21547 VDD.t151 VDD.t148 409.875
R21548 VDD.t2673 VDD.t692 397.793
R21549 VDD.n3915 VDD.t2502 396.406
R21550 VDD.n4142 VDD.t2481 396.348
R21551 VDD.n3687 VDD.t2353 396.348
R21552 VDD.n2699 VDD.t2307 392.87
R21553 VDD.t227 VDD.t651 392.757
R21554 VDD.t1136 VDD.t2287 391.079
R21555 VDD.t2091 VDD.t2342 391.079
R21556 VDD.t1857 VDD.t2320 391.079
R21557 VDD.t1595 VDD.t2299 391.079
R21558 VDD.t1284 VDD.t2290 391.079
R21559 VDD.t1303 VDD.t2366 391.079
R21560 VDD.t1062 VDD.t2296 391.079
R21561 VDD.t879 VDD.t2417 391.079
R21562 VDD.t1380 VDD.t2258 391.079
R21563 VDD.t887 VDD.t2517 391.079
R21564 VDD.n3914 VDD.t2501 391.005
R21565 VDD.n667 VDD.t2371 390.875
R21566 VDD.n4242 VDD.t2408 389.521
R21567 VDD.n3959 VDD.t2402 389.521
R21568 VDD.n1125 VDD.t2531 389.521
R21569 VDD.t675 VDD.t1232 389.399
R21570 VDD.t2520 VDD.t2675 389.399
R21571 VDD.t1926 VDD.t1935 389.399
R21572 VDD.t2634 VDD.t603 389.399
R21573 VDD.t1985 VDD.n875 389.399
R21574 VDD.t94 VDD.t2348 389.399
R21575 VDD.n3795 VDD.t2505 389.046
R21576 VDD.n4060 VDD.t2381 388.851
R21577 VDD.n911 VDD.t2416 388.776
R21578 VDD.n4192 VDD.t2594 388.656
R21579 VDD.n4196 VDD.t2595 388.656
R21580 VDD.n4128 VDD.t2324 388.656
R21581 VDD.n3723 VDD.t2325 388.656
R21582 VDD.n4071 VDD.t2377 388.656
R21583 VDD.n4082 VDD.t2378 388.656
R21584 VDD.n4310 VDD.t2539 388.656
R21585 VDD.n4315 VDD.t2540 388.656
R21586 VDD.n4253 VDD.t2438 388.656
R21587 VDD.n4261 VDD.t2439 388.656
R21588 VDD.n4015 VDD.t2554 388.656
R21589 VDD.n3766 VDD.t2555 388.656
R21590 VDD.n4055 VDD.t2303 388.656
R21591 VDD.n4065 VDD.t2304 388.656
R21592 VDD.n3969 VDD.t2427 388.656
R21593 VDD.n3802 VDD.t2401 388.656
R21594 VDD.n2847 VDD.t2603 388.656
R21595 VDD.n2693 VDD.t2306 388.656
R21596 VDD.n2606 VDD.t2390 388.656
R21597 VDD.n2565 VDD.t2411 388.656
R21598 VDD.n2547 VDD.t2641 388.656
R21599 VDD.n2378 VDD.t2642 388.656
R21600 VDD.n1962 VDD.t2542 388.656
R21601 VDD.n1443 VDD.t2543 388.656
R21602 VDD.n1466 VDD.t2611 388.656
R21603 VDD.n1931 VDD.t2612 388.656
R21604 VDD.n1849 VDD.t2386 388.656
R21605 VDD.n1855 VDD.t2387 388.656
R21606 VDD.n1626 VDD.t2557 388.656
R21607 VDD.n1590 VDD.t2558 388.656
R21608 VDD.n1330 VDD.t2574 388.656
R21609 VDD.n623 VDD.t2475 388.656
R21610 VDD.n749 VDD.t2262 388.656
R21611 VDD.n919 VDD.t2263 388.656
R21612 VDD.n819 VDD.t2638 388.656
R21613 VDD.n804 VDD.t2639 388.656
R21614 VDD.n522 VDD.t2472 388.656
R21615 VDD.n4230 VDD.t2633 388.656
R21616 VDD.n4140 VDD.t2480 388.656
R21617 VDD.n3885 VDD.t2489 388.656
R21618 VDD.n4268 VDD.t2352 388.656
R21619 VDD.n3764 VDD.t2278 388.656
R21620 VDD.n4039 VDD.t2279 388.656
R21621 VDD.n3926 VDD.t2362 388.656
R21622 VDD.n3352 VDD.t2521 388.656
R21623 VDD.n3407 VDD.t2522 388.656
R21624 VDD.n3255 VDD.t2483 388.656
R21625 VDD.n3247 VDD.t2484 388.656
R21626 VDD.n3136 VDD.t2545 388.656
R21627 VDD.n3145 VDD.t2546 388.656
R21628 VDD.n3189 VDD.t2294 388.656
R21629 VDD.n3195 VDD.t2295 388.656
R21630 VDD.n2816 VDD.t2374 388.656
R21631 VDD.n2822 VDD.t2375 388.656
R21632 VDD.n2784 VDD.t2392 388.656
R21633 VDD.n2792 VDD.t2393 388.656
R21634 VDD.n2723 VDD.t2533 388.656
R21635 VDD.n2729 VDD.t2534 388.656
R21636 VDD.n2701 VDD.t2315 388.656
R21637 VDD.n2708 VDD.t2316 388.656
R21638 VDD.n2306 VDD.t2492 388.656
R21639 VDD.n2656 VDD.t2493 388.656
R21640 VDD.n2407 VDD.t2551 388.656
R21641 VDD.n2411 VDD.t2552 388.656
R21642 VDD.n2157 VDD.t2424 388.656
R21643 VDD.n2067 VDD.t2281 388.656
R21644 VDD.n1270 VDD.t2282 388.656
R21645 VDD.n532 VDD.t2318 388.656
R21646 VDD.n582 VDD.t2319 388.656
R21647 VDD.n1167 VDD.t2340 388.656
R21648 VDD.n619 VDD.t2341 388.656
R21649 VDD.n1133 VDD.t2609 388.656
R21650 VDD.n1107 VDD.t2370 388.656
R21651 VDD.n1052 VDD.t2329 388.656
R21652 VDD.n1059 VDD.t2330 388.656
R21653 VDD.n1015 VDD.t2355 388.656
R21654 VDD.n1024 VDD.t2356 388.656
R21655 VDD.n994 VDD.t2272 388.656
R21656 VDD.n719 VDD.t2273 388.656
R21657 VDD.n968 VDD.t2564 388.656
R21658 VDD.n972 VDD.t2565 388.656
R21659 VDD.n950 VDD.t2605 388.656
R21660 VDD.n955 VDD.t2606 388.656
R21661 VDD.n925 VDD.t2450 388.656
R21662 VDD.n742 VDD.t2451 388.656
R21663 VDD.n383 VDD.t58 387.856
R21664 VDD.n3577 VDD.t2334 387.682
R21665 VDD.n3580 VDD.t2453 387.682
R21666 VDD.n2494 VDD.t2268 386.043
R21667 VDD.n2376 VDD.t2590 386.043
R21668 VDD.t2613 VDD.t2491 386.043
R21669 VDD.n2287 VDD.t2314 386.043
R21670 VDD.t2336 VDD.t2357 386.043
R21671 VDD.t1305 VDD.t2271 386.043
R21672 VDD.t2686 VDD.t2794 384.365
R21673 VDD.t726 VDD.t64 384.365
R21674 VDD.n1684 VDD.t2525 382.673
R21675 VDD.n446 VDD.t2309 381.443
R21676 VDD.n1239 VDD.t2310 381.443
R21677 VDD.n1145 VDD.t2570 381.443
R21678 VDD.n642 VDD.t2571 381.443
R21679 VDD.n2031 VDD.t2576 381.443
R21680 VDD.n2036 VDD.t2577 381.443
R21681 VDD.n1346 VDD.t2621 381.44
R21682 VDD.n3691 VDD.t2582 380.193
R21683 VDD.n3737 VDD.t2432 380.193
R21684 VDD.n3828 VDD.t2447 380.193
R21685 VDD.n3848 VDD.t2288 380.193
R21686 VDD.n3851 VDD.t2512 380.193
R21687 VDD.n3673 VDD.t2346 380.193
R21688 VDD.n4390 VDD.t2498 380.193
R21689 VDD.n4393 VDD.t2343 380.193
R21690 VDD.n2922 VDD.t2496 380.193
R21691 VDD.n3048 VDD.t2412 380.193
R21692 VDD.n3051 VDD.t2321 380.193
R21693 VDD.n3040 VDD.t2404 380.193
R21694 VDD.n3068 VDD.t2585 380.193
R21695 VDD.n3599 VDD.t2300 380.193
R21696 VDD.n3602 VDD.t2420 380.193
R21697 VDD.n2227 VDD.t2644 380.193
R21698 VDD.n2356 VDD.t2548 380.193
R21699 VDD.n2474 VDD.t2291 380.193
R21700 VDD.n2477 VDD.t2485 380.193
R21701 VDD.n2102 VDD.t2337 380.193
R21702 VDD.n2127 VDD.t2367 380.193
R21703 VDD.n2130 VDD.t2561 380.193
R21704 VDD.n1452 VDD.t2265 380.193
R21705 VDD.n1746 VDD.t2312 380.193
R21706 VDD.n1656 VDD.t2331 380.193
R21707 VDD.n1659 VDD.t2297 380.193
R21708 VDD.n1293 VDD.t2418 380.193
R21709 VDD.n1296 VDD.t2599 380.193
R21710 VDD.n795 VDD.t2635 380.193
R21711 VDD.n591 VDD.t2349 380.193
R21712 VDD.n648 VDD.t2395 380.193
R21713 VDD.n771 VDD.t2536 380.193
R21714 VDD.n852 VDD.t2326 380.193
R21715 VDD.n855 VDD.t2259 380.193
R21716 VDD.n483 VDD.t2518 380.193
R21717 VDD.n486 VDD.t2578 380.193
R21718 VDD.t893 VDD.t975 379.329
R21719 VDD.t1499 VDD.t1495 360.866
R21720 VDD.t793 VDD.t557 359.188
R21721 VDD.t3099 VDD.t2024 359.188
R21722 VDD.t269 VDD.t1307 359.188
R21723 VDD.n3217 VDD.t732 355.392
R21724 VDD.n2851 VDD.t1872 355.392
R21725 VDD.n351 VDD.n348 353.156
R21726 VDD.n1051 VDD.t1108 350.841
R21727 VDD.n1349 VDD.t1560 350.582
R21728 VDD.n1998 VDD.t1411 350.582
R21729 VDD.n1949 VDD.t1664 350.582
R21730 VDD.n1902 VDD.t912 350.582
R21731 VDD.n1520 VDD.t1239 350.582
R21732 VDD.n1572 VDD.t1570 350.582
R21733 VDD.n3459 VDD.t1760 350.582
R21734 VDD.n1686 VDD.t1824 350.582
R21735 VDD.n1001 VDD.t1184 350.582
R21736 VDD.n1173 VDD.t2170 350.582
R21737 VDD.n927 VDD.t1907 350.582
R21738 VDD.n2554 VDD.t1921 349.507
R21739 VDD.n695 VDD.t1102 348.312
R21740 VDD.n1354 VDD.t1556 347.572
R21741 VDD.n2008 VDD.t1409 347.572
R21742 VDD.n1957 VDD.t1660 347.572
R21743 VDD.n1911 VDD.t906 347.572
R21744 VDD.n1515 VDD.t1241 347.572
R21745 VDD.n1698 VDD.t1568 347.572
R21746 VDD.n2944 VDD.t1758 347.57
R21747 VDD.n1568 VDD.t1820 347.57
R21748 VDD.n1182 VDD.t2174 347.57
R21749 VDD.n716 VDD.t1182 347.57
R21750 VDD.n937 VDD.t1905 347.57
R21751 VDD.t731 VDD.t402 347.438
R21752 VDD.n901 VDD.t495 345.884
R21753 VDD.n894 VDD.t1337 345.884
R21754 VDD.n4212 VDD.t1349 344.06
R21755 VDD.n4164 VDD.t1168 344.06
R21756 VDD.n4119 VDD.t1001 344.06
R21757 VDD.n4334 VDD.t803 344.06
R21758 VDD.n3451 VDD.t942 343.579
R21759 VDD.n3558 VDD.t1625 343.579
R21760 VDD.n3152 VDD.t637 343.579
R21761 VDD.n2746 VDD.t2195 343.579
R21762 VDD.n3354 VDD.t1331 343.577
R21763 VDD.n3307 VDD.t866 343.577
R21764 VDD.n3187 VDD.t821 343.577
R21765 VDD.n2246 VDD.t1275 343.577
R21766 VDD.n569 VDD.t753 343.577
R21767 VDD.n324 VDD.n184 343.467
R21768 VDD.t1442 VDD.t3019 342.404
R21769 VDD.n2238 VDD.t1776 341.43
R21770 VDD.n3676 VDD.t2186 340.536
R21771 VDD.n2926 VDD.t1388 340.45
R21772 VDD.n4157 VDD.t1149 340.243
R21773 VDD.n4081 VDD.t2749 340.243
R21774 VDD.n1606 VDD.t138 340.243
R21775 VDD.n851 VDD.t2785 340.243
R21776 VDD.n482 VDD.t932 340.243
R21777 VDD.n4186 VDD.t1862 340.241
R21778 VDD.n4295 VDD.t2002 340.241
R21779 VDD.n4372 VDD.t1948 340.241
R21780 VDD.n4389 VDD.t1311 340.241
R21781 VDD.n4117 VDD.t1970 340.012
R21782 VDD.n3312 VDD.t1014 340.012
R21783 VDD.n1751 VDD.t1500 340.012
R21784 VDD.n3553 VDD.t1069 340.01
R21785 VDD.n1917 VDD.t1223 340.01
R21786 VDD.t1783 VDD.t2339 339.046
R21787 VDD.n2585 VDD.t1833 338.08
R21788 VDD.n325 VDD.n324 337.423
R21789 VDD.n1736 VDD.t1321 336.567
R21790 VDD.n2592 VDD.t37 336.267
R21791 VDD.n3936 VDD.t1897 333.368
R21792 VDD.n2936 VDD.t1510 333.368
R21793 VDD.t2748 VDD.t26 330.654
R21794 VDD.t1977 VDD.t1811 330.654
R21795 VDD.t3023 VDD.t2694 330.654
R21796 VDD.t2112 VDD.t300 330.654
R21797 VDD.n3015 VDD.t493 329.938
R21798 VDD.n3887 VDD.t3121 328.036
R21799 VDD.n2433 VDD.t3133 327.947
R21800 VDD.t1947 VDD.t2440 327.298
R21801 VDD.t1659 VDD.t1163 327.298
R21802 VDD.n1007 VDD.n1006 326.279
R21803 VDD.n59 VDD.n54 326.158
R21804 VDD.n20 VDD.n19 326.158
R21805 VDD.n4103 VDD.n4102 325.627
R21806 VDD.n2686 VDD.n2293 325.627
R21807 VDD.n1487 VDD.n1486 325.627
R21808 VDD.n893 VDD.n758 325.627
R21809 VDD.n1398 VDD.n1350 323.988
R21810 VDD.n1426 VDD.n1425 323.988
R21811 VDD.n1449 VDD.n1448 323.988
R21812 VDD.n1908 VDD.n1473 323.988
R21813 VDD.n1825 VDD.n1517 323.988
R21814 VDD.n1693 VDD.n1570 323.988
R21815 VDD.n3466 VDD.n2946 323.986
R21816 VDD.n1691 VDD.n1571 323.986
R21817 VDD.n1057 VDD.n697 323.986
R21818 VDD.n1176 VDD.n1175 323.986
R21819 VDD.n930 VDD.n929 323.986
R21820 VDD.n4166 VDD.n3710 322.329
R21821 VDD.n4460 VDD.n3665 322.329
R21822 VDD.n2184 VDD.n2179 322.329
R21823 VDD.n2098 VDD.n2097 322.329
R21824 VDD.n2762 VDD.n2260 322.329
R21825 VDD.n2052 VDD.n2051 322.329
R21826 VDD.n1546 VDD.n1545 322.329
R21827 VDD.n877 VDD.n770 322.329
R21828 VDD.t1579 VDD.t356 322.262
R21829 VDD.t1775 VDD.n2237 322.262
R21830 VDD.t70 VDD.t278 322.262
R21831 VDD.t280 VDD.t2870 322.262
R21832 VDD.t129 VDD.t262 322.262
R21833 VDD.t260 VDD.t3027 322.262
R21834 VDD.n2806 VDD.n2240 320.976
R21835 VDD.n2242 VDD.n2241 320.976
R21836 VDD.n2799 VDD.n2245 320.976
R21837 VDD.n412 VDD.n411 320.976
R21838 VDD.n427 VDD.n415 320.976
R21839 VDD.n52 VDD.n48 320.976
R21840 VDD.n23 VDD.n22 320.976
R21841 VDD.t117 VDD.t1280 318.906
R21842 VDD.t2293 VDD.t548 318.906
R21843 VDD.t2016 VDD.t1786 318.906
R21844 VDD.t2873 VDD.t1422 318.906
R21845 VDD.t1364 VDD.t1320 318.906
R21846 VDD.t3029 VDD.t1140 318.906
R21847 VDD.n94 VDD.n92 318.303
R21848 VDD.n3448 VDD.n2953 317.755
R21849 VDD.t1539 VDD.t1372 317.226
R21850 VDD.t195 VDD.t923 317.226
R21851 VDD.t2043 VDD.t321 317.226
R21852 VDD.t1023 VDD.t125 317.226
R21853 VDD.t1453 VDD.t368 317.226
R21854 VDD.t2151 VDD.t538 317.226
R21855 VDD.t957 VDD.t2305 317.226
R21856 VDD.t671 VDD.t306 317.226
R21857 VDD.t1941 VDD.t873 317.226
R21858 VDD.t735 VDD.t2122 317.226
R21859 VDD.n3395 VDD.n3394 317.104
R21860 VDD.n3204 VDD.n3014 317.104
R21861 VDD.n2213 VDD.n2212 317.104
R21862 VDD.n2738 VDD.n2270 317.104
R21863 VDD.n2692 VDD.n2290 317.104
R21864 VDD.n3212 VDD.n3010 317.103
R21865 VDD.n2207 VDD.n2205 317.103
R21866 VDD.t3081 VDD.t314 315.548
R21867 VDD.t276 VDD.t107 315.548
R21868 VDD.t2625 VDD.t1896 315.548
R21869 VDD.t1896 VDD.t1895 315.548
R21870 VDD.t20 VDD.t270 315.548
R21871 VDD.t3025 VDD.t1481 315.548
R21872 VDD.t1827 VDD.t2967 315.548
R21873 VDD.t22 VDD.t2701 315.548
R21874 VDD.t197 VDD.t1134 315.548
R21875 VDD.t364 VDD.t1387 315.548
R21876 VDD.t2704 VDD.t1975 315.548
R21877 VDD.t1711 VDD.t1047 315.548
R21878 VDD.t496 VDD.t1813 315.548
R21879 VDD.t1837 VDD.t1196 315.548
R21880 VDD.t2824 VDD.t1117 315.548
R21881 VDD.t1118 VDD.t17 315.548
R21882 VDD.t2422 VDD.t72 315.548
R21883 VDD.t592 VDD.t691 315.548
R21884 VDD.t12 VDD.t2663 315.548
R21885 VDD.t1278 VDD.t681 315.548
R21886 VDD.t972 VDD.t1475 315.548
R21887 VDD.t1366 VDD.t474 315.548
R21888 VDD.t901 VDD.t486 315.548
R21889 VDD.t1541 VDD.t466 315.548
R21890 VDD.t358 VDD.t335 315.548
R21891 VDD.t478 VDD.t344 315.548
R21892 VDD.t66 VDD.t897 315.548
R21893 VDD.n3996 VDD.n3776 315.406
R21894 VDD.n1937 VDD.n1460 315.406
R21895 VDD.n2221 VDD.n2220 315.221
R21896 VDD.n595 VDD.n594 315.221
R21897 VDD.n1085 VDD.n683 315.221
R21898 VDD.n1985 VDD.n1434 315.221
R21899 VDD.n1504 VDD.n1503 315.221
R21900 VDD.n1777 VDD.n1540 315.221
R21901 VDD.n598 VDD.n597 315.221
R21902 VDD.n1153 VDD.n638 315.221
R21903 VDD.n4361 VDD.n4309 313.942
R21904 VDD.t2222 VDD.t2637 313.87
R21905 VDD.n2573 VDD.n2361 313.591
R21906 VDD.n2529 VDD.n2385 313.591
R21907 VDD.n755 VDD.n754 313.574
R21908 VDD.n3248 VDD.n3246 313.217
R21909 VDD.n2659 VDD.n2658 313.217
R21910 VDD.n1355 VDD.n1353 313.217
R21911 VDD.n1789 VDD.n1788 313.217
R21912 VDD.n3210 VDD.n3011 312.981
R21913 VDD.n4003 VDD.n3773 312.978
R21914 VDD.n4278 VDD.t3212 312.89
R21915 VDD.n4348 VDD.n4347 312.829
R21916 VDD.n3805 VDD.n3804 312.827
R21917 VDD.n3301 VDD.n2989 312.827
R21918 VDD.n426 VDD.n424 312.699
R21919 VDD.t2440 VDD.t617 312.192
R21920 VDD.t1330 VDD.t2520 312.192
R21921 VDD.t2476 VDD.t44 312.192
R21922 VDD.t2391 VDD.t1274 312.192
R21923 VDD.t350 VDD.t2464 312.192
R21924 VDD.t423 VDD.t99 312.192
R21925 VDD.t425 VDD.t3012 312.192
R21926 VDD.t352 VDD.t2509 312.192
R21927 VDD.n3833 VDD.n3832 312.053
R21928 VDD.n3836 VDD.n3835 312.053
R21929 VDD.n3847 VDD.n3846 312.053
R21930 VDD.n3952 VDD.n3951 312.053
R21931 VDD.n4416 VDD.n4379 312.053
R21932 VDD.n4410 VDD.n4383 312.053
R21933 VDD.n3225 VDD.n3003 312.053
R21934 VDD.n3060 VDD.n3059 312.053
R21935 VDD.n3615 VDD.n3593 312.053
R21936 VDD.n3609 VDD.n3597 312.053
R21937 VDD.n2586 VDD.n2351 312.053
R21938 VDD.n2491 VDD.n2467 312.053
R21939 VDD.n2484 VDD.n2472 312.053
R21940 VDD.n2143 VDD.n2121 312.053
R21941 VDD.n2137 VDD.n2125 312.053
R21942 VDD.n1524 VDD.n1523 312.053
R21943 VDD.n1673 VDD.n1649 312.053
R21944 VDD.n1666 VDD.n1654 312.053
R21945 VDD.n1309 VDD.n1287 312.053
R21946 VDD.n1303 VDD.n1291 312.053
R21947 VDD.n451 VDD.n450 312.053
R21948 VDD.n589 VDD.n588 312.053
R21949 VDD.n1201 VDD.n606 312.053
R21950 VDD.n1152 VDD.n640 312.053
R21951 VDD.n1139 VDD.n654 312.053
R21952 VDD.n673 VDD.n672 312.053
R21953 VDD.n1071 VDD.n690 312.053
R21954 VDD.n979 VDD.n727 312.053
R21955 VDD.n962 VDD.n732 312.053
R21956 VDD.n887 VDD.n761 312.053
R21957 VDD.n883 VDD.n767 312.053
R21958 VDD.n840 VDD.n779 312.053
R21959 VDD.n834 VDD.n783 312.053
R21960 VDD.n826 VDD.n789 312.053
R21961 VDD.n517 VDD.n467 312.053
R21962 VDD.n470 VDD.n469 312.053
R21963 VDD.n474 VDD.n473 312.053
R21964 VDD.n3833 VDD.n3831 312.051
R21965 VDD.n3863 VDD.n3844 312.051
R21966 VDD.n3847 VDD.n3845 312.051
R21967 VDD.n4010 VDD.n4009 312.051
R21968 VDD.n3758 VDD.n3757 312.051
R21969 VDD.n3975 VDD.n3786 312.051
R21970 VDD.n4381 VDD.n4380 312.051
R21971 VDD.n3060 VDD.n3058 312.051
R21972 VDD.n3615 VDD.n3591 312.051
R21973 VDD.n3609 VDD.n3596 312.051
R21974 VDD.n2462 VDD.n2401 312.051
R21975 VDD.n2484 VDD.n2470 312.051
R21976 VDD.n2143 VDD.n2120 312.051
R21977 VDD.n2137 VDD.n2124 312.051
R21978 VDD.n1642 VDD.n1580 312.051
R21979 VDD.n1797 VDD.n1533 312.051
R21980 VDD.n1666 VDD.n1652 312.051
R21981 VDD.n1309 VDD.n1286 312.051
R21982 VDD.n1303 VDD.n1290 312.051
R21983 VDD.n840 VDD.n778 312.051
R21984 VDD.n835 VDD.n782 312.051
R21985 VDD.n786 VDD.n785 312.051
R21986 VDD.n509 VDD.n472 312.051
R21987 VDD.n503 VDD.n476 312.051
R21988 VDD.n1142 VDD.n646 311.767
R21989 VDD.n847 VDD.n846 311.659
R21990 VDD.n478 VDD.n477 311.659
R21991 VDD.n4205 VDD.n4201 311.659
R21992 VDD.n4190 VDD.n4189 311.659
R21993 VDD.n4171 VDD.n3706 311.659
R21994 VDD.n4342 VDD.n4341 311.659
R21995 VDD.n4304 VDD.n4303 311.659
R21996 VDD.n4385 VDD.n4384 311.659
R21997 VDD.n3441 VDD.n2959 311.519
R21998 VDD.n1833 VDD.n1514 310.868
R21999 VDD.n3928 VDD.t3150 310.842
R22000 VDD.t1734 VDD.t2656 310.512
R22001 VDD.n2628 VDD.n2321 310.486
R22002 VDD.n1357 VDD.n1356 310.486
R22003 VDD.n1411 VDD.n1410 310.486
R22004 VDD.n1869 VDD.n1499 310.486
R22005 VDD.n1739 VDD.n1738 310.486
R22006 VDD.n3480 VDD.n2939 309.726
R22007 VDD.n1552 VDD.n1551 309.726
R22008 VDD.n3874 VDD.n3826 309.654
R22009 VDD.n3699 VDD.n3697 309.531
R22010 VDD.n3415 VDD.n3348 309.531
R22011 VDD.n2539 VDD.n2382 309.531
R22012 VDD.n1899 VDD.n1476 309.531
R22013 VDD.n4092 VDD.n3743 309.531
R22014 VDD.n3905 VDD.n3816 309.531
R22015 VDD.n2859 VDD.n2857 309.526
R22016 VDD.n4419 VDD.n4418 309.483
R22017 VDD.n3875 VDD.n3825 309.399
R22018 VDD.t2500 VDD.t2360 308.834
R22019 VDD.t1340 VDD.t1264 308.834
R22020 VDD.n4251 VDD.t2581 308.834
R22021 VDD.t2981 VDD.t391 308.834
R22022 VDD.t2363 VDD.t2550 308.834
R22023 VDD.n2311 VDD.t2613 308.834
R22024 VDD.n2867 VDD.t2336 308.834
R22025 VDD.n1676 VDD.t2523 308.834
R22026 VDD.t2523 VDD.t1823 308.834
R22027 VDD.t1918 VDD.t2535 308.834
R22028 VDD.t2652 VDD.t1297 308.834
R22029 VDD.n875 VDD.t1906 308.834
R22030 VDD.n701 VDD.t1107 308.834
R22031 VDD.t2394 VDD.n645 308.834
R22032 VDD.t2509 VDD.t2470 308.834
R22033 VDD.n357 VDD.n353 308.8
R22034 VDD.n1480 VDD.n1479 308.767
R22035 VDD.n4402 VDD.n4388 308.755
R22036 VDD.n3044 VDD.n3043 308.755
R22037 VDD.n523 VDD.n464 308.755
R22038 VDD.n576 VDD.n538 308.755
R22039 VDD.n1193 VDD.n610 308.755
R22040 VDD.n1183 VDD.n618 308.755
R22041 VDD.n1124 VDD.n664 308.755
R22042 VDD.n1065 VDD.n694 308.755
R22043 VDD.n1045 VDD.n705 308.755
R22044 VDD.n1009 VDD.n718 308.755
R22045 VDD.n917 VDD.n746 308.755
R22046 VDD.n552 VDD.n550 308.755
R22047 VDD.n1160 VDD.n625 308.755
R22048 VDD.n1032 VDD.n710 308.755
R22049 VDD.n740 VDD.n739 308.755
R22050 VDD.n801 VDD.n800 308.755
R22051 VDD.n4425 VDD.n4375 308.755
R22052 VDD.n4087 VDD.n3746 308.755
R22053 VDD.n3066 VDD.n3065 308.755
R22054 VDD.n864 VDD.n850 308.755
R22055 VDD.n495 VDD.n481 308.755
R22056 VDD.n4149 VDD.n3716 308.151
R22057 VDD.n4073 VDD.n3752 308.151
R22058 VDD.n1599 VDD.n1597 308.151
R22059 VDD.n4111 VDD.n3732 308.149
R22060 VDD.n4368 VDD.n4367 308.149
R22061 VDD.n2327 VDD.n2326 307.204
R22062 VDD.n423 VDD.n416 307.204
R22063 VDD.n1819 VDD.n1522 307.204
R22064 VDD.n2707 VDD.n2284 306.976
R22065 VDD.n2612 VDD.n2331 306.976
R22066 VDD.n2503 VDD.n2502 306.976
R22067 VDD.n1997 VDD.n1428 306.976
R22068 VDD.n3717 VDD.t3221 306.735
R22069 VDD.n3893 VDD.t3119 306.735
R22070 VDD.n4325 VDD.t3159 306.735
R22071 VDD.n3683 VDD.t3126 306.735
R22072 VDD.n4032 VDD.t3114 306.735
R22073 VDD.n4370 VDD.t3191 306.735
R22074 VDD.n3119 VDD.t3143 306.735
R22075 VDD.n3073 VDD.t3220 306.735
R22076 VDD.n3081 VDD.t3199 306.735
R22077 VDD.n3099 VDD.t3238 306.735
R22078 VDD.n3585 VDD.t3217 306.735
R22079 VDD.n3585 VDD.t3128 306.735
R22080 VDD.n2181 VDD.t3149 306.735
R22081 VDD.n2231 VDD.t3195 306.735
R22082 VDD.n2667 VDD.t3235 306.735
R22083 VDD.n2334 VDD.t3219 306.735
R22084 VDD.n2394 VDD.t3139 306.735
R22085 VDD.n2425 VDD.t3138 306.735
R22086 VDD.n2409 VDD.t3209 306.735
R22087 VDD.n1586 VDD.t3236 306.735
R22088 VDD.n1605 VDD.t3182 306.735
R22089 VDD.n1278 VDD.t3225 306.735
R22090 VDD.n3456 VDD.n2949 306.541
R22091 VDD.n3968 VDD.n3789 306.428
R22092 VDD.n4126 VDD.n4125 304.731
R22093 VDD.t2703 VDD.t411 300.442
R22094 VDD.n794 VDD.n792 298.538
R22095 VDD.t298 VDD.t2945 297.086
R22096 VDD.t2538 VDD.t2191 295.406
R22097 VDD.n4126 VDD.n3726 295.255
R22098 VDD.n794 VDD.n793 295.051
R22099 VDD.n3945 VDD.n3944 294.281
R22100 VDD.t1216 VDD.t630 293.728
R22101 VDD.t1058 VDD.n3839 292.05
R22102 VDD.t2495 VDD.t2683 287.014
R22103 VDD.t1025 VDD.t213 278.623
R22104 VDD.t1501 VDD.t2899 278.623
R22105 VDD.t562 VDD.t802 276.943
R22106 VDD.t1240 VDD.t1483 275.265
R22107 VDD.t1101 VDD.t377 275.265
R22108 VDD.t1511 VDD.t2856 271.909
R22109 VDD.t1408 VDD.t1992 270.231
R22110 VDD.t2941 VDD.n219 265.26
R22111 VDD.t145 VDD.n219 265.26
R22112 VDD.t2738 VDD.t1535 265.195
R22113 VDD.t852 VDD.t764 265.195
R22114 VDD.t2919 VDD.n193 265.195
R22115 VDD.n418 VDD.t463 262.932
R22116 VDD.n119 VDD.n103 262.401
R22117 VDD.t1530 VDD.t1601 260.159
R22118 VDD.n95 VDD.t1538 256.884
R22119 VDD.t1503 VDD.t1841 256.803
R22120 VDD.n3220 VDD.t546 255.905
R22121 VDD.n2399 VDD.t273 255.905
R22122 VDD.n2150 VDD.t281 255.905
R22123 VDD.n2118 VDD.t2936 255.905
R22124 VDD.n1579 VDD.t2955 255.905
R22125 VDD.n1284 VDD.t3030 255.905
R22126 VDD.n162 VDD.t1473 255.905
R22127 VDD.n93 VDD.t1805 255.905
R22128 VDD.n101 VDD.t2132 255.905
R22129 VDD.n4176 VDD.t1552 255.904
R22130 VDD.n4316 VDD.t1956 255.904
R22131 VDD.n3430 VDD.t1446 255.904
R22132 VDD.n3220 VDD.t407 255.904
R22133 VDD.n2459 VDD.t3066 255.904
R22134 VDD.n2150 VDD.t312 255.904
R22135 VDD.n2118 VDD.t2874 255.904
R22136 VDD.n1632 VDD.t2649 255.904
R22137 VDD.n1638 VDD.t112 255.904
R22138 VDD.n1284 VDD.t3104 255.904
R22139 VDD.n805 VDD.t476 255.904
R22140 VDD.n516 VDD.t543 255.904
R22141 VDD.n162 VDD.t727 255.904
R22142 VDD.n99 VDD.t2687 255.904
R22143 VDD.n59 VDD.t827 255.904
R22144 VDD.n20 VDD.t1317 255.904
R22145 VDD.t2194 VDD.t2045 255.125
R22146 VDD.n2460 VDD.t472 254.907
R22147 VDD.n4190 VDD.t2019 254.232
R22148 VDD.n4304 VDD.t2099 254.232
R22149 VDD.n847 VDD.t2869 254.232
R22150 VDD.n2387 VDD.t1808 254.019
R22151 VDD.n826 VDD.t1031 254.019
R22152 VDD.n470 VDD.t608 254.019
R22153 VDD.n2268 VDD.t1472 253.202
R22154 VDD.n4224 VDD.t2021 252.95
R22155 VDD.n3218 VDD.t552 252.95
R22156 VDD.n2461 VDD.t275 252.95
R22157 VDD.n2458 VDD.t468 252.95
R22158 VDD.n2115 VDD.t279 252.95
R22159 VDD.n2149 VDD.t2934 252.95
R22160 VDD.n1631 VDD.t311 252.95
R22161 VDD.n1637 VDD.t2952 252.95
R22162 VDD.n1315 VDD.t3028 252.95
R22163 VDD.n3701 VDD.t1550 252.948
R22164 VDD.n4349 VDD.t1958 252.948
R22165 VDD.n3218 VDD.t403 252.948
R22166 VDD.n2457 VDD.t3064 252.948
R22167 VDD.n2115 VDD.t313 252.948
R22168 VDD.n2149 VDD.t2871 252.948
R22169 VDD.n1315 VDD.t3106 252.948
R22170 VDD.n790 VDD.t1033 252.948
R22171 VDD.n872 VDD.t2866 252.948
R22172 VDD.n465 VDD.t541 252.948
R22173 VDD.n515 VDD.t606 252.403
R22174 VDD.t1646 VDD.t2604 251.768
R22175 VDD.n1642 VDD.t371 251.516
R22176 VDD.n2491 VDD.t382 251.516
R22177 VDD.n1673 VDD.t3077 251.516
R22178 VDD.n3672 VDD.t892 250.724
R22179 VDD.n3689 VDD.t1518 250.724
R22180 VDD.n1582 VDD.t309 250.724
R22181 VDD.n1644 VDD.t373 250.724
R22182 VDD.n234 VDD.t2918 250.724
R22183 VDD.n2785 VDD.t1787 250.722
R22184 VDD.n2468 VDD.t384 250.722
R22185 VDD.n2156 VDD.t71 250.722
R22186 VDD.n1650 VDD.t3073 250.722
R22187 VDD.n1324 VDD.t130 250.722
R22188 VDD.n1317 VDD.t261 250.722
R22189 VDD.n1630 VDD.t2651 250.609
R22190 VDD.t1000 VDD.n3837 250.089
R22191 VDD.n3134 VDD.t1029 250.089
R22192 VDD.t2142 VDD.n1230 250.089
R22193 VDD.n2960 VDD.t1250 249.451
R22194 VDD.n3868 VDD.t2798 249.363
R22195 VDD.n3862 VDD.t1688 249.363
R22196 VDD.n3856 VDD.t1137 249.363
R22197 VDD.n3047 VDD.t1858 249.363
R22198 VDD.n3594 VDD.t1454 249.363
R22199 VDD.n3598 VDD.t1596 249.363
R22200 VDD.n2584 VDD.t2084 249.363
R22201 VDD.n2473 VDD.t2726 249.363
R22202 VDD.n2122 VDD.t672 249.363
R22203 VDD.n2126 VDD.t1304 249.363
R22204 VDD.n1655 VDD.t2073 249.363
R22205 VDD.n1288 VDD.t736 249.363
R22206 VDD.n1292 VDD.t1522 249.363
R22207 VDD.n1141 VDD.t1876 249.363
R22208 VDD.n1099 VDD.t2233 249.363
R22209 VDD.n691 VDD.t654 249.363
R22210 VDD.n885 VDD.t2657 249.363
R22211 VDD.n776 VDD.t870 249.363
R22212 VDD.n780 VDD.t1480 249.363
R22213 VDD.n828 VDD.t2700 249.363
R22214 VDD.n515 VDD.t2659 249.363
R22215 VDD.n165 VDD.t2929 249.363
R22216 VDD.n3868 VDD.t971 249.362
R22217 VDD.n3856 VDD.t1705 249.362
R22218 VDD.n3017 VDD.t397 249.362
R22219 VDD.n3047 VDD.t2730 249.362
R22220 VDD.n3594 VDD.t1609 249.362
R22221 VDD.n3598 VDD.t2256 249.362
R22222 VDD.n2460 VDD.t815 249.362
R22223 VDD.n2473 VDD.t1285 249.362
R22224 VDD.n2122 VDD.t1378 249.362
R22225 VDD.n2126 VDD.t2068 249.362
R22226 VDD.n1655 VDD.t1063 249.362
R22227 VDD.n1288 VDD.t988 249.362
R22228 VDD.n1292 VDD.t880 249.362
R22229 VDD.n776 VDD.t666 249.362
R22230 VDD.n833 VDD.t1966 249.362
R22231 VDD.n827 VDD.t1892 249.362
R22232 VDD.n165 VDD.t65 249.362
R22233 VDD.n2246 VDD.t251 249.202
R22234 VDD.n774 VDD.t481 249.118
R22235 VDD.n53 VDD.t3051 248.843
R22236 VDD.n24 VDD.t3047 248.843
R22237 VDD.n60 VDD.t2757 248.843
R22238 VDD.n21 VDD.t2723 248.843
R22239 VDD.n4385 VDD.t2747 248.688
R22240 VDD.n478 VDD.t2141 248.686
R22241 VDD.t1719 VDD.t1713 248.599
R22242 VDD.t1713 VDD.t1715 248.599
R22243 VDD.t1715 VDD.t1717 248.599
R22244 VDD.n4381 VDD.t664 248.475
R22245 VDD.n509 VDD.t2164 248.475
R22246 VDD.n503 VDD.t700 248.475
R22247 VDD.n4416 VDD.t2775 248.475
R22248 VDD.n4410 VDD.t1176 248.475
R22249 VDD.n474 VDD.t768 248.475
R22250 VDD.n4447 VDD.t894 248.219
R22251 VDD.n4260 VDD.t1516 248.219
R22252 VDD.n3676 VDD.t2101 248.219
R22253 VDD.n2963 VDD.t1441 248.219
R22254 VDD.n2790 VDD.t1772 248.219
R22255 VDD.n2522 VDD.t1812 248.219
R22256 VDD.n2159 VDD.t73 248.219
R22257 VDD.n1636 VDD.t110 248.219
R22258 VDD.n1279 VDD.t128 248.219
R22259 VDD.n1281 VDD.t263 248.219
R22260 VDD.n56 VDD.t825 248.219
R22261 VDD.n16 VDD.t1319 248.219
R22262 VDD.n1343 VDD.t3172 247.744
R22263 VDD.n1682 VDD.t3155 247.744
R22264 VDD.n163 VDD.t1806 247.394
R22265 VDD.n163 VDD.t1803 247.394
R22266 VDD.n264 VDD.n251 247.387
R22267 VDD.n262 VDD.n255 247.316
R22268 VDD.n3784 VDD.t1341 246.946
R22269 VDD.n884 VDD.t1735 246.946
R22270 VDD.t2046 VDD.t2905 246.732
R22271 VDD.n132 VDD.t726 246.732
R22272 VDD.n3995 VDD.t2984 246.512
R22273 VDD.n1223 VDD.t1255 246.077
R22274 VDD.n3692 VDD.t3239 245.667
R22275 VDD.n3738 VDD.t3198 245.667
R22276 VDD.n3829 VDD.t3227 245.667
R22277 VDD.n3849 VDD.t3226 245.667
R22278 VDD.n3852 VDD.t3116 245.667
R22279 VDD.n3674 VDD.t3129 245.667
R22280 VDD.n4391 VDD.t3211 245.667
R22281 VDD.n4394 VDD.t3131 245.667
R22282 VDD.n2923 VDD.t3165 245.667
R22283 VDD.n3049 VDD.t3207 245.667
R22284 VDD.n3052 VDD.t3201 245.667
R22285 VDD.n3041 VDD.t3125 245.667
R22286 VDD.n3069 VDD.t3203 245.667
R22287 VDD.n3600 VDD.t3168 245.667
R22288 VDD.n3603 VDD.t3170 245.667
R22289 VDD.n2228 VDD.t3153 245.667
R22290 VDD.n2357 VDD.t3218 245.667
R22291 VDD.n2475 VDD.t3122 245.667
R22292 VDD.n2478 VDD.t3214 245.667
R22293 VDD.n2103 VDD.t3123 245.667
R22294 VDD.n2128 VDD.t3190 245.667
R22295 VDD.n2131 VDD.t3113 245.667
R22296 VDD.n1453 VDD.t3167 245.667
R22297 VDD.n1747 VDD.t3158 245.667
R22298 VDD.n1657 VDD.t3151 245.667
R22299 VDD.n1660 VDD.t3206 245.667
R22300 VDD.n1294 VDD.t3202 245.667
R22301 VDD.n1297 VDD.t3162 245.667
R22302 VDD.n796 VDD.t3177 245.667
R22303 VDD.n592 VDD.t3223 245.667
R22304 VDD.n649 VDD.t3132 245.667
R22305 VDD.n772 VDD.t3194 245.667
R22306 VDD.n853 VDD.t3140 245.667
R22307 VDD.n856 VDD.t3233 245.667
R22308 VDD.n484 VDD.t3231 245.667
R22309 VDD.n487 VDD.t3135 245.667
R22310 VDD.n4397 VDD.t2092 245.178
R22311 VDD.n3044 VDD.t1024 245.178
R22312 VDD.n2486 VDD.t2152 245.178
R22313 VDD.n1818 VDD.t1649 245.178
R22314 VDD.n1668 VDD.t1942 245.178
R22315 VDD.n1250 VDD.t878 245.178
R22316 VDD.n1196 VDD.t1641 245.178
R22317 VDD.n626 VDD.t840 245.178
R22318 VDD.n712 VDD.t1842 245.178
R22319 VDD.n981 VDD.t2802 245.178
R22320 VDD.n935 VDD.t848 245.178
R22321 VDD.n811 VDD.t2223 245.178
R22322 VDD.n3066 VDD.t1077 245.178
R22323 VDD.n1577 VDD.t1458 245.178
R22324 VDD.n859 VDD.t1381 245.178
R22325 VDD.n490 VDD.t888 245.178
R22326 VDD.n410 VDD.t1720 244.737
R22327 VDD.n421 VDD.t1732 244.737
R22328 VDD.n570 VDD.t96 243.512
R22329 VDD.n1208 VDD.t2892 243.512
R22330 VDD.n1079 VDD.t216 243.512
R22331 VDD.n735 VDD.t2964 243.512
R22332 VDD.n752 VDD.t612 243.512
R22333 VDD.n1224 VDD.t347 243.512
R22334 VDD.n980 VDD.t2820 243.512
R22335 VDD.n3196 VDD.t549 243.508
R22336 VDD.n1413 VDD.t3175 242.282
R22337 VDD.n449 VDD.t3154 242.282
R22338 VDD.n1146 VDD.t3112 242.282
R22339 VDD.t1601 VDD.t2839 241.696
R22340 VDD.t181 VDD.t756 241.696
R22341 VDD.n2546 VDD.t1814 240.792
R22342 VDD.n4218 VDD.t1527 240.215
R22343 VDD.n3929 VDD.t1810 240.215
R22344 VDD.n1039 VDD.t9 240.215
R22345 VDD.n417 VDD.t2769 240.215
R22346 VDD.n2540 VDD.t1672 240.214
R22347 VDD.n1166 VDD.t1784 240.214
R22348 VDD.n1132 VDD.t1443 240.214
R22349 VDD.n1113 VDD.t3011 240.214
R22350 VDD.n3296 VDD.t1338 240.018
R22351 VDD.n2207 VDD.n2206 239.132
R22352 VDD.n3307 VDD.n2986 238.815
R22353 VDD.n3558 VDD.n3525 238.815
R22354 VDD.n3344 VDD.n2969 238.544
R22355 VDD.t2100 VDD.t2345 238.339
R22356 VDD.n4364 VDD.t891 238.339
R22357 VDD.n874 VDD.t2865 238.339
R22358 VDD.n201 VDD.n198 238.169
R22359 VDD.n3842 VDD.t970 236.661
R22360 VDD.n3838 VDD.t76 236.661
R22361 VDD.n3837 VDD.t1981 236.661
R22362 VDD.n4251 VDD.t738 236.661
R22363 VDD.n4364 VDD.t895 236.661
R22364 VDD.t1076 VDD.n3132 236.661
R22365 VDD.t1457 VDD.n1675 236.661
R22366 VDD.n1676 VDD.t56 236.661
R22367 VDD.t665 VDD.n874 236.661
R22368 VDD.t702 VDD.t191 236.661
R22369 VDD.t2348 VDD.t1254 236.661
R22370 VDD.n132 VDD.t2131 236.661
R22371 VDD.n2645 VDD.t3204 236.231
R22372 VDD.n3699 VDD.n3698 235.248
R22373 VDD.n4328 VDD.n4324 235.248
R22374 VDD.n3515 VDD.n2916 235.248
R22375 VDD.n3474 VDD.n2943 235.248
R22376 VDD.n3378 VDD.n3365 235.248
R22377 VDD.n2190 VDD.n2176 235.248
R22378 VDD.n2782 VDD.n2250 235.248
R22379 VDD.n2753 VDD.n2265 235.248
R22380 VDD.n2679 VDD.n2296 235.248
R22381 VDD.n2068 VDD.n1267 235.248
R22382 VDD.n1795 VDD.n1534 235.248
R22383 VDD.n1106 VDD.n671 235.248
R22384 VDD.t1034 VDD.n3841 234.982
R22385 VDD.n3839 VDD.t1332 234.982
R22386 VDD.t2133 VDD.t1114 234.982
R22387 VDD.t820 VDD.n3133 234.982
R22388 VDD.t1218 VDD.n3295 234.982
R22389 VDD.t1898 VDD.t2218 234.982
R22390 VDD.t1463 VDD.n3421 234.982
R22391 VDD.t1211 VDD.t1230 234.982
R22392 VDD.n3423 VDD.t360 234.982
R22393 VDD.t2239 VDD.t1027 234.982
R22394 VDD.t2681 VDD.t690 234.982
R22395 VDD.t979 VDD.t830 234.982
R22396 VDD.t1251 VDD.n2493 234.982
R22397 VDD.t1920 VDD.n2376 234.982
R22398 VDD.t806 VDD.t1546 234.982
R22399 VDD.n1556 VDD.t1988 234.982
R22400 VDD.t706 VDD.t953 234.982
R22401 VDD.t203 VDD.n1482 234.982
R22402 VDD.t2830 VDD.n1481 234.982
R22403 VDD.t1154 VDD.t2062 234.982
R22404 VDD.t342 VDD.n2058 234.982
R22405 VDD.t34 VDD.n701 234.982
R22406 VDD.n645 VDD.t1444 234.982
R22407 VDD.n1230 VDD.t479 234.982
R22408 VDD.t2229 VDD.t1707 234.982
R22409 VDD.n405 VDD.t60 234.042
R22410 VDD.n397 VDD.t63 234.042
R22411 VDD.n5 VDD.t487 233.349
R22412 VDD.n82 VDD.t374 233.347
R22413 VDD.t2610 VDD.t2204 233.304
R22414 VDD.n405 VDD.t59 232.798
R22415 VDD.n397 VDD.t62 232.798
R22416 VDD.n3840 VDD.t2503 231.625
R22417 VDD.t2379 VDD.n3838 231.625
R22418 VDD.t2581 VDD.t2437 231.625
R22419 VDD.t744 VDD.n2345 231.625
R22420 VDD.t2805 VDD.t2596 231.625
R22421 VDD.t2619 VDD.t2280 231.625
R22422 VDD.t2271 VDD.t1183 231.625
R22423 VDD.n329 VDD.t2920 230.201
R22424 VDD.t2311 VDD.t1202 229.947
R22425 VDD.n3295 VDD.t1851 228.269
R22426 VDD.n2866 VDD.t105 228.269
R22427 VDD.t2734 VDD.t509 228.269
R22428 VDD.n133 VDD.t146 227.642
R22429 VDD.n136 VDD.t148 227.642
R22430 VDD.t1629 VDD.t760 226.59
R22431 VDD.t2120 VDD.t318 224.912
R22432 VDD.t1916 VDD.t123 224.912
R22433 VDD.n3228 VDD.n2997 223.868
R22434 VDD.n1529 VDD.n1528 223.868
R22435 VDD.t2801 VDD.t3095 223.233
R22436 VDD.n4205 VDD.n4204 223.025
R22437 VDD.n318 VDD.n182 222.655
R22438 VDD.t740 VDD.t2373 221.555
R22439 VDD.t1467 VDD.t2385 221.555
R22440 VDD.t1695 VDD.t1004 221.555
R22441 VDD.n230 VDD.n225 220.613
R22442 VDD.n225 VDD.n224 220.613
R22443 VDD.t2596 VDD.t1626 218.198
R22444 VDD.n118 VDD.n105 215.041
R22445 VDD.n909 VDD.t3179 214.929
R22446 VDD.n4062 VDD.t3136 213.977
R22447 VDD.t1794 VDD.t1900 213.163
R22448 VDD.t2153 VDD.t810 213.163
R22449 VDD.t1830 VDD.t781 213.163
R22450 VDD.n3578 VDD.t3173 213.148
R22451 VDD.n3581 VDD.t3127 213.148
R22452 VDD.n3867 VDD.n3842 213.119
R22453 VDD.n4250 VDD.n4249 213.119
R22454 VDD.n3132 VDD.n3131 213.119
R22455 VDD.n3297 VDD.n3296 213.119
R22456 VDD.n3424 VDD.n3423 213.119
R22457 VDD.n3573 VDD.n3572 213.119
R22458 VDD.n2555 VDD.n2376 213.119
R22459 VDD.n2641 VDD.n2311 213.119
R22460 VDD.n2756 VDD.n2263 213.119
R22461 VDD.n2866 VDD.n2865 213.119
R22462 VDD.n2493 VDD.n2492 213.119
R22463 VDD.n2058 VDD.n2057 213.119
R22464 VDD.n1675 VDD.n1674 213.119
R22465 VDD.n3422 VDD.n2940 213.119
R22466 VDD.n3421 VDD.n3420 213.119
R22467 VDD.n3295 VDD.n3294 213.119
R22468 VDD.n2868 VDD.n2867 213.119
R22469 VDD.n2593 VDD.n2345 213.119
R22470 VDD.n1481 VDD.n1429 213.119
R22471 VDD.n1891 VDD.n1483 213.119
R22472 VDD.n1188 VDD.n613 213.119
R22473 VDD.n1098 VDD.n676 213.119
R22474 VDD.n3575 VDD.n3574 212.665
R22475 VDD.n1232 VDD.n1231 212.665
R22476 VDD.n1736 VDD.n1556 212.567
R22477 VDD.n3838 VDD.n3753 211.732
R22478 VDD.n3135 VDD.n3134 211.732
R22479 VDD.n2060 VDD.n2059 211.732
R22480 VDD.n4129 VDD.t3130 210.964
R22481 VDD.n4016 VDD.t3160 210.964
R22482 VDD.n3755 VDD.t3215 210.964
R22483 VDD.n3914 VDD.t3142 210.964
R22484 VDD.n3353 VDD.t3144 210.964
R22485 VDD.n3254 VDD.t3111 210.964
R22486 VDD.n3188 VDD.t3169 210.964
R22487 VDD.n2815 VDD.t3228 210.964
R22488 VDD.n2248 VDD.t3108 210.964
R22489 VDD.n2722 VDD.t3124 210.964
R22490 VDD.n2700 VDD.t3210 210.964
R22491 VDD.n2288 VDD.t3166 210.964
R22492 VDD.n2548 VDD.t3163 210.964
R22493 VDD.n2066 VDD.t3200 210.964
R22494 VDD.n1963 VDD.t3232 210.964
R22495 VDD.n1848 VDD.t3205 210.964
R22496 VDD.n533 VDD.t3107 210.964
R22497 VDD.n698 VDD.t3161 210.964
R22498 VDD.n969 VDD.t3171 210.964
R22499 VDD.n952 VDD.t3157 210.964
R22500 VDD.n926 VDD.t3243 210.964
R22501 VDD.n3840 VDD.n3794 210.524
R22502 VDD.n272 VDD.n271 209.963
R22503 VDD.n1482 VDD.n1480 209.55
R22504 VDD.n4363 VDD.n4362 209.368
R22505 VDD.n3133 VDD.n3019 209.368
R22506 VDD.n2812 VDD.n2237 209.368
R22507 VDD.n2698 VDD.n2287 209.368
R22508 VDD.n2495 VDD.n2494 209.368
R22509 VDD.n1555 VDD.n1535 209.368
R22510 VDD.n1677 VDD.n1676 209.368
R22511 VDD.n1844 VDD.n1508 209.368
R22512 VDD.n985 VDD.n723 209.368
R22513 VDD.n876 VDD.t1918 209.368
R22514 VDD.n2373 VDD.t3145 208.409
R22515 VDD.n456 VDD.t3184 208.409
R22516 VDD.t2425 VDD.t984 208.127
R22517 VDD.t2494 VDD.n256 206.778
R22518 VDD.t2646 VDD.n253 206.778
R22519 VDD.n393 VDD.n333 206.683
R22520 VDD.n368 VDD.n333 206.683
R22521 VDD.n3720 VDD.t3213 206.546
R22522 VDD.n4266 VDD.t3192 206.546
R22523 VDD.t837 VDD.t219 206.45
R22524 VDD.n3423 VDD.t1945 206.45
R22525 VDD.n9 VDD.t3185 204.755
R22526 VDD.n81 VDD.t3189 204.751
R22527 VDD.n6 VDD.t3216 202.582
R22528 VDD.n83 VDD.t3174 202.581
R22529 VDD.n84 VDD.t3188 202.576
R22530 VDD.n7 VDD.t3120 202.573
R22531 VDD.n50 VDD.n49 201.373
R22532 VDD.n12 VDD.n11 201.373
R22533 VDD.t215 VDD.t2148 198.058
R22534 VDD.t2891 VDD.t2070 194.701
R22535 VDD.t1299 VDD.t731 193.022
R22536 VDD.n212 VDD.n211 190.494
R22537 VDD.n213 VDD.n212 190.494
R22538 VDD.t752 VDD.t95 187.987
R22539 VDD.n361 VDD.n360 187.482
R22540 VDD.n360 VDD.n342 187.482
R22541 VDD.n388 VDD.n370 187.482
R22542 VDD.n129 VDD.n117 187.107
R22543 VDD.n126 VDD.n125 187.107
R22544 VDD.n388 VDD.n335 186.73
R22545 VDD.n358 VDD.n352 185.882
R22546 VDD.n358 VDD.n347 185.882
R22547 VDD.t964 VDD.t762 184.63
R22548 VDD.t559 VDD.t2845 184.63
R22549 VDD.n233 VDD.n232 184.056
R22550 VDD.t2580 VDD.n258 183.653
R22551 VDD.n258 VDD.t2286 183.653
R22552 VDD.t923 VDD.t2843 182.952
R22553 VDD.t1232 VDD.t1402 182.952
R22554 VDD.t981 VDD.t590 182.952
R22555 VDD.t44 VDD.t2826 182.952
R22556 VDD.t694 VDD.t1118 182.952
R22557 VDD.t533 VDD.t3017 182.952
R22558 VDD.t1935 VDD.t962 182.952
R22559 VDD.t1089 VDD.t2885 182.952
R22560 VDD.t1131 VDD.t338 182.952
R22561 VDD.t851 VDD.t1591 182.952
R22562 VDD.t1845 VDD.t1006 182.952
R22563 VDD.t649 VDD.t901 182.952
R22564 VDD.n389 VDD.n341 182.309
R22565 VDD.n377 VDD.n341 182.309
R22566 VDD.t1967 VDD.t294 181.273
R22567 VDD.t282 VDD.t634 181.273
R22568 VDD.t818 VDD.t573 181.273
R22569 VDD.t286 VDD.t867 181.273
R22570 VDD.t939 VDD.t2200 181.273
R22571 VDD.t179 VDD.t1755 181.273
R22572 VDD.t1622 VDD.t2857 181.273
R22573 VDD.t791 VDD.t1291 181.273
R22574 VDD.t1520 VDD.t417 181.273
R22575 VDD.t2895 VDD.t2776 181.273
R22576 VDD.t389 VDD.t1926 181.273
R22577 VDD.t413 VDD.t2805 181.273
R22578 VDD.t2208 VDD.t903 181.273
R22579 VDD.t2903 VDD.t1414 181.273
R22580 VDD.t1918 VDD.t304 181.273
R22581 VDD.t1697 VDD.t1693 181.273
R22582 VDD.t80 VDD.t1908 181.273
R22583 VDD.t1294 VDD.t1305 181.273
R22584 VDD.t296 VDD.t1177 181.273
R22585 VDD.t284 VDD.t1109 181.273
R22586 VDD.t175 VDD.t2171 181.273
R22587 VDD.n138 VDD.n103 179.327
R22588 VDD.n373 VDD.n371 178.008
R22589 VDD.n362 VDD.n349 178.008
R22590 VDD.t1002 VDD.t716 177.916
R22591 VDD.t1491 VDD.t1228 177.916
R22592 VDD.t1887 VDD.t302 176.238
R22593 VDD.t610 VDD.t2414 176.238
R22594 VDD.t613 VDD.t2083 174.559
R22595 VDD.t2914 VDD.t101 174.559
R22596 VDD.t722 VDD.n1508 174.559
R22597 VDD.t737 VDD.t951 174.559
R22598 VDD.t1402 VDD.t562 172.881
R22599 VDD.t558 VDD.t1583 172.881
R22600 VDD.t2677 VDD.t560 172.881
R22601 VDD.t1389 VDD.t2849 172.881
R22602 VDD.t1628 VDD.t2837 172.881
R22603 VDD.t2851 VDD.t974 172.881
R22604 VDD.t557 VDD.t694 172.881
R22605 VDD.t762 VDD.t2833 172.881
R22606 VDD.t962 VDD.t559 172.881
R22607 VDD.t1567 VDD.t2782 172.881
R22608 VDD.t490 VDD.t1497 172.881
R22609 VDD.t2665 VDD.t40 172.881
R22610 VDD.t1785 VDD.t1530 171.202
R22611 VDD.t1051 VDD.t1095 171.202
R22612 VDD.t2663 VDD.t696 169.524
R22613 VDD.n3966 VDD.n3790 169.398
R22614 VDD.n2842 VDD.n2841 169.398
R22615 VDD.n627 VDD.n626 169.296
R22616 VDD.t2988 VDD.t153 167.845
R22617 VDD.t13 VDD.t537 167.845
R22618 VDD.t308 VDD.t109 167.845
R22619 VDD.t24 VDD.t424 167.845
R22620 VDD.t201 VDD.t430 167.845
R22621 VDD.t32 VDD.t432 167.845
R22622 VDD.t2227 VDD.t3040 167.845
R22623 VDD.n268 VDD.n251 166.901
R22624 VDD.n255 VDD.n249 166.611
R22625 VDD.t1220 VDD.t1599 166.167
R22626 VDD.t2219 VDD.t2118 166.167
R22627 VDD.t2669 VDD.t1488 166.167
R22628 VDD.t1228 VDD.t1210 166.167
R22629 VDD.t687 VDD.t3089 166.167
R22630 VDD.t622 VDD.t980 166.167
R22631 VDD.t1075 VDD.t1578 166.167
R22632 VDD.t471 VDD.t814 166.167
R22633 VDD.t1745 VDD.t2728 166.167
R22634 VDD.t1543 VDD.t871 166.167
R22635 VDD.t2117 VDD.t2124 166.167
R22636 VDD.t1880 VDD.t1416 166.167
R22637 VDD.t669 VDD.t704 166.167
R22638 VDD.t1612 VDD.t1465 166.167
R22639 VDD.t1050 VDD.t2737 166.167
R22640 VDD.t1581 VDD.t2736 166.167
R22641 VDD.t950 VDD.t954 166.167
R22642 VDD.t945 VDD.t1162 166.167
R22643 VDD.t883 VDD.t851 166.167
R22644 VDD.t1370 VDD.t1646 166.167
R22645 VDD.t1098 VDD.t1503 166.167
R22646 VDD.t2148 VDD.t1939 166.167
R22647 VDD.t2069 VDD.t1611 166.167
R22648 VDD.t718 VDD.t2226 166.167
R22649 VDD.t2658 VDD.t605 166.167
R22650 VDD.t863 VDD.t117 164.488
R22651 VDD.t1743 VDD.t1765 164.488
R22652 VDD.t1424 VDD.t1064 164.488
R22653 VDD.t1426 VDD.t626 164.488
R22654 VDD.t554 VDD.t395 164.488
R22655 VDD.t1338 VDD.t2817 164.488
R22656 VDD.t1669 VDD.t1681 164.488
R22657 VDD.t3102 VDD.t1701 164.488
R22658 VDD.t1691 VDD.t1997 164.488
R22659 VDD.t10 VDD.t2673 164.488
R22660 VDD.t223 VDD.t957 164.488
R22661 VDD.t1528 VDD.t2128 164.488
R22662 VDD.t1524 VDD.t1469 164.488
R22663 VDD.t1157 VDD.t2973 164.488
R22664 VDD.t2954 VDD.t1709 164.488
R22665 VDD.t1979 VDD.t97 164.488
R22666 VDD.t624 VDD.t1032 164.488
R22667 VDD.t475 VDD.t1226 164.488
R22668 VDD.t2010 VDD.t1631 164.488
R22669 VDD.n123 VDD.t642 164.072
R22670 VDD.t1959 VDD.t1086 162.81
R22671 VDD.t2065 VDD.t594 162.81
R22672 VDD.t1064 VDD.t288 162.81
R22673 VDD.t575 VDD.t1426 162.81
R22674 VDD.t411 VDD.t3088 162.81
R22675 VDD.t1027 VDD.t2214 162.81
R22676 VDD.t320 VDD.t941 162.81
R22677 VDD.t1703 VDD.t2971 162.81
R22678 VDD.t1867 VDD.t6 162.81
R22679 VDD.t2716 VDD.t3023 162.81
R22680 VDD.t2863 VDD.t740 162.81
R22681 VDD.t49 VDD.t1418 162.81
R22682 VDD.t290 VDD.t1467 162.81
R22683 VDD.t1723 VDD.t221 162.81
R22684 VDD.t2204 VDD.t706 162.81
R22685 VDD.t645 VDD.t2022 162.81
R22686 VDD.t42 VDD.t1916 162.81
R22687 VDD.t1055 VDD.t90 162.81
R22688 VDD.t2036 VDD.t1340 161.131
R22689 VDD.t2034 VDD.t783 161.131
R22690 VDD.t76 VDD.t2750 161.131
R22691 VDD.t1169 VDD.t1553 161.131
R22692 VDD.t2847 VDD.t1683 161.131
R22693 VDD.t899 VDD.t1865 161.131
R22694 VDD.t738 VDD.t1350 161.131
R22695 VDD.t2437 VDD.t1515 161.131
R22696 VDD.t1999 VDD.t1322 161.131
R22697 VDD.t798 VDD.t1959 161.131
R22698 VDD.t895 VDD.t1951 161.131
R22699 VDD.t2049 VDD.t1314 161.131
R22700 VDD.t594 VDD.t636 161.131
R22701 VDD.t1207 VDD.t326 161.131
R22702 VDD.t716 VDD.t1124 161.131
R22703 VDD.t2967 VDD.t333 161.131
R22704 VDD.t1585 VDD.t1587 161.131
R22705 VDD.t712 VDD.t2841 161.131
R22706 VDD.t2161 VDD.t2028 161.131
R22707 VDD.t2943 VDD.t748 161.131
R22708 VDD.t692 VDD.t1129 161.131
R22709 VDD.t164 VDD.t657 161.131
R22710 VDD.t566 VDD.t2855 161.131
R22711 VDD.t1122 VDD.t964 161.131
R22712 VDD.t2845 VDD.t638 161.131
R22713 VDD.t56 VDD.t139 161.131
R22714 VDD.t773 VDD.t1043 161.131
R22715 VDD.t1043 VDD.t170 161.131
R22716 VDD.t2428 VDD.t127 161.131
R22717 VDD.t1432 VDD.t2786 161.131
R22718 VDD.t2977 VDD.t929 161.131
R22719 VDD.n3987 VDD.n3986 159.476
R22720 VDD.n2532 VDD.n2531 159.476
R22721 VDD.n2576 VDD.n2575 159.476
R22722 VDD.t314 VDD.t1138 159.452
R22723 VDD.t968 VDD.t276 159.452
R22724 VDD.t155 VDD.t1036 159.452
R22725 VDD.t783 VDD.t550 159.452
R22726 VDD.t1981 VDD.t1189 159.452
R22727 VDD.t270 VDD.t2772 159.452
R22728 VDD.t3074 VDD.t661 159.452
R22729 VDD.t379 VDD.t1173 159.452
R22730 VDD.t469 VDD.t2744 159.452
R22731 VDD.t125 VDD.t1855 159.452
R22732 VDD.t3031 VDD.t1021 159.452
R22733 VDD.t264 VDD.t1078 159.452
R22734 VDD.t113 VDD.t1451 159.452
R22735 VDD.t368 VDD.t1597 159.452
R22736 VDD.t538 VDD.t1286 159.452
R22737 VDD.t503 VDD.t1679 159.452
R22738 VDD.t1047 VDD.t1288 159.452
R22739 VDD.t2912 VDD.t488 159.452
R22740 VDD.t167 VDD.t10 159.452
R22741 VDD.t169 VDD.t223 159.452
R22742 VDD.t336 VDD.t330 159.452
R22743 VDD.t1422 VDD.t673 159.452
R22744 VDD.t306 VDD.t1301 159.452
R22745 VDD.t873 VDD.t1060 159.452
R22746 VDD.t1198 VDD.t1650 159.452
R22747 VDD.t2179 VDD.t47 159.452
R22748 VDD.t1140 VDD.t733 159.452
R22749 VDD.t2122 VDD.t881 159.452
R22750 VDD.t681 VDD.t667 159.452
R22751 VDD.t1889 VDD.t972 159.452
R22752 VDD.t2695 VDD.t2697 159.452
R22753 VDD.t1226 VDD.t2224 159.452
R22754 VDD.t494 VDD.t485 159.452
R22755 VDD.t1398 VDD.t1873 159.452
R22756 VDD.t2473 VDD.t839 159.452
R22757 VDD.t841 VDD.t1541 159.452
R22758 VDD.t1642 VDD.t1994 159.452
R22759 VDD.t875 VDD.t966 159.452
R22760 VDD.t2732 VDD.t2165 159.452
R22761 VDD.t765 VDD.t769 159.452
R22762 VDD.t3083 VDD.t697 159.452
R22763 VDD.t1636 VDD.t2138 159.452
R22764 VDD.t1685 VDD.t2487 157.774
R22765 VDD.t2983 VDD.t409 157.774
R22766 VDD.t1881 VDD.t381 157.774
R22767 VDD.t2601 VDD.t2911 157.774
R22768 VDD.t99 VDD.t228 157.774
R22769 VDD.t1326 VDD.t3076 157.774
R22770 VDD.t1709 VDD.t370 157.774
R22771 VDD.t598 VDD.t54 157.774
R22772 VDD.t2921 VDD.t773 157.774
R22773 VDD.t238 VDD.t2813 157.774
R22774 VDD.t234 VDD.t1790 157.774
R22775 VDD.t2280 VDD.t1845 157.774
R22776 VDD.t230 VDD.t0 157.774
R22777 VDD.t232 VDD.t340 157.774
R22778 VDD.t2889 VDD.t240 157.774
R22779 VDD.t2470 VDD.t2742 157.774
R22780 VDD.t2544 VDD.t2063 156.095
R22781 VDD.t1832 VDD.t2161 156.095
R22782 VDD.n1508 VDD.t290 156.095
R22783 VDD.t1875 VDD.t242 156.095
R22784 VDD.t68 VDD.t1815 154.417
R22785 VDD.t121 VDD.t2881 154.417
R22786 VDD.t2277 VDD.t2455 154.417
R22787 VDD.t2014 VDD.t2811 154.417
R22788 VDD.t2302 VDD.t2379 154.417
R22789 VDD.t2526 VDD.t2628 154.417
R22790 VDD.t2622 VDD.t2274 154.417
R22791 VDD.t636 VDD.t1362 154.417
R22792 VDD.t38 VDD.t820 154.417
R22793 VDD.t219 VDD.t1330 154.417
R22794 VDD.t2778 VDD.t2679 154.417
R22795 VDD.t1196 VDD.t2987 154.417
R22796 VDD.t2028 VDD.t1206 154.417
R22797 VDD.t199 VDD.t2016 154.417
R22798 VDD.t1274 VDD.t250 154.417
R22799 VDD.t2124 VDD.t1192 154.417
R22800 VDD.t2506 VDD.t2556 154.417
R22801 VDD.t920 VDD.t1887 154.417
R22802 VDD.t302 VDD.t74 154.417
R22803 VDD.t1902 VDD.t724 154.417
R22804 VDD.t632 VDD.t1886 154.417
R22805 VDD.t2780 VDD.t1070 154.417
R22806 VDD.t1070 VDD.t1216 154.417
R22807 VDD.t861 VDD.t1120 154.417
R22808 VDD.t704 VDD.t2159 154.417
R22809 VDD.t1465 VDD.t943 154.417
R22810 VDD.t960 VDD.t238 154.417
R22811 VDD.n1482 VDD.t2264 154.417
R22812 VDD.t1162 VDD.t2012 154.417
R22813 VDD.t1792 VDD.t234 154.417
R22814 VDD.t1160 VDD.t1342 154.417
R22815 VDD.n2058 VDD.t794 154.417
R22816 VDD.n2059 VDD.t2619 154.417
R22817 VDD.t1645 VDD.t710 154.417
R22818 VDD.t1939 VDD.t1041 154.417
R22819 VDD.t1638 VDD.t230 154.417
R22820 VDD.t242 VDD.t1932 154.417
R22821 VDD.t246 VDD.t1971 154.417
R22822 VDD.t1611 VDD.t1268 154.417
R22823 VDD.t90 VDD.t752 154.417
R22824 VDD.t1847 VDD.t1700 154.417
R22825 VDD.n355 VDD.n354 153.225
R22826 VDD.n385 VDD.n372 153.225
R22827 VDD.t153 VDD.t205 152.739
R22828 VDD.t2431 VDD.t298 152.739
R22829 VDD.t1460 VDD.t535 152.739
R22830 VDD.t2859 VDD.t1491 152.739
R22831 VDD.t1930 VDD.t322 152.739
R22832 VDD.t2839 VDD.t1759 151.06
R22833 VDD.t2640 VDD.t1920 151.06
R22834 VDD.t2691 VDD.t806 151.06
R22835 VDD.t651 VDD.n676 151.06
R22836 VDD.t84 VDD.t2467 149.382
R22837 VDD.t2406 VDD.t195 149.382
R22838 VDD.t544 VDD.t3006 149.382
R22839 VDD.t2728 VDD.t915 149.382
R22840 VDD.t953 VDD.t1262 149.382
R22841 VDD.n142 VDD.n106 149.249
R22842 VDD.t2828 VDD.t1685 147.703
R22843 VDD.t1420 VDD.t2036 147.703
R22844 VDD.t2879 VDD.t863 147.703
R22845 VDD.t1332 VDD.t2034 147.703
R22846 VDD.t617 VDD.t20 147.703
R22847 VDD.t537 VDD.t404 147.703
R22848 VDD.t865 VDD.t1794 147.703
R22849 VDD.t1445 VDD.t2239 147.703
R22850 VDD.t810 VDD.t1624 147.703
R22851 VDD.t1011 VDD.t1781 147.703
R22852 VDD.t1534 VDD.t1438 147.703
R22853 VDD.t603 VDD.t624 147.703
R22854 VDD.t1004 VDD.t256 147.703
R22855 VDD.t3085 VDD.t1985 147.703
R22856 VDD.t1150 VDD.t2032 147.703
R22857 VDD.t2979 VDD.t246 147.703
R22858 VDD.t258 VDD.t1983 147.703
R22859 VDD.t344 VDD.t2807 147.703
R22860 VDD.t3040 VDD.t1961 147.703
R22861 VDD.t2742 VDD.t66 147.703
R22862 VDD.n144 VDD.n143 147.328
R22863 VDD.t550 VDD.t2553 146.025
R22864 VDD.t1428 VDD.t2988 144.346
R22865 VDD.t984 VDD.t771 144.346
R22866 VDD.t771 VDD.t121 144.346
R22867 VDD.t1266 VDD.t1606 144.346
R22868 VDD.t2752 VDD.t2754 144.346
R22869 VDD.t2754 VDD.t2748 144.346
R22870 VDD.t1376 VDD.t2133 144.346
R22871 VDD.t996 VDD.t998 144.346
R22872 VDD.t998 VDD.t994 144.346
R22873 VDD.t1144 VDD.t1142 144.346
R22874 VDD.t1142 VDD.t1146 144.346
R22875 VDD.t1146 VDD.t1148 144.346
R22876 VDD.t1171 VDD.t1169 144.346
R22877 VDD.t1863 VDD.t1861 144.346
R22878 VDD.t1859 VDD.t1863 144.346
R22879 VDD.t1865 VDD.t1859 144.346
R22880 VDD.t2001 VDD.t2005 144.346
R22881 VDD.t2005 VDD.t2003 144.346
R22882 VDD.t2003 VDD.t1999 144.346
R22883 VDD.t1951 VDD.t1953 144.346
R22884 VDD.t1953 VDD.t1949 144.346
R22885 VDD.t1949 VDD.t1947 144.346
R22886 VDD.t1314 VDD.t1308 144.346
R22887 VDD.t1487 VDD.t2672 144.346
R22888 VDD.t2680 VDD.t687 144.346
R22889 VDD.t1577 VDD.t1074 144.346
R22890 VDD.t1681 VDD.t497 144.346
R22891 VDD.t1997 VDD.t1675 144.346
R22892 VDD.t501 VDD.t613 144.346
R22893 VDD.t141 VDD.t137 144.346
R22894 VDD.t135 VDD.t141 144.346
R22895 VDD.t1071 VDD.t1885 144.346
R22896 VDD.t862 VDD.t1880 144.346
R22897 VDD.n1483 VDD.t2740 144.346
R22898 VDD.t1533 VDD.t950 144.346
R22899 VDD.t1161 VDD.t948 144.346
R22900 VDD.t2786 VDD.t2790 144.346
R22901 VDD.t1334 VDD.t505 144.346
R22902 VDD.t505 VDD.t494 144.346
R22903 VDD.t2985 VDD.t2986 144.346
R22904 VDD.t2986 VDD.t589 144.346
R22905 VDD.t589 VDD.t610 144.346
R22906 VDD.t813 VDD.t1098 144.346
R22907 VDD.t1095 VDD.t482 144.346
R22908 VDD.t1610 VDD.t2072 144.346
R22909 VDD.t929 VDD.t925 144.346
R22910 VDD.n2928 VDD.t2884 143.06
R22911 VDD.t1895 VDD.t1428 142.668
R22912 VDD.t2750 VDD.t2376 142.668
R22913 VDD.t3061 VDD.t1312 142.668
R22914 VDD.t1039 VDD.t2669 142.668
R22915 VDD.t419 VDD.t320 142.668
R22916 VDD.t2853 VDD.t1385 142.668
R22917 VDD.t1578 VDD.t1937 142.668
R22918 VDD.t1835 VDD.t835 142.668
R22919 VDD.t139 VDD.t2397 142.668
R22920 VDD.t53 VDD.t499 142.668
R22921 VDD.t933 VDD.t2788 142.668
R22922 VDD.t619 VDD.t927 142.668
R22923 VDD.t1138 VDD.t1136 140.989
R22924 VDD.t1689 VDD.t1687 140.989
R22925 VDD.t970 VDD.t968 140.989
R22926 VDD.t1036 VDD.t1034 140.989
R22927 VDD.t1111 VDD.t683 140.989
R22928 VDD.t1606 VDD.t701 140.989
R22929 VDD.t1665 VDD.t1058 140.989
R22930 VDD.t398 VDD.t587 140.989
R22931 VDD.t717 VDD.t46 140.989
R22932 VDD.t46 VDD.t1743 140.989
R22933 VDD.t26 VDD.t2135 140.989
R22934 VDD.t2080 VDD.t1967 140.989
R22935 VDD.t1189 VDD.t1187 140.989
R22936 VDD.t1551 VDD.t1549 140.989
R22937 VDD.t2110 VDD.t2108 140.989
R22938 VDD.t2020 VDD.t2018 140.989
R22939 VDD.t1515 VDD.t1517 140.989
R22940 VDD.t2098 VDD.t2100 140.989
R22941 VDD.t2185 VDD.t2187 140.989
R22942 VDD.t2191 VDD.t2189 140.989
R22943 VDD.t3071 VDD.t2041 140.989
R22944 VDD.t321 VDD.t3071 140.989
R22945 VDD.t1955 VDD.t1957 140.989
R22946 VDD.t1086 VDD.t1084 140.989
R22947 VDD.t975 VDD.t385 140.989
R22948 VDD.t891 VDD.t893 140.989
R22949 VDD.t2772 VDD.t2774 140.989
R22950 VDD.t661 VDD.t663 140.989
R22951 VDD.t1173 VDD.t1175 140.989
R22952 VDD.t2744 VDD.t2746 140.989
R22953 VDD.t1855 VDD.t1857 140.989
R22954 VDD.t1029 VDD.t983 140.989
R22955 VDD.t983 VDD.t2707 140.989
R22956 VDD.t2063 VDD.t2065 140.989
R22957 VDD.t1362 VDD.t1797 140.989
R22958 VDD.t742 VDD.t282 140.989
R22959 VDD.t573 VDD.t1513 140.989
R22960 VDD.t1081 VDD.t38 140.989
R22961 VDD.t548 VDD.t396 140.989
R22962 VDD.t402 VDD.t406 140.989
R22963 VDD.t266 VDD.t1635 140.989
R22964 VDD.t1635 VDD.t949 140.989
R22965 VDD.t225 VDD.t13 140.989
R22966 VDD.t547 VDD.t1460 140.989
R22967 VDD.t3006 VDD.t1788 140.989
R22968 VDD.t395 VDD.t1482 140.989
R22969 VDD.t1459 VDD.t554 140.989
R22970 VDD.t333 VDD.t3025 140.989
R22971 VDD.t2157 VDD.t2155 140.989
R22972 VDD.t867 VDD.t789 140.989
R22973 VDD.t789 VDD.t131 140.989
R22974 VDD.t1015 VDD.t1487 140.989
R22975 VDD.t2670 VDD.t30 140.989
R22976 VDD.t1249 VDD.t1247 140.989
R22977 VDD.t1751 VDD.t1753 140.989
R22978 VDD.t1753 VDD.t1757 140.989
R22979 VDD.t1618 VDD.t364 140.989
R22980 VDD.t2683 VDD.t2925 140.989
R22981 VDD.t354 VDD.t688 140.989
R22982 VDD.t854 VDD.t1622 140.989
R22983 VDD.t189 VDD.t854 140.989
R22984 VDD.t1074 VDD.t1066 140.989
R22985 VDD.t1451 VDD.t1453 140.989
R22986 VDD.t1597 VDD.t1595 140.989
R22987 VDD.t1286 VDD.t1284 140.989
R22988 VDD.t274 VDD.t272 140.989
R22989 VDD.t814 VDD.t816 140.989
R22990 VDD.t467 VDD.t471 140.989
R22991 VDD.t3063 VDD.t3065 140.989
R22992 VDD.t590 VDD.t600 140.989
R22993 VDD.t2709 VDD.t2704 140.989
R22994 VDD.t1975 VDD.t1977 140.989
R22995 VDD.t1811 VDD.t1807 140.989
R22996 VDD.t2007 VDD.t1987 140.989
R22997 VDD.t1987 VDD.t3102 140.989
R22998 VDD.t1701 VDD.t1703 140.989
R22999 VDD.t2083 VDD.t2085 140.989
R23000 VDD.t2826 VDD.t2815 140.989
R23001 VDD.t2815 VDD.t1740 140.989
R23002 VDD.t1740 VDD.t1745 140.989
R23003 VDD.t2 VDD.t15 140.989
R23004 VDD.t15 VDD.t2947 140.989
R23005 VDD.t1010 VDD.t2943 140.989
R23006 VDD.t3017 VDD.t3020 140.989
R23007 VDD.t3020 VDD.t160 140.989
R23008 VDD.t532 VDD.t164 140.989
R23009 VDD.t2231 VDD.t1528 140.989
R23010 VDD.t2128 VDD.t2126 140.989
R23011 VDD.t2196 VDD.t1547 140.989
R23012 VDD.t1786 VDD.t1771 140.989
R23013 VDD.t250 VDD.t248 140.989
R23014 VDD.t2114 VDD.t350 140.989
R23015 VDD.t2911 VDD.t423 140.989
R23016 VDD.t2855 VDD.t2895 140.989
R23017 VDD.t1626 VDD.t389 140.989
R23018 VDD.t267 VDD.t413 140.989
R23019 VDD.t72 VDD.t70 140.989
R23020 VDD.t278 VDD.t280 140.989
R23021 VDD.t2870 VDD.t2873 140.989
R23022 VDD.t673 VDD.t671 140.989
R23023 VDD.t1301 VDD.t1303 140.989
R23024 VDD.t1060 VDD.t1062 140.989
R23025 VDD.t2951 VDD.t2954 140.989
R23026 VDD.t109 VDD.t111 140.989
R23027 VDD.t310 VDD.t308 140.989
R23028 VDD.t2650 VDD.t2648 140.989
R23029 VDD.t1823 VDD.t1821 140.989
R23030 VDD.t1571 VDD.t1567 140.989
R23031 VDD.t2782 VDD.t569 140.989
R23032 VDD.t1072 VDD.t78 140.989
R23033 VDD.t1825 VDD.t2781 140.989
R23034 VDD.t630 VDD.t1358 140.989
R23035 VDD.t1883 VDD.t1364 140.989
R23036 VDD.t2965 VDD.t3097 140.989
R23037 VDD.t3097 VDD.t3100 140.989
R23038 VDD.t1202 VDD.t1200 140.989
R23039 VDD.t2960 VDD.t1197 140.989
R23040 VDD.t1650 VDD.t1648 140.989
R23041 VDD.t1242 VDD.t1466 140.989
R23042 VDD.t1614 VDD.t24 140.989
R23043 VDD.t424 VDD.t12 140.989
R23044 VDD.t507 VDD.t513 140.989
R23045 VDD.t1721 VDD.t1723 140.989
R23046 VDD.t2667 VDD.t2665 140.989
R23047 VDD.t40 VDD.t2734 140.989
R23048 VDD.t509 VDD.t415 140.989
R23049 VDD.t903 VDD.t1533 140.989
R23050 VDD.t951 VDD.t203 140.989
R23051 VDD.t1163 VDD.t2206 140.989
R23052 VDD.t1655 VDD.t1161 140.989
R23053 VDD.t918 VDD.t1354 140.989
R23054 VDD.t946 VDD.t201 140.989
R23055 VDD.t430 VDD.t2830 140.989
R23056 VDD.t1093 VDD.t1091 140.989
R23057 VDD.t1633 VDD.t1629 140.989
R23058 VDD.t1557 VDD.t1559 140.989
R23059 VDD.t2861 VDD.t796 140.989
R23060 VDD.t127 VDD.t129 140.989
R23061 VDD.t262 VDD.t260 140.989
R23062 VDD.t3027 VDD.t3029 140.989
R23063 VDD.t733 VDD.t735 140.989
R23064 VDD.t881 VDD.t879 140.989
R23065 VDD.t2865 VDD.t2868 140.989
R23066 VDD.t667 VDD.t665 140.989
R23067 VDD.t1477 VDD.t1479 140.989
R23068 VDD.t1965 VDD.t1963 140.989
R23069 VDD.t1891 VDD.t1889 140.989
R23070 VDD.t2697 VDD.t2699 140.989
R23071 VDD.t1032 VDD.t1030 140.989
R23072 VDD.t2224 VDD.t2222 140.989
R23073 VDD.t480 VDD.t475 140.989
R23074 VDD.t304 VDD.t1695 140.989
R23075 VDD.t3008 VDD.t1733 140.989
R23076 VDD.t1910 VDD.t1912 140.989
R23077 VDD.t1912 VDD.t1904 140.989
R23078 VDD.t847 VDD.t845 140.989
R23079 VDD.t1368 VDD.t1366 140.989
R23080 VDD.t2799 VDD.t2801 140.989
R23081 VDD.t1183 VDD.t1179 140.989
R23082 VDD.t1179 VDD.t1185 140.989
R23083 VDD.t781 VDD.t296 140.989
R23084 VDD.t1096 VDD.t34 140.989
R23085 VDD.t1107 VDD.t1103 140.989
R23086 VDD.t1105 VDD.t1101 140.989
R23087 VDD.t2145 VDD.t32 140.989
R23088 VDD.t432 VDD.t227 140.989
R23089 VDD.t2232 VDD.t2234 140.989
R23090 VDD.t3019 VDD.t426 140.989
R23091 VDD.t839 VDD.t841 140.989
R23092 VDD.t2169 VDD.t2175 140.989
R23093 VDD.t2175 VDD.t2177 140.989
R23094 VDD.t2177 VDD.t2173 140.989
R23095 VDD.t2183 VDD.t175 140.989
R23096 VDD.t2070 VDD.t358 140.989
R23097 VDD.t335 VDD.t429 140.989
R23098 VDD.t340 VDD.t2889 140.989
R23099 VDD.t433 VDD.t94 140.989
R23100 VDD.t1254 VDD.t1256 140.989
R23101 VDD.t1631 VDD.t1133 140.989
R23102 VDD.t2008 VDD.t2010 140.989
R23103 VDD.t540 VDD.t542 140.989
R23104 VDD.t2660 VDD.t2658 140.989
R23105 VDD.t605 VDD.t607 140.989
R23106 VDD.t2165 VDD.t2163 140.989
R23107 VDD.t769 VDD.t767 140.989
R23108 VDD.t697 VDD.t699 140.989
R23109 VDD.t2138 VDD.t2140 140.989
R23110 VDD.t2087 VDD.t1537 140.989
R23111 VDD.t64 VDD.t1802 140.989
R23112 VDD.t2760 VDD.t2758 140.989
R23113 VDD.t2758 VDD.t2756 140.989
R23114 VDD.t3050 VDD.t3042 140.989
R23115 VDD.t3042 VDD.t3048 140.989
R23116 VDD.t3054 VDD.t3044 140.989
R23117 VDD.t3046 VDD.t3054 140.989
R23118 VDD.t2718 VDD.t2722 140.989
R23119 VDD.t2724 VDD.t2718 140.989
R23120 VDD.n199 VDD.n196 140.702
R23121 VDD.n199 VDD.n195 140.048
R23122 VDD.t3059 VDD.t1767 139.311
R23123 VDD.t1969 VDD.t1000 139.311
R23124 VDD.t564 VDD.t1344 139.311
R23125 VDD.t1488 VDD.t2220 139.311
R23126 VDD.t977 VDD.t1075 139.311
R23127 VDD.t2149 VDD.t383 139.311
R23128 VDD.t1679 VDD.t2093 139.311
R23129 VDD.t488 VDD.t1204 139.311
R23130 VDD.t2688 VDD.t1524 139.311
R23131 VDD.t1943 VDD.t3072 139.311
R23132 VDD.t1455 VDD.t372 139.311
R23133 VDD.t1360 VDD.t2958 139.311
R23134 VDD.t1873 VDD.t209 139.311
R23135 VDD.t1869 VDD.t746 137.633
R23136 VDD.t2714 VDD.t659 137.633
R23137 VDD.t1878 VDD.t708 137.633
R23138 VDD.t1371 VDD.t2803 137.633
R23139 VDD.t492 VDD.t1002 135.954
R23140 VDD.t2817 VDD.t2482 135.954
R23141 VDD.t600 VDD.t2587 135.954
R23142 VDD.t119 VDD.t329 135.954
R23143 VDD.t2694 VDD.t2532 135.954
R23144 VDD.t2317 VDD.t2142 135.954
R23145 VDD.t400 VDD.t28 134.276
R23146 VDD.t2821 VDD.t408 134.276
R23147 VDD.t2236 VDD.t1208 134.276
R23148 VDD.t1773 VDD.t1914 134.276
R23149 VDD.t236 VDD.t2654 134.276
R23150 VDD.n461 VDD.t3137 133.512
R23151 VDD.n4356 VDD.n4312 133.382
R23152 VDD.t571 VDD.t1489 132.597
R23153 VDD.n3422 VDD.t1828 132.597
R23154 VDD.t1258 VDD.t2901 132.597
R23155 VDD.t913 VDD.t2914 132.597
R23156 VDD.t2973 VDD.t2887 132.597
R23157 VDD.t1677 VDD.t82 132.597
R23158 VDD.t1194 VDD.t862 132.597
R23159 VDD.t1120 VDD.t592 132.597
R23160 VDD.t943 VDD.t960 132.597
R23161 VDD.t2012 VDD.t1792 132.597
R23162 VDD.t1342 VDD.t1131 132.597
R23163 VDD.t338 VDD.t2059 132.597
R23164 VDD.t331 VDD.t362 132.597
R23165 VDD.t1041 VDD.t1638 132.597
R23166 VDD.n613 VDD.t1610 132.597
R23167 VDD.t1268 VDD.t477 132.597
R23168 VDD.t1961 VDD.t1847 132.597
R23169 VDD.n319 VDD.t453 132.355
R23170 VDD.n269 VDD.n250 131.388
R23171 VDD.n263 VDD.n250 131.388
R23172 VDD.t640 VDD.t553 130.919
R23173 VDD.t2345 VDD.t2185 130.919
R23174 VDD.t1621 VDD.t1396 130.919
R23175 VDD.t1575 VDD.t633 130.919
R23176 VDD.n4357 VDD.t3147 129.344
R23177 VDD.n3694 VDD.t3164 129.344
R23178 VDD.n4220 VDD.t3134 129.344
R23179 VDD.n4072 VDD.t3141 129.344
R23180 VDD.n3957 VDD.t3237 129.344
R23181 VDD.n3037 VDD.t3230 129.344
R23182 VDD.n2649 VDD.t3181 129.344
R23183 VDD.n621 VDD.t3183 129.344
R23184 VDD.n669 VDD.t3152 129.344
R23185 VDD.n1018 VDD.t3234 129.344
R23186 VDD.n721 VDD.t3176 129.344
R23187 VDD.n913 VDD.t3178 129.344
R23188 VDD.t915 VDD.t596 129.24
R23189 VDD.t417 VDD.t2202 129.24
R23190 VDD.n635 VDD.t3196 128.489
R23191 VDD.n4238 VDD.t3193 127.883
R23192 VDD.n659 VDD.t3146 127.883
R23193 VDD.n4250 VDD.t2693 127.562
R23194 VDD.t2089 VDD.t1310 127.562
R23195 VDD.t785 VDD.t2949 127.562
R23196 VDD.t786 VDD.t158 127.562
R23197 VDD.t1569 VDD.t1817 127.562
R23198 VDD.t1573 VDD.t1819 127.562
R23199 VDD.t217 VDD.t2662 127.562
R23200 VDD.t211 VDD.t511 127.562
R23201 VDD.t948 VDD.t860 127.562
R23202 VDD.t1382 VDD.t2784 127.562
R23203 VDD.n723 VDD.t1294 127.562
R23204 VDD.t889 VDD.t931 127.562
R23205 VDD.t826 VDD.t3052 127.562
R23206 VDD.t1316 VDD.t3056 127.562
R23207 VDD.t453 VDD.t440 127.291
R23208 VDD.t440 VDD.t442 127.291
R23209 VDD.t442 VDD.t438 127.291
R23210 VDD.t438 VDD.t460 127.291
R23211 VDD.t460 VDD.t448 127.291
R23212 VDD.t434 VDD.t448 127.291
R23213 VDD.t444 VDD.t434 127.291
R23214 VDD.t458 VDD.t444 127.291
R23215 VDD.t436 VDD.t458 127.291
R23216 VDD.t446 VDD.t456 127.291
R23217 VDD.t450 VDD.t446 127.291
R23218 VDD.n1122 VDD.t3180 125.989
R23219 VDD.t2047 VDD.t1346 125.883
R23220 VDD.t808 VDD.t22 125.883
R23221 VDD.t1134 VDD.t1282 125.883
R23222 VDD.t356 VDD.t1234 125.883
R23223 VDD.t1006 VDD.t348 125.883
R23224 VDD.t2096 VDD.t649 125.883
R23225 VDD.t2764 VDD.n380 124.206
R23226 VDD.t2770 VDD.n379 124.206
R23227 VDD.t2768 VDD.n382 124.206
R23228 VDD.t2766 VDD.n381 124.206
R23229 VDD.t2881 VDD.t1420 124.206
R23230 VDD.t1372 VDD.t1928 124.206
R23231 VDD.t375 VDD.t2875 124.206
R23232 VDD.t170 VDD.t1198 124.206
R23233 VDD.n3698 VDD.t2844 123.507
R23234 VDD.n4324 VDD.t1403 123.507
R23235 VDD.n2943 VDD.t2850 123.507
R23236 VDD.n3365 VDD.t1494 123.507
R23237 VDD.n2986 VDD.t1584 123.507
R23238 VDD.n2206 VDD.t2834 123.507
R23239 VDD.n1534 VDD.t776 123.507
R23240 VDD.n2916 VDD.t2838 123.507
R23241 VDD.n2969 VDD.t2678 123.507
R23242 VDD.n3525 VDD.t2852 123.507
R23243 VDD.n2176 VDD.t963 123.507
R23244 VDD.n2250 VDD.t2832 123.507
R23245 VDD.n2265 VDD.t680 123.507
R23246 VDD.n2296 VDD.t695 123.507
R23247 VDD.n1267 VDD.t1007 123.507
R23248 VDD.n671 VDD.t650 123.507
R23249 VDD.t2134 VDD.t1923 122.526
R23250 VDD.t1440 VDD.t993 122.526
R23251 VDD.n2263 VDD.t1543 122.526
R23252 VDD.t2736 VDD.t911 122.526
R23253 VDD.t1904 VDD.t847 122.526
R23254 VDD.t3035 VDD.n346 122.034
R23255 VDD.n390 VDD.t58 122.034
R23256 VDD.t61 VDD.n346 122.034
R23257 VDD.t464 VDD.n390 122.034
R23258 VDD.t3035 VDD.n339 122.034
R23259 VDD.t464 VDD.n339 122.034
R23260 VDD.t1809 VDD.t1296 120.849
R23261 VDD.t1683 VDD.t2706 120.849
R23262 VDD.t323 VDD.t1526 120.849
R23263 VDD.t326 VDD.t1300 120.849
R23264 VDD.t1434 VDD.t1220 120.849
R23265 VDD.t168 VDD.t1827 120.849
R23266 VDD.t1996 VDD.t1099 120.849
R23267 VDD.t628 VDD.t1742 120.849
R23268 VDD.t2856 VDD.t2883 120.849
R23269 VDD.t1125 VDD.t2942 120.849
R23270 VDD.t166 VDD.t712 120.849
R23271 VDD.t1671 VDD.t496 120.849
R23272 VDD.t1813 VDD.t1293 120.849
R23273 VDD.t1117 VDD.t167 120.849
R23274 VDD.t2230 VDD.t2690 120.849
R23275 VDD.t1505 VDD.t1652 120.849
R23276 VDD.t324 VDD.t1156 120.849
R23277 VDD.t330 VDD.t1834 120.849
R23278 VDD.t691 VDD.t171 120.849
R23279 VDD.t1307 VDD.t779 120.849
R23280 VDD.t322 VDD.t737 120.849
R23281 VDD.t764 VDD.t832 120.849
R23282 VDD.t485 VDD.t611 120.849
R23283 VDD.t474 VDD.t2819 120.849
R23284 VDD.t986 VDD.t1437 120.849
R23285 VDD.t486 VDD.t3010 120.849
R23286 VDD.t484 VDD.t1442 120.849
R23287 VDD.t466 VDD.t1783 120.849
R23288 VDD.t2173 VDD.t258 120.849
R23289 VDD.t477 VDD.t2891 120.849
R23290 VDD.t346 VDD.t479 120.849
R23291 VDD.t95 VDD.t478 120.849
R23292 VDD.t754 VDD.t193 120.849
R23293 VDD.n3798 VDD.t3110 119.624
R23294 VDD.n3734 VDD.t1968 119.608
R23295 VDD.n3502 VDD.t1386 119.608
R23296 VDD.n2942 VDD.t1756 119.608
R23297 VDD.n2956 VDD.t940 119.608
R23298 VDD.n3357 VDD.t1329 119.608
R23299 VDD.n2980 VDD.t1016 119.608
R23300 VDD.n2983 VDD.t868 119.608
R23301 VDD.n3529 VDD.t1623 119.608
R23302 VDD.n3532 VDD.t1067 119.608
R23303 VDD.n3159 VDD.t635 119.608
R23304 VDD.n3180 VDD.t819 119.608
R23305 VDD.n2244 VDD.t1273 119.608
R23306 VDD.n2264 VDD.t2197 119.608
R23307 VDD.n1389 VDD.t1564 119.608
R23308 VDD.n1422 VDD.t1415 119.608
R23309 VDD.n1445 VDD.t1656 119.608
R23310 VDD.n1468 VDD.t904 119.608
R23311 VDD.n1471 VDD.t1225 119.608
R23312 VDD.n1513 VDD.t1243 119.608
R23313 VDD.n1702 VDD.t1826 119.608
R23314 VDD.n1565 VDD.t1576 119.608
R23315 VDD.n1759 VDD.t1498 119.608
R23316 VDD.n1016 VDD.t1178 119.608
R23317 VDD.n547 VDD.t751 119.608
R23318 VDD.n614 VDD.t2172 119.608
R23319 VDD.n693 VDD.t1110 119.608
R23320 VDD.n737 VDD.t1909 119.608
R23321 VDD.t1374 VDD.t2079 119.171
R23322 VDD.t1604 VDD.t115 119.171
R23323 VDD.t1871 VDD.t2075 119.171
R23324 VDD.t775 VDD.t2102 119.171
R23325 VDD.t292 VDD.t2961 119.171
R23326 VDD.t1049 VDD.t909 119.171
R23327 VDD.t1224 VDD.t907 119.171
R23328 VDD.n2113 VDD.t3240 119.007
R23329 VDD.n3791 VDD.t3241 118.919
R23330 VDD.n2226 VDD.t3117 118.919
R23331 VDD.n628 VDD.t3224 118.919
R23332 VDD.n4181 VDD.t3156 118.853
R23333 VDD.n3877 VDD.t3208 118.853
R23334 VDD.n3918 VDD.t3115 118.853
R23335 VDD.n2369 VDD.t3186 118.853
R23336 VDD.t602 VDD.t2976 118.267
R23337 VDD.t3039 VDD.t144 118.267
R23338 VDD.t1853 VDD.t36 117.492
R23339 VDD.t92 VDD.t1563 117.492
R23340 VDD.t103 VDD.t884 117.492
R23341 VDD.n2326 VDD.t597 117.451
R23342 VDD.n1479 VDD.t2900 117.451
R23343 VDD.n1522 VDD.t214 117.451
R23344 VDD.n2850 VDD.n2223 117.334
R23345 VDD.n4030 VDD.t3222 117.294
R23346 VDD.n1923 VDD.t3148 117.294
R23347 VDD.n1624 VDD.t3109 117.294
R23348 VDD.n817 VDD.t3242 117.294
R23349 VDD.t2976 VDD.t172 116.82
R23350 VDD.t172 VDD.t412 116.82
R23351 VDD.t412 VDD.t3070 116.82
R23352 VDD.t3070 VDD.t2975 116.82
R23353 VDD.t2975 VDD.t143 116.82
R23354 VDD.t3087 VDD.t157 116.82
R23355 VDD.t3058 VDD.t3087 116.82
R23356 VDD.t2040 VDD.t3058 116.82
R23357 VDD.t3078 VDD.t2040 116.82
R23358 VDD.t144 VDD.t3078 116.82
R23359 VDD.n3710 VDD.t388 116.341
R23360 VDD.n4102 VDD.t422 116.341
R23361 VDD.n3665 VDD.t386 116.341
R23362 VDD.n2179 VDD.t390 116.341
R23363 VDD.n2097 VDD.t414 116.341
R23364 VDD.n2260 VDD.t418 116.341
R23365 VDD.n2293 VDD.t1292 116.341
R23366 VDD.n2051 VDD.t317 116.341
R23367 VDD.n1486 VDD.t416 116.341
R23368 VDD.n1545 VDD.t491 116.341
R23369 VDD.n758 VDD.t1694 116.341
R23370 VDD.n770 VDD.t305 116.341
R23371 VDD.t1762 VDD.t2861 115.814
R23372 VDD.n263 VDD.n262 115.201
R23373 VDD.n264 VDD.n263 115.201
R23374 VDD.n121 VDD.n120 115.201
R23375 VDD.n2107 VDD.t3118 114.912
R23376 VDD.n2406 VDD.t3187 114.546
R23377 VDD.t2969 VDD.t585 114.135
R23378 VDD.t758 VDD.t850 114.135
R23379 VDD.t1181 VDD.t1830 114.135
R23380 VDD.t387 VDD.t1165 112.457
R23381 VDD.t1544 VDD.t2831 112.457
R23382 VDD.t2206 VDD.t2541 112.457
R23383 VDD.t2234 VDD.t563 112.457
R23384 VDD.t2072 VDD.t3079 112.457
R23385 VDD.n1275 VDD.t3229 112.117
R23386 VDD.n2598 VDD.t3197 111.537
R23387 VDD.t122 VDD.t1877 110.778
R23388 VDD.t2882 VDD.t1665 110.778
R23389 VDD.t1549 VDD.t2693 110.778
R23390 VDD.t2711 VDD.t2157 110.778
R23391 VDD.t2837 VDD.t2923 110.778
R23392 VDD.t688 VDD.t166 110.778
R23393 VDD.n132 VDD.t2792 110.394
R23394 VDD.t2241 VDD.n215 110.284
R23395 VDD.n989 VDD.t1295 110.227
R23396 VDD.t162 VDD.t1167 109.1
R23397 VDD.t1356 VDD.t1348 109.1
R23398 VDD.t1246 VDD.t837 109.1
R23399 VDD.t1471 VDD.t1505 109.1
R23400 VDD.t2212 VDD.t1653 109.1
R23401 VDD.t1779 VDD.t2116 109.1
R23402 VDD.t1466 VDD.t431 109.1
R23403 VDD.t2490 VDD.t2494 108.832
R23404 VDD.t2452 VDD.t2580 108.832
R23405 VDD.t2286 VDD.t2372 108.832
R23406 VDD.t2267 VDD.t2646 108.832
R23407 VDD.n129 VDD.n128 108.8
R23408 VDD.n127 VDD.n120 108.8
R23409 VDD.t1565 VDD.t421 107.421
R23410 VDD.t2706 VDD.t1551 107.421
R23411 VDD.t2155 VDD.t558 107.421
R23412 VDD.t1828 VDD.t427 107.421
R23413 VDD.t1620 VDD.t1777 107.421
R23414 VDD.t974 VDD.t354 107.421
R23415 VDD.t763 VDD.t515 107.421
R23416 VDD.t1185 VDD.t3037 107.421
R23417 VDD.n4442 VDD.n4364 106.561
R23418 VDD.n874 VDD.n873 106.561
R23419 VDD.n4252 VDD.n4251 106.559
R23420 VDD.n3837 VDD.n3727 106.559
R23421 VDD.n3839 VDD.n3771 106.559
R23422 VDD.n3841 VDD.n3814 106.559
R23423 VDD.n1230 VDD.n1229 106.559
R23424 VDD.n1143 VDD.n645 106.559
R23425 VDD.n1049 VDD.n701 106.559
R23426 VDD.n875 VDD.n744 106.559
R23427 VDD.t1829 VDD.t1532 105.743
R23428 VDD.t2045 VDD.t714 105.743
R23429 VDD.t244 VDD.t1272 105.743
R23430 VDD.t1769 VDD.t2125 105.743
R23431 VDD.t1613 VDD.t2823 105.743
R23432 VDD.t2147 VDD.t1507 105.743
R23433 VDD.t1437 VDD.t2232 105.743
R23434 VDD.t2189 VDD.n4363 104.064
R23435 VDD.t385 VDD.t2616 104.064
R23436 VDD.t1652 VDD.t2194 104.064
R23437 VDD.t213 VDD.t1238 104.064
R23438 VDD.t2899 VDD.t1663 104.064
R23439 VDD.t1414 VDD.t621 104.064
R23440 VDD.t1159 VDD.t1088 104.064
R23441 VDD.n432 VDD.n412 103.906
R23442 VDD.t1900 VDD.t1013 102.385
R23443 VDD.t2679 VDD.n3573 102.385
R23444 VDD.t1068 VDD.t2153 102.385
R23445 VDD.t1616 VDD.t51 102.385
R23446 VDD.t828 VDD.t2712 102.385
R23447 VDD.t47 VDD.t1581 102.385
R23448 VDD.t856 VDD.t918 102.385
R23449 VDD.t2575 VDD.t1160 102.385
R23450 VDD.t1700 VDD.t2308 102.385
R23451 VDD.n2284 VDD.t534 101.733
R23452 VDD.n2321 VDD.t1012 101.733
R23453 VDD.n2331 VDD.t45 101.733
R23454 VDD.n2502 VDD.t982 101.733
R23455 VDD.n1356 VDD.t1763 101.733
R23456 VDD.n1410 VDD.t1132 101.733
R23457 VDD.n1428 VDD.t1090 101.733
R23458 VDD.n1499 VDD.t2664 101.733
R23459 VDD.n1738 VDD.t1989 101.733
R23460 VDD.t555 VDD.t393 100.707
R23461 VDD.t133 VDD.t1934 100.707
R23462 VDD.t2214 VDD.t1249 100.707
R23463 VDD.t2193 VDD.t2907 100.707
R23464 VDD.t1416 VDD.t2960 100.707
R23465 VDD.t4 VDD.t1236 100.707
R23466 VDD.t1244 VDD.t2956 100.707
R23467 VDD.t2893 VDD.t1657 100.707
R23468 VDD.t1661 VDD.t3014 100.707
R23469 VDD.t2061 VDD.t1394 100.707
R23470 VDD.t1116 VDD.t1557 100.707
R23471 VDD.t966 VDD.t718 100.707
R23472 VDD.t2835 VDD.t1548 99.0288
R23473 VDD.t1152 VDD.t1093 99.0288
R23474 VDD.t97 VDD.t1555 99.0288
R23475 VDD.t1449 VDD.t1008 99.0288
R23476 VDD.t812 VDD.t8 99.0288
R23477 VDD.n4047 VDD.t1744 98.5005
R23478 VDD.n3394 VDD.t328 98.5005
R23479 VDD.n3246 VDD.t2818 98.5005
R23480 VDD.n3010 VDD.t1674 98.5005
R23481 VDD.n3014 VDD.t29 98.5005
R23482 VDD.n3036 VDD.t2708 98.5005
R23483 VDD.n2205 VDD.t337 98.5005
R23484 VDD.n2212 VDD.t2974 98.5005
R23485 VDD.n2270 VDD.t1525 98.5005
R23486 VDD.n2731 VDD.t1529 98.5005
R23487 VDD.n2278 VDD.t165 98.5005
R23488 VDD.n2290 VDD.t224 98.5005
R23489 VDD.n2658 VDD.t11 98.5005
R23490 VDD.n2315 VDD.t2944 98.5005
R23491 VDD.n2366 VDD.t3103 98.5005
R23492 VDD.n1353 VDD.t98 98.5005
R23493 VDD.n1419 VDD.t1395 98.5005
R23494 VDD.n1440 VDD.t1355 98.5005
R23495 VDD.n1494 VDD.t512 98.5005
R23496 VDD.n1788 VDD.t2959 98.5005
R23497 VDD.n534 VDD.t1632 98.5005
R23498 VDD.t1925 VDD.t1463 97.3503
R23499 VDD.t1493 VDD.t1213 97.3503
R23500 VDD.t777 VDD.t2921 97.3503
R23501 VDD.t954 VDD.t2610 97.3503
R23502 VDD.t1053 VDD.t2081 97.3503
R23503 VDD.t642 VDD.t1474 97.2286
R23504 VDD.t2792 VDD.t2685 97.2286
R23505 VDD.n4052 VDD.t2812 96.1553
R23506 VDD.n3776 VDD.t410 96.1553
R23507 VDD.n3779 VDD.t864 96.1553
R23508 VDD.n2959 VDD.t1353 96.1553
R23509 VDD.n3144 VDD.t595 96.1553
R23510 VDD.n2271 VDD.t2689 96.1553
R23511 VDD.n2277 VDD.t3024 96.1553
R23512 VDD.n2314 VDD.t7 96.1553
R23513 VDD.n2361 VDD.t1676 96.1553
R23514 VDD.n2362 VDD.t1998 96.1553
R23515 VDD.n2365 VDD.t2972 96.1553
R23516 VDD.n2385 VDD.t498 96.1553
R23517 VDD.n2386 VDD.t1682 96.1553
R23518 VDD.n1416 VDD.t2898 96.1553
R23519 VDD.n1438 VDD.t2023 96.1553
R23520 VDD.n1460 VDD.t1439 96.1553
R23521 VDD.n1491 VDD.t222 96.1553
R23522 VDD.n546 VDD.t755 96.1553
R23523 VDD.n543 VDD.t91 96.1553
R23524 VDD.n537 VDD.t345 96.1553
R23525 VDD.n347 VDD.n346 95.9736
R23526 VDD.n390 VDD.n389 95.9736
R23527 VDD.t143 VDD.n72 95.7389
R23528 VDD.t157 VDD.n35 95.7389
R23529 VDD.t1083 VDD.t1799 95.6719
R23530 VDD.t1080 VDD.t1796 95.6719
R23531 VDD.t1673 VDD.t1436 95.6719
R23532 VDD.t2026 VDD.t937 95.6719
R23533 VDD.t1017 VDD.t1749 95.6719
R23534 VDD.t2958 VDD.n1555 95.6719
R23535 VDD.t1535 VDD.t1222 95.6719
R23536 VDD.t1410 VDD.t173 95.6719
R23537 VDD.t1412 VDD.t1390 95.6719
R23538 VDD.t1406 VDD.t1392 95.6719
R23539 VDD.t1324 VDD.t843 95.6719
R23540 VDD.t1839 VDD.t1589 95.6719
R23541 VDD.t1849 VDD.t2167 95.6719
R23542 VDD.n203 VDD.n196 95.0755
R23543 VDD.t3093 VDD.t685 93.9934
R23544 VDD.t919 VDD.t939 93.9934
R23545 VDD.t1509 VDD.t2120 93.9934
R23546 VDD.t556 VDD.t852 93.9934
R23547 VDD.t720 VDD.t702 93.9934
R23548 VDD.n3740 VDD.t1115 93.81
R23549 VDD.n3768 VDD.t551 93.81
R23550 VDD.n2915 VDD.t2682 93.81
R23551 VDD.n2935 VDD.t2121 93.81
R23552 VDD.n3432 VDD.t1028 93.81
R23553 VDD.n3386 VDD.t1231 93.81
R23554 VDD.n2975 VDD.t788 93.81
R23555 VDD.n3322 VDD.t1899 93.81
R23556 VDD.n3536 VDD.t831 93.81
R23557 VDD.n2898 VDD.t1261 93.81
R23558 VDD.n3168 VDD.t1065 93.81
R23559 VDD.n3026 VDD.t1427 93.81
R23560 VDD.n2813 VDD.t741 93.81
R23561 VDD.n2764 VDD.t807 93.81
R23562 VDD.n2348 VDD.t120 93.81
R23563 VDD.n1846 VDD.t1468 93.81
R23564 VDD.n1363 VDD.t823 93.81
R23565 VDD.n1415 VDD.t1155 93.81
R23566 VDD.n1439 VDD.t859 93.81
R23567 VDD.n1463 VDD.t707 93.81
R23568 VDD.n1892 VDD.t2741 93.81
R23569 VDD.n1714 VDD.t1903 93.81
R23570 VDD.n1717 VDD.t725 93.81
R23571 VDD.n1542 VDD.t1419 93.81
R23572 VDD.n444 VDD.t1708 93.81
R23573 VDD.n607 VDD.t1668 93.81
R23574 VDD.n687 VDD.t2105 93.81
R23575 VDD.n711 VDD.t1590 93.81
R23576 VDD.n954 VDD.t1917 93.81
R23577 VDD.n354 VDD.n350 93.7417
R23578 VDD.n386 VDD.n385 93.7417
R23579 VDD.n350 VDD.n349 93.7417
R23580 VDD.n75 VDD.t517 93.3253
R23581 VDD.n38 VDD.t3002 93.3253
R23582 VDD.n386 VDD.n371 92.9887
R23583 VDD.n387 VDD.n341 92.5005
R23584 VDD.n341 VDD.t58 92.5005
R23585 VDD.n378 VDD.n372 92.5005
R23586 VDD.n378 VDD.t58 92.5005
R23587 VDD.n369 VDD.n338 92.5005
R23588 VDD.t464 VDD.n338 92.5005
R23589 VDD.n367 VDD.n366 92.5005
R23590 VDD.n366 VDD.t3035 92.5005
R23591 VDD.n356 VDD.n355 92.5005
R23592 VDD.n359 VDD.n358 92.5005
R23593 VDD.n358 VDD.t61 92.5005
R23594 VDD.n363 VDD.n362 92.5005
R23595 VDD.n365 VDD.n334 92.5005
R23596 VDD.t3035 VDD.n365 92.5005
R23597 VDD.n392 VDD.n391 92.5005
R23598 VDD.n391 VDD.t464 92.5005
R23599 VDD.n374 VDD.n373 92.5005
R23600 VDD.n374 VDD.t58 92.5005
R23601 VDD.n200 VDD.n199 92.5005
R23602 VDD.t2919 VDD.n200 92.5005
R23603 VDD.n203 VDD.n202 92.5005
R23604 VDD.n3983 VDD.n3982 92.4449
R23605 VDD.t729 VDD.t1299 92.315
R23606 VDD.t787 VDD.t1039 92.315
R23607 VDD.t1328 VDD.t3016 92.315
R23608 VDD.t1937 VDD.t1260 92.315
R23609 VDD.t1127 VDD.t1973 92.315
R23610 VDD.t779 VDD.t1843 92.315
R23611 VDD.t1738 VDD.t794 92.315
R23612 VDD.t1707 VDD.t877 92.315
R23613 VDD.t1804 VDD.t2087 92.315
R23614 VDD.n232 VDD.n231 91.4829
R23615 VDD.n321 VDD.t436 91.2567
R23616 VDD.t935 VDD.t1212 90.6365
R23617 VDD.t561 VDD.t1211 90.6365
R23618 VDD.t1352 VDD.t2238 90.6365
R23619 VDD.t2143 VDD.t2681 90.6365
R23620 VDD.t2737 VDD.n1483 90.6365
R23621 VDD.t2740 VDD.t2181 90.6365
R23622 VDD.t1091 VDD.t183 90.6365
R23623 VDD.t2897 VDD.t1154 90.6365
R23624 VDD.t1103 VDD.t2328 90.6365
R23625 VDD.t1109 VDD.t653 90.6365
R23626 VDD.t1940 VDD.t655 90.6365
R23627 VDD.n322 VDD.t450 90.3212
R23628 VDD.n317 VDD.n222 90.2911
R23629 VDD.t2253 VDD.t2248 89.8654
R23630 VDD.t2248 VDD.t2245 89.8654
R23631 VDD.t2245 VDD.t2242 89.8654
R23632 VDD.t3016 VDD.t177 88.9581
R23633 VDD.t1247 VDD.t2077 88.9581
R23634 VDD.t1469 VDD.t677 88.9581
R23635 VDD.t1197 VDD.t49 88.9581
R23636 VDD.t760 VDD.t1736 88.9581
R23637 VDD.t316 VDD.t1738 88.9581
R23638 VDD.t756 VDD.t885 88.9581
R23639 VDD.t822 VDD.t1593 88.9581
R23640 VDD.t1908 VDD.t473 88.9581
R23641 VDD.t2849 VDD.t1017 87.2797
R23642 VDD.t1156 VDD.n2866 87.2797
R23643 VDD.t1354 VDD.t2198 87.2797
R23644 VDD.n3703 VDD.t1684 86.7743
R23645 VDD.n4318 VDD.t1405 86.7743
R23646 VDD.n3987 VDD.t2880 86.7743
R23647 VDD.n2919 VDD.t1126 86.7743
R23648 VDD.n3458 VDD.t629 86.7743
R23649 VDD.n3361 VDD.t1100 86.7743
R23650 VDD.n3349 VDD.t3092 86.7743
R23651 VDD.n2990 VDD.t1588 86.7743
R23652 VDD.n3521 VDD.t713 86.7743
R23653 VDD.n2531 VDD.t504 86.7743
R23654 VDD.n2575 VDD.t2913 86.7743
R23655 VDD.n2171 VDD.t1123 86.7743
R23656 VDD.n2173 VDD.t639 86.7743
R23657 VDD.n2255 VDD.t1128 86.7743
R23658 VDD.n2739 VDD.t1506 86.7743
R23659 VDD.n2299 VDD.t1130 86.7743
R23660 VDD.n2324 VDD.t2915 86.7743
R23661 VDD.n2324 VDD.t102 86.7743
R23662 VDD.n1366 VDD.t833 86.7743
R23663 VDD.n1451 VDD.t2894 86.7743
R23664 VDD.n1451 VDD.t1448 86.7743
R23665 VDD.n1518 VDD.t5 86.7743
R23666 VDD.n1518 VDD.t2810 86.7743
R23667 VDD.n1803 VDD.t780 86.7743
R23668 VDD.n677 VDD.t987 86.7743
R23669 VDD.t1553 VDD.t2847 85.6012
R23670 VDD.t1404 VDD.t804 85.6012
R23671 VDD.t3100 VDD.t2311 85.6012
R23672 VDD.t647 VDD.t858 85.6012
R23673 VDD.t1177 VDD.t2354 85.6012
R23674 VDD.n326 VDD.n182 85.5545
R23675 VDD.n362 VDD.n361 84.2672
R23676 VDD.n361 VDD.n334 84.2672
R23677 VDD.n393 VDD.n334 84.2672
R23678 VDD.n393 VDD.n392 84.2672
R23679 VDD.n392 VDD.n335 84.2672
R23680 VDD.n373 VDD.n335 84.2672
R23681 VDD.t2106 VDD.t2046 83.9228
R23682 VDD.t615 VDD.t1990 83.9228
R23683 VDD.t2535 VDD.t480 83.9228
R23684 VDD.t483 VDD.t2104 83.9228
R23685 VDD.t1306 VDD.n989 82.5275
R23686 VDD.t802 VDD.t2031 82.2443
R23687 VDD.t207 VDD.t3091 82.2443
R23688 VDD.t2909 VDD.t1334 82.2443
R23689 VDD.t1640 VDD.t1667 82.2443
R23690 VDD.n3842 VDD.t68 80.5659
R23691 VDD.n3132 VDD.t3031 80.5659
R23692 VDD.t1214 VDD.t1431 80.5659
R23693 VDD.t1800 VDD.t1893 80.5659
R23694 VDD.t990 VDD.t555 80.5659
R23695 VDD.n2493 VDD.t1881 80.5659
R23696 VDD.t6 VDD.n2311 80.5659
R23697 VDD.t956 VDD.t1747 80.5659
R23698 VDD.n1675 VDD.t1326 80.5659
R23699 VDD.t724 VDD.t632 80.5659
R23700 VDD.t2264 VDD.t1501 80.5659
R23701 VDD.n1481 VDD.t1089 80.5659
R23702 VDD.t325 VDD.t1561 80.5659
R23703 VDD.t1297 VDD.t1697 80.5659
R23704 VDD.t1932 VDD.t2394 80.5659
R23705 VDD.t191 VDD.t1640 80.5659
R23706 VDD.t1764 VDD.t750 80.5659
R23707 VDD.t834 VDD.t1699 80.5659
R23708 VDD.n204 VDD.n195 80.5652
R23709 VDD.n231 VDD.n230 80.5652
R23710 VDD.n4312 VDD.t2042 79.0034
R23711 VDD.t2675 VDD.t207 78.8874
R23712 VDD.t415 VDD.t828 78.8874
R23713 VDD.t2210 VDD.t905 78.8874
R23714 VDD.t1693 VDD.t1336 78.8874
R23715 VDD.t2604 VDD.t42 78.8874
R23716 VDD.t300 VDD.t483 78.8874
R23717 VDD.n49 VDD.t2760 78.8874
R23718 VDD.n11 VDD.t2724 78.8874
R23719 VDD.t2616 VDD.t675 77.209
R23720 VDD.n3133 VDD.t2293 77.209
R23721 VDD.t3091 VDD.t1461 77.209
R23722 VDD.t2305 VDD.n2287 77.209
R23723 VDD.t2464 VDD.t2643 77.209
R23724 VDD.t2198 VDD.t647 77.209
R23725 VDD.t2637 VDD.t2634 77.209
R23726 VDD.t1906 VDD.t2449 77.209
R23727 VDD.t2339 VDD.t2169 77.209
R23728 VDD.t1276 VDD.t1171 75.5305
R23729 VDD.t804 VDD.t1400 75.5305
R23730 VDD.t1213 VDD.t561 75.5305
R23731 VDD.t2077 VDD.t1352 75.5305
R23732 VDD.t1270 VDD.t252 75.5305
R23733 VDD.t187 VDD.t244 75.5305
R23734 VDD.t2963 VDD.t1370 75.5305
R23735 VDD.n322 VDD.t2253 75.3458
R23736 VDD.t107 VDD.t2446 73.8521
R23737 VDD.t2446 VDD.t1019 73.8521
R23738 VDD.t1431 VDD.t1801 73.8521
R23739 VDD.t1430 VDD.t1800 73.8521
R23740 VDD.t1212 VDD.t327 73.8521
R23741 VDD.t2025 VDD.t992 73.8521
R23742 VDD.t1387 VDD.t2495 73.8521
R23743 VDD.n3574 VDD.t366 73.8521
R23744 VDD.n2345 VDD.t2877 73.8521
R23745 VDD.t17 VDD.t791 73.8521
R23746 VDD.t679 VDD.t2212 73.8521
R23747 VDD.t2075 VDD.t566 73.8521
R23748 VDD.t1236 VDD.t2809 73.8521
R23749 VDD.t1657 VDD.t1447 73.8521
R23750 VDD.t1559 VDD.t342 73.8521
R23751 VDD.t1593 VDD.t181 73.8521
R23752 VDD.t1841 VDD.t567 73.8521
R23753 VDD.t1444 VDD.t2569 73.8521
R23754 VDD.n1231 VDD.t352 73.8521
R23755 VDD.t2403 VDD.t1023 72.1736
R23756 VDD.t2584 VDD.t1076 72.1736
R23757 VDD.t1587 VDD.t1045 72.1736
R23758 VDD.t2923 VDD.t2143 72.1736
R23759 VDD.t2987 VDD.t2547 72.1736
R23760 VDD.t2547 VDD.t501 72.1736
R23761 VDD.t1653 VDD.t2196 72.1736
R23762 VDD.t2181 VDD.t2216 72.1736
R23763 VDD.t183 VDD.t2897 72.1736
R23764 VDD.n121 VDD.n117 71.9064
R23765 VDD.n125 VDD.n121 71.9064
R23766 VDD.n202 VDD.n201 70.7378
R23767 VDD.t1057 VDD.t122 70.4952
R23768 VDD.t1801 VDD.t1083 70.4952
R23769 VDD.t1799 VDD.t1424 70.4952
R23770 VDD.t626 VDD.t1080 70.4952
R23771 VDD.t1796 VDD.t1430 70.4952
R23772 VDD.t2238 VDD.t2025 70.4952
R23773 VDD.t1320 VDD.n1556 70.4952
R23774 VDD.t185 VDD.t875 70.4952
R23775 VDD.t877 VDD.t185 70.4952
R23776 VDD.n2949 VDD.t1531 69.9355
R23777 VDD.t1165 VDD.t1276 68.8168
R23778 VDD.t1400 VDD.t798 68.8168
R23779 VDD.t1021 VDD.t2403 68.8168
R23780 VDD.t1078 VDD.t2584 68.8168
R23781 VDD.t1436 VDD.t729 68.8168
R23782 VDD.t2905 VDD.t1509 68.8168
R23783 VDD.n1555 VDD.t669 68.8168
R23784 VDD.t1843 VDD.t777 68.8168
R23785 VDD.t2216 VDD.t2179 68.8168
R23786 VDD.t2541 VDD.t1655 68.8168
R23787 VDD.t1644 VDD.t2963 68.8168
R23788 VDD.t2794 VDD.t1804 68.8168
R23789 VDD.n357 VDD.n356 68.2232
R23790 VDD.n3703 VDD.t2848 68.0124
R23791 VDD.n4318 VDD.t1401 68.0124
R23792 VDD.n2919 VDD.t2854 68.0124
R23793 VDD.n3458 VDD.t2840 68.0124
R23794 VDD.n3361 VDD.t1492 68.0124
R23795 VDD.n3349 VDD.t2676 68.0124
R23796 VDD.n2990 VDD.t1586 68.0124
R23797 VDD.n3521 VDD.t2842 68.0124
R23798 VDD.n2171 VDD.t965 68.0124
R23799 VDD.n2173 VDD.t2846 68.0124
R23800 VDD.n2255 VDD.t2836 68.0124
R23801 VDD.n2739 VDD.t678 68.0124
R23802 VDD.n2299 VDD.t693 68.0124
R23803 VDD.n1366 VDD.t1009 68.0124
R23804 VDD.n1803 VDD.t778 68.0124
R23805 VDD.n677 VDD.t652 68.0124
R23806 VDD.t685 VDD.t996 67.1383
R23807 VDD.t327 VDD.t1328 67.1383
R23808 VDD.t1757 VDD.t1389 67.1383
R23809 VDD.n3574 VDD.t1579 67.1383
R23810 VDD.t1129 VDD.t2458 67.1383
R23811 VDD.t714 VDD.t679 67.1383
R23812 VDD.t1546 VDD.t2835 67.1383
R23813 VDD.t2776 VDD.t105 67.1383
R23814 VDD.t2809 VDD.t1244 67.1383
R23815 VDD.t1447 VDD.t1661 67.1383
R23816 VDD.t567 VDD.t1839 67.1383
R23817 VDD.t2569 VDD.t425 67.1383
R23818 VDD.n1231 VDD.t2227 67.1383
R23819 VDD.n3986 VDD.t1265 66.8398
R23820 VDD.n2532 VDD.t2094 66.8398
R23821 VDD.n2576 VDD.t1205 66.8398
R23822 VDD.n4312 VDD.t2192 66.1981
R23823 VDD.n363 VDD.n348 65.5397
R23824 VDD.t1797 VDD.t742 65.4599
R23825 VDD.t1513 VDD.t1081 65.4599
R23826 VDD.t2218 VDD.t133 65.4599
R23827 VDD.t2907 VDD.t979 65.4599
R23828 VDD.t248 VDD.t1270 65.4599
R23829 VDD.t252 VDD.t187 65.4599
R23830 VDD.t1394 VDD.t1152 65.4599
R23831 VDD.t1563 VDD.t1762 65.4599
R23832 VDD.n402 VDD.t465 63.8266
R23833 VDD.n3573 VDD.t690 63.7814
R23834 VDD.t2062 VDD.t2575 63.7814
R23835 VDD.t796 VDD.t1979 63.7814
R23836 VDD.t2449 VDD.t1910 63.7814
R23837 VDD.t845 VDD.t1324 63.7814
R23838 VDD.t1589 VDD.t1051 63.7814
R23839 VDD.t2226 VDD.t834 63.7814
R23840 VDD.t2308 VDD.t2229 63.7814
R23841 VDD.n396 VDD.t3036 63.7312
R23842 VDD.n3734 VDD.t295 63.3219
R23843 VDD.n3740 VDD.t299 63.3219
R23844 VDD.n4018 VDD.t399 63.3219
R23845 VDD.n4018 VDD.t588 63.3219
R23846 VDD.n3779 VDD.t118 63.3219
R23847 VDD.n2915 VDD.t2924 63.3219
R23848 VDD.n3502 VDD.t2926 63.3219
R23849 VDD.n2932 VDD.t319 63.3219
R23850 VDD.n2932 VDD.t1397 63.3219
R23851 VDD.n2935 VDD.t2906 63.3219
R23852 VDD.n2942 VDD.t180 63.3219
R23853 VDD.n2956 VDD.t2201 63.3219
R23854 VDD.n3432 VDD.t2215 63.3219
R23855 VDD.n3386 VDD.t2860 63.3219
R23856 VDD.n3357 VDD.t178 63.3219
R23857 VDD.n2975 VDD.t134 63.3219
R23858 VDD.n3322 VDD.t572 63.3219
R23859 VDD.n2980 VDD.t132 63.3219
R23860 VDD.n2983 VDD.t287 63.3219
R23861 VDD.n3261 VDD.t3026 63.3219
R23862 VDD.n3261 VDD.t334 63.3219
R23863 VDD.n3240 VDD.t2982 63.3219
R23864 VDD.n3240 VDD.t2822 63.3219
R23865 VDD.n3276 VDD.t1789 63.3219
R23866 VDD.n3276 VDD.t3007 63.3219
R23867 VDD.n3282 VDD.t14 63.3219
R23868 VDD.n3282 VDD.t226 63.3219
R23869 VDD.n3529 VDD.t2858 63.3219
R23870 VDD.n3532 VDD.t190 63.3219
R23871 VDD.n3536 VDD.t2902 63.3219
R23872 VDD.n2898 VDD.t2908 63.3219
R23873 VDD.n3015 VDD.t401 63.3219
R23874 VDD.n3159 VDD.t283 63.3219
R23875 VDD.n3168 VDD.t289 63.3219
R23876 VDD.n3026 VDD.t576 63.3219
R23877 VDD.n3180 VDD.t574 63.3219
R23878 VDD.n2813 VDD.t2864 63.3219
R23879 VDD.n2244 VDD.t188 63.3219
R23880 VDD.n2764 VDD.t2203 63.3219
R23881 VDD.n2264 VDD.t2213 63.3219
R23882 VDD.n2346 VDD.t1854 63.3219
R23883 VDD.n2346 VDD.t745 63.3219
R23884 VDD.n2362 VDD.t1692 63.3219
R23885 VDD.n2386 VDD.t1670 63.3219
R23886 VDD.n1846 VDD.t291 63.3219
R23887 VDD.n1363 VDD.t182 63.3219
R23888 VDD.n1389 VDD.t2862 63.3219
R23889 VDD.n1415 VDD.t184 63.3219
R23890 VDD.n1422 VDD.t2904 63.3219
R23891 VDD.n1439 VDD.t2199 63.3219
R23892 VDD.n1445 VDD.t2207 63.3219
R23893 VDD.n1463 VDD.t2205 63.3219
R23894 VDD.n1468 VDD.t2209 63.3219
R23895 VDD.n1471 VDD.t2211 63.3219
R23896 VDD.n1892 VDD.t2217 63.3219
R23897 VDD.n1513 VDD.t293 63.3219
R23898 VDD.n1702 VDD.t570 63.3219
R23899 VDD.n1565 VDD.t79 63.3219
R23900 VDD.n1714 VDD.t303 63.3219
R23901 VDD.n1717 VDD.t75 63.3219
R23902 VDD.n1759 VDD.t83 63.3219
R23903 VDD.n1542 VDD.t50 63.3219
R23904 VDD.n1016 VDD.t297 63.3219
R23905 VDD.n444 VDD.t186 63.3219
R23906 VDD.n547 VDD.t194 63.3219
R23907 VDD.n607 VDD.t192 63.3219
R23908 VDD.n614 VDD.t176 63.3219
R23909 VDD.n687 VDD.t301 63.3219
R23910 VDD.n693 VDD.t285 63.3219
R23911 VDD.n711 VDD.t568 63.3219
R23912 VDD.n954 VDD.t43 63.3219
R23913 VDD.n737 VDD.t81 63.3219
R23914 VDD.n2646 VDD.n2645 63.0618
R23915 VDD.t2031 VDD.t800 62.103
R23916 VDD.t1934 VDD.t787 62.103
R23917 VDD.t1260 VDD.t2193 62.103
R23918 VDD.t1548 VDD.t1127 62.103
R23919 VDD.t2961 VDD.t1242 62.103
R23920 VDD.t907 VDD.t2210 62.103
R23921 VDD.t905 VDD.t2738 62.103
R23922 VDD.t832 VDD.t1449 62.103
R23923 VDD.t1336 VDD.t2909 62.103
R23924 VDD.n49 VDD.t2762 62.103
R23925 VDD.n11 VDD.t2720 62.103
R23926 VDD.t517 VDD.t525 61.7891
R23927 VDD.t525 VDD.t519 61.7891
R23928 VDD.t519 VDD.t523 61.7891
R23929 VDD.t523 VDD.t527 61.7891
R23930 VDD.t527 VDD.t531 61.7891
R23931 VDD.t531 VDD.t526 61.7891
R23932 VDD.t526 VDD.t530 61.7891
R23933 VDD.t530 VDD.t524 61.7891
R23934 VDD.t524 VDD.t516 61.7891
R23935 VDD.t516 VDD.t520 61.7891
R23936 VDD.t520 VDD.t518 61.7891
R23937 VDD.t518 VDD.t528 61.7891
R23938 VDD.t528 VDD.t522 61.7891
R23939 VDD.t522 VDD.t529 61.7891
R23940 VDD.t529 VDD.t521 61.7891
R23941 VDD.t521 VDD.t2052 61.7891
R23942 VDD.t2052 VDD.t2054 61.7891
R23943 VDD.t2054 VDD.t2058 61.7891
R23944 VDD.t2058 VDD.t2051 61.7891
R23945 VDD.t2051 VDD.t2056 61.7891
R23946 VDD.t2055 VDD.t2057 61.7891
R23947 VDD.t2057 VDD.t2053 61.7891
R23948 VDD.t2053 VDD.t2931 61.7891
R23949 VDD.t2931 VDD.t2930 61.7891
R23950 VDD.t2930 VDD.t2932 61.7891
R23951 VDD.t2932 VDD.t2933 61.7891
R23952 VDD.t2933 VDD.t255 61.7891
R23953 VDD.t255 VDD.t254 61.7891
R23954 VDD.t254 VDD.t602 61.7891
R23955 VDD.t2039 VDD.t3039 61.7891
R23956 VDD.t2038 VDD.t2039 61.7891
R23957 VDD.t88 VDD.t2038 61.7891
R23958 VDD.t86 VDD.t88 61.7891
R23959 VDD.t89 VDD.t86 61.7891
R23960 VDD.t87 VDD.t89 61.7891
R23961 VDD.t579 VDD.t87 61.7891
R23962 VDD.t578 VDD.t579 61.7891
R23963 VDD.t583 VDD.t578 61.7891
R23964 VDD.t581 VDD.t584 61.7891
R23965 VDD.t582 VDD.t581 61.7891
R23966 VDD.t577 VDD.t582 61.7891
R23967 VDD.t580 VDD.t577 61.7891
R23968 VDD.t3003 VDD.t580 61.7891
R23969 VDD.t3005 VDD.t3003 61.7891
R23970 VDD.t2991 VDD.t3005 61.7891
R23971 VDD.t2998 VDD.t2991 61.7891
R23972 VDD.t3000 VDD.t2998 61.7891
R23973 VDD.t3004 VDD.t3000 61.7891
R23974 VDD.t2992 VDD.t3004 61.7891
R23975 VDD.t2997 VDD.t2992 61.7891
R23976 VDD.t2990 VDD.t2997 61.7891
R23977 VDD.t2993 VDD.t2990 61.7891
R23978 VDD.t2999 VDD.t2993 61.7891
R23979 VDD.t3001 VDD.t2999 61.7891
R23980 VDD.t2995 VDD.t3001 61.7891
R23981 VDD.t2996 VDD.t2995 61.7891
R23982 VDD.t2994 VDD.t2996 61.7891
R23983 VDD.t3002 VDD.t2994 61.7891
R23984 VDD.t634 VDD.t1214 60.4245
R23985 VDD.t1893 VDD.t818 60.4245
R23986 VDD.t1291 VDD.t956 60.4245
R23987 VDD.t2024 VDD.t1544 60.4245
R23988 VDD.t1418 VDD.t598 60.4245
R23989 VDD.t2823 VDD.t722 60.4245
R23990 VDD.t1555 VDD.t325 60.4245
R23991 VDD.t1507 VDD.t2112 60.4245
R23992 VDD.t750 VDD.t754 60.4245
R23993 VDD.t1699 VDD.t1764 60.4245
R23994 VDD.n355 VDD.n342 59.4829
R23995 VDD.n367 VDD.n342 59.4829
R23996 VDD.n368 VDD.n367 59.4829
R23997 VDD.n369 VDD.n368 59.4829
R23998 VDD.n370 VDD.n369 59.4829
R23999 VDD.n372 VDD.n370 59.4829
R24000 VDD.t421 VDD.t2134 58.7461
R24001 VDD.t800 VDD.t1404 58.7461
R24002 VDD.t1777 VDD.t2106 58.7461
R24003 VDD.t1983 VDD.t2183 58.7461
R24004 VDD.t1667 VDD.t1642 58.7461
R24005 VDD.t1282 VDD.t1493 57.0676
R24006 VDD.t1992 VDD.t615 57.0676
R24007 VDD.t1990 VDD.t2903 57.0676
R24008 VDD.n3831 VDD.t2935 55.4067
R24009 VDD.n3832 VDD.t277 55.4067
R24010 VDD.n3835 VDD.t69 55.4067
R24011 VDD.n3845 VDD.t2872 55.4067
R24012 VDD.n3846 VDD.t315 55.4067
R24013 VDD.n4418 VDD.t271 55.4067
R24014 VDD.n4379 VDD.t3075 55.4067
R24015 VDD.n4380 VDD.t380 55.4067
R24016 VDD.n4383 VDD.t470 55.4067
R24017 VDD.n4388 VDD.t3062 55.4067
R24018 VDD.n3058 VDD.t126 55.4067
R24019 VDD.n3059 VDD.t3105 55.4067
R24020 VDD.n3043 VDD.t3032 55.4067
R24021 VDD.n3065 VDD.t265 55.4067
R24022 VDD.n3591 VDD.t114 55.4067
R24023 VDD.n3593 VDD.t2953 55.4067
R24024 VDD.n3596 VDD.t2647 55.4067
R24025 VDD.n3597 VDD.t369 55.4067
R24026 VDD.n2351 VDD.t2162 55.4067
R24027 VDD.n2401 VDD.t1252 55.4067
R24028 VDD.n2467 VDD.t1882 55.4067
R24029 VDD.n2470 VDD.t609 55.4067
R24030 VDD.n2472 VDD.t539 55.4067
R24031 VDD.n2120 VDD.t2867 55.4067
R24032 VDD.n2121 VDD.t1423 55.4067
R24033 VDD.n2124 VDD.t307 55.4067
R24034 VDD.n2125 VDD.t849 55.4067
R24035 VDD.n1580 VDD.t1710 55.4067
R24036 VDD.n1523 VDD.t1199 55.4067
R24037 VDD.n1649 VDD.t1327 55.4067
R24038 VDD.n1652 VDD.t874 55.4067
R24039 VDD.n1654 VDD.t2130 55.4067
R24040 VDD.n1286 VDD.t2095 55.4067
R24041 VDD.n1287 VDD.t1141 55.4067
R24042 VDD.n1290 VDD.t2137 55.4067
R24043 VDD.n1291 VDD.t2123 55.4067
R24044 VDD.n550 VDD.t967 55.4067
R24045 VDD.n588 VDD.t1253 55.4067
R24046 VDD.n606 VDD.t1995 55.4067
R24047 VDD.n625 VDD.t1542 55.4067
R24048 VDD.n654 VDD.t1399 55.4067
R24049 VDD.n672 VDD.t2097 55.4067
R24050 VDD.n690 VDD.t1508 55.4067
R24051 VDD.n710 VDD.t1052 55.4067
R24052 VDD.n727 VDD.t1191 55.4067
R24053 VDD.n739 VDD.t844 55.4067
R24054 VDD.n761 VDD.t2653 55.4067
R24055 VDD.n778 VDD.t682 55.4067
R24056 VDD.n779 VDD.t959 55.4067
R24057 VDD.n782 VDD.t1279 55.4067
R24058 VDD.n783 VDD.t1476 55.4067
R24059 VDD.n785 VDD.t973 55.4067
R24060 VDD.n789 VDD.t2696 55.4067
R24061 VDD.n800 VDD.t1227 55.4067
R24062 VDD.n850 VDD.t934 55.4067
R24063 VDD.n467 VDD.t898 55.4067
R24064 VDD.n469 VDD.t2733 55.4067
R24065 VDD.n472 VDD.t766 55.4067
R24066 VDD.n473 VDD.t3084 55.4067
R24067 VDD.n476 VDD.t1637 55.4067
R24068 VDD.n481 VDD.t620 55.4067
R24069 VDD.t937 VDD.t419 55.3892
R24070 VDD.t2883 VDD.t1618 55.3892
R24071 VDD.t2841 VDD.t2778 55.3892
R24072 VDD.t858 VDD.t645 55.3892
R24073 VDD.t1008 VDD.t883 55.3892
R24074 VDD.t2354 VDD.t813 55.3892
R24075 VDD.t8 VDD.t1485 55.3892
R24076 VDD.n260 VDD.t2490 54.4158
R24077 VDD.n260 VDD.t2452 54.4158
R24078 VDD.n266 VDD.t2372 54.4158
R24079 VDD.n266 VDD.t2267 54.4158
R24080 VDD.t1210 VDD.t935 53.7107
R24081 VDD.t2458 VDD.t793 53.7107
R24082 VDD.t2102 VDD.t269 53.7107
R24083 VDD.t655 VDD.t2147 53.7107
R24084 VDD.t3079 VDD.t720 53.7107
R24085 VDD.n2949 VDD.t1602 53.1905
R24086 VDD.t1348 VDD.t1603 52.0323
R24087 VDD.t677 VDD.t1471 52.0323
R24088 VDD.t1483 VDD.t1616 52.0323
R24089 VDD.t2712 VDD.t1050 52.0323
R24090 VDD.t1736 VDD.t316 52.0323
R24091 VDD.t885 VDD.t758 52.0323
R24092 VDD.t1591 VDD.t822 52.0323
R24093 VDD.t473 VDD.t1644 52.0323
R24094 VDD.t377 VDD.t1849 52.0323
R24095 VDD.n217 VDD.t2247 50.3754
R24096 VDD.t2244 VDD.n217 50.3754
R24097 VDD.t553 VDD.t1057 50.3539
R24098 VDD.t1877 VDD.t2882 50.3539
R24099 VDD.t2328 VDD.t1105 50.3539
R24100 VDD.t653 VDD.t1940 50.3539
R24101 VDD.n233 VDD.n224 48.9417
R24102 VDD.t1045 VDD.t2711 48.6754
R24103 VDD.t1532 VDD.t1511 48.6754
R24104 VDD.n326 VDD.n325 48.6258
R24105 VDD.n131 VDD.t1474 48.6146
R24106 VDD.t2685 VDD.n131 48.6146
R24107 VDD.n990 VDD.t1306 47.7312
R24108 VDD.t294 VDD.t3093 46.997
R24109 VDD.t992 VDD.t919 46.997
R24110 VDD.t3089 VDD.t1628 46.997
R24111 VDD.t348 VDD.t556 46.997
R24112 VDD.t563 VDD.t2096 46.997
R24113 VDD.n198 VDD.n196 46.2505
R24114 VDD.n197 VDD.n195 46.2505
R24115 VDD.n197 VDD.n193 46.2505
R24116 VDD.n230 VDD.n229 46.2505
R24117 VDD.n227 VDD.n224 46.2505
R24118 VDD.n117 VDD.n113 46.2505
R24119 VDD.n123 VDD.n113 46.2505
R24120 VDD.n125 VDD.n124 46.2505
R24121 VDD.n124 VDD.n123 46.2505
R24122 VDD.n993 VDD.n992 46.0805
R24123 VDD.t2253 VDD.t2248 45.6825
R24124 VDD.t2248 VDD.t2245 45.6825
R24125 VDD.t2245 VDD.t2242 45.6825
R24126 VDD.t2843 VDD.n4250 45.3185
R24127 VDD.t393 VDD.t1673 45.3185
R24128 VDD.t2200 VDD.t2026 45.3185
R24129 VDD.t1749 VDD.t179 45.3185
R24130 VDD.t1222 VDD.t2208 45.3185
R24131 VDD.t2885 VDD.t1410 45.3185
R24132 VDD.t173 VDD.t1412 45.3185
R24133 VDD.t1390 VDD.t1406 45.3185
R24134 VDD.t1392 VDD.t1408 45.3185
R24135 VDD.t843 VDD.t80 45.3185
R24136 VDD.t2167 VDD.t284 45.3185
R24137 VDD.t2242 VDD.n187 44.9329
R24138 VDD.t2251 VDD.n187 44.9329
R24139 VDD.t2249 VDD.n190 44.9329
R24140 VDD.t2255 VDD.n190 44.9329
R24141 VDD.n218 VDD.n188 43.9332
R24142 VDD.n216 VDD.n192 43.9332
R24143 VDD.t1461 VDD.t1925 43.6401
R24144 VDD.t2081 VDD.t1055 43.6401
R24145 VDD.t193 VDD.t1053 43.6401
R24146 VDD.n138 VDD.n134 43.1501
R24147 VDD.n2326 VDD.t2729 42.3555
R24148 VDD.n1479 VDD.t1502 42.3555
R24149 VDD.n1522 VDD.t1026 42.3555
R24150 VDD.t2030 VDD.t1604 41.9616
R24151 VDD.n3747 VDD.t27 41.5552
R24152 VDD.n3747 VDD.t2136 41.5552
R24153 VDD.n2927 VDD.t1619 41.5552
R24154 VDD.n2927 VDD.t365 41.5552
R24155 VDD.n3370 VDD.t1209 41.5552
R24156 VDD.n3370 VDD.t361 41.5552
R24157 VDD.n3368 VDD.t198 41.5552
R24158 VDD.n3368 VDD.t2237 41.5552
R24159 VDD.n2970 VDD.t2671 41.5552
R24160 VDD.n2970 VDD.t31 41.5552
R24161 VDD.n3337 VDD.t2221 41.5552
R24162 VDD.n3337 VDD.t23 41.5552
R24163 VDD.n3522 VDD.t689 41.5552
R24164 VDD.n3522 VDD.t355 41.5552
R24165 VDD.n2910 VDD.t978 41.5552
R24166 VDD.n2910 VDD.t357 41.5552
R24167 VDD.n2911 VDD.t1580 41.5552
R24168 VDD.n2911 VDD.t367 41.5552
R24169 VDD.n3033 VDD.t1363 41.5552
R24170 VDD.n3033 VDD.t1798 41.5552
R24171 VDD.n3021 VDD.t1082 41.5552
R24172 VDD.n3021 VDD.t39 41.5552
R24173 VDD.n2830 VDD.t2115 41.5552
R24174 VDD.n2830 VDD.t351 41.5552
R24175 VDD.n2251 VDD.t1545 41.5552
R24176 VDD.n2251 VDD.t200 41.5552
R24177 VDD.n2079 VDD.t853 41.5552
R24178 VDD.n2079 VDD.t349 41.5552
R24179 VDD.n1409 VDD.t2060 41.5552
R24180 VDD.n1409 VDD.t363 41.5552
R24181 VDD.n1431 VDD.t947 41.5552
R24182 VDD.n1431 VDD.t202 41.5552
R24183 VDD.n1457 VDD.t952 41.5552
R24184 VDD.n1457 VDD.t204 41.5552
R24185 VDD.n1488 VDD.t41 41.5552
R24186 VDD.n1488 VDD.t2735 41.5552
R24187 VDD.n1502 VDD.t1615 41.5552
R24188 VDD.n1502 VDD.t25 41.5552
R24189 VDD.n1559 VDD.t631 41.5552
R24190 VDD.n1559 VDD.t1359 41.5552
R24191 VDD.n1730 VDD.t1884 41.5552
R24192 VDD.n1730 VDD.t1365 41.5552
R24193 VDD.n1786 VDD.t1879 41.5552
R24194 VDD.n1786 VDD.t1361 41.5552
R24195 VDD.n529 VDD.t2228 41.5552
R24196 VDD.n529 VDD.t353 41.5552
R24197 VDD.n600 VDD.t2071 41.5552
R24198 VDD.n600 VDD.t359 41.5552
R24199 VDD.n680 VDD.t2146 41.5552
R24200 VDD.n680 VDD.t33 41.5552
R24201 VDD.n702 VDD.t1097 41.5552
R24202 VDD.n702 VDD.t35 41.5552
R24203 VDD.n971 VDD.t1369 41.5552
R24204 VDD.n971 VDD.t1367 41.5552
R24205 VDD.t1124 VDD.t990 40.2832
R24206 VDD.t1747 VDD.t169 40.2832
R24207 VDD.t2833 VDD.t1835 40.2832
R24208 VDD.t1238 VDD.t4 40.2832
R24209 VDD.t2956 VDD.t1240 40.2832
R24210 VDD.t1663 VDD.t2893 40.2832
R24211 VDD.t3014 VDD.t1659 40.2832
R24212 VDD.t1088 VDD.t2061 40.2832
R24213 VDD.t1561 VDD.t1116 40.2832
R24214 VDD.t2756 VDD.t3050 40.2832
R24215 VDD.t2722 VDD.t3046 40.2832
R24216 VDD.n2284 VDD.t3018 39.7937
R24217 VDD.n2321 VDD.t3 39.7937
R24218 VDD.n2331 VDD.t2827 39.7937
R24219 VDD.n2502 VDD.t591 39.7937
R24220 VDD.n1356 VDD.t93 39.7937
R24221 VDD.n1410 VDD.t339 39.7937
R24222 VDD.n1428 VDD.t2886 39.7937
R24223 VDD.n1499 VDD.t218 39.7937
R24224 VDD.n1738 VDD.t2970 39.7937
R24225 VDD.t1013 VDD.t286 38.6047
R24226 VDD.t2925 VDD.t2853 38.6047
R24227 VDD.t2857 VDD.t1068 38.6047
R24228 VDD.t51 VDD.t292 38.6047
R24229 VDD.t860 VDD.t856 38.6047
R24230 VDD.t611 VDD.t2985 38.6047
R24231 VDD.t2819 VDD.t2799 38.6047
R24232 VDD.t1256 VDD.t346 38.6047
R24233 VDD.n3011 VDD.t991 38.4155
R24234 VDD.n3011 VDD.t394 38.4155
R24235 VDD.n2857 VDD.t2896 38.4155
R24236 VDD.n2857 VDD.t2777 38.4155
R24237 VDD.n92 VDD.t2795 38.4155
R24238 VDD.n4201 VDD.t1351 37.4305
R24239 VDD.n4189 VDD.t1866 37.4305
R24240 VDD.n3706 VDD.t1170 37.4305
R24241 VDD.n3716 VDD.t1145 37.4305
R24242 VDD.n3732 VDD.t997 37.4305
R24243 VDD.n3752 VDD.t2751 37.4305
R24244 VDD.n4367 VDD.t1952 37.4305
R24245 VDD.n4341 VDD.t799 37.4305
R24246 VDD.n4303 VDD.t2000 37.4305
R24247 VDD.n4384 VDD.t1315 37.4305
R24248 VDD.n1597 VDD.t140 37.4305
R24249 VDD.n846 VDD.t2787 37.4305
R24250 VDD.n477 VDD.t930 37.4305
R24251 VDD.n207 VDD.n183 37.2235
R24252 VDD.n207 VDD.n206 37.2235
R24253 VDD.n206 VDD.n205 37.2235
R24254 VDD.n325 VDD.n183 37.1499
R24255 VDD.n4363 VDD.t2187 36.9263
R24256 VDD.t115 VDD.t375 36.9263
R24257 VDD.t2875 VDD.t1434 36.9263
R24258 VDD.t427 VDD.t1620 36.9263
R24259 VDD.t621 VDD.t1159 36.9263
R24260 VDD.t2104 VDD.t215 36.9263
R24261 VDD.n394 VDD.n393 36.4805
R24262 VDD.n3697 VDD.t2109 36.4455
R24263 VDD.n3726 VDD.t1190 36.4455
R24264 VDD.n3743 VDD.t1375 36.4455
R24265 VDD.n3816 VDD.t1037 36.4455
R24266 VDD.n4347 VDD.t1085 36.4455
R24267 VDD.n3804 VDD.t1112 36.4455
R24268 VDD.n3348 VDD.t1462 36.4455
R24269 VDD.n2989 VDD.t2158 36.4455
R24270 VDD.n2382 VDD.t1289 36.4455
R24271 VDD.n1476 VDD.t2180 36.4455
R24272 VDD.t2056 VDD.n74 36.2048
R24273 VDD.t584 VDD.n37 36.2048
R24274 VDD.n4375 VDD.t618 36.1587
R24275 VDD.n4375 VDD.t21 36.1587
R24276 VDD.n3746 VDD.t2916 36.1587
R24277 VDD.n3746 VDD.t1540 36.1587
R24278 VDD.n3825 VDD.t2829 36.1587
R24279 VDD.n3825 VDD.t1686 36.1587
R24280 VDD.n3826 VDD.t108 36.1587
R24281 VDD.n3826 VDD.t1020 36.1587
R24282 VDD.n3844 VDD.t3082 36.1587
R24283 VDD.n3844 VDD.t1816 36.1587
R24284 VDD.n4009 VDD.t1333 36.1587
R24285 VDD.n4009 VDD.t2035 36.1587
R24286 VDD.n3757 VDD.t3060 36.1587
R24287 VDD.n3757 VDD.t2015 36.1587
R24288 VDD.n3786 VDD.t1421 36.1587
R24289 VDD.n3786 VDD.t2037 36.1587
R24290 VDD.n3951 VDD.t206 36.1587
R24291 VDD.n3951 VDD.t684 36.1587
R24292 VDD.n1533 VDD.t2160 36.1587
R24293 VDD.n1533 VDD.t2103 36.1587
R24294 VDD.n464 VDD.t2743 36.1587
R24295 VDD.n464 VDD.t67 36.1587
R24296 VDD.n538 VDD.t2808 36.1587
R24297 VDD.n538 VDD.t1761 36.1587
R24298 VDD.n610 VDD.t3080 36.1587
R24299 VDD.n610 VDD.t703 36.1587
R24300 VDD.n618 VDD.t259 36.1587
R24301 VDD.n618 VDD.t1984 36.1587
R24302 VDD.n664 VDD.t1151 36.1587
R24303 VDD.n664 VDD.t2033 36.1587
R24304 VDD.n694 VDD.t378 36.1587
R24305 VDD.n694 VDD.t2168 36.1587
R24306 VDD.n705 VDD.t3068 36.1587
R24307 VDD.n705 VDD.t644 36.1587
R24308 VDD.n718 VDD.t3038 36.1587
R24309 VDD.n718 VDD.t1831 36.1587
R24310 VDD.n746 VDD.t3086 36.1587
R24311 VDD.n746 VDD.t1986 36.1587
R24312 VDD.n450 VDD.t1962 36.1587
R24313 VDD.n450 VDD.t3041 36.1587
R24314 VDD.n640 VDD.t2980 36.1587
R24315 VDD.n640 VDD.t917 36.1587
R24316 VDD.n732 VDD.t124 36.1587
R24317 VDD.n732 VDD.t2804 36.1587
R24318 VDD.n767 VDD.t1005 36.1587
R24319 VDD.n767 VDD.t257 36.1587
R24320 VDD.n793 VDD.t625 36.1587
R24321 VDD.n793 VDD.t604 36.1587
R24322 VDD.t456 VDD.n321 36.035
R24323 VDD.n3003 VDD.t376 35.4605
R24324 VDD.t1928 VDD.t1374 35.2479
R24325 VDD.t1346 VDD.t1356 35.2479
R24326 VDD.t1583 VDD.t865 35.2479
R24327 VDD.t30 VDD.t2677 35.2479
R24328 VDD.t1396 VDD.t1829 35.2479
R24329 VDD.t1624 VDD.t2851 35.2479
R24330 VDD.t1781 VDD.t2 35.2479
R24331 VDD.t1272 VDD.t1769 35.2479
R24332 VDD.t2125 VDD.t1779 35.2479
R24333 VDD.t228 VDD.t1871 35.2479
R24334 VDD.t431 VDD.t1613 35.2479
R24335 VDD.n235 VDD.n233 34.7055
R24336 VDD.n4093 VDD.n4092 34.6358
R24337 VDD.n4088 VDD.n4087 34.6358
R24338 VDD.n3416 VDD.n3415 34.6358
R24339 VDD.n2539 VDD.n2538 34.6358
R24340 VDD.n1899 VDD.n1477 34.6358
R24341 VDD.n1773 VDD.n1539 34.6358
R24342 VDD.n576 VDD.n575 34.6358
R24343 VDD.n1216 VDD.n1215 34.6358
R24344 VDD.n1193 VDD.n611 34.6358
R24345 VDD.n1045 VDD.n1044 34.6358
R24346 VDD.n1009 VDD.n1008 34.6358
R24347 VDD.n4108 VDD.n3735 34.6358
R24348 VDD.n4104 VDD.n4101 34.6358
R24349 VDD.n4089 VDD.n4088 34.6358
R24350 VDD.n3998 VDD.n3997 34.6358
R24351 VDD.n3998 VDD.n3774 34.6358
R24352 VDD.n4002 VDD.n3774 34.6358
R24353 VDD.n3517 VDD.n2912 34.6358
R24354 VDD.n3514 VDD.n3513 34.6358
R24355 VDD.n3504 VDD.n3501 34.6358
R24356 VDD.n3508 VDD.n3507 34.6358
R24357 VDD.n3509 VDD.n3508 34.6358
R24358 VDD.n3495 VDD.n3494 34.6358
R24359 VDD.n3488 VDD.n3487 34.6358
R24360 VDD.n3461 VDD.n3457 34.6358
R24361 VDD.n3465 VDD.n2947 34.6358
R24362 VDD.n3468 VDD.n3467 34.6358
R24363 VDD.n3455 VDD.n2951 34.6358
R24364 VDD.n3442 VDD.n2957 34.6358
R24365 VDD.n3446 VDD.n2957 34.6358
R24366 VDD.n3438 VDD.n2960 34.6358
R24367 VDD.n3434 VDD.n3431 34.6358
R24368 VDD.n3376 VDD.n3366 34.6358
R24369 VDD.n3385 VDD.n3384 34.6358
R24370 VDD.n3384 VDD.n3363 34.6358
R24371 VDD.n3380 VDD.n3363 34.6358
R24372 VDD.n3380 VDD.n3379 34.6358
R24373 VDD.n3343 VDD.n3342 34.6358
R24374 VDD.n3339 VDD.n3336 34.6358
R24375 VDD.n3336 VDD.n3335 34.6358
R24376 VDD.n3329 VDD.n3328 34.6358
R24377 VDD.n3324 VDD.n3321 34.6358
R24378 VDD.n3264 VDD.n3263 34.6358
R24379 VDD.n3269 VDD.n3268 34.6358
R24380 VDD.n3274 VDD.n3238 34.6358
R24381 VDD.n3289 VDD.n3288 34.6358
R24382 VDD.n3568 VDD.n2913 34.6358
R24383 VDD.n3565 VDD.n3564 34.6358
R24384 VDD.n3560 VDD.n3559 34.6358
R24385 VDD.n3544 VDD.n3534 34.6358
R24386 VDD.n3539 VDD.n3538 34.6358
R24387 VDD.n3650 VDD.n2901 34.6358
R24388 VDD.n3646 VDD.n2901 34.6358
R24389 VDD.n3643 VDD.n3642 34.6358
R24390 VDD.n3230 VDD.n3229 34.6358
R24391 VDD.n3224 VDD.n3004 34.6358
R24392 VDD.n3216 VDD.n3008 34.6358
R24393 VDD.n3205 VDD.n3012 34.6358
R24394 VDD.n3209 VDD.n3012 34.6358
R24395 VDD.n3162 VDD.n3029 34.6358
R24396 VDD.n3175 VDD.n3024 34.6358
R24397 VDD.n2204 VDD.n2203 34.6358
R24398 VDD.n2203 VDD.n2169 34.6358
R24399 VDD.n2199 VDD.n2198 34.6358
R24400 VDD.n2196 VDD.n2174 34.6358
R24401 VDD.n2192 VDD.n2174 34.6358
R24402 VDD.n2192 VDD.n2191 34.6358
R24403 VDD.n2211 VDD.n2167 34.6358
R24404 VDD.n2864 VDD.n2218 34.6358
R24405 VDD.n2856 VDD.n2855 34.6358
R24406 VDD.n2860 VDD.n2856 34.6358
R24407 VDD.n2812 VDD.n2811 34.6358
R24408 VDD.n2805 VDD.n2804 34.6358
R24409 VDD.n2777 VDD.n2776 34.6358
R24410 VDD.n2770 VDD.n2769 34.6358
R24411 VDD.n2771 VDD.n2770 34.6358
R24412 VDD.n2766 VDD.n2763 34.6358
R24413 VDD.n2760 VDD.n2261 34.6358
R24414 VDD.n2752 VDD.n2266 34.6358
R24415 VDD.n2688 VDD.n2687 34.6358
R24416 VDD.n2081 VDD.n1263 34.6358
R24417 VDD.n1371 VDD.n1370 34.6358
R24418 VDD.n1385 VDD.n1384 34.6358
R24419 VDD.n1400 VDD.n1399 34.6358
R24420 VDD.n1397 VDD.n1351 34.6358
R24421 VDD.n2053 VDD.n2050 34.6358
R24422 VDD.n2022 VDD.n2021 34.6358
R24423 VDD.n2017 VDD.n1420 34.6358
R24424 VDD.n2021 VDD.n1420 34.6358
R24425 VDD.n2002 VDD.n1999 34.6358
R24426 VDD.n1991 VDD.n1990 34.6358
R24427 VDD.n1992 VDD.n1991 34.6358
R24428 VDD.n1983 VDD.n1436 34.6358
R24429 VDD.n1975 VDD.n1441 34.6358
R24430 VDD.n1942 VDD.n1458 34.6358
R24431 VDD.n1903 VDD.n1901 34.6358
R24432 VDD.n1907 VDD.n1474 34.6358
R24433 VDD.n1890 VDD.n1484 34.6358
R24434 VDD.n1873 VDD.n1497 34.6358
R24435 VDD.n1863 VDD.n1500 34.6358
R24436 VDD.n1867 VDD.n1500 34.6358
R24437 VDD.n1868 VDD.n1867 34.6358
R24438 VDD.n1845 VDD.n1844 34.6358
R24439 VDD.n1841 VDD.n1840 34.6358
R24440 VDD.n1840 VDD.n1839 34.6358
R24441 VDD.n1817 VDD.n1816 34.6358
R24442 VDD.n1812 VDD.n1811 34.6358
R24443 VDD.n1801 VDD.n1531 34.6358
R24444 VDD.n1802 VDD.n1801 34.6358
R24445 VDD.n1805 VDD.n1802 34.6358
R24446 VDD.n1794 VDD.n1535 34.6358
R24447 VDD.n1708 VDD.n1707 34.6358
R24448 VDD.n1719 VDD.n1561 34.6358
R24449 VDD.n1723 VDD.n1561 34.6358
R24450 VDD.n1732 VDD.n1554 34.6358
R24451 VDD.n1756 VDD.n1548 34.6358
R24452 VDD.n1761 VDD.n1758 34.6358
R24453 VDD.n1765 VDD.n1764 34.6358
R24454 VDD.n1766 VDD.n1765 34.6358
R24455 VDD.n1771 VDD.n1770 34.6358
R24456 VDD.n1785 VDD.n1537 34.6358
R24457 VDD.n557 VDD.n556 34.6358
R24458 VDD.n561 VDD.n548 34.6358
R24459 VDD.n557 VDD.n548 34.6358
R24460 VDD.n575 VDD.n539 34.6358
R24461 VDD.n571 VDD.n539 34.6358
R24462 VDD.n1211 VDD.n1210 34.6358
R24463 VDD.n1203 VDD.n1202 34.6358
R24464 VDD.n1189 VDD.n611 34.6358
R24465 VDD.n1105 VDD.n1104 34.6358
R24466 VDD.n1091 VDD.n1090 34.6358
R24467 VDD.n1092 VDD.n1091 34.6358
R24468 VDD.n1092 VDD.n678 34.6358
R24469 VDD.n1096 VDD.n678 34.6358
R24470 VDD.n1083 VDD.n685 34.6358
R24471 VDD.n1076 VDD.n688 34.6358
R24472 VDD.n1044 VDD.n1043 34.6358
R24473 VDD.n1033 VDD.n708 34.6358
R24474 VDD.n1037 VDD.n708 34.6358
R24475 VDD.n1038 VDD.n1037 34.6358
R24476 VDD.n1030 VDD.n1029 34.6358
R24477 VDD.n986 VDD.n985 34.6358
R24478 VDD.n945 VDD.n944 34.6358
R24479 VDD.n879 VDD.n878 34.6358
R24480 VDD.n98 VDD.n91 34.6358
R24481 VDD.n4204 VDD.t565 34.4755
R24482 VDD.n2997 VDD.t1221 34.4755
R24483 VDD.n2220 VDD.t229 34.4755
R24484 VDD.n1434 VDD.t235 34.4755
R24485 VDD.n1503 VDD.t239 34.4755
R24486 VDD.n1514 VDD.t52 34.4755
R24487 VDD.n1528 VDD.t2922 34.4755
R24488 VDD.n1540 VDD.t55 34.4755
R24489 VDD.n594 VDD.t241 34.4755
R24490 VDD.n597 VDD.t233 34.4755
R24491 VDD.n638 VDD.t247 34.4755
R24492 VDD.n646 VDD.t243 34.4755
R24493 VDD.n683 VDD.t231 34.4755
R24494 VDD.n4052 VDD.t1768 34.3058
R24495 VDD.n3144 VDD.t2066 34.3058
R24496 VDD.n2271 VDD.t2127 34.3058
R24497 VDD.n2277 VDD.t2717 34.3058
R24498 VDD.n2314 VDD.t1868 34.3058
R24499 VDD.n2365 VDD.t1704 34.3058
R24500 VDD.n1416 VDD.t1092 34.3058
R24501 VDD.n1438 VDD.t646 34.3058
R24502 VDD.n1491 VDD.t1724 34.3058
R24503 VDD.n543 VDD.t1056 34.3058
R24504 VDD.n537 VDD.t2009 34.3058
R24505 VDD.n4113 VDD.n3730 34.2593
R24506 VDD.n4004 VDD.n4003 34.2593
R24507 VDD.n4405 VDD.n4404 34.2593
R24508 VDD.n3482 VDD.n2936 34.2593
R24509 VDD.n2044 VDD.n1406 34.2593
R24510 VDD.n2014 VDD.n2013 34.2593
R24511 VDD.n2006 VDD.n2005 34.2593
R24512 VDD.n1218 VDD.n1217 34.2593
R24513 VDD.n498 VDD.n497 34.2593
R24514 VDD.n3831 VDD.t969 34.0906
R24515 VDD.n3832 VDD.t2797 34.0906
R24516 VDD.n3835 VDD.t1690 34.0906
R24517 VDD.n3845 VDD.t1706 34.0906
R24518 VDD.n3846 VDD.t1139 34.0906
R24519 VDD.n4418 VDD.t2773 34.0906
R24520 VDD.n4379 VDD.t662 34.0906
R24521 VDD.n4380 VDD.t1174 34.0906
R24522 VDD.n4383 VDD.t2745 34.0906
R24523 VDD.n4388 VDD.t2090 34.0906
R24524 VDD.n3058 VDD.t2731 34.0906
R24525 VDD.n3059 VDD.t1856 34.0906
R24526 VDD.n3043 VDD.t1022 34.0906
R24527 VDD.n3065 VDD.t1079 34.0906
R24528 VDD.n3591 VDD.t1608 34.0906
R24529 VDD.n3593 VDD.t1452 34.0906
R24530 VDD.n3596 VDD.t2257 34.0906
R24531 VDD.n3597 VDD.t1598 34.0906
R24532 VDD.n2351 VDD.t2086 34.0906
R24533 VDD.n2401 VDD.t817 34.0906
R24534 VDD.n2467 VDD.t2150 34.0906
R24535 VDD.n2470 VDD.t1287 34.0906
R24536 VDD.n2472 VDD.t2727 34.0906
R24537 VDD.n2120 VDD.t1379 34.0906
R24538 VDD.n2121 VDD.t674 34.0906
R24539 VDD.n2124 VDD.t2067 34.0906
R24540 VDD.n2125 VDD.t1302 34.0906
R24541 VDD.n1580 VDD.t1456 34.0906
R24542 VDD.n1523 VDD.t1651 34.0906
R24543 VDD.n1649 VDD.t1944 34.0906
R24544 VDD.n1652 VDD.t1061 34.0906
R24545 VDD.n1654 VDD.t2074 34.0906
R24546 VDD.n1286 VDD.t989 34.0906
R24547 VDD.n1287 VDD.t734 34.0906
R24548 VDD.n1290 VDD.t882 34.0906
R24549 VDD.n1291 VDD.t1523 34.0906
R24550 VDD.n550 VDD.t876 34.0906
R24551 VDD.n588 VDD.t1257 34.0906
R24552 VDD.n606 VDD.t1643 34.0906
R24553 VDD.n625 VDD.t842 34.0906
R24554 VDD.n654 VDD.t1874 34.0906
R24555 VDD.n672 VDD.t2235 34.0906
R24556 VDD.n690 VDD.t656 34.0906
R24557 VDD.n710 VDD.t1840 34.0906
R24558 VDD.n727 VDD.t2800 34.0906
R24559 VDD.n739 VDD.t846 34.0906
R24560 VDD.n761 VDD.t2655 34.0906
R24561 VDD.n778 VDD.t668 34.0906
R24562 VDD.n779 VDD.t869 34.0906
R24563 VDD.n782 VDD.t1964 34.0906
R24564 VDD.n783 VDD.t1478 34.0906
R24565 VDD.n785 VDD.t1890 34.0906
R24566 VDD.n789 VDD.t2698 34.0906
R24567 VDD.n800 VDD.t2225 34.0906
R24568 VDD.n850 VDD.t1383 34.0906
R24569 VDD.n467 VDD.t2661 34.0906
R24570 VDD.n469 VDD.t2166 34.0906
R24571 VDD.n472 VDD.t770 34.0906
R24572 VDD.n473 VDD.t698 34.0906
R24573 VDD.n476 VDD.t2139 34.0906
R24574 VDD.n481 VDD.t890 34.0906
R24575 VDD.n4207 VDD.n4206 33.8829
R24576 VDD.n4170 VDD.n3708 33.8829
R24577 VDD.n4084 VDD.n3748 33.8829
R24578 VDD.n3429 VDD.n2963 33.8829
R24579 VDD.n3371 VDD.n2965 33.8829
R24580 VDD.n3369 VDD.n3366 33.8829
R24581 VDD.n2783 VDD.n2782 33.8829
R24582 VDD.n2592 VDD.n2591 33.8829
R24583 VDD.n2486 VDD.n2485 33.8829
R24584 VDD.n1795 VDD.n1794 33.8829
R24585 VDD.n1668 VDD.n1667 33.8829
R24586 VDD.n1196 VDD.n1195 33.8829
R24587 VDD.n1048 VDD.n703 33.8829
R24588 VDD.n867 VDD.n866 33.8829
R24589 VDD.t2945 VDD.t1565 33.5694
R24590 VDD.t2672 VDD.t571 33.5694
R24591 VDD.t1230 VDD.t1996 33.5694
R24592 VDD.t2901 VDD.t1577 33.5694
R24593 VDD.t3037 VDD.t1181 33.5694
R24594 VDD.n1779 VDD.n1778 33.5064
R24595 VDD.n4204 VDD.t739 33.4905
R24596 VDD.n2997 VDD.t1600 33.4905
R24597 VDD.n1528 VDD.t1844 33.4905
R24598 VDD.n3312 VDD.n3311 33.1299
R24599 VDD.n3554 VDD.n3553 33.1299
R24600 VDD.n2719 VDD.n2279 33.1299
R24601 VDD.n2639 VDD.n2316 33.1299
R24602 VDD.n1752 VDD.n1751 33.1299
R24603 VDD.n565 VDD.n564 33.1299
R24604 VDD.n3442 VDD.n3441 33.1299
R24605 VDD.n2490 VDD.n2468 33.1299
R24606 VDD.n1644 VDD.n1643 33.1299
R24607 VDD.n1790 VDD.n1789 33.1299
R24608 VDD.n1672 VDD.n1650 33.1299
R24609 VDD.n271 VDD.t3069 33.0605
R24610 VDD.n271 VDD.t19 33.0605
R24611 VDD.n4118 VDD.n4117 32.7534
R24612 VDD.n1379 VDD.n1378 32.7534
R24613 VDD.n1955 VDD.n1954 32.7534
R24614 VDD.n1827 VDD.n1826 32.7534
R24615 VDD.n427 VDD.n426 32.7534
R24616 VDD.n269 VDD.n268 32.6405
R24617 VDD.n4197 VDD.t1357 32.5055
R24618 VDD.n4197 VDD.t2048 32.5055
R24619 VDD.n3000 VDD.t116 32.5055
R24620 VDD.n3000 VDD.t2876 32.5055
R24621 VDD.n1526 VDD.t774 32.5055
R24622 VDD.n1526 VDD.t1044 32.5055
R24623 VDD.n3493 VDD.n3492 32.377
R24624 VDD.n3331 VDD.n2973 32.377
R24625 VDD.n3652 VDD.n3651 32.377
R24626 VDD.n3162 VDD.n3161 32.377
R24627 VDD.n3179 VDD.n3024 32.377
R24628 VDD.n2775 VDD.n2774 32.377
R24629 VDD.n2541 VDD.n2540 32.377
R24630 VDD.n1984 VDD.n1983 32.377
R24631 VDD.n1724 VDD.n1723 32.377
R24632 VDD.n1203 VDD.n603 32.377
R24633 VDD.n1084 VDD.n1083 32.377
R24634 VDD.n1039 VDD.n1038 32.377
R24635 VDD.n963 VDD.n730 32.377
R24636 VDD.n217 VDD.n189 32.2119
R24637 VDD.n4402 VDD.n4401 32.0005
R24638 VDD.n3509 VDD.n2917 32.0005
R24639 VDD.n3393 VDD.n3392 32.0005
R24640 VDD.n3166 VDD.n3029 32.0005
R24641 VDD.n3175 VDD.n3174 32.0005
R24642 VDD.n2807 VDD.n2238 32.0005
R24643 VDD.n2713 VDD.n2282 32.0005
R24644 VDD.n2633 VDD.n2319 32.0005
R24645 VDD.n1383 VDD.n1382 32.0005
R24646 VDD.n1971 VDD.n1970 32.0005
R24647 VDD.n1709 VDD.n1708 32.0005
R24648 VDD.n1766 VDD.n1543 32.0005
R24649 VDD.n552 VDD.n551 32.0005
R24650 VDD.n864 VDD.n863 32.0005
R24651 VDD.n495 VDD.n494 32.0005
R24652 VDD.n422 VDD.n421 32.0005
R24653 VDD.n1122 VDD.n1121 31.9622
R24654 VDD.t1167 VDD.t387 31.891
R24655 VDD.t177 VDD.t1246 31.891
R24656 VDD.t1945 VDD.t1440 31.891
R24657 VDD.t2116 VDD.t1773 31.891
R24658 VDD.n2025 VDD.n1417 31.624
R24659 VDD.n578 VDD.n577 31.624
R24660 VDD.n900 VDD.n755 31.624
R24661 VDD.n270 VDD.n249 31.4672
R24662 VDD.n180 VDD.t455 31.2992
R24663 VDD.n179 VDD.t451 31.2448
R24664 VDD.n180 VDD.t454 30.9042
R24665 VDD.n4401 VDD.n4389 30.8711
R24666 VDD.n494 VDD.n482 30.8711
R24667 VDD.n179 VDD.t452 30.8498
R24668 VDD.n376 VDD.n371 30.8338
R24669 VDD.n376 VDD.n375 30.8338
R24670 VDD.n385 VDD.n384 30.8338
R24671 VDD.n384 VDD.n383 30.8338
R24672 VDD.n354 VDD.n353 30.8338
R24673 VDD.n351 VDD.n349 30.8338
R24674 VDD.n863 VDD.n851 30.4946
R24675 VDD.t2251 VDD.t2250 30.2868
R24676 VDD.t2250 VDD.t2240 30.2868
R24677 VDD.t2240 VDD.t2244 30.2868
R24678 VDD.t2247 VDD.t2252 30.2868
R24679 VDD.t2252 VDD.t2246 30.2868
R24680 VDD.t2246 VDD.t2249 30.2868
R24681 VDD.t2255 VDD.t2254 30.2868
R24682 VDD.t2254 VDD.t2243 30.2868
R24683 VDD.t2243 VDD.t2241 30.2868
R24684 VDD.t409 VDD.t640 30.2125
R24685 VDD.t1526 VDD.t2593 30.2125
R24686 VDD.t1489 VDD.t1898 30.2125
R24687 VDD.t830 VDD.t1258 30.2125
R24688 VDD.t1293 VDD.t2640 30.2125
R24689 VDD.t499 VDD.t2969 30.2125
R24690 VDD.t3010 VDD.t2369 30.2125
R24691 VDD.n4110 VDD.n4109 30.1181
R24692 VDD.n943 VDD.n942 30.1181
R24693 VDD.n58 VDD.n55 30.1181
R24694 VDD.n15 VDD.n14 30.1181
R24695 VDD.n3400 VDD.n3399 30.1181
R24696 VDD.n3319 VDD.n3318 30.1181
R24697 VDD.n3547 VDD.n3546 30.1181
R24698 VDD.n3160 VDD.n3031 30.1181
R24699 VDD.n3182 VDD.n3181 30.1181
R24700 VDD.n2801 VDD.n2800 30.1181
R24701 VDD.n1391 VDD.n1390 30.1181
R24702 VDD.n1910 VDD.n1909 30.1181
R24703 VDD.n1835 VDD.n1834 30.1181
R24704 VDD.n1187 VDD.n1186 30.1181
R24705 VDD.n1066 VDD.n1065 30.1181
R24706 VDD.n3315 VDD.n3314 29.7417
R24707 VDD.n3551 VDD.n3550 29.7417
R24708 VDD.n2755 VDD.n2754 29.7417
R24709 VDD.n2017 VDD.n2016 29.7417
R24710 VDD.n562 VDD.n561 29.7417
R24711 VDD.n2953 VDD.t2027 29.5505
R24712 VDD.n2953 VDD.t420 29.5505
R24713 VDD.n313 VDD.t441 29.4286
R24714 VDD.n248 VDD.t447 29.4286
R24715 VDD.n277 VDD.t457 29.4286
R24716 VDD.n280 VDD.t437 29.4286
R24717 VDD.n284 VDD.t459 29.4286
R24718 VDD.n289 VDD.t445 29.4286
R24719 VDD.n292 VDD.t435 29.4286
R24720 VDD.n296 VDD.t449 29.4286
R24721 VDD.n301 VDD.t461 29.4286
R24722 VDD.n304 VDD.t439 29.4286
R24723 VDD.n308 VDD.t443 29.4286
R24724 VDD.n4211 VDD.n4198 29.3652
R24725 VDD.n3475 VDD.n3474 29.3652
R24726 VDD.n2625 VDD.n2327 29.3652
R24727 VDD.n1820 VDD.n1819 29.3652
R24728 VDD.n432 VDD.n410 29.3652
R24729 VDD.n3492 VDD.n2933 28.9887
R24730 VDD.n1986 VDD.n1985 28.9887
R24731 VDD.n1861 VDD.n1504 28.9887
R24732 VDD.n1777 VDD.n1539 28.9887
R24733 VDD.n1218 VDD.n595 28.9887
R24734 VDD.n1215 VDD.n598 28.9887
R24735 VDD.n1086 VDD.n1085 28.9887
R24736 VDD.n3698 VDD.t924 28.752
R24737 VDD.n4324 VDD.t1233 28.752
R24738 VDD.n2916 VDD.t2144 28.752
R24739 VDD.n2943 VDD.t1750 28.752
R24740 VDD.n3365 VDD.t1135 28.752
R24741 VDD.n2969 VDD.t2702 28.752
R24742 VDD.n2986 VDD.t1795 28.752
R24743 VDD.n3525 VDD.t811 28.752
R24744 VDD.n2176 VDD.t1936 28.752
R24745 VDD.n2206 VDD.t836 28.752
R24746 VDD.n2250 VDD.t2017 28.752
R24747 VDD.n2265 VDD.t1654 28.752
R24748 VDD.n2296 VDD.t1119 28.752
R24749 VDD.n1267 VDD.t1846 28.752
R24750 VDD.n1534 VDD.t705 28.752
R24751 VDD.n671 VDD.t902 28.752
R24752 VDD.t28 VDD.t492 28.5341
R24753 VDD.t1599 VDD.t266 28.5341
R24754 VDD.t941 VDD.t1785 28.5341
R24755 VDD.t1973 VDD.t3099 28.5341
R24756 VDD.t2831 VDD.t199 28.5341
R24757 VDD.t708 VDD.t861 28.5341
R24758 VDD.t2159 VDD.t775 28.5341
R24759 VDD.t2803 VDD.t1645 28.5341
R24760 VDD.n2348 VDD.t2029 28.5169
R24761 VDD.n3665 VDD.t676 28.4453
R24762 VDD.n2179 VDD.t1927 28.4453
R24763 VDD.n2097 VDD.t2806 28.4453
R24764 VDD.n2260 VDD.t1521 28.4453
R24765 VDD.n2293 VDD.t792 28.4453
R24766 VDD.n758 VDD.t1698 28.4453
R24767 VDD.n770 VDD.t1919 28.4453
R24768 VDD.n3710 VDD.t1277 28.4453
R24769 VDD.n4102 VDD.t1924 28.4453
R24770 VDD.n2051 VDD.t795 28.4453
R24771 VDD.n1486 VDD.t2713 28.4453
R24772 VDD.n1545 VDD.t1195 28.4453
R24773 VDD.n4176 VDD.n4175 28.2358
R24774 VDD.n3457 VDD.n3456 28.2358
R24775 VDD.n3431 VDD.n3430 28.2358
R24776 VDD.n3220 VDD.n3004 28.2358
R24777 VDD.n2144 VDD.n2118 28.2358
R24778 VDD.n1310 VDD.n1284 28.2358
R24779 VDD.n1918 VDD.n1917 28.2358
R24780 VDD.n3471 VDD.n2944 27.8593
R24781 VDD.n1958 VDD.n1957 27.8593
R24782 VDD.n1831 VDD.n1515 27.8593
R24783 VDD.n1697 VDD.n1568 27.8593
R24784 VDD.n1183 VDD.n1182 27.8593
R24785 VDD.n1012 VDD.n716 27.8593
R24786 VDD.n939 VDD.n937 27.8593
R24787 VDD.n427 VDD.n423 27.8593
R24788 VDD.n3990 VDD.n3989 27.724
R24789 VDD.n2572 VDD.n2571 27.724
R24790 VDD.n2528 VDD.n2527 27.724
R24791 VDD.n4201 VDD.t1519 27.5805
R24792 VDD.n4200 VDD.t1347 27.5805
R24793 VDD.n4200 VDD.t1345 27.5805
R24794 VDD.n4189 VDD.t900 27.5805
R24795 VDD.n4188 VDD.t1864 27.5805
R24796 VDD.n4188 VDD.t1860 27.5805
R24797 VDD.n3697 VDD.t196 27.5805
R24798 VDD.n3726 VDD.t1982 27.5805
R24799 VDD.n3706 VDD.t1554 27.5805
R24800 VDD.n3707 VDD.t1166 27.5805
R24801 VDD.n3707 VDD.t1172 27.5805
R24802 VDD.n4150 VDD.t1143 27.5805
R24803 VDD.n4150 VDD.t1147 27.5805
R24804 VDD.n3716 VDD.t85 27.5805
R24805 VDD.n3743 VDD.t1373 27.5805
R24806 VDD.n3729 VDD.t999 27.5805
R24807 VDD.n3729 VDD.t995 27.5805
R24808 VDD.n3732 VDD.t3094 27.5805
R24809 VDD.n4074 VDD.t2753 27.5805
R24810 VDD.n4074 VDD.t2755 27.5805
R24811 VDD.n3752 VDD.t77 27.5805
R24812 VDD.n3816 VDD.t156 27.5805
R24813 VDD.n4367 VDD.t896 27.5805
R24814 VDD.n4336 VDD.t805 27.5805
R24815 VDD.n4336 VDD.t801 27.5805
R24816 VDD.n4341 VDD.t1960 27.5805
R24817 VDD.n4347 VDD.t2044 27.5805
R24818 VDD.n4297 VDD.t2006 27.5805
R24819 VDD.n4297 VDD.t2004 27.5805
R24820 VDD.n4303 VDD.t1323 27.5805
R24821 VDD.n3783 VDD.t1267 27.5805
R24822 VDD.n3783 VDD.t1607 27.5805
R24823 VDD.n3789 VDD.t985 27.5805
R24824 VDD.n3789 VDD.t772 27.5805
R24825 VDD.n3944 VDD.t1429 27.5805
R24826 VDD.n3944 VDD.t2989 27.5805
R24827 VDD.n3804 VDD.t154 27.5805
R24828 VDD.n4369 VDD.t1954 27.5805
R24829 VDD.n4369 VDD.t1950 27.5805
R24830 VDD.n4384 VDD.t2050 27.5805
R24831 VDD.n4387 VDD.t1309 27.5805
R24832 VDD.n4387 VDD.t1313 27.5805
R24833 VDD.n2939 VDD.t428 27.5805
R24834 VDD.n2939 VDD.t1778 27.5805
R24835 VDD.n3348 VDD.t208 27.5805
R24836 VDD.n2989 VDD.t1046 27.5805
R24837 VDD.n2382 VDD.t1048 27.5805
R24838 VDD.n2354 VDD.t502 27.5805
R24839 VDD.n2354 VDD.t614 27.5805
R24840 VDD.n1476 VDD.t48 27.5805
R24841 VDD.n1551 VDD.t500 27.5805
R24842 VDD.n1551 VDD.t586 27.5805
R24843 VDD.n1597 VDD.t57 27.5805
R24844 VDD.n1595 VDD.t142 27.5805
R24845 VDD.n1595 VDD.t136 27.5805
R24846 VDD.n754 VDD.t1335 27.5805
R24847 VDD.n754 VDD.t506 27.5805
R24848 VDD.n762 VDD.t237 27.5805
R24849 VDD.n762 VDD.t3009 27.5805
R24850 VDD.n846 VDD.t1433 27.5805
R24851 VDD.n849 VDD.t2789 27.5805
R24852 VDD.n849 VDD.t2791 27.5805
R24853 VDD.n477 VDD.t2978 27.5805
R24854 VDD.n480 VDD.t926 27.5805
R24855 VDD.n480 VDD.t928 27.5805
R24856 VDD.n3229 VDD.n3228 27.4829
R24857 VDD.n2591 VDD.n2349 27.4829
R24858 VDD.n1810 VDD.n1809 27.4829
R24859 VDD.n902 VDD.n901 27.4829
R24860 VDD.n4089 VDD.n3744 27.4829
R24861 VDD.n3377 VDD.n3376 27.4829
R24862 VDD.n3342 VDD.n2971 27.4829
R24863 VDD.n3644 VDD.n3643 27.4829
R24864 VDD.n1780 VDD.n1537 27.4829
R24865 VDD.n1043 VDD.n706 27.4829
R24866 VDD.n3277 VDD.n3236 27.1064
R24867 VDD.n3284 VDD.n3283 27.1064
R24868 VDD.n53 VDD.n52 27.1064
R24869 VDD.n24 VDD.n23 27.1064
R24870 VDD.n4441 VDD.n4365 27.0566
R24871 VDD.n3768 VDD.t784 26.9729
R24872 VDD.t1300 VDD.t400 26.8556
R24873 VDD.n3421 VDD.t560 26.8556
R24874 VDD.t2887 VDD.t324 26.8556
R24875 VDD.t78 VDD.t1825 26.8556
R24876 VDD.t585 VDD.t2965 26.8556
R24877 VDD.t850 VDD.t103 26.8556
R24878 VDD.n2582 VDD.n2359 26.7299
R24879 VDD.n2538 VDD.n2383 26.7299
R24880 VDD.n1632 VDD.n1582 26.7299
R24881 VDD.n3776 VDD.t1281 26.5955
R24882 VDD.n2959 VDD.t1248 26.5955
R24883 VDD.n1460 VDD.t1263 26.5955
R24884 VDD.n546 VDD.t1054 26.5955
R24885 VDD.n4309 VDD.t2188 26.5955
R24886 VDD.n4309 VDD.t2190 26.5955
R24887 VDD.n3773 VDD.t1666 26.5955
R24888 VDD.n3773 VDD.t1059 26.5955
R24889 VDD.n2946 VDD.t1752 26.5955
R24890 VDD.n2946 VDD.t1754 26.5955
R24891 VDD.n3003 VDD.t1605 26.5955
R24892 VDD.n2220 VDD.t2076 26.5955
R24893 VDD.n2240 VDD.t1780 26.5955
R24894 VDD.n2240 VDD.t1774 26.5955
R24895 VDD.n2241 VDD.t245 26.5955
R24896 VDD.n2241 VDD.t1770 26.5955
R24897 VDD.n2245 VDD.t249 26.5955
R24898 VDD.n2245 VDD.t253 26.5955
R24899 VDD.n2281 VDD.t3021 26.5955
R24900 VDD.n2281 VDD.t161 26.5955
R24901 VDD.n2318 VDD.t16 26.5955
R24902 VDD.n2318 VDD.t2948 26.5955
R24903 VDD.n2614 VDD.t2816 26.5955
R24904 VDD.n2614 VDD.t1741 26.5955
R24905 VDD.n2393 VDD.t601 26.5955
R24906 VDD.n2393 VDD.t2710 26.5955
R24907 VDD.n1359 VDD.t104 26.5955
R24908 VDD.n1359 VDD.t759 26.5955
R24909 VDD.n1350 VDD.t1558 26.5955
R24910 VDD.n1350 VDD.t1562 26.5955
R24911 VDD.n1408 VDD.t332 26.5955
R24912 VDD.n1408 VDD.t1634 26.5955
R24913 VDD.n2000 VDD.t174 26.5955
R24914 VDD.n2000 VDD.t1391 26.5955
R24915 VDD.n1425 VDD.t1413 26.5955
R24916 VDD.n1425 VDD.t1407 26.5955
R24917 VDD.n1434 VDD.t1793 26.5955
R24918 VDD.n1448 VDD.t1658 26.5955
R24919 VDD.n1448 VDD.t1662 26.5955
R24920 VDD.n1473 VDD.t910 26.5955
R24921 VDD.n1473 VDD.t908 26.5955
R24922 VDD.n1496 VDD.t212 26.5955
R24923 VDD.n1496 VDD.t508 26.5955
R24924 VDD.n1503 VDD.t961 26.5955
R24925 VDD.n1514 VDD.t1484 26.5955
R24926 VDD.n1517 VDD.t1237 26.5955
R24927 VDD.n1517 VDD.t1245 26.5955
R24928 VDD.n1571 VDD.t1822 26.5955
R24929 VDD.n1571 VDD.t1818 26.5955
R24930 VDD.n1570 VDD.t1574 26.5955
R24931 VDD.n1570 VDD.t1572 26.5955
R24932 VDD.n1550 VDD.t2966 26.5955
R24933 VDD.n1550 VDD.t3098 26.5955
R24934 VDD.n1540 VDD.t709 26.5955
R24935 VDD.n1006 VDD.t1180 26.5955
R24936 VDD.n1006 VDD.t1186 26.5955
R24937 VDD.n697 VDD.t1104 26.5955
R24938 VDD.n697 VDD.t1106 26.5955
R24939 VDD.n594 VDD.t1384 26.5955
R24940 VDD.n597 VDD.t1038 26.5955
R24941 VDD.n1175 VDD.t2176 26.5955
R24942 VDD.n1175 VDD.t2178 26.5955
R24943 VDD.n638 VDD.t1972 26.5955
R24944 VDD.n646 VDD.t1933 26.5955
R24945 VDD.n683 VDD.t1639 26.5955
R24946 VDD.n929 VDD.t1911 26.5955
R24947 VDD.n929 VDD.t1913 26.5955
R24948 VDD.n415 VDD.t1730 26.5955
R24949 VDD.n415 VDD.t1726 26.5955
R24950 VDD.n424 VDD.t2771 26.5955
R24951 VDD.n424 VDD.t2928 26.5955
R24952 VDD.n416 VDD.t2767 26.5955
R24953 VDD.n416 VDD.t2765 26.5955
R24954 VDD.n411 VDD.t1714 26.5955
R24955 VDD.n411 VDD.t1716 26.5955
R24956 VDD.n92 VDD.t2088 26.5955
R24957 VDD.n48 VDD.t2761 26.5955
R24958 VDD.n48 VDD.t2759 26.5955
R24959 VDD.n54 VDD.t3043 26.5955
R24960 VDD.n54 VDD.t3049 26.5955
R24961 VDD.n22 VDD.t2719 26.5955
R24962 VDD.n22 VDD.t2725 26.5955
R24963 VDD.n19 VDD.t3045 26.5955
R24964 VDD.n19 VDD.t3055 26.5955
R24965 VDD.n2523 VDD.n2522 26.5743
R24966 VDD.n265 VDD.n264 26.4291
R24967 VDD.n266 VDD.n265 26.4291
R24968 VDD.n262 VDD.n261 26.4291
R24969 VDD.n261 VDD.n260 26.4291
R24970 VDD.n259 VDD.n249 26.4291
R24971 VDD.n260 VDD.n259 26.4291
R24972 VDD.n268 VDD.n267 26.4291
R24973 VDD.n267 VDD.n266 26.4291
R24974 VDD.n130 VDD.n129 26.4291
R24975 VDD.n131 VDD.n130 26.4291
R24976 VDD.n120 VDD.n111 26.4291
R24977 VDD.n131 VDD.n111 26.4291
R24978 VDD.n126 VDD.n112 26.4291
R24979 VDD.n131 VDD.n112 26.4291
R24980 VDD.n1355 VDD.n1354 26.3534
R24981 VDD.n1869 VDD.n1868 26.3534
R24982 VDD.n1739 VDD.n1737 26.3534
R24983 VDD.n2190 VDD.n2189 26.3037
R24984 VDD.n3257 VDD.n3243 25.977
R24985 VDD.n3270 VDD.n3238 25.977
R24986 VDD.n3198 VDD.n3017 25.977
R24987 VDD.n2214 VDD.n2165 25.977
R24988 VDD.n2685 VDD.n2294 25.977
R24989 VDD.n1637 VDD.n1636 25.977
R24990 VDD.n2009 VDD.n2008 25.977
R24991 VDD.n4047 VDD.t1766 25.6105
R24992 VDD.n2928 VDD.t922 25.6105
R24993 VDD.n3394 VDD.t936 25.6105
R24994 VDD.n3246 VDD.t1339 25.6105
R24995 VDD.n3010 VDD.t730 25.6105
R24996 VDD.n3014 VDD.t1003 25.6105
R24997 VDD.n3036 VDD.t2064 25.6105
R24998 VDD.n2205 VDD.t1836 25.6105
R24999 VDD.n2212 VDD.t1158 25.6105
R25000 VDD.n2270 VDD.t1470 25.6105
R25001 VDD.n2731 VDD.t2129 25.6105
R25002 VDD.n2278 VDD.t2715 25.6105
R25003 VDD.n2290 VDD.t958 25.6105
R25004 VDD.n2658 VDD.t2674 25.6105
R25005 VDD.n2315 VDD.t1870 25.6105
R25006 VDD.n2361 VDD.t489 25.6105
R25007 VDD.n2366 VDD.t1702 25.6105
R25008 VDD.n2385 VDD.t1680 25.6105
R25009 VDD.n1353 VDD.t1980 25.6105
R25010 VDD.n1419 VDD.t1094 25.6105
R25011 VDD.n1440 VDD.t648 25.6105
R25012 VDD.n1494 VDD.t1722 25.6105
R25013 VDD.n1788 VDD.t670 25.6105
R25014 VDD.n534 VDD.t2011 25.6105
R25015 VDD.n3869 VDD.n3868 25.6005
R25016 VDD.n3857 VDD.n3856 25.6005
R25017 VDD.n4337 VDD.n4335 25.6005
R25018 VDD.n3976 VDD.n3784 25.6005
R25019 VDD.n3395 VDD.n3393 25.6005
R25020 VDD.n3288 VDD.n3234 25.6005
R25021 VDD.n3212 VDD.n3008 25.6005
R25022 VDD.n3057 VDD.n3047 25.6005
R25023 VDD.n3614 VDD.n3594 25.6005
R25024 VDD.n3608 VDD.n3598 25.6005
R25025 VDD.n2207 VDD.n2204 25.6005
R25026 VDD.n2213 VDD.n2211 25.6005
R25027 VDD.n2741 VDD.n2738 25.6005
R25028 VDD.n2587 VDD.n2349 25.6005
R25029 VDD.n2483 VDD.n2473 25.6005
R25030 VDD.n2142 VDD.n2122 25.6005
R25031 VDD.n2136 VDD.n2126 25.6005
R25032 VDD.n1937 VDD.n1936 25.6005
R25033 VDD.n1665 VDD.n1655 25.6005
R25034 VDD.n1308 VDD.n1288 25.6005
R25035 VDD.n1302 VDD.n1292 25.6005
R25036 VDD.n1100 VDD.n1099 25.6005
R25037 VDD.n1070 VDD.n691 25.6005
R25038 VDD.n841 VDD.n776 25.6005
R25039 VDD.n3617 VDD.n3616 25.5028
R25040 VDD.n4205 VDD.n3696 25.224
R25041 VDD.n4225 VDD.n4190 25.224
R25042 VDD.n4225 VDD.n4224 25.224
R25043 VDD.n4177 VDD.n4176 25.224
R25044 VDD.n4177 VDD.n3701 25.224
R25045 VDD.n4172 VDD.n4171 25.224
R25046 VDD.n4305 VDD.n4304 25.224
R25047 VDD.n4409 VDD.n4385 25.224
R25048 VDD.n3430 VDD.n3429 25.224
R25049 VDD.n3219 VDD.n3218 25.224
R25050 VDD.n3220 VDD.n3219 25.224
R25051 VDD.n3205 VDD.n3204 25.224
R25052 VDD.n2151 VDD.n2115 25.224
R25053 VDD.n2151 VDD.n2150 25.224
R25054 VDD.n2149 VDD.n2148 25.224
R25055 VDD.n2148 VDD.n2118 25.224
R25056 VDD.n1315 VDD.n1314 25.224
R25057 VDD.n1314 VDD.n1284 25.224
R25058 VDD.n825 VDD.n790 25.224
R25059 VDD.n871 VDD.n847 25.224
R25060 VDD.n872 VDD.n871 25.224
R25061 VDD.n502 VDD.n478 25.224
R25062 VDD.n59 VDD.n58 25.224
R25063 VDD.n20 VDD.n14 25.224
R25064 VDD.n4084 VDD.n4083 25.1912
R25065 VDD.n4056 VDD.n4054 25.1912
R25066 VDD.n3974 VDD.n3787 25.1912
R25067 VDD.n3413 VDD.n3350 25.1912
R25068 VDD.n3249 VDD.n2993 25.1912
R25069 VDD.n3257 VDD.n3256 25.1912
R25070 VDD.n3198 VDD.n3197 25.1912
R25071 VDD.n3151 VDD.n3034 25.1912
R25072 VDD.n2786 VDD.n2783 25.1912
R25073 VDD.n2724 VDD.n2721 25.1912
R25074 VDD.n2710 VDD.n2709 25.1912
R25075 VDD.n2069 VDD.n1264 25.1912
R25076 VDD.n2032 VDD.n2030 25.1912
R25077 VDD.n1970 VDD.n1969 25.1912
R25078 VDD.n1936 VDD.n1461 25.1912
R25079 VDD.n1181 VDD.n1180 25.1912
R25080 VDD.n1168 VDD.n1165 25.1912
R25081 VDD.n1165 VDD.n1164 25.1912
R25082 VDD.n1138 VDD.n655 25.1912
R25083 VDD.n978 VDD.n728 25.1912
R25084 VDD.n961 VDD.n733 25.1912
R25085 VDD.n3873 VDD.n3833 24.8476
R25086 VDD.n3861 VDD.n3847 24.8476
R25087 VDD.n4417 VDD.n4416 24.8476
R25088 VDD.n4415 VDD.n4381 24.8476
R25089 VDD.n4411 VDD.n4410 24.8476
R25090 VDD.n3451 VDD.n3450 24.8476
R25091 VDD.n3402 VDD.n3354 24.8476
R25092 VDD.n3308 VDD.n3307 24.8476
R25093 VDD.n3558 VDD.n3557 24.8476
R25094 VDD.n3061 VDD.n3060 24.8476
R25095 VDD.n3616 VDD.n3615 24.8476
R25096 VDD.n3610 VDD.n3609 24.8476
R25097 VDD.n2797 VDD.n2246 24.8476
R25098 VDD.n2748 VDD.n2746 24.8476
R25099 VDD.n2714 VDD.n2713 24.8476
R25100 VDD.n2634 VDD.n2633 24.8476
R25101 VDD.n2587 VDD.n2586 24.8476
R25102 VDD.n2485 VDD.n2484 24.8476
R25103 VDD.n2144 VDD.n2143 24.8476
R25104 VDD.n2138 VDD.n2137 24.8476
R25105 VDD.n1812 VDD.n1524 24.8476
R25106 VDD.n1667 VDD.n1666 24.8476
R25107 VDD.n1310 VDD.n1309 24.8476
R25108 VDD.n1304 VDD.n1303 24.8476
R25109 VDD.n569 VDD.n541 24.8476
R25110 VDD.n1228 VDD.n589 24.8476
R25111 VDD.n1202 VDD.n1201 24.8476
R25112 VDD.n1139 VDD.n1138 24.8476
R25113 VDD.n1104 VDD.n673 24.8476
R25114 VDD.n979 VDD.n978 24.8476
R25115 VDD.n888 VDD.n887 24.8476
R25116 VDD.n840 VDD.n839 24.8476
R25117 VDD.n832 VDD.n786 24.8476
R25118 VDD.n826 VDD.n825 24.8476
R25119 VDD.n514 VDD.n470 24.8476
R25120 VDD.n510 VDD.n509 24.8476
R25121 VDD.n508 VDD.n474 24.8476
R25122 VDD.n504 VDD.n503 24.8476
R25123 VDD.n2598 VDD.n2597 24.5135
R25124 VDD.n1079 VDD.n685 24.4711
R25125 VDD.n982 VDD.n980 24.4711
R25126 VDD.n906 VDD.n752 24.4711
R25127 VDD.n901 VDD.n900 24.4711
R25128 VDD.n1250 VDD.n1249 24.4382
R25129 VDD.n935 VDD.n934 24.4382
R25130 VDD.n1108 VDD.n1106 24.4382
R25131 VDD.n1063 VDD.n695 24.1679
R25132 VDD.n3862 VDD.n3861 24.0946
R25133 VDD.n4054 VDD.n4053 24.0946
R25134 VDD.n3306 VDD.n2987 24.0946
R25135 VDD.n3153 VDD.n3152 24.0946
R25136 VDD.n3187 VDD.n3186 24.0946
R25137 VDD.n3610 VDD.n3594 24.0946
R25138 VDD.n2737 VDD.n2272 24.0946
R25139 VDD.n2721 VDD.n2720 24.0946
R25140 VDD.n2630 VDD.n2629 24.0946
R25141 VDD.n2138 VDD.n2122 24.0946
R25142 VDD.n1371 VDD.n1364 24.0946
R25143 VDD.n1979 VDD.n1436 24.0946
R25144 VDD.n1878 VDD.n1877 24.0946
R25145 VDD.n1304 VDD.n1288 24.0946
R25146 VDD.n839 VDD.n780 24.0946
R25147 VDD.n833 VDD.n832 24.0946
R25148 VDD.n515 VDD.n514 24.0946
R25149 VDD.n4011 VDD.n3769 23.7483
R25150 VDD.n4362 VDD.n3677 23.7181
R25151 VDD.n2715 VDD.n2714 23.7181
R25152 VDD.n2635 VDD.n2634 23.7181
R25153 VDD.n2621 VDD.n2620 23.7181
R25154 VDD.n2057 VDD.n2056 23.7181
R25155 VDD.n1895 VDD.n1891 23.7181
R25156 VDD.n876 VDD.n774 23.7181
R25157 VDD.n4252 VDD.n3696 23.7181
R25158 VDD.n4124 VDD.n3727 23.7181
R25159 VDD.n4098 VDD.n3741 23.7181
R25160 VDD.n3913 VDD.n3814 23.7181
R25161 VDD.n3916 VDD.n3913 23.7181
R25162 VDD.n3874 VDD.n3873 23.7181
R25163 VDD.n4305 VDD.n3677 23.7181
R25164 VDD.n4008 VDD.n3771 23.7181
R25165 VDD.n4004 VDD.n3771 23.7181
R25166 VDD.n3995 VDD.n3994 23.7181
R25167 VDD.n3982 VDD.n3981 23.7181
R25168 VDD.n4442 VDD.n4441 23.7181
R25169 VDD.n3572 VDD.n2912 23.7181
R25170 VDD.n3500 VDD.n3499 23.7181
R25171 VDD.n3479 VDD.n2940 23.7181
R25172 VDD.n3424 VDD.n2965 23.7181
R25173 VDD.n3420 VDD.n2967 23.7181
R25174 VDD.n3297 VDD.n2993 23.7181
R25175 VDD.n3294 VDD.n2994 23.7181
R25176 VDD.n3572 VDD.n2913 23.7181
R25177 VDD.n3202 VDD.n3017 23.7181
R25178 VDD.n3061 VDD.n3045 23.7181
R25179 VDD.n3638 VDD.n3637 23.7181
R25180 VDD.n2865 VDD.n2864 23.7181
R25181 VDD.n2756 VDD.n2261 23.7181
R25182 VDD.n2756 VDD.n2755 23.7181
R25183 VDD.n2745 VDD.n2268 23.7181
R25184 VDD.n2583 VDD.n2582 23.7181
R25185 VDD.n1996 VDD.n1429 23.7181
R25186 VDD.n1992 VDD.n1429 23.7181
R25187 VDD.n1891 VDD.n1890 23.7181
R25188 VDD.n1752 VDD.n1749 23.7181
R25189 VDD.n1229 VDD.n1228 23.7181
R25190 VDD.n1223 VDD.n1222 23.7181
R25191 VDD.n1189 VDD.n1188 23.7181
R25192 VDD.n1050 VDD.n1049 23.7181
R25193 VDD.n1049 VDD.n1048 23.7181
R25194 VDD.n907 VDD.n906 23.7181
R25195 VDD.n166 VDD.n165 23.7181
R25196 VDD.t2041 VDD.t2538 23.4987
R25197 VDD.t2482 VDD.t168 23.4987
R25198 VDD.t329 VDD.t1853 23.4987
R25199 VDD.t36 VDD.t744 23.4987
R25200 VDD.t884 VDD.t92 23.4987
R25201 VDD.n175 VDD.t150 23.3739
R25202 VDD.t147 VDD.n171 23.3739
R25203 VDD.n151 VDD.t2940 23.3739
R25204 VDD.n155 VDD.t2938 23.3739
R25205 VDD.n3439 VDD.n3438 23.3417
R25206 VDD.n2626 VDD.n2625 23.3417
R25207 VDD.n1375 VDD.n1364 23.3417
R25208 VDD.n2025 VDD.n2024 23.3417
R25209 VDD.n1900 VDD.n1899 23.3417
R25210 VDD.n1879 VDD.n1878 23.3417
R25211 VDD.n1844 VDD.n1509 23.3417
R25212 VDD.n555 VDD.n554 23.3417
R25213 VDD.n1195 VDD.n1194 23.3417
R25214 VDD.n256 VDD.n255 23.1255
R25215 VDD.n257 VDD.n250 23.1255
R25216 VDD.n258 VDD.n257 23.1255
R25217 VDD.n253 VDD.n251 23.1255
R25218 VDD.n323 VDD.n322 22.9976
R25219 VDD.n4397 VDD.n4396 22.9652
R25220 VDD.n1674 VDD.n1577 22.9652
R25221 VDD.n859 VDD.n858 22.9652
R25222 VDD.n490 VDD.n489 22.9652
R25223 VDD.n3997 VDD.n3996 22.9652
R25224 VDD.n3947 VDD.n3946 22.9652
R25225 VDD.n3495 VDD.n2929 22.9652
R25226 VDD.n3480 VDD.n3479 22.9652
R25227 VDD.n3344 VDD.n3343 22.9652
R25228 VDD.n3263 VDD.n3262 22.9652
R25229 VDD.n3268 VDD.n3241 22.9652
R25230 VDD.n3290 VDD.n3289 22.9652
R25231 VDD.n3564 VDD.n3523 22.9652
R25232 VDD.n3642 VDD.n3575 22.9652
R25233 VDD.n2777 VDD.n2252 22.9652
R25234 VDD.n2571 VDD.n2363 22.9652
R25235 VDD.n2527 VDD.n2387 22.9652
R25236 VDD.n2081 VDD.n2080 22.9652
R25237 VDD.n1362 VDD.n1360 22.9652
R25238 VDD.n2043 VDD.n2042 22.9652
R25239 VDD.n1943 VDD.n1942 22.9652
R25240 VDD.n1883 VDD.n1489 22.9652
R25241 VDD.n1809 VDD.n1529 22.9652
R25242 VDD.n1729 VDD.n1558 22.9652
R25243 VDD.n1743 VDD.n1552 22.9652
R25244 VDD.n1787 VDD.n1785 22.9652
R25245 VDD.n1233 VDD.n1232 22.9652
R25246 VDD.n2038 VDD.n2037 22.9323
R25247 VDD.n1857 VDD.n1856 22.9323
R25248 VDD.n1238 VDD.n1237 22.9323
R25249 VDD.t2242 VDD.n218 22.842
R25250 VDD.t2249 VDD.n216 22.842
R25251 VDD.n218 VDD.t2251 22.842
R25252 VDD.n216 VDD.t2255 22.842
R25253 VDD.t61 VDD.n348 22.742
R25254 VDD.n3395 VDD.n3356 22.5887
R25255 VDD.n3225 VDD.n3224 22.5887
R25256 VDD.n3212 VDD.n3211 22.5887
R25257 VDD.n2207 VDD.n2167 22.5887
R25258 VDD.n2214 VDD.n2213 22.5887
R25259 VDD.n2738 VDD.n2737 22.5887
R25260 VDD.n2692 VDD.n2691 22.5887
R25261 VDD.n4125 VDD.n4124 22.2123
R25262 VDD.n4010 VDD.n4008 22.2123
R25263 VDD.n4011 VDD.n4010 22.2123
R25264 VDD.n3981 VDD.n3784 22.2123
R25265 VDD.n3976 VDD.n3975 22.2123
R25266 VDD.n3975 VDD.n3974 22.2123
R25267 VDD.n3947 VDD.n3805 22.2123
R25268 VDD.n3302 VDD.n3301 22.2123
R25269 VDD.n3301 VDD.n3300 22.2123
R25270 VDD.n2860 VDD.n2859 22.2123
R25271 VDD.n1797 VDD.n1531 22.2123
R25272 VDD.n1797 VDD.n1796 22.2123
R25273 VDD.n1736 VDD.n1554 22.2123
R25274 VDD.n1233 VDD.n451 22.2123
R25275 VDD.n1072 VDD.n1071 22.2123
R25276 VDD.n963 VDD.n962 22.2123
R25277 VDD.n962 VDD.n961 22.2123
R25278 VDD.n883 VDD.n882 22.2123
R25279 VDD.n2733 VDD.n2732 22.0294
R25280 VDD.n578 VDD.n535 22.0294
R25281 VDD.n4419 VDD.n4417 22.0015
R25282 VDD.n408 VDD.n394 22.0005
R25283 VDD.n3467 VDD.n3466 21.8358
R25284 VDD.n1398 VDD.n1397 21.8358
R25285 VDD.n2005 VDD.n1426 21.8358
R25286 VDD.n1954 VDD.n1449 21.8358
R25287 VDD.n1826 VDD.n1825 21.8358
R25288 VDD.n1692 VDD.n1691 21.8358
R25289 VDD.n1694 VDD.n1693 21.8358
R25290 VDD.n420 VDD.n417 21.8358
R25291 VDD.t2079 VDD.t1376 21.8203
R25292 VDD.t1923 VDD.t2080 21.8203
R25293 VDD.t1788 VDD.t547 21.8203
R25294 VDD.t2690 VDD.t2688 21.8203
R25295 VDD.t1547 VDD.n2263 21.8203
R25296 VDD.t835 VDD.t336 21.8203
R25297 VDD.t911 VDD.t1049 21.8203
R25298 VDD.t909 VDD.t1224 21.8203
R25299 VDD.t482 VDD.t812 21.8203
R25300 VDD.n3994 VDD.n3780 21.4593
R25301 VDD.n3990 VDD.n3780 21.4593
R25302 VDD.n3499 VDD.n2929 21.4593
R25303 VDD.n3488 VDD.n2933 21.4593
R25304 VDD.n3451 VDD.n2951 21.4593
R25305 VDD.n3344 VDD.n2967 21.4593
R25306 VDD.n3307 VDD.n3306 21.4593
R25307 VDD.n3264 VDD.n3241 21.4593
R25308 VDD.n3290 VDD.n2994 21.4593
R25309 VDD.n3560 VDD.n3523 21.4593
R25310 VDD.n3559 VDD.n3558 21.4593
R25311 VDD.n3230 VDD.n2995 21.4593
R25312 VDD.n3203 VDD.n3202 21.4593
R25313 VDD.n3152 VDD.n3151 21.4593
R25314 VDD.n3154 VDD.n3031 21.4593
R25315 VDD.n3182 VDD.n3022 21.4593
R25316 VDD.n3638 VDD.n3575 21.4593
R25317 VDD.n2855 VDD.n2221 21.4593
R25318 VDD.n2781 VDD.n2252 21.4593
R25319 VDD.n2746 VDD.n2745 21.4593
R25320 VDD.n2523 VDD.n2387 21.4593
R25321 VDD.n2080 VDD.n1264 21.4593
R25322 VDD.n1392 VDD.n1391 21.4593
R25323 VDD.n2044 VDD.n2043 21.4593
R25324 VDD.n2013 VDD.n1423 21.4593
R25325 VDD.n1986 VDD.n1432 21.4593
R25326 VDD.n1916 VDD.n1469 21.4593
R25327 VDD.n1862 VDD.n1861 21.4593
R25328 VDD.n1700 VDD.n1699 21.4593
R25329 VDD.n1732 VDD.n1731 21.4593
R25330 VDD.n1737 VDD.n1736 21.4593
R25331 VDD.n1778 VDD.n1777 21.4593
R25332 VDD.n1790 VDD.n1787 21.4593
R25333 VDD.n565 VDD.n545 21.4593
R25334 VDD.n1222 VDD.n595 21.4593
R25335 VDD.n1210 VDD.n1209 21.4593
R25336 VDD.n1211 VDD.n598 21.4593
R25337 VDD.n1186 VDD.n616 21.4593
R25338 VDD.n1086 VDD.n681 21.4593
R25339 VDD.n1065 VDD.n1064 21.4593
R25340 VDD.n892 VDD.n759 21.4593
R25341 VDD.n888 VDD.n759 21.4593
R25342 VDD.n991 VDD.n987 21.1483
R25343 VDD.n1990 VDD.n1432 21.0829
R25344 VDD.n1875 VDD.n1874 21.0829
R25345 VDD.n1863 VDD.n1862 21.0829
R25346 VDD.n1839 VDD.n1511 21.0829
R25347 VDD.n1749 VDD.n1744 21.0829
R25348 VDD.n1090 VDD.n681 21.0829
R25349 VDD.n1008 VDD.n1007 20.9397
R25350 VDD.n2578 VDD.n2359 20.824
R25351 VDD.n2534 VDD.n2383 20.824
R25352 VDD.n4206 VDD.n4205 20.7064
R25353 VDD.n4171 VDD.n4170 20.7064
R25354 VDD.n4342 VDD.n4340 20.7064
R25355 VDD.n4405 VDD.n4385 20.7064
R25356 VDD.n867 VDD.n847 20.7064
R25357 VDD.n498 VDD.n478 20.7064
R25358 VDD.n60 VDD.n59 20.7064
R25359 VDD.n21 VDD.n20 20.7064
R25360 VDD.n228 VDD.n225 20.5561
R25361 VDD.n228 VDD.n219 20.5561
R25362 VDD.n174 VDD.n173 20.5174
R25363 VDD.n172 VDD.n89 20.5174
R25364 VDD.n153 VDD.n152 20.5174
R25365 VDD.n154 VDD.n104 20.5174
R25366 VDD.n1119 VDD.n667 20.4852
R25367 VDD.n4109 VDD.n4108 20.3299
R25368 VDD.n3447 VDD.n3446 20.3299
R25369 VDD.n3399 VDD.n3356 20.3299
R25370 VDD.n2150 VDD.n2149 20.3299
R25371 VDD.n1938 VDD.n1937 20.3299
R25372 VDD.n1707 VDD.n1566 20.3299
R25373 VDD.n944 VDD.n943 20.3299
R25374 VDD.n4334 VDD.n4321 20.2801
R25375 VDD.t1288 VDD.t1671 20.1418
R25376 VDD.t101 VDD.t1011 20.1418
R25377 VDD.t2126 VDD.t2230 20.1418
R25378 VDD.t871 VDD.t1520 20.1418
R25379 VDD.t171 VDD.t1360 20.1418
R25380 VDD.n4212 VDD.n4211 19.9534
R25381 VDD.n4165 VDD.n4164 19.9534
R25382 VDD.n4119 VDD.n4118 19.9534
R25383 VDD.n4094 VDD.n4093 19.9534
R25384 VDD.n4335 VDD.n4334 19.9534
R25385 VDD.n3416 VDD.n2966 19.9534
R25386 VDD.n3302 VDD.n2987 19.9534
R25387 VDD.n3217 VDD.n3216 19.9534
R25388 VDD.n2628 VDD.n2627 19.9534
R25389 VDD.n2541 VDD.n2380 19.9534
R25390 VDD.n571 VDD.n570 19.9534
R25391 VDD.n1208 VDD.n1207 19.9534
R25392 VDD.n1079 VDD.n1078 19.9534
R25393 VDD.n985 VDD.n724 19.9534
R25394 VDD.n945 VDD.n735 19.9534
R25395 VDD.n902 VDD.n752 19.9534
R25396 VDD.n896 VDD.n895 19.9534
R25397 VDD.t61 VDD.n357 19.8857
R25398 VDD.n359 VDD.n350 19.828
R25399 VDD.n360 VDD.n359 19.828
R25400 VDD.n418 VDD.n417 19.6052
R25401 VDD.n3869 VDD.n3833 19.577
R25402 VDD.n3857 VDD.n3847 19.577
R25403 VDD.n4416 VDD.n4415 19.577
R25404 VDD.n4411 VDD.n4381 19.577
R25405 VDD.n4410 VDD.n4409 19.577
R25406 VDD.n3060 VDD.n3057 19.577
R25407 VDD.n3615 VDD.n3614 19.577
R25408 VDD.n3609 VDD.n3608 19.577
R25409 VDD.n2491 VDD.n2490 19.577
R25410 VDD.n2484 VDD.n2483 19.577
R25411 VDD.n2143 VDD.n2142 19.577
R25412 VDD.n2137 VDD.n2136 19.577
R25413 VDD.n1643 VDD.n1642 19.577
R25414 VDD.n1385 VDD.n1357 19.577
R25415 VDD.n2042 VDD.n1411 19.577
R25416 VDD.n1869 VDD.n1497 19.577
R25417 VDD.n1816 VDD.n1524 19.577
R25418 VDD.n1673 VDD.n1672 19.577
R25419 VDD.n1666 VDD.n1665 19.577
R25420 VDD.n1309 VDD.n1308 19.577
R25421 VDD.n1303 VDD.n1302 19.577
R25422 VDD.n1201 VDD.n1200 19.577
R25423 VDD.n1100 VDD.n673 19.577
R25424 VDD.n1071 VDD.n1070 19.577
R25425 VDD.n841 VDD.n840 19.577
R25426 VDD.n510 VDD.n470 19.577
R25427 VDD.n509 VDD.n508 19.577
R25428 VDD.n504 VDD.n474 19.577
R25429 VDD.n503 VDD.n502 19.577
R25430 VDD.n388 VDD.n387 19.4467
R25431 VDD.n387 VDD.n386 19.4467
R25432 VDD.n4112 VDD.n4111 19.2005
R25433 VDD.n3448 VDD.n3447 19.2005
R25434 VDD.n516 VDD.n515 19.2005
R25435 VDD.n1025 VDD.n712 18.9442
R25436 VDD.n1316 VDD.n1315 18.88
R25437 VDD.n4166 VDD.n4165 18.824
R25438 VDD.n3481 VDD.n3480 18.824
R25439 VDD.n2806 VDD.n2805 18.824
R25440 VDD.n2763 VDD.n2762 18.824
R25441 VDD.n1638 VDD.n1579 18.824
R25442 VDD.n2053 VDD.n2052 18.824
R25443 VDD.n1949 VDD.n1948 18.824
R25444 VDD.n1903 VDD.n1902 18.824
R25445 VDD.n1820 VDD.n1520 18.824
R25446 VDD.n1687 VDD.n1572 18.824
R25447 VDD.n938 VDD.n740 18.824
R25448 VDD.n878 VDD.n877 18.824
R25449 VDD.n806 VDD.n805 18.7912
R25450 VDD.n1051 VDD.n1050 18.6667
R25451 VDD.t1861 VDD.t2631 18.4634
R25452 VDD.t1344 VDD.t2047 18.4634
R25453 VDD.t993 VDD.t1445 18.4634
R25454 VDD.t1385 VDD.t1125 18.4634
R25455 VDD.t2409 VDD.t2007 18.4634
R25456 VDD.t1834 VDD.t1157 18.4634
R25457 VDD.t1200 VDD.t1499 18.4634
R25458 VDD.n3517 VDD.n3516 18.4476
R25459 VDD.n3487 VDD.n3486 18.4476
R25460 VDD.n3434 VDD.n3433 18.4476
R25461 VDD.n3270 VDD.n3269 18.4476
R25462 VDD.n3275 VDD.n3274 18.4476
R25463 VDD.n1642 VDD.n1579 18.4476
R25464 VDD.n1376 VDD.n1375 18.4476
R25465 VDD.n2030 VDD.n2029 18.4476
R25466 VDD.n1978 VDD.n1977 18.4476
R25467 VDD.n1773 VDD.n1772 18.4476
R25468 VDD.n1251 VDD.n445 18.4476
R25469 VDD.n1200 VDD.n608 18.4476
R25470 VDD.n895 VDD.n894 18.4476
R25471 VDD.n4213 VDD.n4212 18.4147
R25472 VDD.n168 VDD.n162 18.2003
R25473 VDD.n3494 VDD.n3493 18.0711
R25474 VDD.n3335 VDD.n2973 18.0711
R25475 VDD.n3651 VDD.n3650 18.0711
R25476 VDD.n2776 VDD.n2775 18.0711
R25477 VDD.n2733 VDD.n2272 18.0711
R25478 VDD.n2720 VDD.n2719 18.0711
R25479 VDD.n2640 VDD.n2639 18.0711
R25480 VDD.n1368 VDD.n1263 18.0711
R25481 VDD.n2049 VDD.n2048 18.0711
R25482 VDD.n1979 VDD.n1978 18.0711
R25483 VDD.n1938 VDD.n1458 18.0711
R25484 VDD.n1886 VDD.n1885 18.0711
R25485 VDD.n1725 VDD.n1558 18.0711
R25486 VDD.n1207 VDD.n603 18.0711
R25487 VDD.n3320 VDD.n3319 17.6946
R25488 VDD.n3546 VDD.n3545 17.6946
R25489 VDD.n2799 VDD.n2798 17.6946
R25490 VDD.n2461 VDD.n2460 17.6946
R25491 VDD.n2460 VDD.n2459 17.6946
R25492 VDD.n1833 VDD.n1832 17.6946
R25493 VDD.n4361 VDD.n4360 17.6618
R25494 VDD.n4024 VDD.n4023 17.612
R25495 VDD.n2825 VDD.n2823 17.612
R25496 VDD.n2661 VDD.n2657 17.612
R25497 VDD.n102 VDD.n101 17.5829
R25498 VDD.n4172 VDD.n3704 17.3181
R25499 VDD.n4175 VDD.n3704 17.3181
R25500 VDD.n4340 VDD.n4319 17.3181
R25501 VDD.n3507 VDD.n2920 17.3181
R25502 VDD.n3461 VDD.n3460 17.3181
R25503 VDD.n3362 VDD.n3359 17.3181
R25504 VDD.n3388 VDD.n3362 17.3181
R25505 VDD.n3415 VDD.n3414 17.3181
R25506 VDD.n3414 VDD.n3413 17.3181
R25507 VDD.n3300 VDD.n2991 17.3181
R25508 VDD.n3281 VDD.n3236 17.3181
R25509 VDD.n3284 VDD.n3234 17.3181
R25510 VDD.n3566 VDD.n3565 17.3181
R25511 VDD.n2172 VDD.n2169 17.3181
R25512 VDD.n2199 VDD.n2172 17.3181
R25513 VDD.n2198 VDD.n2197 17.3181
R25514 VDD.n2197 VDD.n2196 17.3181
R25515 VDD.n2771 VDD.n2256 17.3181
R25516 VDD.n2774 VDD.n2256 17.3181
R25517 VDD.n2741 VDD.n2740 17.3181
R25518 VDD.n2492 VDD.n2399 17.3181
R25519 VDD.n2458 VDD.n2457 17.3181
R25520 VDD.n1370 VDD.n1369 17.3181
R25521 VDD.n1805 VDD.n1804 17.3181
R25522 VDD.n1097 VDD.n1096 17.3181
R25523 VDD.n4224 VDD.n4223 17.2853
R25524 VDD.n4350 VDD.n4349 17.2853
R25525 VDD.n2155 VDD.n2115 17.2853
R25526 VDD.n521 VDD.n465 17.2853
R25527 VDD.n2620 VDD.n2619 16.9977
R25528 VDD.n4119 VDD.n3727 16.9417
R25529 VDD.n1948 VDD.n1455 16.9417
R25530 VDD.n1811 VDD.n1810 16.9417
R25531 VDD.n382 VDD.t2766 16.7855
R25532 VDD.n381 VDD.t2764 16.7855
R25533 VDD.n380 VDD.t2770 16.7855
R25534 VDD.n379 VDD.t2927 16.7855
R25535 VDD.t1084 VDD.t1955 16.785
R25536 VDD.t1312 VDD.t2089 16.785
R25537 VDD.t54 VDD.t1878 16.785
R25538 VDD.t1262 VDD.t1534 16.785
R25539 VDD.t2022 VDD.t945 16.785
R25540 VDD.t2788 VDD.t1382 16.785
R25541 VDD.t1963 VDD.t1477 16.785
R25542 VDD.t1994 VDD.t2069 16.785
R25543 VDD.t927 VDD.t889 16.785
R25544 VDD.n201 VDD.t2919 16.7806
R25545 VDD.n1120 VDD.n1119 16.7729
R25546 VDD.n3425 VDD.n3424 16.5652
R25547 VDD.n3218 VDD.n3217 16.5652
R25548 VDD.n1153 VDD.n1152 16.5652
R25549 VDD.n828 VDD.n827 16.5652
R25550 VDD.n2645 VDD.n2644 16.4179
R25551 VDD.n3486 VDD.n3485 16.1887
R25552 VDD.n3433 VDD.n2960 16.1887
R25553 VDD.n2766 VDD.n2765 16.1887
R25554 VDD.n1631 VDD.n1630 16.1887
R25555 VDD.n1377 VDD.n1376 16.1887
R25556 VDD.n2029 VDD.n2028 16.1887
R25557 VDD.n1951 VDD.n1950 16.1887
R25558 VDD.n1893 VDD.n1477 16.1887
R25559 VDD.n1894 VDD.n1893 16.1887
R25560 VDD.n1824 VDD.n1823 16.1887
R25561 VDD.n1772 VDD.n1771 16.1887
R25562 VDD.n551 VDD.n445 16.1887
R25563 VDD.n1197 VDD.n608 16.1887
R25564 VDD.n1031 VDD.n1030 16.1887
R25565 VDD.n2694 VDD.n2692 16.1559
R25566 VDD.n3130 VDD.n3129 16.139
R25567 VDD.n3909 VDD.n3814 15.8683
R25568 VDD.n4443 VDD.n4442 15.8683
R25569 VDD.n4048 VDD.n4046 15.8683
R25570 VDD.n2869 VDD.n2868 15.8683
R25571 VDD.n2681 VDD.n2294 15.8683
R25572 VDD.n4249 VDD.n3701 15.8123
R25573 VDD.n4167 VDD.n4166 15.8123
R25574 VDD.n3459 VDD.n2947 15.8123
R25575 VDD.n2807 VDD.n2806 15.8123
R25576 VDD.n2459 VDD.n2458 15.8123
R25577 VDD.n1632 VDD.n1631 15.8123
R25578 VDD.n1638 VDD.n1637 15.8123
R25579 VDD.n1400 VDD.n1349 15.8123
R25580 VDD.n1999 VDD.n1998 15.8123
R25581 VDD.n1950 VDD.n1949 15.8123
R25582 VDD.n1902 VDD.n1474 15.8123
R25583 VDD.n1823 VDD.n1520 15.8123
R25584 VDD.n1687 VDD.n1686 15.8123
R25585 VDD.n1690 VDD.n1572 15.8123
R25586 VDD.n1703 VDD.n1566 15.8123
R25587 VDD.n1725 VDD.n1724 15.8123
R25588 VDD.n1764 VDD.n1546 15.8123
R25589 VDD.n1032 VDD.n1031 15.8123
R25590 VDD.n835 VDD.n780 15.8123
R25591 VDD.n834 VDD.n833 15.8123
R25592 VDD.n877 VDD.n876 15.8123
R25593 VDD.n873 VDD.n872 15.8123
R25594 VDD.n2814 VDD.n2812 15.606
R25595 VDD.n3516 VDD.n3515 15.4358
R25596 VDD.n3227 VDD.n3226 15.4358
R25597 VDD.n2462 VDD.n2399 15.4358
R25598 VDD.n2052 VDD.n1404 15.4358
R25599 VDD.n1998 VDD.n1997 15.4358
R25600 VDD.n517 VDD.n465 15.4358
R25601 VDD.n4127 VDD.n4126 15.3731
R25602 VDD.n1121 VDD.n666 15.2281
R25603 VDD.n2374 VDD.n2373 15.1657
R25604 VDD.n456 VDD.n455 15.1657
R25605 VDD.t404 VDD.t2703 15.1065
R25606 VDD.t2220 VDD.t808 15.1065
R25607 VDD.t1234 VDD.t977 15.1065
R25608 VDD.t816 VDD.t274 15.1065
R25609 VDD.t2807 VDD.t2008 15.1065
R25610 VDD.t542 VDD.t2660 15.1065
R25611 VDD.n2594 VDD.n2593 15.0593
R25612 VDD.n1369 VDD.n1368 15.0593
R25613 VDD.n949 VDD.n735 15.0265
R25614 VDD.n3637 VDD.n3636 14.9
R25615 VDD.n820 VDD.n794 14.7513
R25616 VDD.n64 VDD.n63 14.7184
R25617 VDD.n42 VDD.n28 14.7184
R25618 VDD.n4099 VDD.n4098 14.6829
R25619 VDD.n2769 VDD.n2258 14.6829
R25620 VDD.n4343 VDD.n4342 14.6829
R25621 VDD.n2048 VDD.n2047 14.6829
R25622 VDD.n1977 VDD.n1976 14.6829
R25623 VDD.n1912 VDD.n1911 14.6829
R25624 VDD.n897 VDD.n896 14.6829
R25625 VDD.n886 VDD.n885 14.6829
R25626 VDD.n3954 VDD.n3953 14.65
R25627 VDD.n2545 VDD.n2380 14.65
R25628 VDD.n2373 VDD.n2372 14.4912
R25629 VDD.n457 VDD.n456 14.4912
R25630 VDD.n74 VDD.n73 14.4822
R25631 VDD.n37 VDD.n36 14.4822
R25632 VDD.n3996 VDD.n3995 14.3064
R25633 VDD.n2851 VDD.n2221 14.3064
R25634 VDD.n792 VDD.n790 14.3064
R25635 VDD.n805 VDD.n774 14.3064
R25636 VDD.n4138 VDD.n4137 14.2735
R25637 VDD.n4070 VDD.n3753 14.2735
R25638 VDD.n4254 VDD.n4252 14.2735
R25639 VDD.n4270 VDD.n4265 14.2735
R25640 VDD.n3137 VDD.n3135 14.2735
R25641 VDD.n1229 VDD.n530 14.2735
R25642 VDD.n1144 VDD.n1143 14.2735
R25643 VDD.n924 VDD.n744 14.2735
R25644 VDD.n920 VDD.n744 14.2735
R25645 VDD.n188 VDD.n183 14.2313
R25646 VDD.n206 VDD.n192 14.2313
R25647 VDD.n213 VDD.n194 14.2313
R25648 VDD.n194 VDD.n190 14.2313
R25649 VDD.n211 VDD.n210 14.2313
R25650 VDD.n210 VDD.n187 14.2313
R25651 VDD.n2060 VDD.n1346 14.2027
R25652 VDD.n4060 VDD.n3753 14.1392
R25653 VDD.n2555 VDD.n2554 14.1211
R25654 VDD.n3867 VDD.n3836 13.9299
R25655 VDD.n2492 VDD.n2491 13.9299
R25656 VDD.n1760 VDD.n1546 13.9299
R25657 VDD.n1674 VDD.n1673 13.9299
R25658 VDD.n981 VDD.n724 13.9299
R25659 VDD.n635 VDD.n634 13.6608
R25660 VDD.n4343 VDD.n4316 13.5534
R25661 VDD.n1224 VDD.n1223 13.5534
R25662 VDD.t1310 VDD.t2091 13.4281
R25663 VDD.t3065 VDD.t467 13.4281
R25664 VDD.t2947 VDD.t785 13.4281
R25665 VDD.t2949 VDD.t1010 13.4281
R25666 VDD.t160 VDD.t786 13.4281
R25667 VDD.t158 VDD.t532 13.4281
R25668 VDD.t2373 VDD.t2117 13.4281
R25669 VDD.t515 VDD.t1122 13.4281
R25670 VDD.t638 VDD.t763 13.4281
R25671 VDD.t111 VDD.t2951 13.4281
R25672 VDD.t2648 VDD.t310 13.4281
R25673 VDD.t1821 VDD.t1569 13.4281
R25674 VDD.t1817 VDD.t1573 13.4281
R25675 VDD.t1819 VDD.t1571 13.4281
R25676 VDD.t569 VDD.t1072 13.4281
R25677 VDD.t2781 VDD.t1575 13.4281
R25678 VDD.t1358 VDD.t1883 13.4281
R25679 VDD.t2385 VDD.t1612 13.4281
R25680 VDD.t696 VDD.t217 13.4281
R25681 VDD.t2662 VDD.t211 13.4281
R25682 VDD.t511 VDD.t507 13.4281
R25683 VDD.t2784 VDD.t1380 13.4281
R25684 VDD.t3095 VDD.n723 13.4281
R25685 VDD.t426 VDD.t1398 13.4281
R25686 VDD.t429 VDD.t232 13.4281
R25687 VDD.t240 VDD.t433 13.4281
R25688 VDD.t931 VDD.t887 13.4281
R25689 VDD.t3048 VDD.t826 13.4281
R25690 VDD.t3052 VDD.t824 13.4281
R25691 VDD.t3056 VDD.t1318 13.4281
R25692 VDD.t3044 VDD.t1316 13.4281
R25693 VDD.n389 VDD.n388 13.2148
R25694 VDD.n344 VDD.n333 13.2148
R25695 VDD.n344 VDD.n339 13.2148
R25696 VDD.n360 VDD.n347 13.2148
R25697 VDD.n4113 VDD.n4112 13.177
R25698 VDD.n4094 VDD.n3741 13.177
R25699 VDD.n3868 VDD.n3867 13.177
R25700 VDD.n3863 VDD.n3862 13.177
R25701 VDD.n4003 VDD.n4002 13.177
R25702 VDD.n3420 VDD.n2966 13.177
R25703 VDD.n3155 VDD.n3154 13.177
R25704 VDD.n3185 VDD.n3022 13.177
R25705 VDD.n2798 VDD.n2797 13.177
R25706 VDD.n2641 VDD.n2640 13.177
R25707 VDD.n2585 VDD.n2584 13.177
R25708 VDD.n2584 VDD.n2583 13.177
R25709 VDD.n1393 VDD.n1392 13.177
R25710 VDD.n2010 VDD.n1423 13.177
R25711 VDD.n1913 VDD.n1469 13.177
R25712 VDD.n1913 VDD.n1912 13.177
R25713 VDD.n1832 VDD.n1831 13.177
R25714 VDD.n1183 VDD.n616 13.177
R25715 VDD.n1142 VDD.n1141 13.177
R25716 VDD.n1099 VDD.n1098 13.177
R25717 VDD.n1064 VDD.n1063 13.177
R25718 VDD.n939 VDD.n938 13.177
R25719 VDD.n884 VDD.n883 13.177
R25720 VDD.n873 VDD.n776 13.177
R25721 VDD.n1685 VDD.n1684 12.9693
R25722 VDD.n4304 VDD.n4302 12.8565
R25723 VDD.n4249 VDD.n3700 12.8005
R25724 VDD.n3875 VDD.n3874 12.8005
R25725 VDD.n4348 VDD.n4316 12.8005
R25726 VDD.n4349 VDD.n4348 12.8005
R25727 VDD.n3466 VDD.n3465 12.8005
R25728 VDD.n3131 VDD.n3045 12.8005
R25729 VDD.n3131 VDD.n3130 12.8005
R25730 VDD.n2868 VDD.n2164 12.8005
R25731 VDD.n2865 VDD.n2165 12.8005
R25732 VDD.n2642 VDD.n2641 12.8005
R25733 VDD.n2595 VDD.n2594 12.8005
R25734 VDD.n2593 VDD.n2592 12.8005
R25735 VDD.n2556 VDD.n2555 12.8005
R25736 VDD.n2060 VDD.n1342 12.8005
R25737 VDD.n1399 VDD.n1398 12.8005
R25738 VDD.n2057 VDD.n1347 12.8005
R25739 VDD.n1944 VDD.n1455 12.8005
R25740 VDD.n1944 VDD.n1943 12.8005
R25741 VDD.n1908 VDD.n1907 12.8005
R25742 VDD.n1691 VDD.n1690 12.8005
R25743 VDD.n1693 VDD.n1692 12.8005
R25744 VDD.n1209 VDD.n1208 12.8005
R25745 VDD.n1143 VDD.n1142 12.8005
R25746 VDD.n3945 VDD.n3943 12.5826
R25747 VDD.n2108 VDD.n2107 12.4487
R25748 VDD.n3503 VDD.n2920 12.424
R25749 VDD.n1141 VDD.n1140 12.424
R25750 VDD.n3294 VDD.n2995 12.0476
R25751 VDD.n1390 VDD.n1357 12.0476
R25752 VDD.n3406 VDD.n3354 12.0147
R25753 VDD.n3190 VDD.n3187 12.0147
R25754 VDD.n2793 VDD.n2246 12.0147
R25755 VDD.n204 VDD.n203 11.7586
R25756 VDD.t2467 VDD.t1144 11.7496
R25757 VDD.t2018 VDD.t899 11.7496
R25758 VDD.t1322 VDD.t2098 11.7496
R25759 VDD.t2118 VDD.t1015 11.7496
R25760 VDD.t1066 VDD.t622 11.7496
R25761 VDD.t596 VDD.t913 11.7496
R25762 VDD.t2202 VDD.t2691 11.7496
R25763 VDD.t1885 VDD.t920 11.7496
R25764 VDD.t1886 VDD.t2780 11.7496
R25765 VDD.t2868 VDD.t1432 11.7496
R25766 VDD.n885 VDD.n884 11.6711
R25767 VDD.n1151 VDD.n1150 11.6382
R25768 VDD.n235 VDD.n234 11.4643
R25769 VDD.n4101 VDD.n4100 11.2946
R25770 VDD.n3440 VDD.n3439 11.2946
R25771 VDD.n3204 VDD.n3203 11.2946
R25772 VDD.n2859 VDD.n2858 11.2946
R25773 VDD.n2851 VDD.n2850 11.2946
R25774 VDD.n2761 VDD.n2760 11.2946
R25775 VDD.n1382 VDD.n1360 11.2946
R25776 VDD.n1901 VDD.n1900 11.2946
R25777 VDD.n1841 VDD.n1509 11.2946
R25778 VDD.n556 VDD.n555 11.2946
R25779 VDD.n570 VDD.n569 11.2946
R25780 VDD.n1194 VDD.n1193 11.2946
R25781 VDD.n4229 VDD.n4190 11.2618
R25782 VDD.n1275 VDD.n1274 11.1615
R25783 VDD.n73 VDD.t2055 11.1031
R25784 VDD.n36 VDD.t583 11.1031
R25785 VDD.n80 VDD.n79 10.969
R25786 VDD.n44 VDD.n43 10.9682
R25787 VDD.n2567 VDD.n2363 10.9181
R25788 VDD.n1879 VDD.n1489 10.9181
R25789 VDD.n1876 VDD.n1875 10.9181
R25790 VDD.n1919 VDD.n1918 10.8853
R25791 VDD.n158 VDD.n157 10.8443
R25792 VDD.n3984 VDD.n3983 10.7794
R25793 VDD.n2643 VDD.n2642 10.5744
R25794 VDD.n2556 VDD.n2375 10.5744
R25795 VDD.n528 VDD.n453 10.5744
R25796 VDD.n133 VDD.n132 10.5561
R25797 VDD.n3456 VDD.n3455 10.5417
R25798 VDD.n3262 VDD.n3243 10.5417
R25799 VDD.n2801 VDD.n2242 10.5417
R25800 VDD.n1232 VDD.n528 10.5417
R25801 VDD.n1154 VDD.n1153 10.5417
R25802 VDD.n100 VDD.n99 10.5417
R25803 VDD.n101 VDD.n100 10.5417
R25804 VDD.n2596 VDD.n2595 10.4607
R25805 VDD.n57 VDD.n56 10.1732
R25806 VDD.n17 VDD.n16 10.1732
R25807 VDD.n3567 VDD.n3566 10.1652
R25808 VDD.n3211 VDD.n3210 10.1652
R25809 VDD.n2462 VDD.n2461 10.1652
R25810 VDD.n1349 VDD.n1347 10.1652
R25811 VDD.n2001 VDD.n1426 10.1652
R25812 VDD.n1804 VDD.n1529 10.1652
R25813 VDD.n545 VDD.n544 10.1652
R25814 VDD.n517 VDD.n516 10.1652
R25815 VDD.n272 VDD.n270 10.1337
R25816 VDD.t2553 VDD.t398 10.0712
R25817 VDD.t1114 VDD.t2431 10.0712
R25818 VDD.t2108 VDD.t2406 10.0712
R25819 VDD.t2746 VDD.t2049 10.0712
R25820 VDD.t1482 VDD.t544 10.0712
R25821 VDD.t1759 VDD.t628 10.0712
R25822 VDD.t1742 VDD.t1751 10.0712
R25823 VDD.t318 VDD.t1621 10.0712
R25824 VDD.t1807 VDD.t1669 10.0712
R25825 VDD.t633 VDD.t1071 10.0712
R25826 VDD.t1988 VDD.t53 10.0712
R25827 VDD.t513 VDD.t1721 10.0712
R25828 VDD.t2699 VDD.t1891 10.0712
R25829 VDD.t1030 VDD.t2695 10.0712
R25830 VDD.t2654 VDD.t3008 10.0712
R25831 VDD.t123 VDD.t1371 10.0712
R25832 VDD.t2563 VDD.t1368 10.0712
R25833 VDD.n676 VDD.t986 10.0712
R25834 VDD.t3012 VDD.t2979 10.0712
R25835 VDD.t607 VDD.t2732 10.0712
R25836 VDD.t2140 VDD.t2977 10.0712
R25837 VDD.t2131 VDD.t2686 10.0712
R25838 VDD.n3106 VDD.n3105 9.8812
R25839 VDD.n3952 VDD.n3805 9.78874
R25840 VDD.n2804 VDD.n2242 9.78874
R25841 VDD.n2038 VDD.n1411 9.78874
R25842 VDD.n2024 VDD.n2023 9.78874
R25843 VDD.n1731 VDD.n1729 9.78874
R25844 VDD.n1066 VDD.n691 9.78874
R25845 VDD.n60 VDD.n53 9.78874
R25846 VDD.n24 VDD.n21 9.78874
R25847 VDD.n4144 VDD.n4143 9.73273
R25848 VDD.n4148 VDD.n4147 9.73273
R25849 VDD.n4156 VDD.n3714 9.73273
R25850 VDD.n4159 VDD.n4158 9.73273
R25851 VDD.n3905 VDD.n3817 9.73273
R25852 VDD.n3906 VDD.n3905 9.73273
R25853 VDD.n4330 VDD.n4329 9.73273
R25854 VDD.n4461 VDD.n3664 9.73273
R25855 VDD.n4459 VDD.n3666 9.73273
R25856 VDD.n4449 VDD.n4448 9.73273
R25857 VDD.n4277 VDD.n4276 9.73273
R25858 VDD.n4299 VDD.n4296 9.73273
R25859 VDD.n4044 VDD.n3760 9.73273
R25860 VDD.n3934 VDD.n3810 9.73273
R25861 VDD.n3935 VDD.n3934 9.73273
R25862 VDD.n3937 VDD.n3935 9.73273
R25863 VDD.n3941 VDD.n3808 9.73273
R25864 VDD.n4435 VDD.n4434 9.73273
R25865 VDD.n4431 VDD.n4430 9.73273
R25866 VDD.n4430 VDD.n4429 9.73273
R25867 VDD.n4429 VDD.n4373 9.73273
R25868 VDD.n4425 VDD.n4373 9.73273
R25869 VDD.n4425 VDD.n4424 9.73273
R25870 VDD.n4424 VDD.n4423 9.73273
R25871 VDD.n2186 VDD.n2185 9.73273
R25872 VDD.n2886 VDD.n2885 9.73273
R25873 VDD.n2885 VDD.n2094 9.73273
R25874 VDD.n2875 VDD.n2874 9.73273
R25875 VDD.n2829 VDD.n2828 9.73273
R25876 VDD.n2832 VDD.n2829 9.73273
R25877 VDD.n2665 VDD.n2302 9.73273
R25878 VDD.n2666 VDD.n2665 9.73273
R25879 VDD.n2672 VDD.n2671 9.73273
R25880 VDD.n2673 VDD.n2672 9.73273
R25881 VDD.n2673 VDD.n2297 9.73273
R25882 VDD.n2677 VDD.n2297 9.73273
R25883 VDD.n2678 VDD.n2677 9.73273
R25884 VDD.n2611 VDD.n2332 9.73273
R25885 VDD.n2616 VDD.n2613 9.73273
R25886 VDD.n2504 VDD.n2501 9.73273
R25887 VDD.n2508 VDD.n2507 9.73273
R25888 VDD.n2516 VDD.n2515 9.73273
R25889 VDD.n2496 VDD.n2495 9.73273
R25890 VDD.n1604 VDD.n1593 9.73273
R25891 VDD.n1598 VDD.n1576 9.73273
R25892 VDD.n1677 VDD.n1576 9.73273
R25893 VDD.n1323 VDD.n1322 9.73273
R25894 VDD.n3107 VDD.n3106 9.65664
R25895 VDD.n4152 VDD.n4151 9.62695
R25896 VDD.n3936 VDD.n3808 9.62695
R25897 VDD.n4437 VDD.n4436 9.62695
R25898 VDD.n2510 VDD.n2391 9.62695
R25899 VDD.n2516 VDD.n2389 9.62695
R25900 VDD.n455 VDD.n454 9.6005
R25901 VDD.n4328 VDD.n4327 9.52116
R25902 VDD.n4447 VDD.n4446 9.52116
R25903 VDD.n1600 VDD.n1596 9.52116
R25904 VDD.n1325 VDD.n1279 9.52116
R25905 VDD.n1319 VDD.n1281 9.52116
R25906 VDD.n2597 VDD.n2337 9.49727
R25907 VDD.n3513 VDD.n2917 9.41227
R25908 VDD.n3482 VDD.n3481 9.41227
R25909 VDD.n3475 VDD.n2940 9.41227
R25910 VDD.n3392 VDD.n3359 9.41227
R25911 VDD.n3328 VDD.n2976 9.41227
R25912 VDD.n3321 VDD.n3320 9.41227
R25913 VDD.n3545 VDD.n3544 9.41227
R25914 VDD.n3540 VDD.n3539 9.41227
R25915 VDD.n3167 VDD.n3166 9.41227
R25916 VDD.n3174 VDD.n3173 9.41227
R25917 VDD.n2811 VDD.n2238 9.41227
R25918 VDD.n2688 VDD.n2291 9.41227
R25919 VDD.n1971 VDD.n1441 9.41227
R25920 VDD.n1885 VDD.n1884 9.41227
R25921 VDD.n1713 VDD.n1563 9.41227
R25922 VDD.n1770 VDD.n1543 9.41227
R25923 VDD.n1188 VDD.n1187 9.41227
R25924 VDD.n1072 VDD.n688 9.41227
R25925 VDD.n879 VDD.n768 9.41227
R25926 VDD.n989 VDD.n988 9.38145
R25927 VDD.n1325 VDD.n1324 9.30959
R25928 VDD.n4239 VDD.n4238 9.30183
R25929 VDD.n660 VDD.n659 9.30183
R25930 VDD.n3858 VDD.n3857 9.3005
R25931 VDD.n3859 VDD.n3847 9.3005
R25932 VDD.n3861 VDD.n3860 9.3005
R25933 VDD.n3862 VDD.n3843 9.3005
R25934 VDD.n3864 VDD.n3863 9.3005
R25935 VDD.n3865 VDD.n3836 9.3005
R25936 VDD.n3867 VDD.n3866 9.3005
R25937 VDD.n3868 VDD.n3834 9.3005
R25938 VDD.n3870 VDD.n3869 9.3005
R25939 VDD.n3871 VDD.n3833 9.3005
R25940 VDD.n3873 VDD.n3872 9.3005
R25941 VDD.n3881 VDD.n3880 9.3005
R25942 VDD.n3882 VDD.n3823 9.3005
R25943 VDD.n3884 VDD.n3883 9.3005
R25944 VDD.n3886 VDD.n3822 9.3005
R25945 VDD.n3889 VDD.n3888 9.3005
R25946 VDD.n3891 VDD.n3890 9.3005
R25947 VDD.n3892 VDD.n3820 9.3005
R25948 VDD.n3895 VDD.n3894 9.3005
R25949 VDD.n3896 VDD.n3819 9.3005
R25950 VDD.n3898 VDD.n3897 9.3005
R25951 VDD.n3899 VDD.n3818 9.3005
R25952 VDD.n3902 VDD.n3901 9.3005
R25953 VDD.n3903 VDD.n3817 9.3005
R25954 VDD.n3905 VDD.n3904 9.3005
R25955 VDD.n3906 VDD.n3815 9.3005
R25956 VDD.n3910 VDD.n3909 9.3005
R25957 VDD.n3911 VDD.n3814 9.3005
R25958 VDD.n3913 VDD.n3912 9.3005
R25959 VDD.n3922 VDD.n3921 9.3005
R25960 VDD.n3923 VDD.n3812 9.3005
R25961 VDD.n3925 VDD.n3924 9.3005
R25962 VDD.n3927 VDD.n3811 9.3005
R25963 VDD.n3931 VDD.n3930 9.3005
R25964 VDD.n3932 VDD.n3810 9.3005
R25965 VDD.n3934 VDD.n3933 9.3005
R25966 VDD.n3935 VDD.n3809 9.3005
R25967 VDD.n3938 VDD.n3937 9.3005
R25968 VDD.n3939 VDD.n3808 9.3005
R25969 VDD.n3941 VDD.n3940 9.3005
R25970 VDD.n3807 VDD.n3806 9.3005
R25971 VDD.n3948 VDD.n3947 9.3005
R25972 VDD.n3949 VDD.n3805 9.3005
R25973 VDD.n3952 VDD.n3950 9.3005
R25974 VDD.n3953 VDD.n3803 9.3005
R25975 VDD.n3955 VDD.n3954 9.3005
R25976 VDD.n3957 VDD.n3956 9.3005
R25977 VDD.n3958 VDD.n3801 9.3005
R25978 VDD.n3961 VDD.n3960 9.3005
R25979 VDD.n3966 VDD.n3965 9.3005
R25980 VDD.n3967 VDD.n3788 9.3005
R25981 VDD.n3971 VDD.n3970 9.3005
R25982 VDD.n3972 VDD.n3787 9.3005
R25983 VDD.n3974 VDD.n3973 9.3005
R25984 VDD.n3975 VDD.n3785 9.3005
R25985 VDD.n3977 VDD.n3976 9.3005
R25986 VDD.n3978 VDD.n3784 9.3005
R25987 VDD.n3981 VDD.n3980 9.3005
R25988 VDD.n3979 VDD.n3782 9.3005
R25989 VDD.n3989 VDD.n3781 9.3005
R25990 VDD.n3991 VDD.n3990 9.3005
R25991 VDD.n3992 VDD.n3780 9.3005
R25992 VDD.n3994 VDD.n3993 9.3005
R25993 VDD.n3995 VDD.n3778 9.3005
R25994 VDD.n3996 VDD.n3777 9.3005
R25995 VDD.n3997 VDD.n3775 9.3005
R25996 VDD.n3999 VDD.n3998 9.3005
R25997 VDD.n4000 VDD.n3774 9.3005
R25998 VDD.n4002 VDD.n4001 9.3005
R25999 VDD.n4003 VDD.n3772 9.3005
R26000 VDD.n4005 VDD.n4004 9.3005
R26001 VDD.n4006 VDD.n3771 9.3005
R26002 VDD.n4008 VDD.n4007 9.3005
R26003 VDD.n4010 VDD.n3770 9.3005
R26004 VDD.n4012 VDD.n4011 9.3005
R26005 VDD.n4014 VDD.n4013 9.3005
R26006 VDD.n4017 VDD.n3767 9.3005
R26007 VDD.n4021 VDD.n4020 9.3005
R26008 VDD.n4023 VDD.n4022 9.3005
R26009 VDD.n4024 VDD.n3765 9.3005
R26010 VDD.n4027 VDD.n4026 9.3005
R26011 VDD.n4029 VDD.n4028 9.3005
R26012 VDD.n4031 VDD.n3763 9.3005
R26013 VDD.n4034 VDD.n4033 9.3005
R26014 VDD.n4035 VDD.n3762 9.3005
R26015 VDD.n4037 VDD.n4036 9.3005
R26016 VDD.n4038 VDD.n3761 9.3005
R26017 VDD.n4041 VDD.n4040 9.3005
R26018 VDD.n4042 VDD.n3760 9.3005
R26019 VDD.n4044 VDD.n4043 9.3005
R26020 VDD.n4046 VDD.n3759 9.3005
R26021 VDD.n4049 VDD.n4048 9.3005
R26022 VDD.n4050 VDD.n3758 9.3005
R26023 VDD.n4053 VDD.n4051 9.3005
R26024 VDD.n4054 VDD.n3756 9.3005
R26025 VDD.n4057 VDD.n4056 9.3005
R26026 VDD.n4059 VDD.n4058 9.3005
R26027 VDD.n4064 VDD.n3754 9.3005
R26028 VDD.n4067 VDD.n4066 9.3005
R26029 VDD.n4068 VDD.n3753 9.3005
R26030 VDD.n4070 VDD.n4069 9.3005
R26031 VDD.n4072 VDD.n3751 9.3005
R26032 VDD.n4077 VDD.n4076 9.3005
R26033 VDD.n4078 VDD.n3750 9.3005
R26034 VDD.n4080 VDD.n4079 9.3005
R26035 VDD.n4083 VDD.n3749 9.3005
R26036 VDD.n4085 VDD.n4084 9.3005
R26037 VDD.n4087 VDD.n4086 9.3005
R26038 VDD.n4088 VDD.n3745 9.3005
R26039 VDD.n4090 VDD.n4089 9.3005
R26040 VDD.n4092 VDD.n4091 9.3005
R26041 VDD.n4093 VDD.n3742 9.3005
R26042 VDD.n4095 VDD.n4094 9.3005
R26043 VDD.n4098 VDD.n4097 9.3005
R26044 VDD.n4101 VDD.n3736 9.3005
R26045 VDD.n4105 VDD.n4104 9.3005
R26046 VDD.n4106 VDD.n3735 9.3005
R26047 VDD.n4108 VDD.n4107 9.3005
R26048 VDD.n4109 VDD.n3733 9.3005
R26049 VDD.n4110 VDD.n3731 9.3005
R26050 VDD.n4114 VDD.n4113 9.3005
R26051 VDD.n4116 VDD.n4115 9.3005
R26052 VDD.n4118 VDD.n3728 9.3005
R26053 VDD.n4120 VDD.n4119 9.3005
R26054 VDD.n4121 VDD.n3727 9.3005
R26055 VDD.n4124 VDD.n4123 9.3005
R26056 VDD.n4122 VDD.n3725 9.3005
R26057 VDD.n4130 VDD.n3724 9.3005
R26058 VDD.n4133 VDD.n4132 9.3005
R26059 VDD.n4137 VDD.n4136 9.3005
R26060 VDD.n4135 VDD.n3722 9.3005
R26061 VDD.n4134 VDD.n3719 9.3005
R26062 VDD.n4143 VDD.n3718 9.3005
R26063 VDD.n4145 VDD.n4144 9.3005
R26064 VDD.n4147 VDD.n4146 9.3005
R26065 VDD.n4148 VDD.n3715 9.3005
R26066 VDD.n4153 VDD.n4152 9.3005
R26067 VDD.n4154 VDD.n3714 9.3005
R26068 VDD.n4156 VDD.n4155 9.3005
R26069 VDD.n4158 VDD.n3713 9.3005
R26070 VDD.n4160 VDD.n4159 9.3005
R26071 VDD.n4162 VDD.n4161 9.3005
R26072 VDD.n4164 VDD.n3711 9.3005
R26073 VDD.n4165 VDD.n3709 9.3005
R26074 VDD.n4168 VDD.n4167 9.3005
R26075 VDD.n4170 VDD.n4169 9.3005
R26076 VDD.n4171 VDD.n3705 9.3005
R26077 VDD.n4173 VDD.n4172 9.3005
R26078 VDD.n4175 VDD.n4174 9.3005
R26079 VDD.n4176 VDD.n3702 9.3005
R26080 VDD.n4178 VDD.n4177 9.3005
R26081 VDD.n4179 VDD.n3701 9.3005
R26082 VDD.n4249 VDD.n4248 9.3005
R26083 VDD.n4246 VDD.n4245 9.3005
R26084 VDD.n4243 VDD.n4180 9.3005
R26085 VDD.n4236 VDD.n4235 9.3005
R26086 VDD.n4234 VDD.n4233 9.3005
R26087 VDD.n4232 VDD.n4187 9.3005
R26088 VDD.n4229 VDD.n4228 9.3005
R26089 VDD.n4227 VDD.n4190 9.3005
R26090 VDD.n4226 VDD.n4225 9.3005
R26091 VDD.n4224 VDD.n4191 9.3005
R26092 VDD.n4223 VDD.n4222 9.3005
R26093 VDD.n4221 VDD.n4220 9.3005
R26094 VDD.n4219 VDD.n4193 9.3005
R26095 VDD.n4217 VDD.n4216 9.3005
R26096 VDD.n4215 VDD.n4194 9.3005
R26097 VDD.n4214 VDD.n4213 9.3005
R26098 VDD.n4212 VDD.n4195 9.3005
R26099 VDD.n4211 VDD.n4210 9.3005
R26100 VDD.n4209 VDD.n4208 9.3005
R26101 VDD.n4206 VDD.n4199 9.3005
R26102 VDD.n4205 VDD.n4203 9.3005
R26103 VDD.n4202 VDD.n3696 9.3005
R26104 VDD.n4252 VDD.n3695 9.3005
R26105 VDD.n4255 VDD.n4254 9.3005
R26106 VDD.n4256 VDD.n3694 9.3005
R26107 VDD.n4258 VDD.n4257 9.3005
R26108 VDD.n4259 VDD.n3690 9.3005
R26109 VDD.n4263 VDD.n4262 9.3005
R26110 VDD.n4265 VDD.n4264 9.3005
R26111 VDD.n4271 VDD.n3688 9.3005
R26112 VDD.n4274 VDD.n4273 9.3005
R26113 VDD.n4276 VDD.n4275 9.3005
R26114 VDD.n4277 VDD.n3686 9.3005
R26115 VDD.n4280 VDD.n4279 9.3005
R26116 VDD.n4282 VDD.n4281 9.3005
R26117 VDD.n4283 VDD.n3684 9.3005
R26118 VDD.n4285 VDD.n4284 9.3005
R26119 VDD.n4287 VDD.n4286 9.3005
R26120 VDD.n4288 VDD.n3682 9.3005
R26121 VDD.n4291 VDD.n4290 9.3005
R26122 VDD.n4292 VDD.n3681 9.3005
R26123 VDD.n4294 VDD.n4293 9.3005
R26124 VDD.n4296 VDD.n3680 9.3005
R26125 VDD.n4300 VDD.n4299 9.3005
R26126 VDD.n4302 VDD.n4301 9.3005
R26127 VDD.n4304 VDD.n3678 9.3005
R26128 VDD.n4306 VDD.n4305 9.3005
R26129 VDD.n4362 VDD.n4308 9.3005
R26130 VDD.n4360 VDD.n4359 9.3005
R26131 VDD.n4358 VDD.n4357 9.3005
R26132 VDD.n4355 VDD.n4311 9.3005
R26133 VDD.n4354 VDD.n4353 9.3005
R26134 VDD.n4352 VDD.n4313 9.3005
R26135 VDD.n4351 VDD.n4350 9.3005
R26136 VDD.n4349 VDD.n4314 9.3005
R26137 VDD.n4348 VDD.n4346 9.3005
R26138 VDD.n4345 VDD.n4316 9.3005
R26139 VDD.n4344 VDD.n4343 9.3005
R26140 VDD.n4342 VDD.n4317 9.3005
R26141 VDD.n4340 VDD.n4339 9.3005
R26142 VDD.n4338 VDD.n4337 9.3005
R26143 VDD.n4335 VDD.n4320 9.3005
R26144 VDD.n4334 VDD.n4333 9.3005
R26145 VDD.n4332 VDD.n4321 9.3005
R26146 VDD.n4331 VDD.n4330 9.3005
R26147 VDD.n4329 VDD.n4322 9.3005
R26148 VDD.n4327 VDD.n4326 9.3005
R26149 VDD.n3664 VDD.n3662 9.3005
R26150 VDD.n4462 VDD.n4461 9.3005
R26151 VDD.n4459 VDD.n4458 9.3005
R26152 VDD.n4451 VDD.n3666 9.3005
R26153 VDD.n4450 VDD.n4449 9.3005
R26154 VDD.n4448 VDD.n3668 9.3005
R26155 VDD.n4446 VDD.n4445 9.3005
R26156 VDD.n4444 VDD.n4443 9.3005
R26157 VDD.n4442 VDD.n3671 9.3005
R26158 VDD.n4441 VDD.n4440 9.3005
R26159 VDD.n4439 VDD.n4365 9.3005
R26160 VDD.n4438 VDD.n4437 9.3005
R26161 VDD.n4435 VDD.n4366 9.3005
R26162 VDD.n4434 VDD.n4433 9.3005
R26163 VDD.n4432 VDD.n4431 9.3005
R26164 VDD.n4430 VDD.n4371 9.3005
R26165 VDD.n4429 VDD.n4428 9.3005
R26166 VDD.n4427 VDD.n4373 9.3005
R26167 VDD.n4426 VDD.n4425 9.3005
R26168 VDD.n4424 VDD.n4374 9.3005
R26169 VDD.n4423 VDD.n4422 9.3005
R26170 VDD.n4421 VDD.n4420 9.3005
R26171 VDD.n4417 VDD.n4377 9.3005
R26172 VDD.n4416 VDD.n4378 9.3005
R26173 VDD.n4415 VDD.n4414 9.3005
R26174 VDD.n4413 VDD.n4381 9.3005
R26175 VDD.n4412 VDD.n4411 9.3005
R26176 VDD.n4410 VDD.n4382 9.3005
R26177 VDD.n4409 VDD.n4408 9.3005
R26178 VDD.n4407 VDD.n4385 9.3005
R26179 VDD.n4406 VDD.n4405 9.3005
R26180 VDD.n4403 VDD.n4386 9.3005
R26181 VDD.n4401 VDD.n4400 9.3005
R26182 VDD.n4399 VDD.n4398 9.3005
R26183 VDD.n3057 VDD.n3056 9.3005
R26184 VDD.n3060 VDD.n3046 9.3005
R26185 VDD.n3062 VDD.n3061 9.3005
R26186 VDD.n3131 VDD.n3064 9.3005
R26187 VDD.n3129 VDD.n3128 9.3005
R26188 VDD.n3127 VDD.n3126 9.3005
R26189 VDD.n3124 VDD.n3072 9.3005
R26190 VDD.n3123 VDD.n3122 9.3005
R26191 VDD.n3121 VDD.n3120 9.3005
R26192 VDD.n3118 VDD.n3074 9.3005
R26193 VDD.n3117 VDD.n3116 9.3005
R26194 VDD.n3115 VDD.n3075 9.3005
R26195 VDD.n3114 VDD.n3113 9.3005
R26196 VDD.n3112 VDD.n3076 9.3005
R26197 VDD.n3111 VDD.n3110 9.3005
R26198 VDD.n3109 VDD.n3108 9.3005
R26199 VDD.n3106 VDD.n3078 9.3005
R26200 VDD.n3104 VDD.n3103 9.3005
R26201 VDD.n3102 VDD.n3101 9.3005
R26202 VDD.n3100 VDD.n3080 9.3005
R26203 VDD.n3098 VDD.n3097 9.3005
R26204 VDD.n3096 VDD.n3095 9.3005
R26205 VDD.n3094 VDD.n3082 9.3005
R26206 VDD.n3093 VDD.n3092 9.3005
R26207 VDD.n3091 VDD.n3083 9.3005
R26208 VDD.n3090 VDD.n3089 9.3005
R26209 VDD.n3088 VDD.n3084 9.3005
R26210 VDD.n3086 VDD.n3085 9.3005
R26211 VDD.n3135 VDD.n3038 9.3005
R26212 VDD.n3138 VDD.n3137 9.3005
R26213 VDD.n3139 VDD.n3037 9.3005
R26214 VDD.n3141 VDD.n3140 9.3005
R26215 VDD.n3142 VDD.n3035 9.3005
R26216 VDD.n3148 VDD.n3147 9.3005
R26217 VDD.n3149 VDD.n3034 9.3005
R26218 VDD.n3151 VDD.n3150 9.3005
R26219 VDD.n3152 VDD.n3032 9.3005
R26220 VDD.n3156 VDD.n3155 9.3005
R26221 VDD.n3157 VDD.n3031 9.3005
R26222 VDD.n3160 VDD.n3158 9.3005
R26223 VDD.n3161 VDD.n3030 9.3005
R26224 VDD.n3163 VDD.n3162 9.3005
R26225 VDD.n3164 VDD.n3029 9.3005
R26226 VDD.n3166 VDD.n3165 9.3005
R26227 VDD.n3167 VDD.n3028 9.3005
R26228 VDD.n3171 VDD.n3170 9.3005
R26229 VDD.n3173 VDD.n3172 9.3005
R26230 VDD.n3174 VDD.n3025 9.3005
R26231 VDD.n3176 VDD.n3175 9.3005
R26232 VDD.n3177 VDD.n3024 9.3005
R26233 VDD.n3179 VDD.n3178 9.3005
R26234 VDD.n3181 VDD.n3023 9.3005
R26235 VDD.n3183 VDD.n3182 9.3005
R26236 VDD.n3185 VDD.n3184 9.3005
R26237 VDD.n3187 VDD.n3020 9.3005
R26238 VDD.n3191 VDD.n3190 9.3005
R26239 VDD.n3192 VDD.n3019 9.3005
R26240 VDD.n3194 VDD.n3193 9.3005
R26241 VDD.n3197 VDD.n3018 9.3005
R26242 VDD.n3199 VDD.n3198 9.3005
R26243 VDD.n3200 VDD.n3017 9.3005
R26244 VDD.n3202 VDD.n3201 9.3005
R26245 VDD.n3203 VDD.n3016 9.3005
R26246 VDD.n3204 VDD.n3013 9.3005
R26247 VDD.n3206 VDD.n3205 9.3005
R26248 VDD.n3207 VDD.n3012 9.3005
R26249 VDD.n3209 VDD.n3208 9.3005
R26250 VDD.n3211 VDD.n3009 9.3005
R26251 VDD.n3213 VDD.n3212 9.3005
R26252 VDD.n3214 VDD.n3008 9.3005
R26253 VDD.n3216 VDD.n3215 9.3005
R26254 VDD.n3217 VDD.n3007 9.3005
R26255 VDD.n3218 VDD.n3006 9.3005
R26256 VDD.n3219 VDD.n3005 9.3005
R26257 VDD.n3221 VDD.n3220 9.3005
R26258 VDD.n3222 VDD.n3004 9.3005
R26259 VDD.n3224 VDD.n3223 9.3005
R26260 VDD.n3225 VDD.n3002 9.3005
R26261 VDD.n3226 VDD.n3001 9.3005
R26262 VDD.n3227 VDD.n2999 9.3005
R26263 VDD.n3228 VDD.n2998 9.3005
R26264 VDD.n3229 VDD.n2996 9.3005
R26265 VDD.n3231 VDD.n3230 9.3005
R26266 VDD.n3232 VDD.n2995 9.3005
R26267 VDD.n3294 VDD.n3293 9.3005
R26268 VDD.n3292 VDD.n2994 9.3005
R26269 VDD.n3291 VDD.n3290 9.3005
R26270 VDD.n3289 VDD.n3233 9.3005
R26271 VDD.n3288 VDD.n3287 9.3005
R26272 VDD.n3286 VDD.n3234 9.3005
R26273 VDD.n3285 VDD.n3284 9.3005
R26274 VDD.n3283 VDD.n3235 9.3005
R26275 VDD.n3281 VDD.n3280 9.3005
R26276 VDD.n3279 VDD.n3236 9.3005
R26277 VDD.n3278 VDD.n3277 9.3005
R26278 VDD.n3275 VDD.n3237 9.3005
R26279 VDD.n3274 VDD.n3273 9.3005
R26280 VDD.n3272 VDD.n3238 9.3005
R26281 VDD.n3271 VDD.n3270 9.3005
R26282 VDD.n3269 VDD.n3239 9.3005
R26283 VDD.n3268 VDD.n3267 9.3005
R26284 VDD.n3266 VDD.n3241 9.3005
R26285 VDD.n3265 VDD.n3264 9.3005
R26286 VDD.n3263 VDD.n3242 9.3005
R26287 VDD.n3262 VDD.n3260 9.3005
R26288 VDD.n3259 VDD.n3243 9.3005
R26289 VDD.n3258 VDD.n3257 9.3005
R26290 VDD.n3256 VDD.n3244 9.3005
R26291 VDD.n3253 VDD.n3252 9.3005
R26292 VDD.n3251 VDD.n3245 9.3005
R26293 VDD.n3250 VDD.n3249 9.3005
R26294 VDD.n2993 VDD.n2992 9.3005
R26295 VDD.n3298 VDD.n3297 9.3005
R26296 VDD.n3300 VDD.n3299 9.3005
R26297 VDD.n3301 VDD.n2988 9.3005
R26298 VDD.n3303 VDD.n3302 9.3005
R26299 VDD.n3304 VDD.n2987 9.3005
R26300 VDD.n3306 VDD.n3305 9.3005
R26301 VDD.n3307 VDD.n2985 9.3005
R26302 VDD.n3309 VDD.n3308 9.3005
R26303 VDD.n3311 VDD.n3310 9.3005
R26304 VDD.n3313 VDD.n2982 9.3005
R26305 VDD.n3316 VDD.n3315 9.3005
R26306 VDD.n3318 VDD.n3317 9.3005
R26307 VDD.n3319 VDD.n2979 9.3005
R26308 VDD.n3320 VDD.n2978 9.3005
R26309 VDD.n3321 VDD.n2977 9.3005
R26310 VDD.n3325 VDD.n3324 9.3005
R26311 VDD.n3326 VDD.n2976 9.3005
R26312 VDD.n3328 VDD.n3327 9.3005
R26313 VDD.n3329 VDD.n2974 9.3005
R26314 VDD.n3332 VDD.n3331 9.3005
R26315 VDD.n3333 VDD.n2973 9.3005
R26316 VDD.n3335 VDD.n3334 9.3005
R26317 VDD.n3336 VDD.n2972 9.3005
R26318 VDD.n3340 VDD.n3339 9.3005
R26319 VDD.n3342 VDD.n3341 9.3005
R26320 VDD.n3343 VDD.n2968 9.3005
R26321 VDD.n3345 VDD.n3344 9.3005
R26322 VDD.n3346 VDD.n2967 9.3005
R26323 VDD.n3420 VDD.n3419 9.3005
R26324 VDD.n3418 VDD.n2966 9.3005
R26325 VDD.n3417 VDD.n3416 9.3005
R26326 VDD.n3415 VDD.n3347 9.3005
R26327 VDD.n3413 VDD.n3412 9.3005
R26328 VDD.n3411 VDD.n3350 9.3005
R26329 VDD.n3410 VDD.n3409 9.3005
R26330 VDD.n3408 VDD.n3351 9.3005
R26331 VDD.n3406 VDD.n3405 9.3005
R26332 VDD.n3404 VDD.n3354 9.3005
R26333 VDD.n3403 VDD.n3402 9.3005
R26334 VDD.n3400 VDD.n3355 9.3005
R26335 VDD.n3399 VDD.n3398 9.3005
R26336 VDD.n3397 VDD.n3356 9.3005
R26337 VDD.n3396 VDD.n3395 9.3005
R26338 VDD.n3393 VDD.n3358 9.3005
R26339 VDD.n3392 VDD.n3391 9.3005
R26340 VDD.n3390 VDD.n3359 9.3005
R26341 VDD.n3389 VDD.n3388 9.3005
R26342 VDD.n3385 VDD.n3360 9.3005
R26343 VDD.n3384 VDD.n3383 9.3005
R26344 VDD.n3382 VDD.n3363 9.3005
R26345 VDD.n3381 VDD.n3380 9.3005
R26346 VDD.n3379 VDD.n3364 9.3005
R26347 VDD.n3376 VDD.n3375 9.3005
R26348 VDD.n3374 VDD.n3366 9.3005
R26349 VDD.n3373 VDD.n3372 9.3005
R26350 VDD.n3367 VDD.n2965 9.3005
R26351 VDD.n3424 VDD.n2964 9.3005
R26352 VDD.n3427 VDD.n3426 9.3005
R26353 VDD.n3429 VDD.n3428 9.3005
R26354 VDD.n3430 VDD.n2962 9.3005
R26355 VDD.n3431 VDD.n2961 9.3005
R26356 VDD.n3435 VDD.n3434 9.3005
R26357 VDD.n3436 VDD.n2960 9.3005
R26358 VDD.n3438 VDD.n3437 9.3005
R26359 VDD.n3440 VDD.n2958 9.3005
R26360 VDD.n3443 VDD.n3442 9.3005
R26361 VDD.n3444 VDD.n2957 9.3005
R26362 VDD.n3446 VDD.n3445 9.3005
R26363 VDD.n3447 VDD.n2955 9.3005
R26364 VDD.n3448 VDD.n2954 9.3005
R26365 VDD.n3450 VDD.n2952 9.3005
R26366 VDD.n3452 VDD.n3451 9.3005
R26367 VDD.n3453 VDD.n2951 9.3005
R26368 VDD.n3455 VDD.n3454 9.3005
R26369 VDD.n3456 VDD.n2950 9.3005
R26370 VDD.n3457 VDD.n2948 9.3005
R26371 VDD.n3462 VDD.n3461 9.3005
R26372 VDD.n3463 VDD.n2947 9.3005
R26373 VDD.n3465 VDD.n3464 9.3005
R26374 VDD.n3467 VDD.n2945 9.3005
R26375 VDD.n3469 VDD.n3468 9.3005
R26376 VDD.n3471 VDD.n3470 9.3005
R26377 VDD.n3473 VDD.n2941 9.3005
R26378 VDD.n3476 VDD.n3475 9.3005
R26379 VDD.n3477 VDD.n2940 9.3005
R26380 VDD.n3479 VDD.n3478 9.3005
R26381 VDD.n3480 VDD.n2938 9.3005
R26382 VDD.n3481 VDD.n2937 9.3005
R26383 VDD.n3483 VDD.n3482 9.3005
R26384 VDD.n3485 VDD.n3484 9.3005
R26385 VDD.n3487 VDD.n2934 9.3005
R26386 VDD.n3489 VDD.n3488 9.3005
R26387 VDD.n3490 VDD.n2933 9.3005
R26388 VDD.n3492 VDD.n3491 9.3005
R26389 VDD.n3493 VDD.n2931 9.3005
R26390 VDD.n3494 VDD.n2930 9.3005
R26391 VDD.n3496 VDD.n3495 9.3005
R26392 VDD.n3497 VDD.n2929 9.3005
R26393 VDD.n3499 VDD.n3498 9.3005
R26394 VDD.n3501 VDD.n2921 9.3005
R26395 VDD.n3505 VDD.n3504 9.3005
R26396 VDD.n3507 VDD.n3506 9.3005
R26397 VDD.n3508 VDD.n2918 9.3005
R26398 VDD.n3510 VDD.n3509 9.3005
R26399 VDD.n3511 VDD.n2917 9.3005
R26400 VDD.n3513 VDD.n3512 9.3005
R26401 VDD.n3514 VDD.n2914 9.3005
R26402 VDD.n3518 VDD.n3517 9.3005
R26403 VDD.n3519 VDD.n2912 9.3005
R26404 VDD.n3572 VDD.n3571 9.3005
R26405 VDD.n3570 VDD.n2913 9.3005
R26406 VDD.n3569 VDD.n3568 9.3005
R26407 VDD.n3565 VDD.n3520 9.3005
R26408 VDD.n3564 VDD.n3563 9.3005
R26409 VDD.n3562 VDD.n3523 9.3005
R26410 VDD.n3561 VDD.n3560 9.3005
R26411 VDD.n3559 VDD.n3524 9.3005
R26412 VDD.n3558 VDD.n3526 9.3005
R26413 VDD.n3557 VDD.n3556 9.3005
R26414 VDD.n3555 VDD.n3554 9.3005
R26415 VDD.n3552 VDD.n3528 9.3005
R26416 VDD.n3550 VDD.n3549 9.3005
R26417 VDD.n3548 VDD.n3547 9.3005
R26418 VDD.n3546 VDD.n3531 9.3005
R26419 VDD.n3545 VDD.n3533 9.3005
R26420 VDD.n3544 VDD.n3543 9.3005
R26421 VDD.n3542 VDD.n3534 9.3005
R26422 VDD.n3541 VDD.n3540 9.3005
R26423 VDD.n3539 VDD.n3535 9.3005
R26424 VDD.n3538 VDD.n2896 9.3005
R26425 VDD.n3653 VDD.n3652 9.3005
R26426 VDD.n3651 VDD.n2900 9.3005
R26427 VDD.n3650 VDD.n3649 9.3005
R26428 VDD.n3648 VDD.n2901 9.3005
R26429 VDD.n3647 VDD.n3646 9.3005
R26430 VDD.n3643 VDD.n2909 9.3005
R26431 VDD.n3642 VDD.n3641 9.3005
R26432 VDD.n3640 VDD.n3575 9.3005
R26433 VDD.n3639 VDD.n3638 9.3005
R26434 VDD.n3636 VDD.n3635 9.3005
R26435 VDD.n3634 VDD.n3633 9.3005
R26436 VDD.n3632 VDD.n3584 9.3005
R26437 VDD.n3631 VDD.n3630 9.3005
R26438 VDD.n3629 VDD.n3628 9.3005
R26439 VDD.n3627 VDD.n3586 9.3005
R26440 VDD.n3626 VDD.n3625 9.3005
R26441 VDD.n3624 VDD.n3587 9.3005
R26442 VDD.n3623 VDD.n3622 9.3005
R26443 VDD.n3621 VDD.n3588 9.3005
R26444 VDD.n3620 VDD.n3619 9.3005
R26445 VDD.n3618 VDD.n3617 9.3005
R26446 VDD.n3616 VDD.n3590 9.3005
R26447 VDD.n3615 VDD.n3592 9.3005
R26448 VDD.n3614 VDD.n3613 9.3005
R26449 VDD.n3612 VDD.n3594 9.3005
R26450 VDD.n3611 VDD.n3610 9.3005
R26451 VDD.n3609 VDD.n3595 9.3005
R26452 VDD.n3608 VDD.n3607 9.3005
R26453 VDD.n2483 VDD.n2482 9.3005
R26454 VDD.n2484 VDD.n2471 9.3005
R26455 VDD.n2485 VDD.n2469 9.3005
R26456 VDD.n2488 VDD.n2487 9.3005
R26457 VDD.n2490 VDD.n2489 9.3005
R26458 VDD.n2491 VDD.n2466 9.3005
R26459 VDD.n2492 VDD.n2465 9.3005
R26460 VDD.n2464 VDD.n2399 9.3005
R26461 VDD.n2463 VDD.n2462 9.3005
R26462 VDD.n2461 VDD.n2400 9.3005
R26463 VDD.n2460 VDD.n2402 9.3005
R26464 VDD.n2459 VDD.n2403 9.3005
R26465 VDD.n2458 VDD.n2404 9.3005
R26466 VDD.n2457 VDD.n2405 9.3005
R26467 VDD.n2455 VDD.n2454 9.3005
R26468 VDD.n2453 VDD.n2452 9.3005
R26469 VDD.n2450 VDD.n2408 9.3005
R26470 VDD.n2449 VDD.n2448 9.3005
R26471 VDD.n2447 VDD.n2446 9.3005
R26472 VDD.n2445 VDD.n2410 9.3005
R26473 VDD.n2444 VDD.n2443 9.3005
R26474 VDD.n2442 VDD.n2441 9.3005
R26475 VDD.n2440 VDD.n2412 9.3005
R26476 VDD.n2438 VDD.n2437 9.3005
R26477 VDD.n2436 VDD.n2413 9.3005
R26478 VDD.n2435 VDD.n2434 9.3005
R26479 VDD.n2432 VDD.n2414 9.3005
R26480 VDD.n2430 VDD.n2429 9.3005
R26481 VDD.n2428 VDD.n2416 9.3005
R26482 VDD.n2427 VDD.n2426 9.3005
R26483 VDD.n2424 VDD.n2417 9.3005
R26484 VDD.n2423 VDD.n2422 9.3005
R26485 VDD.n2421 VDD.n2419 9.3005
R26486 VDD.n2420 VDD.n2398 9.3005
R26487 VDD.n2495 VDD.n2397 9.3005
R26488 VDD.n2497 VDD.n2496 9.3005
R26489 VDD.n2501 VDD.n2395 9.3005
R26490 VDD.n2505 VDD.n2504 9.3005
R26491 VDD.n2507 VDD.n2506 9.3005
R26492 VDD.n2508 VDD.n2392 9.3005
R26493 VDD.n2511 VDD.n2510 9.3005
R26494 VDD.n2513 VDD.n2512 9.3005
R26495 VDD.n2515 VDD.n2390 9.3005
R26496 VDD.n2517 VDD.n2516 9.3005
R26497 VDD.n2519 VDD.n2518 9.3005
R26498 VDD.n2521 VDD.n2388 9.3005
R26499 VDD.n2524 VDD.n2523 9.3005
R26500 VDD.n2525 VDD.n2387 9.3005
R26501 VDD.n2527 VDD.n2526 9.3005
R26502 VDD.n2528 VDD.n2384 9.3005
R26503 VDD.n2535 VDD.n2534 9.3005
R26504 VDD.n2536 VDD.n2383 9.3005
R26505 VDD.n2538 VDD.n2537 9.3005
R26506 VDD.n2539 VDD.n2381 9.3005
R26507 VDD.n2542 VDD.n2541 9.3005
R26508 VDD.n2543 VDD.n2380 9.3005
R26509 VDD.n2545 VDD.n2544 9.3005
R26510 VDD.n2549 VDD.n2379 9.3005
R26511 VDD.n2551 VDD.n2550 9.3005
R26512 VDD.n2553 VDD.n2552 9.3005
R26513 VDD.n2555 VDD.n2377 9.3005
R26514 VDD.n2560 VDD.n2559 9.3005
R26515 VDD.n2561 VDD.n2367 9.3005
R26516 VDD.n2563 VDD.n2562 9.3005
R26517 VDD.n2566 VDD.n2364 9.3005
R26518 VDD.n2568 VDD.n2567 9.3005
R26519 VDD.n2569 VDD.n2363 9.3005
R26520 VDD.n2571 VDD.n2570 9.3005
R26521 VDD.n2572 VDD.n2360 9.3005
R26522 VDD.n2579 VDD.n2578 9.3005
R26523 VDD.n2580 VDD.n2359 9.3005
R26524 VDD.n2582 VDD.n2581 9.3005
R26525 VDD.n2584 VDD.n2353 9.3005
R26526 VDD.n2585 VDD.n2352 9.3005
R26527 VDD.n2586 VDD.n2350 9.3005
R26528 VDD.n2588 VDD.n2587 9.3005
R26529 VDD.n2589 VDD.n2349 9.3005
R26530 VDD.n2591 VDD.n2590 9.3005
R26531 VDD.n2593 VDD.n2344 9.3005
R26532 VDD.n2594 VDD.n2343 9.3005
R26533 VDD.n2595 VDD.n2342 9.3005
R26534 VDD.n2341 VDD.n2340 9.3005
R26535 VDD.n2338 VDD.n2336 9.3005
R26536 VDD.n2600 VDD.n2335 9.3005
R26537 VDD.n2602 VDD.n2601 9.3005
R26538 VDD.n2604 VDD.n2603 9.3005
R26539 VDD.n2605 VDD.n2333 9.3005
R26540 VDD.n2608 VDD.n2607 9.3005
R26541 VDD.n2609 VDD.n2332 9.3005
R26542 VDD.n2611 VDD.n2610 9.3005
R26543 VDD.n2613 VDD.n2330 9.3005
R26544 VDD.n2617 VDD.n2616 9.3005
R26545 VDD.n2619 VDD.n2618 9.3005
R26546 VDD.n2620 VDD.n2328 9.3005
R26547 VDD.n2623 VDD.n2622 9.3005
R26548 VDD.n2625 VDD.n2624 9.3005
R26549 VDD.n2626 VDD.n2325 9.3005
R26550 VDD.n2627 VDD.n2323 9.3005
R26551 VDD.n2628 VDD.n2322 9.3005
R26552 VDD.n2629 VDD.n2320 9.3005
R26553 VDD.n2631 VDD.n2630 9.3005
R26554 VDD.n2633 VDD.n2632 9.3005
R26555 VDD.n2634 VDD.n2317 9.3005
R26556 VDD.n2637 VDD.n2636 9.3005
R26557 VDD.n2639 VDD.n2638 9.3005
R26558 VDD.n2640 VDD.n2313 9.3005
R26559 VDD.n2641 VDD.n2312 9.3005
R26560 VDD.n2642 VDD.n2310 9.3005
R26561 VDD.n2309 VDD.n2308 9.3005
R26562 VDD.n2649 VDD.n2305 9.3005
R26563 VDD.n2652 VDD.n2651 9.3005
R26564 VDD.n2653 VDD.n2304 9.3005
R26565 VDD.n2655 VDD.n2654 9.3005
R26566 VDD.n2657 VDD.n2303 9.3005
R26567 VDD.n2662 VDD.n2661 9.3005
R26568 VDD.n2663 VDD.n2302 9.3005
R26569 VDD.n2665 VDD.n2664 9.3005
R26570 VDD.n2666 VDD.n2301 9.3005
R26571 VDD.n2669 VDD.n2668 9.3005
R26572 VDD.n2671 VDD.n2670 9.3005
R26573 VDD.n2672 VDD.n2298 9.3005
R26574 VDD.n2674 VDD.n2673 9.3005
R26575 VDD.n2675 VDD.n2297 9.3005
R26576 VDD.n2677 VDD.n2676 9.3005
R26577 VDD.n2678 VDD.n2295 9.3005
R26578 VDD.n2682 VDD.n2681 9.3005
R26579 VDD.n2683 VDD.n2294 9.3005
R26580 VDD.n2685 VDD.n2684 9.3005
R26581 VDD.n2687 VDD.n2292 9.3005
R26582 VDD.n2689 VDD.n2688 9.3005
R26583 VDD.n2691 VDD.n2690 9.3005
R26584 VDD.n2692 VDD.n2289 9.3005
R26585 VDD.n2695 VDD.n2694 9.3005
R26586 VDD.n2697 VDD.n2696 9.3005
R26587 VDD.n2698 VDD.n2286 9.3005
R26588 VDD.n2703 VDD.n2702 9.3005
R26589 VDD.n2704 VDD.n2285 9.3005
R26590 VDD.n2706 VDD.n2705 9.3005
R26591 VDD.n2709 VDD.n2283 9.3005
R26592 VDD.n2711 VDD.n2710 9.3005
R26593 VDD.n2713 VDD.n2712 9.3005
R26594 VDD.n2714 VDD.n2280 9.3005
R26595 VDD.n2717 VDD.n2716 9.3005
R26596 VDD.n2719 VDD.n2718 9.3005
R26597 VDD.n2720 VDD.n2276 9.3005
R26598 VDD.n2721 VDD.n2275 9.3005
R26599 VDD.n2725 VDD.n2724 9.3005
R26600 VDD.n2726 VDD.n2274 9.3005
R26601 VDD.n2728 VDD.n2727 9.3005
R26602 VDD.n2730 VDD.n2273 9.3005
R26603 VDD.n2734 VDD.n2733 9.3005
R26604 VDD.n2735 VDD.n2272 9.3005
R26605 VDD.n2737 VDD.n2736 9.3005
R26606 VDD.n2738 VDD.n2269 9.3005
R26607 VDD.n2742 VDD.n2741 9.3005
R26608 VDD.n2743 VDD.n2268 9.3005
R26609 VDD.n2745 VDD.n2744 9.3005
R26610 VDD.n2746 VDD.n2267 9.3005
R26611 VDD.n2749 VDD.n2748 9.3005
R26612 VDD.n2750 VDD.n2266 9.3005
R26613 VDD.n2752 VDD.n2751 9.3005
R26614 VDD.n2755 VDD.n2262 9.3005
R26615 VDD.n2757 VDD.n2756 9.3005
R26616 VDD.n2758 VDD.n2261 9.3005
R26617 VDD.n2760 VDD.n2759 9.3005
R26618 VDD.n2763 VDD.n2259 9.3005
R26619 VDD.n2767 VDD.n2766 9.3005
R26620 VDD.n2769 VDD.n2768 9.3005
R26621 VDD.n2770 VDD.n2257 9.3005
R26622 VDD.n2772 VDD.n2771 9.3005
R26623 VDD.n2774 VDD.n2773 9.3005
R26624 VDD.n2775 VDD.n2254 9.3005
R26625 VDD.n2776 VDD.n2253 9.3005
R26626 VDD.n2778 VDD.n2777 9.3005
R26627 VDD.n2779 VDD.n2252 9.3005
R26628 VDD.n2781 VDD.n2780 9.3005
R26629 VDD.n2783 VDD.n2249 9.3005
R26630 VDD.n2787 VDD.n2786 9.3005
R26631 VDD.n2789 VDD.n2788 9.3005
R26632 VDD.n2791 VDD.n2247 9.3005
R26633 VDD.n2794 VDD.n2793 9.3005
R26634 VDD.n2795 VDD.n2246 9.3005
R26635 VDD.n2797 VDD.n2796 9.3005
R26636 VDD.n2800 VDD.n2243 9.3005
R26637 VDD.n2802 VDD.n2801 9.3005
R26638 VDD.n2804 VDD.n2803 9.3005
R26639 VDD.n2805 VDD.n2239 9.3005
R26640 VDD.n2808 VDD.n2807 9.3005
R26641 VDD.n2809 VDD.n2238 9.3005
R26642 VDD.n2811 VDD.n2810 9.3005
R26643 VDD.n2812 VDD.n2236 9.3005
R26644 VDD.n2818 VDD.n2817 9.3005
R26645 VDD.n2819 VDD.n2235 9.3005
R26646 VDD.n2821 VDD.n2820 9.3005
R26647 VDD.n2823 VDD.n2234 9.3005
R26648 VDD.n2826 VDD.n2825 9.3005
R26649 VDD.n2828 VDD.n2827 9.3005
R26650 VDD.n2829 VDD.n2232 9.3005
R26651 VDD.n2833 VDD.n2832 9.3005
R26652 VDD.n2836 VDD.n2835 9.3005
R26653 VDD.n2843 VDD.n2842 9.3005
R26654 VDD.n2844 VDD.n2224 9.3005
R26655 VDD.n2846 VDD.n2845 9.3005
R26656 VDD.n2849 VDD.n2222 9.3005
R26657 VDD.n2852 VDD.n2851 9.3005
R26658 VDD.n2853 VDD.n2221 9.3005
R26659 VDD.n2855 VDD.n2854 9.3005
R26660 VDD.n2856 VDD.n2219 9.3005
R26661 VDD.n2861 VDD.n2860 9.3005
R26662 VDD.n2862 VDD.n2218 9.3005
R26663 VDD.n2864 VDD.n2863 9.3005
R26664 VDD.n2865 VDD.n2217 9.3005
R26665 VDD.n2216 VDD.n2165 9.3005
R26666 VDD.n2215 VDD.n2214 9.3005
R26667 VDD.n2213 VDD.n2166 9.3005
R26668 VDD.n2211 VDD.n2210 9.3005
R26669 VDD.n2209 VDD.n2167 9.3005
R26670 VDD.n2208 VDD.n2207 9.3005
R26671 VDD.n2204 VDD.n2168 9.3005
R26672 VDD.n2203 VDD.n2202 9.3005
R26673 VDD.n2201 VDD.n2169 9.3005
R26674 VDD.n2200 VDD.n2199 9.3005
R26675 VDD.n2198 VDD.n2170 9.3005
R26676 VDD.n2196 VDD.n2195 9.3005
R26677 VDD.n2194 VDD.n2174 9.3005
R26678 VDD.n2193 VDD.n2192 9.3005
R26679 VDD.n2191 VDD.n2175 9.3005
R26680 VDD.n2189 VDD.n2188 9.3005
R26681 VDD.n2187 VDD.n2186 9.3005
R26682 VDD.n2185 VDD.n2178 9.3005
R26683 VDD.n2183 VDD.n2182 9.3005
R26684 VDD.n2180 VDD.n2091 9.3005
R26685 VDD.n2887 VDD.n2886 9.3005
R26686 VDD.n2885 VDD.n2884 9.3005
R26687 VDD.n2877 VDD.n2094 9.3005
R26688 VDD.n2876 VDD.n2875 9.3005
R26689 VDD.n2874 VDD.n2096 9.3005
R26690 VDD.n2872 VDD.n2871 9.3005
R26691 VDD.n2870 VDD.n2869 9.3005
R26692 VDD.n2868 VDD.n2100 9.3005
R26693 VDD.n2161 VDD.n2160 9.3005
R26694 VDD.n2158 VDD.n2111 9.3005
R26695 VDD.n2155 VDD.n2154 9.3005
R26696 VDD.n2153 VDD.n2115 9.3005
R26697 VDD.n2152 VDD.n2151 9.3005
R26698 VDD.n2150 VDD.n2116 9.3005
R26699 VDD.n2149 VDD.n2117 9.3005
R26700 VDD.n2148 VDD.n2147 9.3005
R26701 VDD.n2146 VDD.n2118 9.3005
R26702 VDD.n2145 VDD.n2144 9.3005
R26703 VDD.n2143 VDD.n2119 9.3005
R26704 VDD.n2142 VDD.n2141 9.3005
R26705 VDD.n2140 VDD.n2122 9.3005
R26706 VDD.n2139 VDD.n2138 9.3005
R26707 VDD.n2137 VDD.n2123 9.3005
R26708 VDD.n2136 VDD.n2135 9.3005
R26709 VDD.n1665 VDD.n1664 9.3005
R26710 VDD.n1666 VDD.n1653 9.3005
R26711 VDD.n1667 VDD.n1651 9.3005
R26712 VDD.n1670 VDD.n1669 9.3005
R26713 VDD.n1672 VDD.n1671 9.3005
R26714 VDD.n1673 VDD.n1648 9.3005
R26715 VDD.n1674 VDD.n1647 9.3005
R26716 VDD.n1646 VDD.n1645 9.3005
R26717 VDD.n1643 VDD.n1578 9.3005
R26718 VDD.n1642 VDD.n1641 9.3005
R26719 VDD.n1640 VDD.n1579 9.3005
R26720 VDD.n1639 VDD.n1638 9.3005
R26721 VDD.n1637 VDD.n1581 9.3005
R26722 VDD.n1635 VDD.n1634 9.3005
R26723 VDD.n1633 VDD.n1632 9.3005
R26724 VDD.n1631 VDD.n1583 9.3005
R26725 VDD.n1630 VDD.n1629 9.3005
R26726 VDD.n1628 VDD.n1627 9.3005
R26727 VDD.n1625 VDD.n1585 9.3005
R26728 VDD.n1623 VDD.n1622 9.3005
R26729 VDD.n1621 VDD.n1620 9.3005
R26730 VDD.n1619 VDD.n1587 9.3005
R26731 VDD.n1618 VDD.n1617 9.3005
R26732 VDD.n1616 VDD.n1588 9.3005
R26733 VDD.n1615 VDD.n1614 9.3005
R26734 VDD.n1613 VDD.n1589 9.3005
R26735 VDD.n1611 VDD.n1610 9.3005
R26736 VDD.n1609 VDD.n1608 9.3005
R26737 VDD.n1607 VDD.n1592 9.3005
R26738 VDD.n1604 VDD.n1603 9.3005
R26739 VDD.n1602 VDD.n1593 9.3005
R26740 VDD.n1601 VDD.n1600 9.3005
R26741 VDD.n1598 VDD.n1594 9.3005
R26742 VDD.n1576 VDD.n1575 9.3005
R26743 VDD.n1678 VDD.n1677 9.3005
R26744 VDD.n1685 VDD.n1573 9.3005
R26745 VDD.n1688 VDD.n1687 9.3005
R26746 VDD.n1690 VDD.n1689 9.3005
R26747 VDD.n1692 VDD.n1569 9.3005
R26748 VDD.n1695 VDD.n1694 9.3005
R26749 VDD.n1697 VDD.n1696 9.3005
R26750 VDD.n1700 VDD.n1567 9.3005
R26751 VDD.n1704 VDD.n1703 9.3005
R26752 VDD.n1705 VDD.n1566 9.3005
R26753 VDD.n1707 VDD.n1706 9.3005
R26754 VDD.n1708 VDD.n1564 9.3005
R26755 VDD.n1710 VDD.n1709 9.3005
R26756 VDD.n1711 VDD.n1563 9.3005
R26757 VDD.n1713 VDD.n1712 9.3005
R26758 VDD.n1716 VDD.n1562 9.3005
R26759 VDD.n1720 VDD.n1719 9.3005
R26760 VDD.n1721 VDD.n1561 9.3005
R26761 VDD.n1723 VDD.n1722 9.3005
R26762 VDD.n1724 VDD.n1560 9.3005
R26763 VDD.n1726 VDD.n1725 9.3005
R26764 VDD.n1727 VDD.n1558 9.3005
R26765 VDD.n1729 VDD.n1728 9.3005
R26766 VDD.n1731 VDD.n1557 9.3005
R26767 VDD.n1733 VDD.n1732 9.3005
R26768 VDD.n1734 VDD.n1554 9.3005
R26769 VDD.n1736 VDD.n1735 9.3005
R26770 VDD.n1737 VDD.n1553 9.3005
R26771 VDD.n1740 VDD.n1739 9.3005
R26772 VDD.n1741 VDD.n1552 9.3005
R26773 VDD.n1743 VDD.n1742 9.3005
R26774 VDD.n1753 VDD.n1752 9.3005
R26775 VDD.n1754 VDD.n1548 9.3005
R26776 VDD.n1756 VDD.n1755 9.3005
R26777 VDD.n1758 VDD.n1547 9.3005
R26778 VDD.n1762 VDD.n1761 9.3005
R26779 VDD.n1764 VDD.n1763 9.3005
R26780 VDD.n1765 VDD.n1544 9.3005
R26781 VDD.n1767 VDD.n1766 9.3005
R26782 VDD.n1768 VDD.n1543 9.3005
R26783 VDD.n1770 VDD.n1769 9.3005
R26784 VDD.n1771 VDD.n1541 9.3005
R26785 VDD.n1774 VDD.n1773 9.3005
R26786 VDD.n1775 VDD.n1539 9.3005
R26787 VDD.n1777 VDD.n1776 9.3005
R26788 VDD.n1778 VDD.n1538 9.3005
R26789 VDD.n1782 VDD.n1781 9.3005
R26790 VDD.n1783 VDD.n1537 9.3005
R26791 VDD.n1785 VDD.n1784 9.3005
R26792 VDD.n1787 VDD.n1536 9.3005
R26793 VDD.n1791 VDD.n1790 9.3005
R26794 VDD.n1792 VDD.n1535 9.3005
R26795 VDD.n1794 VDD.n1793 9.3005
R26796 VDD.n1796 VDD.n1532 9.3005
R26797 VDD.n1798 VDD.n1797 9.3005
R26798 VDD.n1799 VDD.n1531 9.3005
R26799 VDD.n1801 VDD.n1800 9.3005
R26800 VDD.n1802 VDD.n1530 9.3005
R26801 VDD.n1806 VDD.n1805 9.3005
R26802 VDD.n1807 VDD.n1529 9.3005
R26803 VDD.n1809 VDD.n1808 9.3005
R26804 VDD.n1810 VDD.n1527 9.3005
R26805 VDD.n1811 VDD.n1525 9.3005
R26806 VDD.n1813 VDD.n1812 9.3005
R26807 VDD.n1814 VDD.n1524 9.3005
R26808 VDD.n1816 VDD.n1815 9.3005
R26809 VDD.n1817 VDD.n1521 9.3005
R26810 VDD.n1821 VDD.n1820 9.3005
R26811 VDD.n1823 VDD.n1822 9.3005
R26812 VDD.n1824 VDD.n1519 9.3005
R26813 VDD.n1826 VDD.n1516 9.3005
R26814 VDD.n1829 VDD.n1828 9.3005
R26815 VDD.n1831 VDD.n1830 9.3005
R26816 VDD.n1834 VDD.n1512 9.3005
R26817 VDD.n1836 VDD.n1835 9.3005
R26818 VDD.n1837 VDD.n1511 9.3005
R26819 VDD.n1839 VDD.n1838 9.3005
R26820 VDD.n1840 VDD.n1510 9.3005
R26821 VDD.n1842 VDD.n1841 9.3005
R26822 VDD.n1844 VDD.n1843 9.3005
R26823 VDD.n1845 VDD.n1507 9.3005
R26824 VDD.n1851 VDD.n1850 9.3005
R26825 VDD.n1852 VDD.n1506 9.3005
R26826 VDD.n1854 VDD.n1853 9.3005
R26827 VDD.n1856 VDD.n1505 9.3005
R26828 VDD.n1858 VDD.n1857 9.3005
R26829 VDD.n1859 VDD.n1504 9.3005
R26830 VDD.n1861 VDD.n1860 9.3005
R26831 VDD.n1862 VDD.n1501 9.3005
R26832 VDD.n1864 VDD.n1863 9.3005
R26833 VDD.n1865 VDD.n1500 9.3005
R26834 VDD.n1867 VDD.n1866 9.3005
R26835 VDD.n1868 VDD.n1498 9.3005
R26836 VDD.n1870 VDD.n1869 9.3005
R26837 VDD.n1871 VDD.n1497 9.3005
R26838 VDD.n1873 VDD.n1872 9.3005
R26839 VDD.n1875 VDD.n1495 9.3005
R26840 VDD.n1876 VDD.n1493 9.3005
R26841 VDD.n1877 VDD.n1492 9.3005
R26842 VDD.n1878 VDD.n1490 9.3005
R26843 VDD.n1880 VDD.n1879 9.3005
R26844 VDD.n1881 VDD.n1489 9.3005
R26845 VDD.n1883 VDD.n1882 9.3005
R26846 VDD.n1885 VDD.n1485 9.3005
R26847 VDD.n1887 VDD.n1886 9.3005
R26848 VDD.n1888 VDD.n1484 9.3005
R26849 VDD.n1890 VDD.n1889 9.3005
R26850 VDD.n1891 VDD.n1478 9.3005
R26851 VDD.n1896 VDD.n1895 9.3005
R26852 VDD.n1897 VDD.n1477 9.3005
R26853 VDD.n1899 VDD.n1898 9.3005
R26854 VDD.n1901 VDD.n1475 9.3005
R26855 VDD.n1904 VDD.n1903 9.3005
R26856 VDD.n1905 VDD.n1474 9.3005
R26857 VDD.n1907 VDD.n1906 9.3005
R26858 VDD.n1909 VDD.n1472 9.3005
R26859 VDD.n1910 VDD.n1470 9.3005
R26860 VDD.n1914 VDD.n1913 9.3005
R26861 VDD.n1916 VDD.n1915 9.3005
R26862 VDD.n1918 VDD.n1467 9.3005
R26863 VDD.n1920 VDD.n1919 9.3005
R26864 VDD.n1922 VDD.n1921 9.3005
R26865 VDD.n1924 VDD.n1465 9.3005
R26866 VDD.n1926 VDD.n1925 9.3005
R26867 VDD.n1928 VDD.n1927 9.3005
R26868 VDD.n1929 VDD.n1462 9.3005
R26869 VDD.n1933 VDD.n1932 9.3005
R26870 VDD.n1934 VDD.n1461 9.3005
R26871 VDD.n1936 VDD.n1935 9.3005
R26872 VDD.n1937 VDD.n1459 9.3005
R26873 VDD.n1939 VDD.n1938 9.3005
R26874 VDD.n1940 VDD.n1458 9.3005
R26875 VDD.n1942 VDD.n1941 9.3005
R26876 VDD.n1943 VDD.n1456 9.3005
R26877 VDD.n1945 VDD.n1944 9.3005
R26878 VDD.n1948 VDD.n1947 9.3005
R26879 VDD.n1950 VDD.n1450 9.3005
R26880 VDD.n1952 VDD.n1951 9.3005
R26881 VDD.n1954 VDD.n1953 9.3005
R26882 VDD.n1956 VDD.n1447 9.3005
R26883 VDD.n1959 VDD.n1958 9.3005
R26884 VDD.n1961 VDD.n1960 9.3005
R26885 VDD.n1964 VDD.n1444 9.3005
R26886 VDD.n1967 VDD.n1966 9.3005
R26887 VDD.n1969 VDD.n1968 9.3005
R26888 VDD.n1970 VDD.n1442 9.3005
R26889 VDD.n1972 VDD.n1971 9.3005
R26890 VDD.n1973 VDD.n1441 9.3005
R26891 VDD.n1975 VDD.n1974 9.3005
R26892 VDD.n1978 VDD.n1437 9.3005
R26893 VDD.n1980 VDD.n1979 9.3005
R26894 VDD.n1981 VDD.n1436 9.3005
R26895 VDD.n1983 VDD.n1982 9.3005
R26896 VDD.n1984 VDD.n1435 9.3005
R26897 VDD.n1985 VDD.n1433 9.3005
R26898 VDD.n1987 VDD.n1986 9.3005
R26899 VDD.n1988 VDD.n1432 9.3005
R26900 VDD.n1990 VDD.n1989 9.3005
R26901 VDD.n1991 VDD.n1430 9.3005
R26902 VDD.n1993 VDD.n1992 9.3005
R26903 VDD.n1994 VDD.n1429 9.3005
R26904 VDD.n1996 VDD.n1995 9.3005
R26905 VDD.n1999 VDD.n1427 9.3005
R26906 VDD.n2003 VDD.n2002 9.3005
R26907 VDD.n2005 VDD.n2004 9.3005
R26908 VDD.n2007 VDD.n1424 9.3005
R26909 VDD.n2011 VDD.n2010 9.3005
R26910 VDD.n2013 VDD.n2012 9.3005
R26911 VDD.n2015 VDD.n1421 9.3005
R26912 VDD.n2018 VDD.n2017 9.3005
R26913 VDD.n2019 VDD.n1420 9.3005
R26914 VDD.n2021 VDD.n2020 9.3005
R26915 VDD.n2022 VDD.n1418 9.3005
R26916 VDD.n2026 VDD.n2025 9.3005
R26917 VDD.n2028 VDD.n2027 9.3005
R26918 VDD.n2030 VDD.n1414 9.3005
R26919 VDD.n2033 VDD.n2032 9.3005
R26920 VDD.n2035 VDD.n2034 9.3005
R26921 VDD.n2037 VDD.n1412 9.3005
R26922 VDD.n2039 VDD.n2038 9.3005
R26923 VDD.n2040 VDD.n1411 9.3005
R26924 VDD.n2042 VDD.n2041 9.3005
R26925 VDD.n2043 VDD.n1407 9.3005
R26926 VDD.n2045 VDD.n2044 9.3005
R26927 VDD.n2047 VDD.n2046 9.3005
R26928 VDD.n2050 VDD.n1405 9.3005
R26929 VDD.n2054 VDD.n2053 9.3005
R26930 VDD.n2056 VDD.n2055 9.3005
R26931 VDD.n2057 VDD.n1403 9.3005
R26932 VDD.n1402 VDD.n1347 9.3005
R26933 VDD.n1401 VDD.n1400 9.3005
R26934 VDD.n1399 VDD.n1348 9.3005
R26935 VDD.n1397 VDD.n1396 9.3005
R26936 VDD.n1395 VDD.n1351 9.3005
R26937 VDD.n1394 VDD.n1393 9.3005
R26938 VDD.n1391 VDD.n1352 9.3005
R26939 VDD.n1390 VDD.n1388 9.3005
R26940 VDD.n1387 VDD.n1357 9.3005
R26941 VDD.n1386 VDD.n1385 9.3005
R26942 VDD.n1384 VDD.n1358 9.3005
R26943 VDD.n1382 VDD.n1381 9.3005
R26944 VDD.n1380 VDD.n1379 9.3005
R26945 VDD.n1377 VDD.n1361 9.3005
R26946 VDD.n1375 VDD.n1374 9.3005
R26947 VDD.n1373 VDD.n1364 9.3005
R26948 VDD.n1372 VDD.n1371 9.3005
R26949 VDD.n1370 VDD.n1365 9.3005
R26950 VDD.n1368 VDD.n1367 9.3005
R26951 VDD.n1263 VDD.n1261 9.3005
R26952 VDD.n2082 VDD.n2081 9.3005
R26953 VDD.n2080 VDD.n2078 9.3005
R26954 VDD.n2071 VDD.n1264 9.3005
R26955 VDD.n2070 VDD.n2069 9.3005
R26956 VDD.n2065 VDD.n1266 9.3005
R26957 VDD.n2064 VDD.n2063 9.3005
R26958 VDD.n2062 VDD.n2061 9.3005
R26959 VDD.n2060 VDD.n1269 9.3005
R26960 VDD.n1340 VDD.n1339 9.3005
R26961 VDD.n1336 VDD.n1272 9.3005
R26962 VDD.n1335 VDD.n1334 9.3005
R26963 VDD.n1333 VDD.n1276 9.3005
R26964 VDD.n1332 VDD.n1331 9.3005
R26965 VDD.n1329 VDD.n1277 9.3005
R26966 VDD.n1328 VDD.n1327 9.3005
R26967 VDD.n1326 VDD.n1325 9.3005
R26968 VDD.n1323 VDD.n1280 9.3005
R26969 VDD.n1322 VDD.n1321 9.3005
R26970 VDD.n1320 VDD.n1319 9.3005
R26971 VDD.n1316 VDD.n1282 9.3005
R26972 VDD.n1315 VDD.n1283 9.3005
R26973 VDD.n1314 VDD.n1313 9.3005
R26974 VDD.n1312 VDD.n1284 9.3005
R26975 VDD.n1311 VDD.n1310 9.3005
R26976 VDD.n1309 VDD.n1285 9.3005
R26977 VDD.n1308 VDD.n1307 9.3005
R26978 VDD.n1306 VDD.n1288 9.3005
R26979 VDD.n1305 VDD.n1304 9.3005
R26980 VDD.n1303 VDD.n1289 9.3005
R26981 VDD.n1302 VDD.n1301 9.3005
R26982 VDD.n861 VDD.n860 9.3005
R26983 VDD.n863 VDD.n862 9.3005
R26984 VDD.n865 VDD.n848 9.3005
R26985 VDD.n868 VDD.n867 9.3005
R26986 VDD.n869 VDD.n847 9.3005
R26987 VDD.n871 VDD.n870 9.3005
R26988 VDD.n872 VDD.n845 9.3005
R26989 VDD.n873 VDD.n844 9.3005
R26990 VDD.n843 VDD.n776 9.3005
R26991 VDD.n842 VDD.n841 9.3005
R26992 VDD.n840 VDD.n777 9.3005
R26993 VDD.n839 VDD.n838 9.3005
R26994 VDD.n837 VDD.n780 9.3005
R26995 VDD.n836 VDD.n835 9.3005
R26996 VDD.n834 VDD.n781 9.3005
R26997 VDD.n833 VDD.n784 9.3005
R26998 VDD.n832 VDD.n831 9.3005
R26999 VDD.n830 VDD.n786 9.3005
R27000 VDD.n829 VDD.n828 9.3005
R27001 VDD.n827 VDD.n787 9.3005
R27002 VDD.n826 VDD.n788 9.3005
R27003 VDD.n825 VDD.n824 9.3005
R27004 VDD.n823 VDD.n790 9.3005
R27005 VDD.n822 VDD.n821 9.3005
R27006 VDD.n818 VDD.n791 9.3005
R27007 VDD.n816 VDD.n815 9.3005
R27008 VDD.n814 VDD.n798 9.3005
R27009 VDD.n813 VDD.n812 9.3005
R27010 VDD.n810 VDD.n799 9.3005
R27011 VDD.n809 VDD.n808 9.3005
R27012 VDD.n807 VDD.n806 9.3005
R27013 VDD.n805 VDD.n803 9.3005
R27014 VDD.n876 VDD.n775 9.3005
R27015 VDD.n878 VDD.n769 9.3005
R27016 VDD.n880 VDD.n879 9.3005
R27017 VDD.n882 VDD.n881 9.3005
R27018 VDD.n883 VDD.n766 9.3005
R27019 VDD.n884 VDD.n765 9.3005
R27020 VDD.n885 VDD.n764 9.3005
R27021 VDD.n886 VDD.n763 9.3005
R27022 VDD.n887 VDD.n760 9.3005
R27023 VDD.n889 VDD.n888 9.3005
R27024 VDD.n890 VDD.n759 9.3005
R27025 VDD.n892 VDD.n891 9.3005
R27026 VDD.n894 VDD.n757 9.3005
R27027 VDD.n895 VDD.n756 9.3005
R27028 VDD.n898 VDD.n897 9.3005
R27029 VDD.n900 VDD.n899 9.3005
R27030 VDD.n901 VDD.n753 9.3005
R27031 VDD.n903 VDD.n902 9.3005
R27032 VDD.n904 VDD.n752 9.3005
R27033 VDD.n906 VDD.n905 9.3005
R27034 VDD.n750 VDD.n748 9.3005
R27035 VDD.n914 VDD.n913 9.3005
R27036 VDD.n915 VDD.n747 9.3005
R27037 VDD.n917 VDD.n916 9.3005
R27038 VDD.n918 VDD.n745 9.3005
R27039 VDD.n921 VDD.n920 9.3005
R27040 VDD.n922 VDD.n744 9.3005
R27041 VDD.n924 VDD.n923 9.3005
R27042 VDD.n928 VDD.n743 9.3005
R27043 VDD.n932 VDD.n931 9.3005
R27044 VDD.n934 VDD.n933 9.3005
R27045 VDD.n936 VDD.n741 9.3005
R27046 VDD.n940 VDD.n939 9.3005
R27047 VDD.n942 VDD.n941 9.3005
R27048 VDD.n943 VDD.n738 9.3005
R27049 VDD.n944 VDD.n736 9.3005
R27050 VDD.n946 VDD.n945 9.3005
R27051 VDD.n947 VDD.n735 9.3005
R27052 VDD.n949 VDD.n948 9.3005
R27053 VDD.n953 VDD.n734 9.3005
R27054 VDD.n958 VDD.n957 9.3005
R27055 VDD.n959 VDD.n733 9.3005
R27056 VDD.n961 VDD.n960 9.3005
R27057 VDD.n962 VDD.n731 9.3005
R27058 VDD.n964 VDD.n963 9.3005
R27059 VDD.n965 VDD.n730 9.3005
R27060 VDD.n967 VDD.n966 9.3005
R27061 VDD.n970 VDD.n729 9.3005
R27062 VDD.n975 VDD.n974 9.3005
R27063 VDD.n976 VDD.n728 9.3005
R27064 VDD.n978 VDD.n977 9.3005
R27065 VDD.n979 VDD.n726 9.3005
R27066 VDD.n980 VDD.n725 9.3005
R27067 VDD.n983 VDD.n982 9.3005
R27068 VDD.n985 VDD.n984 9.3005
R27069 VDD.n986 VDD.n722 9.3005
R27070 VDD.n996 VDD.n995 9.3005
R27071 VDD.n997 VDD.n721 9.3005
R27072 VDD.n999 VDD.n998 9.3005
R27073 VDD.n1000 VDD.n720 9.3005
R27074 VDD.n1003 VDD.n1002 9.3005
R27075 VDD.n1005 VDD.n1004 9.3005
R27076 VDD.n1008 VDD.n717 9.3005
R27077 VDD.n1010 VDD.n1009 9.3005
R27078 VDD.n1012 VDD.n1011 9.3005
R27079 VDD.n1014 VDD.n715 9.3005
R27080 VDD.n1019 VDD.n1018 9.3005
R27081 VDD.n1020 VDD.n714 9.3005
R27082 VDD.n1022 VDD.n1021 9.3005
R27083 VDD.n1023 VDD.n713 9.3005
R27084 VDD.n1027 VDD.n1026 9.3005
R27085 VDD.n1029 VDD.n1028 9.3005
R27086 VDD.n1030 VDD.n709 9.3005
R27087 VDD.n1034 VDD.n1033 9.3005
R27088 VDD.n1035 VDD.n708 9.3005
R27089 VDD.n1037 VDD.n1036 9.3005
R27090 VDD.n1038 VDD.n707 9.3005
R27091 VDD.n1041 VDD.n1040 9.3005
R27092 VDD.n1043 VDD.n1042 9.3005
R27093 VDD.n1044 VDD.n704 9.3005
R27094 VDD.n1046 VDD.n1045 9.3005
R27095 VDD.n1048 VDD.n1047 9.3005
R27096 VDD.n1049 VDD.n700 9.3005
R27097 VDD.n1050 VDD.n699 9.3005
R27098 VDD.n1054 VDD.n1053 9.3005
R27099 VDD.n1056 VDD.n1055 9.3005
R27100 VDD.n1058 VDD.n696 9.3005
R27101 VDD.n1061 VDD.n1060 9.3005
R27102 VDD.n1063 VDD.n1062 9.3005
R27103 VDD.n1065 VDD.n692 9.3005
R27104 VDD.n1067 VDD.n1066 9.3005
R27105 VDD.n1068 VDD.n691 9.3005
R27106 VDD.n1070 VDD.n1069 9.3005
R27107 VDD.n1071 VDD.n689 9.3005
R27108 VDD.n1073 VDD.n1072 9.3005
R27109 VDD.n1074 VDD.n688 9.3005
R27110 VDD.n1076 VDD.n1075 9.3005
R27111 VDD.n1078 VDD.n686 9.3005
R27112 VDD.n1080 VDD.n1079 9.3005
R27113 VDD.n1081 VDD.n685 9.3005
R27114 VDD.n1083 VDD.n1082 9.3005
R27115 VDD.n1084 VDD.n684 9.3005
R27116 VDD.n1085 VDD.n682 9.3005
R27117 VDD.n1087 VDD.n1086 9.3005
R27118 VDD.n1088 VDD.n681 9.3005
R27119 VDD.n1090 VDD.n1089 9.3005
R27120 VDD.n1091 VDD.n679 9.3005
R27121 VDD.n1093 VDD.n1092 9.3005
R27122 VDD.n1094 VDD.n678 9.3005
R27123 VDD.n1096 VDD.n1095 9.3005
R27124 VDD.n1098 VDD.n675 9.3005
R27125 VDD.n1099 VDD.n674 9.3005
R27126 VDD.n1101 VDD.n1100 9.3005
R27127 VDD.n1102 VDD.n673 9.3005
R27128 VDD.n1104 VDD.n1103 9.3005
R27129 VDD.n1105 VDD.n670 9.3005
R27130 VDD.n1109 VDD.n1108 9.3005
R27131 VDD.n1110 VDD.n669 9.3005
R27132 VDD.n1112 VDD.n1111 9.3005
R27133 VDD.n1114 VDD.n668 9.3005
R27134 VDD.n1116 VDD.n1115 9.3005
R27135 VDD.n1119 VDD.n1118 9.3005
R27136 VDD.n1117 VDD.n665 9.3005
R27137 VDD.n1124 VDD.n663 9.3005
R27138 VDD.n1127 VDD.n1126 9.3005
R27139 VDD.n1130 VDD.n1129 9.3005
R27140 VDD.n1131 VDD.n656 9.3005
R27141 VDD.n1135 VDD.n1134 9.3005
R27142 VDD.n1136 VDD.n655 9.3005
R27143 VDD.n1138 VDD.n1137 9.3005
R27144 VDD.n1139 VDD.n653 9.3005
R27145 VDD.n1140 VDD.n652 9.3005
R27146 VDD.n1141 VDD.n651 9.3005
R27147 VDD.n1143 VDD.n644 9.3005
R27148 VDD.n1144 VDD.n643 9.3005
R27149 VDD.n1148 VDD.n1147 9.3005
R27150 VDD.n1150 VDD.n1149 9.3005
R27151 VDD.n1151 VDD.n641 9.3005
R27152 VDD.n1152 VDD.n639 9.3005
R27153 VDD.n1153 VDD.n631 9.3005
R27154 VDD.n1158 VDD.n1157 9.3005
R27155 VDD.n1159 VDD.n624 9.3005
R27156 VDD.n1162 VDD.n1161 9.3005
R27157 VDD.n1164 VDD.n1163 9.3005
R27158 VDD.n1165 VDD.n622 9.3005
R27159 VDD.n1169 VDD.n1168 9.3005
R27160 VDD.n1170 VDD.n621 9.3005
R27161 VDD.n1172 VDD.n1171 9.3005
R27162 VDD.n1174 VDD.n620 9.3005
R27163 VDD.n1178 VDD.n1177 9.3005
R27164 VDD.n1180 VDD.n1179 9.3005
R27165 VDD.n1181 VDD.n617 9.3005
R27166 VDD.n1184 VDD.n1183 9.3005
R27167 VDD.n1186 VDD.n1185 9.3005
R27168 VDD.n1187 VDD.n615 9.3005
R27169 VDD.n1188 VDD.n612 9.3005
R27170 VDD.n1190 VDD.n1189 9.3005
R27171 VDD.n1191 VDD.n611 9.3005
R27172 VDD.n1193 VDD.n1192 9.3005
R27173 VDD.n1195 VDD.n609 9.3005
R27174 VDD.n1198 VDD.n1197 9.3005
R27175 VDD.n1200 VDD.n1199 9.3005
R27176 VDD.n1201 VDD.n605 9.3005
R27177 VDD.n1202 VDD.n604 9.3005
R27178 VDD.n1204 VDD.n1203 9.3005
R27179 VDD.n1205 VDD.n603 9.3005
R27180 VDD.n1207 VDD.n1206 9.3005
R27181 VDD.n1208 VDD.n602 9.3005
R27182 VDD.n1209 VDD.n601 9.3005
R27183 VDD.n1210 VDD.n599 9.3005
R27184 VDD.n1212 VDD.n1211 9.3005
R27185 VDD.n1213 VDD.n598 9.3005
R27186 VDD.n1215 VDD.n1214 9.3005
R27187 VDD.n1216 VDD.n596 9.3005
R27188 VDD.n1219 VDD.n1218 9.3005
R27189 VDD.n1220 VDD.n595 9.3005
R27190 VDD.n1222 VDD.n1221 9.3005
R27191 VDD.n1225 VDD.n1224 9.3005
R27192 VDD.n1226 VDD.n589 9.3005
R27193 VDD.n1228 VDD.n1227 9.3005
R27194 VDD.n1229 VDD.n587 9.3005
R27195 VDD.n586 VDD.n530 9.3005
R27196 VDD.n585 VDD.n584 9.3005
R27197 VDD.n583 VDD.n531 9.3005
R27198 VDD.n581 VDD.n580 9.3005
R27199 VDD.n579 VDD.n578 9.3005
R27200 VDD.n576 VDD.n536 9.3005
R27201 VDD.n575 VDD.n574 9.3005
R27202 VDD.n573 VDD.n539 9.3005
R27203 VDD.n572 VDD.n571 9.3005
R27204 VDD.n570 VDD.n540 9.3005
R27205 VDD.n569 VDD.n568 9.3005
R27206 VDD.n567 VDD.n541 9.3005
R27207 VDD.n566 VDD.n565 9.3005
R27208 VDD.n563 VDD.n542 9.3005
R27209 VDD.n561 VDD.n560 9.3005
R27210 VDD.n559 VDD.n548 9.3005
R27211 VDD.n558 VDD.n557 9.3005
R27212 VDD.n556 VDD.n549 9.3005
R27213 VDD.n554 VDD.n553 9.3005
R27214 VDD.n551 VDD.n442 9.3005
R27215 VDD.n1252 VDD.n1251 9.3005
R27216 VDD.n1249 VDD.n1248 9.3005
R27217 VDD.n1241 VDD.n1240 9.3005
R27218 VDD.n1238 VDD.n448 9.3005
R27219 VDD.n1237 VDD.n1236 9.3005
R27220 VDD.n1235 VDD.n451 9.3005
R27221 VDD.n1234 VDD.n1233 9.3005
R27222 VDD.n1232 VDD.n452 9.3005
R27223 VDD.n528 VDD.n527 9.3005
R27224 VDD.n525 VDD.n524 9.3005
R27225 VDD.n523 VDD.n460 9.3005
R27226 VDD.n521 VDD.n520 9.3005
R27227 VDD.n519 VDD.n465 9.3005
R27228 VDD.n518 VDD.n517 9.3005
R27229 VDD.n516 VDD.n466 9.3005
R27230 VDD.n515 VDD.n468 9.3005
R27231 VDD.n514 VDD.n513 9.3005
R27232 VDD.n512 VDD.n470 9.3005
R27233 VDD.n511 VDD.n510 9.3005
R27234 VDD.n509 VDD.n471 9.3005
R27235 VDD.n508 VDD.n507 9.3005
R27236 VDD.n506 VDD.n474 9.3005
R27237 VDD.n505 VDD.n504 9.3005
R27238 VDD.n503 VDD.n475 9.3005
R27239 VDD.n502 VDD.n501 9.3005
R27240 VDD.n500 VDD.n478 9.3005
R27241 VDD.n499 VDD.n498 9.3005
R27242 VDD.n496 VDD.n479 9.3005
R27243 VDD.n494 VDD.n493 9.3005
R27244 VDD.n492 VDD.n491 9.3005
R27245 VDD.n428 VDD.n427 9.3005
R27246 VDD.n422 VDD.n414 9.3005
R27247 VDD.n420 VDD.n419 9.3005
R27248 VDD.n433 VDD.n332 9.3005
R27249 VDD.n435 VDD.n434 9.3005
R27250 VDD.n409 VDD.n331 9.3005
R27251 VDD.n408 VDD.n407 9.3005
R27252 VDD.n236 VDD.n222 9.3005
R27253 VDD.n167 VDD.n166 9.3005
R27254 VDD.n100 VDD.n90 9.3005
R27255 VDD.n96 VDD.n91 9.3005
R27256 VDD.n98 VDD.n97 9.3005
R27257 VDD.n53 VDD.n46 9.3005
R27258 VDD.n61 VDD.n60 9.3005
R27259 VDD.n59 VDD.n47 9.3005
R27260 VDD.n58 VDD.n57 9.3005
R27261 VDD.n25 VDD.n24 9.3005
R27262 VDD.n21 VDD.n10 9.3005
R27263 VDD.n17 VDD.n14 9.3005
R27264 VDD.n20 VDD.n18 9.3005
R27265 VDD.n2514 VDD.n2513 9.20381
R27266 VDD.n3721 VDD.n3719 9.09802
R27267 VDD.n4152 VDD.n4149 9.09802
R27268 VDD.n4159 VDD.n3712 9.09802
R27269 VDD.n3907 VDD.n3906 9.09802
R27270 VDD.n4330 VDD.n4323 9.09802
R27271 VDD.n4446 VDD.n3670 9.09802
R27272 VDD.n4273 VDD.n4272 9.09802
R27273 VDD.n4045 VDD.n4044 9.09802
R27274 VDD.n3929 VDD.n3810 9.09802
R27275 VDD.n3942 VDD.n3941 9.09802
R27276 VDD.n4437 VDD.n4368 9.09802
R27277 VDD.n4423 VDD.n4376 9.09802
R27278 VDD.n2186 VDD.n2177 9.09802
R27279 VDD.n2872 VDD.n2099 9.09802
R27280 VDD.n2520 VDD.n2519 9.09802
R27281 VDD.n1600 VDD.n1599 9.09802
R27282 VDD.n1319 VDD.n1318 9.09802
R27283 VDD.n432 VDD.n431 9.0663
R27284 VDD.n3501 VDD.n3500 9.03579
R27285 VDD.n3473 VDD.n3472 9.03579
R27286 VDD.n3401 VDD.n3400 9.03579
R27287 VDD.n3318 VDD.n2981 9.03579
R27288 VDD.n3311 VDD.n2984 9.03579
R27289 VDD.n3554 VDD.n3527 9.03579
R27290 VDD.n3547 VDD.n3530 9.03579
R27291 VDD.n2747 VDD.n2266 9.03579
R27292 VDD.n1877 VDD.n1876 9.03579
R27293 VDD.n1758 VDD.n1757 9.03579
R27294 VDD.n1152 VDD.n1151 9.03579
R27295 VDD.n828 VDD.n786 9.03579
R27296 VDD.n827 VDD.n826 9.03579
R27297 VDD.n2510 VDD.n2509 8.99224
R27298 VDD.n4298 VDD.n3679 8.88645
R27299 VDD.n2680 VDD.n2679 8.88645
R27300 VDD.n2613 VDD.n2612 8.78066
R27301 VDD.n4157 VDD.n4156 8.67488
R27302 VDD.n2660 VDD.n2659 8.67488
R27303 VDD.n4100 VDD.n4099 8.65932
R27304 VDD.n3277 VDD.n3275 8.65932
R27305 VDD.n2567 VDD.n2566 8.62646
R27306 VDD.n967 VDD.n730 8.62646
R27307 VDD.n4296 VDD.n4295 8.56909
R27308 VDD.n3901 VDD.n3817 8.44958
R27309 VDD.n4294 VDD.n3681 8.44958
R27310 VDD.n2495 VDD.n2398 8.44958
R27311 VDD.n1608 VDD.n1607 8.44958
R27312 VDD.t1264 VDD.t1266 8.39273
R27313 VDD.t1767 VDD.t2014 8.39273
R27314 VDD.t2774 VDD.t3074 8.39273
R27315 VDD.t663 VDD.t379 8.39273
R27316 VDD.t1175 VDD.t469 8.39273
R27317 VDD.t2707 VDD.t2544 8.39273
R27318 VDD.t1099 VDD.t2859 8.39273
R27319 VDD.t1755 VDD.n3422 8.39273
R27320 VDD.t74 VDD.t1902 8.39273
R27321 VDD.t1495 VDD.t1677 8.39273
R27322 VDD.t82 VDD.t490 8.39273
R27323 VDD.t1497 VDD.t1194 8.39273
R27324 VDD.t1648 VDD.t1025 8.39273
R27325 VDD.t2059 VDD.t331 8.39273
R27326 VDD.t362 VDD.t1633 8.39273
R27327 VDD.t1733 VDD.t2652 8.39273
R27328 VDD.t2171 VDD.n613 8.39273
R27329 VDD.t2163 VDD.t765 8.39273
R27330 VDD.t767 VDD.t3083 8.39273
R27331 VDD.t699 VDD.t1636 8.39273
R27332 VDD.n2615 VDD.n2329 8.35752
R27333 VDD.n4048 VDD.n3758 8.28285
R27334 VDD.n3283 VDD.n3281 8.28285
R27335 VDD.n3228 VDD.n3227 8.28285
R27336 VDD.n166 VDD.n162 8.28285
R27337 VDD.n93 VDD.n91 8.28285
R27338 VDD.n99 VDD.n98 8.28285
R27339 VDD.n205 VDD.n204 8.27619
R27340 VDD.n69 VDD.n65 8.22907
R27341 VDD.n41 VDD.n29 8.22907
R27342 VDD.n2817 VDD.n2814 7.94989
R27343 VDD.n4242 VDD.n4241 7.93422
R27344 VDD.n3959 VDD.n3800 7.93422
R27345 VDD.n1125 VDD.n662 7.93422
R27346 VDD.n1686 VDD.n1685 7.90638
R27347 VDD.n3126 VDD.n3071 7.85911
R27348 VDD.n4040 VDD.n3760 7.75995
R27349 VDD.n2607 VDD.n2332 7.75995
R27350 VDD.n1329 VDD.n1328 7.75995
R27351 VDD.n2828 VDD.n2233 7.72281
R27352 VDD.n636 VDD.n635 7.58311
R27353 VDD.n4362 VDD.n4361 7.52991
R27354 VDD.n3953 VDD.n3952 7.52991
R27355 VDD.n1909 VDD.n1908 7.52991
R27356 VDD.n2848 VDD.n2223 7.48358
R27357 VDD.n3796 VDD.n3794 7.42178
R27358 VDD.n72 VDD.n71 7.4005
R27359 VDD.n76 VDD.n75 7.4005
R27360 VDD.n39 VDD.n38 7.4005
R27361 VDD.n35 VDD.n34 7.4005
R27362 VDD.n409 VDD.n408 7.3605
R27363 VDD.n434 VDD.n409 7.3605
R27364 VDD.n434 VDD.n433 7.3605
R27365 VDD.n1120 VDD.n666 7.28326
R27366 VDD.n3799 VDD.n3797 7.25383
R27367 VDD.n4238 VDD.n4237 7.23528
R27368 VDD.n2374 VDD.n2371 7.23528
R27369 VDD.n659 VDD.n657 7.23528
R27370 VDD.n912 VDD.n911 7.22943
R27371 VDD.n4092 VDD.n3744 7.15344
R27372 VDD.n3863 VDD.n3836 7.15344
R27373 VDD.n4337 VDD.n4319 7.15344
R27374 VDD.n3426 VDD.n3425 7.15344
R27375 VDD.n3568 VDD.n3567 7.15344
R27376 VDD.n2586 VDD.n2585 7.15344
R27377 VDD.n1835 VDD.n1511 7.15344
R27378 VDD.n1781 VDD.n1780 7.15344
R27379 VDD.n1040 VDD.n706 7.15344
R27380 VDD.n426 VDD.n425 7.13298
R27381 VDD.n4026 VDD.n4025 7.12524
R27382 VDD.n319 VDD.n318 7.11588
R27383 VDD.n324 VDD.n323 7.11588
R27384 VDD.n2643 VDD.n2307 6.95702
R27385 VDD.n2375 VDD.n2371 6.95702
R27386 VDD.n164 VDD.n163 6.91098
R27387 VDD.n150 VDD.n149 6.9065
R27388 VDD.n382 VDD.t1731 6.84014
R27389 VDD.n380 VDD.t1725 6.84014
R27390 VDD.n379 VDD.t1727 6.84014
R27391 VDD.n165 VDD.n164 6.8072
R27392 VDD.n3988 VDD.n3985 6.8005
R27393 VDD.n2577 VDD.n2574 6.8005
R27394 VDD.n2533 VDD.n2530 6.8005
R27395 VDD.n3468 VDD.n2944 6.77697
R27396 VDD.n1354 VDD.n1351 6.77697
R27397 VDD.n2008 VDD.n2007 6.77697
R27398 VDD.n1957 VDD.n1956 6.77697
R27399 VDD.n1911 VDD.n1910 6.77697
R27400 VDD.n1828 VDD.n1515 6.77697
R27401 VDD.n1694 VDD.n1568 6.77697
R27402 VDD.n1698 VDD.n1697 6.77697
R27403 VDD.n1709 VDD.n1563 6.77697
R27404 VDD.n1182 VDD.n1181 6.77697
R27405 VDD.n1009 VDD.n716 6.77697
R27406 VDD.n937 VDD.n936 6.77697
R27407 VDD.n423 VDD.n422 6.77697
R27408 VDD.n2496 VDD.n2396 6.77075
R27409 VDD.n1115 VDD.n667 6.73838
R27410 VDD.n95 VDD.n94 6.73566
R27411 VDD.t205 VDD.t1111 6.71428
R27412 VDD.t1280 VDD.t2983 6.71428
R27413 VDD.t2135 VDD.t1539 6.71428
R27414 VDD.t396 VDD.t1207 6.71428
R27415 VDD.t949 VDD.t1851 6.71428
R27416 VDD.t535 VDD.t225 6.71428
R27417 VDD.t391 VDD.t1459 6.71428
R27418 VDD.t408 VDD.t2981 6.71428
R27419 VDD.t1481 VDD.t2821 6.71428
R27420 VDD.t2701 VDD.t2670 6.71428
R27421 VDD.t1208 VDD.t197 6.71428
R27422 VDD.t360 VDD.t2236 6.71428
R27423 VDD.t2971 VDD.t1691 6.71428
R27424 VDD.t1771 VDD.t2391 6.71428
R27425 VDD.t1914 VDD.t1775 6.71428
R27426 VDD.t1438 VDD.t1930 6.71428
R27427 VDD.t256 VDD.t1734 6.71428
R27428 VDD.t2656 VDD.t236 6.71428
R27429 VDD.t3067 VDD.t1096 6.71428
R27430 VDD.n2837 VDD.n2836 6.66496
R27431 VDD.n2501 VDD.n2500 6.66496
R27432 VDD.n1677 VDD.n1574 6.66496
R27433 VDD.n2441 VDD.n2440 6.52104
R27434 VDD.n1614 VDD.n1613 6.52104
R27435 VDD.n78 VDD.n64 6.49269
R27436 VDD.n28 VDD.n27 6.49269
R27437 VDD.n4241 VDD.n4240 6.48583
R27438 VDD.n3800 VDD.n3799 6.48583
R27439 VDD.n1681 VDD.n1680 6.48583
R27440 VDD.n662 VDD.n661 6.48583
R27441 VDD.n1053 VDD.n1051 6.41951
R27442 VDD.n4104 VDD.n4103 6.4005
R27443 VDD.n3378 VDD.n3377 6.4005
R27444 VDD.n3338 VDD.n2971 6.4005
R27445 VDD.n3297 VDD.n2991 6.4005
R27446 VDD.n3645 VDD.n3644 6.4005
R27447 VDD.n2740 VDD.n2268 6.4005
R27448 VDD.n2687 VDD.n2686 6.4005
R27449 VDD.n1951 VDD.n1449 6.4005
R27450 VDD.n1825 VDD.n1824 6.4005
R27451 VDD.n1699 VDD.n1698 6.4005
R27452 VDD.n1739 VDD.n1552 6.4005
R27453 VDD.n1098 VDD.n1097 6.4005
R27454 VDD.n987 VDD.n986 6.4005
R27455 VDD.n278 VDD.n248 6.28433
R27456 VDD.n2644 VDD.n2307 6.26137
R27457 VDD.n1630 VDD.n1584 6.18951
R27458 VDD.n3387 VDD.n3385 6.02403
R27459 VDD.n3331 VDD.n3330 6.02403
R27460 VDD.n3652 VDD.n2899 6.02403
R27461 VDD.n3169 VDD.n3167 6.02403
R27462 VDD.n3173 VDD.n3027 6.02403
R27463 VDD.n1716 VDD.n1715 6.02403
R27464 VDD.n1719 VDD.n1718 6.02403
R27465 VDD.n1140 VDD.n1139 6.02403
R27466 VDD.n1078 VDD.n1077 6.02403
R27467 VDD.n3135 VDD.n3039 5.98311
R27468 VDD.n278 VDD.n277 5.94683
R27469 VDD.n280 VDD.n279 5.94683
R27470 VDD.n284 VDD.n245 5.94683
R27471 VDD.n290 VDD.n289 5.94683
R27472 VDD.n292 VDD.n291 5.94683
R27473 VDD.n296 VDD.n242 5.94683
R27474 VDD.n302 VDD.n301 5.94683
R27475 VDD.n304 VDD.n303 5.94683
R27476 VDD.n308 VDD.n237 5.94683
R27477 VDD.n314 VDD.n313 5.94683
R27478 VDD.n4239 VDD.n4185 5.8885
R27479 VDD.n660 VDD.n658 5.8885
R27480 VDD.n79 VDD.n63 5.80439
R27481 VDD.n43 VDD.n42 5.80403
R27482 VDD.n169 VDD.n87 5.80248
R27483 VDD.n274 VDD.n273 5.78447
R27484 VDD.n276 VDD.n247 5.78447
R27485 VDD.n282 VDD.n281 5.78447
R27486 VDD.n285 VDD.n283 5.78447
R27487 VDD.n288 VDD.n244 5.78447
R27488 VDD.n294 VDD.n293 5.78447
R27489 VDD.n297 VDD.n295 5.78447
R27490 VDD.n300 VDD.n241 5.78447
R27491 VDD.n306 VDD.n305 5.78447
R27492 VDD.n309 VDD.n307 5.78447
R27493 VDD.n312 VDD.n239 5.78447
R27494 VDD.n144 VDD.n137 5.78175
R27495 VDD.n137 VDD.n136 5.78175
R27496 VDD.n108 VDD.n106 5.78175
R27497 VDD.n136 VDD.n108 5.78175
R27498 VDD.n118 VDD.n107 5.78175
R27499 VDD.n133 VDD.n107 5.78175
R27500 VDD.n134 VDD.n133 5.78175
R27501 VDD.n3892 VDD.n3891 5.66204
R27502 VDD.n3894 VDD.n3892 5.66204
R27503 VDD.n3898 VDD.n3819 5.66204
R27504 VDD.n3899 VDD.n3898 5.66204
R27505 VDD.n4283 VDD.n4282 5.66204
R27506 VDD.n4284 VDD.n4283 5.66204
R27507 VDD.n4288 VDD.n4287 5.66204
R27508 VDD.n4290 VDD.n4288 5.66204
R27509 VDD.n3124 VDD.n3123 5.66204
R27510 VDD.n3118 VDD.n3117 5.66204
R27511 VDD.n3117 VDD.n3075 5.66204
R27512 VDD.n3113 VDD.n3075 5.66204
R27513 VDD.n3113 VDD.n3112 5.66204
R27514 VDD.n3112 VDD.n3111 5.66204
R27515 VDD.n3101 VDD.n3100 5.66204
R27516 VDD.n3095 VDD.n3094 5.66204
R27517 VDD.n3094 VDD.n3093 5.66204
R27518 VDD.n3093 VDD.n3083 5.66204
R27519 VDD.n3089 VDD.n3083 5.66204
R27520 VDD.n3089 VDD.n3088 5.66204
R27521 VDD.n3633 VDD.n3632 5.66204
R27522 VDD.n3632 VDD.n3631 5.66204
R27523 VDD.n3628 VDD.n3627 5.66204
R27524 VDD.n3627 VDD.n3626 5.66204
R27525 VDD.n3626 VDD.n3587 5.66204
R27526 VDD.n3622 VDD.n3587 5.66204
R27527 VDD.n3622 VDD.n3621 5.66204
R27528 VDD.n3621 VDD.n3620 5.66204
R27529 VDD.n2438 VDD.n2413 5.66204
R27530 VDD.n2430 VDD.n2416 5.66204
R27531 VDD.n2426 VDD.n2416 5.66204
R27532 VDD.n2424 VDD.n2423 5.66204
R27533 VDD.n2423 VDD.n2419 5.66204
R27534 VDD.n4053 VDD.n3758 5.64756
R27535 VDD.n2627 VDD.n2626 5.64756
R27536 VDD.n1237 VDD.n451 5.64756
R27537 VDD.n887 VDD.n886 5.64756
R27538 VDD.n3669 VDD.n3666 5.60711
R27539 VDD.n2180 VDD.n2093 5.60711
R27540 VDD.n2874 VDD.n2873 5.60711
R27541 VDD.n1337 VDD.n1275 5.60687
R27542 VDD.n3108 VDD.n3107 5.48759
R27543 VDD.n3105 VDD.n3104 5.42606
R27544 VDD.n4142 VDD.n4141 5.40233
R27545 VDD.n4267 VDD.n3687 5.40233
R27546 VDD.n3915 VDD.n3914 5.40233
R27547 VDD.n398 VDD.n397 5.34555
R27548 VDD.n3891 VDD.n3821 5.29281
R27549 VDD.n3900 VDD.n3899 5.29281
R27550 VDD.n4282 VDD.n3685 5.29281
R27551 VDD.n4290 VDD.n4289 5.29281
R27552 VDD.n3125 VDD.n3124 5.29281
R27553 VDD.n3111 VDD.n3077 5.29281
R27554 VDD.n3101 VDD.n3079 5.29281
R27555 VDD.n3088 VDD.n3087 5.29281
R27556 VDD.n3633 VDD.n3583 5.29281
R27557 VDD.n3620 VDD.n3589 5.29281
R27558 VDD.n2439 VDD.n2438 5.29281
R27559 VDD.n2415 VDD.n2413 5.29281
R27560 VDD.n2431 VDD.n2430 5.29281
R27561 VDD.n2419 VDD.n2418 5.29281
R27562 VDD.n1612 VDD.n1611 5.29281
R27563 VDD.n1611 VDD.n1591 5.29281
R27564 VDD.n1683 VDD.n1682 5.29117
R27565 VDD.n4460 VDD.n4459 5.28976
R27566 VDD.n2184 VDD.n2183 5.28976
R27567 VDD.n2875 VDD.n2098 5.28976
R27568 VDD.n1154 VDD.n637 5.28746
R27569 VDD.n908 VDD.n907 5.28746
R27570 VDD.n4208 VDD.n4198 5.27109
R27571 VDD.n2622 VDD.n2327 5.27109
R27572 VDD.n894 VDD.n893 5.27109
R27573 VDD.n1342 VDD.n1271 5.25888
R27574 VDD.n4144 VDD.n3717 5.18397
R27575 VDD.n4327 VDD.n4325 5.18397
R27576 VDD.n4434 VDD.n4370 5.18397
R27577 VDD.n2183 VDD.n2181 5.18397
R27578 VDD.n2667 VDD.n2666 5.18397
R27579 VDD.n406 VDD.n405 5.14633
R27580 VDD.n239 VDD.n238 5.063
R27581 VDD.n311 VDD.n223 5.058
R27582 VDD.n315 VDD.n314 5.05712
R27583 VDD.n2107 VDD.n2106 5.05557
R27584 VDD.t1815 VDD.t1689 5.03584
R27585 VDD.t701 VDD.t2879 5.03584
R27586 VDD.t994 VDD.t1969 5.03584
R27587 VDD.t1350 VDD.t564 5.03584
R27588 VDD.t2587 VDD.t2709 5.03584
R27589 VDD.t1206 VDD.t119 5.03584
R27590 VDD.t2532 VDD.t2231 5.03584
R27591 VDD.t1133 VDD.t2317 5.03584
R27592 VDD.n2648 VDD.n2647 5.03517
R27593 VDD.n1344 VDD.n1268 5.03517
R27594 VDD.n4278 VDD.n4277 5.03171
R27595 VDD.n2599 VDD.n2598 5.00648
R27596 VDD.n4142 VDD.n3719 4.9724
R27597 VDD.n4273 VDD.n3687 4.9724
R27598 VDD.n2831 VDD.n2231 4.9724
R27599 VDD.n3504 VDD.n3503 4.89462
R27600 VDD.n3314 VDD.n3313 4.89462
R27601 VDD.n3552 VDD.n3551 4.89462
R27602 VDD.n2629 VDD.n2628 4.89462
R27603 VDD.n2016 VDD.n2015 4.89462
R27604 VDD.n1985 VDD.n1984 4.89462
R27605 VDD.n1857 VDD.n1504 4.89462
R27606 VDD.n1761 VDD.n1760 4.89462
R27607 VDD.n563 VDD.n562 4.89462
R27608 VDD.n1224 VDD.n589 4.89462
R27609 VDD.n1085 VDD.n1084 4.89462
R27610 VDD.n980 VDD.n979 4.89462
R27611 VDD.n2668 VDD.n2300 4.86662
R27612 VDD.n2671 VDD.n2300 4.86662
R27613 VDD.n275 VDD.n274 4.838
R27614 VDD.n273 VDD.n272 4.813
R27615 VDD.n636 VDD.n632 4.8005
R27616 VDD.n1274 VDD.n1273 4.77455
R27617 VDD.n4143 VDD.n4142 4.76083
R27618 VDD.n4276 VDD.n3687 4.76083
R27619 VDD.n3055 VDD.n3047 4.75752
R27620 VDD.n3856 VDD.n3855 4.75748
R27621 VDD.n3606 VDD.n3598 4.75748
R27622 VDD.n2481 VDD.n2473 4.75748
R27623 VDD.n2134 VDD.n2126 4.75748
R27624 VDD.n1663 VDD.n1655 4.75748
R27625 VDD.n1300 VDD.n1292 4.75748
R27626 VDD.n234 VDD.n222 4.70477
R27627 VDD.n4220 VDD.n4219 4.67352
R27628 VDD.n4217 VDD.n4194 4.67352
R27629 VDD.n4233 VDD.n4232 4.67352
R27630 VDD.n4080 VDD.n3750 4.67352
R27631 VDD.n4355 VDD.n4354 4.67352
R27632 VDD.n4354 VDD.n4313 4.67352
R27633 VDD.n4258 VDD.n3694 4.67352
R27634 VDD.n4259 VDD.n4258 4.67352
R27635 VDD.n4020 VDD.n4017 4.67352
R27636 VDD.n4064 VDD.n4059 4.67352
R27637 VDD.n3967 VDD.n3966 4.67352
R27638 VDD.n3958 VDD.n3957 4.67352
R27639 VDD.n3960 VDD.n3958 4.67352
R27640 VDD.n3409 VDD.n3408 4.67352
R27641 VDD.n3253 VDD.n3245 4.67352
R27642 VDD.n3141 VDD.n3037 4.67352
R27643 VDD.n3142 VDD.n3141 4.67352
R27644 VDD.n3194 VDD.n3019 4.67352
R27645 VDD.n2842 VDD.n2224 4.67352
R27646 VDD.n2846 VDD.n2224 4.67352
R27647 VDD.n2821 VDD.n2235 4.67352
R27648 VDD.n2728 VDD.n2274 4.67352
R27649 VDD.n2706 VDD.n2285 4.67352
R27650 VDD.n2698 VDD.n2697 4.67352
R27651 VDD.n2651 VDD.n2304 4.67352
R27652 VDD.n2655 VDD.n2304 4.67352
R27653 VDD.n2559 VDD.n2367 4.67352
R27654 VDD.n2563 VDD.n2367 4.67352
R27655 VDD.n2550 VDD.n2549 4.67352
R27656 VDD.n2065 VDD.n2064 4.67352
R27657 VDD.n1925 VDD.n1924 4.67352
R27658 VDD.n1929 VDD.n1928 4.67352
R27659 VDD.n1854 VDD.n1506 4.67352
R27660 VDD.n584 VDD.n583 4.67352
R27661 VDD.n1172 VDD.n621 4.67352
R27662 VDD.n1177 VDD.n1174 4.67352
R27663 VDD.n1159 VDD.n1158 4.67352
R27664 VDD.n1131 VDD.n1130 4.67352
R27665 VDD.n1126 VDD.n1124 4.67352
R27666 VDD.n1112 VDD.n669 4.67352
R27667 VDD.n1115 VDD.n1114 4.67352
R27668 VDD.n1022 VDD.n714 4.67352
R27669 VDD.n1023 VDD.n1022 4.67352
R27670 VDD.n999 VDD.n721 4.67352
R27671 VDD.n1000 VDD.n999 4.67352
R27672 VDD.n974 VDD.n970 4.67352
R27673 VDD.n957 VDD.n953 4.67352
R27674 VDD.n931 VDD.n928 4.67352
R27675 VDD.n913 VDD.n747 4.67352
R27676 VDD.n917 VDD.n747 4.67352
R27677 VDD.n918 VDD.n917 4.67352
R27678 VDD.n816 VDD.n798 4.67352
R27679 VDD.n812 VDD.n798 4.67352
R27680 VDD.n810 VDD.n809 4.67352
R27681 VDD.n524 VDD.n523 4.67352
R27682 VDD.n4076 VDD.n4075 4.62272
R27683 VDD.n2592 VDD.n2347 4.62124
R27684 VDD.n907 VDD.n751 4.62124
R27685 VDD.n1155 VDD.n1154 4.62124
R27686 VDD.n3962 VDD.n3800 4.62124
R27687 VDD.n3963 VDD.n3794 4.62124
R27688 VDD.n4241 VDD.n4184 4.62124
R27689 VDD.n2499 VDD.n2498 4.62124
R27690 VDD.n1680 VDD.n1679 4.62124
R27691 VDD.n1342 VDD.n1341 4.62124
R27692 VDD.n1128 VDD.n662 4.62124
R27693 VDD.n398 VDD.n396 4.60988
R27694 VDD.n403 VDD.n402 4.60206
R27695 VDD.n454 VDD.n453 4.5918
R27696 VDD.n4262 VDD.n4260 4.57193
R27697 VDD.n2790 VDD.n2789 4.57193
R27698 VDD.n2159 VDD.n2158 4.57193
R27699 VDD.n812 VDD.n811 4.57193
R27700 VDD.n4243 VDD.n4242 4.56405
R27701 VDD.n3960 VDD.n3959 4.56405
R27702 VDD.n1126 VDD.n1125 4.56405
R27703 VDD.n4147 VDD.n3717 4.54926
R27704 VDD.n4325 VDD.n3664 4.54926
R27705 VDD.n2181 VDD.n2180 4.54926
R27706 VDD.n2836 VDD.n2231 4.54926
R27707 VDD.n2668 VDD.n2667 4.54926
R27708 VDD.n2507 VDD.n2394 4.54926
R27709 VDD.n1605 VDD.n1604 4.54926
R27710 VDD.n2596 VDD.n2337 4.54244
R27711 VDD.n2650 VDD.n2649 4.52113
R27712 VDD.n2762 VDD.n2761 4.51815
R27713 VDD.n1819 VDD.n1818 4.51815
R27714 VDD.n1703 VDD.n1701 4.51815
R27715 VDD.n835 VDD.n834 4.51815
R27716 VDD.n4465 VDD.n3660 4.51401
R27717 VDD.n4457 VDD.n4456 4.51401
R27718 VDD.n3656 VDD.n2894 4.51401
R27719 VDD.n2908 VDD.n2907 4.51401
R27720 VDD.n2890 VDD.n2089 4.51401
R27721 VDD.n2883 VDD.n2882 4.51401
R27722 VDD.n2085 VDD.n1259 4.51401
R27723 VDD.n2077 VDD.n2076 4.51401
R27724 VDD.n1255 VDD.n440 4.51401
R27725 VDD.n1247 VDD.n1246 4.51401
R27726 VDD.n208 VDD.n189 4.5127
R27727 VDD.n215 VDD.n214 4.5127
R27728 VDD.n4464 VDD.n4463 4.5005
R27729 VDD.n4452 VDD.n3663 4.5005
R27730 VDD.n4455 VDD.n3667 4.5005
R27731 VDD.n3655 VDD.n3654 4.5005
R27732 VDD.n2902 VDD.n2897 4.5005
R27733 VDD.n2906 VDD.n2905 4.5005
R27734 VDD.n2889 VDD.n2888 4.5005
R27735 VDD.n2878 VDD.n2092 4.5005
R27736 VDD.n2881 VDD.n2095 4.5005
R27737 VDD.n2084 VDD.n2083 4.5005
R27738 VDD.n2072 VDD.n1262 4.5005
R27739 VDD.n2075 VDD.n1265 4.5005
R27740 VDD.n1254 VDD.n1253 4.5005
R27741 VDD.n1242 VDD.n443 4.5005
R27742 VDD.n1245 VDD.n447 4.5005
R27743 VDD.n430 VDD.n413 4.5005
R27744 VDD.n430 VDD.n429 4.5005
R27745 VDD.n400 VDD.n399 4.5005
R27746 VDD.n401 VDD.n395 4.5005
R27747 VDD.n305 VDD.n240 4.5005
R27748 VDD.n300 VDD.n299 4.5005
R27749 VDD.n298 VDD.n297 4.5005
R27750 VDD.n293 VDD.n243 4.5005
R27751 VDD.n288 VDD.n287 4.5005
R27752 VDD.n286 VDD.n285 4.5005
R27753 VDD.n281 VDD.n246 4.5005
R27754 VDD.n276 VDD.n275 4.5005
R27755 VDD.n310 VDD.n309 4.5005
R27756 VDD.n312 VDD.n311 4.5005
R27757 VDD.n83 VDD.n82 4.5005
R27758 VDD.n85 VDD.n84 4.5005
R27759 VDD.n8 VDD.n7 4.5005
R27760 VDD.n6 VDD.n5 4.5005
R27761 VDD.n3147 VDD.n3143 4.47034
R27762 VDD.n4141 VDD.n3720 4.46761
R27763 VDD.n4267 VDD.n4266 4.46761
R27764 VDD.n4461 VDD.n4460 4.44348
R27765 VDD.n2185 VDD.n2184 4.44348
R27766 VDD.n2098 VDD.n2094 4.44348
R27767 VDD.n4245 VDD.n4244 4.41955
R27768 VDD.n4131 VDD.n4130 4.41955
R27769 VDD.n3930 VDD.n3928 4.37878
R27770 VDD.n4220 VDD.n4192 4.36875
R27771 VDD.n4218 VDD.n4217 4.36875
R27772 VDD.n4196 VDD.n4194 4.36875
R27773 VDD.n4132 VDD.n3723 4.36875
R27774 VDD.n4072 VDD.n4071 4.36875
R27775 VDD.n4076 VDD.n4073 4.36875
R27776 VDD.n4357 VDD.n4310 4.36875
R27777 VDD.n4315 VDD.n4313 4.36875
R27778 VDD.n4253 VDD.n3694 4.36875
R27779 VDD.n4262 VDD.n4261 4.36875
R27780 VDD.n4065 VDD.n4064 4.36875
R27781 VDD.n3970 VDD.n3969 4.36875
R27782 VDD.n3957 VDD.n3802 4.36875
R27783 VDD.n3408 VDD.n3407 4.36875
R27784 VDD.n3247 VDD.n3245 4.36875
R27785 VDD.n3136 VDD.n3037 4.36875
R27786 VDD.n3195 VDD.n3194 4.36875
R27787 VDD.n2847 VDD.n2846 4.36875
R27788 VDD.n2822 VDD.n2821 4.36875
R27789 VDD.n2792 VDD.n2791 4.36875
R27790 VDD.n2729 VDD.n2728 4.36875
R27791 VDD.n2656 VDD.n2655 4.36875
R27792 VDD.n2550 VDD.n2378 4.36875
R27793 VDD.n2158 VDD.n2157 4.36875
R27794 VDD.n2036 VDD.n2035 4.36875
R27795 VDD.n1966 VDD.n1443 4.36875
R27796 VDD.n1922 VDD.n1466 4.36875
R27797 VDD.n1932 VDD.n1931 4.36875
R27798 VDD.n1855 VDD.n1854 4.36875
R27799 VDD.n1240 VDD.n1239 4.36875
R27800 VDD.n583 VDD.n582 4.36875
R27801 VDD.n1161 VDD.n623 4.36875
R27802 VDD.n1147 VDD.n642 4.36875
R27803 VDD.n1132 VDD.n1131 4.36875
R27804 VDD.n1134 VDD.n1133 4.36875
R27805 VDD.n1107 VDD.n669 4.36875
R27806 VDD.n1113 VDD.n1112 4.36875
R27807 VDD.n1059 VDD.n1058 4.36875
R27808 VDD.n1018 VDD.n1015 4.36875
R27809 VDD.n1024 VDD.n1023 4.36875
R27810 VDD.n994 VDD.n721 4.36875
R27811 VDD.n1002 VDD.n719 4.36875
R27812 VDD.n919 VDD.n918 4.36875
R27813 VDD.n819 VDD.n818 4.36875
R27814 VDD.n523 VDD.n522 4.36875
R27815 VDD.n1160 VDD.n1159 4.31796
R27816 VDD.n809 VDD.n801 4.31796
R27817 VDD.n4231 VDD.n4230 4.26717
R27818 VDD.n3147 VDD.n3146 4.26717
R27819 VDD.n2647 VDD.n2307 4.26717
R27820 VDD.n1345 VDD.n1344 4.26717
R27821 VDD.n973 VDD.n972 4.26717
R27822 VDD.n2503 VDD.n2394 4.2319
R27823 VDD.n4081 VDD.n4080 4.16558
R27824 VDD.n2565 VDD.n2564 4.16558
R27825 VDD.n3226 VDD.n3225 4.14168
R27826 VDD.n2754 VDD.n2753 4.14168
R27827 VDD.n2691 VDD.n2291 4.14168
R27828 VDD.n1886 VDD.n1487 4.14168
R27829 VDD.n1884 VDD.n1883 4.14168
R27830 VDD.n882 VDD.n768 4.14168
R27831 VDD.n860 VDD.n851 4.14168
R27832 VDD.n4449 VDD.n3669 4.12612
R27833 VDD.n2886 VDD.n2093 4.12612
R27834 VDD.n2873 VDD.n2872 4.12612
R27835 VDD.n4233 VDD.n4186 4.11479
R27836 VDD.n1007 VDD.n1005 4.11457
R27837 VDD.n1167 VDD.n1166 4.06399
R27838 VDD.n3741 VDD.n3739 4.02033
R27839 VDD.n3874 VDD.n3830 4.02033
R27840 VDD.n3854 VDD.n3850 4.02033
R27841 VDD.n3854 VDD.n3853 4.02033
R27842 VDD.n3677 VDD.n3675 4.02033
R27843 VDD.n4396 VDD.n4392 4.02033
R27844 VDD.n4396 VDD.n4395 4.02033
R27845 VDD.n3500 VDD.n2924 4.02033
R27846 VDD.n3054 VDD.n3050 4.02033
R27847 VDD.n3054 VDD.n3053 4.02033
R27848 VDD.n3045 VDD.n3042 4.02033
R27849 VDD.n3130 VDD.n3070 4.02033
R27850 VDD.n3605 VDD.n3601 4.02033
R27851 VDD.n3605 VDD.n3604 4.02033
R27852 VDD.n2230 VDD.n2229 4.02033
R27853 VDD.n2583 VDD.n2358 4.02033
R27854 VDD.n2480 VDD.n2476 4.02033
R27855 VDD.n2480 VDD.n2479 4.02033
R27856 VDD.n2133 VDD.n2129 4.02033
R27857 VDD.n2133 VDD.n2132 4.02033
R27858 VDD.n1455 VDD.n1454 4.02033
R27859 VDD.n1749 VDD.n1748 4.02033
R27860 VDD.n1606 VDD.n1605 4.02033
R27861 VDD.n1662 VDD.n1658 4.02033
R27862 VDD.n1662 VDD.n1661 4.02033
R27863 VDD.n1299 VDD.n1295 4.02033
R27864 VDD.n1299 VDD.n1298 4.02033
R27865 VDD.n1223 VDD.n593 4.02033
R27866 VDD.n1142 VDD.n650 4.02033
R27867 VDD.n774 VDD.n773 4.02033
R27868 VDD.n858 VDD.n854 4.02033
R27869 VDD.n858 VDD.n857 4.02033
R27870 VDD.n462 VDD.n459 4.02033
R27871 VDD.n459 VDD.n458 4.02033
R27872 VDD.n489 VDD.n485 4.02033
R27873 VDD.n489 VDD.n488 4.02033
R27874 VDD.n1966 VDD.n1965 4.0132
R27875 VDD.n1017 VDD.n714 4.0132
R27876 VDD.n2708 VDD.n2707 3.91161
R27877 VDD.n2164 VDD.n2104 3.90957
R27878 VDD.n1026 VDD.n1025 3.86515
R27879 VDD.n1847 VDD.n1845 3.8558
R27880 VDD.n2646 VDD.n2307 3.8405
R27881 VDD.n1345 VDD.n1343 3.8405
R27882 VDD.n2500 VDD.n2499 3.78037
R27883 VDD.n4398 VDD.n4389 3.76521
R27884 VDD.n3388 VDD.n3387 3.76521
R27885 VDD.n3330 VDD.n3329 3.76521
R27886 VDD.n3324 VDD.n3323 3.76521
R27887 VDD.n3537 VDD.n3534 3.76521
R27888 VDD.n3538 VDD.n2899 3.76521
R27889 VDD.n3161 VDD.n3160 3.76521
R27890 VDD.n3170 VDD.n3169 3.76521
R27891 VDD.n3170 VDD.n3027 3.76521
R27892 VDD.n3181 VDD.n3179 3.76521
R27893 VDD.n2800 VDD.n2799 3.76521
R27894 VDD.n2765 VDD.n2258 3.76521
R27895 VDD.n1834 VDD.n1833 3.76521
R27896 VDD.n1715 VDD.n1713 3.76521
R27897 VDD.n1718 VDD.n1716 3.76521
R27898 VDD.n1077 VDD.n1076 3.76521
R27899 VDD.n491 VDD.n482 3.76521
R27900 VDD.n56 VDD.n55 3.76521
R27901 VDD.n16 VDD.n15 3.76521
R27902 VDD.n2556 VDD.n2370 3.76495
R27903 VDD.n2499 VDD.n2396 3.69446
R27904 VDD.n433 VDD.n432 3.6805
R27905 VDD.n1680 VDD.n1574 3.66983
R27906 VDD.n463 VDD.n461 3.65009
R27907 VDD.n457 VDD.n454 3.65009
R27908 VDD.n52 VDD.n51 3.63311
R27909 VDD.n23 VDD.n13 3.63295
R27910 VDD.n320 VDD.n182 3.62795
R27911 VDD.t434 VDD.n320 3.62795
R27912 VDD.n232 VDD.n220 3.62795
R27913 VDD.t434 VDD.n220 3.62795
R27914 VDD.n992 VDD.n991 3.61789
R27915 VDD.n910 VDD.n909 3.61789
R27916 VDD.n2838 VDD.n2837 3.59719
R27917 VDD.n3795 VDD.n3793 3.56582
R27918 VDD.n3797 VDD.n3796 3.54093
R27919 VDD.n2164 VDD.n2101 3.52514
R27920 VDD.n2699 VDD.n2698 3.50992
R27921 VDD.n2035 VDD.n1413 3.50526
R27922 VDD.n1240 VDD.n449 3.50526
R27923 VDD.n1147 VDD.n1146 3.50526
R27924 VDD.n4372 VDD.n4370 3.49141
R27925 VDD.n910 VDD.n908 3.47876
R27926 VDD.n3884 VDD.n3823 3.47425
R27927 VDD.n4033 VDD.n3762 3.47425
R27928 VDD.n4037 VDD.n3762 3.47425
R27929 VDD.n4038 VDD.n4037 3.47425
R27930 VDD.n3925 VDD.n3812 3.47425
R27931 VDD.n2601 VDD.n2600 3.47425
R27932 VDD.n2605 VDD.n2604 3.47425
R27933 VDD.n2450 VDD.n2449 3.47425
R27934 VDD.n2446 VDD.n2445 3.47425
R27935 VDD.n2445 VDD.n2444 3.47425
R27936 VDD.n1620 VDD.n1619 3.47425
R27937 VDD.n1619 VDD.n1618 3.47425
R27938 VDD.n1618 VDD.n1588 3.47425
R27939 VDD.n1336 VDD.n1335 3.47425
R27940 VDD.n1335 VDD.n1276 3.47425
R27941 VDD.n4456 VDD.n0 3.43925
R27942 VDD.n4466 VDD.n4465 3.43925
R27943 VDD.n2907 VDD.n1 3.43925
R27944 VDD.n3657 VDD.n3656 3.43925
R27945 VDD.n2882 VDD.n2 3.43925
R27946 VDD.n2891 VDD.n2890 3.43925
R27947 VDD.n2076 VDD.n3 3.43925
R27948 VDD.n2086 VDD.n2085 3.43925
R27949 VDD.n1246 VDD.n4 3.43925
R27950 VDD.n1256 VDD.n1255 3.43925
R27951 VDD.n3661 VDD.n3659 3.4105
R27952 VDD.n4454 VDD.n4453 3.4105
R27953 VDD.n2895 VDD.n2893 3.4105
R27954 VDD.n2904 VDD.n2903 3.4105
R27955 VDD.n2090 VDD.n2088 3.4105
R27956 VDD.n2880 VDD.n2879 3.4105
R27957 VDD.n1260 VDD.n1258 3.4105
R27958 VDD.n2074 VDD.n2073 3.4105
R27959 VDD.n441 VDD.n439 3.4105
R27960 VDD.n1244 VDD.n1243 3.4105
R27961 VDD.n4103 VDD.n3735 3.38874
R27962 VDD.n3323 VDD.n2976 3.38874
R27963 VDD.n3540 VDD.n3537 3.38874
R27964 VDD.n2686 VDD.n2685 3.38874
R27965 VDD.n1997 VDD.n1996 3.38874
R27966 VDD.n1487 VDD.n1484 3.38874
R27967 VDD.n893 VDD.n892 3.38874
R27968 VDD.n94 VDD.n93 3.38874
R27969 VDD.n4279 VDD.n4278 3.37141
R27970 VDD.n4061 VDD.n4060 3.36242
R27971 VDD.n2600 VDD.n2599 3.36097
R27972 VDD.t1296 VDD.t2625 3.35739
R27973 VDD.t1187 VDD.t2323 3.35739
R27974 VDD.t288 VDD.t575 3.35739
R27975 VDD.t3088 VDD.t1218 3.35739
R27976 VDD.n3296 VDD.t1585 3.35739
R27977 VDD.t131 VDD.t2219 3.35739
R27978 VDD.t980 VDD.t189 3.35739
R27979 VDD.t272 VDD.t1251 3.35739
R27980 VDD.t497 VDD.t503 3.35739
R27981 VDD.t1675 VDD.t2912 3.35739
R27982 VDD.t2085 VDD.t1832 3.35739
R27983 VDD.t748 VDD.t1869 3.35739
R27984 VDD.t746 VDD.t1867 3.35739
R27985 VDD.t2491 VDD.t2824 3.35739
R27986 VDD.t2314 VDD.t533 3.35739
R27987 VDD.t657 VDD.t2714 3.35739
R27988 VDD.t659 VDD.t2716 3.35739
R27989 VDD.t2813 VDD.t1614 3.35739
R27990 VDD.t1790 VDD.t946 3.35739
R27991 VDD.t2261 VDD.t3085 3.35739
R27992 VDD.t0 VDD.t2145 3.35739
R27993 VDD.t2032 VDD.t2529 3.35739
R27994 VDD.t2607 VDD.t484 3.35739
R27995 VDD.t897 VDD.t540 3.35739
R27996 VDD.n3928 VDD.n3927 3.30778
R27997 VDD.n1346 VDD.n1345 3.29837
R27998 VDD.n1123 VDD.n1122 3.29403
R27999 VDD.n4399 VDD.n4396 3.28705
R28000 VDD.n861 VDD.n858 3.28705
R28001 VDD.n492 VDD.n489 3.28705
R28002 VDD.n3792 VDD.n3790 3.25799
R28003 VDD.n2841 VDD.n2840 3.25799
R28004 VDD.n629 VDD.n627 3.25799
R28005 VDD.n3879 VDD.n3823 3.2477
R28006 VDD.n3885 VDD.n3884 3.2477
R28007 VDD.n4029 VDD.n3764 3.2477
R28008 VDD.n4039 VDD.n4038 3.2477
R28009 VDD.n3920 VDD.n3812 3.2477
R28010 VDD.n3926 VDD.n3925 3.2477
R28011 VDD.n2339 VDD.n2336 3.2477
R28012 VDD.n2606 VDD.n2605 3.2477
R28013 VDD.n2452 VDD.n2407 3.2477
R28014 VDD.n2444 VDD.n2411 3.2477
R28015 VDD.n1626 VDD.n1625 3.2477
R28016 VDD.n1590 VDD.n1588 3.2477
R28017 VDD.n1331 VDD.n1330 3.2477
R28018 VDD.n3970 VDD.n3968 3.2005
R28019 VDD.n2106 VDD.n2105 3.2005
R28020 VDD.n2160 VDD.n2114 3.2005
R28021 VDD.n666 VDD.n665 3.2005
R28022 VDD.n1124 VDD.n1123 3.2005
R28023 VDD.n524 VDD.n463 3.2005
R28024 VDD.n431 VDD.n430 3.18667
R28025 VDD.n1928 VDD.n1464 3.14971
R28026 VDD.n3694 VDD.n3693 3.12116
R28027 VDD.n4064 VDD.n4063 3.12116
R28028 VDD.n798 VDD.n797 3.12116
R28029 VDD.n4020 VDD.n4019 3.09891
R28030 VDD.n3946 VDD.n3807 3.06827
R28031 VDD.n177 VDD.n176 3.04961
R28032 VDD.n3874 VDD.n3827 3.04861
R28033 VDD.n4096 VDD.n3741 3.04861
R28034 VDD.n4307 VDD.n3677 3.04861
R28035 VDD.n3063 VDD.n3045 3.04861
R28036 VDD.n3130 VDD.n3067 3.04861
R28037 VDD.n3500 VDD.n2925 3.04861
R28038 VDD.n2583 VDD.n2355 3.04861
R28039 VDD.n1749 VDD.n1549 3.04861
R28040 VDD.n1946 VDD.n1455 3.04861
R28041 VDD.n802 VDD.n774 3.04861
R28042 VDD.n1142 VDD.n647 3.04861
R28043 VDD.n1223 VDD.n590 3.04861
R28044 VDD.n2834 VDD.n2230 3.04861
R28045 VDD.n2164 VDD.n2163 3.04861
R28046 VDD.n526 VDD.n459 3.04861
R28047 VDD.n3894 VDD.n3893 3.01588
R28048 VDD.n4284 VDD.n3683 3.01588
R28049 VDD.n3123 VDD.n3073 3.01588
R28050 VDD.n3120 VDD.n3119 3.01588
R28051 VDD.n3100 VDD.n3099 3.01588
R28052 VDD.n3098 VDD.n3081 3.01588
R28053 VDD.n3631 VDD.n3585 3.01588
R28054 VDD.n2426 VDD.n2425 3.01588
R28055 VDD.n2028 VDD.n1417 3.01226
R28056 VDD.n544 VDD.n541 3.01226
R28057 VDD.n577 VDD.n576 3.01226
R28058 VDD.n897 VDD.n755 3.01226
R28059 VDD.n4245 VDD.n4183 2.99733
R28060 VDD.n2559 VDD.n2558 2.99733
R28061 VDD.n4164 VDD.n4163 2.98664
R28062 VDD.n4138 VDD.n3722 2.96248
R28063 VDD.n4271 VDD.n4270 2.96248
R28064 VDD.n1058 VDD.n1057 2.94653
R28065 VDD.n3793 VDD.n3792 2.91308
R28066 VDD.n3637 VDD.n3579 2.91308
R28067 VDD.n3637 VDD.n3582 2.91308
R28068 VDD.n2840 VDD.n2839 2.91308
R28069 VDD.n630 VDD.n629 2.91308
R28070 VDD.n633 VDD.n630 2.91308
R28071 VDD.n4357 VDD.n4356 2.89574
R28072 VDD.n4182 VDD.n3700 2.87861
R28073 VDD.n3876 VDD.n3875 2.87861
R28074 VDD.n3917 VDD.n3916 2.87861
R28075 VDD.n2557 VDD.n2556 2.87861
R28076 VDD.n173 VDD.t152 2.857
R28077 VDD.n173 VDD.t149 2.857
R28078 VDD.n172 VDD.t147 2.857
R28079 VDD.t152 VDD.n172 2.857
R28080 VDD.t2937 VDD.n153 2.857
R28081 VDD.n153 VDD.t2939 2.857
R28082 VDD.t2938 VDD.n154 2.857
R28083 VDD.n154 VDD.t2937 2.857
R28084 VDD.n4240 VDD.n4185 2.8165
R28085 VDD.n1683 VDD.n1681 2.8165
R28086 VDD.n661 VDD.n658 2.8165
R28087 VDD.n327 VDD.n181 2.76312
R28088 VDD.n4062 VDD.n4061 2.75091
R28089 VDD.n2372 VDD.n2371 2.75091
R28090 VDD.n4163 VDD.n4162 2.70664
R28091 VDD.n2451 VDD.n2406 2.6965
R28092 VDD.n70 VDD.n66 2.66717
R28093 VDD.n33 VDD.n30 2.66717
R28094 VDD.n3893 VDD.n3819 2.64665
R28095 VDD.n4287 VDD.n3683 2.64665
R28096 VDD.n3120 VDD.n3073 2.64665
R28097 VDD.n3119 VDD.n3118 2.64665
R28098 VDD.n3099 VDD.n3098 2.64665
R28099 VDD.n3095 VDD.n3081 2.64665
R28100 VDD.n3628 VDD.n3585 2.64665
R28101 VDD.n2425 VDD.n2424 2.64665
R28102 VDD.n4063 VDD.n4061 2.64513
R28103 VDD.n2371 VDD.n2370 2.64513
R28104 VDD.n634 VDD.n632 2.64481
R28105 VDD.n1176 VDD.n619 2.64177
R28106 VDD.n930 VDD.n742 2.64177
R28107 VDD.n4403 VDD.n4402 2.63579
R28108 VDD.n2710 VDD.n2282 2.63579
R28109 VDD.n2630 VDD.n2319 2.63579
R28110 VDD.n1384 VDD.n1383 2.63579
R28111 VDD.n2002 VDD.n2001 2.63579
R28112 VDD.n1874 VDD.n1873 2.63579
R28113 VDD.n1744 VDD.n1743 2.63579
R28114 VDD.n554 VDD.n552 2.63579
R28115 VDD.n1033 VDD.n1032 2.63579
R28116 VDD.n942 VDD.n740 2.63579
R28117 VDD.n865 VDD.n864 2.63579
R28118 VDD.n496 VDD.n495 2.63579
R28119 VDD.n421 VDD.n420 2.63579
R28120 VDD.n3693 VDD.n3691 2.63539
R28121 VDD.n3739 VDD.n3737 2.63539
R28122 VDD.n3830 VDD.n3828 2.63539
R28123 VDD.n3850 VDD.n3848 2.63539
R28124 VDD.n3853 VDD.n3851 2.63539
R28125 VDD.n3675 VDD.n3673 2.63539
R28126 VDD.n4392 VDD.n4390 2.63539
R28127 VDD.n4395 VDD.n4393 2.63539
R28128 VDD.n2924 VDD.n2922 2.63539
R28129 VDD.n3050 VDD.n3048 2.63539
R28130 VDD.n3053 VDD.n3051 2.63539
R28131 VDD.n3042 VDD.n3040 2.63539
R28132 VDD.n3070 VDD.n3068 2.63539
R28133 VDD.n3601 VDD.n3599 2.63539
R28134 VDD.n3604 VDD.n3602 2.63539
R28135 VDD.n2229 VDD.n2227 2.63539
R28136 VDD.n2358 VDD.n2356 2.63539
R28137 VDD.n2476 VDD.n2474 2.63539
R28138 VDD.n2479 VDD.n2477 2.63539
R28139 VDD.n2104 VDD.n2102 2.63539
R28140 VDD.n2129 VDD.n2127 2.63539
R28141 VDD.n2132 VDD.n2130 2.63539
R28142 VDD.n1454 VDD.n1452 2.63539
R28143 VDD.n1748 VDD.n1746 2.63539
R28144 VDD.n1658 VDD.n1656 2.63539
R28145 VDD.n1661 VDD.n1659 2.63539
R28146 VDD.n1295 VDD.n1293 2.63539
R28147 VDD.n1298 VDD.n1296 2.63539
R28148 VDD.n797 VDD.n795 2.63539
R28149 VDD.n593 VDD.n591 2.63539
R28150 VDD.n650 VDD.n648 2.63539
R28151 VDD.n773 VDD.n771 2.63539
R28152 VDD.n854 VDD.n852 2.63539
R28153 VDD.n857 VDD.n855 2.63539
R28154 VDD.n485 VDD.n483 2.63539
R28155 VDD.n488 VDD.n486 2.63539
R28156 VDD.n3880 VDD.n3878 2.63233
R28157 VDD.n3921 VDD.n3919 2.63233
R28158 VDD.n4183 VDD.n4181 2.61352
R28159 VDD.n3878 VDD.n3877 2.61352
R28160 VDD.n3919 VDD.n3918 2.61352
R28161 VDD.n2558 VDD.n2369 2.61352
R28162 VDD.n177 VDD.n87 2.61002
R28163 VDD.n1173 VDD.n1172 2.54018
R28164 VDD.n1001 VDD.n1000 2.54018
R28165 VDD.n1932 VDD.n1930 2.48939
R28166 VDD.n425 VDD.n413 2.48504
R28167 VDD.n1923 VDD.n1922 2.4386
R28168 VDD.n818 VDD.n817 2.4386
R28169 VDD.n4141 VDD.n4140 2.40784
R28170 VDD.n4268 VDD.n4267 2.40784
R28171 VDD.n3692 VDD.n3691 2.37495
R28172 VDD.n3738 VDD.n3737 2.37495
R28173 VDD.n3829 VDD.n3828 2.37495
R28174 VDD.n3852 VDD.n3851 2.37495
R28175 VDD.n3849 VDD.n3848 2.37495
R28176 VDD.n3674 VDD.n3673 2.37495
R28177 VDD.n4394 VDD.n4393 2.37495
R28178 VDD.n4391 VDD.n4390 2.37495
R28179 VDD.n2923 VDD.n2922 2.37495
R28180 VDD.n3052 VDD.n3051 2.37495
R28181 VDD.n3049 VDD.n3048 2.37495
R28182 VDD.n3041 VDD.n3040 2.37495
R28183 VDD.n3069 VDD.n3068 2.37495
R28184 VDD.n3603 VDD.n3602 2.37495
R28185 VDD.n3600 VDD.n3599 2.37495
R28186 VDD.n2228 VDD.n2227 2.37495
R28187 VDD.n2357 VDD.n2356 2.37495
R28188 VDD.n2478 VDD.n2477 2.37495
R28189 VDD.n2475 VDD.n2474 2.37495
R28190 VDD.n2103 VDD.n2102 2.37495
R28191 VDD.n2131 VDD.n2130 2.37495
R28192 VDD.n2128 VDD.n2127 2.37495
R28193 VDD.n1453 VDD.n1452 2.37495
R28194 VDD.n1747 VDD.n1746 2.37495
R28195 VDD.n1660 VDD.n1659 2.37495
R28196 VDD.n1657 VDD.n1656 2.37495
R28197 VDD.n1297 VDD.n1296 2.37495
R28198 VDD.n1294 VDD.n1293 2.37495
R28199 VDD.n796 VDD.n795 2.37495
R28200 VDD.n592 VDD.n591 2.37495
R28201 VDD.n649 VDD.n648 2.37495
R28202 VDD.n772 VDD.n771 2.37495
R28203 VDD.n856 VDD.n855 2.37495
R28204 VDD.n853 VDD.n852 2.37495
R28205 VDD.n487 VDD.n486 2.37495
R28206 VDD.n484 VDD.n483 2.37495
R28207 VDD.n990 VDD.n988 2.34574
R28208 VDD.n4237 VDD.n4185 2.33701
R28209 VDD.n4130 VDD.n4129 2.33701
R28210 VDD.n4017 VDD.n4016 2.33701
R28211 VDD.n4059 VDD.n3755 2.33701
R28212 VDD.n3409 VDD.n3353 2.33701
R28213 VDD.n3254 VDD.n3253 2.33701
R28214 VDD.n3188 VDD.n3019 2.33701
R28215 VDD.n2815 VDD.n2235 2.33701
R28216 VDD.n2789 VDD.n2248 2.33701
R28217 VDD.n2722 VDD.n2274 2.33701
R28218 VDD.n2700 VDD.n2285 2.33701
R28219 VDD.n2697 VDD.n2288 2.33701
R28220 VDD.n2649 VDD.n2648 2.33701
R28221 VDD.n2549 VDD.n2548 2.33701
R28222 VDD.n2066 VDD.n2065 2.33701
R28223 VDD.n2064 VDD.n1268 2.33701
R28224 VDD.n1964 VDD.n1963 2.33701
R28225 VDD.n1848 VDD.n1506 2.33701
R28226 VDD.n584 VDD.n533 2.33701
R28227 VDD.n658 VDD.n657 2.33701
R28228 VDD.n1056 VDD.n698 2.33701
R28229 VDD.n970 VDD.n969 2.33701
R28230 VDD.n953 VDD.n952 2.33701
R28231 VDD.n913 VDD.n912 2.33701
R28232 VDD.n2837 VDD.n2230 2.32777
R28233 VDD.n68 VDD.n66 2.313
R28234 VDD.n74 VDD.n68 2.313
R28235 VDD.n32 VDD.n30 2.313
R28236 VDD.n37 VDD.n32 2.313
R28237 VDD.n637 VDD.n632 2.29615
R28238 VDD.n69 VDD.n67 2.28445
R28239 VDD.n73 VDD.n67 2.28445
R28240 VDD.n31 VDD.n29 2.28445
R28241 VDD.n36 VDD.n31 2.28445
R28242 VDD.n160 VDD.n159 2.28415
R28243 VDD.n2110 VDD.n2109 2.28407
R28244 VDD.n2112 VDD.n2110 2.28407
R28245 VDD.n1273 VDD.n1271 2.28374
R28246 VDD.n4111 VDD.n4110 2.25932
R28247 VDD.n3449 VDD.n3448 2.25932
R28248 VDD.n2540 VDD.n2539 2.25932
R28249 VDD.n1895 VDD.n1894 2.25932
R28250 VDD.n1040 VDD.n1039 2.25932
R28251 VDD.n3916 VDD.n3813 2.25312
R28252 VDD.n3964 VDD.n3793 2.25312
R28253 VDD.n2839 VDD.n2225 2.25312
R28254 VDD.n1156 VDD.n630 2.25312
R28255 VDD.n3875 VDD.n3824 2.25293
R28256 VDD.n4247 VDD.n3700 2.25293
R28257 VDD.n3637 VDD.n3576 2.25293
R28258 VDD.n1924 VDD.n1923 2.23542
R28259 VDD.n817 VDD.n816 2.23542
R28260 VDD.n381 VDD.t1729 2.2191
R28261 VDD.n1930 VDD.n1929 2.18463
R28262 VDD.n957 VDD.n956 2.18463
R28263 VDD.n956 VDD.n955 2.18463
R28264 VDD.n1684 VDD.n1683 2.1843
R28265 VDD.n3796 VDD.n3795 2.13621
R28266 VDD.n1174 VDD.n1173 2.13383
R28267 VDD.n1002 VDD.n1001 2.13383
R28268 VDD.n928 VDD.n927 2.13383
R28269 VDD.n2108 VDD.n2105 2.07374
R28270 VDD.n2114 VDD.n2113 2.07374
R28271 VDD.n911 VDD.n910 2.06227
R28272 VDD.n25 VDD.n13 2.05049
R28273 VDD.n51 VDD.n46 2.05017
R28274 VDD.n4129 VDD.n4128 2.03225
R28275 VDD.n4016 VDD.n4015 2.03225
R28276 VDD.n4055 VDD.n3755 2.03225
R28277 VDD.n3353 VDD.n3352 2.03225
R28278 VDD.n3255 VDD.n3254 2.03225
R28279 VDD.n3189 VDD.n3188 2.03225
R28280 VDD.n2816 VDD.n2815 2.03225
R28281 VDD.n2784 VDD.n2248 2.03225
R28282 VDD.n2723 VDD.n2722 2.03225
R28283 VDD.n2701 VDD.n2700 2.03225
R28284 VDD.n2693 VDD.n2288 2.03225
R28285 VDD.n2648 VDD.n2306 2.03225
R28286 VDD.n2548 VDD.n2547 2.03225
R28287 VDD.n2067 VDD.n2066 2.03225
R28288 VDD.n1270 VDD.n1268 2.03225
R28289 VDD.n1963 VDD.n1962 2.03225
R28290 VDD.n1849 VDD.n1848 2.03225
R28291 VDD.n533 VDD.n532 2.03225
R28292 VDD.n1052 VDD.n698 2.03225
R28293 VDD.n969 VDD.n968 2.03225
R28294 VDD.n926 VDD.n925 2.03225
R28295 VDD.n912 VDD.n749 2.03225
R28296 VDD.n3579 VDD.n3577 2.01703
R28297 VDD.n3582 VDD.n3580 2.01703
R28298 VDD.n141 VDD.n109 2.01137
R28299 VDD.t151 VDD.n109 2.01137
R28300 VDD.n148 VDD.n147 2.01137
R28301 VDD.n147 VDD.t151 2.01137
R28302 VDD.n146 VDD.n145 2.01137
R28303 VDD.t151 VDD.n146 2.01137
R28304 VDD.n3982 VDD.n3782 2.0005
R28305 VDD.n4140 VDD.n4139 1.99683
R28306 VDD.n4269 VDD.n4268 1.99683
R28307 VDD.n143 VDD.n142 1.9205
R28308 VDD.n3581 VDD.n3580 1.88416
R28309 VDD.n3578 VDD.n3577 1.88416
R28310 VDD.n4117 VDD.n4116 1.88285
R28311 VDD.n2716 VDD.n2715 1.88285
R28312 VDD.n2636 VDD.n2635 1.88285
R28313 VDD.n2622 VDD.n2621 1.88285
R28314 VDD.n1378 VDD.n1377 1.88285
R28315 VDD.n2050 VDD.n2049 1.88285
R28316 VDD.n2010 VDD.n2009 1.88285
R28317 VDD.n1956 VDD.n1955 1.88285
R28318 VDD.n1917 VDD.n1916 1.88285
R28319 VDD.n1828 VDD.n1827 1.88285
R28320 VDD.n2434 VDD.n2433 1.88273
R28321 VDD.n13 VDD.n12 1.87577
R28322 VDD.n51 VDD.n50 1.87546
R28323 VDD.n4032 VDD.n4031 1.85065
R28324 VDD.n2601 VDD.n2334 1.85065
R28325 VDD.n2452 VDD.n2451 1.85065
R28326 VDD.n2449 VDD.n2409 1.85065
R28327 VDD.n1623 VDD.n1586 1.85065
R28328 VDD.n1278 VDD.n1276 1.85065
R28329 VDD.n4030 VDD.n4029 1.81289
R28330 VDD.n1625 VDD.n1624 1.81289
R28331 VDD.n3086 VDD.n3039 1.78512
R28332 VDD.n4356 VDD.n4355 1.77828
R28333 VDD.n2556 VDD.n2368 1.76897
R28334 VDD.n2162 VDD.n2110 1.76897
R28335 VDD.n463 VDD.n462 1.74595
R28336 VDD.n458 VDD.n454 1.74595
R28337 VDD.n1177 VDD.n1176 1.72748
R28338 VDD.n1057 VDD.n1056 1.72748
R28339 VDD.n931 VDD.n930 1.72748
R28340 VDD.n1257 VDD.n4 1.69188
R28341 VDD.n1257 VDD.n1256 1.69188
R28342 VDD.n2087 VDD.n3 1.69188
R28343 VDD.n2087 VDD.n2086 1.69188
R28344 VDD.n2892 VDD.n2 1.69188
R28345 VDD.n2892 VDD.n2891 1.69188
R28346 VDD.n3658 VDD.n1 1.69188
R28347 VDD.n3658 VDD.n3657 1.69188
R28348 VDD.n4467 VDD.n0 1.69188
R28349 VDD.n4467 VDD.n4466 1.69188
R28350 VDD.n2839 VDD.n2838 1.68673
R28351 VDD.n3855 VDD.n3854 1.6819
R28352 VDD.n3606 VDD.n3605 1.6819
R28353 VDD.n2481 VDD.n2480 1.6819
R28354 VDD.n2134 VDD.n2133 1.6819
R28355 VDD.n1663 VDD.n1662 1.6819
R28356 VDD.n1300 VDD.n1299 1.6819
R28357 VDD.n3055 VDD.n3054 1.68181
R28358 VDD.t1687 VDD.t3081 1.67895
R28359 VDD.t1765 VDD.t3059 1.67895
R28360 VDD.t2376 VDD.t2752 1.67895
R28361 VDD.t1957 VDD.t2043 1.67895
R28362 VDD.t1308 VDD.t3061 1.67895
R28363 VDD.t2942 VDD.t2680 1.67895
R28364 VDD.t383 VDD.t2151 1.67895
R28365 VDD.t381 VDD.t2149 1.67895
R28366 VDD.t2093 VDD.t1711 1.67895
R28367 VDD.t1204 VDD.t1837 1.67895
R28368 VDD.n2237 VDD.t2863 1.67895
R28369 VDD.t3072 VDD.t1941 1.67895
R28370 VDD.t3076 VDD.t1943 1.67895
R28371 VDD.t372 VDD.t1457 1.67895
R28372 VDD.t370 VDD.t1455 1.67895
R28373 VDD.t2397 VDD.t135 1.67895
R28374 VDD.t221 VDD.t2667 1.67895
R28375 VDD.t2790 VDD.t933 1.67895
R28376 VDD.t1479 VDD.t1278 1.67895
R28377 VDD.t1475 VDD.t1965 1.67895
R28378 VDD.t209 VDD.t1875 1.67895
R28379 VDD.t925 VDD.t619 1.67895
R28380 VDD.n4031 VDD.n4030 1.66186
R28381 VDD.n1624 VDD.n1623 1.66186
R28382 VDD.n178 VDD.n86 1.6358
R28383 VDD.n4033 VDD.n4032 1.6241
R28384 VDD.n2604 VDD.n2334 1.6241
R28385 VDD.n2451 VDD.n2450 1.6241
R28386 VDD.n2446 VDD.n2409 1.6241
R28387 VDD.n1620 VDD.n1586 1.6241
R28388 VDD.n1338 VDD.n1337 1.6241
R28389 VDD.n1337 VDD.n1336 1.6241
R28390 VDD.n1331 VDD.n1278 1.6241
R28391 VDD.n2433 VDD.n2432 1.62188
R28392 VDD.n81 VDD.n80 1.58787
R28393 VDD.n3888 VDD.n3887 1.5792
R28394 VDD.n2105 VDD.n2101 1.53093
R28395 VDD.n1925 VDD.n1464 1.52431
R28396 VDD.n3460 VDD.n3459 1.50638
R28397 VDD.n3441 VDD.n3440 1.50638
R28398 VDD.n3313 VDD.n3312 1.50638
R28399 VDD.n3553 VDD.n3552 1.50638
R28400 VDD.n2716 VDD.n2279 1.50638
R28401 VDD.n2636 VDD.n2316 1.50638
R28402 VDD.n2487 VDD.n2468 1.50638
R28403 VDD.n1635 VDD.n1582 1.50638
R28404 VDD.n1645 VDD.n1644 1.50638
R28405 VDD.n1393 VDD.n1355 1.50638
R28406 VDD.n2023 VDD.n2022 1.50638
R28407 VDD.n1976 VDD.n1975 1.50638
R28408 VDD.n1789 VDD.n1535 1.50638
R28409 VDD.n1669 VDD.n1650 1.50638
R28410 VDD.n564 VDD.n563 1.50638
R28411 VDD.n80 VDD.n62 1.49911
R28412 VDD.n44 VDD.n26 1.49911
R28413 VDD.n178 VDD.n177 1.49369
R28414 VDD.n4125 VDD.n3725 1.47352
R28415 VDD.n4066 VDD.n3753 1.47352
R28416 VDD.n3968 VDD.n3967 1.47352
R28417 VDD.n2850 VDD.n2849 1.47352
R28418 VDD.n2642 VDD.n2308 1.47352
R28419 VDD.n2061 VDD.n2060 1.47352
R28420 VDD.n1123 VDD.n665 1.47352
R28421 VDD.n907 VDD.n750 1.47352
R28422 VDD.n821 VDD.n792 1.47352
R28423 VDD.n1961 VDD.n1446 1.45766
R28424 VDD.n1014 VDD.n1013 1.45766
R28425 VDD.n328 VDD.n179 1.41175
R28426 VDD.n145 VDD.n139 1.4085
R28427 VDD.n2578 VDD.n2577 1.4005
R28428 VDD.n2534 VDD.n2533 1.4005
R28429 VDD.n1850 VDD.n1847 1.38171
R28430 VDD.n2824 VDD.n2233 1.37571
R28431 VDD.n150 VDD.n88 1.3755
R28432 VDD.n45 VDD.n44 1.37105
R28433 VDD.n3858 VDD.n3855 1.30718
R28434 VDD.n3607 VDD.n3606 1.30718
R28435 VDD.n2482 VDD.n2481 1.30718
R28436 VDD.n2135 VDD.n2134 1.30718
R28437 VDD.n1664 VDD.n1663 1.30718
R28438 VDD.n1301 VDD.n1300 1.30718
R28439 VDD.n3056 VDD.n3055 1.30711
R28440 VDD.n4019 VDD.n3766 1.27034
R28441 VDD.n633 VDD.n632 1.26517
R28442 VDD.n176 VDD.n88 1.2505
R28443 VDD.n4183 VDD.n4182 1.2502
R28444 VDD.n3878 VDD.n3876 1.2502
R28445 VDD.n3919 VDD.n3917 1.2502
R28446 VDD.n2558 VDD.n2557 1.2502
R28447 VDD.n3887 VDD.n3886 1.23724
R28448 VDD.n951 VDD.n950 1.21955
R28449 VDD.n438 VDD.n45 1.21856
R28450 VDD.n437 VDD.n436 1.2116
R28451 VDD.n270 VDD.n269 1.17383
R28452 VDD.n4295 VDD.n4294 1.16414
R28453 VDD.n1607 VDD.n1606 1.16414
R28454 VDD.n2858 VDD.n2218 1.12991
R28455 VDD.n1751 VDD.n1750 1.12991
R28456 VDD.n1781 VDD.n1779 1.12991
R28457 VDD.n149 VDD.n148 1.09764
R28458 VDD.n1627 VDD.n1584 1.09549
R28459 VDD.n2702 VDD.n2699 1.08084
R28460 VDD.n330 VDD.n178 1.07996
R28461 VDD.n437 VDD.n330 1.06614
R28462 VDD.n4158 VDD.n4157 1.05835
R28463 VDD.n4431 VDD.n4372 1.05835
R28464 VDD.n2340 VDD.n2337 1.05773
R28465 VDD.n2456 VDD.n2455 1.05773
R28466 VDD.n1339 VDD.n1273 1.05773
R28467 VDD.n329 VDD.n328 1.03946
R28468 VDD.n1060 VDD.n695 1.01251
R28469 VDD.n3989 VDD.n3988 1.0005
R28470 VDD.n2109 VDD.n2105 0.992049
R28471 VDD.n2114 VDD.n2112 0.992049
R28472 VDD.n995 VDD.n993 0.965579
R28473 VDD.n2612 VDD.n2611 0.952566
R28474 VDD.n2504 VDD.n2503 0.952566
R28475 VDD.n419 VDD.n418 0.944798
R28476 VDD.n170 VDD.n169 0.904346
R28477 VDD.n3984 VDD.n3782 0.9005
R28478 VDD.n3677 VDD.n3676 0.899674
R28479 VDD.n3045 VDD.n3044 0.899674
R28480 VDD.n3130 VDD.n3066 0.899674
R28481 VDD.n1749 VDD.n1745 0.899674
R28482 VDD.n4237 VDD.n4236 0.863992
R28483 VDD.n2031 VDD.n1413 0.863992
R28484 VDD.n449 VDD.n446 0.863992
R28485 VDD.n1146 VDD.n1145 0.863992
R28486 VDD.n1130 VDD.n657 0.863992
R28487 VDD.n952 VDD.n951 0.813198
R28488 VDD.n170 VDD.n161 0.808192
R28489 VDD.n1958 VDD.n1446 0.770079
R28490 VDD.n1013 VDD.n1012 0.770079
R28491 VDD.n155 VDD.n104 0.757118
R28492 VDD.n152 VDD.n104 0.757118
R28493 VDD.n152 VDD.n151 0.757118
R28494 VDD.n171 VDD.n89 0.757118
R28495 VDD.n174 VDD.n89 0.757118
R28496 VDD.n175 VDD.n174 0.757118
R28497 VDD.n4208 VDD.n4207 0.753441
R28498 VDD.n4167 VDD.n3708 0.753441
R28499 VDD.n4087 VDD.n3748 0.753441
R28500 VDD.n4398 VDD.n4397 0.753441
R28501 VDD.n3515 VDD.n3514 0.753441
R28502 VDD.n3474 VDD.n3473 0.753441
R28503 VDD.n3472 VDD.n3471 0.753441
R28504 VDD.n3450 VDD.n3449 0.753441
R28505 VDD.n3426 VDD.n2963 0.753441
R28506 VDD.n3372 VDD.n3369 0.753441
R28507 VDD.n3372 VDD.n3371 0.753441
R28508 VDD.n3379 VDD.n3378 0.753441
R28509 VDD.n3402 VDD.n3401 0.753441
R28510 VDD.n3339 VDD.n3338 0.753441
R28511 VDD.n3315 VDD.n2981 0.753441
R28512 VDD.n3308 VDD.n2984 0.753441
R28513 VDD.n3557 VDD.n3527 0.753441
R28514 VDD.n3550 VDD.n3530 0.753441
R28515 VDD.n3646 VDD.n3645 0.753441
R28516 VDD.n3210 VDD.n3209 0.753441
R28517 VDD.n3155 VDD.n3153 0.753441
R28518 VDD.n3186 VDD.n3185 0.753441
R28519 VDD.n2191 VDD.n2190 0.753441
R28520 VDD.n2782 VDD.n2781 0.753441
R28521 VDD.n2753 VDD.n2752 0.753441
R28522 VDD.n2748 VDD.n2747 0.753441
R28523 VDD.n2487 VDD.n2486 0.753441
R28524 VDD.n1636 VDD.n1635 0.753441
R28525 VDD.n1645 VDD.n1577 0.753441
R28526 VDD.n1818 VDD.n1817 0.753441
R28527 VDD.n1796 VDD.n1795 0.753441
R28528 VDD.n1701 VDD.n1700 0.753441
R28529 VDD.n1757 VDD.n1756 0.753441
R28530 VDD.n1669 VDD.n1668 0.753441
R28531 VDD.n1251 VDD.n1250 0.753441
R28532 VDD.n1197 VDD.n1196 0.753441
R28533 VDD.n1106 VDD.n1105 0.753441
R28534 VDD.n1045 VDD.n703 0.753441
R28535 VDD.n1029 VDD.n712 0.753441
R28536 VDD.n982 VDD.n981 0.753441
R28537 VDD.n936 VDD.n935 0.753441
R28538 VDD.n866 VDD.n865 0.753441
R28539 VDD.n860 VDD.n859 0.753441
R28540 VDD.n491 VDD.n490 0.753441
R28541 VDD.n2616 VDD.n2615 0.740996
R28542 VDD.n2509 VDD.n2508 0.740996
R28543 VDD.n1480 VDD.n1455 0.708966
R28544 VDD.n2574 VDD.n2573 0.7005
R28545 VDD.n2530 VDD.n2529 0.7005
R28546 VDD.n1965 VDD.n1964 0.660817
R28547 VDD.n1018 VDD.n1017 0.660817
R28548 VDD.n3791 VDD.n3790 0.651997
R28549 VDD.n2841 VDD.n2226 0.651997
R28550 VDD.n628 VDD.n627 0.651997
R28551 VDD.n3700 VDD.n3699 0.644287
R28552 VDD.n3916 VDD.n3915 0.644287
R28553 VDD.n77 VDD.n76 0.6405
R28554 VDD.n40 VDD.n39 0.6405
R28555 VDD.n3722 VDD.n3721 0.635211
R28556 VDD.n4149 VDD.n4148 0.635211
R28557 VDD.n4162 VDD.n3712 0.635211
R28558 VDD.n4323 VDD.n4321 0.635211
R28559 VDD.n4272 VDD.n4271 0.635211
R28560 VDD.n4302 VDD.n3679 0.635211
R28561 VDD.n4025 VDD.n4024 0.635211
R28562 VDD.n4046 VDD.n4045 0.635211
R28563 VDD.n3930 VDD.n3929 0.635211
R28564 VDD.n4368 VDD.n4365 0.635211
R28565 VDD.n4420 VDD.n4376 0.635211
R28566 VDD.n3129 VDD.n3071 0.635211
R28567 VDD.n2189 VDD.n2177 0.635211
R28568 VDD.n2869 VDD.n2099 0.635211
R28569 VDD.n2825 VDD.n2824 0.635211
R28570 VDD.n2661 VDD.n2660 0.635211
R28571 VDD.n2681 VDD.n2680 0.635211
R28572 VDD.n2619 VDD.n2329 0.635211
R28573 VDD.n2521 VDD.n2520 0.635211
R28574 VDD.n1599 VDD.n1598 0.635211
R28575 VDD.n318 VDD.n317 0.622722
R28576 VDD.n43 VDD.n27 0.600153
R28577 VDD.n79 VDD.n78 0.599785
R28578 VDD.n156 VDD.n155 0.590759
R28579 VDD.n96 VDD.n95 0.589728
R28580 VDD.n167 VDD.n164 0.588815
R28581 VDD.n4420 VDD.n4419 0.581389
R28582 VDD.n4236 VDD.n4186 0.55923
R28583 VDD.n3909 VDD.n3908 0.529426
R28584 VDD.n2515 VDD.n2514 0.529426
R28585 VDD.n316 VDD.n315 0.519731
R28586 VDD.n993 VDD.n987 0.508436
R28587 VDD.n3985 VDD.n3984 0.5005
R28588 VDD.n315 VDD.n236 0.491846
R28589 VDD.n328 VDD.n327 0.488781
R28590 VDD.n238 VDD.n223 0.481269
R28591 VDD.n2163 VDD.n2162 0.474085
R28592 VDD.n2707 VDD.n2706 0.457643
R28593 VDD.n438 VDD.n437 0.440923
R28594 VDD.n3500 VDD.n2926 0.440094
R28595 VDD.n401 VDD.n400 0.438
R28596 VDD.n3798 VDD.n3797 0.435058
R28597 VDD.n9 VDD.n8 0.433948
R28598 VDD.n4443 VDD.n3672 0.42364
R28599 VDD.n2659 VDD.n2302 0.42364
R28600 VDD.n1324 VDD.n1323 0.42364
R28601 VDD.n1317 VDD.n1316 0.42364
R28602 VDD.n2834 VDD.n2225 0.417164
R28603 VDD.n3827 VDD.n3824 0.417114
R28604 VDD.n330 VDD.n329 0.393625
R28605 VDD.n78 VDD.n77 0.388
R28606 VDD.n40 VDD.n27 0.388
R28607 VDD.n158 VDD.n156 0.383913
R28608 VDD.n1257 VDD.n438 0.376992
R28609 VDD.n4116 VDD.n3730 0.376971
R28610 VDD.n4404 VDD.n4403 0.376971
R28611 VDD.n3485 VDD.n2936 0.376971
R28612 VDD.n1379 VDD.n1362 0.376971
R28613 VDD.n2056 VDD.n1404 0.376971
R28614 VDD.n2047 VDD.n1406 0.376971
R28615 VDD.n2015 VDD.n2014 0.376971
R28616 VDD.n2007 VDD.n2006 0.376971
R28617 VDD.n1750 VDD.n1548 0.376971
R28618 VDD.n1217 VDD.n1216 0.376971
R28619 VDD.n497 VDD.n496 0.376971
R28620 VDD.n3888 VDD.n3821 0.369731
R28621 VDD.n3901 VDD.n3900 0.369731
R28622 VDD.n4279 VDD.n3685 0.369731
R28623 VDD.n4289 VDD.n3681 0.369731
R28624 VDD.n3126 VDD.n3125 0.369731
R28625 VDD.n3108 VDD.n3077 0.369731
R28626 VDD.n3104 VDD.n3079 0.369731
R28627 VDD.n3087 VDD.n3086 0.369731
R28628 VDD.n3636 VDD.n3583 0.369731
R28629 VDD.n3617 VDD.n3589 0.369731
R28630 VDD.n2440 VDD.n2439 0.369731
R28631 VDD.n2434 VDD.n2415 0.369731
R28632 VDD.n2432 VDD.n2431 0.369731
R28633 VDD.n2418 VDD.n2398 0.369731
R28634 VDD.n1613 VDD.n1612 0.369731
R28635 VDD.n1608 VDD.n1591 0.369731
R28636 VDD.n159 VDD.n158 0.359875
R28637 VDD.n3964 VDD.n3963 0.358087
R28638 VDD.n1156 VDD.n1155 0.358087
R28639 VDD.n1161 VDD.n1160 0.356056
R28640 VDD.n2377 VDD.n2368 0.354995
R28641 VDD.n2560 VDD.n2368 0.353728
R28642 VDD.n2162 VDD.n2161 0.353728
R28643 VDD.n310 VDD.n240 0.3505
R28644 VDD.n287 VDD.n286 0.3505
R28645 VDD.n307 VDD.n306 0.3505
R28646 VDD.n283 VDD.n244 0.3505
R28647 VDD.n303 VDD.n237 0.3505
R28648 VDD.n290 VDD.n245 0.3505
R28649 VDD.n311 VDD.n310 0.338
R28650 VDD.n299 VDD.n240 0.338
R28651 VDD.n299 VDD.n298 0.338
R28652 VDD.n298 VDD.n243 0.338
R28653 VDD.n287 VDD.n243 0.338
R28654 VDD.n286 VDD.n246 0.338
R28655 VDD.n275 VDD.n246 0.338
R28656 VDD.n307 VDD.n239 0.338
R28657 VDD.n306 VDD.n241 0.338
R28658 VDD.n295 VDD.n241 0.338
R28659 VDD.n295 VDD.n294 0.338
R28660 VDD.n294 VDD.n244 0.338
R28661 VDD.n283 VDD.n282 0.338
R28662 VDD.n282 VDD.n247 0.338
R28663 VDD.n273 VDD.n247 0.338
R28664 VDD.n314 VDD.n237 0.338
R28665 VDD.n303 VDD.n302 0.338
R28666 VDD.n302 VDD.n242 0.338
R28667 VDD.n291 VDD.n242 0.338
R28668 VDD.n291 VDD.n290 0.338
R28669 VDD.n279 VDD.n245 0.338
R28670 VDD.n279 VDD.n278 0.338
R28671 VDD.n317 VDD.n316 0.332643
R28672 VDD.n3943 VDD.n3942 0.317855
R28673 VDD.n3943 VDD.n3807 0.317855
R28674 VDD.n404 VDD.n394 0.3105
R28675 VDD.n4014 VDD.n3769 0.310308
R28676 VDD.n4223 VDD.n4192 0.305262
R28677 VDD.n4219 VDD.n4218 0.305262
R28678 VDD.n4213 VDD.n4196 0.305262
R28679 VDD.n4230 VDD.n4229 0.305262
R28680 VDD.n4137 VDD.n3723 0.305262
R28681 VDD.n4071 VDD.n4070 0.305262
R28682 VDD.n4073 VDD.n4072 0.305262
R28683 VDD.n4083 VDD.n4082 0.305262
R28684 VDD.n4360 VDD.n4310 0.305262
R28685 VDD.n4350 VDD.n4315 0.305262
R28686 VDD.n4254 VDD.n4253 0.305262
R28687 VDD.n4015 VDD.n4014 0.305262
R28688 VDD.n4023 VDD.n3766 0.305262
R28689 VDD.n4056 VDD.n4055 0.305262
R28690 VDD.n4066 VDD.n4065 0.305262
R28691 VDD.n3969 VDD.n3787 0.305262
R28692 VDD.n3954 VDD.n3802 0.305262
R28693 VDD.n3352 VDD.n3350 0.305262
R28694 VDD.n3407 VDD.n3406 0.305262
R28695 VDD.n3256 VDD.n3255 0.305262
R28696 VDD.n3137 VDD.n3136 0.305262
R28697 VDD.n3145 VDD.n3034 0.305262
R28698 VDD.n3190 VDD.n3189 0.305262
R28699 VDD.n2817 VDD.n2816 0.305262
R28700 VDD.n2823 VDD.n2822 0.305262
R28701 VDD.n2793 VDD.n2792 0.305262
R28702 VDD.n2724 VDD.n2723 0.305262
R28703 VDD.n2730 VDD.n2729 0.305262
R28704 VDD.n2702 VDD.n2701 0.305262
R28705 VDD.n2709 VDD.n2708 0.305262
R28706 VDD.n2694 VDD.n2693 0.305262
R28707 VDD.n2308 VDD.n2306 0.305262
R28708 VDD.n2657 VDD.n2656 0.305262
R28709 VDD.n2566 VDD.n2565 0.305262
R28710 VDD.n2553 VDD.n2378 0.305262
R28711 VDD.n2061 VDD.n1270 0.305262
R28712 VDD.n2032 VDD.n2031 0.305262
R28713 VDD.n2037 VDD.n2036 0.305262
R28714 VDD.n1962 VDD.n1961 0.305262
R28715 VDD.n1969 VDD.n1443 0.305262
R28716 VDD.n1919 VDD.n1466 0.305262
R28717 VDD.n1931 VDD.n1461 0.305262
R28718 VDD.n1850 VDD.n1849 0.305262
R28719 VDD.n1856 VDD.n1855 0.305262
R28720 VDD.n1249 VDD.n446 0.305262
R28721 VDD.n1239 VDD.n1238 0.305262
R28722 VDD.n532 VDD.n530 0.305262
R28723 VDD.n582 VDD.n581 0.305262
R28724 VDD.n1168 VDD.n1167 0.305262
R28725 VDD.n1166 VDD.n621 0.305262
R28726 VDD.n1180 VDD.n619 0.305262
R28727 VDD.n1164 VDD.n623 0.305262
R28728 VDD.n1145 VDD.n1144 0.305262
R28729 VDD.n1150 VDD.n642 0.305262
R28730 VDD.n1134 VDD.n1132 0.305262
R28731 VDD.n1133 VDD.n655 0.305262
R28732 VDD.n1108 VDD.n1107 0.305262
R28733 VDD.n1114 VDD.n1113 0.305262
R28734 VDD.n1053 VDD.n1052 0.305262
R28735 VDD.n1060 VDD.n1059 0.305262
R28736 VDD.n1015 VDD.n1014 0.305262
R28737 VDD.n1026 VDD.n1024 0.305262
R28738 VDD.n995 VDD.n994 0.305262
R28739 VDD.n1005 VDD.n719 0.305262
R28740 VDD.n968 VDD.n967 0.305262
R28741 VDD.n972 VDD.n728 0.305262
R28742 VDD.n950 VDD.n949 0.305262
R28743 VDD.n955 VDD.n733 0.305262
R28744 VDD.n925 VDD.n924 0.305262
R28745 VDD.n934 VDD.n742 0.305262
R28746 VDD.n750 VDD.n749 0.305262
R28747 VDD.n920 VDD.n919 0.305262
R28748 VDD.n806 VDD.n804 0.305262
R28749 VDD.n522 VDD.n521 0.305262
R28750 VDD.n2573 VDD.n2572 0.3005
R28751 VDD.n2529 VDD.n2528 0.3005
R28752 VDD.n3912 VDD.n3813 0.298074
R28753 VDD.n3881 VDD.n3824 0.29768
R28754 VDD.n4248 VDD.n4247 0.29768
R28755 VDD.n4247 VDD.n4246 0.29768
R28756 VDD.n3639 VDD.n3576 0.29768
R28757 VDD.n3635 VDD.n3576 0.29768
R28758 VDD.n3922 VDD.n3813 0.297291
R28759 VDD.n3965 VDD.n3964 0.297291
R28760 VDD.n2843 VDD.n2225 0.297291
R28761 VDD.n1157 VDD.n1156 0.297291
R28762 VDD.n181 VDD.n180 0.278
R28763 VDD.n4244 VDD.n4243 0.254468
R28764 VDD.n4132 VDD.n4131 0.254468
R28765 VDD.n3196 VDD.n3195 0.254468
R28766 VDD.n3963 VDD.n3962 0.240317
R28767 VDD.n4097 VDD.n4096 0.239726
R28768 VDD.n4308 VDD.n4307 0.239726
R28769 VDD.n3064 VDD.n3063 0.239726
R28770 VDD.n3128 VDD.n3067 0.239726
R28771 VDD.n2925 VDD.n2921 0.239726
R28772 VDD.n2355 VDD.n2353 0.239726
R28773 VDD.n1753 VDD.n1549 0.239726
R28774 VDD.n1947 VDD.n1946 0.239726
R28775 VDD.n802 VDD.n775 0.239726
R28776 VDD.n647 VDD.n644 0.239726
R28777 VDD.n1225 VDD.n590 0.239726
R28778 VDD.n2835 VDD.n2834 0.239726
R28779 VDD.n2163 VDD.n2100 0.239726
R28780 VDD.n527 VDD.n526 0.239726
R28781 VDD.n3872 VDD.n3827 0.239381
R28782 VDD.n4096 VDD.n4095 0.239381
R28783 VDD.n4307 VDD.n4306 0.239381
R28784 VDD.n3063 VDD.n3062 0.239381
R28785 VDD.n3067 VDD.n3064 0.239381
R28786 VDD.n3498 VDD.n2925 0.239381
R28787 VDD.n2581 VDD.n2355 0.239381
R28788 VDD.n1742 VDD.n1549 0.239381
R28789 VDD.n1946 VDD.n1945 0.239381
R28790 VDD.n803 VDD.n802 0.239381
R28791 VDD.n651 VDD.n647 0.239381
R28792 VDD.n1221 VDD.n590 0.239381
R28793 VDD.n526 VDD.n525 0.239381
R28794 VDD.n3880 VDD.n3879 0.227049
R28795 VDD.n3886 VDD.n3885 0.227049
R28796 VDD.n4026 VDD.n3764 0.227049
R28797 VDD.n4040 VDD.n4039 0.227049
R28798 VDD.n3921 VDD.n3920 0.227049
R28799 VDD.n3927 VDD.n3926 0.227049
R28800 VDD.n2340 VDD.n2339 0.227049
R28801 VDD.n2607 VDD.n2606 0.227049
R28802 VDD.n2455 VDD.n2407 0.227049
R28803 VDD.n2441 VDD.n2411 0.227049
R28804 VDD.n1627 VDD.n1626 0.227049
R28805 VDD.n1614 VDD.n1590 0.227049
R28806 VDD.n1339 VDD.n1338 0.227049
R28807 VDD.n1330 VDD.n1329 0.227049
R28808 VDD.n399 VDD.n395 0.21925
R28809 VDD.n4329 VDD.n4328 0.21207
R28810 VDD.n4448 VDD.n4447 0.21207
R28811 VDD.n3672 VDD.n3670 0.21207
R28812 VDD.n4299 VDD.n4298 0.21207
R28813 VDD.n2832 VDD.n2831 0.21207
R28814 VDD.n2679 VDD.n2678 0.21207
R28815 VDD.n2522 VDD.n2521 0.21207
R28816 VDD.n1596 VDD.n1593 0.21207
R28817 VDD.n1328 VDD.n1279 0.21207
R28818 VDD.n1322 VDD.n1281 0.21207
R28819 VDD.n1318 VDD.n1317 0.21207
R28820 VDD.n4128 VDD.n4127 0.203675
R28821 VDD.n4082 VDD.n4081 0.203675
R28822 VDD.n4265 VDD.n3689 0.203675
R28823 VDD.n3249 VDD.n3248 0.203675
R28824 VDD.n3143 VDD.n3142 0.203675
R28825 VDD.n2786 VDD.n2785 0.203675
R28826 VDD.n2564 VDD.n2563 0.203675
R28827 VDD.n2546 VDD.n2545 0.203675
R28828 VDD.n2156 VDD.n2155 0.203675
R28829 VDD.n2068 VDD.n2067 0.203675
R28830 VDD.n927 VDD.n926 0.203675
R28831 VDD.n820 VDD.n819 0.203675
R28832 VDD.n160 VDD.n103 0.202674
R28833 VDD.n236 VDD.n235 0.184982
R28834 VDD.n2590 VDD.n2347 0.180304
R28835 VDD.n2347 VDD.n2344 0.180304
R28836 VDD.n905 VDD.n751 0.180304
R28837 VDD.n751 VDD.n748 0.180304
R28838 VDD.n1155 VDD.n631 0.180304
R28839 VDD.n3962 VDD.n3961 0.180304
R28840 VDD.n4184 VDD.n4180 0.180304
R28841 VDD.n4235 VDD.n4184 0.180304
R28842 VDD.n2498 VDD.n2497 0.180304
R28843 VDD.n2498 VDD.n2395 0.180304
R28844 VDD.n1679 VDD.n1678 0.180304
R28845 VDD.n1679 VDD.n1573 0.180304
R28846 VDD.n1341 VDD.n1269 0.180304
R28847 VDD.n1341 VDD.n1340 0.180304
R28848 VDD.n1128 VDD.n1127 0.180304
R28849 VDD.n1129 VDD.n1128 0.180304
R28850 VDD VDD.n4467 0.175722
R28851 VDD.n4467 VDD.n3658 0.1603
R28852 VDD.n3658 VDD.n2892 0.1603
R28853 VDD.n2892 VDD.n2087 0.1603
R28854 VDD.n2087 VDD.n1257 0.1603
R28855 VDD.n169 VDD.n168 0.159538
R28856 VDD.n86 VDD.n85 0.15831
R28857 VDD.n2848 VDD.n2847 0.152881
R28858 VDD.n2849 VDD.n2848 0.152881
R28859 VDD.n2651 VDD.n2650 0.152881
R28860 VDD.n2554 VDD.n2553 0.152881
R28861 VDD.n407 VDD.n406 0.148457
R28862 VDD.n143 VDD.n88 0.148119
R28863 VDD.n274 VDD.n248 0.142484
R28864 VDD.n277 VDD.n276 0.142484
R28865 VDD.n281 VDD.n280 0.142484
R28866 VDD.n285 VDD.n284 0.142484
R28867 VDD.n289 VDD.n288 0.142484
R28868 VDD.n293 VDD.n292 0.142484
R28869 VDD.n297 VDD.n296 0.142484
R28870 VDD.n301 VDD.n300 0.142484
R28871 VDD.n305 VDD.n304 0.142484
R28872 VDD.n309 VDD.n308 0.142484
R28873 VDD.n313 VDD.n312 0.142484
R28874 VDD.n168 VDD.n167 0.141672
R28875 VDD.n404 VDD.n403 0.141125
R28876 VDD.n86 VDD.n81 0.132625
R28877 VDD.n2732 VDD.n2730 0.130856
R28878 VDD.n581 VDD.n535 0.130856
R28879 VDD.n70 VDD.n64 0.122868
R28880 VDD.n33 VDD.n28 0.122868
R28881 VDD.n7 VDD.n6 0.120751
R28882 VDD.n84 VDD.n83 0.120751
R28883 VDD.n3859 VDD.n3858 0.120292
R28884 VDD.n3860 VDD.n3859 0.120292
R28885 VDD.n3860 VDD.n3843 0.120292
R28886 VDD.n3864 VDD.n3843 0.120292
R28887 VDD.n3865 VDD.n3864 0.120292
R28888 VDD.n3866 VDD.n3865 0.120292
R28889 VDD.n3866 VDD.n3834 0.120292
R28890 VDD.n3870 VDD.n3834 0.120292
R28891 VDD.n3871 VDD.n3870 0.120292
R28892 VDD.n3872 VDD.n3871 0.120292
R28893 VDD.n3882 VDD.n3881 0.120292
R28894 VDD.n3883 VDD.n3882 0.120292
R28895 VDD.n3883 VDD.n3822 0.120292
R28896 VDD.n3889 VDD.n3822 0.120292
R28897 VDD.n3890 VDD.n3889 0.120292
R28898 VDD.n3890 VDD.n3820 0.120292
R28899 VDD.n3895 VDD.n3820 0.120292
R28900 VDD.n3896 VDD.n3895 0.120292
R28901 VDD.n3897 VDD.n3896 0.120292
R28902 VDD.n3897 VDD.n3818 0.120292
R28903 VDD.n3902 VDD.n3818 0.120292
R28904 VDD.n3903 VDD.n3902 0.120292
R28905 VDD.n3904 VDD.n3903 0.120292
R28906 VDD.n3904 VDD.n3815 0.120292
R28907 VDD.n3910 VDD.n3815 0.120292
R28908 VDD.n3911 VDD.n3910 0.120292
R28909 VDD.n3912 VDD.n3911 0.120292
R28910 VDD.n3923 VDD.n3922 0.120292
R28911 VDD.n3924 VDD.n3923 0.120292
R28912 VDD.n3924 VDD.n3811 0.120292
R28913 VDD.n3931 VDD.n3811 0.120292
R28914 VDD.n3932 VDD.n3931 0.120292
R28915 VDD.n3933 VDD.n3932 0.120292
R28916 VDD.n3933 VDD.n3809 0.120292
R28917 VDD.n3938 VDD.n3809 0.120292
R28918 VDD.n3939 VDD.n3938 0.120292
R28919 VDD.n3940 VDD.n3939 0.120292
R28920 VDD.n3940 VDD.n3806 0.120292
R28921 VDD.n3948 VDD.n3806 0.120292
R28922 VDD.n3949 VDD.n3948 0.120292
R28923 VDD.n3950 VDD.n3949 0.120292
R28924 VDD.n3950 VDD.n3803 0.120292
R28925 VDD.n3955 VDD.n3803 0.120292
R28926 VDD.n3956 VDD.n3955 0.120292
R28927 VDD.n3956 VDD.n3801 0.120292
R28928 VDD.n3961 VDD.n3801 0.120292
R28929 VDD.n3965 VDD.n3788 0.120292
R28930 VDD.n3971 VDD.n3788 0.120292
R28931 VDD.n3972 VDD.n3971 0.120292
R28932 VDD.n3973 VDD.n3972 0.120292
R28933 VDD.n3973 VDD.n3785 0.120292
R28934 VDD.n3977 VDD.n3785 0.120292
R28935 VDD.n3978 VDD.n3977 0.120292
R28936 VDD.n3980 VDD.n3978 0.120292
R28937 VDD.n3980 VDD.n3979 0.120292
R28938 VDD.n3979 VDD.n3781 0.120292
R28939 VDD.n3991 VDD.n3781 0.120292
R28940 VDD.n3992 VDD.n3991 0.120292
R28941 VDD.n3993 VDD.n3992 0.120292
R28942 VDD.n3993 VDD.n3778 0.120292
R28943 VDD.n3778 VDD.n3777 0.120292
R28944 VDD.n3777 VDD.n3775 0.120292
R28945 VDD.n3999 VDD.n3775 0.120292
R28946 VDD.n4000 VDD.n3999 0.120292
R28947 VDD.n4001 VDD.n4000 0.120292
R28948 VDD.n4001 VDD.n3772 0.120292
R28949 VDD.n4005 VDD.n3772 0.120292
R28950 VDD.n4006 VDD.n4005 0.120292
R28951 VDD.n4007 VDD.n4006 0.120292
R28952 VDD.n4007 VDD.n3770 0.120292
R28953 VDD.n4012 VDD.n3770 0.120292
R28954 VDD.n4013 VDD.n4012 0.120292
R28955 VDD.n4013 VDD.n3767 0.120292
R28956 VDD.n4021 VDD.n3767 0.120292
R28957 VDD.n4022 VDD.n4021 0.120292
R28958 VDD.n4022 VDD.n3765 0.120292
R28959 VDD.n4027 VDD.n3765 0.120292
R28960 VDD.n4028 VDD.n4027 0.120292
R28961 VDD.n4028 VDD.n3763 0.120292
R28962 VDD.n4034 VDD.n3763 0.120292
R28963 VDD.n4035 VDD.n4034 0.120292
R28964 VDD.n4036 VDD.n4035 0.120292
R28965 VDD.n4036 VDD.n3761 0.120292
R28966 VDD.n4041 VDD.n3761 0.120292
R28967 VDD.n4042 VDD.n4041 0.120292
R28968 VDD.n4043 VDD.n4042 0.120292
R28969 VDD.n4043 VDD.n3759 0.120292
R28970 VDD.n4049 VDD.n3759 0.120292
R28971 VDD.n4050 VDD.n4049 0.120292
R28972 VDD.n4051 VDD.n4050 0.120292
R28973 VDD.n4051 VDD.n3756 0.120292
R28974 VDD.n4057 VDD.n3756 0.120292
R28975 VDD.n4058 VDD.n4057 0.120292
R28976 VDD.n4058 VDD.n3754 0.120292
R28977 VDD.n4067 VDD.n3754 0.120292
R28978 VDD.n4068 VDD.n4067 0.120292
R28979 VDD.n4069 VDD.n4068 0.120292
R28980 VDD.n4069 VDD.n3751 0.120292
R28981 VDD.n4077 VDD.n3751 0.120292
R28982 VDD.n4078 VDD.n4077 0.120292
R28983 VDD.n4079 VDD.n4078 0.120292
R28984 VDD.n4079 VDD.n3749 0.120292
R28985 VDD.n4085 VDD.n3749 0.120292
R28986 VDD.n4086 VDD.n4085 0.120292
R28987 VDD.n4086 VDD.n3745 0.120292
R28988 VDD.n4090 VDD.n3745 0.120292
R28989 VDD.n4091 VDD.n4090 0.120292
R28990 VDD.n4091 VDD.n3742 0.120292
R28991 VDD.n4095 VDD.n3742 0.120292
R28992 VDD.n4097 VDD.n3736 0.120292
R28993 VDD.n4105 VDD.n3736 0.120292
R28994 VDD.n4106 VDD.n4105 0.120292
R28995 VDD.n4107 VDD.n4106 0.120292
R28996 VDD.n4107 VDD.n3733 0.120292
R28997 VDD.n3733 VDD.n3731 0.120292
R28998 VDD.n4114 VDD.n3731 0.120292
R28999 VDD.n4115 VDD.n4114 0.120292
R29000 VDD.n4115 VDD.n3728 0.120292
R29001 VDD.n4120 VDD.n3728 0.120292
R29002 VDD.n4121 VDD.n4120 0.120292
R29003 VDD.n4123 VDD.n4121 0.120292
R29004 VDD.n4123 VDD.n4122 0.120292
R29005 VDD.n4122 VDD.n3724 0.120292
R29006 VDD.n4133 VDD.n3724 0.120292
R29007 VDD.n4136 VDD.n4133 0.120292
R29008 VDD.n4136 VDD.n4135 0.120292
R29009 VDD.n4135 VDD.n4134 0.120292
R29010 VDD.n4134 VDD.n3718 0.120292
R29011 VDD.n4145 VDD.n3718 0.120292
R29012 VDD.n4146 VDD.n4145 0.120292
R29013 VDD.n4146 VDD.n3715 0.120292
R29014 VDD.n4153 VDD.n3715 0.120292
R29015 VDD.n4154 VDD.n4153 0.120292
R29016 VDD.n4155 VDD.n4154 0.120292
R29017 VDD.n4155 VDD.n3713 0.120292
R29018 VDD.n4160 VDD.n3713 0.120292
R29019 VDD.n4161 VDD.n4160 0.120292
R29020 VDD.n4161 VDD.n3711 0.120292
R29021 VDD.n3711 VDD.n3709 0.120292
R29022 VDD.n4168 VDD.n3709 0.120292
R29023 VDD.n4169 VDD.n4168 0.120292
R29024 VDD.n4169 VDD.n3705 0.120292
R29025 VDD.n4173 VDD.n3705 0.120292
R29026 VDD.n4174 VDD.n4173 0.120292
R29027 VDD.n4174 VDD.n3702 0.120292
R29028 VDD.n4178 VDD.n3702 0.120292
R29029 VDD.n4179 VDD.n4178 0.120292
R29030 VDD.n4248 VDD.n4179 0.120292
R29031 VDD.n4246 VDD.n4180 0.120292
R29032 VDD.n4235 VDD.n4234 0.120292
R29033 VDD.n4234 VDD.n4187 0.120292
R29034 VDD.n4228 VDD.n4187 0.120292
R29035 VDD.n4228 VDD.n4227 0.120292
R29036 VDD.n4227 VDD.n4226 0.120292
R29037 VDD.n4226 VDD.n4191 0.120292
R29038 VDD.n4222 VDD.n4191 0.120292
R29039 VDD.n4222 VDD.n4221 0.120292
R29040 VDD.n4221 VDD.n4193 0.120292
R29041 VDD.n4216 VDD.n4193 0.120292
R29042 VDD.n4216 VDD.n4215 0.120292
R29043 VDD.n4215 VDD.n4214 0.120292
R29044 VDD.n4214 VDD.n4195 0.120292
R29045 VDD.n4210 VDD.n4195 0.120292
R29046 VDD.n4210 VDD.n4209 0.120292
R29047 VDD.n4209 VDD.n4199 0.120292
R29048 VDD.n4203 VDD.n4199 0.120292
R29049 VDD.n4203 VDD.n4202 0.120292
R29050 VDD.n4202 VDD.n3695 0.120292
R29051 VDD.n4255 VDD.n3695 0.120292
R29052 VDD.n4256 VDD.n4255 0.120292
R29053 VDD.n4257 VDD.n4256 0.120292
R29054 VDD.n4257 VDD.n3690 0.120292
R29055 VDD.n4263 VDD.n3690 0.120292
R29056 VDD.n4264 VDD.n4263 0.120292
R29057 VDD.n4264 VDD.n3688 0.120292
R29058 VDD.n4274 VDD.n3688 0.120292
R29059 VDD.n4275 VDD.n4274 0.120292
R29060 VDD.n4275 VDD.n3686 0.120292
R29061 VDD.n4280 VDD.n3686 0.120292
R29062 VDD.n4281 VDD.n4280 0.120292
R29063 VDD.n4281 VDD.n3684 0.120292
R29064 VDD.n4285 VDD.n3684 0.120292
R29065 VDD.n4286 VDD.n4285 0.120292
R29066 VDD.n4286 VDD.n3682 0.120292
R29067 VDD.n4291 VDD.n3682 0.120292
R29068 VDD.n4292 VDD.n4291 0.120292
R29069 VDD.n4293 VDD.n4292 0.120292
R29070 VDD.n4293 VDD.n3680 0.120292
R29071 VDD.n4300 VDD.n3680 0.120292
R29072 VDD.n4301 VDD.n4300 0.120292
R29073 VDD.n4301 VDD.n3678 0.120292
R29074 VDD.n4306 VDD.n3678 0.120292
R29075 VDD.n4359 VDD.n4308 0.120292
R29076 VDD.n4359 VDD.n4358 0.120292
R29077 VDD.n4358 VDD.n4311 0.120292
R29078 VDD.n4353 VDD.n4311 0.120292
R29079 VDD.n4353 VDD.n4352 0.120292
R29080 VDD.n4352 VDD.n4351 0.120292
R29081 VDD.n4351 VDD.n4314 0.120292
R29082 VDD.n4346 VDD.n4314 0.120292
R29083 VDD.n4346 VDD.n4345 0.120292
R29084 VDD.n4345 VDD.n4344 0.120292
R29085 VDD.n4344 VDD.n4317 0.120292
R29086 VDD.n4339 VDD.n4317 0.120292
R29087 VDD.n4339 VDD.n4338 0.120292
R29088 VDD.n4338 VDD.n4320 0.120292
R29089 VDD.n4333 VDD.n4320 0.120292
R29090 VDD.n4333 VDD.n4332 0.120292
R29091 VDD.n4332 VDD.n4331 0.120292
R29092 VDD.n4331 VDD.n4322 0.120292
R29093 VDD.n4326 VDD.n4322 0.120292
R29094 VDD.n4451 VDD.n4450 0.120292
R29095 VDD.n4450 VDD.n3668 0.120292
R29096 VDD.n4445 VDD.n3668 0.120292
R29097 VDD.n4445 VDD.n4444 0.120292
R29098 VDD.n4444 VDD.n3671 0.120292
R29099 VDD.n4440 VDD.n3671 0.120292
R29100 VDD.n4440 VDD.n4439 0.120292
R29101 VDD.n4439 VDD.n4438 0.120292
R29102 VDD.n4438 VDD.n4366 0.120292
R29103 VDD.n4433 VDD.n4366 0.120292
R29104 VDD.n4433 VDD.n4432 0.120292
R29105 VDD.n4432 VDD.n4371 0.120292
R29106 VDD.n4428 VDD.n4371 0.120292
R29107 VDD.n4428 VDD.n4427 0.120292
R29108 VDD.n4427 VDD.n4426 0.120292
R29109 VDD.n4426 VDD.n4374 0.120292
R29110 VDD.n4422 VDD.n4374 0.120292
R29111 VDD.n4422 VDD.n4421 0.120292
R29112 VDD.n4421 VDD.n4377 0.120292
R29113 VDD.n4378 VDD.n4377 0.120292
R29114 VDD.n4414 VDD.n4378 0.120292
R29115 VDD.n4414 VDD.n4413 0.120292
R29116 VDD.n4413 VDD.n4412 0.120292
R29117 VDD.n4412 VDD.n4382 0.120292
R29118 VDD.n4408 VDD.n4382 0.120292
R29119 VDD.n4408 VDD.n4407 0.120292
R29120 VDD.n4407 VDD.n4406 0.120292
R29121 VDD.n4406 VDD.n4386 0.120292
R29122 VDD.n4400 VDD.n4386 0.120292
R29123 VDD.n4400 VDD.n4399 0.120292
R29124 VDD.n3056 VDD.n3046 0.120292
R29125 VDD.n3062 VDD.n3046 0.120292
R29126 VDD.n3128 VDD.n3127 0.120292
R29127 VDD.n3127 VDD.n3072 0.120292
R29128 VDD.n3122 VDD.n3072 0.120292
R29129 VDD.n3122 VDD.n3121 0.120292
R29130 VDD.n3121 VDD.n3074 0.120292
R29131 VDD.n3116 VDD.n3074 0.120292
R29132 VDD.n3116 VDD.n3115 0.120292
R29133 VDD.n3115 VDD.n3114 0.120292
R29134 VDD.n3114 VDD.n3076 0.120292
R29135 VDD.n3110 VDD.n3076 0.120292
R29136 VDD.n3110 VDD.n3109 0.120292
R29137 VDD.n3109 VDD.n3078 0.120292
R29138 VDD.n3103 VDD.n3078 0.120292
R29139 VDD.n3103 VDD.n3102 0.120292
R29140 VDD.n3102 VDD.n3080 0.120292
R29141 VDD.n3097 VDD.n3080 0.120292
R29142 VDD.n3097 VDD.n3096 0.120292
R29143 VDD.n3096 VDD.n3082 0.120292
R29144 VDD.n3092 VDD.n3082 0.120292
R29145 VDD.n3092 VDD.n3091 0.120292
R29146 VDD.n3091 VDD.n3090 0.120292
R29147 VDD.n3090 VDD.n3084 0.120292
R29148 VDD.n3085 VDD.n3084 0.120292
R29149 VDD.n3085 VDD.n3038 0.120292
R29150 VDD.n3138 VDD.n3038 0.120292
R29151 VDD.n3139 VDD.n3138 0.120292
R29152 VDD.n3140 VDD.n3139 0.120292
R29153 VDD.n3140 VDD.n3035 0.120292
R29154 VDD.n3148 VDD.n3035 0.120292
R29155 VDD.n3149 VDD.n3148 0.120292
R29156 VDD.n3150 VDD.n3149 0.120292
R29157 VDD.n3150 VDD.n3032 0.120292
R29158 VDD.n3156 VDD.n3032 0.120292
R29159 VDD.n3157 VDD.n3156 0.120292
R29160 VDD.n3158 VDD.n3157 0.120292
R29161 VDD.n3158 VDD.n3030 0.120292
R29162 VDD.n3163 VDD.n3030 0.120292
R29163 VDD.n3164 VDD.n3163 0.120292
R29164 VDD.n3165 VDD.n3164 0.120292
R29165 VDD.n3165 VDD.n3028 0.120292
R29166 VDD.n3171 VDD.n3028 0.120292
R29167 VDD.n3172 VDD.n3171 0.120292
R29168 VDD.n3172 VDD.n3025 0.120292
R29169 VDD.n3176 VDD.n3025 0.120292
R29170 VDD.n3177 VDD.n3176 0.120292
R29171 VDD.n3178 VDD.n3177 0.120292
R29172 VDD.n3178 VDD.n3023 0.120292
R29173 VDD.n3183 VDD.n3023 0.120292
R29174 VDD.n3184 VDD.n3183 0.120292
R29175 VDD.n3184 VDD.n3020 0.120292
R29176 VDD.n3191 VDD.n3020 0.120292
R29177 VDD.n3192 VDD.n3191 0.120292
R29178 VDD.n3193 VDD.n3192 0.120292
R29179 VDD.n3193 VDD.n3018 0.120292
R29180 VDD.n3199 VDD.n3018 0.120292
R29181 VDD.n3200 VDD.n3199 0.120292
R29182 VDD.n3201 VDD.n3200 0.120292
R29183 VDD.n3201 VDD.n3016 0.120292
R29184 VDD.n3016 VDD.n3013 0.120292
R29185 VDD.n3206 VDD.n3013 0.120292
R29186 VDD.n3207 VDD.n3206 0.120292
R29187 VDD.n3208 VDD.n3207 0.120292
R29188 VDD.n3208 VDD.n3009 0.120292
R29189 VDD.n3213 VDD.n3009 0.120292
R29190 VDD.n3214 VDD.n3213 0.120292
R29191 VDD.n3215 VDD.n3214 0.120292
R29192 VDD.n3215 VDD.n3007 0.120292
R29193 VDD.n3007 VDD.n3006 0.120292
R29194 VDD.n3006 VDD.n3005 0.120292
R29195 VDD.n3221 VDD.n3005 0.120292
R29196 VDD.n3222 VDD.n3221 0.120292
R29197 VDD.n3223 VDD.n3222 0.120292
R29198 VDD.n3223 VDD.n3002 0.120292
R29199 VDD.n3002 VDD.n3001 0.120292
R29200 VDD.n3001 VDD.n2999 0.120292
R29201 VDD.n2999 VDD.n2998 0.120292
R29202 VDD.n2998 VDD.n2996 0.120292
R29203 VDD.n3231 VDD.n2996 0.120292
R29204 VDD.n3232 VDD.n3231 0.120292
R29205 VDD.n3293 VDD.n3232 0.120292
R29206 VDD.n3293 VDD.n3292 0.120292
R29207 VDD.n3292 VDD.n3291 0.120292
R29208 VDD.n3291 VDD.n3233 0.120292
R29209 VDD.n3287 VDD.n3233 0.120292
R29210 VDD.n3287 VDD.n3286 0.120292
R29211 VDD.n3286 VDD.n3285 0.120292
R29212 VDD.n3285 VDD.n3235 0.120292
R29213 VDD.n3280 VDD.n3235 0.120292
R29214 VDD.n3280 VDD.n3279 0.120292
R29215 VDD.n3279 VDD.n3278 0.120292
R29216 VDD.n3278 VDD.n3237 0.120292
R29217 VDD.n3273 VDD.n3237 0.120292
R29218 VDD.n3273 VDD.n3272 0.120292
R29219 VDD.n3272 VDD.n3271 0.120292
R29220 VDD.n3271 VDD.n3239 0.120292
R29221 VDD.n3267 VDD.n3239 0.120292
R29222 VDD.n3267 VDD.n3266 0.120292
R29223 VDD.n3266 VDD.n3265 0.120292
R29224 VDD.n3265 VDD.n3242 0.120292
R29225 VDD.n3260 VDD.n3242 0.120292
R29226 VDD.n3260 VDD.n3259 0.120292
R29227 VDD.n3259 VDD.n3258 0.120292
R29228 VDD.n3258 VDD.n3244 0.120292
R29229 VDD.n3252 VDD.n3244 0.120292
R29230 VDD.n3252 VDD.n3251 0.120292
R29231 VDD.n3251 VDD.n3250 0.120292
R29232 VDD.n3250 VDD.n2992 0.120292
R29233 VDD.n3298 VDD.n2992 0.120292
R29234 VDD.n3299 VDD.n3298 0.120292
R29235 VDD.n3299 VDD.n2988 0.120292
R29236 VDD.n3303 VDD.n2988 0.120292
R29237 VDD.n3304 VDD.n3303 0.120292
R29238 VDD.n3305 VDD.n3304 0.120292
R29239 VDD.n3305 VDD.n2985 0.120292
R29240 VDD.n3309 VDD.n2985 0.120292
R29241 VDD.n3310 VDD.n3309 0.120292
R29242 VDD.n3310 VDD.n2982 0.120292
R29243 VDD.n3316 VDD.n2982 0.120292
R29244 VDD.n3317 VDD.n3316 0.120292
R29245 VDD.n3317 VDD.n2979 0.120292
R29246 VDD.n2979 VDD.n2978 0.120292
R29247 VDD.n2978 VDD.n2977 0.120292
R29248 VDD.n3325 VDD.n2977 0.120292
R29249 VDD.n3326 VDD.n3325 0.120292
R29250 VDD.n3327 VDD.n3326 0.120292
R29251 VDD.n3327 VDD.n2974 0.120292
R29252 VDD.n3332 VDD.n2974 0.120292
R29253 VDD.n3333 VDD.n3332 0.120292
R29254 VDD.n3334 VDD.n3333 0.120292
R29255 VDD.n3334 VDD.n2972 0.120292
R29256 VDD.n3340 VDD.n2972 0.120292
R29257 VDD.n3341 VDD.n3340 0.120292
R29258 VDD.n3341 VDD.n2968 0.120292
R29259 VDD.n3345 VDD.n2968 0.120292
R29260 VDD.n3346 VDD.n3345 0.120292
R29261 VDD.n3419 VDD.n3346 0.120292
R29262 VDD.n3419 VDD.n3418 0.120292
R29263 VDD.n3418 VDD.n3417 0.120292
R29264 VDD.n3417 VDD.n3347 0.120292
R29265 VDD.n3412 VDD.n3347 0.120292
R29266 VDD.n3412 VDD.n3411 0.120292
R29267 VDD.n3411 VDD.n3410 0.120292
R29268 VDD.n3410 VDD.n3351 0.120292
R29269 VDD.n3405 VDD.n3351 0.120292
R29270 VDD.n3405 VDD.n3404 0.120292
R29271 VDD.n3404 VDD.n3403 0.120292
R29272 VDD.n3403 VDD.n3355 0.120292
R29273 VDD.n3398 VDD.n3355 0.120292
R29274 VDD.n3398 VDD.n3397 0.120292
R29275 VDD.n3397 VDD.n3396 0.120292
R29276 VDD.n3396 VDD.n3358 0.120292
R29277 VDD.n3391 VDD.n3358 0.120292
R29278 VDD.n3391 VDD.n3390 0.120292
R29279 VDD.n3390 VDD.n3389 0.120292
R29280 VDD.n3389 VDD.n3360 0.120292
R29281 VDD.n3383 VDD.n3360 0.120292
R29282 VDD.n3383 VDD.n3382 0.120292
R29283 VDD.n3382 VDD.n3381 0.120292
R29284 VDD.n3381 VDD.n3364 0.120292
R29285 VDD.n3375 VDD.n3364 0.120292
R29286 VDD.n3375 VDD.n3374 0.120292
R29287 VDD.n3374 VDD.n3373 0.120292
R29288 VDD.n3373 VDD.n3367 0.120292
R29289 VDD.n3367 VDD.n2964 0.120292
R29290 VDD.n3427 VDD.n2964 0.120292
R29291 VDD.n3428 VDD.n3427 0.120292
R29292 VDD.n3428 VDD.n2962 0.120292
R29293 VDD.n2962 VDD.n2961 0.120292
R29294 VDD.n3435 VDD.n2961 0.120292
R29295 VDD.n3436 VDD.n3435 0.120292
R29296 VDD.n3437 VDD.n3436 0.120292
R29297 VDD.n3437 VDD.n2958 0.120292
R29298 VDD.n3443 VDD.n2958 0.120292
R29299 VDD.n3444 VDD.n3443 0.120292
R29300 VDD.n3445 VDD.n3444 0.120292
R29301 VDD.n3445 VDD.n2955 0.120292
R29302 VDD.n2955 VDD.n2954 0.120292
R29303 VDD.n2954 VDD.n2952 0.120292
R29304 VDD.n3452 VDD.n2952 0.120292
R29305 VDD.n3453 VDD.n3452 0.120292
R29306 VDD.n3454 VDD.n3453 0.120292
R29307 VDD.n3454 VDD.n2950 0.120292
R29308 VDD.n2950 VDD.n2948 0.120292
R29309 VDD.n3462 VDD.n2948 0.120292
R29310 VDD.n3463 VDD.n3462 0.120292
R29311 VDD.n3464 VDD.n3463 0.120292
R29312 VDD.n3464 VDD.n2945 0.120292
R29313 VDD.n3469 VDD.n2945 0.120292
R29314 VDD.n3470 VDD.n3469 0.120292
R29315 VDD.n3470 VDD.n2941 0.120292
R29316 VDD.n3476 VDD.n2941 0.120292
R29317 VDD.n3477 VDD.n3476 0.120292
R29318 VDD.n3478 VDD.n3477 0.120292
R29319 VDD.n3478 VDD.n2938 0.120292
R29320 VDD.n2938 VDD.n2937 0.120292
R29321 VDD.n3483 VDD.n2937 0.120292
R29322 VDD.n3484 VDD.n3483 0.120292
R29323 VDD.n3484 VDD.n2934 0.120292
R29324 VDD.n3489 VDD.n2934 0.120292
R29325 VDD.n3490 VDD.n3489 0.120292
R29326 VDD.n3491 VDD.n3490 0.120292
R29327 VDD.n3491 VDD.n2931 0.120292
R29328 VDD.n2931 VDD.n2930 0.120292
R29329 VDD.n3496 VDD.n2930 0.120292
R29330 VDD.n3497 VDD.n3496 0.120292
R29331 VDD.n3498 VDD.n3497 0.120292
R29332 VDD.n3505 VDD.n2921 0.120292
R29333 VDD.n3506 VDD.n3505 0.120292
R29334 VDD.n3506 VDD.n2918 0.120292
R29335 VDD.n3510 VDD.n2918 0.120292
R29336 VDD.n3511 VDD.n3510 0.120292
R29337 VDD.n3512 VDD.n3511 0.120292
R29338 VDD.n3512 VDD.n2914 0.120292
R29339 VDD.n3518 VDD.n2914 0.120292
R29340 VDD.n3519 VDD.n3518 0.120292
R29341 VDD.n3571 VDD.n3519 0.120292
R29342 VDD.n3571 VDD.n3570 0.120292
R29343 VDD.n3570 VDD.n3569 0.120292
R29344 VDD.n3569 VDD.n3520 0.120292
R29345 VDD.n3563 VDD.n3520 0.120292
R29346 VDD.n3563 VDD.n3562 0.120292
R29347 VDD.n3562 VDD.n3561 0.120292
R29348 VDD.n3561 VDD.n3524 0.120292
R29349 VDD.n3526 VDD.n3524 0.120292
R29350 VDD.n3556 VDD.n3526 0.120292
R29351 VDD.n3556 VDD.n3555 0.120292
R29352 VDD.n3555 VDD.n3528 0.120292
R29353 VDD.n3549 VDD.n3528 0.120292
R29354 VDD.n3549 VDD.n3548 0.120292
R29355 VDD.n3548 VDD.n3531 0.120292
R29356 VDD.n3533 VDD.n3531 0.120292
R29357 VDD.n3543 VDD.n3533 0.120292
R29358 VDD.n3543 VDD.n3542 0.120292
R29359 VDD.n3542 VDD.n3541 0.120292
R29360 VDD.n3541 VDD.n3535 0.120292
R29361 VDD.n3649 VDD.n3648 0.120292
R29362 VDD.n3648 VDD.n3647 0.120292
R29363 VDD.n3647 VDD.n2909 0.120292
R29364 VDD.n3641 VDD.n2909 0.120292
R29365 VDD.n3641 VDD.n3640 0.120292
R29366 VDD.n3640 VDD.n3639 0.120292
R29367 VDD.n3635 VDD.n3634 0.120292
R29368 VDD.n3634 VDD.n3584 0.120292
R29369 VDD.n3630 VDD.n3584 0.120292
R29370 VDD.n3630 VDD.n3629 0.120292
R29371 VDD.n3629 VDD.n3586 0.120292
R29372 VDD.n3625 VDD.n3586 0.120292
R29373 VDD.n3625 VDD.n3624 0.120292
R29374 VDD.n3624 VDD.n3623 0.120292
R29375 VDD.n3623 VDD.n3588 0.120292
R29376 VDD.n3619 VDD.n3588 0.120292
R29377 VDD.n3619 VDD.n3618 0.120292
R29378 VDD.n3618 VDD.n3590 0.120292
R29379 VDD.n3592 VDD.n3590 0.120292
R29380 VDD.n3613 VDD.n3592 0.120292
R29381 VDD.n3613 VDD.n3612 0.120292
R29382 VDD.n3612 VDD.n3611 0.120292
R29383 VDD.n3611 VDD.n3595 0.120292
R29384 VDD.n3607 VDD.n3595 0.120292
R29385 VDD.n2482 VDD.n2471 0.120292
R29386 VDD.n2471 VDD.n2469 0.120292
R29387 VDD.n2488 VDD.n2469 0.120292
R29388 VDD.n2489 VDD.n2488 0.120292
R29389 VDD.n2489 VDD.n2466 0.120292
R29390 VDD.n2466 VDD.n2465 0.120292
R29391 VDD.n2465 VDD.n2464 0.120292
R29392 VDD.n2464 VDD.n2463 0.120292
R29393 VDD.n2463 VDD.n2400 0.120292
R29394 VDD.n2402 VDD.n2400 0.120292
R29395 VDD.n2403 VDD.n2402 0.120292
R29396 VDD.n2404 VDD.n2403 0.120292
R29397 VDD.n2405 VDD.n2404 0.120292
R29398 VDD.n2454 VDD.n2405 0.120292
R29399 VDD.n2454 VDD.n2453 0.120292
R29400 VDD.n2453 VDD.n2408 0.120292
R29401 VDD.n2448 VDD.n2408 0.120292
R29402 VDD.n2448 VDD.n2447 0.120292
R29403 VDD.n2447 VDD.n2410 0.120292
R29404 VDD.n2443 VDD.n2410 0.120292
R29405 VDD.n2443 VDD.n2442 0.120292
R29406 VDD.n2442 VDD.n2412 0.120292
R29407 VDD.n2437 VDD.n2412 0.120292
R29408 VDD.n2437 VDD.n2436 0.120292
R29409 VDD.n2436 VDD.n2435 0.120292
R29410 VDD.n2435 VDD.n2414 0.120292
R29411 VDD.n2429 VDD.n2414 0.120292
R29412 VDD.n2429 VDD.n2428 0.120292
R29413 VDD.n2428 VDD.n2427 0.120292
R29414 VDD.n2427 VDD.n2417 0.120292
R29415 VDD.n2422 VDD.n2417 0.120292
R29416 VDD.n2422 VDD.n2421 0.120292
R29417 VDD.n2421 VDD.n2420 0.120292
R29418 VDD.n2420 VDD.n2397 0.120292
R29419 VDD.n2497 VDD.n2397 0.120292
R29420 VDD.n2505 VDD.n2395 0.120292
R29421 VDD.n2506 VDD.n2505 0.120292
R29422 VDD.n2506 VDD.n2392 0.120292
R29423 VDD.n2511 VDD.n2392 0.120292
R29424 VDD.n2512 VDD.n2511 0.120292
R29425 VDD.n2512 VDD.n2390 0.120292
R29426 VDD.n2517 VDD.n2390 0.120292
R29427 VDD.n2518 VDD.n2517 0.120292
R29428 VDD.n2518 VDD.n2388 0.120292
R29429 VDD.n2524 VDD.n2388 0.120292
R29430 VDD.n2525 VDD.n2524 0.120292
R29431 VDD.n2526 VDD.n2525 0.120292
R29432 VDD.n2526 VDD.n2384 0.120292
R29433 VDD.n2535 VDD.n2384 0.120292
R29434 VDD.n2536 VDD.n2535 0.120292
R29435 VDD.n2537 VDD.n2536 0.120292
R29436 VDD.n2537 VDD.n2381 0.120292
R29437 VDD.n2542 VDD.n2381 0.120292
R29438 VDD.n2543 VDD.n2542 0.120292
R29439 VDD.n2544 VDD.n2543 0.120292
R29440 VDD.n2544 VDD.n2379 0.120292
R29441 VDD.n2551 VDD.n2379 0.120292
R29442 VDD.n2552 VDD.n2551 0.120292
R29443 VDD.n2552 VDD.n2377 0.120292
R29444 VDD.n2561 VDD.n2560 0.120292
R29445 VDD.n2562 VDD.n2561 0.120292
R29446 VDD.n2562 VDD.n2364 0.120292
R29447 VDD.n2568 VDD.n2364 0.120292
R29448 VDD.n2569 VDD.n2568 0.120292
R29449 VDD.n2570 VDD.n2569 0.120292
R29450 VDD.n2570 VDD.n2360 0.120292
R29451 VDD.n2579 VDD.n2360 0.120292
R29452 VDD.n2580 VDD.n2579 0.120292
R29453 VDD.n2581 VDD.n2580 0.120292
R29454 VDD.n2353 VDD.n2352 0.120292
R29455 VDD.n2352 VDD.n2350 0.120292
R29456 VDD.n2588 VDD.n2350 0.120292
R29457 VDD.n2589 VDD.n2588 0.120292
R29458 VDD.n2590 VDD.n2589 0.120292
R29459 VDD.n2344 VDD.n2343 0.120292
R29460 VDD.n2343 VDD.n2342 0.120292
R29461 VDD.n2342 VDD.n2341 0.120292
R29462 VDD.n2341 VDD.n2338 0.120292
R29463 VDD.n2338 VDD.n2335 0.120292
R29464 VDD.n2602 VDD.n2335 0.120292
R29465 VDD.n2603 VDD.n2602 0.120292
R29466 VDD.n2603 VDD.n2333 0.120292
R29467 VDD.n2608 VDD.n2333 0.120292
R29468 VDD.n2609 VDD.n2608 0.120292
R29469 VDD.n2610 VDD.n2609 0.120292
R29470 VDD.n2610 VDD.n2330 0.120292
R29471 VDD.n2617 VDD.n2330 0.120292
R29472 VDD.n2618 VDD.n2617 0.120292
R29473 VDD.n2618 VDD.n2328 0.120292
R29474 VDD.n2623 VDD.n2328 0.120292
R29475 VDD.n2624 VDD.n2623 0.120292
R29476 VDD.n2624 VDD.n2325 0.120292
R29477 VDD.n2325 VDD.n2323 0.120292
R29478 VDD.n2323 VDD.n2322 0.120292
R29479 VDD.n2322 VDD.n2320 0.120292
R29480 VDD.n2631 VDD.n2320 0.120292
R29481 VDD.n2632 VDD.n2631 0.120292
R29482 VDD.n2632 VDD.n2317 0.120292
R29483 VDD.n2637 VDD.n2317 0.120292
R29484 VDD.n2638 VDD.n2637 0.120292
R29485 VDD.n2638 VDD.n2313 0.120292
R29486 VDD.n2313 VDD.n2312 0.120292
R29487 VDD.n2312 VDD.n2310 0.120292
R29488 VDD.n2310 VDD.n2309 0.120292
R29489 VDD.n2309 VDD.n2305 0.120292
R29490 VDD.n2652 VDD.n2305 0.120292
R29491 VDD.n2653 VDD.n2652 0.120292
R29492 VDD.n2654 VDD.n2653 0.120292
R29493 VDD.n2654 VDD.n2303 0.120292
R29494 VDD.n2662 VDD.n2303 0.120292
R29495 VDD.n2663 VDD.n2662 0.120292
R29496 VDD.n2664 VDD.n2663 0.120292
R29497 VDD.n2664 VDD.n2301 0.120292
R29498 VDD.n2669 VDD.n2301 0.120292
R29499 VDD.n2670 VDD.n2669 0.120292
R29500 VDD.n2670 VDD.n2298 0.120292
R29501 VDD.n2674 VDD.n2298 0.120292
R29502 VDD.n2675 VDD.n2674 0.120292
R29503 VDD.n2676 VDD.n2675 0.120292
R29504 VDD.n2676 VDD.n2295 0.120292
R29505 VDD.n2682 VDD.n2295 0.120292
R29506 VDD.n2683 VDD.n2682 0.120292
R29507 VDD.n2684 VDD.n2683 0.120292
R29508 VDD.n2684 VDD.n2292 0.120292
R29509 VDD.n2689 VDD.n2292 0.120292
R29510 VDD.n2690 VDD.n2689 0.120292
R29511 VDD.n2690 VDD.n2289 0.120292
R29512 VDD.n2695 VDD.n2289 0.120292
R29513 VDD.n2696 VDD.n2695 0.120292
R29514 VDD.n2696 VDD.n2286 0.120292
R29515 VDD.n2703 VDD.n2286 0.120292
R29516 VDD.n2704 VDD.n2703 0.120292
R29517 VDD.n2705 VDD.n2704 0.120292
R29518 VDD.n2705 VDD.n2283 0.120292
R29519 VDD.n2711 VDD.n2283 0.120292
R29520 VDD.n2712 VDD.n2711 0.120292
R29521 VDD.n2712 VDD.n2280 0.120292
R29522 VDD.n2717 VDD.n2280 0.120292
R29523 VDD.n2718 VDD.n2717 0.120292
R29524 VDD.n2718 VDD.n2276 0.120292
R29525 VDD.n2276 VDD.n2275 0.120292
R29526 VDD.n2725 VDD.n2275 0.120292
R29527 VDD.n2726 VDD.n2725 0.120292
R29528 VDD.n2727 VDD.n2726 0.120292
R29529 VDD.n2727 VDD.n2273 0.120292
R29530 VDD.n2734 VDD.n2273 0.120292
R29531 VDD.n2735 VDD.n2734 0.120292
R29532 VDD.n2736 VDD.n2735 0.120292
R29533 VDD.n2736 VDD.n2269 0.120292
R29534 VDD.n2742 VDD.n2269 0.120292
R29535 VDD.n2743 VDD.n2742 0.120292
R29536 VDD.n2744 VDD.n2743 0.120292
R29537 VDD.n2744 VDD.n2267 0.120292
R29538 VDD.n2749 VDD.n2267 0.120292
R29539 VDD.n2750 VDD.n2749 0.120292
R29540 VDD.n2751 VDD.n2750 0.120292
R29541 VDD.n2751 VDD.n2262 0.120292
R29542 VDD.n2757 VDD.n2262 0.120292
R29543 VDD.n2758 VDD.n2757 0.120292
R29544 VDD.n2759 VDD.n2758 0.120292
R29545 VDD.n2759 VDD.n2259 0.120292
R29546 VDD.n2767 VDD.n2259 0.120292
R29547 VDD.n2768 VDD.n2767 0.120292
R29548 VDD.n2768 VDD.n2257 0.120292
R29549 VDD.n2772 VDD.n2257 0.120292
R29550 VDD.n2773 VDD.n2772 0.120292
R29551 VDD.n2773 VDD.n2254 0.120292
R29552 VDD.n2254 VDD.n2253 0.120292
R29553 VDD.n2778 VDD.n2253 0.120292
R29554 VDD.n2779 VDD.n2778 0.120292
R29555 VDD.n2780 VDD.n2779 0.120292
R29556 VDD.n2780 VDD.n2249 0.120292
R29557 VDD.n2787 VDD.n2249 0.120292
R29558 VDD.n2788 VDD.n2787 0.120292
R29559 VDD.n2788 VDD.n2247 0.120292
R29560 VDD.n2794 VDD.n2247 0.120292
R29561 VDD.n2795 VDD.n2794 0.120292
R29562 VDD.n2796 VDD.n2795 0.120292
R29563 VDD.n2796 VDD.n2243 0.120292
R29564 VDD.n2802 VDD.n2243 0.120292
R29565 VDD.n2803 VDD.n2802 0.120292
R29566 VDD.n2803 VDD.n2239 0.120292
R29567 VDD.n2808 VDD.n2239 0.120292
R29568 VDD.n2809 VDD.n2808 0.120292
R29569 VDD.n2810 VDD.n2809 0.120292
R29570 VDD.n2810 VDD.n2236 0.120292
R29571 VDD.n2818 VDD.n2236 0.120292
R29572 VDD.n2819 VDD.n2818 0.120292
R29573 VDD.n2820 VDD.n2819 0.120292
R29574 VDD.n2820 VDD.n2234 0.120292
R29575 VDD.n2826 VDD.n2234 0.120292
R29576 VDD.n2827 VDD.n2826 0.120292
R29577 VDD.n2827 VDD.n2232 0.120292
R29578 VDD.n2833 VDD.n2232 0.120292
R29579 VDD.n2835 VDD.n2833 0.120292
R29580 VDD.n2844 VDD.n2843 0.120292
R29581 VDD.n2845 VDD.n2844 0.120292
R29582 VDD.n2845 VDD.n2222 0.120292
R29583 VDD.n2852 VDD.n2222 0.120292
R29584 VDD.n2853 VDD.n2852 0.120292
R29585 VDD.n2854 VDD.n2853 0.120292
R29586 VDD.n2854 VDD.n2219 0.120292
R29587 VDD.n2861 VDD.n2219 0.120292
R29588 VDD.n2862 VDD.n2861 0.120292
R29589 VDD.n2863 VDD.n2862 0.120292
R29590 VDD.n2863 VDD.n2217 0.120292
R29591 VDD.n2217 VDD.n2216 0.120292
R29592 VDD.n2216 VDD.n2215 0.120292
R29593 VDD.n2215 VDD.n2166 0.120292
R29594 VDD.n2210 VDD.n2166 0.120292
R29595 VDD.n2210 VDD.n2209 0.120292
R29596 VDD.n2209 VDD.n2208 0.120292
R29597 VDD.n2208 VDD.n2168 0.120292
R29598 VDD.n2202 VDD.n2168 0.120292
R29599 VDD.n2202 VDD.n2201 0.120292
R29600 VDD.n2201 VDD.n2200 0.120292
R29601 VDD.n2200 VDD.n2170 0.120292
R29602 VDD.n2195 VDD.n2170 0.120292
R29603 VDD.n2195 VDD.n2194 0.120292
R29604 VDD.n2194 VDD.n2193 0.120292
R29605 VDD.n2193 VDD.n2175 0.120292
R29606 VDD.n2188 VDD.n2175 0.120292
R29607 VDD.n2188 VDD.n2187 0.120292
R29608 VDD.n2187 VDD.n2178 0.120292
R29609 VDD.n2182 VDD.n2178 0.120292
R29610 VDD.n2877 VDD.n2876 0.120292
R29611 VDD.n2876 VDD.n2096 0.120292
R29612 VDD.n2871 VDD.n2096 0.120292
R29613 VDD.n2871 VDD.n2870 0.120292
R29614 VDD.n2870 VDD.n2100 0.120292
R29615 VDD.n2161 VDD.n2111 0.120292
R29616 VDD.n2154 VDD.n2111 0.120292
R29617 VDD.n2154 VDD.n2153 0.120292
R29618 VDD.n2153 VDD.n2152 0.120292
R29619 VDD.n2152 VDD.n2116 0.120292
R29620 VDD.n2117 VDD.n2116 0.120292
R29621 VDD.n2147 VDD.n2117 0.120292
R29622 VDD.n2147 VDD.n2146 0.120292
R29623 VDD.n2146 VDD.n2145 0.120292
R29624 VDD.n2145 VDD.n2119 0.120292
R29625 VDD.n2141 VDD.n2119 0.120292
R29626 VDD.n2141 VDD.n2140 0.120292
R29627 VDD.n2140 VDD.n2139 0.120292
R29628 VDD.n2139 VDD.n2123 0.120292
R29629 VDD.n2135 VDD.n2123 0.120292
R29630 VDD.n1664 VDD.n1653 0.120292
R29631 VDD.n1653 VDD.n1651 0.120292
R29632 VDD.n1670 VDD.n1651 0.120292
R29633 VDD.n1671 VDD.n1670 0.120292
R29634 VDD.n1671 VDD.n1648 0.120292
R29635 VDD.n1648 VDD.n1647 0.120292
R29636 VDD.n1647 VDD.n1646 0.120292
R29637 VDD.n1646 VDD.n1578 0.120292
R29638 VDD.n1641 VDD.n1578 0.120292
R29639 VDD.n1641 VDD.n1640 0.120292
R29640 VDD.n1640 VDD.n1639 0.120292
R29641 VDD.n1639 VDD.n1581 0.120292
R29642 VDD.n1634 VDD.n1581 0.120292
R29643 VDD.n1634 VDD.n1633 0.120292
R29644 VDD.n1633 VDD.n1583 0.120292
R29645 VDD.n1629 VDD.n1583 0.120292
R29646 VDD.n1629 VDD.n1628 0.120292
R29647 VDD.n1628 VDD.n1585 0.120292
R29648 VDD.n1622 VDD.n1585 0.120292
R29649 VDD.n1622 VDD.n1621 0.120292
R29650 VDD.n1621 VDD.n1587 0.120292
R29651 VDD.n1617 VDD.n1587 0.120292
R29652 VDD.n1617 VDD.n1616 0.120292
R29653 VDD.n1616 VDD.n1615 0.120292
R29654 VDD.n1615 VDD.n1589 0.120292
R29655 VDD.n1610 VDD.n1589 0.120292
R29656 VDD.n1610 VDD.n1609 0.120292
R29657 VDD.n1609 VDD.n1592 0.120292
R29658 VDD.n1603 VDD.n1592 0.120292
R29659 VDD.n1603 VDD.n1602 0.120292
R29660 VDD.n1602 VDD.n1601 0.120292
R29661 VDD.n1601 VDD.n1594 0.120292
R29662 VDD.n1594 VDD.n1575 0.120292
R29663 VDD.n1678 VDD.n1575 0.120292
R29664 VDD.n1688 VDD.n1573 0.120292
R29665 VDD.n1689 VDD.n1688 0.120292
R29666 VDD.n1689 VDD.n1569 0.120292
R29667 VDD.n1695 VDD.n1569 0.120292
R29668 VDD.n1696 VDD.n1695 0.120292
R29669 VDD.n1696 VDD.n1567 0.120292
R29670 VDD.n1704 VDD.n1567 0.120292
R29671 VDD.n1705 VDD.n1704 0.120292
R29672 VDD.n1706 VDD.n1705 0.120292
R29673 VDD.n1706 VDD.n1564 0.120292
R29674 VDD.n1710 VDD.n1564 0.120292
R29675 VDD.n1711 VDD.n1710 0.120292
R29676 VDD.n1712 VDD.n1711 0.120292
R29677 VDD.n1712 VDD.n1562 0.120292
R29678 VDD.n1720 VDD.n1562 0.120292
R29679 VDD.n1721 VDD.n1720 0.120292
R29680 VDD.n1722 VDD.n1721 0.120292
R29681 VDD.n1722 VDD.n1560 0.120292
R29682 VDD.n1726 VDD.n1560 0.120292
R29683 VDD.n1727 VDD.n1726 0.120292
R29684 VDD.n1728 VDD.n1727 0.120292
R29685 VDD.n1728 VDD.n1557 0.120292
R29686 VDD.n1733 VDD.n1557 0.120292
R29687 VDD.n1734 VDD.n1733 0.120292
R29688 VDD.n1735 VDD.n1734 0.120292
R29689 VDD.n1735 VDD.n1553 0.120292
R29690 VDD.n1740 VDD.n1553 0.120292
R29691 VDD.n1741 VDD.n1740 0.120292
R29692 VDD.n1742 VDD.n1741 0.120292
R29693 VDD.n1754 VDD.n1753 0.120292
R29694 VDD.n1755 VDD.n1754 0.120292
R29695 VDD.n1755 VDD.n1547 0.120292
R29696 VDD.n1762 VDD.n1547 0.120292
R29697 VDD.n1763 VDD.n1762 0.120292
R29698 VDD.n1763 VDD.n1544 0.120292
R29699 VDD.n1767 VDD.n1544 0.120292
R29700 VDD.n1768 VDD.n1767 0.120292
R29701 VDD.n1769 VDD.n1768 0.120292
R29702 VDD.n1769 VDD.n1541 0.120292
R29703 VDD.n1774 VDD.n1541 0.120292
R29704 VDD.n1775 VDD.n1774 0.120292
R29705 VDD.n1776 VDD.n1775 0.120292
R29706 VDD.n1776 VDD.n1538 0.120292
R29707 VDD.n1782 VDD.n1538 0.120292
R29708 VDD.n1783 VDD.n1782 0.120292
R29709 VDD.n1784 VDD.n1783 0.120292
R29710 VDD.n1784 VDD.n1536 0.120292
R29711 VDD.n1791 VDD.n1536 0.120292
R29712 VDD.n1792 VDD.n1791 0.120292
R29713 VDD.n1793 VDD.n1792 0.120292
R29714 VDD.n1793 VDD.n1532 0.120292
R29715 VDD.n1798 VDD.n1532 0.120292
R29716 VDD.n1799 VDD.n1798 0.120292
R29717 VDD.n1800 VDD.n1799 0.120292
R29718 VDD.n1800 VDD.n1530 0.120292
R29719 VDD.n1806 VDD.n1530 0.120292
R29720 VDD.n1807 VDD.n1806 0.120292
R29721 VDD.n1808 VDD.n1807 0.120292
R29722 VDD.n1808 VDD.n1527 0.120292
R29723 VDD.n1527 VDD.n1525 0.120292
R29724 VDD.n1813 VDD.n1525 0.120292
R29725 VDD.n1814 VDD.n1813 0.120292
R29726 VDD.n1815 VDD.n1814 0.120292
R29727 VDD.n1815 VDD.n1521 0.120292
R29728 VDD.n1821 VDD.n1521 0.120292
R29729 VDD.n1822 VDD.n1821 0.120292
R29730 VDD.n1822 VDD.n1519 0.120292
R29731 VDD.n1519 VDD.n1516 0.120292
R29732 VDD.n1829 VDD.n1516 0.120292
R29733 VDD.n1830 VDD.n1829 0.120292
R29734 VDD.n1830 VDD.n1512 0.120292
R29735 VDD.n1836 VDD.n1512 0.120292
R29736 VDD.n1837 VDD.n1836 0.120292
R29737 VDD.n1838 VDD.n1837 0.120292
R29738 VDD.n1838 VDD.n1510 0.120292
R29739 VDD.n1842 VDD.n1510 0.120292
R29740 VDD.n1843 VDD.n1842 0.120292
R29741 VDD.n1843 VDD.n1507 0.120292
R29742 VDD.n1851 VDD.n1507 0.120292
R29743 VDD.n1852 VDD.n1851 0.120292
R29744 VDD.n1853 VDD.n1852 0.120292
R29745 VDD.n1853 VDD.n1505 0.120292
R29746 VDD.n1858 VDD.n1505 0.120292
R29747 VDD.n1859 VDD.n1858 0.120292
R29748 VDD.n1860 VDD.n1859 0.120292
R29749 VDD.n1860 VDD.n1501 0.120292
R29750 VDD.n1864 VDD.n1501 0.120292
R29751 VDD.n1865 VDD.n1864 0.120292
R29752 VDD.n1866 VDD.n1865 0.120292
R29753 VDD.n1866 VDD.n1498 0.120292
R29754 VDD.n1870 VDD.n1498 0.120292
R29755 VDD.n1871 VDD.n1870 0.120292
R29756 VDD.n1872 VDD.n1871 0.120292
R29757 VDD.n1872 VDD.n1495 0.120292
R29758 VDD.n1495 VDD.n1493 0.120292
R29759 VDD.n1493 VDD.n1492 0.120292
R29760 VDD.n1492 VDD.n1490 0.120292
R29761 VDD.n1880 VDD.n1490 0.120292
R29762 VDD.n1881 VDD.n1880 0.120292
R29763 VDD.n1882 VDD.n1881 0.120292
R29764 VDD.n1882 VDD.n1485 0.120292
R29765 VDD.n1887 VDD.n1485 0.120292
R29766 VDD.n1888 VDD.n1887 0.120292
R29767 VDD.n1889 VDD.n1888 0.120292
R29768 VDD.n1889 VDD.n1478 0.120292
R29769 VDD.n1896 VDD.n1478 0.120292
R29770 VDD.n1897 VDD.n1896 0.120292
R29771 VDD.n1898 VDD.n1897 0.120292
R29772 VDD.n1898 VDD.n1475 0.120292
R29773 VDD.n1904 VDD.n1475 0.120292
R29774 VDD.n1905 VDD.n1904 0.120292
R29775 VDD.n1906 VDD.n1905 0.120292
R29776 VDD.n1906 VDD.n1472 0.120292
R29777 VDD.n1472 VDD.n1470 0.120292
R29778 VDD.n1914 VDD.n1470 0.120292
R29779 VDD.n1915 VDD.n1914 0.120292
R29780 VDD.n1915 VDD.n1467 0.120292
R29781 VDD.n1920 VDD.n1467 0.120292
R29782 VDD.n1921 VDD.n1920 0.120292
R29783 VDD.n1921 VDD.n1465 0.120292
R29784 VDD.n1926 VDD.n1465 0.120292
R29785 VDD.n1927 VDD.n1926 0.120292
R29786 VDD.n1927 VDD.n1462 0.120292
R29787 VDD.n1933 VDD.n1462 0.120292
R29788 VDD.n1934 VDD.n1933 0.120292
R29789 VDD.n1935 VDD.n1934 0.120292
R29790 VDD.n1935 VDD.n1459 0.120292
R29791 VDD.n1939 VDD.n1459 0.120292
R29792 VDD.n1940 VDD.n1939 0.120292
R29793 VDD.n1941 VDD.n1940 0.120292
R29794 VDD.n1941 VDD.n1456 0.120292
R29795 VDD.n1945 VDD.n1456 0.120292
R29796 VDD.n1947 VDD.n1450 0.120292
R29797 VDD.n1952 VDD.n1450 0.120292
R29798 VDD.n1953 VDD.n1952 0.120292
R29799 VDD.n1953 VDD.n1447 0.120292
R29800 VDD.n1959 VDD.n1447 0.120292
R29801 VDD.n1960 VDD.n1959 0.120292
R29802 VDD.n1960 VDD.n1444 0.120292
R29803 VDD.n1967 VDD.n1444 0.120292
R29804 VDD.n1968 VDD.n1967 0.120292
R29805 VDD.n1968 VDD.n1442 0.120292
R29806 VDD.n1972 VDD.n1442 0.120292
R29807 VDD.n1973 VDD.n1972 0.120292
R29808 VDD.n1974 VDD.n1973 0.120292
R29809 VDD.n1974 VDD.n1437 0.120292
R29810 VDD.n1980 VDD.n1437 0.120292
R29811 VDD.n1981 VDD.n1980 0.120292
R29812 VDD.n1982 VDD.n1981 0.120292
R29813 VDD.n1982 VDD.n1435 0.120292
R29814 VDD.n1435 VDD.n1433 0.120292
R29815 VDD.n1987 VDD.n1433 0.120292
R29816 VDD.n1988 VDD.n1987 0.120292
R29817 VDD.n1989 VDD.n1988 0.120292
R29818 VDD.n1989 VDD.n1430 0.120292
R29819 VDD.n1993 VDD.n1430 0.120292
R29820 VDD.n1994 VDD.n1993 0.120292
R29821 VDD.n1995 VDD.n1994 0.120292
R29822 VDD.n1995 VDD.n1427 0.120292
R29823 VDD.n2003 VDD.n1427 0.120292
R29824 VDD.n2004 VDD.n2003 0.120292
R29825 VDD.n2004 VDD.n1424 0.120292
R29826 VDD.n2011 VDD.n1424 0.120292
R29827 VDD.n2012 VDD.n2011 0.120292
R29828 VDD.n2012 VDD.n1421 0.120292
R29829 VDD.n2018 VDD.n1421 0.120292
R29830 VDD.n2019 VDD.n2018 0.120292
R29831 VDD.n2020 VDD.n2019 0.120292
R29832 VDD.n2020 VDD.n1418 0.120292
R29833 VDD.n2026 VDD.n1418 0.120292
R29834 VDD.n2027 VDD.n2026 0.120292
R29835 VDD.n2027 VDD.n1414 0.120292
R29836 VDD.n2033 VDD.n1414 0.120292
R29837 VDD.n2034 VDD.n2033 0.120292
R29838 VDD.n2034 VDD.n1412 0.120292
R29839 VDD.n2039 VDD.n1412 0.120292
R29840 VDD.n2040 VDD.n2039 0.120292
R29841 VDD.n2041 VDD.n2040 0.120292
R29842 VDD.n2041 VDD.n1407 0.120292
R29843 VDD.n2045 VDD.n1407 0.120292
R29844 VDD.n2046 VDD.n2045 0.120292
R29845 VDD.n2046 VDD.n1405 0.120292
R29846 VDD.n2054 VDD.n1405 0.120292
R29847 VDD.n2055 VDD.n2054 0.120292
R29848 VDD.n2055 VDD.n1403 0.120292
R29849 VDD.n1403 VDD.n1402 0.120292
R29850 VDD.n1402 VDD.n1401 0.120292
R29851 VDD.n1401 VDD.n1348 0.120292
R29852 VDD.n1396 VDD.n1348 0.120292
R29853 VDD.n1396 VDD.n1395 0.120292
R29854 VDD.n1395 VDD.n1394 0.120292
R29855 VDD.n1394 VDD.n1352 0.120292
R29856 VDD.n1388 VDD.n1352 0.120292
R29857 VDD.n1388 VDD.n1387 0.120292
R29858 VDD.n1387 VDD.n1386 0.120292
R29859 VDD.n1386 VDD.n1358 0.120292
R29860 VDD.n1381 VDD.n1358 0.120292
R29861 VDD.n1381 VDD.n1380 0.120292
R29862 VDD.n1380 VDD.n1361 0.120292
R29863 VDD.n1374 VDD.n1361 0.120292
R29864 VDD.n1374 VDD.n1373 0.120292
R29865 VDD.n1373 VDD.n1372 0.120292
R29866 VDD.n1372 VDD.n1365 0.120292
R29867 VDD.n1367 VDD.n1365 0.120292
R29868 VDD.n2071 VDD.n2070 0.120292
R29869 VDD.n2070 VDD.n1266 0.120292
R29870 VDD.n2063 VDD.n1266 0.120292
R29871 VDD.n2063 VDD.n2062 0.120292
R29872 VDD.n2062 VDD.n1269 0.120292
R29873 VDD.n1340 VDD.n1272 0.120292
R29874 VDD.n1334 VDD.n1272 0.120292
R29875 VDD.n1334 VDD.n1333 0.120292
R29876 VDD.n1333 VDD.n1332 0.120292
R29877 VDD.n1332 VDD.n1277 0.120292
R29878 VDD.n1327 VDD.n1277 0.120292
R29879 VDD.n1327 VDD.n1326 0.120292
R29880 VDD.n1326 VDD.n1280 0.120292
R29881 VDD.n1321 VDD.n1280 0.120292
R29882 VDD.n1321 VDD.n1320 0.120292
R29883 VDD.n1320 VDD.n1282 0.120292
R29884 VDD.n1283 VDD.n1282 0.120292
R29885 VDD.n1313 VDD.n1283 0.120292
R29886 VDD.n1313 VDD.n1312 0.120292
R29887 VDD.n1312 VDD.n1311 0.120292
R29888 VDD.n1311 VDD.n1285 0.120292
R29889 VDD.n1307 VDD.n1285 0.120292
R29890 VDD.n1307 VDD.n1306 0.120292
R29891 VDD.n1306 VDD.n1305 0.120292
R29892 VDD.n1305 VDD.n1289 0.120292
R29893 VDD.n1301 VDD.n1289 0.120292
R29894 VDD.n862 VDD.n861 0.120292
R29895 VDD.n862 VDD.n848 0.120292
R29896 VDD.n868 VDD.n848 0.120292
R29897 VDD.n869 VDD.n868 0.120292
R29898 VDD.n870 VDD.n869 0.120292
R29899 VDD.n870 VDD.n845 0.120292
R29900 VDD.n845 VDD.n844 0.120292
R29901 VDD.n844 VDD.n843 0.120292
R29902 VDD.n843 VDD.n842 0.120292
R29903 VDD.n842 VDD.n777 0.120292
R29904 VDD.n838 VDD.n777 0.120292
R29905 VDD.n838 VDD.n837 0.120292
R29906 VDD.n837 VDD.n836 0.120292
R29907 VDD.n836 VDD.n781 0.120292
R29908 VDD.n784 VDD.n781 0.120292
R29909 VDD.n831 VDD.n784 0.120292
R29910 VDD.n831 VDD.n830 0.120292
R29911 VDD.n830 VDD.n829 0.120292
R29912 VDD.n829 VDD.n787 0.120292
R29913 VDD.n788 VDD.n787 0.120292
R29914 VDD.n824 VDD.n788 0.120292
R29915 VDD.n824 VDD.n823 0.120292
R29916 VDD.n823 VDD.n822 0.120292
R29917 VDD.n822 VDD.n791 0.120292
R29918 VDD.n815 VDD.n791 0.120292
R29919 VDD.n815 VDD.n814 0.120292
R29920 VDD.n814 VDD.n813 0.120292
R29921 VDD.n813 VDD.n799 0.120292
R29922 VDD.n808 VDD.n799 0.120292
R29923 VDD.n808 VDD.n807 0.120292
R29924 VDD.n807 VDD.n803 0.120292
R29925 VDD.n775 VDD.n769 0.120292
R29926 VDD.n880 VDD.n769 0.120292
R29927 VDD.n881 VDD.n880 0.120292
R29928 VDD.n881 VDD.n766 0.120292
R29929 VDD.n766 VDD.n765 0.120292
R29930 VDD.n765 VDD.n764 0.120292
R29931 VDD.n764 VDD.n763 0.120292
R29932 VDD.n763 VDD.n760 0.120292
R29933 VDD.n889 VDD.n760 0.120292
R29934 VDD.n890 VDD.n889 0.120292
R29935 VDD.n891 VDD.n890 0.120292
R29936 VDD.n891 VDD.n757 0.120292
R29937 VDD.n757 VDD.n756 0.120292
R29938 VDD.n898 VDD.n756 0.120292
R29939 VDD.n899 VDD.n898 0.120292
R29940 VDD.n899 VDD.n753 0.120292
R29941 VDD.n903 VDD.n753 0.120292
R29942 VDD.n904 VDD.n903 0.120292
R29943 VDD.n905 VDD.n904 0.120292
R29944 VDD.n914 VDD.n748 0.120292
R29945 VDD.n915 VDD.n914 0.120292
R29946 VDD.n916 VDD.n915 0.120292
R29947 VDD.n916 VDD.n745 0.120292
R29948 VDD.n921 VDD.n745 0.120292
R29949 VDD.n922 VDD.n921 0.120292
R29950 VDD.n923 VDD.n922 0.120292
R29951 VDD.n923 VDD.n743 0.120292
R29952 VDD.n932 VDD.n743 0.120292
R29953 VDD.n933 VDD.n932 0.120292
R29954 VDD.n933 VDD.n741 0.120292
R29955 VDD.n940 VDD.n741 0.120292
R29956 VDD.n941 VDD.n940 0.120292
R29957 VDD.n941 VDD.n738 0.120292
R29958 VDD.n738 VDD.n736 0.120292
R29959 VDD.n946 VDD.n736 0.120292
R29960 VDD.n947 VDD.n946 0.120292
R29961 VDD.n948 VDD.n947 0.120292
R29962 VDD.n948 VDD.n734 0.120292
R29963 VDD.n958 VDD.n734 0.120292
R29964 VDD.n959 VDD.n958 0.120292
R29965 VDD.n960 VDD.n959 0.120292
R29966 VDD.n960 VDD.n731 0.120292
R29967 VDD.n964 VDD.n731 0.120292
R29968 VDD.n965 VDD.n964 0.120292
R29969 VDD.n966 VDD.n965 0.120292
R29970 VDD.n966 VDD.n729 0.120292
R29971 VDD.n975 VDD.n729 0.120292
R29972 VDD.n976 VDD.n975 0.120292
R29973 VDD.n977 VDD.n976 0.120292
R29974 VDD.n977 VDD.n726 0.120292
R29975 VDD.n726 VDD.n725 0.120292
R29976 VDD.n983 VDD.n725 0.120292
R29977 VDD.n984 VDD.n983 0.120292
R29978 VDD.n984 VDD.n722 0.120292
R29979 VDD.n996 VDD.n722 0.120292
R29980 VDD.n997 VDD.n996 0.120292
R29981 VDD.n998 VDD.n997 0.120292
R29982 VDD.n998 VDD.n720 0.120292
R29983 VDD.n1003 VDD.n720 0.120292
R29984 VDD.n1004 VDD.n1003 0.120292
R29985 VDD.n1004 VDD.n717 0.120292
R29986 VDD.n1010 VDD.n717 0.120292
R29987 VDD.n1011 VDD.n1010 0.120292
R29988 VDD.n1011 VDD.n715 0.120292
R29989 VDD.n1019 VDD.n715 0.120292
R29990 VDD.n1020 VDD.n1019 0.120292
R29991 VDD.n1021 VDD.n1020 0.120292
R29992 VDD.n1021 VDD.n713 0.120292
R29993 VDD.n1027 VDD.n713 0.120292
R29994 VDD.n1028 VDD.n1027 0.120292
R29995 VDD.n1028 VDD.n709 0.120292
R29996 VDD.n1034 VDD.n709 0.120292
R29997 VDD.n1035 VDD.n1034 0.120292
R29998 VDD.n1036 VDD.n1035 0.120292
R29999 VDD.n1036 VDD.n707 0.120292
R30000 VDD.n1041 VDD.n707 0.120292
R30001 VDD.n1042 VDD.n1041 0.120292
R30002 VDD.n1042 VDD.n704 0.120292
R30003 VDD.n1046 VDD.n704 0.120292
R30004 VDD.n1047 VDD.n1046 0.120292
R30005 VDD.n1047 VDD.n700 0.120292
R30006 VDD.n700 VDD.n699 0.120292
R30007 VDD.n1054 VDD.n699 0.120292
R30008 VDD.n1055 VDD.n1054 0.120292
R30009 VDD.n1055 VDD.n696 0.120292
R30010 VDD.n1061 VDD.n696 0.120292
R30011 VDD.n1062 VDD.n1061 0.120292
R30012 VDD.n1062 VDD.n692 0.120292
R30013 VDD.n1067 VDD.n692 0.120292
R30014 VDD.n1068 VDD.n1067 0.120292
R30015 VDD.n1069 VDD.n1068 0.120292
R30016 VDD.n1069 VDD.n689 0.120292
R30017 VDD.n1073 VDD.n689 0.120292
R30018 VDD.n1074 VDD.n1073 0.120292
R30019 VDD.n1075 VDD.n1074 0.120292
R30020 VDD.n1075 VDD.n686 0.120292
R30021 VDD.n1080 VDD.n686 0.120292
R30022 VDD.n1081 VDD.n1080 0.120292
R30023 VDD.n1082 VDD.n1081 0.120292
R30024 VDD.n1082 VDD.n684 0.120292
R30025 VDD.n684 VDD.n682 0.120292
R30026 VDD.n1087 VDD.n682 0.120292
R30027 VDD.n1088 VDD.n1087 0.120292
R30028 VDD.n1089 VDD.n1088 0.120292
R30029 VDD.n1089 VDD.n679 0.120292
R30030 VDD.n1093 VDD.n679 0.120292
R30031 VDD.n1094 VDD.n1093 0.120292
R30032 VDD.n1095 VDD.n1094 0.120292
R30033 VDD.n1095 VDD.n675 0.120292
R30034 VDD.n675 VDD.n674 0.120292
R30035 VDD.n1101 VDD.n674 0.120292
R30036 VDD.n1102 VDD.n1101 0.120292
R30037 VDD.n1103 VDD.n1102 0.120292
R30038 VDD.n1103 VDD.n670 0.120292
R30039 VDD.n1109 VDD.n670 0.120292
R30040 VDD.n1110 VDD.n1109 0.120292
R30041 VDD.n1111 VDD.n1110 0.120292
R30042 VDD.n1111 VDD.n668 0.120292
R30043 VDD.n1116 VDD.n668 0.120292
R30044 VDD.n1118 VDD.n1116 0.120292
R30045 VDD.n1118 VDD.n1117 0.120292
R30046 VDD.n1117 VDD.n663 0.120292
R30047 VDD.n1127 VDD.n663 0.120292
R30048 VDD.n1129 VDD.n656 0.120292
R30049 VDD.n1135 VDD.n656 0.120292
R30050 VDD.n1136 VDD.n1135 0.120292
R30051 VDD.n1137 VDD.n1136 0.120292
R30052 VDD.n1137 VDD.n653 0.120292
R30053 VDD.n653 VDD.n652 0.120292
R30054 VDD.n652 VDD.n651 0.120292
R30055 VDD.n644 VDD.n643 0.120292
R30056 VDD.n1148 VDD.n643 0.120292
R30057 VDD.n1149 VDD.n1148 0.120292
R30058 VDD.n1149 VDD.n641 0.120292
R30059 VDD.n641 VDD.n639 0.120292
R30060 VDD.n639 VDD.n631 0.120292
R30061 VDD.n1157 VDD.n624 0.120292
R30062 VDD.n1162 VDD.n624 0.120292
R30063 VDD.n1163 VDD.n1162 0.120292
R30064 VDD.n1163 VDD.n622 0.120292
R30065 VDD.n1169 VDD.n622 0.120292
R30066 VDD.n1170 VDD.n1169 0.120292
R30067 VDD.n1171 VDD.n1170 0.120292
R30068 VDD.n1171 VDD.n620 0.120292
R30069 VDD.n1178 VDD.n620 0.120292
R30070 VDD.n1179 VDD.n1178 0.120292
R30071 VDD.n1179 VDD.n617 0.120292
R30072 VDD.n1184 VDD.n617 0.120292
R30073 VDD.n1185 VDD.n1184 0.120292
R30074 VDD.n1185 VDD.n615 0.120292
R30075 VDD.n615 VDD.n612 0.120292
R30076 VDD.n1190 VDD.n612 0.120292
R30077 VDD.n1191 VDD.n1190 0.120292
R30078 VDD.n1192 VDD.n1191 0.120292
R30079 VDD.n1192 VDD.n609 0.120292
R30080 VDD.n1198 VDD.n609 0.120292
R30081 VDD.n1199 VDD.n1198 0.120292
R30082 VDD.n1199 VDD.n605 0.120292
R30083 VDD.n605 VDD.n604 0.120292
R30084 VDD.n1204 VDD.n604 0.120292
R30085 VDD.n1205 VDD.n1204 0.120292
R30086 VDD.n1206 VDD.n1205 0.120292
R30087 VDD.n1206 VDD.n602 0.120292
R30088 VDD.n602 VDD.n601 0.120292
R30089 VDD.n601 VDD.n599 0.120292
R30090 VDD.n1212 VDD.n599 0.120292
R30091 VDD.n1213 VDD.n1212 0.120292
R30092 VDD.n1214 VDD.n1213 0.120292
R30093 VDD.n1214 VDD.n596 0.120292
R30094 VDD.n1219 VDD.n596 0.120292
R30095 VDD.n1220 VDD.n1219 0.120292
R30096 VDD.n1221 VDD.n1220 0.120292
R30097 VDD.n1226 VDD.n1225 0.120292
R30098 VDD.n1227 VDD.n1226 0.120292
R30099 VDD.n1227 VDD.n587 0.120292
R30100 VDD.n587 VDD.n586 0.120292
R30101 VDD.n586 VDD.n585 0.120292
R30102 VDD.n585 VDD.n531 0.120292
R30103 VDD.n580 VDD.n531 0.120292
R30104 VDD.n580 VDD.n579 0.120292
R30105 VDD.n579 VDD.n536 0.120292
R30106 VDD.n574 VDD.n536 0.120292
R30107 VDD.n574 VDD.n573 0.120292
R30108 VDD.n573 VDD.n572 0.120292
R30109 VDD.n572 VDD.n540 0.120292
R30110 VDD.n568 VDD.n540 0.120292
R30111 VDD.n568 VDD.n567 0.120292
R30112 VDD.n567 VDD.n566 0.120292
R30113 VDD.n566 VDD.n542 0.120292
R30114 VDD.n560 VDD.n542 0.120292
R30115 VDD.n560 VDD.n559 0.120292
R30116 VDD.n559 VDD.n558 0.120292
R30117 VDD.n558 VDD.n549 0.120292
R30118 VDD.n553 VDD.n549 0.120292
R30119 VDD.n1241 VDD.n448 0.120292
R30120 VDD.n1236 VDD.n448 0.120292
R30121 VDD.n1236 VDD.n1235 0.120292
R30122 VDD.n1235 VDD.n1234 0.120292
R30123 VDD.n1234 VDD.n452 0.120292
R30124 VDD.n527 VDD.n452 0.120292
R30125 VDD.n525 VDD.n460 0.120292
R30126 VDD.n520 VDD.n460 0.120292
R30127 VDD.n520 VDD.n519 0.120292
R30128 VDD.n519 VDD.n518 0.120292
R30129 VDD.n518 VDD.n466 0.120292
R30130 VDD.n468 VDD.n466 0.120292
R30131 VDD.n513 VDD.n468 0.120292
R30132 VDD.n513 VDD.n512 0.120292
R30133 VDD.n512 VDD.n511 0.120292
R30134 VDD.n511 VDD.n471 0.120292
R30135 VDD.n507 VDD.n471 0.120292
R30136 VDD.n507 VDD.n506 0.120292
R30137 VDD.n506 VDD.n505 0.120292
R30138 VDD.n505 VDD.n475 0.120292
R30139 VDD.n501 VDD.n475 0.120292
R30140 VDD.n501 VDD.n500 0.120292
R30141 VDD.n500 VDD.n499 0.120292
R30142 VDD.n499 VDD.n479 0.120292
R30143 VDD.n493 VDD.n479 0.120292
R30144 VDD.n493 VDD.n492 0.120292
R30145 VDD.n419 VDD.n414 0.120292
R30146 VDD.n97 VDD.n96 0.120292
R30147 VDD.n97 VDD.n90 0.120292
R30148 VDD.n102 VDD.n90 0.120292
R30149 VDD.n61 VDD.n47 0.120292
R30150 VDD.n57 VDD.n47 0.120292
R30151 VDD.n18 VDD.n17 0.120292
R30152 VDD.n18 VDD.n10 0.120292
R30153 VDD.n65 VDD.n63 0.119731
R30154 VDD.n42 VDD.n41 0.119731
R30155 VDD.n2599 VDD.n2336 0.113774
R30156 VDD.n327 VDD.n326 0.111214
R30157 VDD.n400 VDD.n396 0.109875
R30158 VDD.n399 VDD.n398 0.109875
R30159 VDD.n139 VDD.n87 0.107397
R30160 VDD.n4151 VDD.n3714 0.106285
R30161 VDD.n3908 VDD.n3907 0.106285
R30162 VDD.n3937 VDD.n3936 0.106285
R30163 VDD.n4436 VDD.n4435 0.106285
R30164 VDD.n2513 VDD.n2391 0.106285
R30165 VDD.n2519 VDD.n2389 0.106285
R30166 VDD.n4232 VDD.n4231 0.102087
R30167 VDD.n4127 VDD.n3725 0.102087
R30168 VDD.n4260 VDD.n4259 0.102087
R30169 VDD.n4261 VDD.n3689 0.102087
R30170 VDD.n3248 VDD.n3247 0.102087
R30171 VDD.n3146 VDD.n3145 0.102087
R30172 VDD.n2785 VDD.n2784 0.102087
R30173 VDD.n2791 VDD.n2790 0.102087
R30174 VDD.n2547 VDD.n2546 0.102087
R30175 VDD.n2160 VDD.n2159 0.102087
R30176 VDD.n2157 VDD.n2156 0.102087
R30177 VDD.n2069 VDD.n2068 0.102087
R30178 VDD.n1158 VDD.n626 0.102087
R30179 VDD.n974 VDD.n973 0.102087
R30180 VDD.n821 VDD.n820 0.102087
R30181 VDD.n811 VDD.n810 0.102087
R30182 VDD.n402 VDD.n401 0.102062
R30183 VDD.n403 VDD.n395 0.102062
R30184 VDD.n4465 VDD.n4464 0.0950946
R30185 VDD.n4456 VDD.n4455 0.0950946
R30186 VDD.n3656 VDD.n3655 0.0950946
R30187 VDD.n2907 VDD.n2906 0.0950946
R30188 VDD.n2890 VDD.n2889 0.0950946
R30189 VDD.n2882 VDD.n2881 0.0950946
R30190 VDD.n2085 VDD.n2084 0.0950946
R30191 VDD.n2076 VDD.n2075 0.0950946
R30192 VDD.n1255 VDD.n1254 0.0950946
R30193 VDD.n1246 VDD.n1245 0.0950946
R30194 VDD.n62 VDD.n46 0.0890417
R30195 VDD.n26 VDD.n25 0.0877396
R30196 VDD.n3667 VDD.n3663 0.0838333
R30197 VDD.n2905 VDD.n2897 0.0838333
R30198 VDD.n2095 VDD.n2092 0.0838333
R30199 VDD.n1265 VDD.n1262 0.0838333
R30200 VDD.n447 VDD.n443 0.0838333
R30201 VDD.n4463 VDD.n4462 0.0812292
R30202 VDD.n3654 VDD.n3653 0.0812292
R30203 VDD.n2888 VDD.n2887 0.0812292
R30204 VDD.n2083 VDD.n2082 0.0812292
R30205 VDD.n1253 VDD.n1252 0.0812292
R30206 VDD.n4326 VDD.n3660 0.0760208
R30207 VDD.n3535 VDD.n2894 0.0760208
R30208 VDD.n2182 VDD.n2089 0.0760208
R30209 VDD.n1367 VDD.n1259 0.0760208
R30210 VDD.n553 VDD.n440 0.0760208
R30211 VDD.n431 VDD.n332 0.0759845
R30212 VDD.n45 VDD.n9 0.0712087
R30213 VDD.n4457 VDD.n4451 0.0708125
R30214 VDD.n3649 VDD.n2908 0.0708125
R30215 VDD.n2883 VDD.n2877 0.0708125
R30216 VDD.n2077 VDD.n2071 0.0708125
R30217 VDD.n1247 VDD.n1241 0.0708125
R30218 VDD.n4452 VDD.n3661 0.0680676
R30219 VDD.n4454 VDD.n4452 0.0680676
R30220 VDD.n2902 VDD.n2895 0.0680676
R30221 VDD.n2904 VDD.n2902 0.0680676
R30222 VDD.n2878 VDD.n2090 0.0680676
R30223 VDD.n2880 VDD.n2878 0.0680676
R30224 VDD.n2072 VDD.n1260 0.0680676
R30225 VDD.n2074 VDD.n2072 0.0680676
R30226 VDD.n1242 VDD.n441 0.0680676
R30227 VDD.n1244 VDD.n1242 0.0680676
R30228 VDD.n316 VDD.n223 0.0678077
R30229 VDD.n85 VDD.n82 0.0672614
R30230 VDD.n8 VDD.n5 0.0672614
R30231 VDD.n429 VDD.n428 0.0656042
R30232 VDD.n428 VDD.n413 0.0656042
R30233 VDD.n161 VDD.n160 0.063
R30234 VDD.n161 VDD.n102 0.0603958
R30235 VDD.n406 VDD.n404 0.0590938
R30236 VDD.n4453 VDD.n3659 0.0574697
R30237 VDD.n2903 VDD.n2893 0.0574697
R30238 VDD.n2879 VDD.n2088 0.0574697
R30239 VDD.n2073 VDD.n1258 0.0574697
R30240 VDD.n1243 VDD.n439 0.0574697
R30241 VDD.n407 VDD.n331 0.0557885
R30242 VDD.n435 VDD.n332 0.0557885
R30243 VDD.n429 VDD.n414 0.0551875
R30244 VDD.n4075 VDD.n3750 0.0512937
R30245 VDD.n3197 VDD.n3196 0.0512937
R30246 VDD.n804 VDD.n801 0.0512937
R30247 VDD.n4458 VDD.n4457 0.0499792
R30248 VDD.n2908 VDD.n2900 0.0499792
R30249 VDD.n2884 VDD.n2883 0.0499792
R30250 VDD.n2078 VDD.n2077 0.0499792
R30251 VDD.n1248 VDD.n1247 0.0499792
R30252 VDD.n3662 VDD.n3660 0.0447708
R30253 VDD.n2896 VDD.n2894 0.0447708
R30254 VDD.n2091 VDD.n2089 0.0447708
R30255 VDD.n1261 VDD.n1259 0.0447708
R30256 VDD.n442 VDD.n440 0.0447708
R30257 VDD.n151 VDD.n150 0.0435147
R30258 VDD.n176 VDD.n175 0.0435147
R30259 VDD.n436 VDD.n435 0.0419663
R30260 VDD.n4464 VDD.n3661 0.0410405
R30261 VDD.n4455 VDD.n4454 0.0410405
R30262 VDD.n3655 VDD.n2895 0.0410405
R30263 VDD.n2906 VDD.n2904 0.0410405
R30264 VDD.n2889 VDD.n2090 0.0410405
R30265 VDD.n2881 VDD.n2880 0.0410405
R30266 VDD.n2084 VDD.n1260 0.0410405
R30267 VDD.n2075 VDD.n2074 0.0410405
R30268 VDD.n1254 VDD.n441 0.0410405
R30269 VDD.n1245 VDD.n1244 0.0410405
R30270 VDD.n171 VDD.n170 0.0405735
R30271 VDD.n4463 VDD.n3662 0.0395625
R30272 VDD.n3654 VDD.n2896 0.0395625
R30273 VDD.n2888 VDD.n2091 0.0395625
R30274 VDD.n2083 VDD.n1261 0.0395625
R30275 VDD.n1253 VDD.n442 0.0395625
R30276 VDD.n4458 VDD.n3667 0.0343542
R30277 VDD.n2905 VDD.n2900 0.0343542
R30278 VDD.n2884 VDD.n2095 0.0343542
R30279 VDD.n2078 VDD.n1265 0.0343542
R30280 VDD.n1248 VDD.n447 0.0343542
R30281 VDD.n26 VDD.n10 0.0330521
R30282 VDD.n62 VDD.n61 0.03175
R30283 VDD.n1256 VDD.n439 0.0292489
R30284 VDD.n1243 VDD.n4 0.0292489
R30285 VDD.n2086 VDD.n1258 0.0292489
R30286 VDD.n2073 VDD.n3 0.0292489
R30287 VDD.n2891 VDD.n2088 0.0292489
R30288 VDD.n2879 VDD.n2 0.0292489
R30289 VDD.n3657 VDD.n2893 0.0292489
R30290 VDD.n2903 VDD.n1 0.0292489
R30291 VDD.n4466 VDD.n3659 0.0292489
R30292 VDD.n4453 VDD.n0 0.0292489
R30293 VDD.n436 VDD.n331 0.0143221
R30294 VDD.n238 VDD.n181 0.00530769
R30295 VDD.n4462 VDD.n3663 0.00310417
R30296 VDD.n3653 VDD.n2897 0.00310417
R30297 VDD.n2887 VDD.n2092 0.00310417
R30298 VDD.n2082 VDD.n1262 0.00310417
R30299 VDD.n1252 VDD.n443 0.00310417
R30300 C10_P_btm C10_P_btm.n32 92.1047
R30301 C10_P_btm.n2 C10_P_btm.n0 33.0802
R30302 C10_P_btm.n14 C10_P_btm.n13 32.3614
R30303 C10_P_btm.n12 C10_P_btm.n11 32.3614
R30304 C10_P_btm.n10 C10_P_btm.n9 32.3614
R30305 C10_P_btm.n8 C10_P_btm.n7 32.3614
R30306 C10_P_btm.n6 C10_P_btm.n5 32.3614
R30307 C10_P_btm.n4 C10_P_btm.n3 32.3614
R30308 C10_P_btm.n2 C10_P_btm.n1 32.3614
R30309 C10_P_btm.n22 C10_P_btm.n14 29.1203
R30310 C10_P_btm.n24 C10_P_btm.n23 20.3263
R30311 C10_P_btm.n28 C10_P_btm.n26 15.4755
R30312 C10_P_btm.n17 C10_P_btm.n15 15.394
R30313 C10_P_btm.n31 C10_P_btm.n25 14.9755
R30314 C10_P_btm.n28 C10_P_btm.n27 14.9755
R30315 C10_P_btm.n30 C10_P_btm.n29 14.9755
R30316 C10_P_btm.n21 C10_P_btm.n20 14.894
R30317 C10_P_btm.n19 C10_P_btm.n18 14.894
R30318 C10_P_btm.n17 C10_P_btm.n16 14.894
R30319 C10_P_btm C10_P_btm.n3897 6.338
R30320 C10_P_btm.n24 C10_P_btm.n22 6.29217
R30321 C10_P_btm.n22 C10_P_btm.n21 5.43279
R30322 C10_P_btm.n32 C10_P_btm.n31 5.33904
R30323 C10_P_btm.n34 C10_P_btm.t19 5.03712
R30324 C10_P_btm.n35 C10_P_btm.t24 5.03712
R30325 C10_P_btm.n36 C10_P_btm.t21 5.03712
R30326 C10_P_btm.n37 C10_P_btm.t13 5.03712
R30327 C10_P_btm.n38 C10_P_btm.t14 5.03712
R30328 C10_P_btm.n39 C10_P_btm.t20 5.03712
R30329 C10_P_btm.n40 C10_P_btm.t25 5.03712
R30330 C10_P_btm.n41 C10_P_btm.t16 5.03712
R30331 C10_P_btm.n42 C10_P_btm.t23 5.03712
R30332 C10_P_btm.n3866 C10_P_btm.t30 5.03712
R30333 C10_P_btm.n2413 C10_P_btm.t10 5.03712
R30334 C10_P_btm.n2429 C10_P_btm.t11 5.03712
R30335 C10_P_btm.n2428 C10_P_btm.t15 5.03712
R30336 C10_P_btm.n2427 C10_P_btm.t18 5.03712
R30337 C10_P_btm.n2426 C10_P_btm.t31 5.03712
R30338 C10_P_btm.n2425 C10_P_btm.t26 5.03712
R30339 C10_P_btm.n2424 C10_P_btm.t22 5.03712
R30340 C10_P_btm.n2423 C10_P_btm.t28 5.03712
R30341 C10_P_btm.n2422 C10_P_btm.t12 5.03712
R30342 C10_P_btm.n2460 C10_P_btm.t27 5.03712
R30343 C10_P_btm.n2456 C10_P_btm.t29 5.03712
R30344 C10_P_btm.n32 C10_P_btm.n24 4.7505
R30345 C10_P_btm.n3894 C10_P_btm.n3893 4.60698
R30346 C10_P_btm.n3893 C10_P_btm.n3892 4.60698
R30347 C10_P_btm.n3891 C10_P_btm.n3890 4.60698
R30348 C10_P_btm.n3890 C10_P_btm.n3889 4.60698
R30349 C10_P_btm.n3888 C10_P_btm.n3887 4.60698
R30350 C10_P_btm.n3887 C10_P_btm.n3886 4.60698
R30351 C10_P_btm.n3885 C10_P_btm.n3884 4.60698
R30352 C10_P_btm.n3884 C10_P_btm.n3883 4.60698
R30353 C10_P_btm.n3882 C10_P_btm.n3881 4.60698
R30354 C10_P_btm.n3881 C10_P_btm.n3880 4.60698
R30355 C10_P_btm.n3879 C10_P_btm.n3878 4.60698
R30356 C10_P_btm.n3878 C10_P_btm.n3877 4.60698
R30357 C10_P_btm.n3876 C10_P_btm.n3875 4.60698
R30358 C10_P_btm.n3875 C10_P_btm.n3874 4.60698
R30359 C10_P_btm.n3873 C10_P_btm.n3872 4.60698
R30360 C10_P_btm.n3872 C10_P_btm.n3871 4.60698
R30361 C10_P_btm.n3870 C10_P_btm.n3869 4.60698
R30362 C10_P_btm.n3869 C10_P_btm.n3868 4.60698
R30363 C10_P_btm.n3863 C10_P_btm.n3862 4.60698
R30364 C10_P_btm.n3862 C10_P_btm.n3861 4.60698
R30365 C10_P_btm.n3860 C10_P_btm.n3859 4.60698
R30366 C10_P_btm.n3859 C10_P_btm.n3858 4.60698
R30367 C10_P_btm.n3857 C10_P_btm.n3856 4.60698
R30368 C10_P_btm.n3856 C10_P_btm.n3855 4.60698
R30369 C10_P_btm.n3854 C10_P_btm.n3853 4.60698
R30370 C10_P_btm.n3853 C10_P_btm.n3852 4.60698
R30371 C10_P_btm.n3851 C10_P_btm.n3850 4.60698
R30372 C10_P_btm.n3850 C10_P_btm.n3849 4.60698
R30373 C10_P_btm.n3848 C10_P_btm.n3847 4.60698
R30374 C10_P_btm.n3847 C10_P_btm.n3846 4.60698
R30375 C10_P_btm.n3845 C10_P_btm.n3844 4.60698
R30376 C10_P_btm.n3844 C10_P_btm.n3843 4.60698
R30377 C10_P_btm.n3842 C10_P_btm.n3841 4.60698
R30378 C10_P_btm.n3841 C10_P_btm.n3840 4.60698
R30379 C10_P_btm.n3839 C10_P_btm.n3838 4.60698
R30380 C10_P_btm.n3838 C10_P_btm.n3837 4.60698
R30381 C10_P_btm.n3833 C10_P_btm.n3832 4.60698
R30382 C10_P_btm.n3832 C10_P_btm.n53 4.60698
R30383 C10_P_btm.n3830 C10_P_btm.n3829 4.60698
R30384 C10_P_btm.n3831 C10_P_btm.n3830 4.60698
R30385 C10_P_btm.n3827 C10_P_btm.n3826 4.60698
R30386 C10_P_btm.n3828 C10_P_btm.n3827 4.60698
R30387 C10_P_btm.n3824 C10_P_btm.n3823 4.60698
R30388 C10_P_btm.n3825 C10_P_btm.n3824 4.60698
R30389 C10_P_btm.n3821 C10_P_btm.n3820 4.60698
R30390 C10_P_btm.n3822 C10_P_btm.n3821 4.60698
R30391 C10_P_btm.n3818 C10_P_btm.n3817 4.60698
R30392 C10_P_btm.n3819 C10_P_btm.n3818 4.60698
R30393 C10_P_btm.n3815 C10_P_btm.n3814 4.60698
R30394 C10_P_btm.n3816 C10_P_btm.n3815 4.60698
R30395 C10_P_btm.n3812 C10_P_btm.n3811 4.60698
R30396 C10_P_btm.n3813 C10_P_btm.n3812 4.60698
R30397 C10_P_btm.n3809 C10_P_btm.n3808 4.60698
R30398 C10_P_btm.n3810 C10_P_btm.n3809 4.60698
R30399 C10_P_btm.n3804 C10_P_btm.n3803 4.60698
R30400 C10_P_btm.n3803 C10_P_btm.n62 4.60698
R30401 C10_P_btm.n3745 C10_P_btm.n3744 4.60698
R30402 C10_P_btm.n3746 C10_P_btm.n3745 4.60698
R30403 C10_P_btm.n3748 C10_P_btm.n3747 4.60698
R30404 C10_P_btm.n3749 C10_P_btm.n3748 4.60698
R30405 C10_P_btm.n3751 C10_P_btm.n3750 4.60698
R30406 C10_P_btm.n3752 C10_P_btm.n3751 4.60698
R30407 C10_P_btm.n3754 C10_P_btm.n3753 4.60698
R30408 C10_P_btm.n3755 C10_P_btm.n3754 4.60698
R30409 C10_P_btm.n3757 C10_P_btm.n3756 4.60698
R30410 C10_P_btm.n3758 C10_P_btm.n3757 4.60698
R30411 C10_P_btm.n3760 C10_P_btm.n3759 4.60698
R30412 C10_P_btm.n3761 C10_P_btm.n3760 4.60698
R30413 C10_P_btm.n3763 C10_P_btm.n3762 4.60698
R30414 C10_P_btm.n3764 C10_P_btm.n3763 4.60698
R30415 C10_P_btm.n3766 C10_P_btm.n3765 4.60698
R30416 C10_P_btm.n3767 C10_P_btm.n3766 4.60698
R30417 C10_P_btm.n3774 C10_P_btm.n3773 4.60698
R30418 C10_P_btm.n3773 C10_P_btm.n3772 4.60698
R30419 C10_P_btm.n3777 C10_P_btm.n3776 4.60698
R30420 C10_P_btm.n3776 C10_P_btm.n3775 4.60698
R30421 C10_P_btm.n3780 C10_P_btm.n3779 4.60698
R30422 C10_P_btm.n3779 C10_P_btm.n3778 4.60698
R30423 C10_P_btm.n3783 C10_P_btm.n3782 4.60698
R30424 C10_P_btm.n3782 C10_P_btm.n3781 4.60698
R30425 C10_P_btm.n3786 C10_P_btm.n3785 4.60698
R30426 C10_P_btm.n3785 C10_P_btm.n3784 4.60698
R30427 C10_P_btm.n3789 C10_P_btm.n3788 4.60698
R30428 C10_P_btm.n3788 C10_P_btm.n3787 4.60698
R30429 C10_P_btm.n3792 C10_P_btm.n3791 4.60698
R30430 C10_P_btm.n3791 C10_P_btm.n3790 4.60698
R30431 C10_P_btm.n3795 C10_P_btm.n3794 4.60698
R30432 C10_P_btm.n3794 C10_P_btm.n3793 4.60698
R30433 C10_P_btm.n3798 C10_P_btm.n3797 4.60698
R30434 C10_P_btm.n3797 C10_P_btm.n3796 4.60698
R30435 C10_P_btm.n3707 C10_P_btm.n3706 4.60698
R30436 C10_P_btm.n3708 C10_P_btm.n3707 4.60698
R30437 C10_P_btm.n3710 C10_P_btm.n3709 4.60698
R30438 C10_P_btm.n3711 C10_P_btm.n3710 4.60698
R30439 C10_P_btm.n3713 C10_P_btm.n3712 4.60698
R30440 C10_P_btm.n3714 C10_P_btm.n3713 4.60698
R30441 C10_P_btm.n3716 C10_P_btm.n3715 4.60698
R30442 C10_P_btm.n3717 C10_P_btm.n3716 4.60698
R30443 C10_P_btm.n3719 C10_P_btm.n3718 4.60698
R30444 C10_P_btm.n3720 C10_P_btm.n3719 4.60698
R30445 C10_P_btm.n3722 C10_P_btm.n3721 4.60698
R30446 C10_P_btm.n3723 C10_P_btm.n3722 4.60698
R30447 C10_P_btm.n3725 C10_P_btm.n3724 4.60698
R30448 C10_P_btm.n3726 C10_P_btm.n3725 4.60698
R30449 C10_P_btm.n3728 C10_P_btm.n3727 4.60698
R30450 C10_P_btm.n3729 C10_P_btm.n3728 4.60698
R30451 C10_P_btm.n3731 C10_P_btm.n3730 4.60698
R30452 C10_P_btm.n3732 C10_P_btm.n3731 4.60698
R30453 C10_P_btm.n122 C10_P_btm.n121 4.60698
R30454 C10_P_btm.n121 C10_P_btm.n92 4.60698
R30455 C10_P_btm.n119 C10_P_btm.n118 4.60698
R30456 C10_P_btm.n120 C10_P_btm.n119 4.60698
R30457 C10_P_btm.n116 C10_P_btm.n115 4.60698
R30458 C10_P_btm.n117 C10_P_btm.n116 4.60698
R30459 C10_P_btm.n113 C10_P_btm.n112 4.60698
R30460 C10_P_btm.n114 C10_P_btm.n113 4.60698
R30461 C10_P_btm.n110 C10_P_btm.n109 4.60698
R30462 C10_P_btm.n111 C10_P_btm.n110 4.60698
R30463 C10_P_btm.n107 C10_P_btm.n106 4.60698
R30464 C10_P_btm.n108 C10_P_btm.n107 4.60698
R30465 C10_P_btm.n104 C10_P_btm.n103 4.60698
R30466 C10_P_btm.n105 C10_P_btm.n104 4.60698
R30467 C10_P_btm.n101 C10_P_btm.n100 4.60698
R30468 C10_P_btm.n102 C10_P_btm.n101 4.60698
R30469 C10_P_btm.n3702 C10_P_btm.n3701 4.60698
R30470 C10_P_btm.n3701 C10_P_btm.n82 4.60698
R30471 C10_P_btm.n3696 C10_P_btm.n3695 4.60698
R30472 C10_P_btm.n3695 C10_P_btm.n3694 4.60698
R30473 C10_P_btm.n3693 C10_P_btm.n3692 4.60698
R30474 C10_P_btm.n3692 C10_P_btm.n3691 4.60698
R30475 C10_P_btm.n3690 C10_P_btm.n3689 4.60698
R30476 C10_P_btm.n3689 C10_P_btm.n3688 4.60698
R30477 C10_P_btm.n3687 C10_P_btm.n3686 4.60698
R30478 C10_P_btm.n3686 C10_P_btm.n3685 4.60698
R30479 C10_P_btm.n3684 C10_P_btm.n3683 4.60698
R30480 C10_P_btm.n3683 C10_P_btm.n3682 4.60698
R30481 C10_P_btm.n3681 C10_P_btm.n3680 4.60698
R30482 C10_P_btm.n3680 C10_P_btm.n3679 4.60698
R30483 C10_P_btm.n3678 C10_P_btm.n3677 4.60698
R30484 C10_P_btm.n3677 C10_P_btm.n3676 4.60698
R30485 C10_P_btm.n3675 C10_P_btm.n3674 4.60698
R30486 C10_P_btm.n3674 C10_P_btm.n3673 4.60698
R30487 C10_P_btm.n3672 C10_P_btm.n3671 4.60698
R30488 C10_P_btm.n3671 C10_P_btm.n3670 4.60698
R30489 C10_P_btm.n3664 C10_P_btm.n3663 4.60698
R30490 C10_P_btm.n3665 C10_P_btm.n3664 4.60698
R30491 C10_P_btm.n3661 C10_P_btm.n3660 4.60698
R30492 C10_P_btm.n3662 C10_P_btm.n3661 4.60698
R30493 C10_P_btm.n3658 C10_P_btm.n3657 4.60698
R30494 C10_P_btm.n3659 C10_P_btm.n3658 4.60698
R30495 C10_P_btm.n3655 C10_P_btm.n3654 4.60698
R30496 C10_P_btm.n3656 C10_P_btm.n3655 4.60698
R30497 C10_P_btm.n3652 C10_P_btm.n3651 4.60698
R30498 C10_P_btm.n3653 C10_P_btm.n3652 4.60698
R30499 C10_P_btm.n3649 C10_P_btm.n3648 4.60698
R30500 C10_P_btm.n3650 C10_P_btm.n3649 4.60698
R30501 C10_P_btm.n3646 C10_P_btm.n3645 4.60698
R30502 C10_P_btm.n3647 C10_P_btm.n3646 4.60698
R30503 C10_P_btm.n3643 C10_P_btm.n3642 4.60698
R30504 C10_P_btm.n3644 C10_P_btm.n3643 4.60698
R30505 C10_P_btm.n3640 C10_P_btm.n3639 4.60698
R30506 C10_P_btm.n3641 C10_P_btm.n3640 4.60698
R30507 C10_P_btm.n3635 C10_P_btm.n3634 4.60698
R30508 C10_P_btm.n3634 C10_P_btm.n135 4.60698
R30509 C10_P_btm.n154 C10_P_btm.n153 4.60698
R30510 C10_P_btm.n155 C10_P_btm.n154 4.60698
R30511 C10_P_btm.n157 C10_P_btm.n156 4.60698
R30512 C10_P_btm.n158 C10_P_btm.n157 4.60698
R30513 C10_P_btm.n160 C10_P_btm.n159 4.60698
R30514 C10_P_btm.n161 C10_P_btm.n160 4.60698
R30515 C10_P_btm.n163 C10_P_btm.n162 4.60698
R30516 C10_P_btm.n164 C10_P_btm.n163 4.60698
R30517 C10_P_btm.n166 C10_P_btm.n165 4.60698
R30518 C10_P_btm.n167 C10_P_btm.n166 4.60698
R30519 C10_P_btm.n169 C10_P_btm.n168 4.60698
R30520 C10_P_btm.n170 C10_P_btm.n169 4.60698
R30521 C10_P_btm.n172 C10_P_btm.n171 4.60698
R30522 C10_P_btm.n173 C10_P_btm.n172 4.60698
R30523 C10_P_btm.n175 C10_P_btm.n174 4.60698
R30524 C10_P_btm.n174 C10_P_btm.n145 4.60698
R30525 C10_P_btm.n3605 C10_P_btm.n3604 4.60698
R30526 C10_P_btm.n3604 C10_P_btm.n3603 4.60698
R30527 C10_P_btm.n3608 C10_P_btm.n3607 4.60698
R30528 C10_P_btm.n3607 C10_P_btm.n3606 4.60698
R30529 C10_P_btm.n3611 C10_P_btm.n3610 4.60698
R30530 C10_P_btm.n3610 C10_P_btm.n3609 4.60698
R30531 C10_P_btm.n3614 C10_P_btm.n3613 4.60698
R30532 C10_P_btm.n3613 C10_P_btm.n3612 4.60698
R30533 C10_P_btm.n3617 C10_P_btm.n3616 4.60698
R30534 C10_P_btm.n3616 C10_P_btm.n3615 4.60698
R30535 C10_P_btm.n3620 C10_P_btm.n3619 4.60698
R30536 C10_P_btm.n3619 C10_P_btm.n3618 4.60698
R30537 C10_P_btm.n3623 C10_P_btm.n3622 4.60698
R30538 C10_P_btm.n3622 C10_P_btm.n3621 4.60698
R30539 C10_P_btm.n3626 C10_P_btm.n3625 4.60698
R30540 C10_P_btm.n3625 C10_P_btm.n3624 4.60698
R30541 C10_P_btm.n3629 C10_P_btm.n3628 4.60698
R30542 C10_P_btm.n3628 C10_P_btm.n3627 4.60698
R30543 C10_P_btm.n3573 C10_P_btm.n3572 4.60698
R30544 C10_P_btm.n3574 C10_P_btm.n3573 4.60698
R30545 C10_P_btm.n3576 C10_P_btm.n3575 4.60698
R30546 C10_P_btm.n3577 C10_P_btm.n3576 4.60698
R30547 C10_P_btm.n3579 C10_P_btm.n3578 4.60698
R30548 C10_P_btm.n3580 C10_P_btm.n3579 4.60698
R30549 C10_P_btm.n3582 C10_P_btm.n3581 4.60698
R30550 C10_P_btm.n3583 C10_P_btm.n3582 4.60698
R30551 C10_P_btm.n3585 C10_P_btm.n3584 4.60698
R30552 C10_P_btm.n3586 C10_P_btm.n3585 4.60698
R30553 C10_P_btm.n3588 C10_P_btm.n3587 4.60698
R30554 C10_P_btm.n3589 C10_P_btm.n3588 4.60698
R30555 C10_P_btm.n3591 C10_P_btm.n3590 4.60698
R30556 C10_P_btm.n3592 C10_P_btm.n3591 4.60698
R30557 C10_P_btm.n3594 C10_P_btm.n3593 4.60698
R30558 C10_P_btm.n3595 C10_P_btm.n3594 4.60698
R30559 C10_P_btm.n3597 C10_P_btm.n3596 4.60698
R30560 C10_P_btm.n3598 C10_P_btm.n3597 4.60698
R30561 C10_P_btm.n228 C10_P_btm.n227 4.60698
R30562 C10_P_btm.n227 C10_P_btm.n198 4.60698
R30563 C10_P_btm.n225 C10_P_btm.n224 4.60698
R30564 C10_P_btm.n226 C10_P_btm.n225 4.60698
R30565 C10_P_btm.n222 C10_P_btm.n221 4.60698
R30566 C10_P_btm.n223 C10_P_btm.n222 4.60698
R30567 C10_P_btm.n219 C10_P_btm.n218 4.60698
R30568 C10_P_btm.n220 C10_P_btm.n219 4.60698
R30569 C10_P_btm.n216 C10_P_btm.n215 4.60698
R30570 C10_P_btm.n217 C10_P_btm.n216 4.60698
R30571 C10_P_btm.n213 C10_P_btm.n212 4.60698
R30572 C10_P_btm.n214 C10_P_btm.n213 4.60698
R30573 C10_P_btm.n210 C10_P_btm.n209 4.60698
R30574 C10_P_btm.n211 C10_P_btm.n210 4.60698
R30575 C10_P_btm.n207 C10_P_btm.n206 4.60698
R30576 C10_P_btm.n208 C10_P_btm.n207 4.60698
R30577 C10_P_btm.n3568 C10_P_btm.n3567 4.60698
R30578 C10_P_btm.n3567 C10_P_btm.n188 4.60698
R30579 C10_P_btm.n3562 C10_P_btm.n3561 4.60698
R30580 C10_P_btm.n3561 C10_P_btm.n3560 4.60698
R30581 C10_P_btm.n3559 C10_P_btm.n3558 4.60698
R30582 C10_P_btm.n3558 C10_P_btm.n3557 4.60698
R30583 C10_P_btm.n3556 C10_P_btm.n3555 4.60698
R30584 C10_P_btm.n3555 C10_P_btm.n3554 4.60698
R30585 C10_P_btm.n3553 C10_P_btm.n3552 4.60698
R30586 C10_P_btm.n3552 C10_P_btm.n3551 4.60698
R30587 C10_P_btm.n3550 C10_P_btm.n3549 4.60698
R30588 C10_P_btm.n3549 C10_P_btm.n3548 4.60698
R30589 C10_P_btm.n3547 C10_P_btm.n3546 4.60698
R30590 C10_P_btm.n3546 C10_P_btm.n3545 4.60698
R30591 C10_P_btm.n3544 C10_P_btm.n3543 4.60698
R30592 C10_P_btm.n3543 C10_P_btm.n3542 4.60698
R30593 C10_P_btm.n3541 C10_P_btm.n3540 4.60698
R30594 C10_P_btm.n3540 C10_P_btm.n3539 4.60698
R30595 C10_P_btm.n3538 C10_P_btm.n3537 4.60698
R30596 C10_P_btm.n3537 C10_P_btm.n3536 4.60698
R30597 C10_P_btm.n3530 C10_P_btm.n3529 4.60698
R30598 C10_P_btm.n3531 C10_P_btm.n3530 4.60698
R30599 C10_P_btm.n3527 C10_P_btm.n3526 4.60698
R30600 C10_P_btm.n3528 C10_P_btm.n3527 4.60698
R30601 C10_P_btm.n3524 C10_P_btm.n3523 4.60698
R30602 C10_P_btm.n3525 C10_P_btm.n3524 4.60698
R30603 C10_P_btm.n3521 C10_P_btm.n3520 4.60698
R30604 C10_P_btm.n3522 C10_P_btm.n3521 4.60698
R30605 C10_P_btm.n3518 C10_P_btm.n3517 4.60698
R30606 C10_P_btm.n3519 C10_P_btm.n3518 4.60698
R30607 C10_P_btm.n3515 C10_P_btm.n3514 4.60698
R30608 C10_P_btm.n3516 C10_P_btm.n3515 4.60698
R30609 C10_P_btm.n3512 C10_P_btm.n3511 4.60698
R30610 C10_P_btm.n3513 C10_P_btm.n3512 4.60698
R30611 C10_P_btm.n3509 C10_P_btm.n3508 4.60698
R30612 C10_P_btm.n3510 C10_P_btm.n3509 4.60698
R30613 C10_P_btm.n3506 C10_P_btm.n3505 4.60698
R30614 C10_P_btm.n3507 C10_P_btm.n3506 4.60698
R30615 C10_P_btm.n3501 C10_P_btm.n3500 4.60698
R30616 C10_P_btm.n3500 C10_P_btm.n241 4.60698
R30617 C10_P_btm.n260 C10_P_btm.n259 4.60698
R30618 C10_P_btm.n261 C10_P_btm.n260 4.60698
R30619 C10_P_btm.n263 C10_P_btm.n262 4.60698
R30620 C10_P_btm.n264 C10_P_btm.n263 4.60698
R30621 C10_P_btm.n266 C10_P_btm.n265 4.60698
R30622 C10_P_btm.n267 C10_P_btm.n266 4.60698
R30623 C10_P_btm.n269 C10_P_btm.n268 4.60698
R30624 C10_P_btm.n270 C10_P_btm.n269 4.60698
R30625 C10_P_btm.n272 C10_P_btm.n271 4.60698
R30626 C10_P_btm.n273 C10_P_btm.n272 4.60698
R30627 C10_P_btm.n275 C10_P_btm.n274 4.60698
R30628 C10_P_btm.n276 C10_P_btm.n275 4.60698
R30629 C10_P_btm.n278 C10_P_btm.n277 4.60698
R30630 C10_P_btm.n279 C10_P_btm.n278 4.60698
R30631 C10_P_btm.n281 C10_P_btm.n280 4.60698
R30632 C10_P_btm.n280 C10_P_btm.n251 4.60698
R30633 C10_P_btm.n3471 C10_P_btm.n3470 4.60698
R30634 C10_P_btm.n3470 C10_P_btm.n3469 4.60698
R30635 C10_P_btm.n3474 C10_P_btm.n3473 4.60698
R30636 C10_P_btm.n3473 C10_P_btm.n3472 4.60698
R30637 C10_P_btm.n3477 C10_P_btm.n3476 4.60698
R30638 C10_P_btm.n3476 C10_P_btm.n3475 4.60698
R30639 C10_P_btm.n3480 C10_P_btm.n3479 4.60698
R30640 C10_P_btm.n3479 C10_P_btm.n3478 4.60698
R30641 C10_P_btm.n3483 C10_P_btm.n3482 4.60698
R30642 C10_P_btm.n3482 C10_P_btm.n3481 4.60698
R30643 C10_P_btm.n3486 C10_P_btm.n3485 4.60698
R30644 C10_P_btm.n3485 C10_P_btm.n3484 4.60698
R30645 C10_P_btm.n3489 C10_P_btm.n3488 4.60698
R30646 C10_P_btm.n3488 C10_P_btm.n3487 4.60698
R30647 C10_P_btm.n3492 C10_P_btm.n3491 4.60698
R30648 C10_P_btm.n3491 C10_P_btm.n3490 4.60698
R30649 C10_P_btm.n3495 C10_P_btm.n3494 4.60698
R30650 C10_P_btm.n3494 C10_P_btm.n3493 4.60698
R30651 C10_P_btm.n3439 C10_P_btm.n3438 4.60698
R30652 C10_P_btm.n3440 C10_P_btm.n3439 4.60698
R30653 C10_P_btm.n3442 C10_P_btm.n3441 4.60698
R30654 C10_P_btm.n3443 C10_P_btm.n3442 4.60698
R30655 C10_P_btm.n3445 C10_P_btm.n3444 4.60698
R30656 C10_P_btm.n3446 C10_P_btm.n3445 4.60698
R30657 C10_P_btm.n3448 C10_P_btm.n3447 4.60698
R30658 C10_P_btm.n3449 C10_P_btm.n3448 4.60698
R30659 C10_P_btm.n3451 C10_P_btm.n3450 4.60698
R30660 C10_P_btm.n3452 C10_P_btm.n3451 4.60698
R30661 C10_P_btm.n3454 C10_P_btm.n3453 4.60698
R30662 C10_P_btm.n3455 C10_P_btm.n3454 4.60698
R30663 C10_P_btm.n3457 C10_P_btm.n3456 4.60698
R30664 C10_P_btm.n3458 C10_P_btm.n3457 4.60698
R30665 C10_P_btm.n3460 C10_P_btm.n3459 4.60698
R30666 C10_P_btm.n3461 C10_P_btm.n3460 4.60698
R30667 C10_P_btm.n3463 C10_P_btm.n3462 4.60698
R30668 C10_P_btm.n3464 C10_P_btm.n3463 4.60698
R30669 C10_P_btm.n334 C10_P_btm.n333 4.60698
R30670 C10_P_btm.n333 C10_P_btm.n304 4.60698
R30671 C10_P_btm.n331 C10_P_btm.n330 4.60698
R30672 C10_P_btm.n332 C10_P_btm.n331 4.60698
R30673 C10_P_btm.n328 C10_P_btm.n327 4.60698
R30674 C10_P_btm.n329 C10_P_btm.n328 4.60698
R30675 C10_P_btm.n325 C10_P_btm.n324 4.60698
R30676 C10_P_btm.n326 C10_P_btm.n325 4.60698
R30677 C10_P_btm.n322 C10_P_btm.n321 4.60698
R30678 C10_P_btm.n323 C10_P_btm.n322 4.60698
R30679 C10_P_btm.n319 C10_P_btm.n318 4.60698
R30680 C10_P_btm.n320 C10_P_btm.n319 4.60698
R30681 C10_P_btm.n316 C10_P_btm.n315 4.60698
R30682 C10_P_btm.n317 C10_P_btm.n316 4.60698
R30683 C10_P_btm.n313 C10_P_btm.n312 4.60698
R30684 C10_P_btm.n314 C10_P_btm.n313 4.60698
R30685 C10_P_btm.n3434 C10_P_btm.n3433 4.60698
R30686 C10_P_btm.n3433 C10_P_btm.n294 4.60698
R30687 C10_P_btm.n3428 C10_P_btm.n3427 4.60698
R30688 C10_P_btm.n3427 C10_P_btm.n3426 4.60698
R30689 C10_P_btm.n3425 C10_P_btm.n3424 4.60698
R30690 C10_P_btm.n3424 C10_P_btm.n3423 4.60698
R30691 C10_P_btm.n3422 C10_P_btm.n3421 4.60698
R30692 C10_P_btm.n3421 C10_P_btm.n3420 4.60698
R30693 C10_P_btm.n3419 C10_P_btm.n3418 4.60698
R30694 C10_P_btm.n3418 C10_P_btm.n3417 4.60698
R30695 C10_P_btm.n3416 C10_P_btm.n3415 4.60698
R30696 C10_P_btm.n3415 C10_P_btm.n3414 4.60698
R30697 C10_P_btm.n3413 C10_P_btm.n3412 4.60698
R30698 C10_P_btm.n3412 C10_P_btm.n3411 4.60698
R30699 C10_P_btm.n3410 C10_P_btm.n3409 4.60698
R30700 C10_P_btm.n3409 C10_P_btm.n3408 4.60698
R30701 C10_P_btm.n3407 C10_P_btm.n3406 4.60698
R30702 C10_P_btm.n3406 C10_P_btm.n3405 4.60698
R30703 C10_P_btm.n3404 C10_P_btm.n3403 4.60698
R30704 C10_P_btm.n3403 C10_P_btm.n3402 4.60698
R30705 C10_P_btm.n3396 C10_P_btm.n3395 4.60698
R30706 C10_P_btm.n3397 C10_P_btm.n3396 4.60698
R30707 C10_P_btm.n3393 C10_P_btm.n3392 4.60698
R30708 C10_P_btm.n3394 C10_P_btm.n3393 4.60698
R30709 C10_P_btm.n3390 C10_P_btm.n3389 4.60698
R30710 C10_P_btm.n3391 C10_P_btm.n3390 4.60698
R30711 C10_P_btm.n3387 C10_P_btm.n3386 4.60698
R30712 C10_P_btm.n3388 C10_P_btm.n3387 4.60698
R30713 C10_P_btm.n3384 C10_P_btm.n3383 4.60698
R30714 C10_P_btm.n3385 C10_P_btm.n3384 4.60698
R30715 C10_P_btm.n3381 C10_P_btm.n3380 4.60698
R30716 C10_P_btm.n3382 C10_P_btm.n3381 4.60698
R30717 C10_P_btm.n3378 C10_P_btm.n3377 4.60698
R30718 C10_P_btm.n3379 C10_P_btm.n3378 4.60698
R30719 C10_P_btm.n3375 C10_P_btm.n3374 4.60698
R30720 C10_P_btm.n3376 C10_P_btm.n3375 4.60698
R30721 C10_P_btm.n3372 C10_P_btm.n3371 4.60698
R30722 C10_P_btm.n3373 C10_P_btm.n3372 4.60698
R30723 C10_P_btm.n3367 C10_P_btm.n3366 4.60698
R30724 C10_P_btm.n3366 C10_P_btm.n347 4.60698
R30725 C10_P_btm.n366 C10_P_btm.n365 4.60698
R30726 C10_P_btm.n367 C10_P_btm.n366 4.60698
R30727 C10_P_btm.n369 C10_P_btm.n368 4.60698
R30728 C10_P_btm.n370 C10_P_btm.n369 4.60698
R30729 C10_P_btm.n372 C10_P_btm.n371 4.60698
R30730 C10_P_btm.n373 C10_P_btm.n372 4.60698
R30731 C10_P_btm.n375 C10_P_btm.n374 4.60698
R30732 C10_P_btm.n376 C10_P_btm.n375 4.60698
R30733 C10_P_btm.n378 C10_P_btm.n377 4.60698
R30734 C10_P_btm.n379 C10_P_btm.n378 4.60698
R30735 C10_P_btm.n381 C10_P_btm.n380 4.60698
R30736 C10_P_btm.n382 C10_P_btm.n381 4.60698
R30737 C10_P_btm.n384 C10_P_btm.n383 4.60698
R30738 C10_P_btm.n385 C10_P_btm.n384 4.60698
R30739 C10_P_btm.n387 C10_P_btm.n386 4.60698
R30740 C10_P_btm.n386 C10_P_btm.n357 4.60698
R30741 C10_P_btm.n3337 C10_P_btm.n3336 4.60698
R30742 C10_P_btm.n3336 C10_P_btm.n3335 4.60698
R30743 C10_P_btm.n3340 C10_P_btm.n3339 4.60698
R30744 C10_P_btm.n3339 C10_P_btm.n3338 4.60698
R30745 C10_P_btm.n3343 C10_P_btm.n3342 4.60698
R30746 C10_P_btm.n3342 C10_P_btm.n3341 4.60698
R30747 C10_P_btm.n3346 C10_P_btm.n3345 4.60698
R30748 C10_P_btm.n3345 C10_P_btm.n3344 4.60698
R30749 C10_P_btm.n3349 C10_P_btm.n3348 4.60698
R30750 C10_P_btm.n3348 C10_P_btm.n3347 4.60698
R30751 C10_P_btm.n3352 C10_P_btm.n3351 4.60698
R30752 C10_P_btm.n3351 C10_P_btm.n3350 4.60698
R30753 C10_P_btm.n3355 C10_P_btm.n3354 4.60698
R30754 C10_P_btm.n3354 C10_P_btm.n3353 4.60698
R30755 C10_P_btm.n3358 C10_P_btm.n3357 4.60698
R30756 C10_P_btm.n3357 C10_P_btm.n3356 4.60698
R30757 C10_P_btm.n3361 C10_P_btm.n3360 4.60698
R30758 C10_P_btm.n3360 C10_P_btm.n3359 4.60698
R30759 C10_P_btm.n3305 C10_P_btm.n3304 4.60698
R30760 C10_P_btm.n3306 C10_P_btm.n3305 4.60698
R30761 C10_P_btm.n3308 C10_P_btm.n3307 4.60698
R30762 C10_P_btm.n3309 C10_P_btm.n3308 4.60698
R30763 C10_P_btm.n3311 C10_P_btm.n3310 4.60698
R30764 C10_P_btm.n3312 C10_P_btm.n3311 4.60698
R30765 C10_P_btm.n3314 C10_P_btm.n3313 4.60698
R30766 C10_P_btm.n3315 C10_P_btm.n3314 4.60698
R30767 C10_P_btm.n3317 C10_P_btm.n3316 4.60698
R30768 C10_P_btm.n3318 C10_P_btm.n3317 4.60698
R30769 C10_P_btm.n3320 C10_P_btm.n3319 4.60698
R30770 C10_P_btm.n3321 C10_P_btm.n3320 4.60698
R30771 C10_P_btm.n3323 C10_P_btm.n3322 4.60698
R30772 C10_P_btm.n3324 C10_P_btm.n3323 4.60698
R30773 C10_P_btm.n3326 C10_P_btm.n3325 4.60698
R30774 C10_P_btm.n3327 C10_P_btm.n3326 4.60698
R30775 C10_P_btm.n3329 C10_P_btm.n3328 4.60698
R30776 C10_P_btm.n3330 C10_P_btm.n3329 4.60698
R30777 C10_P_btm.n469 C10_P_btm.n468 4.60698
R30778 C10_P_btm.n468 C10_P_btm.n467 4.60698
R30779 C10_P_btm.n465 C10_P_btm.n464 4.60698
R30780 C10_P_btm.n466 C10_P_btm.n465 4.60698
R30781 C10_P_btm.n462 C10_P_btm.n461 4.60698
R30782 C10_P_btm.n463 C10_P_btm.n462 4.60698
R30783 C10_P_btm.n459 C10_P_btm.n458 4.60698
R30784 C10_P_btm.n460 C10_P_btm.n459 4.60698
R30785 C10_P_btm.n456 C10_P_btm.n455 4.60698
R30786 C10_P_btm.n457 C10_P_btm.n456 4.60698
R30787 C10_P_btm.n453 C10_P_btm.n452 4.60698
R30788 C10_P_btm.n454 C10_P_btm.n453 4.60698
R30789 C10_P_btm.n450 C10_P_btm.n449 4.60698
R30790 C10_P_btm.n451 C10_P_btm.n450 4.60698
R30791 C10_P_btm.n447 C10_P_btm.n446 4.60698
R30792 C10_P_btm.n448 C10_P_btm.n447 4.60698
R30793 C10_P_btm.n444 C10_P_btm.n443 4.60698
R30794 C10_P_btm.n445 C10_P_btm.n444 4.60698
R30795 C10_P_btm.n3300 C10_P_btm.n3299 4.60698
R30796 C10_P_btm.n3299 C10_P_btm.n400 4.60698
R30797 C10_P_btm.n3294 C10_P_btm.n3293 4.60698
R30798 C10_P_btm.n3293 C10_P_btm.n3292 4.60698
R30799 C10_P_btm.n3291 C10_P_btm.n3290 4.60698
R30800 C10_P_btm.n3290 C10_P_btm.n3289 4.60698
R30801 C10_P_btm.n3288 C10_P_btm.n3287 4.60698
R30802 C10_P_btm.n3287 C10_P_btm.n3286 4.60698
R30803 C10_P_btm.n3285 C10_P_btm.n3284 4.60698
R30804 C10_P_btm.n3284 C10_P_btm.n3283 4.60698
R30805 C10_P_btm.n3282 C10_P_btm.n3281 4.60698
R30806 C10_P_btm.n3281 C10_P_btm.n3280 4.60698
R30807 C10_P_btm.n3279 C10_P_btm.n3278 4.60698
R30808 C10_P_btm.n3278 C10_P_btm.n3277 4.60698
R30809 C10_P_btm.n3276 C10_P_btm.n3275 4.60698
R30810 C10_P_btm.n3275 C10_P_btm.n3274 4.60698
R30811 C10_P_btm.n3273 C10_P_btm.n3272 4.60698
R30812 C10_P_btm.n3272 C10_P_btm.n3271 4.60698
R30813 C10_P_btm.n3270 C10_P_btm.n3269 4.60698
R30814 C10_P_btm.n3269 C10_P_btm.n3268 4.60698
R30815 C10_P_btm.n3267 C10_P_btm.n3266 4.60698
R30816 C10_P_btm.n3266 C10_P_btm.n3265 4.60698
R30817 C10_P_btm.n3264 C10_P_btm.n3263 4.60698
R30818 C10_P_btm.n3263 C10_P_btm.n3262 4.60698
R30819 C10_P_btm.n3261 C10_P_btm.n3260 4.60698
R30820 C10_P_btm.n3260 C10_P_btm.n3259 4.60698
R30821 C10_P_btm.n3258 C10_P_btm.n3257 4.60698
R30822 C10_P_btm.n3257 C10_P_btm.n3256 4.60698
R30823 C10_P_btm.n3255 C10_P_btm.n3254 4.60698
R30824 C10_P_btm.n3254 C10_P_btm.n3253 4.60698
R30825 C10_P_btm.n3252 C10_P_btm.n3251 4.60698
R30826 C10_P_btm.n3251 C10_P_btm.n3250 4.60698
R30827 C10_P_btm.n3249 C10_P_btm.n3248 4.60698
R30828 C10_P_btm.n3248 C10_P_btm.n3247 4.60698
R30829 C10_P_btm.n3246 C10_P_btm.n3245 4.60698
R30830 C10_P_btm.n3245 C10_P_btm.n3244 4.60698
R30831 C10_P_btm.n3243 C10_P_btm.n3242 4.60698
R30832 C10_P_btm.n3242 C10_P_btm.n3241 4.60698
R30833 C10_P_btm.n3240 C10_P_btm.n3239 4.60698
R30834 C10_P_btm.n3239 C10_P_btm.n3238 4.60698
R30835 C10_P_btm.n3237 C10_P_btm.n3236 4.60698
R30836 C10_P_btm.n3236 C10_P_btm.n3235 4.60698
R30837 C10_P_btm.n3234 C10_P_btm.n3233 4.60698
R30838 C10_P_btm.n3233 C10_P_btm.n3232 4.60698
R30839 C10_P_btm.n3231 C10_P_btm.n3230 4.60698
R30840 C10_P_btm.n3230 C10_P_btm.n3229 4.60698
R30841 C10_P_btm.n3227 C10_P_btm.n3226 4.60698
R30842 C10_P_btm.n3228 C10_P_btm.n3227 4.60698
R30843 C10_P_btm.n505 C10_P_btm.n504 4.60698
R30844 C10_P_btm.n504 C10_P_btm.n503 4.60698
R30845 C10_P_btm.n502 C10_P_btm.n501 4.60698
R30846 C10_P_btm.n501 C10_P_btm.n500 4.60698
R30847 C10_P_btm.n499 C10_P_btm.n498 4.60698
R30848 C10_P_btm.n498 C10_P_btm.n497 4.60698
R30849 C10_P_btm.n496 C10_P_btm.n495 4.60698
R30850 C10_P_btm.n495 C10_P_btm.n494 4.60698
R30851 C10_P_btm.n493 C10_P_btm.n492 4.60698
R30852 C10_P_btm.n492 C10_P_btm.n491 4.60698
R30853 C10_P_btm.n490 C10_P_btm.n489 4.60698
R30854 C10_P_btm.n489 C10_P_btm.n488 4.60698
R30855 C10_P_btm.n487 C10_P_btm.n486 4.60698
R30856 C10_P_btm.n486 C10_P_btm.n485 4.60698
R30857 C10_P_btm.n484 C10_P_btm.n483 4.60698
R30858 C10_P_btm.n483 C10_P_btm.n482 4.60698
R30859 C10_P_btm.n481 C10_P_btm.n480 4.60698
R30860 C10_P_btm.n480 C10_P_btm.n479 4.60698
R30861 C10_P_btm.n478 C10_P_btm.n477 4.60698
R30862 C10_P_btm.n477 C10_P_btm.n476 4.60698
R30863 C10_P_btm.n475 C10_P_btm.n474 4.60698
R30864 C10_P_btm.n474 C10_P_btm.n473 4.60698
R30865 C10_P_btm.n472 C10_P_btm.n471 4.60698
R30866 C10_P_btm.n471 C10_P_btm.n470 4.60698
R30867 C10_P_btm.n3224 C10_P_btm.n3223 4.60698
R30868 C10_P_btm.n3225 C10_P_btm.n3224 4.60698
R30869 C10_P_btm.n3221 C10_P_btm.n3220 4.60698
R30870 C10_P_btm.n3222 C10_P_btm.n3221 4.60698
R30871 C10_P_btm.n3218 C10_P_btm.n3217 4.60698
R30872 C10_P_btm.n3219 C10_P_btm.n3218 4.60698
R30873 C10_P_btm.n3215 C10_P_btm.n3214 4.60698
R30874 C10_P_btm.n3216 C10_P_btm.n3215 4.60698
R30875 C10_P_btm.n3212 C10_P_btm.n3211 4.60698
R30876 C10_P_btm.n3213 C10_P_btm.n3212 4.60698
R30877 C10_P_btm.n3209 C10_P_btm.n3208 4.60698
R30878 C10_P_btm.n3210 C10_P_btm.n3209 4.60698
R30879 C10_P_btm.n3206 C10_P_btm.n3205 4.60698
R30880 C10_P_btm.n3207 C10_P_btm.n3206 4.60698
R30881 C10_P_btm.n3203 C10_P_btm.n3202 4.60698
R30882 C10_P_btm.n3204 C10_P_btm.n3203 4.60698
R30883 C10_P_btm.n3200 C10_P_btm.n3199 4.60698
R30884 C10_P_btm.n3201 C10_P_btm.n3200 4.60698
R30885 C10_P_btm.n3197 C10_P_btm.n3196 4.60698
R30886 C10_P_btm.n3198 C10_P_btm.n3197 4.60698
R30887 C10_P_btm.n3194 C10_P_btm.n3193 4.60698
R30888 C10_P_btm.n3195 C10_P_btm.n3194 4.60698
R30889 C10_P_btm.n3191 C10_P_btm.n3190 4.60698
R30890 C10_P_btm.n3192 C10_P_btm.n3191 4.60698
R30891 C10_P_btm.n3188 C10_P_btm.n3187 4.60698
R30892 C10_P_btm.n3189 C10_P_btm.n3188 4.60698
R30893 C10_P_btm.n3185 C10_P_btm.n3184 4.60698
R30894 C10_P_btm.n3186 C10_P_btm.n3185 4.60698
R30895 C10_P_btm.n3182 C10_P_btm.n3181 4.60698
R30896 C10_P_btm.n3183 C10_P_btm.n3182 4.60698
R30897 C10_P_btm.n3179 C10_P_btm.n3178 4.60698
R30898 C10_P_btm.n3180 C10_P_btm.n3179 4.60698
R30899 C10_P_btm.n3177 C10_P_btm.n3176 4.60698
R30900 C10_P_btm.n3176 C10_P_btm.n3175 4.60698
R30901 C10_P_btm.n3174 C10_P_btm.n3173 4.60698
R30902 C10_P_btm.n3173 C10_P_btm.n3172 4.60698
R30903 C10_P_btm.n3171 C10_P_btm.n3170 4.60698
R30904 C10_P_btm.n3170 C10_P_btm.n3169 4.60698
R30905 C10_P_btm.n3168 C10_P_btm.n3167 4.60698
R30906 C10_P_btm.n3167 C10_P_btm.n3166 4.60698
R30907 C10_P_btm.n3165 C10_P_btm.n3164 4.60698
R30908 C10_P_btm.n3164 C10_P_btm.n3163 4.60698
R30909 C10_P_btm.n3162 C10_P_btm.n3161 4.60698
R30910 C10_P_btm.n3161 C10_P_btm.n3160 4.60698
R30911 C10_P_btm.n3159 C10_P_btm.n3158 4.60698
R30912 C10_P_btm.n3158 C10_P_btm.n3157 4.60698
R30913 C10_P_btm.n3156 C10_P_btm.n3155 4.60698
R30914 C10_P_btm.n3155 C10_P_btm.n3154 4.60698
R30915 C10_P_btm.n3153 C10_P_btm.n3152 4.60698
R30916 C10_P_btm.n3152 C10_P_btm.n3151 4.60698
R30917 C10_P_btm.n3150 C10_P_btm.n3149 4.60698
R30918 C10_P_btm.n3149 C10_P_btm.n3148 4.60698
R30919 C10_P_btm.n3147 C10_P_btm.n3146 4.60698
R30920 C10_P_btm.n3146 C10_P_btm.n3145 4.60698
R30921 C10_P_btm.n3144 C10_P_btm.n3143 4.60698
R30922 C10_P_btm.n3143 C10_P_btm.n3142 4.60698
R30923 C10_P_btm.n3141 C10_P_btm.n3140 4.60698
R30924 C10_P_btm.n3140 C10_P_btm.n3139 4.60698
R30925 C10_P_btm.n3138 C10_P_btm.n3137 4.60698
R30926 C10_P_btm.n3137 C10_P_btm.n3136 4.60698
R30927 C10_P_btm.n3135 C10_P_btm.n3134 4.60698
R30928 C10_P_btm.n3134 C10_P_btm.n3133 4.60698
R30929 C10_P_btm.n3132 C10_P_btm.n3131 4.60698
R30930 C10_P_btm.n3131 C10_P_btm.n3130 4.60698
R30931 C10_P_btm.n3129 C10_P_btm.n3128 4.60698
R30932 C10_P_btm.n3128 C10_P_btm.n3127 4.60698
R30933 C10_P_btm.n3126 C10_P_btm.n3125 4.60698
R30934 C10_P_btm.n3125 C10_P_btm.n3124 4.60698
R30935 C10_P_btm.n3123 C10_P_btm.n3122 4.60698
R30936 C10_P_btm.n3122 C10_P_btm.n3121 4.60698
R30937 C10_P_btm.n3120 C10_P_btm.n3119 4.60698
R30938 C10_P_btm.n3119 C10_P_btm.n3118 4.60698
R30939 C10_P_btm.n3117 C10_P_btm.n3116 4.60698
R30940 C10_P_btm.n3116 C10_P_btm.n3115 4.60698
R30941 C10_P_btm.n3114 C10_P_btm.n3113 4.60698
R30942 C10_P_btm.n3113 C10_P_btm.n3112 4.60698
R30943 C10_P_btm.n3111 C10_P_btm.n3110 4.60698
R30944 C10_P_btm.n3110 C10_P_btm.n3109 4.60698
R30945 C10_P_btm.n3103 C10_P_btm.n3102 4.60698
R30946 C10_P_btm.n3104 C10_P_btm.n3103 4.60698
R30947 C10_P_btm.n3100 C10_P_btm.n3099 4.60698
R30948 C10_P_btm.n3101 C10_P_btm.n3100 4.60698
R30949 C10_P_btm.n3097 C10_P_btm.n3096 4.60698
R30950 C10_P_btm.n3098 C10_P_btm.n3097 4.60698
R30951 C10_P_btm.n3094 C10_P_btm.n3093 4.60698
R30952 C10_P_btm.n3095 C10_P_btm.n3094 4.60698
R30953 C10_P_btm.n3091 C10_P_btm.n3090 4.60698
R30954 C10_P_btm.n3092 C10_P_btm.n3091 4.60698
R30955 C10_P_btm.n3088 C10_P_btm.n3087 4.60698
R30956 C10_P_btm.n3089 C10_P_btm.n3088 4.60698
R30957 C10_P_btm.n3085 C10_P_btm.n3084 4.60698
R30958 C10_P_btm.n3086 C10_P_btm.n3085 4.60698
R30959 C10_P_btm.n3082 C10_P_btm.n3081 4.60698
R30960 C10_P_btm.n3083 C10_P_btm.n3082 4.60698
R30961 C10_P_btm.n3079 C10_P_btm.n3078 4.60698
R30962 C10_P_btm.n3080 C10_P_btm.n3079 4.60698
R30963 C10_P_btm.n3076 C10_P_btm.n3075 4.60698
R30964 C10_P_btm.n3077 C10_P_btm.n3076 4.60698
R30965 C10_P_btm.n3022 C10_P_btm.n3021 4.60698
R30966 C10_P_btm.n3021 C10_P_btm.n3020 4.60698
R30967 C10_P_btm.n3019 C10_P_btm.n3018 4.60698
R30968 C10_P_btm.n3018 C10_P_btm.n3017 4.60698
R30969 C10_P_btm.n3016 C10_P_btm.n3015 4.60698
R30970 C10_P_btm.n3015 C10_P_btm.n3014 4.60698
R30971 C10_P_btm.n3013 C10_P_btm.n3012 4.60698
R30972 C10_P_btm.n3012 C10_P_btm.n3011 4.60698
R30973 C10_P_btm.n3010 C10_P_btm.n3009 4.60698
R30974 C10_P_btm.n3009 C10_P_btm.n3008 4.60698
R30975 C10_P_btm.n3007 C10_P_btm.n3006 4.60698
R30976 C10_P_btm.n3006 C10_P_btm.n3005 4.60698
R30977 C10_P_btm.n3004 C10_P_btm.n3003 4.60698
R30978 C10_P_btm.n3003 C10_P_btm.n3002 4.60698
R30979 C10_P_btm.n3001 C10_P_btm.n3000 4.60698
R30980 C10_P_btm.n3000 C10_P_btm.n2999 4.60698
R30981 C10_P_btm.n2998 C10_P_btm.n2997 4.60698
R30982 C10_P_btm.n2997 C10_P_btm.n2996 4.60698
R30983 C10_P_btm.n2992 C10_P_btm.n2991 4.60698
R30984 C10_P_btm.n2991 C10_P_btm.n2076 4.60698
R30985 C10_P_btm.n2989 C10_P_btm.n2988 4.60698
R30986 C10_P_btm.n2990 C10_P_btm.n2989 4.60698
R30987 C10_P_btm.n2986 C10_P_btm.n2985 4.60698
R30988 C10_P_btm.n2987 C10_P_btm.n2986 4.60698
R30989 C10_P_btm.n2983 C10_P_btm.n2982 4.60698
R30990 C10_P_btm.n2984 C10_P_btm.n2983 4.60698
R30991 C10_P_btm.n2980 C10_P_btm.n2979 4.60698
R30992 C10_P_btm.n2981 C10_P_btm.n2980 4.60698
R30993 C10_P_btm.n2977 C10_P_btm.n2976 4.60698
R30994 C10_P_btm.n2978 C10_P_btm.n2977 4.60698
R30995 C10_P_btm.n2974 C10_P_btm.n2973 4.60698
R30996 C10_P_btm.n2975 C10_P_btm.n2974 4.60698
R30997 C10_P_btm.n2971 C10_P_btm.n2970 4.60698
R30998 C10_P_btm.n2972 C10_P_btm.n2971 4.60698
R30999 C10_P_btm.n2968 C10_P_btm.n2967 4.60698
R31000 C10_P_btm.n2969 C10_P_btm.n2968 4.60698
R31001 C10_P_btm.n2963 C10_P_btm.n2962 4.60698
R31002 C10_P_btm.n2962 C10_P_btm.n2085 4.60698
R31003 C10_P_btm.n2904 C10_P_btm.n2903 4.60698
R31004 C10_P_btm.n2905 C10_P_btm.n2904 4.60698
R31005 C10_P_btm.n2907 C10_P_btm.n2906 4.60698
R31006 C10_P_btm.n2908 C10_P_btm.n2907 4.60698
R31007 C10_P_btm.n2910 C10_P_btm.n2909 4.60698
R31008 C10_P_btm.n2911 C10_P_btm.n2910 4.60698
R31009 C10_P_btm.n2913 C10_P_btm.n2912 4.60698
R31010 C10_P_btm.n2914 C10_P_btm.n2913 4.60698
R31011 C10_P_btm.n2916 C10_P_btm.n2915 4.60698
R31012 C10_P_btm.n2917 C10_P_btm.n2916 4.60698
R31013 C10_P_btm.n2919 C10_P_btm.n2918 4.60698
R31014 C10_P_btm.n2920 C10_P_btm.n2919 4.60698
R31015 C10_P_btm.n2922 C10_P_btm.n2921 4.60698
R31016 C10_P_btm.n2923 C10_P_btm.n2922 4.60698
R31017 C10_P_btm.n2925 C10_P_btm.n2924 4.60698
R31018 C10_P_btm.n2926 C10_P_btm.n2925 4.60698
R31019 C10_P_btm.n2933 C10_P_btm.n2932 4.60698
R31020 C10_P_btm.n2932 C10_P_btm.n2931 4.60698
R31021 C10_P_btm.n2936 C10_P_btm.n2935 4.60698
R31022 C10_P_btm.n2935 C10_P_btm.n2934 4.60698
R31023 C10_P_btm.n2939 C10_P_btm.n2938 4.60698
R31024 C10_P_btm.n2938 C10_P_btm.n2937 4.60698
R31025 C10_P_btm.n2942 C10_P_btm.n2941 4.60698
R31026 C10_P_btm.n2941 C10_P_btm.n2940 4.60698
R31027 C10_P_btm.n2945 C10_P_btm.n2944 4.60698
R31028 C10_P_btm.n2944 C10_P_btm.n2943 4.60698
R31029 C10_P_btm.n2948 C10_P_btm.n2947 4.60698
R31030 C10_P_btm.n2947 C10_P_btm.n2946 4.60698
R31031 C10_P_btm.n2951 C10_P_btm.n2950 4.60698
R31032 C10_P_btm.n2950 C10_P_btm.n2949 4.60698
R31033 C10_P_btm.n2954 C10_P_btm.n2953 4.60698
R31034 C10_P_btm.n2953 C10_P_btm.n2952 4.60698
R31035 C10_P_btm.n2957 C10_P_btm.n2956 4.60698
R31036 C10_P_btm.n2956 C10_P_btm.n2955 4.60698
R31037 C10_P_btm.n2866 C10_P_btm.n2865 4.60698
R31038 C10_P_btm.n2867 C10_P_btm.n2866 4.60698
R31039 C10_P_btm.n2869 C10_P_btm.n2868 4.60698
R31040 C10_P_btm.n2870 C10_P_btm.n2869 4.60698
R31041 C10_P_btm.n2872 C10_P_btm.n2871 4.60698
R31042 C10_P_btm.n2873 C10_P_btm.n2872 4.60698
R31043 C10_P_btm.n2875 C10_P_btm.n2874 4.60698
R31044 C10_P_btm.n2876 C10_P_btm.n2875 4.60698
R31045 C10_P_btm.n2878 C10_P_btm.n2877 4.60698
R31046 C10_P_btm.n2879 C10_P_btm.n2878 4.60698
R31047 C10_P_btm.n2881 C10_P_btm.n2880 4.60698
R31048 C10_P_btm.n2882 C10_P_btm.n2881 4.60698
R31049 C10_P_btm.n2884 C10_P_btm.n2883 4.60698
R31050 C10_P_btm.n2885 C10_P_btm.n2884 4.60698
R31051 C10_P_btm.n2887 C10_P_btm.n2886 4.60698
R31052 C10_P_btm.n2888 C10_P_btm.n2887 4.60698
R31053 C10_P_btm.n2890 C10_P_btm.n2889 4.60698
R31054 C10_P_btm.n2891 C10_P_btm.n2890 4.60698
R31055 C10_P_btm.n2145 C10_P_btm.n2144 4.60698
R31056 C10_P_btm.n2144 C10_P_btm.n2115 4.60698
R31057 C10_P_btm.n2142 C10_P_btm.n2141 4.60698
R31058 C10_P_btm.n2143 C10_P_btm.n2142 4.60698
R31059 C10_P_btm.n2139 C10_P_btm.n2138 4.60698
R31060 C10_P_btm.n2140 C10_P_btm.n2139 4.60698
R31061 C10_P_btm.n2136 C10_P_btm.n2135 4.60698
R31062 C10_P_btm.n2137 C10_P_btm.n2136 4.60698
R31063 C10_P_btm.n2133 C10_P_btm.n2132 4.60698
R31064 C10_P_btm.n2134 C10_P_btm.n2133 4.60698
R31065 C10_P_btm.n2130 C10_P_btm.n2129 4.60698
R31066 C10_P_btm.n2131 C10_P_btm.n2130 4.60698
R31067 C10_P_btm.n2127 C10_P_btm.n2126 4.60698
R31068 C10_P_btm.n2128 C10_P_btm.n2127 4.60698
R31069 C10_P_btm.n2124 C10_P_btm.n2123 4.60698
R31070 C10_P_btm.n2125 C10_P_btm.n2124 4.60698
R31071 C10_P_btm.n2861 C10_P_btm.n2860 4.60698
R31072 C10_P_btm.n2860 C10_P_btm.n2105 4.60698
R31073 C10_P_btm.n2855 C10_P_btm.n2854 4.60698
R31074 C10_P_btm.n2854 C10_P_btm.n2853 4.60698
R31075 C10_P_btm.n2852 C10_P_btm.n2851 4.60698
R31076 C10_P_btm.n2851 C10_P_btm.n2850 4.60698
R31077 C10_P_btm.n2849 C10_P_btm.n2848 4.60698
R31078 C10_P_btm.n2848 C10_P_btm.n2847 4.60698
R31079 C10_P_btm.n2846 C10_P_btm.n2845 4.60698
R31080 C10_P_btm.n2845 C10_P_btm.n2844 4.60698
R31081 C10_P_btm.n2843 C10_P_btm.n2842 4.60698
R31082 C10_P_btm.n2842 C10_P_btm.n2841 4.60698
R31083 C10_P_btm.n2840 C10_P_btm.n2839 4.60698
R31084 C10_P_btm.n2839 C10_P_btm.n2838 4.60698
R31085 C10_P_btm.n2837 C10_P_btm.n2836 4.60698
R31086 C10_P_btm.n2836 C10_P_btm.n2835 4.60698
R31087 C10_P_btm.n2834 C10_P_btm.n2833 4.60698
R31088 C10_P_btm.n2833 C10_P_btm.n2832 4.60698
R31089 C10_P_btm.n2831 C10_P_btm.n2830 4.60698
R31090 C10_P_btm.n2830 C10_P_btm.n2829 4.60698
R31091 C10_P_btm.n2823 C10_P_btm.n2822 4.60698
R31092 C10_P_btm.n2824 C10_P_btm.n2823 4.60698
R31093 C10_P_btm.n2820 C10_P_btm.n2819 4.60698
R31094 C10_P_btm.n2821 C10_P_btm.n2820 4.60698
R31095 C10_P_btm.n2817 C10_P_btm.n2816 4.60698
R31096 C10_P_btm.n2818 C10_P_btm.n2817 4.60698
R31097 C10_P_btm.n2814 C10_P_btm.n2813 4.60698
R31098 C10_P_btm.n2815 C10_P_btm.n2814 4.60698
R31099 C10_P_btm.n2811 C10_P_btm.n2810 4.60698
R31100 C10_P_btm.n2812 C10_P_btm.n2811 4.60698
R31101 C10_P_btm.n2808 C10_P_btm.n2807 4.60698
R31102 C10_P_btm.n2809 C10_P_btm.n2808 4.60698
R31103 C10_P_btm.n2805 C10_P_btm.n2804 4.60698
R31104 C10_P_btm.n2806 C10_P_btm.n2805 4.60698
R31105 C10_P_btm.n2802 C10_P_btm.n2801 4.60698
R31106 C10_P_btm.n2803 C10_P_btm.n2802 4.60698
R31107 C10_P_btm.n2799 C10_P_btm.n2798 4.60698
R31108 C10_P_btm.n2800 C10_P_btm.n2799 4.60698
R31109 C10_P_btm.n2794 C10_P_btm.n2793 4.60698
R31110 C10_P_btm.n2793 C10_P_btm.n2158 4.60698
R31111 C10_P_btm.n2177 C10_P_btm.n2176 4.60698
R31112 C10_P_btm.n2178 C10_P_btm.n2177 4.60698
R31113 C10_P_btm.n2180 C10_P_btm.n2179 4.60698
R31114 C10_P_btm.n2181 C10_P_btm.n2180 4.60698
R31115 C10_P_btm.n2183 C10_P_btm.n2182 4.60698
R31116 C10_P_btm.n2184 C10_P_btm.n2183 4.60698
R31117 C10_P_btm.n2186 C10_P_btm.n2185 4.60698
R31118 C10_P_btm.n2187 C10_P_btm.n2186 4.60698
R31119 C10_P_btm.n2189 C10_P_btm.n2188 4.60698
R31120 C10_P_btm.n2190 C10_P_btm.n2189 4.60698
R31121 C10_P_btm.n2192 C10_P_btm.n2191 4.60698
R31122 C10_P_btm.n2193 C10_P_btm.n2192 4.60698
R31123 C10_P_btm.n2195 C10_P_btm.n2194 4.60698
R31124 C10_P_btm.n2196 C10_P_btm.n2195 4.60698
R31125 C10_P_btm.n2198 C10_P_btm.n2197 4.60698
R31126 C10_P_btm.n2197 C10_P_btm.n2168 4.60698
R31127 C10_P_btm.n2764 C10_P_btm.n2763 4.60698
R31128 C10_P_btm.n2763 C10_P_btm.n2762 4.60698
R31129 C10_P_btm.n2767 C10_P_btm.n2766 4.60698
R31130 C10_P_btm.n2766 C10_P_btm.n2765 4.60698
R31131 C10_P_btm.n2770 C10_P_btm.n2769 4.60698
R31132 C10_P_btm.n2769 C10_P_btm.n2768 4.60698
R31133 C10_P_btm.n2773 C10_P_btm.n2772 4.60698
R31134 C10_P_btm.n2772 C10_P_btm.n2771 4.60698
R31135 C10_P_btm.n2776 C10_P_btm.n2775 4.60698
R31136 C10_P_btm.n2775 C10_P_btm.n2774 4.60698
R31137 C10_P_btm.n2779 C10_P_btm.n2778 4.60698
R31138 C10_P_btm.n2778 C10_P_btm.n2777 4.60698
R31139 C10_P_btm.n2782 C10_P_btm.n2781 4.60698
R31140 C10_P_btm.n2781 C10_P_btm.n2780 4.60698
R31141 C10_P_btm.n2785 C10_P_btm.n2784 4.60698
R31142 C10_P_btm.n2784 C10_P_btm.n2783 4.60698
R31143 C10_P_btm.n2788 C10_P_btm.n2787 4.60698
R31144 C10_P_btm.n2787 C10_P_btm.n2786 4.60698
R31145 C10_P_btm.n2732 C10_P_btm.n2731 4.60698
R31146 C10_P_btm.n2733 C10_P_btm.n2732 4.60698
R31147 C10_P_btm.n2735 C10_P_btm.n2734 4.60698
R31148 C10_P_btm.n2736 C10_P_btm.n2735 4.60698
R31149 C10_P_btm.n2738 C10_P_btm.n2737 4.60698
R31150 C10_P_btm.n2739 C10_P_btm.n2738 4.60698
R31151 C10_P_btm.n2741 C10_P_btm.n2740 4.60698
R31152 C10_P_btm.n2742 C10_P_btm.n2741 4.60698
R31153 C10_P_btm.n2744 C10_P_btm.n2743 4.60698
R31154 C10_P_btm.n2745 C10_P_btm.n2744 4.60698
R31155 C10_P_btm.n2747 C10_P_btm.n2746 4.60698
R31156 C10_P_btm.n2748 C10_P_btm.n2747 4.60698
R31157 C10_P_btm.n2750 C10_P_btm.n2749 4.60698
R31158 C10_P_btm.n2751 C10_P_btm.n2750 4.60698
R31159 C10_P_btm.n2753 C10_P_btm.n2752 4.60698
R31160 C10_P_btm.n2754 C10_P_btm.n2753 4.60698
R31161 C10_P_btm.n2756 C10_P_btm.n2755 4.60698
R31162 C10_P_btm.n2757 C10_P_btm.n2756 4.60698
R31163 C10_P_btm.n2251 C10_P_btm.n2250 4.60698
R31164 C10_P_btm.n2250 C10_P_btm.n2221 4.60698
R31165 C10_P_btm.n2248 C10_P_btm.n2247 4.60698
R31166 C10_P_btm.n2249 C10_P_btm.n2248 4.60698
R31167 C10_P_btm.n2245 C10_P_btm.n2244 4.60698
R31168 C10_P_btm.n2246 C10_P_btm.n2245 4.60698
R31169 C10_P_btm.n2242 C10_P_btm.n2241 4.60698
R31170 C10_P_btm.n2243 C10_P_btm.n2242 4.60698
R31171 C10_P_btm.n2239 C10_P_btm.n2238 4.60698
R31172 C10_P_btm.n2240 C10_P_btm.n2239 4.60698
R31173 C10_P_btm.n2236 C10_P_btm.n2235 4.60698
R31174 C10_P_btm.n2237 C10_P_btm.n2236 4.60698
R31175 C10_P_btm.n2233 C10_P_btm.n2232 4.60698
R31176 C10_P_btm.n2234 C10_P_btm.n2233 4.60698
R31177 C10_P_btm.n2230 C10_P_btm.n2229 4.60698
R31178 C10_P_btm.n2231 C10_P_btm.n2230 4.60698
R31179 C10_P_btm.n2727 C10_P_btm.n2726 4.60698
R31180 C10_P_btm.n2726 C10_P_btm.n2211 4.60698
R31181 C10_P_btm.n2721 C10_P_btm.n2720 4.60698
R31182 C10_P_btm.n2720 C10_P_btm.n2719 4.60698
R31183 C10_P_btm.n2718 C10_P_btm.n2717 4.60698
R31184 C10_P_btm.n2717 C10_P_btm.n2716 4.60698
R31185 C10_P_btm.n2715 C10_P_btm.n2714 4.60698
R31186 C10_P_btm.n2714 C10_P_btm.n2713 4.60698
R31187 C10_P_btm.n2712 C10_P_btm.n2711 4.60698
R31188 C10_P_btm.n2711 C10_P_btm.n2710 4.60698
R31189 C10_P_btm.n2709 C10_P_btm.n2708 4.60698
R31190 C10_P_btm.n2708 C10_P_btm.n2707 4.60698
R31191 C10_P_btm.n2706 C10_P_btm.n2705 4.60698
R31192 C10_P_btm.n2705 C10_P_btm.n2704 4.60698
R31193 C10_P_btm.n2703 C10_P_btm.n2702 4.60698
R31194 C10_P_btm.n2702 C10_P_btm.n2701 4.60698
R31195 C10_P_btm.n2700 C10_P_btm.n2699 4.60698
R31196 C10_P_btm.n2699 C10_P_btm.n2698 4.60698
R31197 C10_P_btm.n2697 C10_P_btm.n2696 4.60698
R31198 C10_P_btm.n2696 C10_P_btm.n2695 4.60698
R31199 C10_P_btm.n2689 C10_P_btm.n2688 4.60698
R31200 C10_P_btm.n2690 C10_P_btm.n2689 4.60698
R31201 C10_P_btm.n2686 C10_P_btm.n2685 4.60698
R31202 C10_P_btm.n2687 C10_P_btm.n2686 4.60698
R31203 C10_P_btm.n2683 C10_P_btm.n2682 4.60698
R31204 C10_P_btm.n2684 C10_P_btm.n2683 4.60698
R31205 C10_P_btm.n2680 C10_P_btm.n2679 4.60698
R31206 C10_P_btm.n2681 C10_P_btm.n2680 4.60698
R31207 C10_P_btm.n2677 C10_P_btm.n2676 4.60698
R31208 C10_P_btm.n2678 C10_P_btm.n2677 4.60698
R31209 C10_P_btm.n2674 C10_P_btm.n2673 4.60698
R31210 C10_P_btm.n2675 C10_P_btm.n2674 4.60698
R31211 C10_P_btm.n2671 C10_P_btm.n2670 4.60698
R31212 C10_P_btm.n2672 C10_P_btm.n2671 4.60698
R31213 C10_P_btm.n2668 C10_P_btm.n2667 4.60698
R31214 C10_P_btm.n2669 C10_P_btm.n2668 4.60698
R31215 C10_P_btm.n2665 C10_P_btm.n2664 4.60698
R31216 C10_P_btm.n2666 C10_P_btm.n2665 4.60698
R31217 C10_P_btm.n2660 C10_P_btm.n2659 4.60698
R31218 C10_P_btm.n2659 C10_P_btm.n2264 4.60698
R31219 C10_P_btm.n2283 C10_P_btm.n2282 4.60698
R31220 C10_P_btm.n2284 C10_P_btm.n2283 4.60698
R31221 C10_P_btm.n2286 C10_P_btm.n2285 4.60698
R31222 C10_P_btm.n2287 C10_P_btm.n2286 4.60698
R31223 C10_P_btm.n2289 C10_P_btm.n2288 4.60698
R31224 C10_P_btm.n2290 C10_P_btm.n2289 4.60698
R31225 C10_P_btm.n2292 C10_P_btm.n2291 4.60698
R31226 C10_P_btm.n2293 C10_P_btm.n2292 4.60698
R31227 C10_P_btm.n2295 C10_P_btm.n2294 4.60698
R31228 C10_P_btm.n2296 C10_P_btm.n2295 4.60698
R31229 C10_P_btm.n2298 C10_P_btm.n2297 4.60698
R31230 C10_P_btm.n2299 C10_P_btm.n2298 4.60698
R31231 C10_P_btm.n2301 C10_P_btm.n2300 4.60698
R31232 C10_P_btm.n2302 C10_P_btm.n2301 4.60698
R31233 C10_P_btm.n2304 C10_P_btm.n2303 4.60698
R31234 C10_P_btm.n2303 C10_P_btm.n2274 4.60698
R31235 C10_P_btm.n2630 C10_P_btm.n2629 4.60698
R31236 C10_P_btm.n2629 C10_P_btm.n2628 4.60698
R31237 C10_P_btm.n2633 C10_P_btm.n2632 4.60698
R31238 C10_P_btm.n2632 C10_P_btm.n2631 4.60698
R31239 C10_P_btm.n2636 C10_P_btm.n2635 4.60698
R31240 C10_P_btm.n2635 C10_P_btm.n2634 4.60698
R31241 C10_P_btm.n2639 C10_P_btm.n2638 4.60698
R31242 C10_P_btm.n2638 C10_P_btm.n2637 4.60698
R31243 C10_P_btm.n2642 C10_P_btm.n2641 4.60698
R31244 C10_P_btm.n2641 C10_P_btm.n2640 4.60698
R31245 C10_P_btm.n2645 C10_P_btm.n2644 4.60698
R31246 C10_P_btm.n2644 C10_P_btm.n2643 4.60698
R31247 C10_P_btm.n2648 C10_P_btm.n2647 4.60698
R31248 C10_P_btm.n2647 C10_P_btm.n2646 4.60698
R31249 C10_P_btm.n2651 C10_P_btm.n2650 4.60698
R31250 C10_P_btm.n2650 C10_P_btm.n2649 4.60698
R31251 C10_P_btm.n2654 C10_P_btm.n2653 4.60698
R31252 C10_P_btm.n2653 C10_P_btm.n2652 4.60698
R31253 C10_P_btm.n2598 C10_P_btm.n2597 4.60698
R31254 C10_P_btm.n2599 C10_P_btm.n2598 4.60698
R31255 C10_P_btm.n2601 C10_P_btm.n2600 4.60698
R31256 C10_P_btm.n2602 C10_P_btm.n2601 4.60698
R31257 C10_P_btm.n2604 C10_P_btm.n2603 4.60698
R31258 C10_P_btm.n2605 C10_P_btm.n2604 4.60698
R31259 C10_P_btm.n2607 C10_P_btm.n2606 4.60698
R31260 C10_P_btm.n2608 C10_P_btm.n2607 4.60698
R31261 C10_P_btm.n2610 C10_P_btm.n2609 4.60698
R31262 C10_P_btm.n2611 C10_P_btm.n2610 4.60698
R31263 C10_P_btm.n2613 C10_P_btm.n2612 4.60698
R31264 C10_P_btm.n2614 C10_P_btm.n2613 4.60698
R31265 C10_P_btm.n2616 C10_P_btm.n2615 4.60698
R31266 C10_P_btm.n2617 C10_P_btm.n2616 4.60698
R31267 C10_P_btm.n2619 C10_P_btm.n2618 4.60698
R31268 C10_P_btm.n2620 C10_P_btm.n2619 4.60698
R31269 C10_P_btm.n2622 C10_P_btm.n2621 4.60698
R31270 C10_P_btm.n2623 C10_P_btm.n2622 4.60698
R31271 C10_P_btm.n2357 C10_P_btm.n2356 4.60698
R31272 C10_P_btm.n2356 C10_P_btm.n2327 4.60698
R31273 C10_P_btm.n2354 C10_P_btm.n2353 4.60698
R31274 C10_P_btm.n2355 C10_P_btm.n2354 4.60698
R31275 C10_P_btm.n2351 C10_P_btm.n2350 4.60698
R31276 C10_P_btm.n2352 C10_P_btm.n2351 4.60698
R31277 C10_P_btm.n2348 C10_P_btm.n2347 4.60698
R31278 C10_P_btm.n2349 C10_P_btm.n2348 4.60698
R31279 C10_P_btm.n2345 C10_P_btm.n2344 4.60698
R31280 C10_P_btm.n2346 C10_P_btm.n2345 4.60698
R31281 C10_P_btm.n2342 C10_P_btm.n2341 4.60698
R31282 C10_P_btm.n2343 C10_P_btm.n2342 4.60698
R31283 C10_P_btm.n2339 C10_P_btm.n2338 4.60698
R31284 C10_P_btm.n2340 C10_P_btm.n2339 4.60698
R31285 C10_P_btm.n2336 C10_P_btm.n2335 4.60698
R31286 C10_P_btm.n2337 C10_P_btm.n2336 4.60698
R31287 C10_P_btm.n2593 C10_P_btm.n2592 4.60698
R31288 C10_P_btm.n2592 C10_P_btm.n2317 4.60698
R31289 C10_P_btm.n2587 C10_P_btm.n2586 4.60698
R31290 C10_P_btm.n2586 C10_P_btm.n2585 4.60698
R31291 C10_P_btm.n2584 C10_P_btm.n2583 4.60698
R31292 C10_P_btm.n2583 C10_P_btm.n2582 4.60698
R31293 C10_P_btm.n2581 C10_P_btm.n2580 4.60698
R31294 C10_P_btm.n2580 C10_P_btm.n2579 4.60698
R31295 C10_P_btm.n2578 C10_P_btm.n2577 4.60698
R31296 C10_P_btm.n2577 C10_P_btm.n2576 4.60698
R31297 C10_P_btm.n2575 C10_P_btm.n2574 4.60698
R31298 C10_P_btm.n2574 C10_P_btm.n2573 4.60698
R31299 C10_P_btm.n2572 C10_P_btm.n2571 4.60698
R31300 C10_P_btm.n2571 C10_P_btm.n2570 4.60698
R31301 C10_P_btm.n2569 C10_P_btm.n2568 4.60698
R31302 C10_P_btm.n2568 C10_P_btm.n2567 4.60698
R31303 C10_P_btm.n2566 C10_P_btm.n2565 4.60698
R31304 C10_P_btm.n2565 C10_P_btm.n2564 4.60698
R31305 C10_P_btm.n2563 C10_P_btm.n2562 4.60698
R31306 C10_P_btm.n2562 C10_P_btm.n2561 4.60698
R31307 C10_P_btm.n2555 C10_P_btm.n2554 4.60698
R31308 C10_P_btm.n2556 C10_P_btm.n2555 4.60698
R31309 C10_P_btm.n2552 C10_P_btm.n2551 4.60698
R31310 C10_P_btm.n2553 C10_P_btm.n2552 4.60698
R31311 C10_P_btm.n2549 C10_P_btm.n2548 4.60698
R31312 C10_P_btm.n2550 C10_P_btm.n2549 4.60698
R31313 C10_P_btm.n2546 C10_P_btm.n2545 4.60698
R31314 C10_P_btm.n2547 C10_P_btm.n2546 4.60698
R31315 C10_P_btm.n2543 C10_P_btm.n2542 4.60698
R31316 C10_P_btm.n2544 C10_P_btm.n2543 4.60698
R31317 C10_P_btm.n2540 C10_P_btm.n2539 4.60698
R31318 C10_P_btm.n2541 C10_P_btm.n2540 4.60698
R31319 C10_P_btm.n2537 C10_P_btm.n2536 4.60698
R31320 C10_P_btm.n2538 C10_P_btm.n2537 4.60698
R31321 C10_P_btm.n2534 C10_P_btm.n2533 4.60698
R31322 C10_P_btm.n2535 C10_P_btm.n2534 4.60698
R31323 C10_P_btm.n2531 C10_P_btm.n2530 4.60698
R31324 C10_P_btm.n2532 C10_P_btm.n2531 4.60698
R31325 C10_P_btm.n2526 C10_P_btm.n2525 4.60698
R31326 C10_P_btm.n2525 C10_P_btm.n2370 4.60698
R31327 C10_P_btm.n2389 C10_P_btm.n2388 4.60698
R31328 C10_P_btm.n2390 C10_P_btm.n2389 4.60698
R31329 C10_P_btm.n2392 C10_P_btm.n2391 4.60698
R31330 C10_P_btm.n2393 C10_P_btm.n2392 4.60698
R31331 C10_P_btm.n2395 C10_P_btm.n2394 4.60698
R31332 C10_P_btm.n2396 C10_P_btm.n2395 4.60698
R31333 C10_P_btm.n2398 C10_P_btm.n2397 4.60698
R31334 C10_P_btm.n2399 C10_P_btm.n2398 4.60698
R31335 C10_P_btm.n2401 C10_P_btm.n2400 4.60698
R31336 C10_P_btm.n2402 C10_P_btm.n2401 4.60698
R31337 C10_P_btm.n2404 C10_P_btm.n2403 4.60698
R31338 C10_P_btm.n2405 C10_P_btm.n2404 4.60698
R31339 C10_P_btm.n2407 C10_P_btm.n2406 4.60698
R31340 C10_P_btm.n2408 C10_P_btm.n2407 4.60698
R31341 C10_P_btm.n2410 C10_P_btm.n2409 4.60698
R31342 C10_P_btm.n2409 C10_P_btm.n2380 4.60698
R31343 C10_P_btm.n2496 C10_P_btm.n2495 4.60698
R31344 C10_P_btm.n2495 C10_P_btm.n2494 4.60698
R31345 C10_P_btm.n2499 C10_P_btm.n2498 4.60698
R31346 C10_P_btm.n2498 C10_P_btm.n2497 4.60698
R31347 C10_P_btm.n2502 C10_P_btm.n2501 4.60698
R31348 C10_P_btm.n2501 C10_P_btm.n2500 4.60698
R31349 C10_P_btm.n2505 C10_P_btm.n2504 4.60698
R31350 C10_P_btm.n2504 C10_P_btm.n2503 4.60698
R31351 C10_P_btm.n2508 C10_P_btm.n2507 4.60698
R31352 C10_P_btm.n2507 C10_P_btm.n2506 4.60698
R31353 C10_P_btm.n2511 C10_P_btm.n2510 4.60698
R31354 C10_P_btm.n2510 C10_P_btm.n2509 4.60698
R31355 C10_P_btm.n2514 C10_P_btm.n2513 4.60698
R31356 C10_P_btm.n2513 C10_P_btm.n2512 4.60698
R31357 C10_P_btm.n2517 C10_P_btm.n2516 4.60698
R31358 C10_P_btm.n2516 C10_P_btm.n2515 4.60698
R31359 C10_P_btm.n2520 C10_P_btm.n2519 4.60698
R31360 C10_P_btm.n2519 C10_P_btm.n2518 4.60698
R31361 C10_P_btm.n2464 C10_P_btm.n2463 4.60698
R31362 C10_P_btm.n2465 C10_P_btm.n2464 4.60698
R31363 C10_P_btm.n2467 C10_P_btm.n2466 4.60698
R31364 C10_P_btm.n2468 C10_P_btm.n2467 4.60698
R31365 C10_P_btm.n2470 C10_P_btm.n2469 4.60698
R31366 C10_P_btm.n2471 C10_P_btm.n2470 4.60698
R31367 C10_P_btm.n2473 C10_P_btm.n2472 4.60698
R31368 C10_P_btm.n2474 C10_P_btm.n2473 4.60698
R31369 C10_P_btm.n2476 C10_P_btm.n2475 4.60698
R31370 C10_P_btm.n2477 C10_P_btm.n2476 4.60698
R31371 C10_P_btm.n2479 C10_P_btm.n2478 4.60698
R31372 C10_P_btm.n2480 C10_P_btm.n2479 4.60698
R31373 C10_P_btm.n2482 C10_P_btm.n2481 4.60698
R31374 C10_P_btm.n2483 C10_P_btm.n2482 4.60698
R31375 C10_P_btm.n2485 C10_P_btm.n2484 4.60698
R31376 C10_P_btm.n2486 C10_P_btm.n2485 4.60698
R31377 C10_P_btm.n2488 C10_P_btm.n2487 4.60698
R31378 C10_P_btm.n2489 C10_P_btm.n2488 4.60698
R31379 C10_P_btm.n2432 C10_P_btm.n2431 4.60698
R31380 C10_P_btm.n2433 C10_P_btm.n2432 4.60698
R31381 C10_P_btm.n2435 C10_P_btm.n2434 4.60698
R31382 C10_P_btm.n2436 C10_P_btm.n2435 4.60698
R31383 C10_P_btm.n2438 C10_P_btm.n2437 4.60698
R31384 C10_P_btm.n2439 C10_P_btm.n2438 4.60698
R31385 C10_P_btm.n2441 C10_P_btm.n2440 4.60698
R31386 C10_P_btm.n2442 C10_P_btm.n2441 4.60698
R31387 C10_P_btm.n2444 C10_P_btm.n2443 4.60698
R31388 C10_P_btm.n2445 C10_P_btm.n2444 4.60698
R31389 C10_P_btm.n2447 C10_P_btm.n2446 4.60698
R31390 C10_P_btm.n2448 C10_P_btm.n2447 4.60698
R31391 C10_P_btm.n2450 C10_P_btm.n2449 4.60698
R31392 C10_P_btm.n2451 C10_P_btm.n2450 4.60698
R31393 C10_P_btm.n2453 C10_P_btm.n2452 4.60698
R31394 C10_P_btm.n2454 C10_P_btm.n2453 4.60698
R31395 C10_P_btm.n2458 C10_P_btm.n2455 4.60698
R31396 C10_P_btm.n2459 C10_P_btm.n2458 4.60698
R31397 C10_P_btm.n3074 C10_P_btm.n3073 4.60698
R31398 C10_P_btm.n3073 C10_P_btm.n3072 4.60698
R31399 C10_P_btm.n3071 C10_P_btm.n3070 4.60698
R31400 C10_P_btm.n3070 C10_P_btm.n3069 4.60698
R31401 C10_P_btm.n3068 C10_P_btm.n3067 4.60698
R31402 C10_P_btm.n3067 C10_P_btm.n3066 4.60698
R31403 C10_P_btm.n3065 C10_P_btm.n3064 4.60698
R31404 C10_P_btm.n3064 C10_P_btm.n3063 4.60698
R31405 C10_P_btm.n3062 C10_P_btm.n3061 4.60698
R31406 C10_P_btm.n3061 C10_P_btm.n3060 4.60698
R31407 C10_P_btm.n3059 C10_P_btm.n3058 4.60698
R31408 C10_P_btm.n3058 C10_P_btm.n3057 4.60698
R31409 C10_P_btm.n3056 C10_P_btm.n3055 4.60698
R31410 C10_P_btm.n3055 C10_P_btm.n3054 4.60698
R31411 C10_P_btm.n3053 C10_P_btm.n3052 4.60698
R31412 C10_P_btm.n3052 C10_P_btm.n3051 4.60698
R31413 C10_P_btm.n3050 C10_P_btm.n3049 4.60698
R31414 C10_P_btm.n3049 C10_P_btm.n3048 4.60698
R31415 C10_P_btm.n3047 C10_P_btm.n3046 4.60698
R31416 C10_P_btm.n3046 C10_P_btm.n3045 4.60698
R31417 C10_P_btm.n3044 C10_P_btm.n3043 4.60698
R31418 C10_P_btm.n3043 C10_P_btm.n3042 4.60698
R31419 C10_P_btm.n3041 C10_P_btm.n3040 4.60698
R31420 C10_P_btm.n3040 C10_P_btm.n3039 4.60698
R31421 C10_P_btm.n2052 C10_P_btm.n2051 4.60698
R31422 C10_P_btm.n2053 C10_P_btm.n2052 4.60698
R31423 C10_P_btm.n2049 C10_P_btm.n2048 4.60698
R31424 C10_P_btm.n2050 C10_P_btm.n2049 4.60698
R31425 C10_P_btm.n2046 C10_P_btm.n2045 4.60698
R31426 C10_P_btm.n2047 C10_P_btm.n2046 4.60698
R31427 C10_P_btm.n2043 C10_P_btm.n2042 4.60698
R31428 C10_P_btm.n2044 C10_P_btm.n2043 4.60698
R31429 C10_P_btm.n2040 C10_P_btm.n2039 4.60698
R31430 C10_P_btm.n2041 C10_P_btm.n2040 4.60698
R31431 C10_P_btm.n2037 C10_P_btm.n2036 4.60698
R31432 C10_P_btm.n2038 C10_P_btm.n2037 4.60698
R31433 C10_P_btm.n2034 C10_P_btm.n2033 4.60698
R31434 C10_P_btm.n2035 C10_P_btm.n2034 4.60698
R31435 C10_P_btm.n2031 C10_P_btm.n2030 4.60698
R31436 C10_P_btm.n2032 C10_P_btm.n2031 4.60698
R31437 C10_P_btm.n2028 C10_P_btm.n2027 4.60698
R31438 C10_P_btm.n2029 C10_P_btm.n2028 4.60698
R31439 C10_P_btm.n2025 C10_P_btm.n2024 4.60698
R31440 C10_P_btm.n2026 C10_P_btm.n2025 4.60698
R31441 C10_P_btm.n2022 C10_P_btm.n2021 4.60698
R31442 C10_P_btm.n2023 C10_P_btm.n2022 4.60698
R31443 C10_P_btm.n2019 C10_P_btm.n2018 4.60698
R31444 C10_P_btm.n2020 C10_P_btm.n2019 4.60698
R31445 C10_P_btm.n2016 C10_P_btm.n2015 4.60698
R31446 C10_P_btm.n2017 C10_P_btm.n2016 4.60698
R31447 C10_P_btm.n2013 C10_P_btm.n2012 4.60698
R31448 C10_P_btm.n2014 C10_P_btm.n2013 4.60698
R31449 C10_P_btm.n2010 C10_P_btm.n2009 4.60698
R31450 C10_P_btm.n2011 C10_P_btm.n2010 4.60698
R31451 C10_P_btm.n2007 C10_P_btm.n2006 4.60698
R31452 C10_P_btm.n2008 C10_P_btm.n2007 4.60698
R31453 C10_P_btm.n2004 C10_P_btm.n2003 4.60698
R31454 C10_P_btm.n2005 C10_P_btm.n2004 4.60698
R31455 C10_P_btm.n2001 C10_P_btm.n2000 4.60698
R31456 C10_P_btm.n2002 C10_P_btm.n2001 4.60698
R31457 C10_P_btm.n1998 C10_P_btm.n1997 4.60698
R31458 C10_P_btm.n1999 C10_P_btm.n1998 4.60698
R31459 C10_P_btm.n1995 C10_P_btm.n1994 4.60698
R31460 C10_P_btm.n1996 C10_P_btm.n1995 4.60698
R31461 C10_P_btm.n1992 C10_P_btm.n1991 4.60698
R31462 C10_P_btm.n1993 C10_P_btm.n1992 4.60698
R31463 C10_P_btm.n1989 C10_P_btm.n1988 4.60698
R31464 C10_P_btm.n1990 C10_P_btm.n1989 4.60698
R31465 C10_P_btm.n1986 C10_P_btm.n1985 4.60698
R31466 C10_P_btm.n1987 C10_P_btm.n1986 4.60698
R31467 C10_P_btm.n1983 C10_P_btm.n1982 4.60698
R31468 C10_P_btm.n1984 C10_P_btm.n1983 4.60698
R31469 C10_P_btm.n1980 C10_P_btm.n1979 4.60698
R31470 C10_P_btm.n1981 C10_P_btm.n1980 4.60698
R31471 C10_P_btm.n1977 C10_P_btm.n1976 4.60698
R31472 C10_P_btm.n1978 C10_P_btm.n1977 4.60698
R31473 C10_P_btm.n1974 C10_P_btm.n1973 4.60698
R31474 C10_P_btm.n1975 C10_P_btm.n1974 4.60698
R31475 C10_P_btm.n1971 C10_P_btm.n1970 4.60698
R31476 C10_P_btm.n1972 C10_P_btm.n1971 4.60698
R31477 C10_P_btm.n1968 C10_P_btm.n1967 4.60698
R31478 C10_P_btm.n1969 C10_P_btm.n1968 4.60698
R31479 C10_P_btm.n1965 C10_P_btm.n1964 4.60698
R31480 C10_P_btm.n1966 C10_P_btm.n1965 4.60698
R31481 C10_P_btm.n1962 C10_P_btm.n1961 4.60698
R31482 C10_P_btm.n1963 C10_P_btm.n1962 4.60698
R31483 C10_P_btm.n1959 C10_P_btm.n1958 4.60698
R31484 C10_P_btm.n1960 C10_P_btm.n1959 4.60698
R31485 C10_P_btm.n1956 C10_P_btm.n1955 4.60698
R31486 C10_P_btm.n1957 C10_P_btm.n1956 4.60698
R31487 C10_P_btm.n1953 C10_P_btm.n1952 4.60698
R31488 C10_P_btm.n1954 C10_P_btm.n1953 4.60698
R31489 C10_P_btm.n1950 C10_P_btm.n1949 4.60698
R31490 C10_P_btm.n1951 C10_P_btm.n1950 4.60698
R31491 C10_P_btm.n1947 C10_P_btm.n1946 4.60698
R31492 C10_P_btm.n1948 C10_P_btm.n1947 4.60698
R31493 C10_P_btm.n1944 C10_P_btm.n1943 4.60698
R31494 C10_P_btm.n1945 C10_P_btm.n1944 4.60698
R31495 C10_P_btm.n1941 C10_P_btm.n1940 4.60698
R31496 C10_P_btm.n1942 C10_P_btm.n1941 4.60698
R31497 C10_P_btm.n1938 C10_P_btm.n1937 4.60698
R31498 C10_P_btm.n1939 C10_P_btm.n1938 4.60698
R31499 C10_P_btm.n1935 C10_P_btm.n1934 4.60698
R31500 C10_P_btm.n1936 C10_P_btm.n1935 4.60698
R31501 C10_P_btm.n1932 C10_P_btm.n1931 4.60698
R31502 C10_P_btm.n1933 C10_P_btm.n1932 4.60698
R31503 C10_P_btm.n1929 C10_P_btm.n1928 4.60698
R31504 C10_P_btm.n1930 C10_P_btm.n1929 4.60698
R31505 C10_P_btm.n1926 C10_P_btm.n1925 4.60698
R31506 C10_P_btm.n1927 C10_P_btm.n1926 4.60698
R31507 C10_P_btm.n1923 C10_P_btm.n1922 4.60698
R31508 C10_P_btm.n1924 C10_P_btm.n1923 4.60698
R31509 C10_P_btm.n1920 C10_P_btm.n1919 4.60698
R31510 C10_P_btm.n1921 C10_P_btm.n1920 4.60698
R31511 C10_P_btm.n1917 C10_P_btm.n1916 4.60698
R31512 C10_P_btm.n1918 C10_P_btm.n1917 4.60698
R31513 C10_P_btm.n1914 C10_P_btm.n1913 4.60698
R31514 C10_P_btm.n1915 C10_P_btm.n1914 4.60698
R31515 C10_P_btm.n1911 C10_P_btm.n1910 4.60698
R31516 C10_P_btm.n1912 C10_P_btm.n1911 4.60698
R31517 C10_P_btm.n1908 C10_P_btm.n1907 4.60698
R31518 C10_P_btm.n1909 C10_P_btm.n1908 4.60698
R31519 C10_P_btm.n1905 C10_P_btm.n1904 4.60698
R31520 C10_P_btm.n1906 C10_P_btm.n1905 4.60698
R31521 C10_P_btm.n1902 C10_P_btm.n1901 4.60698
R31522 C10_P_btm.n1903 C10_P_btm.n1902 4.60698
R31523 C10_P_btm.n1899 C10_P_btm.n1898 4.60698
R31524 C10_P_btm.n1900 C10_P_btm.n1899 4.60698
R31525 C10_P_btm.n1896 C10_P_btm.n1895 4.60698
R31526 C10_P_btm.n1897 C10_P_btm.n1896 4.60698
R31527 C10_P_btm.n1893 C10_P_btm.n1892 4.60698
R31528 C10_P_btm.n1894 C10_P_btm.n1893 4.60698
R31529 C10_P_btm.n1890 C10_P_btm.n1889 4.60698
R31530 C10_P_btm.n1891 C10_P_btm.n1890 4.60698
R31531 C10_P_btm.n1887 C10_P_btm.n1886 4.60698
R31532 C10_P_btm.n1888 C10_P_btm.n1887 4.60698
R31533 C10_P_btm.n1884 C10_P_btm.n1883 4.60698
R31534 C10_P_btm.n1885 C10_P_btm.n1884 4.60698
R31535 C10_P_btm.n1881 C10_P_btm.n1880 4.60698
R31536 C10_P_btm.n1882 C10_P_btm.n1881 4.60698
R31537 C10_P_btm.n1878 C10_P_btm.n1877 4.60698
R31538 C10_P_btm.n1879 C10_P_btm.n1878 4.60698
R31539 C10_P_btm.n1875 C10_P_btm.n1874 4.60698
R31540 C10_P_btm.n1876 C10_P_btm.n1875 4.60698
R31541 C10_P_btm.n1872 C10_P_btm.n1871 4.60698
R31542 C10_P_btm.n1873 C10_P_btm.n1872 4.60698
R31543 C10_P_btm.n1869 C10_P_btm.n1868 4.60698
R31544 C10_P_btm.n1870 C10_P_btm.n1869 4.60698
R31545 C10_P_btm.n1864 C10_P_btm.n1863 4.60698
R31546 C10_P_btm.n1863 C10_P_btm.n610 4.60698
R31547 C10_P_btm.n735 C10_P_btm.n734 4.60698
R31548 C10_P_btm.n736 C10_P_btm.n735 4.60698
R31549 C10_P_btm.n738 C10_P_btm.n737 4.60698
R31550 C10_P_btm.n739 C10_P_btm.n738 4.60698
R31551 C10_P_btm.n741 C10_P_btm.n740 4.60698
R31552 C10_P_btm.n742 C10_P_btm.n741 4.60698
R31553 C10_P_btm.n744 C10_P_btm.n743 4.60698
R31554 C10_P_btm.n745 C10_P_btm.n744 4.60698
R31555 C10_P_btm.n747 C10_P_btm.n746 4.60698
R31556 C10_P_btm.n748 C10_P_btm.n747 4.60698
R31557 C10_P_btm.n750 C10_P_btm.n749 4.60698
R31558 C10_P_btm.n751 C10_P_btm.n750 4.60698
R31559 C10_P_btm.n753 C10_P_btm.n752 4.60698
R31560 C10_P_btm.n754 C10_P_btm.n753 4.60698
R31561 C10_P_btm.n756 C10_P_btm.n755 4.60698
R31562 C10_P_btm.n757 C10_P_btm.n756 4.60698
R31563 C10_P_btm.n759 C10_P_btm.n758 4.60698
R31564 C10_P_btm.n760 C10_P_btm.n759 4.60698
R31565 C10_P_btm.n762 C10_P_btm.n761 4.60698
R31566 C10_P_btm.n763 C10_P_btm.n762 4.60698
R31567 C10_P_btm.n765 C10_P_btm.n764 4.60698
R31568 C10_P_btm.n766 C10_P_btm.n765 4.60698
R31569 C10_P_btm.n768 C10_P_btm.n767 4.60698
R31570 C10_P_btm.n769 C10_P_btm.n768 4.60698
R31571 C10_P_btm.n771 C10_P_btm.n770 4.60698
R31572 C10_P_btm.n772 C10_P_btm.n771 4.60698
R31573 C10_P_btm.n774 C10_P_btm.n773 4.60698
R31574 C10_P_btm.n775 C10_P_btm.n774 4.60698
R31575 C10_P_btm.n777 C10_P_btm.n776 4.60698
R31576 C10_P_btm.n778 C10_P_btm.n777 4.60698
R31577 C10_P_btm.n780 C10_P_btm.n779 4.60698
R31578 C10_P_btm.n781 C10_P_btm.n780 4.60698
R31579 C10_P_btm.n783 C10_P_btm.n782 4.60698
R31580 C10_P_btm.n784 C10_P_btm.n783 4.60698
R31581 C10_P_btm.n786 C10_P_btm.n785 4.60698
R31582 C10_P_btm.n787 C10_P_btm.n786 4.60698
R31583 C10_P_btm.n789 C10_P_btm.n788 4.60698
R31584 C10_P_btm.n790 C10_P_btm.n789 4.60698
R31585 C10_P_btm.n792 C10_P_btm.n791 4.60698
R31586 C10_P_btm.n793 C10_P_btm.n792 4.60698
R31587 C10_P_btm.n795 C10_P_btm.n794 4.60698
R31588 C10_P_btm.n796 C10_P_btm.n795 4.60698
R31589 C10_P_btm.n798 C10_P_btm.n797 4.60698
R31590 C10_P_btm.n799 C10_P_btm.n798 4.60698
R31591 C10_P_btm.n801 C10_P_btm.n800 4.60698
R31592 C10_P_btm.n802 C10_P_btm.n801 4.60698
R31593 C10_P_btm.n804 C10_P_btm.n803 4.60698
R31594 C10_P_btm.n805 C10_P_btm.n804 4.60698
R31595 C10_P_btm.n807 C10_P_btm.n806 4.60698
R31596 C10_P_btm.n808 C10_P_btm.n807 4.60698
R31597 C10_P_btm.n810 C10_P_btm.n809 4.60698
R31598 C10_P_btm.n811 C10_P_btm.n810 4.60698
R31599 C10_P_btm.n813 C10_P_btm.n812 4.60698
R31600 C10_P_btm.n814 C10_P_btm.n813 4.60698
R31601 C10_P_btm.n816 C10_P_btm.n815 4.60698
R31602 C10_P_btm.n817 C10_P_btm.n816 4.60698
R31603 C10_P_btm.n819 C10_P_btm.n818 4.60698
R31604 C10_P_btm.n820 C10_P_btm.n819 4.60698
R31605 C10_P_btm.n822 C10_P_btm.n821 4.60698
R31606 C10_P_btm.n823 C10_P_btm.n822 4.60698
R31607 C10_P_btm.n825 C10_P_btm.n824 4.60698
R31608 C10_P_btm.n826 C10_P_btm.n825 4.60698
R31609 C10_P_btm.n828 C10_P_btm.n827 4.60698
R31610 C10_P_btm.n829 C10_P_btm.n828 4.60698
R31611 C10_P_btm.n831 C10_P_btm.n830 4.60698
R31612 C10_P_btm.n832 C10_P_btm.n831 4.60698
R31613 C10_P_btm.n834 C10_P_btm.n833 4.60698
R31614 C10_P_btm.n835 C10_P_btm.n834 4.60698
R31615 C10_P_btm.n837 C10_P_btm.n836 4.60698
R31616 C10_P_btm.n838 C10_P_btm.n837 4.60698
R31617 C10_P_btm.n840 C10_P_btm.n839 4.60698
R31618 C10_P_btm.n841 C10_P_btm.n840 4.60698
R31619 C10_P_btm.n843 C10_P_btm.n842 4.60698
R31620 C10_P_btm.n844 C10_P_btm.n843 4.60698
R31621 C10_P_btm.n846 C10_P_btm.n845 4.60698
R31622 C10_P_btm.n847 C10_P_btm.n846 4.60698
R31623 C10_P_btm.n849 C10_P_btm.n848 4.60698
R31624 C10_P_btm.n850 C10_P_btm.n849 4.60698
R31625 C10_P_btm.n852 C10_P_btm.n851 4.60698
R31626 C10_P_btm.n853 C10_P_btm.n852 4.60698
R31627 C10_P_btm.n855 C10_P_btm.n854 4.60698
R31628 C10_P_btm.n856 C10_P_btm.n855 4.60698
R31629 C10_P_btm.n858 C10_P_btm.n857 4.60698
R31630 C10_P_btm.n859 C10_P_btm.n858 4.60698
R31631 C10_P_btm.n861 C10_P_btm.n860 4.60698
R31632 C10_P_btm.n862 C10_P_btm.n861 4.60698
R31633 C10_P_btm.n864 C10_P_btm.n863 4.60698
R31634 C10_P_btm.n865 C10_P_btm.n864 4.60698
R31635 C10_P_btm.n867 C10_P_btm.n866 4.60698
R31636 C10_P_btm.n868 C10_P_btm.n867 4.60698
R31637 C10_P_btm.n870 C10_P_btm.n869 4.60698
R31638 C10_P_btm.n871 C10_P_btm.n870 4.60698
R31639 C10_P_btm.n873 C10_P_btm.n872 4.60698
R31640 C10_P_btm.n874 C10_P_btm.n873 4.60698
R31641 C10_P_btm.n876 C10_P_btm.n875 4.60698
R31642 C10_P_btm.n877 C10_P_btm.n876 4.60698
R31643 C10_P_btm.n879 C10_P_btm.n878 4.60698
R31644 C10_P_btm.n880 C10_P_btm.n879 4.60698
R31645 C10_P_btm.n882 C10_P_btm.n881 4.60698
R31646 C10_P_btm.n883 C10_P_btm.n882 4.60698
R31647 C10_P_btm.n885 C10_P_btm.n884 4.60698
R31648 C10_P_btm.n886 C10_P_btm.n885 4.60698
R31649 C10_P_btm.n888 C10_P_btm.n887 4.60698
R31650 C10_P_btm.n889 C10_P_btm.n888 4.60698
R31651 C10_P_btm.n891 C10_P_btm.n890 4.60698
R31652 C10_P_btm.n892 C10_P_btm.n891 4.60698
R31653 C10_P_btm.n894 C10_P_btm.n893 4.60698
R31654 C10_P_btm.n895 C10_P_btm.n894 4.60698
R31655 C10_P_btm.n897 C10_P_btm.n896 4.60698
R31656 C10_P_btm.n898 C10_P_btm.n897 4.60698
R31657 C10_P_btm.n900 C10_P_btm.n899 4.60698
R31658 C10_P_btm.n901 C10_P_btm.n900 4.60698
R31659 C10_P_btm.n903 C10_P_btm.n902 4.60698
R31660 C10_P_btm.n904 C10_P_btm.n903 4.60698
R31661 C10_P_btm.n906 C10_P_btm.n905 4.60698
R31662 C10_P_btm.n907 C10_P_btm.n906 4.60698
R31663 C10_P_btm.n909 C10_P_btm.n908 4.60698
R31664 C10_P_btm.n910 C10_P_btm.n909 4.60698
R31665 C10_P_btm.n912 C10_P_btm.n911 4.60698
R31666 C10_P_btm.n913 C10_P_btm.n912 4.60698
R31667 C10_P_btm.n915 C10_P_btm.n914 4.60698
R31668 C10_P_btm.n914 C10_P_btm.n673 4.60698
R31669 C10_P_btm.n1675 C10_P_btm.n1674 4.60698
R31670 C10_P_btm.n1674 C10_P_btm.n1673 4.60698
R31671 C10_P_btm.n1678 C10_P_btm.n1677 4.60698
R31672 C10_P_btm.n1677 C10_P_btm.n1676 4.60698
R31673 C10_P_btm.n1681 C10_P_btm.n1680 4.60698
R31674 C10_P_btm.n1680 C10_P_btm.n1679 4.60698
R31675 C10_P_btm.n1684 C10_P_btm.n1683 4.60698
R31676 C10_P_btm.n1683 C10_P_btm.n1682 4.60698
R31677 C10_P_btm.n1687 C10_P_btm.n1686 4.60698
R31678 C10_P_btm.n1686 C10_P_btm.n1685 4.60698
R31679 C10_P_btm.n1690 C10_P_btm.n1689 4.60698
R31680 C10_P_btm.n1689 C10_P_btm.n1688 4.60698
R31681 C10_P_btm.n1693 C10_P_btm.n1692 4.60698
R31682 C10_P_btm.n1692 C10_P_btm.n1691 4.60698
R31683 C10_P_btm.n1696 C10_P_btm.n1695 4.60698
R31684 C10_P_btm.n1695 C10_P_btm.n1694 4.60698
R31685 C10_P_btm.n1699 C10_P_btm.n1698 4.60698
R31686 C10_P_btm.n1698 C10_P_btm.n1697 4.60698
R31687 C10_P_btm.n1702 C10_P_btm.n1701 4.60698
R31688 C10_P_btm.n1701 C10_P_btm.n1700 4.60698
R31689 C10_P_btm.n1705 C10_P_btm.n1704 4.60698
R31690 C10_P_btm.n1704 C10_P_btm.n1703 4.60698
R31691 C10_P_btm.n1708 C10_P_btm.n1707 4.60698
R31692 C10_P_btm.n1707 C10_P_btm.n1706 4.60698
R31693 C10_P_btm.n1711 C10_P_btm.n1710 4.60698
R31694 C10_P_btm.n1710 C10_P_btm.n1709 4.60698
R31695 C10_P_btm.n1714 C10_P_btm.n1713 4.60698
R31696 C10_P_btm.n1713 C10_P_btm.n1712 4.60698
R31697 C10_P_btm.n1717 C10_P_btm.n1716 4.60698
R31698 C10_P_btm.n1716 C10_P_btm.n1715 4.60698
R31699 C10_P_btm.n1720 C10_P_btm.n1719 4.60698
R31700 C10_P_btm.n1719 C10_P_btm.n1718 4.60698
R31701 C10_P_btm.n1723 C10_P_btm.n1722 4.60698
R31702 C10_P_btm.n1722 C10_P_btm.n1721 4.60698
R31703 C10_P_btm.n1726 C10_P_btm.n1725 4.60698
R31704 C10_P_btm.n1725 C10_P_btm.n1724 4.60698
R31705 C10_P_btm.n1729 C10_P_btm.n1728 4.60698
R31706 C10_P_btm.n1728 C10_P_btm.n1727 4.60698
R31707 C10_P_btm.n1732 C10_P_btm.n1731 4.60698
R31708 C10_P_btm.n1731 C10_P_btm.n1730 4.60698
R31709 C10_P_btm.n1735 C10_P_btm.n1734 4.60698
R31710 C10_P_btm.n1734 C10_P_btm.n1733 4.60698
R31711 C10_P_btm.n1738 C10_P_btm.n1737 4.60698
R31712 C10_P_btm.n1737 C10_P_btm.n1736 4.60698
R31713 C10_P_btm.n1741 C10_P_btm.n1740 4.60698
R31714 C10_P_btm.n1740 C10_P_btm.n1739 4.60698
R31715 C10_P_btm.n1744 C10_P_btm.n1743 4.60698
R31716 C10_P_btm.n1743 C10_P_btm.n1742 4.60698
R31717 C10_P_btm.n1747 C10_P_btm.n1746 4.60698
R31718 C10_P_btm.n1746 C10_P_btm.n1745 4.60698
R31719 C10_P_btm.n1750 C10_P_btm.n1749 4.60698
R31720 C10_P_btm.n1749 C10_P_btm.n1748 4.60698
R31721 C10_P_btm.n1753 C10_P_btm.n1752 4.60698
R31722 C10_P_btm.n1752 C10_P_btm.n1751 4.60698
R31723 C10_P_btm.n1756 C10_P_btm.n1755 4.60698
R31724 C10_P_btm.n1755 C10_P_btm.n1754 4.60698
R31725 C10_P_btm.n1759 C10_P_btm.n1758 4.60698
R31726 C10_P_btm.n1758 C10_P_btm.n1757 4.60698
R31727 C10_P_btm.n1762 C10_P_btm.n1761 4.60698
R31728 C10_P_btm.n1761 C10_P_btm.n1760 4.60698
R31729 C10_P_btm.n1765 C10_P_btm.n1764 4.60698
R31730 C10_P_btm.n1764 C10_P_btm.n1763 4.60698
R31731 C10_P_btm.n1768 C10_P_btm.n1767 4.60698
R31732 C10_P_btm.n1767 C10_P_btm.n1766 4.60698
R31733 C10_P_btm.n1771 C10_P_btm.n1770 4.60698
R31734 C10_P_btm.n1770 C10_P_btm.n1769 4.60698
R31735 C10_P_btm.n1774 C10_P_btm.n1773 4.60698
R31736 C10_P_btm.n1773 C10_P_btm.n1772 4.60698
R31737 C10_P_btm.n1777 C10_P_btm.n1776 4.60698
R31738 C10_P_btm.n1776 C10_P_btm.n1775 4.60698
R31739 C10_P_btm.n1780 C10_P_btm.n1779 4.60698
R31740 C10_P_btm.n1779 C10_P_btm.n1778 4.60698
R31741 C10_P_btm.n1783 C10_P_btm.n1782 4.60698
R31742 C10_P_btm.n1782 C10_P_btm.n1781 4.60698
R31743 C10_P_btm.n1786 C10_P_btm.n1785 4.60698
R31744 C10_P_btm.n1785 C10_P_btm.n1784 4.60698
R31745 C10_P_btm.n1789 C10_P_btm.n1788 4.60698
R31746 C10_P_btm.n1788 C10_P_btm.n1787 4.60698
R31747 C10_P_btm.n1792 C10_P_btm.n1791 4.60698
R31748 C10_P_btm.n1791 C10_P_btm.n1790 4.60698
R31749 C10_P_btm.n1795 C10_P_btm.n1794 4.60698
R31750 C10_P_btm.n1794 C10_P_btm.n1793 4.60698
R31751 C10_P_btm.n1798 C10_P_btm.n1797 4.60698
R31752 C10_P_btm.n1797 C10_P_btm.n1796 4.60698
R31753 C10_P_btm.n1801 C10_P_btm.n1800 4.60698
R31754 C10_P_btm.n1800 C10_P_btm.n1799 4.60698
R31755 C10_P_btm.n1804 C10_P_btm.n1803 4.60698
R31756 C10_P_btm.n1803 C10_P_btm.n1802 4.60698
R31757 C10_P_btm.n1807 C10_P_btm.n1806 4.60698
R31758 C10_P_btm.n1806 C10_P_btm.n1805 4.60698
R31759 C10_P_btm.n1810 C10_P_btm.n1809 4.60698
R31760 C10_P_btm.n1809 C10_P_btm.n1808 4.60698
R31761 C10_P_btm.n1813 C10_P_btm.n1812 4.60698
R31762 C10_P_btm.n1812 C10_P_btm.n1811 4.60698
R31763 C10_P_btm.n1816 C10_P_btm.n1815 4.60698
R31764 C10_P_btm.n1815 C10_P_btm.n1814 4.60698
R31765 C10_P_btm.n1819 C10_P_btm.n1818 4.60698
R31766 C10_P_btm.n1818 C10_P_btm.n1817 4.60698
R31767 C10_P_btm.n1822 C10_P_btm.n1821 4.60698
R31768 C10_P_btm.n1821 C10_P_btm.n1820 4.60698
R31769 C10_P_btm.n1825 C10_P_btm.n1824 4.60698
R31770 C10_P_btm.n1824 C10_P_btm.n1823 4.60698
R31771 C10_P_btm.n1828 C10_P_btm.n1827 4.60698
R31772 C10_P_btm.n1827 C10_P_btm.n1826 4.60698
R31773 C10_P_btm.n1831 C10_P_btm.n1830 4.60698
R31774 C10_P_btm.n1830 C10_P_btm.n1829 4.60698
R31775 C10_P_btm.n1834 C10_P_btm.n1833 4.60698
R31776 C10_P_btm.n1833 C10_P_btm.n1832 4.60698
R31777 C10_P_btm.n1837 C10_P_btm.n1836 4.60698
R31778 C10_P_btm.n1836 C10_P_btm.n1835 4.60698
R31779 C10_P_btm.n1840 C10_P_btm.n1839 4.60698
R31780 C10_P_btm.n1839 C10_P_btm.n1838 4.60698
R31781 C10_P_btm.n1843 C10_P_btm.n1842 4.60698
R31782 C10_P_btm.n1842 C10_P_btm.n1841 4.60698
R31783 C10_P_btm.n1846 C10_P_btm.n1845 4.60698
R31784 C10_P_btm.n1845 C10_P_btm.n1844 4.60698
R31785 C10_P_btm.n1849 C10_P_btm.n1848 4.60698
R31786 C10_P_btm.n1848 C10_P_btm.n1847 4.60698
R31787 C10_P_btm.n1852 C10_P_btm.n1851 4.60698
R31788 C10_P_btm.n1851 C10_P_btm.n1850 4.60698
R31789 C10_P_btm.n1855 C10_P_btm.n1854 4.60698
R31790 C10_P_btm.n1854 C10_P_btm.n1853 4.60698
R31791 C10_P_btm.n1858 C10_P_btm.n1857 4.60698
R31792 C10_P_btm.n1857 C10_P_btm.n1856 4.60698
R31793 C10_P_btm.n1484 C10_P_btm.n1483 4.60698
R31794 C10_P_btm.n1485 C10_P_btm.n1484 4.60698
R31795 C10_P_btm.n1487 C10_P_btm.n1486 4.60698
R31796 C10_P_btm.n1488 C10_P_btm.n1487 4.60698
R31797 C10_P_btm.n1490 C10_P_btm.n1489 4.60698
R31798 C10_P_btm.n1491 C10_P_btm.n1490 4.60698
R31799 C10_P_btm.n1493 C10_P_btm.n1492 4.60698
R31800 C10_P_btm.n1494 C10_P_btm.n1493 4.60698
R31801 C10_P_btm.n1496 C10_P_btm.n1495 4.60698
R31802 C10_P_btm.n1497 C10_P_btm.n1496 4.60698
R31803 C10_P_btm.n1499 C10_P_btm.n1498 4.60698
R31804 C10_P_btm.n1500 C10_P_btm.n1499 4.60698
R31805 C10_P_btm.n1502 C10_P_btm.n1501 4.60698
R31806 C10_P_btm.n1503 C10_P_btm.n1502 4.60698
R31807 C10_P_btm.n1505 C10_P_btm.n1504 4.60698
R31808 C10_P_btm.n1506 C10_P_btm.n1505 4.60698
R31809 C10_P_btm.n1508 C10_P_btm.n1507 4.60698
R31810 C10_P_btm.n1509 C10_P_btm.n1508 4.60698
R31811 C10_P_btm.n1511 C10_P_btm.n1510 4.60698
R31812 C10_P_btm.n1512 C10_P_btm.n1511 4.60698
R31813 C10_P_btm.n1514 C10_P_btm.n1513 4.60698
R31814 C10_P_btm.n1515 C10_P_btm.n1514 4.60698
R31815 C10_P_btm.n1517 C10_P_btm.n1516 4.60698
R31816 C10_P_btm.n1518 C10_P_btm.n1517 4.60698
R31817 C10_P_btm.n1520 C10_P_btm.n1519 4.60698
R31818 C10_P_btm.n1521 C10_P_btm.n1520 4.60698
R31819 C10_P_btm.n1523 C10_P_btm.n1522 4.60698
R31820 C10_P_btm.n1524 C10_P_btm.n1523 4.60698
R31821 C10_P_btm.n1526 C10_P_btm.n1525 4.60698
R31822 C10_P_btm.n1527 C10_P_btm.n1526 4.60698
R31823 C10_P_btm.n1529 C10_P_btm.n1528 4.60698
R31824 C10_P_btm.n1530 C10_P_btm.n1529 4.60698
R31825 C10_P_btm.n1532 C10_P_btm.n1531 4.60698
R31826 C10_P_btm.n1533 C10_P_btm.n1532 4.60698
R31827 C10_P_btm.n1535 C10_P_btm.n1534 4.60698
R31828 C10_P_btm.n1536 C10_P_btm.n1535 4.60698
R31829 C10_P_btm.n1538 C10_P_btm.n1537 4.60698
R31830 C10_P_btm.n1539 C10_P_btm.n1538 4.60698
R31831 C10_P_btm.n1541 C10_P_btm.n1540 4.60698
R31832 C10_P_btm.n1542 C10_P_btm.n1541 4.60698
R31833 C10_P_btm.n1544 C10_P_btm.n1543 4.60698
R31834 C10_P_btm.n1545 C10_P_btm.n1544 4.60698
R31835 C10_P_btm.n1547 C10_P_btm.n1546 4.60698
R31836 C10_P_btm.n1548 C10_P_btm.n1547 4.60698
R31837 C10_P_btm.n1550 C10_P_btm.n1549 4.60698
R31838 C10_P_btm.n1551 C10_P_btm.n1550 4.60698
R31839 C10_P_btm.n1553 C10_P_btm.n1552 4.60698
R31840 C10_P_btm.n1554 C10_P_btm.n1553 4.60698
R31841 C10_P_btm.n1556 C10_P_btm.n1555 4.60698
R31842 C10_P_btm.n1557 C10_P_btm.n1556 4.60698
R31843 C10_P_btm.n1559 C10_P_btm.n1558 4.60698
R31844 C10_P_btm.n1560 C10_P_btm.n1559 4.60698
R31845 C10_P_btm.n1562 C10_P_btm.n1561 4.60698
R31846 C10_P_btm.n1563 C10_P_btm.n1562 4.60698
R31847 C10_P_btm.n1565 C10_P_btm.n1564 4.60698
R31848 C10_P_btm.n1566 C10_P_btm.n1565 4.60698
R31849 C10_P_btm.n1568 C10_P_btm.n1567 4.60698
R31850 C10_P_btm.n1569 C10_P_btm.n1568 4.60698
R31851 C10_P_btm.n1571 C10_P_btm.n1570 4.60698
R31852 C10_P_btm.n1572 C10_P_btm.n1571 4.60698
R31853 C10_P_btm.n1574 C10_P_btm.n1573 4.60698
R31854 C10_P_btm.n1575 C10_P_btm.n1574 4.60698
R31855 C10_P_btm.n1577 C10_P_btm.n1576 4.60698
R31856 C10_P_btm.n1578 C10_P_btm.n1577 4.60698
R31857 C10_P_btm.n1580 C10_P_btm.n1579 4.60698
R31858 C10_P_btm.n1581 C10_P_btm.n1580 4.60698
R31859 C10_P_btm.n1583 C10_P_btm.n1582 4.60698
R31860 C10_P_btm.n1584 C10_P_btm.n1583 4.60698
R31861 C10_P_btm.n1586 C10_P_btm.n1585 4.60698
R31862 C10_P_btm.n1587 C10_P_btm.n1586 4.60698
R31863 C10_P_btm.n1589 C10_P_btm.n1588 4.60698
R31864 C10_P_btm.n1590 C10_P_btm.n1589 4.60698
R31865 C10_P_btm.n1592 C10_P_btm.n1591 4.60698
R31866 C10_P_btm.n1593 C10_P_btm.n1592 4.60698
R31867 C10_P_btm.n1595 C10_P_btm.n1594 4.60698
R31868 C10_P_btm.n1596 C10_P_btm.n1595 4.60698
R31869 C10_P_btm.n1598 C10_P_btm.n1597 4.60698
R31870 C10_P_btm.n1599 C10_P_btm.n1598 4.60698
R31871 C10_P_btm.n1601 C10_P_btm.n1600 4.60698
R31872 C10_P_btm.n1602 C10_P_btm.n1601 4.60698
R31873 C10_P_btm.n1604 C10_P_btm.n1603 4.60698
R31874 C10_P_btm.n1605 C10_P_btm.n1604 4.60698
R31875 C10_P_btm.n1607 C10_P_btm.n1606 4.60698
R31876 C10_P_btm.n1608 C10_P_btm.n1607 4.60698
R31877 C10_P_btm.n1610 C10_P_btm.n1609 4.60698
R31878 C10_P_btm.n1611 C10_P_btm.n1610 4.60698
R31879 C10_P_btm.n1613 C10_P_btm.n1612 4.60698
R31880 C10_P_btm.n1614 C10_P_btm.n1613 4.60698
R31881 C10_P_btm.n1616 C10_P_btm.n1615 4.60698
R31882 C10_P_btm.n1617 C10_P_btm.n1616 4.60698
R31883 C10_P_btm.n1619 C10_P_btm.n1618 4.60698
R31884 C10_P_btm.n1620 C10_P_btm.n1619 4.60698
R31885 C10_P_btm.n1622 C10_P_btm.n1621 4.60698
R31886 C10_P_btm.n1623 C10_P_btm.n1622 4.60698
R31887 C10_P_btm.n1625 C10_P_btm.n1624 4.60698
R31888 C10_P_btm.n1626 C10_P_btm.n1625 4.60698
R31889 C10_P_btm.n1628 C10_P_btm.n1627 4.60698
R31890 C10_P_btm.n1629 C10_P_btm.n1628 4.60698
R31891 C10_P_btm.n1631 C10_P_btm.n1630 4.60698
R31892 C10_P_btm.n1632 C10_P_btm.n1631 4.60698
R31893 C10_P_btm.n1634 C10_P_btm.n1633 4.60698
R31894 C10_P_btm.n1635 C10_P_btm.n1634 4.60698
R31895 C10_P_btm.n1637 C10_P_btm.n1636 4.60698
R31896 C10_P_btm.n1638 C10_P_btm.n1637 4.60698
R31897 C10_P_btm.n1640 C10_P_btm.n1639 4.60698
R31898 C10_P_btm.n1641 C10_P_btm.n1640 4.60698
R31899 C10_P_btm.n1643 C10_P_btm.n1642 4.60698
R31900 C10_P_btm.n1644 C10_P_btm.n1643 4.60698
R31901 C10_P_btm.n1646 C10_P_btm.n1645 4.60698
R31902 C10_P_btm.n1647 C10_P_btm.n1646 4.60698
R31903 C10_P_btm.n1649 C10_P_btm.n1648 4.60698
R31904 C10_P_btm.n1650 C10_P_btm.n1649 4.60698
R31905 C10_P_btm.n1652 C10_P_btm.n1651 4.60698
R31906 C10_P_btm.n1653 C10_P_btm.n1652 4.60698
R31907 C10_P_btm.n1655 C10_P_btm.n1654 4.60698
R31908 C10_P_btm.n1656 C10_P_btm.n1655 4.60698
R31909 C10_P_btm.n1658 C10_P_btm.n1657 4.60698
R31910 C10_P_btm.n1659 C10_P_btm.n1658 4.60698
R31911 C10_P_btm.n1661 C10_P_btm.n1660 4.60698
R31912 C10_P_btm.n1662 C10_P_btm.n1661 4.60698
R31913 C10_P_btm.n1664 C10_P_btm.n1663 4.60698
R31914 C10_P_btm.n1665 C10_P_btm.n1664 4.60698
R31915 C10_P_btm.n1667 C10_P_btm.n1666 4.60698
R31916 C10_P_btm.n1668 C10_P_btm.n1667 4.60698
R31917 C10_P_btm.n1285 C10_P_btm.n1284 4.60698
R31918 C10_P_btm.n1284 C10_P_btm.n1043 4.60698
R31919 C10_P_btm.n1282 C10_P_btm.n1281 4.60698
R31920 C10_P_btm.n1283 C10_P_btm.n1282 4.60698
R31921 C10_P_btm.n1279 C10_P_btm.n1278 4.60698
R31922 C10_P_btm.n1280 C10_P_btm.n1279 4.60698
R31923 C10_P_btm.n1276 C10_P_btm.n1275 4.60698
R31924 C10_P_btm.n1277 C10_P_btm.n1276 4.60698
R31925 C10_P_btm.n1273 C10_P_btm.n1272 4.60698
R31926 C10_P_btm.n1274 C10_P_btm.n1273 4.60698
R31927 C10_P_btm.n1270 C10_P_btm.n1269 4.60698
R31928 C10_P_btm.n1271 C10_P_btm.n1270 4.60698
R31929 C10_P_btm.n1267 C10_P_btm.n1266 4.60698
R31930 C10_P_btm.n1268 C10_P_btm.n1267 4.60698
R31931 C10_P_btm.n1264 C10_P_btm.n1263 4.60698
R31932 C10_P_btm.n1265 C10_P_btm.n1264 4.60698
R31933 C10_P_btm.n1261 C10_P_btm.n1260 4.60698
R31934 C10_P_btm.n1262 C10_P_btm.n1261 4.60698
R31935 C10_P_btm.n1258 C10_P_btm.n1257 4.60698
R31936 C10_P_btm.n1259 C10_P_btm.n1258 4.60698
R31937 C10_P_btm.n1255 C10_P_btm.n1254 4.60698
R31938 C10_P_btm.n1256 C10_P_btm.n1255 4.60698
R31939 C10_P_btm.n1252 C10_P_btm.n1251 4.60698
R31940 C10_P_btm.n1253 C10_P_btm.n1252 4.60698
R31941 C10_P_btm.n1249 C10_P_btm.n1248 4.60698
R31942 C10_P_btm.n1250 C10_P_btm.n1249 4.60698
R31943 C10_P_btm.n1246 C10_P_btm.n1245 4.60698
R31944 C10_P_btm.n1247 C10_P_btm.n1246 4.60698
R31945 C10_P_btm.n1243 C10_P_btm.n1242 4.60698
R31946 C10_P_btm.n1244 C10_P_btm.n1243 4.60698
R31947 C10_P_btm.n1240 C10_P_btm.n1239 4.60698
R31948 C10_P_btm.n1241 C10_P_btm.n1240 4.60698
R31949 C10_P_btm.n1237 C10_P_btm.n1236 4.60698
R31950 C10_P_btm.n1238 C10_P_btm.n1237 4.60698
R31951 C10_P_btm.n1234 C10_P_btm.n1233 4.60698
R31952 C10_P_btm.n1235 C10_P_btm.n1234 4.60698
R31953 C10_P_btm.n1231 C10_P_btm.n1230 4.60698
R31954 C10_P_btm.n1232 C10_P_btm.n1231 4.60698
R31955 C10_P_btm.n1228 C10_P_btm.n1227 4.60698
R31956 C10_P_btm.n1229 C10_P_btm.n1228 4.60698
R31957 C10_P_btm.n1225 C10_P_btm.n1224 4.60698
R31958 C10_P_btm.n1226 C10_P_btm.n1225 4.60698
R31959 C10_P_btm.n1222 C10_P_btm.n1221 4.60698
R31960 C10_P_btm.n1223 C10_P_btm.n1222 4.60698
R31961 C10_P_btm.n1219 C10_P_btm.n1218 4.60698
R31962 C10_P_btm.n1220 C10_P_btm.n1219 4.60698
R31963 C10_P_btm.n1216 C10_P_btm.n1215 4.60698
R31964 C10_P_btm.n1217 C10_P_btm.n1216 4.60698
R31965 C10_P_btm.n1213 C10_P_btm.n1212 4.60698
R31966 C10_P_btm.n1214 C10_P_btm.n1213 4.60698
R31967 C10_P_btm.n1210 C10_P_btm.n1209 4.60698
R31968 C10_P_btm.n1211 C10_P_btm.n1210 4.60698
R31969 C10_P_btm.n1207 C10_P_btm.n1206 4.60698
R31970 C10_P_btm.n1208 C10_P_btm.n1207 4.60698
R31971 C10_P_btm.n1204 C10_P_btm.n1203 4.60698
R31972 C10_P_btm.n1205 C10_P_btm.n1204 4.60698
R31973 C10_P_btm.n1201 C10_P_btm.n1200 4.60698
R31974 C10_P_btm.n1202 C10_P_btm.n1201 4.60698
R31975 C10_P_btm.n1198 C10_P_btm.n1197 4.60698
R31976 C10_P_btm.n1199 C10_P_btm.n1198 4.60698
R31977 C10_P_btm.n1195 C10_P_btm.n1194 4.60698
R31978 C10_P_btm.n1196 C10_P_btm.n1195 4.60698
R31979 C10_P_btm.n1192 C10_P_btm.n1191 4.60698
R31980 C10_P_btm.n1193 C10_P_btm.n1192 4.60698
R31981 C10_P_btm.n1189 C10_P_btm.n1188 4.60698
R31982 C10_P_btm.n1190 C10_P_btm.n1189 4.60698
R31983 C10_P_btm.n1186 C10_P_btm.n1185 4.60698
R31984 C10_P_btm.n1187 C10_P_btm.n1186 4.60698
R31985 C10_P_btm.n1183 C10_P_btm.n1182 4.60698
R31986 C10_P_btm.n1184 C10_P_btm.n1183 4.60698
R31987 C10_P_btm.n1180 C10_P_btm.n1179 4.60698
R31988 C10_P_btm.n1181 C10_P_btm.n1180 4.60698
R31989 C10_P_btm.n1177 C10_P_btm.n1176 4.60698
R31990 C10_P_btm.n1178 C10_P_btm.n1177 4.60698
R31991 C10_P_btm.n1174 C10_P_btm.n1173 4.60698
R31992 C10_P_btm.n1175 C10_P_btm.n1174 4.60698
R31993 C10_P_btm.n1171 C10_P_btm.n1170 4.60698
R31994 C10_P_btm.n1172 C10_P_btm.n1171 4.60698
R31995 C10_P_btm.n1168 C10_P_btm.n1167 4.60698
R31996 C10_P_btm.n1169 C10_P_btm.n1168 4.60698
R31997 C10_P_btm.n1165 C10_P_btm.n1164 4.60698
R31998 C10_P_btm.n1166 C10_P_btm.n1165 4.60698
R31999 C10_P_btm.n1162 C10_P_btm.n1161 4.60698
R32000 C10_P_btm.n1163 C10_P_btm.n1162 4.60698
R32001 C10_P_btm.n1159 C10_P_btm.n1158 4.60698
R32002 C10_P_btm.n1160 C10_P_btm.n1159 4.60698
R32003 C10_P_btm.n1156 C10_P_btm.n1155 4.60698
R32004 C10_P_btm.n1157 C10_P_btm.n1156 4.60698
R32005 C10_P_btm.n1153 C10_P_btm.n1152 4.60698
R32006 C10_P_btm.n1154 C10_P_btm.n1153 4.60698
R32007 C10_P_btm.n1150 C10_P_btm.n1149 4.60698
R32008 C10_P_btm.n1151 C10_P_btm.n1150 4.60698
R32009 C10_P_btm.n1147 C10_P_btm.n1146 4.60698
R32010 C10_P_btm.n1148 C10_P_btm.n1147 4.60698
R32011 C10_P_btm.n1144 C10_P_btm.n1143 4.60698
R32012 C10_P_btm.n1145 C10_P_btm.n1144 4.60698
R32013 C10_P_btm.n1141 C10_P_btm.n1140 4.60698
R32014 C10_P_btm.n1142 C10_P_btm.n1141 4.60698
R32015 C10_P_btm.n1138 C10_P_btm.n1137 4.60698
R32016 C10_P_btm.n1139 C10_P_btm.n1138 4.60698
R32017 C10_P_btm.n1135 C10_P_btm.n1134 4.60698
R32018 C10_P_btm.n1136 C10_P_btm.n1135 4.60698
R32019 C10_P_btm.n1132 C10_P_btm.n1131 4.60698
R32020 C10_P_btm.n1133 C10_P_btm.n1132 4.60698
R32021 C10_P_btm.n1129 C10_P_btm.n1128 4.60698
R32022 C10_P_btm.n1130 C10_P_btm.n1129 4.60698
R32023 C10_P_btm.n1126 C10_P_btm.n1125 4.60698
R32024 C10_P_btm.n1127 C10_P_btm.n1126 4.60698
R32025 C10_P_btm.n1123 C10_P_btm.n1122 4.60698
R32026 C10_P_btm.n1124 C10_P_btm.n1123 4.60698
R32027 C10_P_btm.n1120 C10_P_btm.n1119 4.60698
R32028 C10_P_btm.n1121 C10_P_btm.n1120 4.60698
R32029 C10_P_btm.n1117 C10_P_btm.n1116 4.60698
R32030 C10_P_btm.n1118 C10_P_btm.n1117 4.60698
R32031 C10_P_btm.n1114 C10_P_btm.n1113 4.60698
R32032 C10_P_btm.n1115 C10_P_btm.n1114 4.60698
R32033 C10_P_btm.n1111 C10_P_btm.n1110 4.60698
R32034 C10_P_btm.n1112 C10_P_btm.n1111 4.60698
R32035 C10_P_btm.n1108 C10_P_btm.n1107 4.60698
R32036 C10_P_btm.n1109 C10_P_btm.n1108 4.60698
R32037 C10_P_btm.n1105 C10_P_btm.n1104 4.60698
R32038 C10_P_btm.n1106 C10_P_btm.n1105 4.60698
R32039 C10_P_btm.n1479 C10_P_btm.n1478 4.60698
R32040 C10_P_btm.n1478 C10_P_btm.n981 4.60698
R32041 C10_P_btm.n1474 C10_P_btm.n1473 4.60698
R32042 C10_P_btm.n1473 C10_P_btm.n1472 4.60698
R32043 C10_P_btm.n1471 C10_P_btm.n1470 4.60698
R32044 C10_P_btm.n1470 C10_P_btm.n1469 4.60698
R32045 C10_P_btm.n1468 C10_P_btm.n1467 4.60698
R32046 C10_P_btm.n1467 C10_P_btm.n1466 4.60698
R32047 C10_P_btm.n1465 C10_P_btm.n1464 4.60698
R32048 C10_P_btm.n1464 C10_P_btm.n1463 4.60698
R32049 C10_P_btm.n1462 C10_P_btm.n1461 4.60698
R32050 C10_P_btm.n1461 C10_P_btm.n1460 4.60698
R32051 C10_P_btm.n1459 C10_P_btm.n1458 4.60698
R32052 C10_P_btm.n1458 C10_P_btm.n1457 4.60698
R32053 C10_P_btm.n1456 C10_P_btm.n1455 4.60698
R32054 C10_P_btm.n1455 C10_P_btm.n1454 4.60698
R32055 C10_P_btm.n1453 C10_P_btm.n1452 4.60698
R32056 C10_P_btm.n1452 C10_P_btm.n1451 4.60698
R32057 C10_P_btm.n1450 C10_P_btm.n1449 4.60698
R32058 C10_P_btm.n1449 C10_P_btm.n1448 4.60698
R32059 C10_P_btm.n1447 C10_P_btm.n1446 4.60698
R32060 C10_P_btm.n1446 C10_P_btm.n1445 4.60698
R32061 C10_P_btm.n1444 C10_P_btm.n1443 4.60698
R32062 C10_P_btm.n1443 C10_P_btm.n1442 4.60698
R32063 C10_P_btm.n1441 C10_P_btm.n1440 4.60698
R32064 C10_P_btm.n1440 C10_P_btm.n1439 4.60698
R32065 C10_P_btm.n1438 C10_P_btm.n1437 4.60698
R32066 C10_P_btm.n1437 C10_P_btm.n1436 4.60698
R32067 C10_P_btm.n1435 C10_P_btm.n1434 4.60698
R32068 C10_P_btm.n1434 C10_P_btm.n1433 4.60698
R32069 C10_P_btm.n1432 C10_P_btm.n1431 4.60698
R32070 C10_P_btm.n1431 C10_P_btm.n1430 4.60698
R32071 C10_P_btm.n1429 C10_P_btm.n1428 4.60698
R32072 C10_P_btm.n1428 C10_P_btm.n1427 4.60698
R32073 C10_P_btm.n1426 C10_P_btm.n1425 4.60698
R32074 C10_P_btm.n1425 C10_P_btm.n1424 4.60698
R32075 C10_P_btm.n1423 C10_P_btm.n1422 4.60698
R32076 C10_P_btm.n1422 C10_P_btm.n1421 4.60698
R32077 C10_P_btm.n1420 C10_P_btm.n1419 4.60698
R32078 C10_P_btm.n1419 C10_P_btm.n1418 4.60698
R32079 C10_P_btm.n1417 C10_P_btm.n1416 4.60698
R32080 C10_P_btm.n1416 C10_P_btm.n1415 4.60698
R32081 C10_P_btm.n1414 C10_P_btm.n1413 4.60698
R32082 C10_P_btm.n1413 C10_P_btm.n1412 4.60698
R32083 C10_P_btm.n1411 C10_P_btm.n1410 4.60698
R32084 C10_P_btm.n1410 C10_P_btm.n1409 4.60698
R32085 C10_P_btm.n1408 C10_P_btm.n1407 4.60698
R32086 C10_P_btm.n1407 C10_P_btm.n1406 4.60698
R32087 C10_P_btm.n1405 C10_P_btm.n1404 4.60698
R32088 C10_P_btm.n1404 C10_P_btm.n1403 4.60698
R32089 C10_P_btm.n1402 C10_P_btm.n1401 4.60698
R32090 C10_P_btm.n1401 C10_P_btm.n1400 4.60698
R32091 C10_P_btm.n1399 C10_P_btm.n1398 4.60698
R32092 C10_P_btm.n1398 C10_P_btm.n1397 4.60698
R32093 C10_P_btm.n1396 C10_P_btm.n1395 4.60698
R32094 C10_P_btm.n1395 C10_P_btm.n1394 4.60698
R32095 C10_P_btm.n1393 C10_P_btm.n1392 4.60698
R32096 C10_P_btm.n1392 C10_P_btm.n1391 4.60698
R32097 C10_P_btm.n1390 C10_P_btm.n1389 4.60698
R32098 C10_P_btm.n1389 C10_P_btm.n1388 4.60698
R32099 C10_P_btm.n1387 C10_P_btm.n1386 4.60698
R32100 C10_P_btm.n1386 C10_P_btm.n1385 4.60698
R32101 C10_P_btm.n1384 C10_P_btm.n1383 4.60698
R32102 C10_P_btm.n1383 C10_P_btm.n1382 4.60698
R32103 C10_P_btm.n1381 C10_P_btm.n1380 4.60698
R32104 C10_P_btm.n1380 C10_P_btm.n1379 4.60698
R32105 C10_P_btm.n1378 C10_P_btm.n1377 4.60698
R32106 C10_P_btm.n1377 C10_P_btm.n1376 4.60698
R32107 C10_P_btm.n1375 C10_P_btm.n1374 4.60698
R32108 C10_P_btm.n1374 C10_P_btm.n1373 4.60698
R32109 C10_P_btm.n1372 C10_P_btm.n1371 4.60698
R32110 C10_P_btm.n1371 C10_P_btm.n1370 4.60698
R32111 C10_P_btm.n1369 C10_P_btm.n1368 4.60698
R32112 C10_P_btm.n1368 C10_P_btm.n1367 4.60698
R32113 C10_P_btm.n1366 C10_P_btm.n1365 4.60698
R32114 C10_P_btm.n1365 C10_P_btm.n1364 4.60698
R32115 C10_P_btm.n1363 C10_P_btm.n1362 4.60698
R32116 C10_P_btm.n1362 C10_P_btm.n1361 4.60698
R32117 C10_P_btm.n1360 C10_P_btm.n1359 4.60698
R32118 C10_P_btm.n1359 C10_P_btm.n1358 4.60698
R32119 C10_P_btm.n1357 C10_P_btm.n1356 4.60698
R32120 C10_P_btm.n1356 C10_P_btm.n1355 4.60698
R32121 C10_P_btm.n1354 C10_P_btm.n1353 4.60698
R32122 C10_P_btm.n1353 C10_P_btm.n1352 4.60698
R32123 C10_P_btm.n1351 C10_P_btm.n1350 4.60698
R32124 C10_P_btm.n1350 C10_P_btm.n1349 4.60698
R32125 C10_P_btm.n1348 C10_P_btm.n1347 4.60698
R32126 C10_P_btm.n1347 C10_P_btm.n1346 4.60698
R32127 C10_P_btm.n1345 C10_P_btm.n1344 4.60698
R32128 C10_P_btm.n1344 C10_P_btm.n1343 4.60698
R32129 C10_P_btm.n1342 C10_P_btm.n1341 4.60698
R32130 C10_P_btm.n1341 C10_P_btm.n1340 4.60698
R32131 C10_P_btm.n1339 C10_P_btm.n1338 4.60698
R32132 C10_P_btm.n1338 C10_P_btm.n1337 4.60698
R32133 C10_P_btm.n1336 C10_P_btm.n1335 4.60698
R32134 C10_P_btm.n1335 C10_P_btm.n1334 4.60698
R32135 C10_P_btm.n1333 C10_P_btm.n1332 4.60698
R32136 C10_P_btm.n1332 C10_P_btm.n1331 4.60698
R32137 C10_P_btm.n1330 C10_P_btm.n1329 4.60698
R32138 C10_P_btm.n1329 C10_P_btm.n1328 4.60698
R32139 C10_P_btm.n1327 C10_P_btm.n1326 4.60698
R32140 C10_P_btm.n1326 C10_P_btm.n1325 4.60698
R32141 C10_P_btm.n1324 C10_P_btm.n1323 4.60698
R32142 C10_P_btm.n1323 C10_P_btm.n1322 4.60698
R32143 C10_P_btm.n1321 C10_P_btm.n1320 4.60698
R32144 C10_P_btm.n1320 C10_P_btm.n1319 4.60698
R32145 C10_P_btm.n1318 C10_P_btm.n1317 4.60698
R32146 C10_P_btm.n1317 C10_P_btm.n1316 4.60698
R32147 C10_P_btm.n1315 C10_P_btm.n1314 4.60698
R32148 C10_P_btm.n1314 C10_P_btm.n1313 4.60698
R32149 C10_P_btm.n1312 C10_P_btm.n1311 4.60698
R32150 C10_P_btm.n1311 C10_P_btm.n1310 4.60698
R32151 C10_P_btm.n1309 C10_P_btm.n1308 4.60698
R32152 C10_P_btm.n1308 C10_P_btm.n1307 4.60698
R32153 C10_P_btm.n1306 C10_P_btm.n1305 4.60698
R32154 C10_P_btm.n1305 C10_P_btm.n1304 4.60698
R32155 C10_P_btm.n1303 C10_P_btm.n1302 4.60698
R32156 C10_P_btm.n1302 C10_P_btm.n1301 4.60698
R32157 C10_P_btm.n1300 C10_P_btm.n1299 4.60698
R32158 C10_P_btm.n1299 C10_P_btm.n1298 4.60698
R32159 C10_P_btm.n1297 C10_P_btm.n1296 4.60698
R32160 C10_P_btm.n1296 C10_P_btm.n1295 4.60698
R32161 C10_P_btm.n1294 C10_P_btm.n1293 4.60698
R32162 C10_P_btm.n1293 C10_P_btm.n1292 4.60698
R32163 C10_P_btm.n1291 C10_P_btm.n1290 4.60698
R32164 C10_P_btm.n1290 C10_P_btm.n1289 4.60698
R32165 C10_P_btm.n3897 C10_P_btm.t17 4.03712
R32166 C10_P_btm.n3895 C10_P_btm.t897 3.98193
R32167 C10_P_btm.n3867 C10_P_btm.t703 3.98193
R32168 C10_P_btm.n3836 C10_P_btm.t385 3.98193
R32169 C10_P_btm.n3735 C10_P_btm.t139 3.98193
R32170 C10_P_btm.n3768 C10_P_btm.t552 3.98193
R32171 C10_P_btm.n3771 C10_P_btm.t174 3.98193
R32172 C10_P_btm.n3733 C10_P_btm.t849 3.98193
R32173 C10_P_btm.n91 C10_P_btm.t340 3.98193
R32174 C10_P_btm.n3669 C10_P_btm.t1014 3.98193
R32175 C10_P_btm.n3666 C10_P_btm.t507 3.98193
R32176 C10_P_btm.n144 C10_P_btm.t122 3.98193
R32177 C10_P_btm.n3602 C10_P_btm.t804 3.98193
R32178 C10_P_btm.n3599 C10_P_btm.t286 3.98193
R32179 C10_P_btm.n197 C10_P_btm.t971 3.98193
R32180 C10_P_btm.n3535 C10_P_btm.t461 3.98193
R32181 C10_P_btm.n3532 C10_P_btm.t79 3.98193
R32182 C10_P_btm.n250 C10_P_btm.t751 3.98193
R32183 C10_P_btm.n3468 C10_P_btm.t868 3.98193
R32184 C10_P_btm.n3465 C10_P_btm.t920 3.98193
R32185 C10_P_btm.n303 C10_P_btm.t328 3.98193
R32186 C10_P_btm.n3401 C10_P_btm.t1008 3.98193
R32187 C10_P_btm.n3398 C10_P_btm.t310 3.98193
R32188 C10_P_btm.n356 C10_P_btm.t602 3.98193
R32189 C10_P_btm.n3334 C10_P_btm.t987 3.98193
R32190 C10_P_btm.n3331 C10_P_btm.t333 3.98193
R32191 C10_P_btm.n506 C10_P_btm.t885 3.98193
R32192 C10_P_btm.n3108 C10_P_btm.t241 3.98193
R32193 C10_P_btm.n3105 C10_P_btm.t129 3.98193
R32194 C10_P_btm.n2995 C10_P_btm.t51 3.98193
R32195 C10_P_btm.n2894 C10_P_btm.t375 3.98193
R32196 C10_P_btm.n2927 C10_P_btm.t277 3.98193
R32197 C10_P_btm.n2930 C10_P_btm.t415 3.98193
R32198 C10_P_btm.n2892 C10_P_btm.t1038 3.98193
R32199 C10_P_btm.n2114 C10_P_btm.t615 3.98193
R32200 C10_P_btm.n2828 C10_P_btm.t754 3.98193
R32201 C10_P_btm.n2825 C10_P_btm.t589 3.98193
R32202 C10_P_btm.n2167 C10_P_btm.t472 3.98193
R32203 C10_P_btm.n2761 C10_P_btm.t321 3.98193
R32204 C10_P_btm.n2758 C10_P_btm.t417 3.98193
R32205 C10_P_btm.n2220 C10_P_btm.t66 3.98193
R32206 C10_P_btm.n2694 C10_P_btm.t163 3.98193
R32207 C10_P_btm.n2691 C10_P_btm.t861 3.98193
R32208 C10_P_btm.n2273 C10_P_btm.t957 3.98193
R32209 C10_P_btm.n2627 C10_P_btm.t664 3.98193
R32210 C10_P_btm.n2624 C10_P_btm.t695 3.98193
R32211 C10_P_btm.n2326 C10_P_btm.t797 3.98193
R32212 C10_P_btm.n2560 C10_P_btm.t427 3.98193
R32213 C10_P_btm.n2557 C10_P_btm.t1054 3.98193
R32214 C10_P_btm.n2379 C10_P_btm.t628 3.98193
R32215 C10_P_btm.n2493 C10_P_btm.t257 3.98193
R32216 C10_P_btm.n2490 C10_P_btm.t353 3.98193
R32217 C10_P_btm.n2430 C10_P_btm.t464 3.98193
R32218 C10_P_btm.n2457 C10_P_btm.t872 3.98193
R32219 C10_P_btm.n2462 C10_P_btm.t170 3.98193
R32220 C10_P_btm.n2521 C10_P_btm.t73 3.98193
R32221 C10_P_btm.n2524 C10_P_btm.t426 3.98193
R32222 C10_P_btm.n2529 C10_P_btm.t329 3.98193
R32223 C10_P_btm.n2588 C10_P_btm.t494 3.98193
R32224 C10_P_btm.n2591 C10_P_btm.t596 3.98193
R32225 C10_P_btm.n2596 C10_P_btm.t1019 3.98193
R32226 C10_P_btm.n2655 C10_P_btm.t860 3.98193
R32227 C10_P_btm.n2658 C10_P_btm.t766 3.98193
R32228 C10_P_btm.n2663 C10_P_btm.t676 3.98193
R32229 C10_P_btm.n2722 C10_P_btm.t1026 3.98193
R32230 C10_P_btm.n2725 C10_P_btm.t933 3.98193
R32231 C10_P_btm.n2730 C10_P_btm.t469 3.98193
R32232 C10_P_btm.n2789 C10_P_btm.t133 3.98193
R32233 C10_P_btm.n2792 C10_P_btm.t107 3.98193
R32234 C10_P_btm.n2797 C10_P_btm.t394 3.98193
R32235 C10_P_btm.n2856 C10_P_btm.t295 3.98193
R32236 C10_P_btm.n2859 C10_P_btm.t413 3.98193
R32237 C10_P_btm.n2864 C10_P_btm.t319 3.98193
R32238 C10_P_btm.n2958 C10_P_btm.t245 3.98193
R32239 C10_P_btm.n2961 C10_P_btm.t98 3.98193
R32240 C10_P_btm.n2966 C10_P_btm.t184 3.98193
R32241 C10_P_btm.n3023 C10_P_btm.t911 3.98193
R32242 C10_P_btm.n3038 C10_P_btm.t592 3.98193
R32243 C10_P_btm.n2054 C10_P_btm.t930 3.98193
R32244 C10_P_btm.n672 C10_P_btm.t1023 3.98193
R32245 C10_P_btm.n1672 C10_P_btm.t672 3.98193
R32246 C10_P_btm.n1669 C10_P_btm.t761 3.98193
R32247 C10_P_btm.n1042 C10_P_btm.t857 3.98193
R32248 C10_P_btm.n1288 C10_P_btm.t859 3.98193
R32249 C10_P_btm.n1475 C10_P_btm.t402 3.98193
R32250 C10_P_btm.n1477 C10_P_btm.t968 3.98193
R32251 C10_P_btm.n1482 C10_P_btm.t576 3.98193
R32252 C10_P_btm.n1859 C10_P_btm.t189 3.98193
R32253 C10_P_btm.n1862 C10_P_btm.t749 3.98193
R32254 C10_P_btm.n1867 C10_P_btm.t360 3.98193
R32255 C10_P_btm.n3295 C10_P_btm.t919 3.98193
R32256 C10_P_btm.n3298 C10_P_btm.t526 3.98193
R32257 C10_P_btm.n3303 C10_P_btm.t145 3.98193
R32258 C10_P_btm.n3362 C10_P_btm.t802 3.98193
R32259 C10_P_btm.n3365 C10_P_btm.t404 3.98193
R32260 C10_P_btm.n3370 C10_P_btm.t432 3.98193
R32261 C10_P_btm.n3429 C10_P_btm.t822 3.98193
R32262 C10_P_btm.n3432 C10_P_btm.t140 3.98193
R32263 C10_P_btm.n3437 C10_P_btm.t734 3.98193
R32264 C10_P_btm.n3496 C10_P_btm.t1032 3.98193
R32265 C10_P_btm.n3499 C10_P_btm.t556 3.98193
R32266 C10_P_btm.n3504 C10_P_btm.t946 3.98193
R32267 C10_P_btm.n3563 C10_P_btm.t273 3.98193
R32268 C10_P_btm.n3566 C10_P_btm.t786 3.98193
R32269 C10_P_btm.n3571 C10_P_btm.t118 3.98193
R32270 C10_P_btm.n3630 C10_P_btm.t614 3.98193
R32271 C10_P_btm.n3633 C10_P_btm.t997 3.98193
R32272 C10_P_btm.n3638 C10_P_btm.t311 3.98193
R32273 C10_P_btm.n3697 C10_P_btm.t828 3.98193
R32274 C10_P_btm.n3700 C10_P_btm.t72 3.98193
R32275 C10_P_btm.n3705 C10_P_btm.t656 3.98193
R32276 C10_P_btm.n3799 C10_P_btm.t37 3.98193
R32277 C10_P_btm.n3802 C10_P_btm.t364 3.98193
R32278 C10_P_btm.n3807 C10_P_btm.t877 3.98193
R32279 C10_P_btm.n3864 C10_P_btm.t196 3.98193
R32280 C10_P_btm.n13 C10_P_btm.t1060 3.57113
R32281 C10_P_btm.n13 C10_P_btm.t1068 3.57113
R32282 C10_P_btm.n11 C10_P_btm.t1061 3.57113
R32283 C10_P_btm.n11 C10_P_btm.t1062 3.57113
R32284 C10_P_btm.n9 C10_P_btm.t1065 3.57113
R32285 C10_P_btm.n9 C10_P_btm.t1067 3.57113
R32286 C10_P_btm.n7 C10_P_btm.t1056 3.57113
R32287 C10_P_btm.n7 C10_P_btm.t1059 3.57113
R32288 C10_P_btm.n5 C10_P_btm.t1058 3.57113
R32289 C10_P_btm.n5 C10_P_btm.t1063 3.57113
R32290 C10_P_btm.n3 C10_P_btm.t1066 3.57113
R32291 C10_P_btm.n3 C10_P_btm.t1070 3.57113
R32292 C10_P_btm.n1 C10_P_btm.t1057 3.57113
R32293 C10_P_btm.n1 C10_P_btm.t1064 3.57113
R32294 C10_P_btm.n0 C10_P_btm.t1069 3.57113
R32295 C10_P_btm.n0 C10_P_btm.t1071 3.57113
R32296 C10_P_btm.n25 C10_P_btm.t1 2.4755
R32297 C10_P_btm.n25 C10_P_btm.t6 2.4755
R32298 C10_P_btm.n23 C10_P_btm.t8 2.4755
R32299 C10_P_btm.n23 C10_P_btm.t9 2.4755
R32300 C10_P_btm.n20 C10_P_btm.t1076 2.4755
R32301 C10_P_btm.n20 C10_P_btm.t1079 2.4755
R32302 C10_P_btm.n18 C10_P_btm.t1075 2.4755
R32303 C10_P_btm.n18 C10_P_btm.t1072 2.4755
R32304 C10_P_btm.n16 C10_P_btm.t1077 2.4755
R32305 C10_P_btm.n16 C10_P_btm.t1078 2.4755
R32306 C10_P_btm.n15 C10_P_btm.t1074 2.4755
R32307 C10_P_btm.n15 C10_P_btm.t1073 2.4755
R32308 C10_P_btm.n27 C10_P_btm.t5 2.4755
R32309 C10_P_btm.n27 C10_P_btm.t2 2.4755
R32310 C10_P_btm.n26 C10_P_btm.t7 2.4755
R32311 C10_P_btm.n26 C10_P_btm.t3 2.4755
R32312 C10_P_btm.n29 C10_P_btm.t0 2.4755
R32313 C10_P_btm.n29 C10_P_btm.t4 2.4755
R32314 C10_P_btm.n3893 C10_P_btm.t669 1.67819
R32315 C10_P_btm.n3890 C10_P_btm.t948 1.67819
R32316 C10_P_btm.n3887 C10_P_btm.t719 1.67819
R32317 C10_P_btm.n3884 C10_P_btm.t509 1.67819
R32318 C10_P_btm.n3881 C10_P_btm.t778 1.67819
R32319 C10_P_btm.n3878 C10_P_btm.t536 1.67819
R32320 C10_P_btm.n3875 C10_P_btm.t301 1.67819
R32321 C10_P_btm.n3872 C10_P_btm.t648 1.67819
R32322 C10_P_btm.n3869 C10_P_btm.t362 1.67819
R32323 C10_P_btm.n3862 C10_P_btm.t924 1.67819
R32324 C10_P_btm.n3859 C10_P_btm.t141 1.67819
R32325 C10_P_btm.n3856 C10_P_btm.t871 1.67819
R32326 C10_P_btm.n3853 C10_P_btm.t55 1.67819
R32327 C10_P_btm.n3850 C10_P_btm.t264 1.67819
R32328 C10_P_btm.n3847 C10_P_btm.t52 1.67819
R32329 C10_P_btm.n3844 C10_P_btm.t211 1.67819
R32330 C10_P_btm.n3841 C10_P_btm.t446 1.67819
R32331 C10_P_btm.n3838 C10_P_btm.t160 1.67819
R32332 C10_P_btm.n3832 C10_P_btm.t839 1.67819
R32333 C10_P_btm.n3830 C10_P_btm.t57 1.67819
R32334 C10_P_btm.n3827 C10_P_btm.t891 1.67819
R32335 C10_P_btm.n3824 C10_P_btm.t661 1.67819
R32336 C10_P_btm.n3821 C10_P_btm.t939 1.67819
R32337 C10_P_btm.n3818 C10_P_btm.t714 1.67819
R32338 C10_P_btm.n3815 C10_P_btm.t492 1.67819
R32339 C10_P_btm.n3812 C10_P_btm.t824 1.67819
R32340 C10_P_btm.n3809 C10_P_btm.t530 1.67819
R32341 C10_P_btm.n3803 C10_P_btm.t40 1.67819
R32342 C10_P_btm.n3745 C10_P_btm.t303 1.67819
R32343 C10_P_btm.n3748 C10_P_btm.t94 1.67819
R32344 C10_P_btm.n3751 C10_P_btm.t205 1.67819
R32345 C10_P_btm.n3754 C10_P_btm.t438 1.67819
R32346 C10_P_btm.n3757 C10_P_btm.t153 1.67819
R32347 C10_P_btm.n3760 C10_P_btm.t381 1.67819
R32348 C10_P_btm.n3763 C10_P_btm.t619 1.67819
R32349 C10_P_btm.n3766 C10_P_btm.t322 1.67819
R32350 C10_P_btm.n3773 C10_P_btm.t1005 1.67819
R32351 C10_P_btm.n3776 C10_P_btm.t240 1.67819
R32352 C10_P_btm.n3779 C10_P_btm.t1010 1.67819
R32353 C10_P_btm.n3782 C10_P_btm.t832 1.67819
R32354 C10_P_btm.n3785 C10_P_btm.t243 1.67819
R32355 C10_P_btm.n3788 C10_P_btm.t884 1.67819
R32356 C10_P_btm.n3791 C10_P_btm.t652 1.67819
R32357 C10_P_btm.n3794 C10_P_btm.t988 1.67819
R32358 C10_P_btm.n3797 C10_P_btm.t706 1.67819
R32359 C10_P_btm.n3707 C10_P_btm.t151 1.67819
R32360 C10_P_btm.n3710 C10_P_btm.t603 1.67819
R32361 C10_P_btm.n3713 C10_P_btm.t260 1.67819
R32362 C10_P_btm.n3716 C10_P_btm.t699 1.67819
R32363 C10_P_btm.n3719 C10_P_btm.t728 1.67819
R32364 C10_P_btm.n3722 C10_P_btm.t444 1.67819
R32365 C10_P_btm.n3725 C10_P_btm.t675 1.67819
R32366 C10_P_btm.n3728 C10_P_btm.t905 1.67819
R32367 C10_P_btm.n3731 C10_P_btm.t625 1.67819
R32368 C10_P_btm.n121 C10_P_btm.t483 1.67819
R32369 C10_P_btm.n119 C10_P_btm.t390 1.67819
R32370 C10_P_btm.n116 C10_P_btm.t169 1.67819
R32371 C10_P_btm.n113 C10_P_btm.t1001 1.67819
R32372 C10_P_btm.n110 C10_P_btm.t230 1.67819
R32373 C10_P_btm.n107 C10_P_btm.t894 1.67819
R32374 C10_P_btm.n104 C10_P_btm.t826 1.67819
R32375 C10_P_btm.n101 C10_P_btm.t111 1.67819
R32376 C10_P_btm.n3701 C10_P_btm.t878 1.67819
R32377 C10_P_btm.n3695 C10_P_btm.t500 1.67819
R32378 C10_P_btm.n3692 C10_P_btm.t775 1.67819
R32379 C10_P_btm.n3689 C10_P_btm.t435 1.67819
R32380 C10_P_btm.n3686 C10_P_btm.t668 1.67819
R32381 C10_P_btm.n3683 C10_P_btm.t896 1.67819
R32382 C10_P_btm.n3680 C10_P_btm.t617 1.67819
R32383 C10_P_btm.n3677 C10_P_btm.t844 1.67819
R32384 C10_P_btm.n3674 C10_P_btm.t64 1.67819
R32385 C10_P_btm.n3671 C10_P_btm.t796 1.67819
R32386 C10_P_btm.n3664 C10_P_btm.t276 1.67819
R32387 C10_P_btm.n3661 C10_P_btm.t562 1.67819
R32388 C10_P_btm.n3658 C10_P_btm.t330 1.67819
R32389 C10_P_btm.n3655 C10_P_btm.t224 1.67819
R32390 C10_P_btm.n3652 C10_P_btm.t1042 1.67819
R32391 C10_P_btm.n3649 C10_P_btm.t159 1.67819
R32392 C10_P_btm.n3646 C10_P_btm.t990 1.67819
R32393 C10_P_btm.n3643 C10_P_btm.t261 1.67819
R32394 C10_P_btm.n3640 C10_P_btm.t49 1.67819
R32395 C10_P_btm.n3634 C10_P_btm.t659 1.67819
R32396 C10_P_btm.n154 C10_P_btm.t938 1.67819
R32397 C10_P_btm.n157 C10_P_btm.t606 1.67819
R32398 C10_P_btm.n160 C10_P_btm.t837 1.67819
R32399 C10_P_btm.n163 C10_P_btm.t266 1.67819
R32400 C10_P_btm.n166 C10_P_btm.t789 1.67819
R32401 C10_P_btm.n169 C10_P_btm.t1012 1.67819
R32402 C10_P_btm.n172 C10_P_btm.t179 1.67819
R32403 C10_P_btm.n174 C10_P_btm.t956 1.67819
R32404 C10_P_btm.n3604 C10_P_btm.t566 1.67819
R32405 C10_P_btm.n3607 C10_P_btm.t854 1.67819
R32406 C10_P_btm.n3610 C10_P_btm.t632 1.67819
R32407 C10_P_btm.n3613 C10_P_btm.t1049 1.67819
R32408 C10_P_btm.n3616 C10_P_btm.t684 1.67819
R32409 C10_P_btm.n3619 C10_P_btm.t452 1.67819
R32410 C10_P_btm.n3622 C10_P_btm.t223 1.67819
R32411 C10_P_btm.n3625 C10_P_btm.t549 1.67819
R32412 C10_P_btm.n3628 C10_P_btm.t271 1.67819
R32413 C10_P_btm.n3573 C10_P_btm.t831 1.67819
R32414 C10_P_btm.n3576 C10_P_btm.t228 1.67819
R32415 C10_P_btm.n3579 C10_P_btm.t779 1.67819
R32416 C10_P_btm.n3582 C10_P_btm.t1004 1.67819
R32417 C10_P_btm.n3585 C10_P_btm.t173 1.67819
R32418 C10_P_btm.n3588 C10_P_btm.t949 1.67819
R32419 C10_P_btm.n3591 C10_P_btm.t631 1.67819
R32420 C10_P_btm.n3594 C10_P_btm.t346 1.67819
R32421 C10_P_btm.n3597 C10_P_btm.t65 1.67819
R32422 C10_P_btm.n227 C10_P_btm.t740 1.67819
R32423 C10_P_btm.n225 C10_P_btm.t1020 1.67819
R32424 C10_P_btm.n222 C10_P_btm.t800 1.67819
R32425 C10_P_btm.n219 C10_P_btm.t558 1.67819
R32426 C10_P_btm.n216 C10_P_btm.t848 1.67819
R32427 C10_P_btm.n213 C10_P_btm.t624 1.67819
R32428 C10_P_btm.n210 C10_P_btm.t1039 1.67819
R32429 C10_P_btm.n207 C10_P_btm.t727 1.67819
R32430 C10_P_btm.n3567 C10_P_btm.t443 1.67819
R32431 C10_P_btm.n3561 C10_P_btm.t999 1.67819
R32432 C10_P_btm.n3558 C10_P_btm.t226 1.67819
R32433 C10_P_btm.n3555 C10_P_btm.t942 1.67819
R32434 C10_P_btm.n3552 C10_P_btm.t473 1.67819
R32435 C10_P_btm.n3549 C10_P_btm.t339 1.67819
R32436 C10_P_btm.n3546 C10_P_btm.t60 1.67819
R32437 C10_P_btm.n3543 C10_P_btm.t282 1.67819
R32438 C10_P_btm.n3540 C10_P_btm.t1044 1.67819
R32439 C10_P_btm.n3537 C10_P_btm.t479 1.67819
R32440 C10_P_btm.n3530 C10_P_btm.t912 1.67819
R32441 C10_P_btm.n3527 C10_P_btm.t127 1.67819
R32442 C10_P_btm.n3524 C10_P_btm.t962 1.67819
R32443 C10_P_btm.n3521 C10_P_btm.t735 1.67819
R32444 C10_P_btm.n3518 C10_P_btm.t1028 1.67819
R32445 C10_P_btm.n3515 C10_P_btm.t795 1.67819
R32446 C10_P_btm.n3512 C10_P_btm.t551 1.67819
R32447 C10_P_btm.n3509 C10_P_btm.t895 1.67819
R32448 C10_P_btm.n3506 C10_P_btm.t616 1.67819
R32449 C10_P_btm.n3500 C10_P_btm.t237 1.67819
R32450 C10_P_btm.n260 C10_P_btm.t503 1.67819
R32451 C10_P_btm.n263 C10_P_btm.t171 1.67819
R32452 C10_P_btm.n266 C10_P_btm.t393 1.67819
R32453 C10_P_btm.n269 C10_P_btm.t637 1.67819
R32454 C10_P_btm.n272 C10_P_btm.t345 1.67819
R32455 C10_P_btm.n275 C10_P_btm.t572 1.67819
R32456 C10_P_btm.n278 C10_P_btm.t812 1.67819
R32457 C10_P_btm.n280 C10_P_btm.t1052 1.67819
R32458 C10_P_btm.n3470 C10_P_btm.t93 1.67819
R32459 C10_P_btm.n3473 C10_P_btm.t290 1.67819
R32460 C10_P_btm.n3476 C10_P_btm.t43 1.67819
R32461 C10_P_btm.n3479 C10_P_btm.t907 1.67819
R32462 C10_P_btm.n3482 C10_P_btm.t121 1.67819
R32463 C10_P_btm.n3485 C10_P_btm.t955 1.67819
R32464 C10_P_btm.n3488 C10_P_btm.t729 1.67819
R32465 C10_P_btm.n3491 C10_P_btm.t420 1.67819
R32466 C10_P_btm.n3494 C10_P_btm.t787 1.67819
R32467 C10_P_btm.n3439 C10_P_btm.t1047 1.67819
R32468 C10_P_btm.n3442 C10_P_btm.t681 1.67819
R32469 C10_P_btm.n3445 C10_P_btm.t336 1.67819
R32470 C10_P_btm.n3448 C10_P_btm.t565 1.67819
R32471 C10_P_btm.n3451 C10_P_btm.t803 1.67819
R32472 C10_P_btm.n3454 C10_P_btm.t1040 1.67819
R32473 C10_P_btm.n3457 C10_P_btm.t743 1.67819
R32474 C10_P_btm.n3460 C10_P_btm.t976 1.67819
R32475 C10_P_btm.n3463 C10_P_btm.t693 1.67819
R32476 C10_P_btm.n333 C10_P_btm.t217 1.67819
R32477 C10_P_btm.n331 C10_P_btm.t1041 1.67819
R32478 C10_P_btm.n328 C10_P_btm.t158 1.67819
R32479 C10_P_btm.n325 C10_P_btm.t989 1.67819
R32480 C10_P_btm.n322 C10_P_btm.t210 1.67819
R32481 C10_P_btm.n319 C10_P_btm.t45 1.67819
R32482 C10_P_btm.n316 C10_P_btm.t817 1.67819
R32483 C10_P_btm.n313 C10_P_btm.t91 1.67819
R32484 C10_P_btm.n3433 C10_P_btm.t870 1.67819
R32485 C10_P_btm.n3427 C10_P_btm.t487 1.67819
R32486 C10_P_btm.n3424 C10_P_btm.t765 1.67819
R32487 C10_P_btm.n3421 C10_P_btm.t424 1.67819
R32488 C10_P_btm.n3418 C10_P_btm.t658 1.67819
R32489 C10_P_btm.n3415 C10_P_btm.t889 1.67819
R32490 C10_P_btm.n3412 C10_P_btm.t605 1.67819
R32491 C10_P_btm.n3409 C10_P_btm.t836 1.67819
R32492 C10_P_btm.n3406 C10_P_btm.t344 1.67819
R32493 C10_P_btm.n3403 C10_P_btm.t788 1.67819
R32494 C10_P_btm.n3396 C10_P_btm.t387 1.67819
R32495 C10_P_btm.n3393 C10_P_btm.t683 1.67819
R32496 C10_P_btm.n3390 C10_P_btm.t451 1.67819
R32497 C10_P_btm.n3387 C10_P_btm.t222 1.67819
R32498 C10_P_btm.n3384 C10_P_btm.t993 1.67819
R32499 C10_P_btm.n3381 C10_P_btm.t270 1.67819
R32500 C10_P_btm.n3378 C10_P_btm.t104 1.67819
R32501 C10_P_btm.n3375 C10_P_btm.t378 1.67819
R32502 C10_P_btm.n3372 C10_P_btm.t110 1.67819
R32503 C10_P_btm.n3366 C10_P_btm.t77 1.67819
R32504 C10_P_btm.n366 C10_P_btm.t354 1.67819
R32505 C10_P_btm.n369 C10_P_btm.t236 1.67819
R32506 C10_P_btm.n372 C10_P_btm.t250 1.67819
R32507 C10_P_btm.n375 C10_P_btm.t484 1.67819
R32508 C10_P_btm.n378 C10_P_btm.t194 1.67819
R32509 C10_P_btm.n381 C10_P_btm.t423 1.67819
R32510 C10_P_btm.n384 C10_P_btm.t655 1.67819
R32511 C10_P_btm.n386 C10_P_btm.t371 1.67819
R32512 C10_P_btm.n3336 C10_P_btm.t758 1.67819
R32513 C10_P_btm.n3339 C10_P_btm.t34 1.67819
R32514 C10_P_btm.n3342 C10_P_btm.t816 1.67819
R32515 C10_P_btm.n3345 C10_P_btm.t582 1.67819
R32516 C10_P_btm.n3348 C10_P_btm.t866 1.67819
R32517 C10_P_btm.n3351 C10_P_btm.t641 1.67819
R32518 C10_P_btm.n3354 C10_P_btm.t398 1.67819
R32519 C10_P_btm.n3357 C10_P_btm.t742 1.67819
R32520 C10_P_btm.n3360 C10_P_btm.t458 1.67819
R32521 C10_P_btm.n3305 C10_P_btm.t874 1.67819
R32522 C10_P_btm.n3308 C10_P_btm.t103 1.67819
R32523 C10_P_btm.n3311 C10_P_btm.t819 1.67819
R32524 C10_P_btm.n3314 C10_P_btm.t974 1.67819
R32525 C10_P_btm.n3317 C10_P_btm.t212 1.67819
R32526 C10_P_btm.n3320 C10_P_btm.t753 1.67819
R32527 C10_P_btm.n3323 C10_P_btm.t164 1.67819
R32528 C10_P_btm.n3326 C10_P_btm.t386 1.67819
R32529 C10_P_btm.n3329 C10_P_btm.t234 1.67819
R32530 C10_P_btm.n468 C10_P_btm.t725 1.67819
R32531 C10_P_btm.n465 C10_P_btm.t629 1.67819
R32532 C10_P_btm.n462 C10_P_btm.t784 1.67819
R32533 C10_P_btm.n459 C10_P_btm.t541 1.67819
R32534 C10_P_btm.n456 C10_P_btm.t308 1.67819
R32535 C10_P_btm.n453 C10_P_btm.t600 1.67819
R32536 C10_P_btm.n450 C10_P_btm.t369 1.67819
R32537 C10_P_btm.n447 C10_P_btm.t138 1.67819
R32538 C10_P_btm.n444 C10_P_btm.t480 1.67819
R32539 C10_P_btm.n3299 C10_P_btm.t191 1.67819
R32540 C10_P_btm.n3293 C10_P_btm.t580 1.67819
R32541 C10_P_btm.n3290 C10_P_btm.t865 1.67819
R32542 C10_P_btm.n3287 C10_P_btm.t520 1.67819
R32543 C10_P_btm.n3284 C10_P_btm.t183 1.67819
R32544 C10_P_btm.n3281 C10_P_btm.t985 1.67819
R32545 C10_P_btm.n3278 C10_P_btm.t702 1.67819
R32546 C10_P_btm.n3275 C10_P_btm.t932 1.67819
R32547 C10_P_btm.n3272 C10_P_btm.t117 1.67819
R32548 C10_P_btm.n3269 C10_P_btm.t882 1.67819
R32549 C10_P_btm.n3266 C10_P_btm.t218 1.67819
R32550 C10_P_btm.n3263 C10_P_btm.t776 1.67819
R32551 C10_P_btm.n3260 C10_P_btm.t579 1.67819
R32552 C10_P_btm.n3257 C10_P_btm.t233 1.67819
R32553 C10_P_btm.n3254 C10_P_btm.t454 1.67819
R32554 C10_P_btm.n3251 C10_P_btm.t686 1.67819
R32555 C10_P_btm.n3248 C10_P_btm.t964 1.67819
R32556 C10_P_btm.n3245 C10_P_btm.t634 1.67819
R32557 C10_P_btm.n3242 C10_P_btm.t856 1.67819
R32558 C10_P_btm.n3239 C10_P_btm.t81 1.67819
R32559 C10_P_btm.n3236 C10_P_btm.t808 1.67819
R32560 C10_P_btm.n3233 C10_P_btm.t1035 1.67819
R32561 C10_P_btm.n3230 C10_P_btm.t747 1.67819
R32562 C10_P_btm.n3227 C10_P_btm.t979 1.67819
R32563 C10_P_btm.n504 C10_P_btm.t653 1.67819
R32564 C10_P_btm.n501 C10_P_btm.t935 1.67819
R32565 C10_P_btm.n498 C10_P_btm.t707 1.67819
R32566 C10_P_btm.n495 C10_P_btm.t41 1.67819
R32567 C10_P_btm.n492 C10_P_btm.t760 1.67819
R32568 C10_P_btm.n489 C10_P_btm.t523 1.67819
R32569 C10_P_btm.n486 C10_P_btm.t869 1.67819
R32570 C10_P_btm.n483 C10_P_btm.t584 1.67819
R32571 C10_P_btm.n480 C10_P_btm.t350 1.67819
R32572 C10_P_btm.n477 C10_P_btm.t904 1.67819
R32573 C10_P_btm.n474 C10_P_btm.t674 1.67819
R32574 C10_P_btm.n471 C10_P_btm.t1037 1.67819
R32575 C10_P_btm.n3224 C10_P_btm.t146 1.67819
R32576 C10_P_btm.n3221 C10_P_btm.t875 1.67819
R32577 C10_P_btm.n3218 C10_P_btm.t105 1.67819
R32578 C10_P_btm.n3215 C10_P_btm.t317 1.67819
R32579 C10_P_btm.n3212 C10_P_btm.t961 1.67819
R32580 C10_P_btm.n3209 C10_P_btm.t267 1.67819
R32581 C10_P_btm.n3206 C10_P_btm.t994 1.67819
R32582 C10_P_btm.n3203 C10_P_btm.t165 1.67819
R32583 C10_P_btm.n3200 C10_P_btm.t448 1.67819
R32584 C10_P_btm.n3197 C10_P_btm.t239 1.67819
R32585 C10_P_btm.n3194 C10_P_btm.t334 1.67819
R32586 C10_P_btm.n3191 C10_P_btm.t563 1.67819
R32587 C10_P_btm.n3188 C10_P_btm.t279 1.67819
R32588 C10_P_btm.n3185 C10_P_btm.t1036 1.67819
R32589 C10_P_btm.n3182 C10_P_btm.t177 1.67819
R32590 C10_P_btm.n3179 C10_P_btm.t457 1.67819
R32591 C10_P_btm.n3176 C10_P_btm.t692 1.67819
R32592 C10_P_btm.n3173 C10_P_btm.t388 1.67819
R32593 C10_P_btm.n3170 C10_P_btm.t682 1.67819
R32594 C10_P_btm.n3167 C10_P_btm.t910 1.67819
R32595 C10_P_btm.n3164 C10_P_btm.t568 1.67819
R32596 C10_P_btm.n3161 C10_P_btm.t805 1.67819
R32597 C10_P_btm.n3158 C10_P_btm.t475 1.67819
R32598 C10_P_btm.n3155 C10_P_btm.t744 1.67819
R32599 C10_P_btm.n3152 C10_P_btm.t977 1.67819
R32600 C10_P_btm.n3149 C10_P_btm.t694 1.67819
R32601 C10_P_btm.n3146 C10_P_btm.t921 1.67819
R32602 C10_P_btm.n3143 C10_P_btm.t96 1.67819
R32603 C10_P_btm.n3140 C10_P_btm.t429 1.67819
R32604 C10_P_btm.n3137 C10_P_btm.t50 1.67819
R32605 C10_P_btm.n3134 C10_P_btm.t262 1.67819
R32606 C10_P_btm.n3131 C10_P_btm.t991 1.67819
R32607 C10_P_btm.n3128 C10_P_btm.t209 1.67819
R32608 C10_P_btm.n3125 C10_P_btm.t934 1.67819
R32609 C10_P_btm.n3122 C10_P_btm.t227 1.67819
R32610 C10_P_btm.n3119 C10_P_btm.t384 1.67819
R32611 C10_P_btm.n3116 C10_P_btm.t474 1.67819
R32612 C10_P_btm.n3113 C10_P_btm.t278 1.67819
R32613 C10_P_btm.n3110 C10_P_btm.t559 1.67819
R32614 C10_P_btm.n3103 C10_P_btm.t465 1.67819
R32615 C10_P_btm.n3100 C10_P_btm.t185 1.67819
R32616 C10_P_btm.n3097 C10_P_btm.t1015 1.67819
R32617 C10_P_btm.n3094 C10_P_btm.t284 1.67819
R32618 C10_P_btm.n3091 C10_P_btm.t48 1.67819
R32619 C10_P_btm.n3088 C10_P_btm.t845 1.67819
R32620 C10_P_btm.n3085 C10_P_btm.t512 1.67819
R32621 C10_P_btm.n3082 C10_P_btm.t899 1.67819
R32622 C10_P_btm.n3079 C10_P_btm.t172 1.67819
R32623 C10_P_btm.n3076 C10_P_btm.t1002 1.67819
R32624 C10_P_btm.n3021 C10_P_btm.t78 1.67819
R32625 C10_P_btm.n3018 C10_P_btm.t806 1.67819
R32626 C10_P_btm.n3015 C10_P_btm.t514 1.67819
R32627 C10_P_btm.n3012 C10_P_btm.t745 1.67819
R32628 C10_P_btm.n3009 C10_P_btm.t978 1.67819
R32629 C10_P_btm.n3006 C10_P_btm.t195 1.67819
R32630 C10_P_btm.n3003 C10_P_btm.t922 1.67819
R32631 C10_P_btm.n3000 C10_P_btm.t99 1.67819
R32632 C10_P_btm.n2997 C10_P_btm.t372 1.67819
R32633 C10_P_btm.n2991 C10_P_btm.t715 1.67819
R32634 C10_P_btm.n2989 C10_P_btm.t428 1.67819
R32635 C10_P_btm.n2986 C10_P_btm.t200 1.67819
R32636 C10_P_btm.n2983 C10_P_btm.t532 1.67819
R32637 C10_P_btm.n2980 C10_P_btm.t252 1.67819
R32638 C10_P_btm.n2977 C10_P_btm.t1033 1.67819
R32639 C10_P_btm.n2974 C10_P_btm.t357 1.67819
R32640 C10_P_btm.n2971 C10_P_btm.t83 1.67819
R32641 C10_P_btm.n2968 C10_P_btm.t409 1.67819
R32642 C10_P_btm.n2962 C10_P_btm.t313 1.67819
R32643 C10_P_btm.n2904 C10_P_btm.t56 1.67819
R32644 C10_P_btm.n2907 C10_P_btm.t263 1.67819
R32645 C10_P_btm.n2910 C10_P_btm.t992 1.67819
R32646 C10_P_btm.n2913 C10_P_btm.t161 1.67819
R32647 C10_P_btm.n2916 C10_P_btm.t445 1.67819
R32648 C10_P_btm.n2919 C10_P_btm.t231 1.67819
R32649 C10_P_btm.n2922 C10_P_btm.t331 1.67819
R32650 C10_P_btm.n2925 C10_P_btm.t626 1.67819
R32651 C10_P_btm.n2932 C10_P_btm.t374 1.67819
R32652 C10_P_btm.n2935 C10_P_btm.t467 1.67819
R32653 C10_P_btm.n2938 C10_P_btm.t518 1.67819
R32654 C10_P_btm.n2941 C10_P_btm.t577 1.67819
R32655 C10_P_btm.n2944 C10_P_btm.t287 1.67819
R32656 C10_P_btm.n2947 C10_P_btm.t70 1.67819
R32657 C10_P_btm.n2950 C10_P_btm.t397 1.67819
R32658 C10_P_btm.n2953 C10_P_btm.t967 1.67819
R32659 C10_P_btm.n2956 C10_P_btm.t456 1.67819
R32660 C10_P_btm.n2866 C10_P_btm.t546 1.67819
R32661 C10_P_btm.n2869 C10_P_btm.t215 1.67819
R32662 C10_P_btm.n2872 C10_P_btm.t929 1.67819
R32663 C10_P_btm.n2875 C10_P_btm.t167 1.67819
R32664 C10_P_btm.n2878 C10_P_btm.t1045 1.67819
R32665 C10_P_btm.n2881 C10_P_btm.t680 1.67819
R32666 C10_P_btm.n2884 C10_P_btm.t335 1.67819
R32667 C10_P_btm.n2887 C10_P_btm.t564 1.67819
R32668 C10_P_btm.n2890 C10_P_btm.t853 1.67819
R32669 C10_P_btm.n2144 C10_P_btm.t944 1.67819
R32670 C10_P_btm.n2142 C10_P_btm.t666 1.67819
R32671 C10_P_btm.n2139 C10_P_btm.t433 1.67819
R32672 C10_P_btm.n2136 C10_P_btm.t773 1.67819
R32673 C10_P_btm.n2133 C10_P_btm.t499 1.67819
R32674 C10_P_btm.n2130 C10_P_btm.t255 1.67819
R32675 C10_P_btm.n2127 C10_P_btm.t593 1.67819
R32676 C10_P_btm.n2124 C10_P_btm.t300 1.67819
R32677 C10_P_btm.n2860 C10_P_btm.t646 1.67819
R32678 C10_P_btm.n2854 C10_P_btm.t528 1.67819
R32679 C10_P_btm.n2851 C10_P_btm.t197 1.67819
R32680 C10_P_btm.n2848 C10_P_btm.t485 1.67819
R32681 C10_P_btm.n2845 C10_P_btm.t142 1.67819
R32682 C10_P_btm.n2842 C10_P_btm.t373 1.67819
R32683 C10_P_btm.n2839 C10_P_btm.t657 1.67819
R32684 C10_P_btm.n2836 C10_P_btm.t312 1.67819
R32685 C10_P_btm.n2833 C10_P_btm.t544 1.67819
R32686 C10_P_btm.n2830 C10_P_btm.t835 1.67819
R32687 C10_P_btm.n2823 C10_P_btm.t928 1.67819
R32688 C10_P_btm.n2820 C10_P_btm.t645 1.67819
R32689 C10_P_btm.n2817 C10_P_btm.t408 1.67819
R32690 C10_P_btm.n2814 C10_P_btm.t752 1.67819
R32691 C10_P_btm.n2811 C10_P_btm.t468 1.67819
R32692 C10_P_btm.n2808 C10_P_btm.t497 1.67819
R32693 C10_P_btm.n2805 C10_P_btm.t573 1.67819
R32694 C10_P_btm.n2802 C10_P_btm.t285 1.67819
R32695 C10_P_btm.n2799 C10_P_btm.t638 1.67819
R32696 C10_P_btm.n2793 C10_P_btm.t272 1.67819
R32697 C10_P_btm.n2177 C10_P_btm.t998 1.67819
R32698 C10_P_btm.n2180 C10_P_btm.t225 1.67819
R32699 C10_P_btm.n2183 C10_P_btm.t940 1.67819
R32700 C10_P_btm.n2186 C10_P_btm.t246 1.67819
R32701 C10_P_btm.n2189 C10_P_btm.t1051 1.67819
R32702 C10_P_btm.n2192 C10_P_btm.t58 1.67819
R32703 C10_P_btm.n2195 C10_P_btm.t281 1.67819
R32704 C10_P_btm.n2197 C10_P_btm.t567 1.67819
R32705 C10_P_btm.n2763 C10_P_btm.t670 1.67819
R32706 C10_P_btm.n2766 C10_P_btm.t380 1.67819
R32707 C10_P_btm.n2769 C10_P_btm.t152 1.67819
R32708 C10_P_btm.n2772 C10_P_btm.t510 1.67819
R32709 C10_P_btm.n2775 C10_P_btm.t204 1.67819
R32710 C10_P_btm.n2778 C10_P_btm.t53 1.67819
R32711 C10_P_btm.n2781 C10_P_btm.t302 1.67819
R32712 C10_P_btm.n2784 C10_P_btm.t36 1.67819
R32713 C10_P_btm.n2787 C10_P_btm.t363 1.67819
R32714 C10_P_btm.n2732 C10_P_btm.t460 1.67819
R32715 C10_P_btm.n2735 C10_P_btm.t125 1.67819
R32716 C10_P_btm.n2738 C10_P_btm.t399 1.67819
R32717 C10_P_btm.n2741 C10_P_btm.t74 1.67819
R32718 C10_P_btm.n2744 C10_P_btm.t293 1.67819
R32719 C10_P_btm.n2747 C10_P_btm.t583 1.67819
R32720 C10_P_btm.n2750 C10_P_btm.t1011 1.67819
R32721 C10_P_btm.n2753 C10_P_btm.t478 1.67819
R32722 C10_P_btm.n2756 C10_P_btm.t759 1.67819
R32723 C10_P_btm.n2250 C10_P_btm.t395 1.67819
R32724 C10_P_btm.n2248 C10_P_btm.t770 1.67819
R32725 C10_P_btm.n2245 C10_P_btm.t950 1.67819
R32726 C10_P_btm.n2242 C10_P_btm.t238 1.67819
R32727 C10_P_btm.n2239 C10_P_btm.t1006 1.67819
R32728 C10_P_btm.n2236 C10_P_btm.t780 1.67819
R32729 C10_P_btm.n2233 C10_P_btm.t235 1.67819
R32730 C10_P_btm.n2230 C10_P_btm.t833 1.67819
R32731 C10_P_btm.n2726 C10_P_btm.t214 1.67819
R32732 C10_P_btm.n2720 C10_P_btm.t198 1.67819
R32733 C10_P_btm.n2717 C10_P_btm.t925 1.67819
R32734 C10_P_btm.n2714 C10_P_btm.t143 1.67819
R32735 C10_P_btm.n2711 C10_P_btm.t873 1.67819
R32736 C10_P_btm.n2708 C10_P_btm.t92 1.67819
R32737 C10_P_btm.n2705 C10_P_btm.t314 1.67819
R32738 C10_P_btm.n2702 C10_P_btm.t220 1.67819
R32739 C10_P_btm.n2699 C10_P_btm.t213 1.67819
R32740 C10_P_btm.n2696 C10_P_btm.t757 1.67819
R32741 C10_P_btm.n2689 C10_P_btm.t134 1.67819
R32742 C10_P_btm.n2686 C10_P_btm.t917 1.67819
R32743 C10_P_btm.n2683 C10_P_btm.t689 1.67819
R32744 C10_P_btm.n2680 C10_P_btm.t1021 1.67819
R32745 C10_P_btm.n2677 C10_P_btm.t741 1.67819
R32746 C10_P_btm.n2674 C10_P_btm.t505 1.67819
R32747 C10_P_btm.n2671 C10_P_btm.t850 1.67819
R32748 C10_P_btm.n2668 C10_P_btm.t560 1.67819
R32749 C10_P_btm.n2665 C10_P_btm.t906 1.67819
R32750 C10_P_btm.n2659 C10_P_btm.t1000 1.67819
R32751 C10_P_btm.n2283 C10_P_btm.t663 1.67819
R32752 C10_P_btm.n2286 C10_P_btm.t941 1.67819
R32753 C10_P_btm.n2289 C10_P_btm.t609 1.67819
R32754 C10_P_btm.n2292 C10_P_btm.t841 1.67819
R32755 C10_P_btm.n2295 C10_P_btm.t59 1.67819
R32756 C10_P_btm.n2298 C10_P_btm.t791 1.67819
R32757 C10_P_btm.n2301 C10_P_btm.t1027 1.67819
R32758 C10_P_btm.n2303 C10_P_btm.t482 1.67819
R32759 C10_P_btm.n2629 C10_P_btm.t323 1.67819
R32760 C10_P_btm.n2632 C10_P_btm.t115 1.67819
R32761 C10_P_btm.n2635 C10_P_btm.t880 1.67819
R32762 C10_P_btm.n2638 C10_P_btm.t154 1.67819
R32763 C10_P_btm.n2641 C10_P_btm.t931 1.67819
R32764 C10_P_btm.n2644 C10_P_btm.t701 1.67819
R32765 C10_P_btm.n2647 C10_P_btm.t109 1.67819
R32766 C10_P_btm.n2650 C10_P_btm.t756 1.67819
R32767 C10_P_btm.n2653 C10_P_btm.t39 1.67819
R32768 C10_P_btm.n2598 C10_P_btm.t736 1.67819
R32769 C10_P_btm.n2601 C10_P_btm.t391 1.67819
R32770 C10_P_btm.n2604 C10_P_btm.t685 1.67819
R32771 C10_P_btm.n2607 C10_P_btm.t341 1.67819
R32772 C10_P_btm.n2610 C10_P_btm.t570 1.67819
R32773 C10_P_btm.n2613 C10_P_btm.t855 1.67819
R32774 C10_P_btm.n2616 C10_P_btm.t1046 1.67819
R32775 C10_P_btm.n2619 C10_P_btm.t748 1.67819
R32776 C10_P_btm.n2622 C10_P_btm.t221 1.67819
R32777 C10_P_btm.n2356 C10_P_btm.t67 1.67819
R32778 C10_P_btm.n2354 C10_P_btm.t847 1.67819
R32779 C10_P_btm.n2351 C10_P_btm.t620 1.67819
R32780 C10_P_btm.n2348 C10_P_btm.t951 1.67819
R32781 C10_P_btm.n2345 C10_P_btm.t673 1.67819
R32782 C10_P_btm.n2342 C10_P_btm.t439 1.67819
R32783 C10_P_btm.n2339 C10_P_btm.t781 1.67819
R32784 C10_P_btm.n2336 C10_P_btm.t522 1.67819
R32785 C10_P_btm.n2592 C10_P_btm.t412 1.67819
R32786 C10_P_btm.n2586 C10_P_btm.t466 1.67819
R32787 C10_P_btm.n2583 C10_P_btm.t131 1.67819
R32788 C10_P_btm.n2580 C10_P_btm.t407 1.67819
R32789 C10_P_btm.n2577 C10_P_btm.t82 1.67819
R32790 C10_P_btm.n2574 C10_P_btm.t298 1.67819
R32791 C10_P_btm.n2571 C10_P_btm.t588 1.67819
R32792 C10_P_btm.n2568 C10_P_btm.t251 1.67819
R32793 C10_P_btm.n2565 C10_P_btm.t496 1.67819
R32794 C10_P_btm.n2562 C10_P_btm.t767 1.67819
R32795 C10_P_btm.n2555 C10_P_btm.t862 1.67819
R32796 C10_P_btm.n2552 C10_P_btm.t575 1.67819
R32797 C10_P_btm.n2549 C10_P_btm.t348 1.67819
R32798 C10_P_btm.n2546 C10_P_btm.t690 1.67819
R32799 C10_P_btm.n2543 C10_P_btm.t396 1.67819
R32800 C10_P_btm.n2540 C10_P_btm.t176 1.67819
R32801 C10_P_btm.n2537 C10_P_btm.t506 1.67819
R32802 C10_P_btm.n2534 C10_P_btm.t244 1.67819
R32803 C10_P_btm.n2531 C10_P_btm.t561 1.67819
R32804 C10_P_btm.n2525 C10_P_btm.t665 1.67819
R32805 C10_P_btm.n2389 C10_P_btm.t318 1.67819
R32806 C10_P_btm.n2392 C10_P_btm.t610 1.67819
R32807 C10_P_btm.n2395 C10_P_btm.t268 1.67819
R32808 C10_P_btm.n2398 C10_P_btm.t867 1.67819
R32809 C10_P_btm.n2401 C10_P_btm.t792 1.67819
R32810 C10_P_btm.n2404 C10_P_btm.t449 1.67819
R32811 C10_P_btm.n2407 C10_P_btm.t679 1.67819
R32812 C10_P_btm.n2409 C10_P_btm.t958 1.67819
R32813 C10_P_btm.n2495 C10_P_btm.t597 1.67819
R32814 C10_P_btm.n2498 C10_P_btm.t307 1.67819
R32815 C10_P_btm.n2501 C10_P_btm.t88 1.67819
R32816 C10_P_btm.n2504 C10_P_btm.t416 1.67819
R32817 C10_P_btm.n2507 C10_P_btm.t137 1.67819
R32818 C10_P_btm.n2510 C10_P_btm.t973 1.67819
R32819 C10_P_btm.n2513 C10_P_btm.t966 1.67819
R32820 C10_P_btm.n2516 C10_P_btm.t1025 1.67819
R32821 C10_P_btm.n2519 C10_P_btm.t292 1.67819
R32822 C10_P_btm.n2464 C10_P_btm.t392 1.67819
R32823 C10_P_btm.n2467 C10_P_btm.t63 1.67819
R32824 C10_P_btm.n2470 C10_P_btm.t342 1.67819
R32825 C10_P_btm.n2473 C10_P_btm.t242 1.67819
R32826 C10_P_btm.n2476 C10_P_btm.t489 1.67819
R32827 C10_P_btm.n2479 C10_P_btm.t1048 1.67819
R32828 C10_P_btm.n2482 C10_P_btm.t182 1.67819
R32829 C10_P_btm.n2485 C10_P_btm.t403 1.67819
R32830 C10_P_btm.n2488 C10_P_btm.t696 1.67819
R32831 C10_P_btm.n2432 C10_P_btm.t332 1.67819
R32832 C10_P_btm.n2435 C10_P_btm.t491 1.67819
R32833 C10_P_btm.n2438 C10_P_btm.t887 1.67819
R32834 C10_P_btm.n2441 C10_P_btm.t162 1.67819
R32835 C10_P_btm.n2444 C10_P_btm.t936 1.67819
R32836 C10_P_btm.n2447 C10_P_btm.t710 1.67819
R32837 C10_P_btm.n2450 C10_P_btm.t1053 1.67819
R32838 C10_P_btm.n2453 C10_P_btm.t763 1.67819
R32839 C10_P_btm.n2458 C10_P_btm.t87 1.67819
R32840 C10_P_btm.n3073 C10_P_btm.t777 1.67819
R32841 C10_P_btm.n3070 C10_P_btm.t578 1.67819
R32842 C10_P_btm.n3067 C10_P_btm.t829 1.67819
R32843 C10_P_btm.n3064 C10_P_btm.t595 1.67819
R32844 C10_P_btm.n3061 C10_P_btm.t883 1.67819
R32845 C10_P_btm.n3058 C10_P_btm.t649 1.67819
R32846 C10_P_btm.n3055 C10_P_btm.t986 1.67819
R32847 C10_P_btm.n3052 C10_P_btm.t704 1.67819
R32848 C10_P_btm.n3049 C10_P_btm.t470 1.67819
R32849 C10_P_btm.n3046 C10_P_btm.t815 1.67819
R32850 C10_P_btm.n3043 C10_P_btm.t581 1.67819
R32851 C10_P_btm.n3040 C10_P_btm.t288 1.67819
R32852 C10_P_btm.n2052 C10_P_btm.t203 1.67819
R32853 C10_P_btm.n2049 C10_P_btm.t982 1.67819
R32854 C10_P_btm.n2046 C10_P_btm.t755 1.67819
R32855 C10_P_btm.n2043 C10_P_btm.t35 1.67819
R32856 C10_P_btm.n2040 C10_P_btm.t813 1.67819
R32857 C10_P_btm.n2037 C10_P_btm.t574 1.67819
R32858 C10_P_btm.n2034 C10_P_btm.t916 1.67819
R32859 C10_P_btm.n2031 C10_P_btm.t639 1.67819
R32860 C10_P_btm.n2028 C10_P_btm.t970 1.67819
R32861 C10_P_btm.n2025 C10_P_btm.t739 1.67819
R32862 C10_P_btm.n2022 C10_P_btm.t504 1.67819
R32863 C10_P_btm.n2019 C10_P_btm.t799 1.67819
R32864 C10_P_btm.n2016 C10_P_btm.t557 1.67819
R32865 C10_P_btm.n2013 C10_P_btm.t327 1.67819
R32866 C10_P_btm.n2010 C10_P_btm.t623 1.67819
R32867 C10_P_btm.n2007 C10_P_btm.t383 1.67819
R32868 C10_P_btm.n2004 C10_P_btm.t726 1.67819
R32869 C10_P_btm.n2001 C10_P_btm.t442 1.67819
R32870 C10_P_btm.n1998 C10_P_btm.t208 1.67819
R32871 C10_P_btm.n1995 C10_P_btm.t543 1.67819
R32872 C10_P_btm.n1992 C10_P_btm.t309 1.67819
R32873 C10_P_btm.n1989 C10_P_btm.t47 1.67819
R32874 C10_P_btm.n1986 C10_P_btm.t325 1.67819
R32875 C10_P_btm.n1983 C10_P_btm.t114 1.67819
R32876 C10_P_btm.n1980 C10_P_btm.t881 1.67819
R32877 C10_P_btm.n1977 C10_P_btm.t156 1.67819
R32878 C10_P_btm.n1974 C10_P_btm.t984 1.67819
R32879 C10_P_btm.n1971 C10_P_btm.t206 1.67819
R32880 C10_P_btm.n1968 C10_P_btm.t476 1.67819
R32881 C10_P_btm.n1965 C10_P_btm.t814 1.67819
R32882 C10_P_btm.n1962 C10_P_btm.t85 1.67819
R32883 C10_P_btm.n1959 C10_P_btm.t863 1.67819
R32884 C10_P_btm.n1956 C10_P_btm.t640 1.67819
R32885 C10_P_btm.n1953 C10_P_btm.t972 1.67819
R32886 C10_P_btm.n1950 C10_P_btm.t691 1.67819
R32887 C10_P_btm.n1947 C10_P_btm.t1024 1.67819
R32888 C10_P_btm.n1944 C10_P_btm.t801 1.67819
R32889 C10_P_btm.n1941 C10_P_btm.t508 1.67819
R32890 C10_P_btm.n1938 C10_P_btm.t852 1.67819
R32891 C10_P_btm.n1935 C10_P_btm.t627 1.67819
R32892 C10_P_btm.n1932 C10_P_btm.t1043 1.67819
R32893 C10_P_btm.n1929 C10_P_btm.t678 1.67819
R32894 C10_P_btm.n1926 C10_P_btm.t447 1.67819
R32895 C10_P_btm.n1923 C10_P_btm.t790 1.67819
R32896 C10_P_btm.n1920 C10_P_btm.t768 1.67819
R32897 C10_P_btm.n1917 C10_P_btm.t265 1.67819
R32898 C10_P_btm.n1914 C10_P_btm.t608 1.67819
R32899 C10_P_btm.n1911 C10_P_btm.t315 1.67819
R32900 C10_P_btm.n1908 C10_P_btm.t102 1.67819
R32901 C10_P_btm.n1905 C10_P_btm.t733 1.67819
R32902 C10_P_btm.n1902 C10_P_btm.t965 1.67819
R32903 C10_P_btm.n1899 C10_P_btm.t216 1.67819
R32904 C10_P_btm.n1896 C10_P_btm.t548 1.67819
R32905 C10_P_btm.n1893 C10_P_btm.t320 1.67819
R32906 C10_P_btm.n1890 C10_P_btm.t613 1.67819
R32907 C10_P_btm.n1887 C10_P_btm.t377 1.67819
R32908 C10_P_btm.n1884 C10_P_btm.t148 1.67819
R32909 C10_P_btm.n1881 C10_P_btm.t431 1.67819
R32910 C10_P_btm.n1878 C10_P_btm.t202 1.67819
R32911 C10_P_btm.n1875 C10_P_btm.t38 1.67819
R32912 C10_P_btm.n1872 C10_P_btm.t299 1.67819
R32913 C10_P_btm.n1869 C10_P_btm.t32 1.67819
R32914 C10_P_btm.n1863 C10_P_btm.t405 1.67819
R32915 C10_P_btm.n735 C10_P_btm.t697 1.67819
R32916 C10_P_btm.n738 C10_P_btm.t355 1.67819
R32917 C10_P_btm.n741 C10_P_btm.t587 1.67819
R32918 C10_P_btm.n744 C10_P_btm.t821 1.67819
R32919 C10_P_btm.n747 C10_P_btm.t527 1.67819
R32920 C10_P_btm.n750 C10_P_btm.t764 1.67819
R32921 C10_P_btm.n753 C10_P_btm.t996 1.67819
R32922 C10_P_btm.n756 C10_P_btm.t711 1.67819
R32923 C10_P_btm.n759 C10_P_btm.t937 1.67819
R32924 C10_P_btm.n762 C10_P_btm.t604 1.67819
R32925 C10_P_btm.n765 C10_P_btm.t888 1.67819
R32926 C10_P_btm.n768 C10_P_btm.t513 1.67819
R32927 C10_P_btm.n771 C10_P_btm.t186 1.67819
R32928 C10_P_btm.n774 C10_P_btm.t410 1.67819
R32929 C10_P_btm.n777 C10_P_btm.t700 1.67819
R32930 C10_P_btm.n780 C10_P_btm.t358 1.67819
R32931 C10_P_btm.n783 C10_P_btm.t590 1.67819
R32932 C10_P_btm.n786 C10_P_btm.t879 1.67819
R32933 C10_P_btm.n789 C10_P_btm.t533 1.67819
R32934 C10_P_btm.n792 C10_P_btm.t772 1.67819
R32935 C10_P_btm.n795 C10_P_btm.t495 1.67819
R32936 C10_P_btm.n798 C10_P_btm.t716 1.67819
R32937 C10_P_btm.n801 C10_P_btm.t943 1.67819
R32938 C10_P_btm.n804 C10_P_btm.t611 1.67819
R32939 C10_P_btm.n807 C10_P_btm.t893 1.67819
R32940 C10_P_btm.n810 C10_P_btm.t62 1.67819
R32941 C10_P_btm.n813 C10_P_btm.t793 1.67819
R32942 C10_P_btm.n816 C10_P_btm.t490 1.67819
R32943 C10_P_btm.n819 C10_P_btm.t731 1.67819
R32944 C10_P_btm.n822 C10_P_btm.t959 1.67819
R32945 C10_P_btm.n825 C10_P_btm.t181 1.67819
R32946 C10_P_btm.n828 C10_P_btm.t909 1.67819
R32947 C10_P_btm.n831 C10_P_btm.t75 1.67819
R32948 C10_P_btm.n834 C10_P_btm.t294 1.67819
R32949 C10_P_btm.n837 C10_P_btm.t116 1.67819
R32950 C10_P_btm.n840 C10_P_btm.t248 1.67819
R32951 C10_P_btm.n843 C10_P_btm.t975 1.67819
R32952 C10_P_btm.n846 C10_P_btm.t192 1.67819
R32953 C10_P_btm.n849 C10_P_btm.t421 1.67819
R32954 C10_P_btm.n852 C10_P_btm.t126 1.67819
R32955 C10_P_btm.n855 C10_P_btm.t406 1.67819
R32956 C10_P_btm.n858 C10_P_btm.t644 1.67819
R32957 C10_P_btm.n861 C10_P_btm.t296 1.67819
R32958 C10_P_btm.n864 C10_P_btm.t529 1.67819
R32959 C10_P_btm.n867 C10_P_btm.t823 1.67819
R32960 C10_P_btm.n870 C10_P_btm.t488 1.67819
R32961 C10_P_btm.n873 C10_P_btm.t713 1.67819
R32962 C10_P_btm.n876 C10_P_btm.t425 1.67819
R32963 C10_P_btm.n879 C10_P_btm.t660 1.67819
R32964 C10_P_btm.n882 C10_P_btm.t890 1.67819
R32965 C10_P_btm.n885 C10_P_btm.t607 1.67819
R32966 C10_P_btm.n888 C10_P_btm.t838 1.67819
R32967 C10_P_btm.n891 C10_P_btm.t147 1.67819
R32968 C10_P_btm.n894 C10_P_btm.t730 1.67819
R32969 C10_P_btm.n897 C10_P_btm.t1018 1.67819
R32970 C10_P_btm.n900 C10_P_btm.t677 1.67819
R32971 C10_P_btm.n903 C10_P_btm.t908 1.67819
R32972 C10_P_btm.n906 C10_P_btm.t123 1.67819
R32973 C10_P_btm.n909 C10_P_btm.t851 1.67819
R32974 C10_P_btm.n912 C10_P_btm.t101 1.67819
R32975 C10_P_btm.n914 C10_P_btm.t291 1.67819
R32976 C10_P_btm.n1674 C10_P_btm.t1003 1.67819
R32977 C10_P_btm.n1677 C10_P_btm.t721 1.67819
R32978 C10_P_btm.n1680 C10_P_btm.t517 1.67819
R32979 C10_P_btm.n1683 C10_P_btm.t830 1.67819
R32980 C10_P_btm.n1686 C10_P_btm.t538 1.67819
R32981 C10_P_btm.n1689 C10_P_btm.t305 1.67819
R32982 C10_P_btm.n1692 C10_P_btm.t651 1.67819
R32983 C10_P_btm.n1695 C10_P_btm.t366 1.67819
R32984 C10_P_btm.n1698 C10_P_btm.t705 1.67819
R32985 C10_P_btm.n1701 C10_P_btm.t477 1.67819
R32986 C10_P_btm.n1704 C10_P_btm.t769 1.67819
R32987 C10_P_btm.n1707 C10_P_btm.t521 1.67819
R32988 C10_P_btm.n1710 C10_P_btm.t289 1.67819
R32989 C10_P_btm.n1713 C10_P_btm.t71 1.67819
R32990 C10_P_btm.n1716 C10_P_btm.t349 1.67819
R32991 C10_P_btm.n1719 C10_P_btm.t120 1.67819
R32992 C10_P_btm.n1722 C10_P_btm.t459 1.67819
R32993 C10_P_btm.n1725 C10_P_btm.t178 1.67819
R32994 C10_P_btm.n1728 C10_P_btm.t1009 1.67819
R32995 C10_P_btm.n1731 C10_P_btm.t280 1.67819
R32996 C10_P_btm.n1734 C10_P_btm.t771 1.67819
R32997 C10_P_btm.n1737 C10_P_btm.t834 1.67819
R32998 C10_P_btm.n1740 C10_P_btm.t69 1.67819
R32999 C10_P_btm.n1743 C10_P_btm.t903 1.67819
R33000 C10_P_btm.n1746 C10_P_btm.t622 1.67819
R33001 C10_P_btm.n1749 C10_P_btm.t954 1.67819
R33002 C10_P_btm.n1752 C10_P_btm.t724 1.67819
R33003 C10_P_btm.n1755 C10_P_btm.t1007 1.67819
R33004 C10_P_btm.n1758 C10_P_btm.t783 1.67819
R33005 C10_P_btm.n1761 C10_P_btm.t540 1.67819
R33006 C10_P_btm.n1764 C10_P_btm.t886 1.67819
R33007 C10_P_btm.n1767 C10_P_btm.t599 1.67819
R33008 C10_P_btm.n1770 C10_P_btm.t368 1.67819
R33009 C10_P_btm.n1773 C10_P_btm.t709 1.67819
R33010 C10_P_btm.n1776 C10_P_btm.t419 1.67819
R33011 C10_P_btm.n1779 C10_P_btm.t762 1.67819
R33012 C10_P_btm.n1782 C10_P_btm.t525 1.67819
R33013 C10_P_btm.n1785 C10_P_btm.t247 1.67819
R33014 C10_P_btm.n1788 C10_P_btm.t586 1.67819
R33015 C10_P_btm.n1791 C10_P_btm.t351 1.67819
R33016 C10_P_btm.n1794 C10_P_btm.t124 1.67819
R33017 C10_P_btm.n1797 C10_P_btm.t401 1.67819
R33018 C10_P_btm.n1800 C10_P_btm.t180 1.67819
R33019 C10_P_btm.n1803 C10_P_btm.t515 1.67819
R33020 C10_P_btm.n1806 C10_P_btm.t486 1.67819
R33021 C10_P_btm.n1809 C10_P_btm.t1031 1.67819
R33022 C10_P_btm.n1812 C10_P_btm.t338 1.67819
R33023 C10_P_btm.n1815 C10_P_btm.t61 1.67819
R33024 C10_P_btm.n1818 C10_P_btm.t892 1.67819
R33025 C10_P_btm.n1821 C10_P_btm.t554 1.67819
R33026 C10_P_btm.n1824 C10_P_btm.t326 1.67819
R33027 C10_P_btm.n1827 C10_P_btm.t119 1.67819
R33028 C10_P_btm.n1830 C10_P_btm.t382 1.67819
R33029 C10_P_btm.n1833 C10_P_btm.t157 1.67819
R33030 C10_P_btm.n1836 C10_P_btm.t440 1.67819
R33031 C10_P_btm.n1839 C10_P_btm.t207 1.67819
R33032 C10_P_btm.n1842 C10_P_btm.t1034 1.67819
R33033 C10_P_btm.n1845 C10_P_btm.t258 1.67819
R33034 C10_P_btm.n1848 C10_P_btm.t42 1.67819
R33035 C10_P_btm.n1851 C10_P_btm.t864 1.67819
R33036 C10_P_btm.n1854 C10_P_btm.t136 1.67819
R33037 C10_P_btm.n1857 C10_P_btm.t918 1.67819
R33038 C10_P_btm.n1484 C10_P_btm.t511 1.67819
R33039 C10_P_btm.n1487 C10_P_btm.t519 1.67819
R33040 C10_P_btm.n1490 C10_P_btm.t188 1.67819
R33041 C10_P_btm.n1493 C10_P_btm.t414 1.67819
R33042 C10_P_btm.n1496 C10_P_btm.t647 1.67819
R33043 C10_P_btm.n1499 C10_P_btm.t361 1.67819
R33044 C10_P_btm.n1502 C10_P_btm.t594 1.67819
R33045 C10_P_btm.n1505 C10_P_btm.t827 1.67819
R33046 C10_P_btm.n1508 C10_P_btm.t535 1.67819
R33047 C10_P_btm.n1511 C10_P_btm.t774 1.67819
R33048 C10_P_btm.n1514 C10_P_btm.t434 1.67819
R33049 C10_P_btm.n1517 C10_P_btm.t718 1.67819
R33050 C10_P_btm.n1520 C10_P_btm.t945 1.67819
R33051 C10_P_btm.n1523 C10_P_btm.t983 1.67819
R33052 C10_P_btm.n1526 C10_P_btm.t155 1.67819
R33053 C10_P_btm.n1529 C10_P_btm.t437 1.67819
R33054 C10_P_btm.n1532 C10_P_btm.t113 1.67819
R33055 C10_P_btm.n1535 C10_P_btm.t324 1.67819
R33056 C10_P_btm.n1538 C10_P_btm.t618 1.67819
R33057 C10_P_btm.n1541 C10_P_btm.t275 1.67819
R33058 C10_P_btm.n1544 C10_P_btm.t502 1.67819
R33059 C10_P_btm.n1547 C10_P_btm.t232 1.67819
R33060 C10_P_btm.n1550 C10_P_btm.t455 1.67819
R33061 C10_P_btm.n1553 C10_P_btm.t688 1.67819
R33062 C10_P_btm.n1556 C10_P_btm.t343 1.67819
R33063 C10_P_btm.n1559 C10_P_btm.t635 1.67819
R33064 C10_P_btm.n1562 C10_P_btm.t858 1.67819
R33065 C10_P_btm.n1565 C10_P_btm.t1050 1.67819
R33066 C10_P_btm.n1568 C10_P_btm.t809 1.67819
R33067 C10_P_btm.n1571 C10_P_btm.t463 1.67819
R33068 C10_P_btm.n1574 C10_P_btm.t698 1.67819
R33069 C10_P_btm.n1577 C10_P_btm.t980 1.67819
R33070 C10_P_btm.n1580 C10_P_btm.t643 1.67819
R33071 C10_P_btm.n1583 C10_P_btm.t876 1.67819
R33072 C10_P_btm.n1586 C10_P_btm.t97 1.67819
R33073 C10_P_btm.n1589 C10_P_btm.t820 1.67819
R33074 C10_P_btm.n1592 C10_P_btm.t898 1.67819
R33075 C10_P_btm.n1595 C10_P_btm.t712 1.67819
R33076 C10_P_btm.n1598 C10_P_btm.t995 1.67819
R33077 C10_P_btm.n1601 C10_P_btm.t166 1.67819
R33078 C10_P_btm.n1604 C10_P_btm.t927 1.67819
R33079 C10_P_btm.n1607 C10_P_btm.t150 1.67819
R33080 C10_P_btm.n1610 C10_P_btm.t379 1.67819
R33081 C10_P_btm.n1613 C10_P_btm.t112 1.67819
R33082 C10_P_btm.n1616 C10_P_btm.t274 1.67819
R33083 C10_P_btm.n1619 C10_P_btm.t550 1.67819
R33084 C10_P_btm.n1622 C10_P_btm.t229 1.67819
R33085 C10_P_btm.n1625 C10_P_btm.t453 1.67819
R33086 C10_P_btm.n1628 C10_P_btm.t168 1.67819
R33087 C10_P_btm.n1631 C10_P_btm.t389 1.67819
R33088 C10_P_btm.n1634 C10_P_btm.t633 1.67819
R33089 C10_P_btm.n1637 C10_P_btm.t337 1.67819
R33090 C10_P_btm.n1640 C10_P_btm.t569 1.67819
R33091 C10_P_btm.n1643 C10_P_btm.t807 1.67819
R33092 C10_P_btm.n1646 C10_P_btm.t462 1.67819
R33093 C10_P_btm.n1649 C10_P_btm.t746 1.67819
R33094 C10_P_btm.n1652 C10_P_btm.t400 1.67819
R33095 C10_P_btm.n1655 C10_P_btm.t642 1.67819
R33096 C10_P_btm.n1658 C10_P_btm.t923 1.67819
R33097 C10_P_btm.n1661 C10_P_btm.t585 1.67819
R33098 C10_P_btm.n1664 C10_P_btm.t818 1.67819
R33099 C10_P_btm.n1667 C10_P_btm.t54 1.67819
R33100 C10_P_btm.n1284 C10_P_btm.t130 1.67819
R33101 C10_P_btm.n1282 C10_P_btm.t913 1.67819
R33102 C10_P_btm.n1279 C10_P_btm.t687 1.67819
R33103 C10_P_btm.n1276 C10_P_btm.t1016 1.67819
R33104 C10_P_btm.n1273 C10_P_btm.t737 1.67819
R33105 C10_P_btm.n1270 C10_P_btm.t1029 1.67819
R33106 C10_P_btm.n1267 C10_P_btm.t846 1.67819
R33107 C10_P_btm.n1264 C10_P_btm.t553 1.67819
R33108 C10_P_btm.n1261 C10_P_btm.t900 1.67819
R33109 C10_P_btm.n1258 C10_P_btm.t671 1.67819
R33110 C10_P_btm.n1255 C10_P_btm.t436 1.67819
R33111 C10_P_btm.n1252 C10_P_btm.t720 1.67819
R33112 C10_P_btm.n1249 C10_P_btm.t516 1.67819
R33113 C10_P_btm.n1246 C10_P_btm.t256 1.67819
R33114 C10_P_btm.n1243 C10_P_btm.t537 1.67819
R33115 C10_P_btm.n1240 C10_P_btm.t304 1.67819
R33116 C10_P_btm.n1237 C10_P_btm.t650 1.67819
R33117 C10_P_btm.n1234 C10_P_btm.t365 1.67819
R33118 C10_P_btm.n1231 C10_P_btm.t135 1.67819
R33119 C10_P_btm.n1228 C10_P_btm.t471 1.67819
R33120 C10_P_btm.n1225 C10_P_btm.t630 1.67819
R33121 C10_P_btm.n1222 C10_P_btm.t1022 1.67819
R33122 C10_P_btm.n1219 C10_P_btm.t254 1.67819
R33123 C10_P_btm.n1216 C10_P_btm.t33 1.67819
R33124 C10_P_btm.n1213 C10_P_btm.t811 1.67819
R33125 C10_P_btm.n1210 C10_P_btm.t86 1.67819
R33126 C10_P_btm.n1207 C10_P_btm.t915 1.67819
R33127 C10_P_btm.n1204 C10_P_btm.t132 1.67819
R33128 C10_P_btm.n1201 C10_P_btm.t969 1.67819
R33129 C10_P_btm.n1198 C10_P_btm.t738 1.67819
R33130 C10_P_btm.n1195 C10_P_btm.t531 1.67819
R33131 C10_P_btm.n1192 C10_P_btm.t798 1.67819
R33132 C10_P_btm.n1189 C10_P_btm.t555 1.67819
R33133 C10_P_btm.n1186 C10_P_btm.t902 1.67819
R33134 C10_P_btm.n1183 C10_P_btm.t621 1.67819
R33135 C10_P_btm.n1180 C10_P_btm.t953 1.67819
R33136 C10_P_btm.n1177 C10_P_btm.t723 1.67819
R33137 C10_P_btm.n1174 C10_P_btm.t441 1.67819
R33138 C10_P_btm.n1171 C10_P_btm.t782 1.67819
R33139 C10_P_btm.n1168 C10_P_btm.t539 1.67819
R33140 C10_P_btm.n1165 C10_P_btm.t306 1.67819
R33141 C10_P_btm.n1162 C10_P_btm.t598 1.67819
R33142 C10_P_btm.n1159 C10_P_btm.t367 1.67819
R33143 C10_P_btm.n1156 C10_P_btm.t708 1.67819
R33144 C10_P_btm.n1153 C10_P_btm.t418 1.67819
R33145 C10_P_btm.n1150 C10_P_btm.t190 1.67819
R33146 C10_P_btm.n1147 C10_P_btm.t524 1.67819
R33147 C10_P_btm.n1144 C10_P_btm.t1030 1.67819
R33148 C10_P_btm.n1141 C10_P_btm.t108 1.67819
R33149 C10_P_btm.n1138 C10_P_btm.t269 1.67819
R33150 C10_P_btm.n1135 C10_P_btm.t100 1.67819
R33151 C10_P_btm.n1132 C10_P_btm.t825 1.67819
R33152 C10_P_btm.n1129 C10_P_btm.t106 1.67819
R33153 C10_P_btm.n1126 C10_P_btm.t926 1.67819
R33154 C10_P_btm.n1123 C10_P_btm.t149 1.67819
R33155 C10_P_btm.n1120 C10_P_btm.t981 1.67819
R33156 C10_P_btm.n1117 C10_P_btm.t750 1.67819
R33157 C10_P_btm.n1114 C10_P_btm.t46 1.67819
R33158 C10_P_btm.n1111 C10_P_btm.t810 1.67819
R33159 C10_P_btm.n1108 C10_P_btm.t571 1.67819
R33160 C10_P_btm.n1105 C10_P_btm.t914 1.67819
R33161 C10_P_btm.n1478 C10_P_btm.t636 1.67819
R33162 C10_P_btm.n1473 C10_P_btm.t76 1.67819
R33163 C10_P_btm.n1470 C10_P_btm.t352 1.67819
R33164 C10_P_btm.n1467 C10_P_btm.t219 1.67819
R33165 C10_P_btm.n1464 C10_P_btm.t249 1.67819
R33166 C10_P_btm.n1461 C10_P_btm.t481 1.67819
R33167 C10_P_btm.n1458 C10_P_btm.t193 1.67819
R33168 C10_P_btm.n1455 C10_P_btm.t422 1.67819
R33169 C10_P_btm.n1452 C10_P_btm.t654 1.67819
R33170 C10_P_btm.n1449 C10_P_btm.t370 1.67819
R33171 C10_P_btm.n1446 C10_P_btm.t601 1.67819
R33172 C10_P_btm.n1443 C10_P_btm.t259 1.67819
R33173 C10_P_btm.n1440 C10_P_btm.t542 1.67819
R33174 C10_P_btm.n1437 C10_P_btm.t785 1.67819
R33175 C10_P_btm.n1434 C10_P_btm.t722 1.67819
R33176 C10_P_btm.n1431 C10_P_btm.t952 1.67819
R33177 C10_P_btm.n1428 C10_P_btm.t175 1.67819
R33178 C10_P_btm.n1425 C10_P_btm.t901 1.67819
R33179 C10_P_btm.n1422 C10_P_btm.t68 1.67819
R33180 C10_P_btm.n1419 C10_P_btm.t347 1.67819
R33181 C10_P_btm.n1416 C10_P_btm.t44 1.67819
R33182 C10_P_btm.n1413 C10_P_btm.t501 1.67819
R33183 C10_P_btm.n1410 C10_P_btm.t1017 1.67819
R33184 C10_P_btm.n1407 C10_P_btm.t187 1.67819
R33185 C10_P_btm.n1404 C10_P_btm.t411 1.67819
R33186 C10_P_btm.n1401 C10_P_btm.t84 1.67819
R33187 C10_P_btm.n1398 C10_P_btm.t359 1.67819
R33188 C10_P_btm.n1395 C10_P_btm.t591 1.67819
R33189 C10_P_btm.n1392 C10_P_btm.t253 1.67819
R33190 C10_P_btm.n1389 C10_P_btm.t534 1.67819
R33191 C10_P_btm.n1386 C10_P_btm.t201 1.67819
R33192 C10_P_btm.n1383 C10_P_btm.t430 1.67819
R33193 C10_P_btm.n1380 C10_P_btm.t717 1.67819
R33194 C10_P_btm.n1377 C10_P_btm.t376 1.67819
R33195 C10_P_btm.n1374 C10_P_btm.t612 1.67819
R33196 C10_P_btm.n1371 C10_P_btm.t842 1.67819
R33197 C10_P_btm.n1368 C10_P_btm.t547 1.67819
R33198 C10_P_btm.n1365 C10_P_btm.t794 1.67819
R33199 C10_P_btm.n1362 C10_P_btm.t450 1.67819
R33200 C10_P_btm.n1359 C10_P_btm.t732 1.67819
R33201 C10_P_btm.n1356 C10_P_btm.t960 1.67819
R33202 C10_P_btm.n1353 C10_P_btm.t667 1.67819
R33203 C10_P_btm.n1350 C10_P_btm.t947 1.67819
R33204 C10_P_btm.n1347 C10_P_btm.t498 1.67819
R33205 C10_P_btm.n1344 C10_P_btm.t843 1.67819
R33206 C10_P_btm.n1341 C10_P_btm.t95 1.67819
R33207 C10_P_btm.n1338 C10_P_btm.t283 1.67819
R33208 C10_P_btm.n1335 C10_P_btm.t1013 1.67819
R33209 C10_P_btm.n1332 C10_P_btm.t90 1.67819
R33210 C10_P_btm.n1329 C10_P_btm.t963 1.67819
R33211 C10_P_btm.n1326 C10_P_btm.t128 1.67819
R33212 C10_P_btm.n1323 C10_P_btm.t356 1.67819
R33213 C10_P_btm.n1320 C10_P_btm.t80 1.67819
R33214 C10_P_btm.n1317 C10_P_btm.t297 1.67819
R33215 C10_P_btm.n1314 C10_P_btm.t1055 1.67819
R33216 C10_P_btm.n1311 C10_P_btm.t199 1.67819
R33217 C10_P_btm.n1308 C10_P_btm.t493 1.67819
R33218 C10_P_btm.n1305 C10_P_btm.t144 1.67819
R33219 C10_P_btm.n1302 C10_P_btm.t89 1.67819
R33220 C10_P_btm.n1299 C10_P_btm.t662 1.67819
R33221 C10_P_btm.n1296 C10_P_btm.t316 1.67819
R33222 C10_P_btm.n1293 C10_P_btm.t545 1.67819
R33223 C10_P_btm.n1290 C10_P_btm.t840 1.67819
R33224 C10_P_btm.n507 C10_P_btm.n506 1.05569
R33225 C10_P_btm.n3038 C10_P_btm.n524 1.05569
R33226 C10_P_btm.n1288 C10_P_btm.n918 1.05569
R33227 C10_P_btm.n1476 C10_P_btm.n1475 1.05569
R33228 C10_P_btm.n44 C10_P_btm.n42 1.0005
R33229 C10_P_btm.n45 C10_P_btm.n41 1.0005
R33230 C10_P_btm.n46 C10_P_btm.n40 1.0005
R33231 C10_P_btm.n47 C10_P_btm.n39 1.0005
R33232 C10_P_btm.n48 C10_P_btm.n38 1.0005
R33233 C10_P_btm.n49 C10_P_btm.n37 1.0005
R33234 C10_P_btm.n50 C10_P_btm.n36 1.0005
R33235 C10_P_btm.n51 C10_P_btm.n35 1.0005
R33236 C10_P_btm.n3835 C10_P_btm.n34 1.0005
R33237 C10_P_btm.n3835 C10_P_btm.n3834 1.0005
R33238 C10_P_btm.n54 C10_P_btm.n51 1.0005
R33239 C10_P_btm.n55 C10_P_btm.n50 1.0005
R33240 C10_P_btm.n56 C10_P_btm.n49 1.0005
R33241 C10_P_btm.n57 C10_P_btm.n48 1.0005
R33242 C10_P_btm.n58 C10_P_btm.n47 1.0005
R33243 C10_P_btm.n59 C10_P_btm.n46 1.0005
R33244 C10_P_btm.n60 C10_P_btm.n45 1.0005
R33245 C10_P_btm.n3806 C10_P_btm.n44 1.0005
R33246 C10_P_btm.n3806 C10_P_btm.n3805 1.0005
R33247 C10_P_btm.n3743 C10_P_btm.n60 1.0005
R33248 C10_P_btm.n3742 C10_P_btm.n59 1.0005
R33249 C10_P_btm.n3741 C10_P_btm.n58 1.0005
R33250 C10_P_btm.n3740 C10_P_btm.n57 1.0005
R33251 C10_P_btm.n3739 C10_P_btm.n56 1.0005
R33252 C10_P_btm.n3738 C10_P_btm.n55 1.0005
R33253 C10_P_btm.n3737 C10_P_btm.n54 1.0005
R33254 C10_P_btm.n3834 C10_P_btm.n52 1.0005
R33255 C10_P_btm.n71 C10_P_btm.n52 1.0005
R33256 C10_P_btm.n3737 C10_P_btm.n70 1.0005
R33257 C10_P_btm.n3738 C10_P_btm.n69 1.0005
R33258 C10_P_btm.n3739 C10_P_btm.n68 1.0005
R33259 C10_P_btm.n3740 C10_P_btm.n67 1.0005
R33260 C10_P_btm.n3741 C10_P_btm.n66 1.0005
R33261 C10_P_btm.n3742 C10_P_btm.n65 1.0005
R33262 C10_P_btm.n3743 C10_P_btm.n64 1.0005
R33263 C10_P_btm.n3805 C10_P_btm.n61 1.0005
R33264 C10_P_btm.n3704 C10_P_btm.n61 1.0005
R33265 C10_P_btm.n80 C10_P_btm.n64 1.0005
R33266 C10_P_btm.n79 C10_P_btm.n65 1.0005
R33267 C10_P_btm.n78 C10_P_btm.n66 1.0005
R33268 C10_P_btm.n77 C10_P_btm.n67 1.0005
R33269 C10_P_btm.n76 C10_P_btm.n68 1.0005
R33270 C10_P_btm.n75 C10_P_btm.n69 1.0005
R33271 C10_P_btm.n74 C10_P_btm.n70 1.0005
R33272 C10_P_btm.n73 C10_P_btm.n71 1.0005
R33273 C10_P_btm.n123 C10_P_btm.n73 1.0005
R33274 C10_P_btm.n93 C10_P_btm.n74 1.0005
R33275 C10_P_btm.n94 C10_P_btm.n75 1.0005
R33276 C10_P_btm.n95 C10_P_btm.n76 1.0005
R33277 C10_P_btm.n96 C10_P_btm.n77 1.0005
R33278 C10_P_btm.n97 C10_P_btm.n78 1.0005
R33279 C10_P_btm.n98 C10_P_btm.n79 1.0005
R33280 C10_P_btm.n99 C10_P_btm.n80 1.0005
R33281 C10_P_btm.n3704 C10_P_btm.n3703 1.0005
R33282 C10_P_btm.n3703 C10_P_btm.n81 1.0005
R33283 C10_P_btm.n99 C10_P_btm.n84 1.0005
R33284 C10_P_btm.n98 C10_P_btm.n85 1.0005
R33285 C10_P_btm.n97 C10_P_btm.n86 1.0005
R33286 C10_P_btm.n96 C10_P_btm.n87 1.0005
R33287 C10_P_btm.n95 C10_P_btm.n88 1.0005
R33288 C10_P_btm.n94 C10_P_btm.n89 1.0005
R33289 C10_P_btm.n93 C10_P_btm.n90 1.0005
R33290 C10_P_btm.n124 C10_P_btm.n123 1.0005
R33291 C10_P_btm.n126 C10_P_btm.n124 1.0005
R33292 C10_P_btm.n127 C10_P_btm.n90 1.0005
R33293 C10_P_btm.n128 C10_P_btm.n89 1.0005
R33294 C10_P_btm.n129 C10_P_btm.n88 1.0005
R33295 C10_P_btm.n130 C10_P_btm.n87 1.0005
R33296 C10_P_btm.n131 C10_P_btm.n86 1.0005
R33297 C10_P_btm.n132 C10_P_btm.n85 1.0005
R33298 C10_P_btm.n133 C10_P_btm.n84 1.0005
R33299 C10_P_btm.n3637 C10_P_btm.n81 1.0005
R33300 C10_P_btm.n3637 C10_P_btm.n3636 1.0005
R33301 C10_P_btm.n152 C10_P_btm.n133 1.0005
R33302 C10_P_btm.n151 C10_P_btm.n132 1.0005
R33303 C10_P_btm.n150 C10_P_btm.n131 1.0005
R33304 C10_P_btm.n149 C10_P_btm.n130 1.0005
R33305 C10_P_btm.n148 C10_P_btm.n129 1.0005
R33306 C10_P_btm.n147 C10_P_btm.n128 1.0005
R33307 C10_P_btm.n146 C10_P_btm.n127 1.0005
R33308 C10_P_btm.n176 C10_P_btm.n126 1.0005
R33309 C10_P_btm.n177 C10_P_btm.n176 1.0005
R33310 C10_P_btm.n146 C10_P_btm.n143 1.0005
R33311 C10_P_btm.n147 C10_P_btm.n142 1.0005
R33312 C10_P_btm.n148 C10_P_btm.n141 1.0005
R33313 C10_P_btm.n149 C10_P_btm.n140 1.0005
R33314 C10_P_btm.n150 C10_P_btm.n139 1.0005
R33315 C10_P_btm.n151 C10_P_btm.n138 1.0005
R33316 C10_P_btm.n152 C10_P_btm.n137 1.0005
R33317 C10_P_btm.n3636 C10_P_btm.n134 1.0005
R33318 C10_P_btm.n3570 C10_P_btm.n134 1.0005
R33319 C10_P_btm.n186 C10_P_btm.n137 1.0005
R33320 C10_P_btm.n185 C10_P_btm.n138 1.0005
R33321 C10_P_btm.n184 C10_P_btm.n139 1.0005
R33322 C10_P_btm.n183 C10_P_btm.n140 1.0005
R33323 C10_P_btm.n182 C10_P_btm.n141 1.0005
R33324 C10_P_btm.n181 C10_P_btm.n142 1.0005
R33325 C10_P_btm.n180 C10_P_btm.n143 1.0005
R33326 C10_P_btm.n179 C10_P_btm.n177 1.0005
R33327 C10_P_btm.n229 C10_P_btm.n179 1.0005
R33328 C10_P_btm.n199 C10_P_btm.n180 1.0005
R33329 C10_P_btm.n200 C10_P_btm.n181 1.0005
R33330 C10_P_btm.n201 C10_P_btm.n182 1.0005
R33331 C10_P_btm.n202 C10_P_btm.n183 1.0005
R33332 C10_P_btm.n203 C10_P_btm.n184 1.0005
R33333 C10_P_btm.n204 C10_P_btm.n185 1.0005
R33334 C10_P_btm.n205 C10_P_btm.n186 1.0005
R33335 C10_P_btm.n3570 C10_P_btm.n3569 1.0005
R33336 C10_P_btm.n3569 C10_P_btm.n187 1.0005
R33337 C10_P_btm.n205 C10_P_btm.n190 1.0005
R33338 C10_P_btm.n204 C10_P_btm.n191 1.0005
R33339 C10_P_btm.n203 C10_P_btm.n192 1.0005
R33340 C10_P_btm.n202 C10_P_btm.n193 1.0005
R33341 C10_P_btm.n201 C10_P_btm.n194 1.0005
R33342 C10_P_btm.n200 C10_P_btm.n195 1.0005
R33343 C10_P_btm.n199 C10_P_btm.n196 1.0005
R33344 C10_P_btm.n230 C10_P_btm.n229 1.0005
R33345 C10_P_btm.n232 C10_P_btm.n230 1.0005
R33346 C10_P_btm.n233 C10_P_btm.n196 1.0005
R33347 C10_P_btm.n234 C10_P_btm.n195 1.0005
R33348 C10_P_btm.n235 C10_P_btm.n194 1.0005
R33349 C10_P_btm.n236 C10_P_btm.n193 1.0005
R33350 C10_P_btm.n237 C10_P_btm.n192 1.0005
R33351 C10_P_btm.n238 C10_P_btm.n191 1.0005
R33352 C10_P_btm.n239 C10_P_btm.n190 1.0005
R33353 C10_P_btm.n3503 C10_P_btm.n187 1.0005
R33354 C10_P_btm.n3503 C10_P_btm.n3502 1.0005
R33355 C10_P_btm.n258 C10_P_btm.n239 1.0005
R33356 C10_P_btm.n257 C10_P_btm.n238 1.0005
R33357 C10_P_btm.n256 C10_P_btm.n237 1.0005
R33358 C10_P_btm.n255 C10_P_btm.n236 1.0005
R33359 C10_P_btm.n254 C10_P_btm.n235 1.0005
R33360 C10_P_btm.n253 C10_P_btm.n234 1.0005
R33361 C10_P_btm.n252 C10_P_btm.n233 1.0005
R33362 C10_P_btm.n282 C10_P_btm.n232 1.0005
R33363 C10_P_btm.n283 C10_P_btm.n282 1.0005
R33364 C10_P_btm.n252 C10_P_btm.n249 1.0005
R33365 C10_P_btm.n253 C10_P_btm.n248 1.0005
R33366 C10_P_btm.n254 C10_P_btm.n247 1.0005
R33367 C10_P_btm.n255 C10_P_btm.n246 1.0005
R33368 C10_P_btm.n256 C10_P_btm.n245 1.0005
R33369 C10_P_btm.n257 C10_P_btm.n244 1.0005
R33370 C10_P_btm.n258 C10_P_btm.n243 1.0005
R33371 C10_P_btm.n3502 C10_P_btm.n240 1.0005
R33372 C10_P_btm.n3436 C10_P_btm.n240 1.0005
R33373 C10_P_btm.n292 C10_P_btm.n243 1.0005
R33374 C10_P_btm.n291 C10_P_btm.n244 1.0005
R33375 C10_P_btm.n290 C10_P_btm.n245 1.0005
R33376 C10_P_btm.n289 C10_P_btm.n246 1.0005
R33377 C10_P_btm.n288 C10_P_btm.n247 1.0005
R33378 C10_P_btm.n287 C10_P_btm.n248 1.0005
R33379 C10_P_btm.n286 C10_P_btm.n249 1.0005
R33380 C10_P_btm.n285 C10_P_btm.n283 1.0005
R33381 C10_P_btm.n335 C10_P_btm.n285 1.0005
R33382 C10_P_btm.n305 C10_P_btm.n286 1.0005
R33383 C10_P_btm.n306 C10_P_btm.n287 1.0005
R33384 C10_P_btm.n307 C10_P_btm.n288 1.0005
R33385 C10_P_btm.n308 C10_P_btm.n289 1.0005
R33386 C10_P_btm.n309 C10_P_btm.n290 1.0005
R33387 C10_P_btm.n310 C10_P_btm.n291 1.0005
R33388 C10_P_btm.n311 C10_P_btm.n292 1.0005
R33389 C10_P_btm.n3436 C10_P_btm.n3435 1.0005
R33390 C10_P_btm.n3435 C10_P_btm.n293 1.0005
R33391 C10_P_btm.n311 C10_P_btm.n296 1.0005
R33392 C10_P_btm.n310 C10_P_btm.n297 1.0005
R33393 C10_P_btm.n309 C10_P_btm.n298 1.0005
R33394 C10_P_btm.n308 C10_P_btm.n299 1.0005
R33395 C10_P_btm.n307 C10_P_btm.n300 1.0005
R33396 C10_P_btm.n306 C10_P_btm.n301 1.0005
R33397 C10_P_btm.n305 C10_P_btm.n302 1.0005
R33398 C10_P_btm.n336 C10_P_btm.n335 1.0005
R33399 C10_P_btm.n338 C10_P_btm.n336 1.0005
R33400 C10_P_btm.n339 C10_P_btm.n302 1.0005
R33401 C10_P_btm.n340 C10_P_btm.n301 1.0005
R33402 C10_P_btm.n341 C10_P_btm.n300 1.0005
R33403 C10_P_btm.n342 C10_P_btm.n299 1.0005
R33404 C10_P_btm.n343 C10_P_btm.n298 1.0005
R33405 C10_P_btm.n344 C10_P_btm.n297 1.0005
R33406 C10_P_btm.n345 C10_P_btm.n296 1.0005
R33407 C10_P_btm.n3369 C10_P_btm.n293 1.0005
R33408 C10_P_btm.n3369 C10_P_btm.n3368 1.0005
R33409 C10_P_btm.n364 C10_P_btm.n345 1.0005
R33410 C10_P_btm.n363 C10_P_btm.n344 1.0005
R33411 C10_P_btm.n362 C10_P_btm.n343 1.0005
R33412 C10_P_btm.n361 C10_P_btm.n342 1.0005
R33413 C10_P_btm.n360 C10_P_btm.n341 1.0005
R33414 C10_P_btm.n359 C10_P_btm.n340 1.0005
R33415 C10_P_btm.n358 C10_P_btm.n339 1.0005
R33416 C10_P_btm.n388 C10_P_btm.n338 1.0005
R33417 C10_P_btm.n389 C10_P_btm.n388 1.0005
R33418 C10_P_btm.n358 C10_P_btm.n355 1.0005
R33419 C10_P_btm.n359 C10_P_btm.n354 1.0005
R33420 C10_P_btm.n360 C10_P_btm.n353 1.0005
R33421 C10_P_btm.n361 C10_P_btm.n352 1.0005
R33422 C10_P_btm.n362 C10_P_btm.n351 1.0005
R33423 C10_P_btm.n363 C10_P_btm.n350 1.0005
R33424 C10_P_btm.n364 C10_P_btm.n349 1.0005
R33425 C10_P_btm.n3368 C10_P_btm.n346 1.0005
R33426 C10_P_btm.n3302 C10_P_btm.n346 1.0005
R33427 C10_P_btm.n398 C10_P_btm.n349 1.0005
R33428 C10_P_btm.n397 C10_P_btm.n350 1.0005
R33429 C10_P_btm.n396 C10_P_btm.n351 1.0005
R33430 C10_P_btm.n395 C10_P_btm.n352 1.0005
R33431 C10_P_btm.n394 C10_P_btm.n353 1.0005
R33432 C10_P_btm.n393 C10_P_btm.n354 1.0005
R33433 C10_P_btm.n392 C10_P_btm.n355 1.0005
R33434 C10_P_btm.n391 C10_P_btm.n389 1.0005
R33435 C10_P_btm.n435 C10_P_btm.n391 1.0005
R33436 C10_P_btm.n436 C10_P_btm.n392 1.0005
R33437 C10_P_btm.n437 C10_P_btm.n393 1.0005
R33438 C10_P_btm.n438 C10_P_btm.n394 1.0005
R33439 C10_P_btm.n439 C10_P_btm.n395 1.0005
R33440 C10_P_btm.n440 C10_P_btm.n396 1.0005
R33441 C10_P_btm.n441 C10_P_btm.n397 1.0005
R33442 C10_P_btm.n442 C10_P_btm.n398 1.0005
R33443 C10_P_btm.n3302 C10_P_btm.n3301 1.0005
R33444 C10_P_btm.n3301 C10_P_btm.n399 1.0005
R33445 C10_P_btm.n442 C10_P_btm.n402 1.0005
R33446 C10_P_btm.n441 C10_P_btm.n403 1.0005
R33447 C10_P_btm.n440 C10_P_btm.n404 1.0005
R33448 C10_P_btm.n439 C10_P_btm.n405 1.0005
R33449 C10_P_btm.n438 C10_P_btm.n406 1.0005
R33450 C10_P_btm.n437 C10_P_btm.n407 1.0005
R33451 C10_P_btm.n436 C10_P_btm.n408 1.0005
R33452 C10_P_btm.n435 C10_P_btm.n409 1.0005
R33453 C10_P_btm.n410 C10_P_btm.n390 1.0005
R33454 C10_P_btm.n423 C10_P_btm.n422 1.0005
R33455 C10_P_btm.n424 C10_P_btm.n421 1.0005
R33456 C10_P_btm.n425 C10_P_btm.n420 1.0005
R33457 C10_P_btm.n426 C10_P_btm.n419 1.0005
R33458 C10_P_btm.n427 C10_P_btm.n418 1.0005
R33459 C10_P_btm.n428 C10_P_btm.n417 1.0005
R33460 C10_P_btm.n429 C10_P_btm.n416 1.0005
R33461 C10_P_btm.n430 C10_P_btm.n415 1.0005
R33462 C10_P_btm.n431 C10_P_btm.n414 1.0005
R33463 C10_P_btm.n432 C10_P_btm.n413 1.0005
R33464 C10_P_btm.n433 C10_P_btm.n412 1.0005
R33465 C10_P_btm.n434 C10_P_btm.n411 1.0005
R33466 C10_P_btm.n2057 C10_P_btm.n546 1.0005
R33467 C10_P_btm.n2058 C10_P_btm.n545 1.0005
R33468 C10_P_btm.n2059 C10_P_btm.n544 1.0005
R33469 C10_P_btm.n2060 C10_P_btm.n543 1.0005
R33470 C10_P_btm.n2061 C10_P_btm.n542 1.0005
R33471 C10_P_btm.n2062 C10_P_btm.n541 1.0005
R33472 C10_P_btm.n2063 C10_P_btm.n540 1.0005
R33473 C10_P_btm.n2064 C10_P_btm.n539 1.0005
R33474 C10_P_btm.n2065 C10_P_btm.n538 1.0005
R33475 C10_P_btm.n2067 C10_P_btm.n2065 1.0005
R33476 C10_P_btm.n2068 C10_P_btm.n2064 1.0005
R33477 C10_P_btm.n2069 C10_P_btm.n2063 1.0005
R33478 C10_P_btm.n2070 C10_P_btm.n2062 1.0005
R33479 C10_P_btm.n2071 C10_P_btm.n2061 1.0005
R33480 C10_P_btm.n2072 C10_P_btm.n2060 1.0005
R33481 C10_P_btm.n2073 C10_P_btm.n2059 1.0005
R33482 C10_P_btm.n2074 C10_P_btm.n2058 1.0005
R33483 C10_P_btm.n2994 C10_P_btm.n2057 1.0005
R33484 C10_P_btm.n2994 C10_P_btm.n2993 1.0005
R33485 C10_P_btm.n2077 C10_P_btm.n2074 1.0005
R33486 C10_P_btm.n2078 C10_P_btm.n2073 1.0005
R33487 C10_P_btm.n2079 C10_P_btm.n2072 1.0005
R33488 C10_P_btm.n2080 C10_P_btm.n2071 1.0005
R33489 C10_P_btm.n2081 C10_P_btm.n2070 1.0005
R33490 C10_P_btm.n2082 C10_P_btm.n2069 1.0005
R33491 C10_P_btm.n2083 C10_P_btm.n2068 1.0005
R33492 C10_P_btm.n2965 C10_P_btm.n2067 1.0005
R33493 C10_P_btm.n2965 C10_P_btm.n2964 1.0005
R33494 C10_P_btm.n2902 C10_P_btm.n2083 1.0005
R33495 C10_P_btm.n2901 C10_P_btm.n2082 1.0005
R33496 C10_P_btm.n2900 C10_P_btm.n2081 1.0005
R33497 C10_P_btm.n2899 C10_P_btm.n2080 1.0005
R33498 C10_P_btm.n2898 C10_P_btm.n2079 1.0005
R33499 C10_P_btm.n2897 C10_P_btm.n2078 1.0005
R33500 C10_P_btm.n2896 C10_P_btm.n2077 1.0005
R33501 C10_P_btm.n2993 C10_P_btm.n2075 1.0005
R33502 C10_P_btm.n2094 C10_P_btm.n2075 1.0005
R33503 C10_P_btm.n2896 C10_P_btm.n2093 1.0005
R33504 C10_P_btm.n2897 C10_P_btm.n2092 1.0005
R33505 C10_P_btm.n2898 C10_P_btm.n2091 1.0005
R33506 C10_P_btm.n2899 C10_P_btm.n2090 1.0005
R33507 C10_P_btm.n2900 C10_P_btm.n2089 1.0005
R33508 C10_P_btm.n2901 C10_P_btm.n2088 1.0005
R33509 C10_P_btm.n2902 C10_P_btm.n2087 1.0005
R33510 C10_P_btm.n2964 C10_P_btm.n2084 1.0005
R33511 C10_P_btm.n2863 C10_P_btm.n2084 1.0005
R33512 C10_P_btm.n2103 C10_P_btm.n2087 1.0005
R33513 C10_P_btm.n2102 C10_P_btm.n2088 1.0005
R33514 C10_P_btm.n2101 C10_P_btm.n2089 1.0005
R33515 C10_P_btm.n2100 C10_P_btm.n2090 1.0005
R33516 C10_P_btm.n2099 C10_P_btm.n2091 1.0005
R33517 C10_P_btm.n2098 C10_P_btm.n2092 1.0005
R33518 C10_P_btm.n2097 C10_P_btm.n2093 1.0005
R33519 C10_P_btm.n2096 C10_P_btm.n2094 1.0005
R33520 C10_P_btm.n2146 C10_P_btm.n2096 1.0005
R33521 C10_P_btm.n2116 C10_P_btm.n2097 1.0005
R33522 C10_P_btm.n2117 C10_P_btm.n2098 1.0005
R33523 C10_P_btm.n2118 C10_P_btm.n2099 1.0005
R33524 C10_P_btm.n2119 C10_P_btm.n2100 1.0005
R33525 C10_P_btm.n2120 C10_P_btm.n2101 1.0005
R33526 C10_P_btm.n2121 C10_P_btm.n2102 1.0005
R33527 C10_P_btm.n2122 C10_P_btm.n2103 1.0005
R33528 C10_P_btm.n2863 C10_P_btm.n2862 1.0005
R33529 C10_P_btm.n2862 C10_P_btm.n2104 1.0005
R33530 C10_P_btm.n2122 C10_P_btm.n2107 1.0005
R33531 C10_P_btm.n2121 C10_P_btm.n2108 1.0005
R33532 C10_P_btm.n2120 C10_P_btm.n2109 1.0005
R33533 C10_P_btm.n2119 C10_P_btm.n2110 1.0005
R33534 C10_P_btm.n2118 C10_P_btm.n2111 1.0005
R33535 C10_P_btm.n2117 C10_P_btm.n2112 1.0005
R33536 C10_P_btm.n2116 C10_P_btm.n2113 1.0005
R33537 C10_P_btm.n2147 C10_P_btm.n2146 1.0005
R33538 C10_P_btm.n2149 C10_P_btm.n2147 1.0005
R33539 C10_P_btm.n2150 C10_P_btm.n2113 1.0005
R33540 C10_P_btm.n2151 C10_P_btm.n2112 1.0005
R33541 C10_P_btm.n2152 C10_P_btm.n2111 1.0005
R33542 C10_P_btm.n2153 C10_P_btm.n2110 1.0005
R33543 C10_P_btm.n2154 C10_P_btm.n2109 1.0005
R33544 C10_P_btm.n2155 C10_P_btm.n2108 1.0005
R33545 C10_P_btm.n2156 C10_P_btm.n2107 1.0005
R33546 C10_P_btm.n2796 C10_P_btm.n2104 1.0005
R33547 C10_P_btm.n2796 C10_P_btm.n2795 1.0005
R33548 C10_P_btm.n2175 C10_P_btm.n2156 1.0005
R33549 C10_P_btm.n2174 C10_P_btm.n2155 1.0005
R33550 C10_P_btm.n2173 C10_P_btm.n2154 1.0005
R33551 C10_P_btm.n2172 C10_P_btm.n2153 1.0005
R33552 C10_P_btm.n2171 C10_P_btm.n2152 1.0005
R33553 C10_P_btm.n2170 C10_P_btm.n2151 1.0005
R33554 C10_P_btm.n2169 C10_P_btm.n2150 1.0005
R33555 C10_P_btm.n2199 C10_P_btm.n2149 1.0005
R33556 C10_P_btm.n2200 C10_P_btm.n2199 1.0005
R33557 C10_P_btm.n2169 C10_P_btm.n2166 1.0005
R33558 C10_P_btm.n2170 C10_P_btm.n2165 1.0005
R33559 C10_P_btm.n2171 C10_P_btm.n2164 1.0005
R33560 C10_P_btm.n2172 C10_P_btm.n2163 1.0005
R33561 C10_P_btm.n2173 C10_P_btm.n2162 1.0005
R33562 C10_P_btm.n2174 C10_P_btm.n2161 1.0005
R33563 C10_P_btm.n2175 C10_P_btm.n2160 1.0005
R33564 C10_P_btm.n2795 C10_P_btm.n2157 1.0005
R33565 C10_P_btm.n2729 C10_P_btm.n2157 1.0005
R33566 C10_P_btm.n2209 C10_P_btm.n2160 1.0005
R33567 C10_P_btm.n2208 C10_P_btm.n2161 1.0005
R33568 C10_P_btm.n2207 C10_P_btm.n2162 1.0005
R33569 C10_P_btm.n2206 C10_P_btm.n2163 1.0005
R33570 C10_P_btm.n2205 C10_P_btm.n2164 1.0005
R33571 C10_P_btm.n2204 C10_P_btm.n2165 1.0005
R33572 C10_P_btm.n2203 C10_P_btm.n2166 1.0005
R33573 C10_P_btm.n2202 C10_P_btm.n2200 1.0005
R33574 C10_P_btm.n2252 C10_P_btm.n2202 1.0005
R33575 C10_P_btm.n2222 C10_P_btm.n2203 1.0005
R33576 C10_P_btm.n2223 C10_P_btm.n2204 1.0005
R33577 C10_P_btm.n2224 C10_P_btm.n2205 1.0005
R33578 C10_P_btm.n2225 C10_P_btm.n2206 1.0005
R33579 C10_P_btm.n2226 C10_P_btm.n2207 1.0005
R33580 C10_P_btm.n2227 C10_P_btm.n2208 1.0005
R33581 C10_P_btm.n2228 C10_P_btm.n2209 1.0005
R33582 C10_P_btm.n2729 C10_P_btm.n2728 1.0005
R33583 C10_P_btm.n2728 C10_P_btm.n2210 1.0005
R33584 C10_P_btm.n2228 C10_P_btm.n2213 1.0005
R33585 C10_P_btm.n2227 C10_P_btm.n2214 1.0005
R33586 C10_P_btm.n2226 C10_P_btm.n2215 1.0005
R33587 C10_P_btm.n2225 C10_P_btm.n2216 1.0005
R33588 C10_P_btm.n2224 C10_P_btm.n2217 1.0005
R33589 C10_P_btm.n2223 C10_P_btm.n2218 1.0005
R33590 C10_P_btm.n2222 C10_P_btm.n2219 1.0005
R33591 C10_P_btm.n2253 C10_P_btm.n2252 1.0005
R33592 C10_P_btm.n2255 C10_P_btm.n2253 1.0005
R33593 C10_P_btm.n2256 C10_P_btm.n2219 1.0005
R33594 C10_P_btm.n2257 C10_P_btm.n2218 1.0005
R33595 C10_P_btm.n2258 C10_P_btm.n2217 1.0005
R33596 C10_P_btm.n2259 C10_P_btm.n2216 1.0005
R33597 C10_P_btm.n2260 C10_P_btm.n2215 1.0005
R33598 C10_P_btm.n2261 C10_P_btm.n2214 1.0005
R33599 C10_P_btm.n2262 C10_P_btm.n2213 1.0005
R33600 C10_P_btm.n2662 C10_P_btm.n2210 1.0005
R33601 C10_P_btm.n2662 C10_P_btm.n2661 1.0005
R33602 C10_P_btm.n2281 C10_P_btm.n2262 1.0005
R33603 C10_P_btm.n2280 C10_P_btm.n2261 1.0005
R33604 C10_P_btm.n2279 C10_P_btm.n2260 1.0005
R33605 C10_P_btm.n2278 C10_P_btm.n2259 1.0005
R33606 C10_P_btm.n2277 C10_P_btm.n2258 1.0005
R33607 C10_P_btm.n2276 C10_P_btm.n2257 1.0005
R33608 C10_P_btm.n2275 C10_P_btm.n2256 1.0005
R33609 C10_P_btm.n2305 C10_P_btm.n2255 1.0005
R33610 C10_P_btm.n2306 C10_P_btm.n2305 1.0005
R33611 C10_P_btm.n2275 C10_P_btm.n2272 1.0005
R33612 C10_P_btm.n2276 C10_P_btm.n2271 1.0005
R33613 C10_P_btm.n2277 C10_P_btm.n2270 1.0005
R33614 C10_P_btm.n2278 C10_P_btm.n2269 1.0005
R33615 C10_P_btm.n2279 C10_P_btm.n2268 1.0005
R33616 C10_P_btm.n2280 C10_P_btm.n2267 1.0005
R33617 C10_P_btm.n2281 C10_P_btm.n2266 1.0005
R33618 C10_P_btm.n2661 C10_P_btm.n2263 1.0005
R33619 C10_P_btm.n2595 C10_P_btm.n2263 1.0005
R33620 C10_P_btm.n2315 C10_P_btm.n2266 1.0005
R33621 C10_P_btm.n2314 C10_P_btm.n2267 1.0005
R33622 C10_P_btm.n2313 C10_P_btm.n2268 1.0005
R33623 C10_P_btm.n2312 C10_P_btm.n2269 1.0005
R33624 C10_P_btm.n2311 C10_P_btm.n2270 1.0005
R33625 C10_P_btm.n2310 C10_P_btm.n2271 1.0005
R33626 C10_P_btm.n2309 C10_P_btm.n2272 1.0005
R33627 C10_P_btm.n2308 C10_P_btm.n2306 1.0005
R33628 C10_P_btm.n2358 C10_P_btm.n2308 1.0005
R33629 C10_P_btm.n2328 C10_P_btm.n2309 1.0005
R33630 C10_P_btm.n2329 C10_P_btm.n2310 1.0005
R33631 C10_P_btm.n2330 C10_P_btm.n2311 1.0005
R33632 C10_P_btm.n2331 C10_P_btm.n2312 1.0005
R33633 C10_P_btm.n2332 C10_P_btm.n2313 1.0005
R33634 C10_P_btm.n2333 C10_P_btm.n2314 1.0005
R33635 C10_P_btm.n2334 C10_P_btm.n2315 1.0005
R33636 C10_P_btm.n2595 C10_P_btm.n2594 1.0005
R33637 C10_P_btm.n2594 C10_P_btm.n2316 1.0005
R33638 C10_P_btm.n2334 C10_P_btm.n2319 1.0005
R33639 C10_P_btm.n2333 C10_P_btm.n2320 1.0005
R33640 C10_P_btm.n2332 C10_P_btm.n2321 1.0005
R33641 C10_P_btm.n2331 C10_P_btm.n2322 1.0005
R33642 C10_P_btm.n2330 C10_P_btm.n2323 1.0005
R33643 C10_P_btm.n2329 C10_P_btm.n2324 1.0005
R33644 C10_P_btm.n2328 C10_P_btm.n2325 1.0005
R33645 C10_P_btm.n2359 C10_P_btm.n2358 1.0005
R33646 C10_P_btm.n2361 C10_P_btm.n2359 1.0005
R33647 C10_P_btm.n2362 C10_P_btm.n2325 1.0005
R33648 C10_P_btm.n2363 C10_P_btm.n2324 1.0005
R33649 C10_P_btm.n2364 C10_P_btm.n2323 1.0005
R33650 C10_P_btm.n2365 C10_P_btm.n2322 1.0005
R33651 C10_P_btm.n2366 C10_P_btm.n2321 1.0005
R33652 C10_P_btm.n2367 C10_P_btm.n2320 1.0005
R33653 C10_P_btm.n2368 C10_P_btm.n2319 1.0005
R33654 C10_P_btm.n2528 C10_P_btm.n2316 1.0005
R33655 C10_P_btm.n2528 C10_P_btm.n2527 1.0005
R33656 C10_P_btm.n2387 C10_P_btm.n2368 1.0005
R33657 C10_P_btm.n2386 C10_P_btm.n2367 1.0005
R33658 C10_P_btm.n2385 C10_P_btm.n2366 1.0005
R33659 C10_P_btm.n2384 C10_P_btm.n2365 1.0005
R33660 C10_P_btm.n2383 C10_P_btm.n2364 1.0005
R33661 C10_P_btm.n2382 C10_P_btm.n2363 1.0005
R33662 C10_P_btm.n2381 C10_P_btm.n2362 1.0005
R33663 C10_P_btm.n2411 C10_P_btm.n2361 1.0005
R33664 C10_P_btm.n2412 C10_P_btm.n2411 1.0005
R33665 C10_P_btm.n2381 C10_P_btm.n2378 1.0005
R33666 C10_P_btm.n2382 C10_P_btm.n2377 1.0005
R33667 C10_P_btm.n2383 C10_P_btm.n2376 1.0005
R33668 C10_P_btm.n2384 C10_P_btm.n2375 1.0005
R33669 C10_P_btm.n2385 C10_P_btm.n2374 1.0005
R33670 C10_P_btm.n2386 C10_P_btm.n2373 1.0005
R33671 C10_P_btm.n2387 C10_P_btm.n2372 1.0005
R33672 C10_P_btm.n2527 C10_P_btm.n2369 1.0005
R33673 C10_P_btm.n2461 C10_P_btm.n2369 1.0005
R33674 C10_P_btm.n2421 C10_P_btm.n2372 1.0005
R33675 C10_P_btm.n2420 C10_P_btm.n2373 1.0005
R33676 C10_P_btm.n2419 C10_P_btm.n2374 1.0005
R33677 C10_P_btm.n2418 C10_P_btm.n2375 1.0005
R33678 C10_P_btm.n2417 C10_P_btm.n2376 1.0005
R33679 C10_P_btm.n2416 C10_P_btm.n2377 1.0005
R33680 C10_P_btm.n2415 C10_P_btm.n2378 1.0005
R33681 C10_P_btm.n2414 C10_P_btm.n2412 1.0005
R33682 C10_P_btm.n2429 C10_P_btm.n2414 1.0005
R33683 C10_P_btm.n2428 C10_P_btm.n2415 1.0005
R33684 C10_P_btm.n2427 C10_P_btm.n2416 1.0005
R33685 C10_P_btm.n2426 C10_P_btm.n2417 1.0005
R33686 C10_P_btm.n2425 C10_P_btm.n2418 1.0005
R33687 C10_P_btm.n2424 C10_P_btm.n2419 1.0005
R33688 C10_P_btm.n2423 C10_P_btm.n2420 1.0005
R33689 C10_P_btm.n2422 C10_P_btm.n2421 1.0005
R33690 C10_P_btm.n2461 C10_P_btm.n2460 1.0005
R33691 C10_P_btm.n2456 C10_P_btm.n2371 1.0005
R33692 C10_P_btm.n2492 C10_P_btm.n2491 1.0005
R33693 C10_P_btm.n2491 C10_P_btm.n2413 1.0005
R33694 C10_P_btm.n2523 C10_P_btm.n2522 1.0005
R33695 C10_P_btm.n2522 C10_P_btm.n2371 1.0005
R33696 C10_P_btm.n2558 C10_P_btm.n2360 1.0005
R33697 C10_P_btm.n2492 C10_P_btm.n2360 1.0005
R33698 C10_P_btm.n2589 C10_P_btm.n2318 1.0005
R33699 C10_P_btm.n2523 C10_P_btm.n2318 1.0005
R33700 C10_P_btm.n2559 C10_P_btm.n2307 1.0005
R33701 C10_P_btm.n2559 C10_P_btm.n2558 1.0005
R33702 C10_P_btm.n2590 C10_P_btm.n2265 1.0005
R33703 C10_P_btm.n2590 C10_P_btm.n2589 1.0005
R33704 C10_P_btm.n2626 C10_P_btm.n2625 1.0005
R33705 C10_P_btm.n2625 C10_P_btm.n2307 1.0005
R33706 C10_P_btm.n2657 C10_P_btm.n2656 1.0005
R33707 C10_P_btm.n2656 C10_P_btm.n2265 1.0005
R33708 C10_P_btm.n2692 C10_P_btm.n2254 1.0005
R33709 C10_P_btm.n2626 C10_P_btm.n2254 1.0005
R33710 C10_P_btm.n2723 C10_P_btm.n2212 1.0005
R33711 C10_P_btm.n2657 C10_P_btm.n2212 1.0005
R33712 C10_P_btm.n2693 C10_P_btm.n2201 1.0005
R33713 C10_P_btm.n2693 C10_P_btm.n2692 1.0005
R33714 C10_P_btm.n2724 C10_P_btm.n2159 1.0005
R33715 C10_P_btm.n2724 C10_P_btm.n2723 1.0005
R33716 C10_P_btm.n2760 C10_P_btm.n2759 1.0005
R33717 C10_P_btm.n2759 C10_P_btm.n2201 1.0005
R33718 C10_P_btm.n2791 C10_P_btm.n2790 1.0005
R33719 C10_P_btm.n2790 C10_P_btm.n2159 1.0005
R33720 C10_P_btm.n2826 C10_P_btm.n2148 1.0005
R33721 C10_P_btm.n2760 C10_P_btm.n2148 1.0005
R33722 C10_P_btm.n2857 C10_P_btm.n2106 1.0005
R33723 C10_P_btm.n2791 C10_P_btm.n2106 1.0005
R33724 C10_P_btm.n2827 C10_P_btm.n2095 1.0005
R33725 C10_P_btm.n2827 C10_P_btm.n2826 1.0005
R33726 C10_P_btm.n2858 C10_P_btm.n2086 1.0005
R33727 C10_P_btm.n2858 C10_P_btm.n2857 1.0005
R33728 C10_P_btm.n2929 C10_P_btm.n2893 1.0005
R33729 C10_P_btm.n2893 C10_P_btm.n2095 1.0005
R33730 C10_P_btm.n2960 C10_P_btm.n2959 1.0005
R33731 C10_P_btm.n2959 C10_P_btm.n2086 1.0005
R33732 C10_P_btm.n2928 C10_P_btm.n2895 1.0005
R33733 C10_P_btm.n2929 C10_P_btm.n2928 1.0005
R33734 C10_P_btm.n3024 C10_P_btm.n2066 1.0005
R33735 C10_P_btm.n2960 C10_P_btm.n2066 1.0005
R33736 C10_P_btm.n3106 C10_P_btm.n2056 1.0005
R33737 C10_P_btm.n2895 C10_P_btm.n2056 1.0005
R33738 C10_P_btm.n3025 C10_P_btm.n537 1.0005
R33739 C10_P_btm.n3025 C10_P_btm.n3024 1.0005
R33740 C10_P_btm.n3026 C10_P_btm.n536 1.0005
R33741 C10_P_btm.n3027 C10_P_btm.n535 1.0005
R33742 C10_P_btm.n3028 C10_P_btm.n534 1.0005
R33743 C10_P_btm.n3029 C10_P_btm.n533 1.0005
R33744 C10_P_btm.n3030 C10_P_btm.n532 1.0005
R33745 C10_P_btm.n3031 C10_P_btm.n531 1.0005
R33746 C10_P_btm.n3032 C10_P_btm.n530 1.0005
R33747 C10_P_btm.n3033 C10_P_btm.n529 1.0005
R33748 C10_P_btm.n3034 C10_P_btm.n528 1.0005
R33749 C10_P_btm.n3035 C10_P_btm.n527 1.0005
R33750 C10_P_btm.n3036 C10_P_btm.n526 1.0005
R33751 C10_P_btm.n3037 C10_P_btm.n525 1.0005
R33752 C10_P_btm.n548 C10_P_btm.n546 1.0005
R33753 C10_P_btm.n549 C10_P_btm.n545 1.0005
R33754 C10_P_btm.n550 C10_P_btm.n544 1.0005
R33755 C10_P_btm.n551 C10_P_btm.n543 1.0005
R33756 C10_P_btm.n552 C10_P_btm.n542 1.0005
R33757 C10_P_btm.n553 C10_P_btm.n541 1.0005
R33758 C10_P_btm.n554 C10_P_btm.n540 1.0005
R33759 C10_P_btm.n555 C10_P_btm.n539 1.0005
R33760 C10_P_btm.n556 C10_P_btm.n538 1.0005
R33761 C10_P_btm.n557 C10_P_btm.n537 1.0005
R33762 C10_P_btm.n558 C10_P_btm.n536 1.0005
R33763 C10_P_btm.n559 C10_P_btm.n535 1.0005
R33764 C10_P_btm.n560 C10_P_btm.n534 1.0005
R33765 C10_P_btm.n561 C10_P_btm.n533 1.0005
R33766 C10_P_btm.n562 C10_P_btm.n532 1.0005
R33767 C10_P_btm.n563 C10_P_btm.n531 1.0005
R33768 C10_P_btm.n564 C10_P_btm.n530 1.0005
R33769 C10_P_btm.n565 C10_P_btm.n529 1.0005
R33770 C10_P_btm.n566 C10_P_btm.n528 1.0005
R33771 C10_P_btm.n567 C10_P_btm.n527 1.0005
R33772 C10_P_btm.n568 C10_P_btm.n526 1.0005
R33773 C10_P_btm.n569 C10_P_btm.n525 1.0005
R33774 C10_P_btm.n570 C10_P_btm.n524 1.0005
R33775 C10_P_btm.n571 C10_P_btm.n523 1.0005
R33776 C10_P_btm.n572 C10_P_btm.n522 1.0005
R33777 C10_P_btm.n573 C10_P_btm.n521 1.0005
R33778 C10_P_btm.n574 C10_P_btm.n520 1.0005
R33779 C10_P_btm.n575 C10_P_btm.n519 1.0005
R33780 C10_P_btm.n576 C10_P_btm.n518 1.0005
R33781 C10_P_btm.n577 C10_P_btm.n517 1.0005
R33782 C10_P_btm.n578 C10_P_btm.n516 1.0005
R33783 C10_P_btm.n579 C10_P_btm.n515 1.0005
R33784 C10_P_btm.n580 C10_P_btm.n514 1.0005
R33785 C10_P_btm.n581 C10_P_btm.n513 1.0005
R33786 C10_P_btm.n582 C10_P_btm.n512 1.0005
R33787 C10_P_btm.n583 C10_P_btm.n511 1.0005
R33788 C10_P_btm.n584 C10_P_btm.n510 1.0005
R33789 C10_P_btm.n585 C10_P_btm.n509 1.0005
R33790 C10_P_btm.n586 C10_P_btm.n508 1.0005
R33791 C10_P_btm.n587 C10_P_btm.n507 1.0005
R33792 C10_P_btm.n588 C10_P_btm.n422 1.0005
R33793 C10_P_btm.n589 C10_P_btm.n421 1.0005
R33794 C10_P_btm.n590 C10_P_btm.n420 1.0005
R33795 C10_P_btm.n591 C10_P_btm.n419 1.0005
R33796 C10_P_btm.n592 C10_P_btm.n418 1.0005
R33797 C10_P_btm.n593 C10_P_btm.n417 1.0005
R33798 C10_P_btm.n594 C10_P_btm.n416 1.0005
R33799 C10_P_btm.n595 C10_P_btm.n415 1.0005
R33800 C10_P_btm.n596 C10_P_btm.n414 1.0005
R33801 C10_P_btm.n597 C10_P_btm.n413 1.0005
R33802 C10_P_btm.n598 C10_P_btm.n412 1.0005
R33803 C10_P_btm.n599 C10_P_btm.n411 1.0005
R33804 C10_P_btm.n600 C10_P_btm.n410 1.0005
R33805 C10_P_btm.n601 C10_P_btm.n409 1.0005
R33806 C10_P_btm.n602 C10_P_btm.n408 1.0005
R33807 C10_P_btm.n603 C10_P_btm.n407 1.0005
R33808 C10_P_btm.n604 C10_P_btm.n406 1.0005
R33809 C10_P_btm.n605 C10_P_btm.n405 1.0005
R33810 C10_P_btm.n606 C10_P_btm.n404 1.0005
R33811 C10_P_btm.n607 C10_P_btm.n403 1.0005
R33812 C10_P_btm.n608 C10_P_btm.n402 1.0005
R33813 C10_P_btm.n1866 C10_P_btm.n399 1.0005
R33814 C10_P_btm.n1866 C10_P_btm.n1865 1.0005
R33815 C10_P_btm.n733 C10_P_btm.n608 1.0005
R33816 C10_P_btm.n732 C10_P_btm.n607 1.0005
R33817 C10_P_btm.n731 C10_P_btm.n606 1.0005
R33818 C10_P_btm.n730 C10_P_btm.n605 1.0005
R33819 C10_P_btm.n729 C10_P_btm.n604 1.0005
R33820 C10_P_btm.n728 C10_P_btm.n603 1.0005
R33821 C10_P_btm.n727 C10_P_btm.n602 1.0005
R33822 C10_P_btm.n726 C10_P_btm.n601 1.0005
R33823 C10_P_btm.n725 C10_P_btm.n600 1.0005
R33824 C10_P_btm.n724 C10_P_btm.n599 1.0005
R33825 C10_P_btm.n723 C10_P_btm.n598 1.0005
R33826 C10_P_btm.n722 C10_P_btm.n597 1.0005
R33827 C10_P_btm.n721 C10_P_btm.n596 1.0005
R33828 C10_P_btm.n720 C10_P_btm.n595 1.0005
R33829 C10_P_btm.n719 C10_P_btm.n594 1.0005
R33830 C10_P_btm.n718 C10_P_btm.n593 1.0005
R33831 C10_P_btm.n717 C10_P_btm.n592 1.0005
R33832 C10_P_btm.n716 C10_P_btm.n591 1.0005
R33833 C10_P_btm.n715 C10_P_btm.n590 1.0005
R33834 C10_P_btm.n714 C10_P_btm.n589 1.0005
R33835 C10_P_btm.n713 C10_P_btm.n588 1.0005
R33836 C10_P_btm.n712 C10_P_btm.n587 1.0005
R33837 C10_P_btm.n711 C10_P_btm.n586 1.0005
R33838 C10_P_btm.n710 C10_P_btm.n585 1.0005
R33839 C10_P_btm.n709 C10_P_btm.n584 1.0005
R33840 C10_P_btm.n708 C10_P_btm.n583 1.0005
R33841 C10_P_btm.n707 C10_P_btm.n582 1.0005
R33842 C10_P_btm.n706 C10_P_btm.n581 1.0005
R33843 C10_P_btm.n705 C10_P_btm.n580 1.0005
R33844 C10_P_btm.n704 C10_P_btm.n579 1.0005
R33845 C10_P_btm.n703 C10_P_btm.n578 1.0005
R33846 C10_P_btm.n702 C10_P_btm.n577 1.0005
R33847 C10_P_btm.n701 C10_P_btm.n576 1.0005
R33848 C10_P_btm.n700 C10_P_btm.n575 1.0005
R33849 C10_P_btm.n699 C10_P_btm.n574 1.0005
R33850 C10_P_btm.n698 C10_P_btm.n573 1.0005
R33851 C10_P_btm.n697 C10_P_btm.n572 1.0005
R33852 C10_P_btm.n696 C10_P_btm.n571 1.0005
R33853 C10_P_btm.n695 C10_P_btm.n570 1.0005
R33854 C10_P_btm.n694 C10_P_btm.n569 1.0005
R33855 C10_P_btm.n693 C10_P_btm.n568 1.0005
R33856 C10_P_btm.n692 C10_P_btm.n567 1.0005
R33857 C10_P_btm.n691 C10_P_btm.n566 1.0005
R33858 C10_P_btm.n690 C10_P_btm.n565 1.0005
R33859 C10_P_btm.n689 C10_P_btm.n564 1.0005
R33860 C10_P_btm.n688 C10_P_btm.n563 1.0005
R33861 C10_P_btm.n687 C10_P_btm.n562 1.0005
R33862 C10_P_btm.n686 C10_P_btm.n561 1.0005
R33863 C10_P_btm.n685 C10_P_btm.n560 1.0005
R33864 C10_P_btm.n684 C10_P_btm.n559 1.0005
R33865 C10_P_btm.n683 C10_P_btm.n558 1.0005
R33866 C10_P_btm.n682 C10_P_btm.n557 1.0005
R33867 C10_P_btm.n681 C10_P_btm.n556 1.0005
R33868 C10_P_btm.n680 C10_P_btm.n555 1.0005
R33869 C10_P_btm.n679 C10_P_btm.n554 1.0005
R33870 C10_P_btm.n678 C10_P_btm.n553 1.0005
R33871 C10_P_btm.n677 C10_P_btm.n552 1.0005
R33872 C10_P_btm.n676 C10_P_btm.n551 1.0005
R33873 C10_P_btm.n675 C10_P_btm.n550 1.0005
R33874 C10_P_btm.n674 C10_P_btm.n549 1.0005
R33875 C10_P_btm.n916 C10_P_btm.n548 1.0005
R33876 C10_P_btm.n917 C10_P_btm.n916 1.0005
R33877 C10_P_btm.n674 C10_P_btm.n671 1.0005
R33878 C10_P_btm.n675 C10_P_btm.n670 1.0005
R33879 C10_P_btm.n676 C10_P_btm.n669 1.0005
R33880 C10_P_btm.n677 C10_P_btm.n668 1.0005
R33881 C10_P_btm.n678 C10_P_btm.n667 1.0005
R33882 C10_P_btm.n679 C10_P_btm.n666 1.0005
R33883 C10_P_btm.n680 C10_P_btm.n665 1.0005
R33884 C10_P_btm.n681 C10_P_btm.n664 1.0005
R33885 C10_P_btm.n682 C10_P_btm.n663 1.0005
R33886 C10_P_btm.n683 C10_P_btm.n662 1.0005
R33887 C10_P_btm.n684 C10_P_btm.n661 1.0005
R33888 C10_P_btm.n685 C10_P_btm.n660 1.0005
R33889 C10_P_btm.n686 C10_P_btm.n659 1.0005
R33890 C10_P_btm.n687 C10_P_btm.n658 1.0005
R33891 C10_P_btm.n688 C10_P_btm.n657 1.0005
R33892 C10_P_btm.n689 C10_P_btm.n656 1.0005
R33893 C10_P_btm.n690 C10_P_btm.n655 1.0005
R33894 C10_P_btm.n691 C10_P_btm.n654 1.0005
R33895 C10_P_btm.n692 C10_P_btm.n653 1.0005
R33896 C10_P_btm.n693 C10_P_btm.n652 1.0005
R33897 C10_P_btm.n694 C10_P_btm.n651 1.0005
R33898 C10_P_btm.n695 C10_P_btm.n650 1.0005
R33899 C10_P_btm.n696 C10_P_btm.n649 1.0005
R33900 C10_P_btm.n697 C10_P_btm.n648 1.0005
R33901 C10_P_btm.n698 C10_P_btm.n647 1.0005
R33902 C10_P_btm.n699 C10_P_btm.n646 1.0005
R33903 C10_P_btm.n700 C10_P_btm.n645 1.0005
R33904 C10_P_btm.n701 C10_P_btm.n644 1.0005
R33905 C10_P_btm.n702 C10_P_btm.n643 1.0005
R33906 C10_P_btm.n703 C10_P_btm.n642 1.0005
R33907 C10_P_btm.n704 C10_P_btm.n641 1.0005
R33908 C10_P_btm.n705 C10_P_btm.n640 1.0005
R33909 C10_P_btm.n706 C10_P_btm.n639 1.0005
R33910 C10_P_btm.n707 C10_P_btm.n638 1.0005
R33911 C10_P_btm.n708 C10_P_btm.n637 1.0005
R33912 C10_P_btm.n709 C10_P_btm.n636 1.0005
R33913 C10_P_btm.n710 C10_P_btm.n635 1.0005
R33914 C10_P_btm.n711 C10_P_btm.n634 1.0005
R33915 C10_P_btm.n712 C10_P_btm.n633 1.0005
R33916 C10_P_btm.n713 C10_P_btm.n632 1.0005
R33917 C10_P_btm.n714 C10_P_btm.n631 1.0005
R33918 C10_P_btm.n715 C10_P_btm.n630 1.0005
R33919 C10_P_btm.n716 C10_P_btm.n629 1.0005
R33920 C10_P_btm.n717 C10_P_btm.n628 1.0005
R33921 C10_P_btm.n718 C10_P_btm.n627 1.0005
R33922 C10_P_btm.n719 C10_P_btm.n626 1.0005
R33923 C10_P_btm.n720 C10_P_btm.n625 1.0005
R33924 C10_P_btm.n721 C10_P_btm.n624 1.0005
R33925 C10_P_btm.n722 C10_P_btm.n623 1.0005
R33926 C10_P_btm.n723 C10_P_btm.n622 1.0005
R33927 C10_P_btm.n724 C10_P_btm.n621 1.0005
R33928 C10_P_btm.n725 C10_P_btm.n620 1.0005
R33929 C10_P_btm.n726 C10_P_btm.n619 1.0005
R33930 C10_P_btm.n727 C10_P_btm.n618 1.0005
R33931 C10_P_btm.n728 C10_P_btm.n617 1.0005
R33932 C10_P_btm.n729 C10_P_btm.n616 1.0005
R33933 C10_P_btm.n730 C10_P_btm.n615 1.0005
R33934 C10_P_btm.n731 C10_P_btm.n614 1.0005
R33935 C10_P_btm.n732 C10_P_btm.n613 1.0005
R33936 C10_P_btm.n733 C10_P_btm.n612 1.0005
R33937 C10_P_btm.n1865 C10_P_btm.n609 1.0005
R33938 C10_P_btm.n1481 C10_P_btm.n609 1.0005
R33939 C10_P_btm.n979 C10_P_btm.n612 1.0005
R33940 C10_P_btm.n978 C10_P_btm.n613 1.0005
R33941 C10_P_btm.n977 C10_P_btm.n614 1.0005
R33942 C10_P_btm.n976 C10_P_btm.n615 1.0005
R33943 C10_P_btm.n975 C10_P_btm.n616 1.0005
R33944 C10_P_btm.n974 C10_P_btm.n617 1.0005
R33945 C10_P_btm.n973 C10_P_btm.n618 1.0005
R33946 C10_P_btm.n972 C10_P_btm.n619 1.0005
R33947 C10_P_btm.n971 C10_P_btm.n620 1.0005
R33948 C10_P_btm.n970 C10_P_btm.n621 1.0005
R33949 C10_P_btm.n969 C10_P_btm.n622 1.0005
R33950 C10_P_btm.n968 C10_P_btm.n623 1.0005
R33951 C10_P_btm.n967 C10_P_btm.n624 1.0005
R33952 C10_P_btm.n966 C10_P_btm.n625 1.0005
R33953 C10_P_btm.n965 C10_P_btm.n626 1.0005
R33954 C10_P_btm.n964 C10_P_btm.n627 1.0005
R33955 C10_P_btm.n963 C10_P_btm.n628 1.0005
R33956 C10_P_btm.n962 C10_P_btm.n629 1.0005
R33957 C10_P_btm.n961 C10_P_btm.n630 1.0005
R33958 C10_P_btm.n960 C10_P_btm.n631 1.0005
R33959 C10_P_btm.n959 C10_P_btm.n632 1.0005
R33960 C10_P_btm.n958 C10_P_btm.n633 1.0005
R33961 C10_P_btm.n957 C10_P_btm.n634 1.0005
R33962 C10_P_btm.n956 C10_P_btm.n635 1.0005
R33963 C10_P_btm.n955 C10_P_btm.n636 1.0005
R33964 C10_P_btm.n954 C10_P_btm.n637 1.0005
R33965 C10_P_btm.n953 C10_P_btm.n638 1.0005
R33966 C10_P_btm.n952 C10_P_btm.n639 1.0005
R33967 C10_P_btm.n951 C10_P_btm.n640 1.0005
R33968 C10_P_btm.n950 C10_P_btm.n641 1.0005
R33969 C10_P_btm.n949 C10_P_btm.n642 1.0005
R33970 C10_P_btm.n948 C10_P_btm.n643 1.0005
R33971 C10_P_btm.n947 C10_P_btm.n644 1.0005
R33972 C10_P_btm.n946 C10_P_btm.n645 1.0005
R33973 C10_P_btm.n945 C10_P_btm.n646 1.0005
R33974 C10_P_btm.n944 C10_P_btm.n647 1.0005
R33975 C10_P_btm.n943 C10_P_btm.n648 1.0005
R33976 C10_P_btm.n942 C10_P_btm.n649 1.0005
R33977 C10_P_btm.n941 C10_P_btm.n650 1.0005
R33978 C10_P_btm.n940 C10_P_btm.n651 1.0005
R33979 C10_P_btm.n939 C10_P_btm.n652 1.0005
R33980 C10_P_btm.n938 C10_P_btm.n653 1.0005
R33981 C10_P_btm.n937 C10_P_btm.n654 1.0005
R33982 C10_P_btm.n936 C10_P_btm.n655 1.0005
R33983 C10_P_btm.n935 C10_P_btm.n656 1.0005
R33984 C10_P_btm.n934 C10_P_btm.n657 1.0005
R33985 C10_P_btm.n933 C10_P_btm.n658 1.0005
R33986 C10_P_btm.n932 C10_P_btm.n659 1.0005
R33987 C10_P_btm.n931 C10_P_btm.n660 1.0005
R33988 C10_P_btm.n930 C10_P_btm.n661 1.0005
R33989 C10_P_btm.n929 C10_P_btm.n662 1.0005
R33990 C10_P_btm.n928 C10_P_btm.n663 1.0005
R33991 C10_P_btm.n927 C10_P_btm.n664 1.0005
R33992 C10_P_btm.n926 C10_P_btm.n665 1.0005
R33993 C10_P_btm.n925 C10_P_btm.n666 1.0005
R33994 C10_P_btm.n924 C10_P_btm.n667 1.0005
R33995 C10_P_btm.n923 C10_P_btm.n668 1.0005
R33996 C10_P_btm.n922 C10_P_btm.n669 1.0005
R33997 C10_P_btm.n921 C10_P_btm.n670 1.0005
R33998 C10_P_btm.n920 C10_P_btm.n671 1.0005
R33999 C10_P_btm.n919 C10_P_btm.n917 1.0005
R34000 C10_P_btm.n1286 C10_P_btm.n919 1.0005
R34001 C10_P_btm.n1044 C10_P_btm.n920 1.0005
R34002 C10_P_btm.n1045 C10_P_btm.n921 1.0005
R34003 C10_P_btm.n1046 C10_P_btm.n922 1.0005
R34004 C10_P_btm.n1047 C10_P_btm.n923 1.0005
R34005 C10_P_btm.n1048 C10_P_btm.n924 1.0005
R34006 C10_P_btm.n1049 C10_P_btm.n925 1.0005
R34007 C10_P_btm.n1050 C10_P_btm.n926 1.0005
R34008 C10_P_btm.n1051 C10_P_btm.n927 1.0005
R34009 C10_P_btm.n1052 C10_P_btm.n928 1.0005
R34010 C10_P_btm.n1053 C10_P_btm.n929 1.0005
R34011 C10_P_btm.n1054 C10_P_btm.n930 1.0005
R34012 C10_P_btm.n1055 C10_P_btm.n931 1.0005
R34013 C10_P_btm.n1056 C10_P_btm.n932 1.0005
R34014 C10_P_btm.n1057 C10_P_btm.n933 1.0005
R34015 C10_P_btm.n1058 C10_P_btm.n934 1.0005
R34016 C10_P_btm.n1059 C10_P_btm.n935 1.0005
R34017 C10_P_btm.n1060 C10_P_btm.n936 1.0005
R34018 C10_P_btm.n1061 C10_P_btm.n937 1.0005
R34019 C10_P_btm.n1062 C10_P_btm.n938 1.0005
R34020 C10_P_btm.n1063 C10_P_btm.n939 1.0005
R34021 C10_P_btm.n1064 C10_P_btm.n940 1.0005
R34022 C10_P_btm.n1065 C10_P_btm.n941 1.0005
R34023 C10_P_btm.n1066 C10_P_btm.n942 1.0005
R34024 C10_P_btm.n1067 C10_P_btm.n943 1.0005
R34025 C10_P_btm.n1068 C10_P_btm.n944 1.0005
R34026 C10_P_btm.n1069 C10_P_btm.n945 1.0005
R34027 C10_P_btm.n1070 C10_P_btm.n946 1.0005
R34028 C10_P_btm.n1071 C10_P_btm.n947 1.0005
R34029 C10_P_btm.n1072 C10_P_btm.n948 1.0005
R34030 C10_P_btm.n1073 C10_P_btm.n949 1.0005
R34031 C10_P_btm.n1074 C10_P_btm.n950 1.0005
R34032 C10_P_btm.n1075 C10_P_btm.n951 1.0005
R34033 C10_P_btm.n1076 C10_P_btm.n952 1.0005
R34034 C10_P_btm.n1077 C10_P_btm.n953 1.0005
R34035 C10_P_btm.n1078 C10_P_btm.n954 1.0005
R34036 C10_P_btm.n1079 C10_P_btm.n955 1.0005
R34037 C10_P_btm.n1080 C10_P_btm.n956 1.0005
R34038 C10_P_btm.n1081 C10_P_btm.n957 1.0005
R34039 C10_P_btm.n1082 C10_P_btm.n958 1.0005
R34040 C10_P_btm.n1083 C10_P_btm.n959 1.0005
R34041 C10_P_btm.n1084 C10_P_btm.n960 1.0005
R34042 C10_P_btm.n1085 C10_P_btm.n961 1.0005
R34043 C10_P_btm.n1086 C10_P_btm.n962 1.0005
R34044 C10_P_btm.n1087 C10_P_btm.n963 1.0005
R34045 C10_P_btm.n1088 C10_P_btm.n964 1.0005
R34046 C10_P_btm.n1089 C10_P_btm.n965 1.0005
R34047 C10_P_btm.n1090 C10_P_btm.n966 1.0005
R34048 C10_P_btm.n1091 C10_P_btm.n967 1.0005
R34049 C10_P_btm.n1092 C10_P_btm.n968 1.0005
R34050 C10_P_btm.n1093 C10_P_btm.n969 1.0005
R34051 C10_P_btm.n1094 C10_P_btm.n970 1.0005
R34052 C10_P_btm.n1095 C10_P_btm.n971 1.0005
R34053 C10_P_btm.n1096 C10_P_btm.n972 1.0005
R34054 C10_P_btm.n1097 C10_P_btm.n973 1.0005
R34055 C10_P_btm.n1098 C10_P_btm.n974 1.0005
R34056 C10_P_btm.n1099 C10_P_btm.n975 1.0005
R34057 C10_P_btm.n1100 C10_P_btm.n976 1.0005
R34058 C10_P_btm.n1101 C10_P_btm.n977 1.0005
R34059 C10_P_btm.n1102 C10_P_btm.n978 1.0005
R34060 C10_P_btm.n1103 C10_P_btm.n979 1.0005
R34061 C10_P_btm.n1481 C10_P_btm.n1480 1.0005
R34062 C10_P_btm.n1480 C10_P_btm.n980 1.0005
R34063 C10_P_btm.n1103 C10_P_btm.n982 1.0005
R34064 C10_P_btm.n1102 C10_P_btm.n983 1.0005
R34065 C10_P_btm.n1101 C10_P_btm.n984 1.0005
R34066 C10_P_btm.n1100 C10_P_btm.n985 1.0005
R34067 C10_P_btm.n1099 C10_P_btm.n986 1.0005
R34068 C10_P_btm.n1098 C10_P_btm.n987 1.0005
R34069 C10_P_btm.n1097 C10_P_btm.n988 1.0005
R34070 C10_P_btm.n1096 C10_P_btm.n989 1.0005
R34071 C10_P_btm.n1095 C10_P_btm.n990 1.0005
R34072 C10_P_btm.n1094 C10_P_btm.n991 1.0005
R34073 C10_P_btm.n1093 C10_P_btm.n992 1.0005
R34074 C10_P_btm.n1092 C10_P_btm.n993 1.0005
R34075 C10_P_btm.n1091 C10_P_btm.n994 1.0005
R34076 C10_P_btm.n1090 C10_P_btm.n995 1.0005
R34077 C10_P_btm.n1089 C10_P_btm.n996 1.0005
R34078 C10_P_btm.n1088 C10_P_btm.n997 1.0005
R34079 C10_P_btm.n1087 C10_P_btm.n998 1.0005
R34080 C10_P_btm.n1086 C10_P_btm.n999 1.0005
R34081 C10_P_btm.n1085 C10_P_btm.n1000 1.0005
R34082 C10_P_btm.n1084 C10_P_btm.n1001 1.0005
R34083 C10_P_btm.n1083 C10_P_btm.n1002 1.0005
R34084 C10_P_btm.n1082 C10_P_btm.n1003 1.0005
R34085 C10_P_btm.n1081 C10_P_btm.n1004 1.0005
R34086 C10_P_btm.n1080 C10_P_btm.n1005 1.0005
R34087 C10_P_btm.n1079 C10_P_btm.n1006 1.0005
R34088 C10_P_btm.n1078 C10_P_btm.n1007 1.0005
R34089 C10_P_btm.n1077 C10_P_btm.n1008 1.0005
R34090 C10_P_btm.n1076 C10_P_btm.n1009 1.0005
R34091 C10_P_btm.n1075 C10_P_btm.n1010 1.0005
R34092 C10_P_btm.n1074 C10_P_btm.n1011 1.0005
R34093 C10_P_btm.n1073 C10_P_btm.n1012 1.0005
R34094 C10_P_btm.n1072 C10_P_btm.n1013 1.0005
R34095 C10_P_btm.n1071 C10_P_btm.n1014 1.0005
R34096 C10_P_btm.n1070 C10_P_btm.n1015 1.0005
R34097 C10_P_btm.n1069 C10_P_btm.n1016 1.0005
R34098 C10_P_btm.n1068 C10_P_btm.n1017 1.0005
R34099 C10_P_btm.n1067 C10_P_btm.n1018 1.0005
R34100 C10_P_btm.n1066 C10_P_btm.n1019 1.0005
R34101 C10_P_btm.n1065 C10_P_btm.n1020 1.0005
R34102 C10_P_btm.n1064 C10_P_btm.n1021 1.0005
R34103 C10_P_btm.n1063 C10_P_btm.n1022 1.0005
R34104 C10_P_btm.n1062 C10_P_btm.n1023 1.0005
R34105 C10_P_btm.n1061 C10_P_btm.n1024 1.0005
R34106 C10_P_btm.n1060 C10_P_btm.n1025 1.0005
R34107 C10_P_btm.n1059 C10_P_btm.n1026 1.0005
R34108 C10_P_btm.n1058 C10_P_btm.n1027 1.0005
R34109 C10_P_btm.n1057 C10_P_btm.n1028 1.0005
R34110 C10_P_btm.n1056 C10_P_btm.n1029 1.0005
R34111 C10_P_btm.n1055 C10_P_btm.n1030 1.0005
R34112 C10_P_btm.n1054 C10_P_btm.n1031 1.0005
R34113 C10_P_btm.n1053 C10_P_btm.n1032 1.0005
R34114 C10_P_btm.n1052 C10_P_btm.n1033 1.0005
R34115 C10_P_btm.n1051 C10_P_btm.n1034 1.0005
R34116 C10_P_btm.n1050 C10_P_btm.n1035 1.0005
R34117 C10_P_btm.n1049 C10_P_btm.n1036 1.0005
R34118 C10_P_btm.n1048 C10_P_btm.n1037 1.0005
R34119 C10_P_btm.n1047 C10_P_btm.n1038 1.0005
R34120 C10_P_btm.n1046 C10_P_btm.n1039 1.0005
R34121 C10_P_btm.n1045 C10_P_btm.n1040 1.0005
R34122 C10_P_btm.n1044 C10_P_btm.n1041 1.0005
R34123 C10_P_btm.n1287 C10_P_btm.n1286 1.0005
R34124 C10_P_btm.n1476 C10_P_btm.n611 1.0005
R34125 C10_P_btm.n1670 C10_P_btm.n918 1.0005
R34126 C10_P_btm.n1671 C10_P_btm.n1670 1.0005
R34127 C10_P_btm.n1860 C10_P_btm.n611 1.0005
R34128 C10_P_btm.n1861 C10_P_btm.n1860 1.0005
R34129 C10_P_btm.n1671 C10_P_btm.n547 1.0005
R34130 C10_P_btm.n2055 C10_P_btm.n547 1.0005
R34131 C10_P_btm.n1861 C10_P_btm.n401 1.0005
R34132 C10_P_btm.n3296 C10_P_btm.n401 1.0005
R34133 C10_P_btm.n3107 C10_P_btm.n2055 1.0005
R34134 C10_P_btm.n3107 C10_P_btm.n3106 1.0005
R34135 C10_P_btm.n3297 C10_P_btm.n3296 1.0005
R34136 C10_P_btm.n3297 C10_P_btm.n348 1.0005
R34137 C10_P_btm.n3332 C10_P_btm.n390 1.0005
R34138 C10_P_btm.n3333 C10_P_btm.n3332 1.0005
R34139 C10_P_btm.n3363 C10_P_btm.n348 1.0005
R34140 C10_P_btm.n3364 C10_P_btm.n3363 1.0005
R34141 C10_P_btm.n3333 C10_P_btm.n337 1.0005
R34142 C10_P_btm.n3399 C10_P_btm.n337 1.0005
R34143 C10_P_btm.n3364 C10_P_btm.n295 1.0005
R34144 C10_P_btm.n3430 C10_P_btm.n295 1.0005
R34145 C10_P_btm.n3400 C10_P_btm.n3399 1.0005
R34146 C10_P_btm.n3400 C10_P_btm.n284 1.0005
R34147 C10_P_btm.n3431 C10_P_btm.n3430 1.0005
R34148 C10_P_btm.n3431 C10_P_btm.n242 1.0005
R34149 C10_P_btm.n3466 C10_P_btm.n284 1.0005
R34150 C10_P_btm.n3467 C10_P_btm.n3466 1.0005
R34151 C10_P_btm.n3497 C10_P_btm.n242 1.0005
R34152 C10_P_btm.n3498 C10_P_btm.n3497 1.0005
R34153 C10_P_btm.n3467 C10_P_btm.n231 1.0005
R34154 C10_P_btm.n3533 C10_P_btm.n231 1.0005
R34155 C10_P_btm.n3498 C10_P_btm.n189 1.0005
R34156 C10_P_btm.n3564 C10_P_btm.n189 1.0005
R34157 C10_P_btm.n3534 C10_P_btm.n3533 1.0005
R34158 C10_P_btm.n3534 C10_P_btm.n178 1.0005
R34159 C10_P_btm.n3565 C10_P_btm.n3564 1.0005
R34160 C10_P_btm.n3565 C10_P_btm.n136 1.0005
R34161 C10_P_btm.n3600 C10_P_btm.n178 1.0005
R34162 C10_P_btm.n3601 C10_P_btm.n3600 1.0005
R34163 C10_P_btm.n3631 C10_P_btm.n136 1.0005
R34164 C10_P_btm.n3632 C10_P_btm.n3631 1.0005
R34165 C10_P_btm.n3601 C10_P_btm.n125 1.0005
R34166 C10_P_btm.n3667 C10_P_btm.n125 1.0005
R34167 C10_P_btm.n3632 C10_P_btm.n83 1.0005
R34168 C10_P_btm.n3698 C10_P_btm.n83 1.0005
R34169 C10_P_btm.n3668 C10_P_btm.n3667 1.0005
R34170 C10_P_btm.n3668 C10_P_btm.n72 1.0005
R34171 C10_P_btm.n3699 C10_P_btm.n3698 1.0005
R34172 C10_P_btm.n3699 C10_P_btm.n63 1.0005
R34173 C10_P_btm.n3734 C10_P_btm.n72 1.0005
R34174 C10_P_btm.n3770 C10_P_btm.n3734 1.0005
R34175 C10_P_btm.n3800 C10_P_btm.n63 1.0005
R34176 C10_P_btm.n3801 C10_P_btm.n3800 1.0005
R34177 C10_P_btm.n3770 C10_P_btm.n3769 1.0005
R34178 C10_P_btm.n3769 C10_P_btm.n3736 1.0005
R34179 C10_P_btm.n3801 C10_P_btm.n43 1.0005
R34180 C10_P_btm.n3865 C10_P_btm.n43 1.0005
R34181 C10_P_btm.n3736 C10_P_btm.n33 1.0005
R34182 C10_P_btm.n3896 C10_P_btm.n33 1.0005
R34183 C10_P_btm.n3866 C10_P_btm.n3865 1.0005
R34184 C10_P_btm.n3897 C10_P_btm.n3896 1.0005
R34185 C10_P_btm.n4 C10_P_btm.n2 0.71925
R34186 C10_P_btm.n8 C10_P_btm.n6 0.71925
R34187 C10_P_btm.n12 C10_P_btm.n10 0.71925
R34188 C10_P_btm.n6 C10_P_btm.n4 0.688
R34189 C10_P_btm.n10 C10_P_btm.n8 0.688
R34190 C10_P_btm.n506 C10_P_btm.n505 0.679419
R34191 C10_P_btm.n2459 C10_P_btm.n2457 0.679419
R34192 C10_P_btm.n2431 C10_P_btm.n2430 0.679419
R34193 C10_P_btm.n2490 C10_P_btm.n2489 0.679419
R34194 C10_P_btm.n2463 C10_P_btm.n2462 0.679419
R34195 C10_P_btm.n2521 C10_P_btm.n2520 0.679419
R34196 C10_P_btm.n2494 C10_P_btm.n2493 0.679419
R34197 C10_P_btm.n2380 C10_P_btm.n2379 0.679419
R34198 C10_P_btm.n2526 C10_P_btm.n2524 0.679419
R34199 C10_P_btm.n2530 C10_P_btm.n2529 0.679419
R34200 C10_P_btm.n2557 C10_P_btm.n2556 0.679419
R34201 C10_P_btm.n2561 C10_P_btm.n2560 0.679419
R34202 C10_P_btm.n2588 C10_P_btm.n2587 0.679419
R34203 C10_P_btm.n2593 C10_P_btm.n2591 0.679419
R34204 C10_P_btm.n2327 C10_P_btm.n2326 0.679419
R34205 C10_P_btm.n2624 C10_P_btm.n2623 0.679419
R34206 C10_P_btm.n2597 C10_P_btm.n2596 0.679419
R34207 C10_P_btm.n2655 C10_P_btm.n2654 0.679419
R34208 C10_P_btm.n2628 C10_P_btm.n2627 0.679419
R34209 C10_P_btm.n2274 C10_P_btm.n2273 0.679419
R34210 C10_P_btm.n2660 C10_P_btm.n2658 0.679419
R34211 C10_P_btm.n2664 C10_P_btm.n2663 0.679419
R34212 C10_P_btm.n2691 C10_P_btm.n2690 0.679419
R34213 C10_P_btm.n2695 C10_P_btm.n2694 0.679419
R34214 C10_P_btm.n2722 C10_P_btm.n2721 0.679419
R34215 C10_P_btm.n2727 C10_P_btm.n2725 0.679419
R34216 C10_P_btm.n2221 C10_P_btm.n2220 0.679419
R34217 C10_P_btm.n2758 C10_P_btm.n2757 0.679419
R34218 C10_P_btm.n2731 C10_P_btm.n2730 0.679419
R34219 C10_P_btm.n2789 C10_P_btm.n2788 0.679419
R34220 C10_P_btm.n2762 C10_P_btm.n2761 0.679419
R34221 C10_P_btm.n2168 C10_P_btm.n2167 0.679419
R34222 C10_P_btm.n2794 C10_P_btm.n2792 0.679419
R34223 C10_P_btm.n2798 C10_P_btm.n2797 0.679419
R34224 C10_P_btm.n2825 C10_P_btm.n2824 0.679419
R34225 C10_P_btm.n2829 C10_P_btm.n2828 0.679419
R34226 C10_P_btm.n2856 C10_P_btm.n2855 0.679419
R34227 C10_P_btm.n2861 C10_P_btm.n2859 0.679419
R34228 C10_P_btm.n2115 C10_P_btm.n2114 0.679419
R34229 C10_P_btm.n2892 C10_P_btm.n2891 0.679419
R34230 C10_P_btm.n2865 C10_P_btm.n2864 0.679419
R34231 C10_P_btm.n2958 C10_P_btm.n2957 0.679419
R34232 C10_P_btm.n2931 C10_P_btm.n2930 0.679419
R34233 C10_P_btm.n2927 C10_P_btm.n2926 0.679419
R34234 C10_P_btm.n2963 C10_P_btm.n2961 0.679419
R34235 C10_P_btm.n2967 C10_P_btm.n2966 0.679419
R34236 C10_P_btm.n2894 C10_P_btm.n2076 0.679419
R34237 C10_P_btm.n2996 C10_P_btm.n2995 0.679419
R34238 C10_P_btm.n3023 C10_P_btm.n3022 0.679419
R34239 C10_P_btm.n3039 C10_P_btm.n3038 0.679419
R34240 C10_P_btm.n3105 C10_P_btm.n3104 0.679419
R34241 C10_P_btm.n1289 C10_P_btm.n1288 0.679419
R34242 C10_P_btm.n1475 C10_P_btm.n1474 0.679419
R34243 C10_P_btm.n1479 C10_P_btm.n1477 0.679419
R34244 C10_P_btm.n1043 C10_P_btm.n1042 0.679419
R34245 C10_P_btm.n1669 C10_P_btm.n1668 0.679419
R34246 C10_P_btm.n1483 C10_P_btm.n1482 0.679419
R34247 C10_P_btm.n1859 C10_P_btm.n1858 0.679419
R34248 C10_P_btm.n1673 C10_P_btm.n1672 0.679419
R34249 C10_P_btm.n673 C10_P_btm.n672 0.679419
R34250 C10_P_btm.n1864 C10_P_btm.n1862 0.679419
R34251 C10_P_btm.n1868 C10_P_btm.n1867 0.679419
R34252 C10_P_btm.n2054 C10_P_btm.n2053 0.679419
R34253 C10_P_btm.n3109 C10_P_btm.n3108 0.679419
R34254 C10_P_btm.n3295 C10_P_btm.n3294 0.679419
R34255 C10_P_btm.n3300 C10_P_btm.n3298 0.679419
R34256 C10_P_btm.n3331 C10_P_btm.n3330 0.679419
R34257 C10_P_btm.n3304 C10_P_btm.n3303 0.679419
R34258 C10_P_btm.n3362 C10_P_btm.n3361 0.679419
R34259 C10_P_btm.n3335 C10_P_btm.n3334 0.679419
R34260 C10_P_btm.n357 C10_P_btm.n356 0.679419
R34261 C10_P_btm.n3367 C10_P_btm.n3365 0.679419
R34262 C10_P_btm.n3371 C10_P_btm.n3370 0.679419
R34263 C10_P_btm.n3398 C10_P_btm.n3397 0.679419
R34264 C10_P_btm.n3402 C10_P_btm.n3401 0.679419
R34265 C10_P_btm.n3429 C10_P_btm.n3428 0.679419
R34266 C10_P_btm.n3434 C10_P_btm.n3432 0.679419
R34267 C10_P_btm.n304 C10_P_btm.n303 0.679419
R34268 C10_P_btm.n3465 C10_P_btm.n3464 0.679419
R34269 C10_P_btm.n3438 C10_P_btm.n3437 0.679419
R34270 C10_P_btm.n3496 C10_P_btm.n3495 0.679419
R34271 C10_P_btm.n3469 C10_P_btm.n3468 0.679419
R34272 C10_P_btm.n251 C10_P_btm.n250 0.679419
R34273 C10_P_btm.n3501 C10_P_btm.n3499 0.679419
R34274 C10_P_btm.n3505 C10_P_btm.n3504 0.679419
R34275 C10_P_btm.n3532 C10_P_btm.n3531 0.679419
R34276 C10_P_btm.n3536 C10_P_btm.n3535 0.679419
R34277 C10_P_btm.n3563 C10_P_btm.n3562 0.679419
R34278 C10_P_btm.n3568 C10_P_btm.n3566 0.679419
R34279 C10_P_btm.n198 C10_P_btm.n197 0.679419
R34280 C10_P_btm.n3599 C10_P_btm.n3598 0.679419
R34281 C10_P_btm.n3572 C10_P_btm.n3571 0.679419
R34282 C10_P_btm.n3630 C10_P_btm.n3629 0.679419
R34283 C10_P_btm.n3603 C10_P_btm.n3602 0.679419
R34284 C10_P_btm.n145 C10_P_btm.n144 0.679419
R34285 C10_P_btm.n3635 C10_P_btm.n3633 0.679419
R34286 C10_P_btm.n3639 C10_P_btm.n3638 0.679419
R34287 C10_P_btm.n3666 C10_P_btm.n3665 0.679419
R34288 C10_P_btm.n3670 C10_P_btm.n3669 0.679419
R34289 C10_P_btm.n3697 C10_P_btm.n3696 0.679419
R34290 C10_P_btm.n3702 C10_P_btm.n3700 0.679419
R34291 C10_P_btm.n92 C10_P_btm.n91 0.679419
R34292 C10_P_btm.n3733 C10_P_btm.n3732 0.679419
R34293 C10_P_btm.n3706 C10_P_btm.n3705 0.679419
R34294 C10_P_btm.n3799 C10_P_btm.n3798 0.679419
R34295 C10_P_btm.n3772 C10_P_btm.n3771 0.679419
R34296 C10_P_btm.n3768 C10_P_btm.n3767 0.679419
R34297 C10_P_btm.n3804 C10_P_btm.n3802 0.679419
R34298 C10_P_btm.n3808 C10_P_btm.n3807 0.679419
R34299 C10_P_btm.n3735 C10_P_btm.n53 0.679419
R34300 C10_P_btm.n3837 C10_P_btm.n3836 0.679419
R34301 C10_P_btm.n3864 C10_P_btm.n3863 0.679419
R34302 C10_P_btm.n3868 C10_P_btm.n3867 0.679419
R34303 C10_P_btm.n3895 C10_P_btm.n3894 0.679419
R34304 C10_P_btm.n14 C10_P_btm.n12 0.672375
R34305 C10_P_btm.n470 C10_P_btm.n469 0.6255
R34306 C10_P_btm.n473 C10_P_btm.n472 0.6255
R34307 C10_P_btm.n476 C10_P_btm.n475 0.6255
R34308 C10_P_btm.n479 C10_P_btm.n478 0.6255
R34309 C10_P_btm.n482 C10_P_btm.n481 0.6255
R34310 C10_P_btm.n485 C10_P_btm.n484 0.6255
R34311 C10_P_btm.n488 C10_P_btm.n487 0.6255
R34312 C10_P_btm.n491 C10_P_btm.n490 0.6255
R34313 C10_P_btm.n494 C10_P_btm.n493 0.6255
R34314 C10_P_btm.n497 C10_P_btm.n496 0.6255
R34315 C10_P_btm.n500 C10_P_btm.n499 0.6255
R34316 C10_P_btm.n503 C10_P_btm.n502 0.6255
R34317 C10_P_btm.n2455 C10_P_btm.n2454 0.6255
R34318 C10_P_btm.n2452 C10_P_btm.n2451 0.6255
R34319 C10_P_btm.n2449 C10_P_btm.n2448 0.6255
R34320 C10_P_btm.n2446 C10_P_btm.n2445 0.6255
R34321 C10_P_btm.n2443 C10_P_btm.n2442 0.6255
R34322 C10_P_btm.n2440 C10_P_btm.n2439 0.6255
R34323 C10_P_btm.n2437 C10_P_btm.n2436 0.6255
R34324 C10_P_btm.n2434 C10_P_btm.n2433 0.6255
R34325 C10_P_btm.n2487 C10_P_btm.n2486 0.6255
R34326 C10_P_btm.n2484 C10_P_btm.n2483 0.6255
R34327 C10_P_btm.n2481 C10_P_btm.n2480 0.6255
R34328 C10_P_btm.n2478 C10_P_btm.n2477 0.6255
R34329 C10_P_btm.n2475 C10_P_btm.n2474 0.6255
R34330 C10_P_btm.n2472 C10_P_btm.n2471 0.6255
R34331 C10_P_btm.n2469 C10_P_btm.n2468 0.6255
R34332 C10_P_btm.n2466 C10_P_btm.n2465 0.6255
R34333 C10_P_btm.n2518 C10_P_btm.n2517 0.6255
R34334 C10_P_btm.n2515 C10_P_btm.n2514 0.6255
R34335 C10_P_btm.n2512 C10_P_btm.n2511 0.6255
R34336 C10_P_btm.n2509 C10_P_btm.n2508 0.6255
R34337 C10_P_btm.n2506 C10_P_btm.n2505 0.6255
R34338 C10_P_btm.n2503 C10_P_btm.n2502 0.6255
R34339 C10_P_btm.n2500 C10_P_btm.n2499 0.6255
R34340 C10_P_btm.n2497 C10_P_btm.n2496 0.6255
R34341 C10_P_btm.n2410 C10_P_btm.n2408 0.6255
R34342 C10_P_btm.n2406 C10_P_btm.n2405 0.6255
R34343 C10_P_btm.n2403 C10_P_btm.n2402 0.6255
R34344 C10_P_btm.n2400 C10_P_btm.n2399 0.6255
R34345 C10_P_btm.n2397 C10_P_btm.n2396 0.6255
R34346 C10_P_btm.n2394 C10_P_btm.n2393 0.6255
R34347 C10_P_btm.n2391 C10_P_btm.n2390 0.6255
R34348 C10_P_btm.n2388 C10_P_btm.n2370 0.6255
R34349 C10_P_btm.n2533 C10_P_btm.n2532 0.6255
R34350 C10_P_btm.n2536 C10_P_btm.n2535 0.6255
R34351 C10_P_btm.n2539 C10_P_btm.n2538 0.6255
R34352 C10_P_btm.n2542 C10_P_btm.n2541 0.6255
R34353 C10_P_btm.n2545 C10_P_btm.n2544 0.6255
R34354 C10_P_btm.n2548 C10_P_btm.n2547 0.6255
R34355 C10_P_btm.n2551 C10_P_btm.n2550 0.6255
R34356 C10_P_btm.n2554 C10_P_btm.n2553 0.6255
R34357 C10_P_btm.n2564 C10_P_btm.n2563 0.6255
R34358 C10_P_btm.n2567 C10_P_btm.n2566 0.6255
R34359 C10_P_btm.n2570 C10_P_btm.n2569 0.6255
R34360 C10_P_btm.n2573 C10_P_btm.n2572 0.6255
R34361 C10_P_btm.n2576 C10_P_btm.n2575 0.6255
R34362 C10_P_btm.n2579 C10_P_btm.n2578 0.6255
R34363 C10_P_btm.n2582 C10_P_btm.n2581 0.6255
R34364 C10_P_btm.n2585 C10_P_btm.n2584 0.6255
R34365 C10_P_btm.n2335 C10_P_btm.n2317 0.6255
R34366 C10_P_btm.n2338 C10_P_btm.n2337 0.6255
R34367 C10_P_btm.n2341 C10_P_btm.n2340 0.6255
R34368 C10_P_btm.n2344 C10_P_btm.n2343 0.6255
R34369 C10_P_btm.n2347 C10_P_btm.n2346 0.6255
R34370 C10_P_btm.n2350 C10_P_btm.n2349 0.6255
R34371 C10_P_btm.n2353 C10_P_btm.n2352 0.6255
R34372 C10_P_btm.n2357 C10_P_btm.n2355 0.6255
R34373 C10_P_btm.n2621 C10_P_btm.n2620 0.6255
R34374 C10_P_btm.n2618 C10_P_btm.n2617 0.6255
R34375 C10_P_btm.n2615 C10_P_btm.n2614 0.6255
R34376 C10_P_btm.n2612 C10_P_btm.n2611 0.6255
R34377 C10_P_btm.n2609 C10_P_btm.n2608 0.6255
R34378 C10_P_btm.n2606 C10_P_btm.n2605 0.6255
R34379 C10_P_btm.n2603 C10_P_btm.n2602 0.6255
R34380 C10_P_btm.n2600 C10_P_btm.n2599 0.6255
R34381 C10_P_btm.n2652 C10_P_btm.n2651 0.6255
R34382 C10_P_btm.n2649 C10_P_btm.n2648 0.6255
R34383 C10_P_btm.n2646 C10_P_btm.n2645 0.6255
R34384 C10_P_btm.n2643 C10_P_btm.n2642 0.6255
R34385 C10_P_btm.n2640 C10_P_btm.n2639 0.6255
R34386 C10_P_btm.n2637 C10_P_btm.n2636 0.6255
R34387 C10_P_btm.n2634 C10_P_btm.n2633 0.6255
R34388 C10_P_btm.n2631 C10_P_btm.n2630 0.6255
R34389 C10_P_btm.n2304 C10_P_btm.n2302 0.6255
R34390 C10_P_btm.n2300 C10_P_btm.n2299 0.6255
R34391 C10_P_btm.n2297 C10_P_btm.n2296 0.6255
R34392 C10_P_btm.n2294 C10_P_btm.n2293 0.6255
R34393 C10_P_btm.n2291 C10_P_btm.n2290 0.6255
R34394 C10_P_btm.n2288 C10_P_btm.n2287 0.6255
R34395 C10_P_btm.n2285 C10_P_btm.n2284 0.6255
R34396 C10_P_btm.n2282 C10_P_btm.n2264 0.6255
R34397 C10_P_btm.n2667 C10_P_btm.n2666 0.6255
R34398 C10_P_btm.n2670 C10_P_btm.n2669 0.6255
R34399 C10_P_btm.n2673 C10_P_btm.n2672 0.6255
R34400 C10_P_btm.n2676 C10_P_btm.n2675 0.6255
R34401 C10_P_btm.n2679 C10_P_btm.n2678 0.6255
R34402 C10_P_btm.n2682 C10_P_btm.n2681 0.6255
R34403 C10_P_btm.n2685 C10_P_btm.n2684 0.6255
R34404 C10_P_btm.n2688 C10_P_btm.n2687 0.6255
R34405 C10_P_btm.n2698 C10_P_btm.n2697 0.6255
R34406 C10_P_btm.n2701 C10_P_btm.n2700 0.6255
R34407 C10_P_btm.n2704 C10_P_btm.n2703 0.6255
R34408 C10_P_btm.n2707 C10_P_btm.n2706 0.6255
R34409 C10_P_btm.n2710 C10_P_btm.n2709 0.6255
R34410 C10_P_btm.n2713 C10_P_btm.n2712 0.6255
R34411 C10_P_btm.n2716 C10_P_btm.n2715 0.6255
R34412 C10_P_btm.n2719 C10_P_btm.n2718 0.6255
R34413 C10_P_btm.n2229 C10_P_btm.n2211 0.6255
R34414 C10_P_btm.n2232 C10_P_btm.n2231 0.6255
R34415 C10_P_btm.n2235 C10_P_btm.n2234 0.6255
R34416 C10_P_btm.n2238 C10_P_btm.n2237 0.6255
R34417 C10_P_btm.n2241 C10_P_btm.n2240 0.6255
R34418 C10_P_btm.n2244 C10_P_btm.n2243 0.6255
R34419 C10_P_btm.n2247 C10_P_btm.n2246 0.6255
R34420 C10_P_btm.n2251 C10_P_btm.n2249 0.6255
R34421 C10_P_btm.n2755 C10_P_btm.n2754 0.6255
R34422 C10_P_btm.n2752 C10_P_btm.n2751 0.6255
R34423 C10_P_btm.n2749 C10_P_btm.n2748 0.6255
R34424 C10_P_btm.n2746 C10_P_btm.n2745 0.6255
R34425 C10_P_btm.n2743 C10_P_btm.n2742 0.6255
R34426 C10_P_btm.n2740 C10_P_btm.n2739 0.6255
R34427 C10_P_btm.n2737 C10_P_btm.n2736 0.6255
R34428 C10_P_btm.n2734 C10_P_btm.n2733 0.6255
R34429 C10_P_btm.n2786 C10_P_btm.n2785 0.6255
R34430 C10_P_btm.n2783 C10_P_btm.n2782 0.6255
R34431 C10_P_btm.n2780 C10_P_btm.n2779 0.6255
R34432 C10_P_btm.n2777 C10_P_btm.n2776 0.6255
R34433 C10_P_btm.n2774 C10_P_btm.n2773 0.6255
R34434 C10_P_btm.n2771 C10_P_btm.n2770 0.6255
R34435 C10_P_btm.n2768 C10_P_btm.n2767 0.6255
R34436 C10_P_btm.n2765 C10_P_btm.n2764 0.6255
R34437 C10_P_btm.n2198 C10_P_btm.n2196 0.6255
R34438 C10_P_btm.n2194 C10_P_btm.n2193 0.6255
R34439 C10_P_btm.n2191 C10_P_btm.n2190 0.6255
R34440 C10_P_btm.n2188 C10_P_btm.n2187 0.6255
R34441 C10_P_btm.n2185 C10_P_btm.n2184 0.6255
R34442 C10_P_btm.n2182 C10_P_btm.n2181 0.6255
R34443 C10_P_btm.n2179 C10_P_btm.n2178 0.6255
R34444 C10_P_btm.n2176 C10_P_btm.n2158 0.6255
R34445 C10_P_btm.n2801 C10_P_btm.n2800 0.6255
R34446 C10_P_btm.n2804 C10_P_btm.n2803 0.6255
R34447 C10_P_btm.n2807 C10_P_btm.n2806 0.6255
R34448 C10_P_btm.n2810 C10_P_btm.n2809 0.6255
R34449 C10_P_btm.n2813 C10_P_btm.n2812 0.6255
R34450 C10_P_btm.n2816 C10_P_btm.n2815 0.6255
R34451 C10_P_btm.n2819 C10_P_btm.n2818 0.6255
R34452 C10_P_btm.n2822 C10_P_btm.n2821 0.6255
R34453 C10_P_btm.n2832 C10_P_btm.n2831 0.6255
R34454 C10_P_btm.n2835 C10_P_btm.n2834 0.6255
R34455 C10_P_btm.n2838 C10_P_btm.n2837 0.6255
R34456 C10_P_btm.n2841 C10_P_btm.n2840 0.6255
R34457 C10_P_btm.n2844 C10_P_btm.n2843 0.6255
R34458 C10_P_btm.n2847 C10_P_btm.n2846 0.6255
R34459 C10_P_btm.n2850 C10_P_btm.n2849 0.6255
R34460 C10_P_btm.n2853 C10_P_btm.n2852 0.6255
R34461 C10_P_btm.n2123 C10_P_btm.n2105 0.6255
R34462 C10_P_btm.n2126 C10_P_btm.n2125 0.6255
R34463 C10_P_btm.n2129 C10_P_btm.n2128 0.6255
R34464 C10_P_btm.n2132 C10_P_btm.n2131 0.6255
R34465 C10_P_btm.n2135 C10_P_btm.n2134 0.6255
R34466 C10_P_btm.n2138 C10_P_btm.n2137 0.6255
R34467 C10_P_btm.n2141 C10_P_btm.n2140 0.6255
R34468 C10_P_btm.n2145 C10_P_btm.n2143 0.6255
R34469 C10_P_btm.n2889 C10_P_btm.n2888 0.6255
R34470 C10_P_btm.n2886 C10_P_btm.n2885 0.6255
R34471 C10_P_btm.n2883 C10_P_btm.n2882 0.6255
R34472 C10_P_btm.n2880 C10_P_btm.n2879 0.6255
R34473 C10_P_btm.n2877 C10_P_btm.n2876 0.6255
R34474 C10_P_btm.n2874 C10_P_btm.n2873 0.6255
R34475 C10_P_btm.n2871 C10_P_btm.n2870 0.6255
R34476 C10_P_btm.n2868 C10_P_btm.n2867 0.6255
R34477 C10_P_btm.n2955 C10_P_btm.n2954 0.6255
R34478 C10_P_btm.n2952 C10_P_btm.n2951 0.6255
R34479 C10_P_btm.n2949 C10_P_btm.n2948 0.6255
R34480 C10_P_btm.n2946 C10_P_btm.n2945 0.6255
R34481 C10_P_btm.n2943 C10_P_btm.n2942 0.6255
R34482 C10_P_btm.n2940 C10_P_btm.n2939 0.6255
R34483 C10_P_btm.n2937 C10_P_btm.n2936 0.6255
R34484 C10_P_btm.n2934 C10_P_btm.n2933 0.6255
R34485 C10_P_btm.n2924 C10_P_btm.n2923 0.6255
R34486 C10_P_btm.n2921 C10_P_btm.n2920 0.6255
R34487 C10_P_btm.n2918 C10_P_btm.n2917 0.6255
R34488 C10_P_btm.n2915 C10_P_btm.n2914 0.6255
R34489 C10_P_btm.n2912 C10_P_btm.n2911 0.6255
R34490 C10_P_btm.n2909 C10_P_btm.n2908 0.6255
R34491 C10_P_btm.n2906 C10_P_btm.n2905 0.6255
R34492 C10_P_btm.n2903 C10_P_btm.n2085 0.6255
R34493 C10_P_btm.n2970 C10_P_btm.n2969 0.6255
R34494 C10_P_btm.n2973 C10_P_btm.n2972 0.6255
R34495 C10_P_btm.n2976 C10_P_btm.n2975 0.6255
R34496 C10_P_btm.n2979 C10_P_btm.n2978 0.6255
R34497 C10_P_btm.n2982 C10_P_btm.n2981 0.6255
R34498 C10_P_btm.n2985 C10_P_btm.n2984 0.6255
R34499 C10_P_btm.n2988 C10_P_btm.n2987 0.6255
R34500 C10_P_btm.n2992 C10_P_btm.n2990 0.6255
R34501 C10_P_btm.n2999 C10_P_btm.n2998 0.6255
R34502 C10_P_btm.n3002 C10_P_btm.n3001 0.6255
R34503 C10_P_btm.n3005 C10_P_btm.n3004 0.6255
R34504 C10_P_btm.n3008 C10_P_btm.n3007 0.6255
R34505 C10_P_btm.n3011 C10_P_btm.n3010 0.6255
R34506 C10_P_btm.n3014 C10_P_btm.n3013 0.6255
R34507 C10_P_btm.n3017 C10_P_btm.n3016 0.6255
R34508 C10_P_btm.n3020 C10_P_btm.n3019 0.6255
R34509 C10_P_btm.n3042 C10_P_btm.n3041 0.6255
R34510 C10_P_btm.n3045 C10_P_btm.n3044 0.6255
R34511 C10_P_btm.n3048 C10_P_btm.n3047 0.6255
R34512 C10_P_btm.n3051 C10_P_btm.n3050 0.6255
R34513 C10_P_btm.n3054 C10_P_btm.n3053 0.6255
R34514 C10_P_btm.n3057 C10_P_btm.n3056 0.6255
R34515 C10_P_btm.n3060 C10_P_btm.n3059 0.6255
R34516 C10_P_btm.n3063 C10_P_btm.n3062 0.6255
R34517 C10_P_btm.n3066 C10_P_btm.n3065 0.6255
R34518 C10_P_btm.n3069 C10_P_btm.n3068 0.6255
R34519 C10_P_btm.n3072 C10_P_btm.n3071 0.6255
R34520 C10_P_btm.n3075 C10_P_btm.n3074 0.6255
R34521 C10_P_btm.n3078 C10_P_btm.n3077 0.6255
R34522 C10_P_btm.n3081 C10_P_btm.n3080 0.6255
R34523 C10_P_btm.n3084 C10_P_btm.n3083 0.6255
R34524 C10_P_btm.n3087 C10_P_btm.n3086 0.6255
R34525 C10_P_btm.n3090 C10_P_btm.n3089 0.6255
R34526 C10_P_btm.n3093 C10_P_btm.n3092 0.6255
R34527 C10_P_btm.n3096 C10_P_btm.n3095 0.6255
R34528 C10_P_btm.n3099 C10_P_btm.n3098 0.6255
R34529 C10_P_btm.n3102 C10_P_btm.n3101 0.6255
R34530 C10_P_btm.n1292 C10_P_btm.n1291 0.6255
R34531 C10_P_btm.n1295 C10_P_btm.n1294 0.6255
R34532 C10_P_btm.n1298 C10_P_btm.n1297 0.6255
R34533 C10_P_btm.n1301 C10_P_btm.n1300 0.6255
R34534 C10_P_btm.n1304 C10_P_btm.n1303 0.6255
R34535 C10_P_btm.n1307 C10_P_btm.n1306 0.6255
R34536 C10_P_btm.n1310 C10_P_btm.n1309 0.6255
R34537 C10_P_btm.n1313 C10_P_btm.n1312 0.6255
R34538 C10_P_btm.n1316 C10_P_btm.n1315 0.6255
R34539 C10_P_btm.n1319 C10_P_btm.n1318 0.6255
R34540 C10_P_btm.n1322 C10_P_btm.n1321 0.6255
R34541 C10_P_btm.n1325 C10_P_btm.n1324 0.6255
R34542 C10_P_btm.n1328 C10_P_btm.n1327 0.6255
R34543 C10_P_btm.n1331 C10_P_btm.n1330 0.6255
R34544 C10_P_btm.n1334 C10_P_btm.n1333 0.6255
R34545 C10_P_btm.n1337 C10_P_btm.n1336 0.6255
R34546 C10_P_btm.n1340 C10_P_btm.n1339 0.6255
R34547 C10_P_btm.n1343 C10_P_btm.n1342 0.6255
R34548 C10_P_btm.n1346 C10_P_btm.n1345 0.6255
R34549 C10_P_btm.n1349 C10_P_btm.n1348 0.6255
R34550 C10_P_btm.n1352 C10_P_btm.n1351 0.6255
R34551 C10_P_btm.n1355 C10_P_btm.n1354 0.6255
R34552 C10_P_btm.n1358 C10_P_btm.n1357 0.6255
R34553 C10_P_btm.n1361 C10_P_btm.n1360 0.6255
R34554 C10_P_btm.n1364 C10_P_btm.n1363 0.6255
R34555 C10_P_btm.n1367 C10_P_btm.n1366 0.6255
R34556 C10_P_btm.n1370 C10_P_btm.n1369 0.6255
R34557 C10_P_btm.n1373 C10_P_btm.n1372 0.6255
R34558 C10_P_btm.n1376 C10_P_btm.n1375 0.6255
R34559 C10_P_btm.n1379 C10_P_btm.n1378 0.6255
R34560 C10_P_btm.n1382 C10_P_btm.n1381 0.6255
R34561 C10_P_btm.n1385 C10_P_btm.n1384 0.6255
R34562 C10_P_btm.n1388 C10_P_btm.n1387 0.6255
R34563 C10_P_btm.n1391 C10_P_btm.n1390 0.6255
R34564 C10_P_btm.n1394 C10_P_btm.n1393 0.6255
R34565 C10_P_btm.n1397 C10_P_btm.n1396 0.6255
R34566 C10_P_btm.n1400 C10_P_btm.n1399 0.6255
R34567 C10_P_btm.n1403 C10_P_btm.n1402 0.6255
R34568 C10_P_btm.n1406 C10_P_btm.n1405 0.6255
R34569 C10_P_btm.n1409 C10_P_btm.n1408 0.6255
R34570 C10_P_btm.n1412 C10_P_btm.n1411 0.6255
R34571 C10_P_btm.n1415 C10_P_btm.n1414 0.6255
R34572 C10_P_btm.n1418 C10_P_btm.n1417 0.6255
R34573 C10_P_btm.n1421 C10_P_btm.n1420 0.6255
R34574 C10_P_btm.n1424 C10_P_btm.n1423 0.6255
R34575 C10_P_btm.n1427 C10_P_btm.n1426 0.6255
R34576 C10_P_btm.n1430 C10_P_btm.n1429 0.6255
R34577 C10_P_btm.n1433 C10_P_btm.n1432 0.6255
R34578 C10_P_btm.n1436 C10_P_btm.n1435 0.6255
R34579 C10_P_btm.n1439 C10_P_btm.n1438 0.6255
R34580 C10_P_btm.n1442 C10_P_btm.n1441 0.6255
R34581 C10_P_btm.n1445 C10_P_btm.n1444 0.6255
R34582 C10_P_btm.n1448 C10_P_btm.n1447 0.6255
R34583 C10_P_btm.n1451 C10_P_btm.n1450 0.6255
R34584 C10_P_btm.n1454 C10_P_btm.n1453 0.6255
R34585 C10_P_btm.n1457 C10_P_btm.n1456 0.6255
R34586 C10_P_btm.n1460 C10_P_btm.n1459 0.6255
R34587 C10_P_btm.n1463 C10_P_btm.n1462 0.6255
R34588 C10_P_btm.n1466 C10_P_btm.n1465 0.6255
R34589 C10_P_btm.n1469 C10_P_btm.n1468 0.6255
R34590 C10_P_btm.n1472 C10_P_btm.n1471 0.6255
R34591 C10_P_btm.n1104 C10_P_btm.n981 0.6255
R34592 C10_P_btm.n1107 C10_P_btm.n1106 0.6255
R34593 C10_P_btm.n1110 C10_P_btm.n1109 0.6255
R34594 C10_P_btm.n1113 C10_P_btm.n1112 0.6255
R34595 C10_P_btm.n1116 C10_P_btm.n1115 0.6255
R34596 C10_P_btm.n1119 C10_P_btm.n1118 0.6255
R34597 C10_P_btm.n1122 C10_P_btm.n1121 0.6255
R34598 C10_P_btm.n1125 C10_P_btm.n1124 0.6255
R34599 C10_P_btm.n1128 C10_P_btm.n1127 0.6255
R34600 C10_P_btm.n1131 C10_P_btm.n1130 0.6255
R34601 C10_P_btm.n1134 C10_P_btm.n1133 0.6255
R34602 C10_P_btm.n1137 C10_P_btm.n1136 0.6255
R34603 C10_P_btm.n1140 C10_P_btm.n1139 0.6255
R34604 C10_P_btm.n1143 C10_P_btm.n1142 0.6255
R34605 C10_P_btm.n1146 C10_P_btm.n1145 0.6255
R34606 C10_P_btm.n1149 C10_P_btm.n1148 0.6255
R34607 C10_P_btm.n1152 C10_P_btm.n1151 0.6255
R34608 C10_P_btm.n1155 C10_P_btm.n1154 0.6255
R34609 C10_P_btm.n1158 C10_P_btm.n1157 0.6255
R34610 C10_P_btm.n1161 C10_P_btm.n1160 0.6255
R34611 C10_P_btm.n1164 C10_P_btm.n1163 0.6255
R34612 C10_P_btm.n1167 C10_P_btm.n1166 0.6255
R34613 C10_P_btm.n1170 C10_P_btm.n1169 0.6255
R34614 C10_P_btm.n1173 C10_P_btm.n1172 0.6255
R34615 C10_P_btm.n1176 C10_P_btm.n1175 0.6255
R34616 C10_P_btm.n1179 C10_P_btm.n1178 0.6255
R34617 C10_P_btm.n1182 C10_P_btm.n1181 0.6255
R34618 C10_P_btm.n1185 C10_P_btm.n1184 0.6255
R34619 C10_P_btm.n1188 C10_P_btm.n1187 0.6255
R34620 C10_P_btm.n1191 C10_P_btm.n1190 0.6255
R34621 C10_P_btm.n1194 C10_P_btm.n1193 0.6255
R34622 C10_P_btm.n1197 C10_P_btm.n1196 0.6255
R34623 C10_P_btm.n1200 C10_P_btm.n1199 0.6255
R34624 C10_P_btm.n1203 C10_P_btm.n1202 0.6255
R34625 C10_P_btm.n1206 C10_P_btm.n1205 0.6255
R34626 C10_P_btm.n1209 C10_P_btm.n1208 0.6255
R34627 C10_P_btm.n1212 C10_P_btm.n1211 0.6255
R34628 C10_P_btm.n1215 C10_P_btm.n1214 0.6255
R34629 C10_P_btm.n1218 C10_P_btm.n1217 0.6255
R34630 C10_P_btm.n1221 C10_P_btm.n1220 0.6255
R34631 C10_P_btm.n1224 C10_P_btm.n1223 0.6255
R34632 C10_P_btm.n1227 C10_P_btm.n1226 0.6255
R34633 C10_P_btm.n1230 C10_P_btm.n1229 0.6255
R34634 C10_P_btm.n1233 C10_P_btm.n1232 0.6255
R34635 C10_P_btm.n1236 C10_P_btm.n1235 0.6255
R34636 C10_P_btm.n1239 C10_P_btm.n1238 0.6255
R34637 C10_P_btm.n1242 C10_P_btm.n1241 0.6255
R34638 C10_P_btm.n1245 C10_P_btm.n1244 0.6255
R34639 C10_P_btm.n1248 C10_P_btm.n1247 0.6255
R34640 C10_P_btm.n1251 C10_P_btm.n1250 0.6255
R34641 C10_P_btm.n1254 C10_P_btm.n1253 0.6255
R34642 C10_P_btm.n1257 C10_P_btm.n1256 0.6255
R34643 C10_P_btm.n1260 C10_P_btm.n1259 0.6255
R34644 C10_P_btm.n1263 C10_P_btm.n1262 0.6255
R34645 C10_P_btm.n1266 C10_P_btm.n1265 0.6255
R34646 C10_P_btm.n1269 C10_P_btm.n1268 0.6255
R34647 C10_P_btm.n1272 C10_P_btm.n1271 0.6255
R34648 C10_P_btm.n1275 C10_P_btm.n1274 0.6255
R34649 C10_P_btm.n1278 C10_P_btm.n1277 0.6255
R34650 C10_P_btm.n1281 C10_P_btm.n1280 0.6255
R34651 C10_P_btm.n1285 C10_P_btm.n1283 0.6255
R34652 C10_P_btm.n1666 C10_P_btm.n1665 0.6255
R34653 C10_P_btm.n1663 C10_P_btm.n1662 0.6255
R34654 C10_P_btm.n1660 C10_P_btm.n1659 0.6255
R34655 C10_P_btm.n1657 C10_P_btm.n1656 0.6255
R34656 C10_P_btm.n1654 C10_P_btm.n1653 0.6255
R34657 C10_P_btm.n1651 C10_P_btm.n1650 0.6255
R34658 C10_P_btm.n1648 C10_P_btm.n1647 0.6255
R34659 C10_P_btm.n1645 C10_P_btm.n1644 0.6255
R34660 C10_P_btm.n1642 C10_P_btm.n1641 0.6255
R34661 C10_P_btm.n1639 C10_P_btm.n1638 0.6255
R34662 C10_P_btm.n1636 C10_P_btm.n1635 0.6255
R34663 C10_P_btm.n1633 C10_P_btm.n1632 0.6255
R34664 C10_P_btm.n1630 C10_P_btm.n1629 0.6255
R34665 C10_P_btm.n1627 C10_P_btm.n1626 0.6255
R34666 C10_P_btm.n1624 C10_P_btm.n1623 0.6255
R34667 C10_P_btm.n1621 C10_P_btm.n1620 0.6255
R34668 C10_P_btm.n1618 C10_P_btm.n1617 0.6255
R34669 C10_P_btm.n1615 C10_P_btm.n1614 0.6255
R34670 C10_P_btm.n1612 C10_P_btm.n1611 0.6255
R34671 C10_P_btm.n1609 C10_P_btm.n1608 0.6255
R34672 C10_P_btm.n1606 C10_P_btm.n1605 0.6255
R34673 C10_P_btm.n1603 C10_P_btm.n1602 0.6255
R34674 C10_P_btm.n1600 C10_P_btm.n1599 0.6255
R34675 C10_P_btm.n1597 C10_P_btm.n1596 0.6255
R34676 C10_P_btm.n1594 C10_P_btm.n1593 0.6255
R34677 C10_P_btm.n1591 C10_P_btm.n1590 0.6255
R34678 C10_P_btm.n1588 C10_P_btm.n1587 0.6255
R34679 C10_P_btm.n1585 C10_P_btm.n1584 0.6255
R34680 C10_P_btm.n1582 C10_P_btm.n1581 0.6255
R34681 C10_P_btm.n1579 C10_P_btm.n1578 0.6255
R34682 C10_P_btm.n1576 C10_P_btm.n1575 0.6255
R34683 C10_P_btm.n1573 C10_P_btm.n1572 0.6255
R34684 C10_P_btm.n1570 C10_P_btm.n1569 0.6255
R34685 C10_P_btm.n1567 C10_P_btm.n1566 0.6255
R34686 C10_P_btm.n1564 C10_P_btm.n1563 0.6255
R34687 C10_P_btm.n1561 C10_P_btm.n1560 0.6255
R34688 C10_P_btm.n1558 C10_P_btm.n1557 0.6255
R34689 C10_P_btm.n1555 C10_P_btm.n1554 0.6255
R34690 C10_P_btm.n1552 C10_P_btm.n1551 0.6255
R34691 C10_P_btm.n1549 C10_P_btm.n1548 0.6255
R34692 C10_P_btm.n1546 C10_P_btm.n1545 0.6255
R34693 C10_P_btm.n1543 C10_P_btm.n1542 0.6255
R34694 C10_P_btm.n1540 C10_P_btm.n1539 0.6255
R34695 C10_P_btm.n1537 C10_P_btm.n1536 0.6255
R34696 C10_P_btm.n1534 C10_P_btm.n1533 0.6255
R34697 C10_P_btm.n1531 C10_P_btm.n1530 0.6255
R34698 C10_P_btm.n1528 C10_P_btm.n1527 0.6255
R34699 C10_P_btm.n1525 C10_P_btm.n1524 0.6255
R34700 C10_P_btm.n1522 C10_P_btm.n1521 0.6255
R34701 C10_P_btm.n1519 C10_P_btm.n1518 0.6255
R34702 C10_P_btm.n1516 C10_P_btm.n1515 0.6255
R34703 C10_P_btm.n1513 C10_P_btm.n1512 0.6255
R34704 C10_P_btm.n1510 C10_P_btm.n1509 0.6255
R34705 C10_P_btm.n1507 C10_P_btm.n1506 0.6255
R34706 C10_P_btm.n1504 C10_P_btm.n1503 0.6255
R34707 C10_P_btm.n1501 C10_P_btm.n1500 0.6255
R34708 C10_P_btm.n1498 C10_P_btm.n1497 0.6255
R34709 C10_P_btm.n1495 C10_P_btm.n1494 0.6255
R34710 C10_P_btm.n1492 C10_P_btm.n1491 0.6255
R34711 C10_P_btm.n1489 C10_P_btm.n1488 0.6255
R34712 C10_P_btm.n1486 C10_P_btm.n1485 0.6255
R34713 C10_P_btm.n1856 C10_P_btm.n1855 0.6255
R34714 C10_P_btm.n1853 C10_P_btm.n1852 0.6255
R34715 C10_P_btm.n1850 C10_P_btm.n1849 0.6255
R34716 C10_P_btm.n1847 C10_P_btm.n1846 0.6255
R34717 C10_P_btm.n1844 C10_P_btm.n1843 0.6255
R34718 C10_P_btm.n1841 C10_P_btm.n1840 0.6255
R34719 C10_P_btm.n1838 C10_P_btm.n1837 0.6255
R34720 C10_P_btm.n1835 C10_P_btm.n1834 0.6255
R34721 C10_P_btm.n1832 C10_P_btm.n1831 0.6255
R34722 C10_P_btm.n1829 C10_P_btm.n1828 0.6255
R34723 C10_P_btm.n1826 C10_P_btm.n1825 0.6255
R34724 C10_P_btm.n1823 C10_P_btm.n1822 0.6255
R34725 C10_P_btm.n1820 C10_P_btm.n1819 0.6255
R34726 C10_P_btm.n1817 C10_P_btm.n1816 0.6255
R34727 C10_P_btm.n1814 C10_P_btm.n1813 0.6255
R34728 C10_P_btm.n1811 C10_P_btm.n1810 0.6255
R34729 C10_P_btm.n1808 C10_P_btm.n1807 0.6255
R34730 C10_P_btm.n1805 C10_P_btm.n1804 0.6255
R34731 C10_P_btm.n1802 C10_P_btm.n1801 0.6255
R34732 C10_P_btm.n1799 C10_P_btm.n1798 0.6255
R34733 C10_P_btm.n1796 C10_P_btm.n1795 0.6255
R34734 C10_P_btm.n1793 C10_P_btm.n1792 0.6255
R34735 C10_P_btm.n1790 C10_P_btm.n1789 0.6255
R34736 C10_P_btm.n1787 C10_P_btm.n1786 0.6255
R34737 C10_P_btm.n1784 C10_P_btm.n1783 0.6255
R34738 C10_P_btm.n1781 C10_P_btm.n1780 0.6255
R34739 C10_P_btm.n1778 C10_P_btm.n1777 0.6255
R34740 C10_P_btm.n1775 C10_P_btm.n1774 0.6255
R34741 C10_P_btm.n1772 C10_P_btm.n1771 0.6255
R34742 C10_P_btm.n1769 C10_P_btm.n1768 0.6255
R34743 C10_P_btm.n1766 C10_P_btm.n1765 0.6255
R34744 C10_P_btm.n1763 C10_P_btm.n1762 0.6255
R34745 C10_P_btm.n1760 C10_P_btm.n1759 0.6255
R34746 C10_P_btm.n1757 C10_P_btm.n1756 0.6255
R34747 C10_P_btm.n1754 C10_P_btm.n1753 0.6255
R34748 C10_P_btm.n1751 C10_P_btm.n1750 0.6255
R34749 C10_P_btm.n1748 C10_P_btm.n1747 0.6255
R34750 C10_P_btm.n1745 C10_P_btm.n1744 0.6255
R34751 C10_P_btm.n1742 C10_P_btm.n1741 0.6255
R34752 C10_P_btm.n1739 C10_P_btm.n1738 0.6255
R34753 C10_P_btm.n1736 C10_P_btm.n1735 0.6255
R34754 C10_P_btm.n1733 C10_P_btm.n1732 0.6255
R34755 C10_P_btm.n1730 C10_P_btm.n1729 0.6255
R34756 C10_P_btm.n1727 C10_P_btm.n1726 0.6255
R34757 C10_P_btm.n1724 C10_P_btm.n1723 0.6255
R34758 C10_P_btm.n1721 C10_P_btm.n1720 0.6255
R34759 C10_P_btm.n1718 C10_P_btm.n1717 0.6255
R34760 C10_P_btm.n1715 C10_P_btm.n1714 0.6255
R34761 C10_P_btm.n1712 C10_P_btm.n1711 0.6255
R34762 C10_P_btm.n1709 C10_P_btm.n1708 0.6255
R34763 C10_P_btm.n1706 C10_P_btm.n1705 0.6255
R34764 C10_P_btm.n1703 C10_P_btm.n1702 0.6255
R34765 C10_P_btm.n1700 C10_P_btm.n1699 0.6255
R34766 C10_P_btm.n1697 C10_P_btm.n1696 0.6255
R34767 C10_P_btm.n1694 C10_P_btm.n1693 0.6255
R34768 C10_P_btm.n1691 C10_P_btm.n1690 0.6255
R34769 C10_P_btm.n1688 C10_P_btm.n1687 0.6255
R34770 C10_P_btm.n1685 C10_P_btm.n1684 0.6255
R34771 C10_P_btm.n1682 C10_P_btm.n1681 0.6255
R34772 C10_P_btm.n1679 C10_P_btm.n1678 0.6255
R34773 C10_P_btm.n1676 C10_P_btm.n1675 0.6255
R34774 C10_P_btm.n915 C10_P_btm.n913 0.6255
R34775 C10_P_btm.n911 C10_P_btm.n910 0.6255
R34776 C10_P_btm.n908 C10_P_btm.n907 0.6255
R34777 C10_P_btm.n905 C10_P_btm.n904 0.6255
R34778 C10_P_btm.n902 C10_P_btm.n901 0.6255
R34779 C10_P_btm.n899 C10_P_btm.n898 0.6255
R34780 C10_P_btm.n896 C10_P_btm.n895 0.6255
R34781 C10_P_btm.n893 C10_P_btm.n892 0.6255
R34782 C10_P_btm.n890 C10_P_btm.n889 0.6255
R34783 C10_P_btm.n887 C10_P_btm.n886 0.6255
R34784 C10_P_btm.n884 C10_P_btm.n883 0.6255
R34785 C10_P_btm.n881 C10_P_btm.n880 0.6255
R34786 C10_P_btm.n878 C10_P_btm.n877 0.6255
R34787 C10_P_btm.n875 C10_P_btm.n874 0.6255
R34788 C10_P_btm.n872 C10_P_btm.n871 0.6255
R34789 C10_P_btm.n869 C10_P_btm.n868 0.6255
R34790 C10_P_btm.n866 C10_P_btm.n865 0.6255
R34791 C10_P_btm.n863 C10_P_btm.n862 0.6255
R34792 C10_P_btm.n860 C10_P_btm.n859 0.6255
R34793 C10_P_btm.n857 C10_P_btm.n856 0.6255
R34794 C10_P_btm.n854 C10_P_btm.n853 0.6255
R34795 C10_P_btm.n851 C10_P_btm.n850 0.6255
R34796 C10_P_btm.n848 C10_P_btm.n847 0.6255
R34797 C10_P_btm.n845 C10_P_btm.n844 0.6255
R34798 C10_P_btm.n842 C10_P_btm.n841 0.6255
R34799 C10_P_btm.n839 C10_P_btm.n838 0.6255
R34800 C10_P_btm.n836 C10_P_btm.n835 0.6255
R34801 C10_P_btm.n833 C10_P_btm.n832 0.6255
R34802 C10_P_btm.n830 C10_P_btm.n829 0.6255
R34803 C10_P_btm.n827 C10_P_btm.n826 0.6255
R34804 C10_P_btm.n824 C10_P_btm.n823 0.6255
R34805 C10_P_btm.n821 C10_P_btm.n820 0.6255
R34806 C10_P_btm.n818 C10_P_btm.n817 0.6255
R34807 C10_P_btm.n815 C10_P_btm.n814 0.6255
R34808 C10_P_btm.n812 C10_P_btm.n811 0.6255
R34809 C10_P_btm.n809 C10_P_btm.n808 0.6255
R34810 C10_P_btm.n806 C10_P_btm.n805 0.6255
R34811 C10_P_btm.n803 C10_P_btm.n802 0.6255
R34812 C10_P_btm.n800 C10_P_btm.n799 0.6255
R34813 C10_P_btm.n797 C10_P_btm.n796 0.6255
R34814 C10_P_btm.n794 C10_P_btm.n793 0.6255
R34815 C10_P_btm.n791 C10_P_btm.n790 0.6255
R34816 C10_P_btm.n788 C10_P_btm.n787 0.6255
R34817 C10_P_btm.n785 C10_P_btm.n784 0.6255
R34818 C10_P_btm.n782 C10_P_btm.n781 0.6255
R34819 C10_P_btm.n779 C10_P_btm.n778 0.6255
R34820 C10_P_btm.n776 C10_P_btm.n775 0.6255
R34821 C10_P_btm.n773 C10_P_btm.n772 0.6255
R34822 C10_P_btm.n770 C10_P_btm.n769 0.6255
R34823 C10_P_btm.n767 C10_P_btm.n766 0.6255
R34824 C10_P_btm.n764 C10_P_btm.n763 0.6255
R34825 C10_P_btm.n761 C10_P_btm.n760 0.6255
R34826 C10_P_btm.n758 C10_P_btm.n757 0.6255
R34827 C10_P_btm.n755 C10_P_btm.n754 0.6255
R34828 C10_P_btm.n752 C10_P_btm.n751 0.6255
R34829 C10_P_btm.n749 C10_P_btm.n748 0.6255
R34830 C10_P_btm.n746 C10_P_btm.n745 0.6255
R34831 C10_P_btm.n743 C10_P_btm.n742 0.6255
R34832 C10_P_btm.n740 C10_P_btm.n739 0.6255
R34833 C10_P_btm.n737 C10_P_btm.n736 0.6255
R34834 C10_P_btm.n734 C10_P_btm.n610 0.6255
R34835 C10_P_btm.n1871 C10_P_btm.n1870 0.6255
R34836 C10_P_btm.n1874 C10_P_btm.n1873 0.6255
R34837 C10_P_btm.n1877 C10_P_btm.n1876 0.6255
R34838 C10_P_btm.n1880 C10_P_btm.n1879 0.6255
R34839 C10_P_btm.n1883 C10_P_btm.n1882 0.6255
R34840 C10_P_btm.n1886 C10_P_btm.n1885 0.6255
R34841 C10_P_btm.n1889 C10_P_btm.n1888 0.6255
R34842 C10_P_btm.n1892 C10_P_btm.n1891 0.6255
R34843 C10_P_btm.n1895 C10_P_btm.n1894 0.6255
R34844 C10_P_btm.n1898 C10_P_btm.n1897 0.6255
R34845 C10_P_btm.n1901 C10_P_btm.n1900 0.6255
R34846 C10_P_btm.n1904 C10_P_btm.n1903 0.6255
R34847 C10_P_btm.n1907 C10_P_btm.n1906 0.6255
R34848 C10_P_btm.n1910 C10_P_btm.n1909 0.6255
R34849 C10_P_btm.n1913 C10_P_btm.n1912 0.6255
R34850 C10_P_btm.n1916 C10_P_btm.n1915 0.6255
R34851 C10_P_btm.n1919 C10_P_btm.n1918 0.6255
R34852 C10_P_btm.n1922 C10_P_btm.n1921 0.6255
R34853 C10_P_btm.n1925 C10_P_btm.n1924 0.6255
R34854 C10_P_btm.n1928 C10_P_btm.n1927 0.6255
R34855 C10_P_btm.n1931 C10_P_btm.n1930 0.6255
R34856 C10_P_btm.n1934 C10_P_btm.n1933 0.6255
R34857 C10_P_btm.n1937 C10_P_btm.n1936 0.6255
R34858 C10_P_btm.n1940 C10_P_btm.n1939 0.6255
R34859 C10_P_btm.n1943 C10_P_btm.n1942 0.6255
R34860 C10_P_btm.n1946 C10_P_btm.n1945 0.6255
R34861 C10_P_btm.n1949 C10_P_btm.n1948 0.6255
R34862 C10_P_btm.n1952 C10_P_btm.n1951 0.6255
R34863 C10_P_btm.n1955 C10_P_btm.n1954 0.6255
R34864 C10_P_btm.n1958 C10_P_btm.n1957 0.6255
R34865 C10_P_btm.n1961 C10_P_btm.n1960 0.6255
R34866 C10_P_btm.n1964 C10_P_btm.n1963 0.6255
R34867 C10_P_btm.n1967 C10_P_btm.n1966 0.6255
R34868 C10_P_btm.n1970 C10_P_btm.n1969 0.6255
R34869 C10_P_btm.n1973 C10_P_btm.n1972 0.6255
R34870 C10_P_btm.n1976 C10_P_btm.n1975 0.6255
R34871 C10_P_btm.n1979 C10_P_btm.n1978 0.6255
R34872 C10_P_btm.n1982 C10_P_btm.n1981 0.6255
R34873 C10_P_btm.n1985 C10_P_btm.n1984 0.6255
R34874 C10_P_btm.n1988 C10_P_btm.n1987 0.6255
R34875 C10_P_btm.n1991 C10_P_btm.n1990 0.6255
R34876 C10_P_btm.n1994 C10_P_btm.n1993 0.6255
R34877 C10_P_btm.n1997 C10_P_btm.n1996 0.6255
R34878 C10_P_btm.n2000 C10_P_btm.n1999 0.6255
R34879 C10_P_btm.n2003 C10_P_btm.n2002 0.6255
R34880 C10_P_btm.n2006 C10_P_btm.n2005 0.6255
R34881 C10_P_btm.n2009 C10_P_btm.n2008 0.6255
R34882 C10_P_btm.n2012 C10_P_btm.n2011 0.6255
R34883 C10_P_btm.n2015 C10_P_btm.n2014 0.6255
R34884 C10_P_btm.n2018 C10_P_btm.n2017 0.6255
R34885 C10_P_btm.n2021 C10_P_btm.n2020 0.6255
R34886 C10_P_btm.n2024 C10_P_btm.n2023 0.6255
R34887 C10_P_btm.n2027 C10_P_btm.n2026 0.6255
R34888 C10_P_btm.n2030 C10_P_btm.n2029 0.6255
R34889 C10_P_btm.n2033 C10_P_btm.n2032 0.6255
R34890 C10_P_btm.n2036 C10_P_btm.n2035 0.6255
R34891 C10_P_btm.n2039 C10_P_btm.n2038 0.6255
R34892 C10_P_btm.n2042 C10_P_btm.n2041 0.6255
R34893 C10_P_btm.n2045 C10_P_btm.n2044 0.6255
R34894 C10_P_btm.n2048 C10_P_btm.n2047 0.6255
R34895 C10_P_btm.n2051 C10_P_btm.n2050 0.6255
R34896 C10_P_btm.n3112 C10_P_btm.n3111 0.6255
R34897 C10_P_btm.n3115 C10_P_btm.n3114 0.6255
R34898 C10_P_btm.n3118 C10_P_btm.n3117 0.6255
R34899 C10_P_btm.n3121 C10_P_btm.n3120 0.6255
R34900 C10_P_btm.n3124 C10_P_btm.n3123 0.6255
R34901 C10_P_btm.n3127 C10_P_btm.n3126 0.6255
R34902 C10_P_btm.n3130 C10_P_btm.n3129 0.6255
R34903 C10_P_btm.n3133 C10_P_btm.n3132 0.6255
R34904 C10_P_btm.n3136 C10_P_btm.n3135 0.6255
R34905 C10_P_btm.n3139 C10_P_btm.n3138 0.6255
R34906 C10_P_btm.n3142 C10_P_btm.n3141 0.6255
R34907 C10_P_btm.n3145 C10_P_btm.n3144 0.6255
R34908 C10_P_btm.n3148 C10_P_btm.n3147 0.6255
R34909 C10_P_btm.n3151 C10_P_btm.n3150 0.6255
R34910 C10_P_btm.n3154 C10_P_btm.n3153 0.6255
R34911 C10_P_btm.n3157 C10_P_btm.n3156 0.6255
R34912 C10_P_btm.n3160 C10_P_btm.n3159 0.6255
R34913 C10_P_btm.n3163 C10_P_btm.n3162 0.6255
R34914 C10_P_btm.n3166 C10_P_btm.n3165 0.6255
R34915 C10_P_btm.n3169 C10_P_btm.n3168 0.6255
R34916 C10_P_btm.n3172 C10_P_btm.n3171 0.6255
R34917 C10_P_btm.n3175 C10_P_btm.n3174 0.6255
R34918 C10_P_btm.n3178 C10_P_btm.n3177 0.6255
R34919 C10_P_btm.n3181 C10_P_btm.n3180 0.6255
R34920 C10_P_btm.n3184 C10_P_btm.n3183 0.6255
R34921 C10_P_btm.n3187 C10_P_btm.n3186 0.6255
R34922 C10_P_btm.n3190 C10_P_btm.n3189 0.6255
R34923 C10_P_btm.n3193 C10_P_btm.n3192 0.6255
R34924 C10_P_btm.n3196 C10_P_btm.n3195 0.6255
R34925 C10_P_btm.n3199 C10_P_btm.n3198 0.6255
R34926 C10_P_btm.n3202 C10_P_btm.n3201 0.6255
R34927 C10_P_btm.n3205 C10_P_btm.n3204 0.6255
R34928 C10_P_btm.n3208 C10_P_btm.n3207 0.6255
R34929 C10_P_btm.n3211 C10_P_btm.n3210 0.6255
R34930 C10_P_btm.n3214 C10_P_btm.n3213 0.6255
R34931 C10_P_btm.n3217 C10_P_btm.n3216 0.6255
R34932 C10_P_btm.n3220 C10_P_btm.n3219 0.6255
R34933 C10_P_btm.n3223 C10_P_btm.n3222 0.6255
R34934 C10_P_btm.n3226 C10_P_btm.n3225 0.6255
R34935 C10_P_btm.n3229 C10_P_btm.n3228 0.6255
R34936 C10_P_btm.n3232 C10_P_btm.n3231 0.6255
R34937 C10_P_btm.n3235 C10_P_btm.n3234 0.6255
R34938 C10_P_btm.n3238 C10_P_btm.n3237 0.6255
R34939 C10_P_btm.n3241 C10_P_btm.n3240 0.6255
R34940 C10_P_btm.n3244 C10_P_btm.n3243 0.6255
R34941 C10_P_btm.n3247 C10_P_btm.n3246 0.6255
R34942 C10_P_btm.n3250 C10_P_btm.n3249 0.6255
R34943 C10_P_btm.n3253 C10_P_btm.n3252 0.6255
R34944 C10_P_btm.n3256 C10_P_btm.n3255 0.6255
R34945 C10_P_btm.n3259 C10_P_btm.n3258 0.6255
R34946 C10_P_btm.n3262 C10_P_btm.n3261 0.6255
R34947 C10_P_btm.n3265 C10_P_btm.n3264 0.6255
R34948 C10_P_btm.n3268 C10_P_btm.n3267 0.6255
R34949 C10_P_btm.n3271 C10_P_btm.n3270 0.6255
R34950 C10_P_btm.n3274 C10_P_btm.n3273 0.6255
R34951 C10_P_btm.n3277 C10_P_btm.n3276 0.6255
R34952 C10_P_btm.n3280 C10_P_btm.n3279 0.6255
R34953 C10_P_btm.n3283 C10_P_btm.n3282 0.6255
R34954 C10_P_btm.n3286 C10_P_btm.n3285 0.6255
R34955 C10_P_btm.n3289 C10_P_btm.n3288 0.6255
R34956 C10_P_btm.n3292 C10_P_btm.n3291 0.6255
R34957 C10_P_btm.n443 C10_P_btm.n400 0.6255
R34958 C10_P_btm.n446 C10_P_btm.n445 0.6255
R34959 C10_P_btm.n449 C10_P_btm.n448 0.6255
R34960 C10_P_btm.n452 C10_P_btm.n451 0.6255
R34961 C10_P_btm.n455 C10_P_btm.n454 0.6255
R34962 C10_P_btm.n458 C10_P_btm.n457 0.6255
R34963 C10_P_btm.n461 C10_P_btm.n460 0.6255
R34964 C10_P_btm.n464 C10_P_btm.n463 0.6255
R34965 C10_P_btm.n467 C10_P_btm.n466 0.6255
R34966 C10_P_btm.n3328 C10_P_btm.n3327 0.6255
R34967 C10_P_btm.n3325 C10_P_btm.n3324 0.6255
R34968 C10_P_btm.n3322 C10_P_btm.n3321 0.6255
R34969 C10_P_btm.n3319 C10_P_btm.n3318 0.6255
R34970 C10_P_btm.n3316 C10_P_btm.n3315 0.6255
R34971 C10_P_btm.n3313 C10_P_btm.n3312 0.6255
R34972 C10_P_btm.n3310 C10_P_btm.n3309 0.6255
R34973 C10_P_btm.n3307 C10_P_btm.n3306 0.6255
R34974 C10_P_btm.n3359 C10_P_btm.n3358 0.6255
R34975 C10_P_btm.n3356 C10_P_btm.n3355 0.6255
R34976 C10_P_btm.n3353 C10_P_btm.n3352 0.6255
R34977 C10_P_btm.n3350 C10_P_btm.n3349 0.6255
R34978 C10_P_btm.n3347 C10_P_btm.n3346 0.6255
R34979 C10_P_btm.n3344 C10_P_btm.n3343 0.6255
R34980 C10_P_btm.n3341 C10_P_btm.n3340 0.6255
R34981 C10_P_btm.n3338 C10_P_btm.n3337 0.6255
R34982 C10_P_btm.n387 C10_P_btm.n385 0.6255
R34983 C10_P_btm.n383 C10_P_btm.n382 0.6255
R34984 C10_P_btm.n380 C10_P_btm.n379 0.6255
R34985 C10_P_btm.n377 C10_P_btm.n376 0.6255
R34986 C10_P_btm.n374 C10_P_btm.n373 0.6255
R34987 C10_P_btm.n371 C10_P_btm.n370 0.6255
R34988 C10_P_btm.n368 C10_P_btm.n367 0.6255
R34989 C10_P_btm.n365 C10_P_btm.n347 0.6255
R34990 C10_P_btm.n3374 C10_P_btm.n3373 0.6255
R34991 C10_P_btm.n3377 C10_P_btm.n3376 0.6255
R34992 C10_P_btm.n3380 C10_P_btm.n3379 0.6255
R34993 C10_P_btm.n3383 C10_P_btm.n3382 0.6255
R34994 C10_P_btm.n3386 C10_P_btm.n3385 0.6255
R34995 C10_P_btm.n3389 C10_P_btm.n3388 0.6255
R34996 C10_P_btm.n3392 C10_P_btm.n3391 0.6255
R34997 C10_P_btm.n3395 C10_P_btm.n3394 0.6255
R34998 C10_P_btm.n3405 C10_P_btm.n3404 0.6255
R34999 C10_P_btm.n3408 C10_P_btm.n3407 0.6255
R35000 C10_P_btm.n3411 C10_P_btm.n3410 0.6255
R35001 C10_P_btm.n3414 C10_P_btm.n3413 0.6255
R35002 C10_P_btm.n3417 C10_P_btm.n3416 0.6255
R35003 C10_P_btm.n3420 C10_P_btm.n3419 0.6255
R35004 C10_P_btm.n3423 C10_P_btm.n3422 0.6255
R35005 C10_P_btm.n3426 C10_P_btm.n3425 0.6255
R35006 C10_P_btm.n312 C10_P_btm.n294 0.6255
R35007 C10_P_btm.n315 C10_P_btm.n314 0.6255
R35008 C10_P_btm.n318 C10_P_btm.n317 0.6255
R35009 C10_P_btm.n321 C10_P_btm.n320 0.6255
R35010 C10_P_btm.n324 C10_P_btm.n323 0.6255
R35011 C10_P_btm.n327 C10_P_btm.n326 0.6255
R35012 C10_P_btm.n330 C10_P_btm.n329 0.6255
R35013 C10_P_btm.n334 C10_P_btm.n332 0.6255
R35014 C10_P_btm.n3462 C10_P_btm.n3461 0.6255
R35015 C10_P_btm.n3459 C10_P_btm.n3458 0.6255
R35016 C10_P_btm.n3456 C10_P_btm.n3455 0.6255
R35017 C10_P_btm.n3453 C10_P_btm.n3452 0.6255
R35018 C10_P_btm.n3450 C10_P_btm.n3449 0.6255
R35019 C10_P_btm.n3447 C10_P_btm.n3446 0.6255
R35020 C10_P_btm.n3444 C10_P_btm.n3443 0.6255
R35021 C10_P_btm.n3441 C10_P_btm.n3440 0.6255
R35022 C10_P_btm.n3493 C10_P_btm.n3492 0.6255
R35023 C10_P_btm.n3490 C10_P_btm.n3489 0.6255
R35024 C10_P_btm.n3487 C10_P_btm.n3486 0.6255
R35025 C10_P_btm.n3484 C10_P_btm.n3483 0.6255
R35026 C10_P_btm.n3481 C10_P_btm.n3480 0.6255
R35027 C10_P_btm.n3478 C10_P_btm.n3477 0.6255
R35028 C10_P_btm.n3475 C10_P_btm.n3474 0.6255
R35029 C10_P_btm.n3472 C10_P_btm.n3471 0.6255
R35030 C10_P_btm.n281 C10_P_btm.n279 0.6255
R35031 C10_P_btm.n277 C10_P_btm.n276 0.6255
R35032 C10_P_btm.n274 C10_P_btm.n273 0.6255
R35033 C10_P_btm.n271 C10_P_btm.n270 0.6255
R35034 C10_P_btm.n268 C10_P_btm.n267 0.6255
R35035 C10_P_btm.n265 C10_P_btm.n264 0.6255
R35036 C10_P_btm.n262 C10_P_btm.n261 0.6255
R35037 C10_P_btm.n259 C10_P_btm.n241 0.6255
R35038 C10_P_btm.n3508 C10_P_btm.n3507 0.6255
R35039 C10_P_btm.n3511 C10_P_btm.n3510 0.6255
R35040 C10_P_btm.n3514 C10_P_btm.n3513 0.6255
R35041 C10_P_btm.n3517 C10_P_btm.n3516 0.6255
R35042 C10_P_btm.n3520 C10_P_btm.n3519 0.6255
R35043 C10_P_btm.n3523 C10_P_btm.n3522 0.6255
R35044 C10_P_btm.n3526 C10_P_btm.n3525 0.6255
R35045 C10_P_btm.n3529 C10_P_btm.n3528 0.6255
R35046 C10_P_btm.n3539 C10_P_btm.n3538 0.6255
R35047 C10_P_btm.n3542 C10_P_btm.n3541 0.6255
R35048 C10_P_btm.n3545 C10_P_btm.n3544 0.6255
R35049 C10_P_btm.n3548 C10_P_btm.n3547 0.6255
R35050 C10_P_btm.n3551 C10_P_btm.n3550 0.6255
R35051 C10_P_btm.n3554 C10_P_btm.n3553 0.6255
R35052 C10_P_btm.n3557 C10_P_btm.n3556 0.6255
R35053 C10_P_btm.n3560 C10_P_btm.n3559 0.6255
R35054 C10_P_btm.n206 C10_P_btm.n188 0.6255
R35055 C10_P_btm.n209 C10_P_btm.n208 0.6255
R35056 C10_P_btm.n212 C10_P_btm.n211 0.6255
R35057 C10_P_btm.n215 C10_P_btm.n214 0.6255
R35058 C10_P_btm.n218 C10_P_btm.n217 0.6255
R35059 C10_P_btm.n221 C10_P_btm.n220 0.6255
R35060 C10_P_btm.n224 C10_P_btm.n223 0.6255
R35061 C10_P_btm.n228 C10_P_btm.n226 0.6255
R35062 C10_P_btm.n3596 C10_P_btm.n3595 0.6255
R35063 C10_P_btm.n3593 C10_P_btm.n3592 0.6255
R35064 C10_P_btm.n3590 C10_P_btm.n3589 0.6255
R35065 C10_P_btm.n3587 C10_P_btm.n3586 0.6255
R35066 C10_P_btm.n3584 C10_P_btm.n3583 0.6255
R35067 C10_P_btm.n3581 C10_P_btm.n3580 0.6255
R35068 C10_P_btm.n3578 C10_P_btm.n3577 0.6255
R35069 C10_P_btm.n3575 C10_P_btm.n3574 0.6255
R35070 C10_P_btm.n3627 C10_P_btm.n3626 0.6255
R35071 C10_P_btm.n3624 C10_P_btm.n3623 0.6255
R35072 C10_P_btm.n3621 C10_P_btm.n3620 0.6255
R35073 C10_P_btm.n3618 C10_P_btm.n3617 0.6255
R35074 C10_P_btm.n3615 C10_P_btm.n3614 0.6255
R35075 C10_P_btm.n3612 C10_P_btm.n3611 0.6255
R35076 C10_P_btm.n3609 C10_P_btm.n3608 0.6255
R35077 C10_P_btm.n3606 C10_P_btm.n3605 0.6255
R35078 C10_P_btm.n175 C10_P_btm.n173 0.6255
R35079 C10_P_btm.n171 C10_P_btm.n170 0.6255
R35080 C10_P_btm.n168 C10_P_btm.n167 0.6255
R35081 C10_P_btm.n165 C10_P_btm.n164 0.6255
R35082 C10_P_btm.n162 C10_P_btm.n161 0.6255
R35083 C10_P_btm.n159 C10_P_btm.n158 0.6255
R35084 C10_P_btm.n156 C10_P_btm.n155 0.6255
R35085 C10_P_btm.n153 C10_P_btm.n135 0.6255
R35086 C10_P_btm.n3642 C10_P_btm.n3641 0.6255
R35087 C10_P_btm.n3645 C10_P_btm.n3644 0.6255
R35088 C10_P_btm.n3648 C10_P_btm.n3647 0.6255
R35089 C10_P_btm.n3651 C10_P_btm.n3650 0.6255
R35090 C10_P_btm.n3654 C10_P_btm.n3653 0.6255
R35091 C10_P_btm.n3657 C10_P_btm.n3656 0.6255
R35092 C10_P_btm.n3660 C10_P_btm.n3659 0.6255
R35093 C10_P_btm.n3663 C10_P_btm.n3662 0.6255
R35094 C10_P_btm.n3673 C10_P_btm.n3672 0.6255
R35095 C10_P_btm.n3676 C10_P_btm.n3675 0.6255
R35096 C10_P_btm.n3679 C10_P_btm.n3678 0.6255
R35097 C10_P_btm.n3682 C10_P_btm.n3681 0.6255
R35098 C10_P_btm.n3685 C10_P_btm.n3684 0.6255
R35099 C10_P_btm.n3688 C10_P_btm.n3687 0.6255
R35100 C10_P_btm.n3691 C10_P_btm.n3690 0.6255
R35101 C10_P_btm.n3694 C10_P_btm.n3693 0.6255
R35102 C10_P_btm.n100 C10_P_btm.n82 0.6255
R35103 C10_P_btm.n103 C10_P_btm.n102 0.6255
R35104 C10_P_btm.n106 C10_P_btm.n105 0.6255
R35105 C10_P_btm.n109 C10_P_btm.n108 0.6255
R35106 C10_P_btm.n112 C10_P_btm.n111 0.6255
R35107 C10_P_btm.n115 C10_P_btm.n114 0.6255
R35108 C10_P_btm.n118 C10_P_btm.n117 0.6255
R35109 C10_P_btm.n122 C10_P_btm.n120 0.6255
R35110 C10_P_btm.n3730 C10_P_btm.n3729 0.6255
R35111 C10_P_btm.n3727 C10_P_btm.n3726 0.6255
R35112 C10_P_btm.n3724 C10_P_btm.n3723 0.6255
R35113 C10_P_btm.n3721 C10_P_btm.n3720 0.6255
R35114 C10_P_btm.n3718 C10_P_btm.n3717 0.6255
R35115 C10_P_btm.n3715 C10_P_btm.n3714 0.6255
R35116 C10_P_btm.n3712 C10_P_btm.n3711 0.6255
R35117 C10_P_btm.n3709 C10_P_btm.n3708 0.6255
R35118 C10_P_btm.n3796 C10_P_btm.n3795 0.6255
R35119 C10_P_btm.n3793 C10_P_btm.n3792 0.6255
R35120 C10_P_btm.n3790 C10_P_btm.n3789 0.6255
R35121 C10_P_btm.n3787 C10_P_btm.n3786 0.6255
R35122 C10_P_btm.n3784 C10_P_btm.n3783 0.6255
R35123 C10_P_btm.n3781 C10_P_btm.n3780 0.6255
R35124 C10_P_btm.n3778 C10_P_btm.n3777 0.6255
R35125 C10_P_btm.n3775 C10_P_btm.n3774 0.6255
R35126 C10_P_btm.n3765 C10_P_btm.n3764 0.6255
R35127 C10_P_btm.n3762 C10_P_btm.n3761 0.6255
R35128 C10_P_btm.n3759 C10_P_btm.n3758 0.6255
R35129 C10_P_btm.n3756 C10_P_btm.n3755 0.6255
R35130 C10_P_btm.n3753 C10_P_btm.n3752 0.6255
R35131 C10_P_btm.n3750 C10_P_btm.n3749 0.6255
R35132 C10_P_btm.n3747 C10_P_btm.n3746 0.6255
R35133 C10_P_btm.n3744 C10_P_btm.n62 0.6255
R35134 C10_P_btm.n3811 C10_P_btm.n3810 0.6255
R35135 C10_P_btm.n3814 C10_P_btm.n3813 0.6255
R35136 C10_P_btm.n3817 C10_P_btm.n3816 0.6255
R35137 C10_P_btm.n3820 C10_P_btm.n3819 0.6255
R35138 C10_P_btm.n3823 C10_P_btm.n3822 0.6255
R35139 C10_P_btm.n3826 C10_P_btm.n3825 0.6255
R35140 C10_P_btm.n3829 C10_P_btm.n3828 0.6255
R35141 C10_P_btm.n3833 C10_P_btm.n3831 0.6255
R35142 C10_P_btm.n3840 C10_P_btm.n3839 0.6255
R35143 C10_P_btm.n3843 C10_P_btm.n3842 0.6255
R35144 C10_P_btm.n3846 C10_P_btm.n3845 0.6255
R35145 C10_P_btm.n3849 C10_P_btm.n3848 0.6255
R35146 C10_P_btm.n3852 C10_P_btm.n3851 0.6255
R35147 C10_P_btm.n3855 C10_P_btm.n3854 0.6255
R35148 C10_P_btm.n3858 C10_P_btm.n3857 0.6255
R35149 C10_P_btm.n3861 C10_P_btm.n3860 0.6255
R35150 C10_P_btm.n3871 C10_P_btm.n3870 0.6255
R35151 C10_P_btm.n3874 C10_P_btm.n3873 0.6255
R35152 C10_P_btm.n3877 C10_P_btm.n3876 0.6255
R35153 C10_P_btm.n3880 C10_P_btm.n3879 0.6255
R35154 C10_P_btm.n3883 C10_P_btm.n3882 0.6255
R35155 C10_P_btm.n3886 C10_P_btm.n3885 0.6255
R35156 C10_P_btm.n3889 C10_P_btm.n3888 0.6255
R35157 C10_P_btm.n3892 C10_P_btm.n3891 0.6255
R35158 C10_P_btm.n19 C10_P_btm.n17 0.5005
R35159 C10_P_btm.n30 C10_P_btm.n28 0.5005
R35160 C10_P_btm.n31 C10_P_btm.n30 0.484875
R35161 C10_P_btm.n21 C10_P_btm.n19 0.453625
R35162 C10_P_btm.n472 C10_P_btm.n434 0.109875
R35163 C10_P_btm.n470 C10_P_btm.n434 0.109875
R35164 C10_P_btm.n475 C10_P_btm.n433 0.109875
R35165 C10_P_btm.n473 C10_P_btm.n433 0.109875
R35166 C10_P_btm.n478 C10_P_btm.n432 0.109875
R35167 C10_P_btm.n476 C10_P_btm.n432 0.109875
R35168 C10_P_btm.n481 C10_P_btm.n431 0.109875
R35169 C10_P_btm.n479 C10_P_btm.n431 0.109875
R35170 C10_P_btm.n484 C10_P_btm.n430 0.109875
R35171 C10_P_btm.n482 C10_P_btm.n430 0.109875
R35172 C10_P_btm.n487 C10_P_btm.n429 0.109875
R35173 C10_P_btm.n485 C10_P_btm.n429 0.109875
R35174 C10_P_btm.n490 C10_P_btm.n428 0.109875
R35175 C10_P_btm.n488 C10_P_btm.n428 0.109875
R35176 C10_P_btm.n493 C10_P_btm.n427 0.109875
R35177 C10_P_btm.n491 C10_P_btm.n427 0.109875
R35178 C10_P_btm.n496 C10_P_btm.n426 0.109875
R35179 C10_P_btm.n494 C10_P_btm.n426 0.109875
R35180 C10_P_btm.n499 C10_P_btm.n425 0.109875
R35181 C10_P_btm.n497 C10_P_btm.n425 0.109875
R35182 C10_P_btm.n502 C10_P_btm.n424 0.109875
R35183 C10_P_btm.n500 C10_P_btm.n424 0.109875
R35184 C10_P_btm.n505 C10_P_btm.n423 0.109875
R35185 C10_P_btm.n503 C10_P_btm.n423 0.109875
R35186 C10_P_btm.n2460 C10_P_btm.n2455 0.109875
R35187 C10_P_btm.n2460 C10_P_btm.n2459 0.109875
R35188 C10_P_btm.n2452 C10_P_btm.n2422 0.109875
R35189 C10_P_btm.n2454 C10_P_btm.n2422 0.109875
R35190 C10_P_btm.n2449 C10_P_btm.n2423 0.109875
R35191 C10_P_btm.n2451 C10_P_btm.n2423 0.109875
R35192 C10_P_btm.n2446 C10_P_btm.n2424 0.109875
R35193 C10_P_btm.n2448 C10_P_btm.n2424 0.109875
R35194 C10_P_btm.n2443 C10_P_btm.n2425 0.109875
R35195 C10_P_btm.n2445 C10_P_btm.n2425 0.109875
R35196 C10_P_btm.n2440 C10_P_btm.n2426 0.109875
R35197 C10_P_btm.n2442 C10_P_btm.n2426 0.109875
R35198 C10_P_btm.n2437 C10_P_btm.n2427 0.109875
R35199 C10_P_btm.n2439 C10_P_btm.n2427 0.109875
R35200 C10_P_btm.n2434 C10_P_btm.n2428 0.109875
R35201 C10_P_btm.n2436 C10_P_btm.n2428 0.109875
R35202 C10_P_btm.n2431 C10_P_btm.n2429 0.109875
R35203 C10_P_btm.n2433 C10_P_btm.n2429 0.109875
R35204 C10_P_btm.n2489 C10_P_btm.n2414 0.109875
R35205 C10_P_btm.n2487 C10_P_btm.n2414 0.109875
R35206 C10_P_btm.n2486 C10_P_btm.n2415 0.109875
R35207 C10_P_btm.n2484 C10_P_btm.n2415 0.109875
R35208 C10_P_btm.n2483 C10_P_btm.n2416 0.109875
R35209 C10_P_btm.n2481 C10_P_btm.n2416 0.109875
R35210 C10_P_btm.n2480 C10_P_btm.n2417 0.109875
R35211 C10_P_btm.n2478 C10_P_btm.n2417 0.109875
R35212 C10_P_btm.n2477 C10_P_btm.n2418 0.109875
R35213 C10_P_btm.n2475 C10_P_btm.n2418 0.109875
R35214 C10_P_btm.n2474 C10_P_btm.n2419 0.109875
R35215 C10_P_btm.n2472 C10_P_btm.n2419 0.109875
R35216 C10_P_btm.n2471 C10_P_btm.n2420 0.109875
R35217 C10_P_btm.n2469 C10_P_btm.n2420 0.109875
R35218 C10_P_btm.n2468 C10_P_btm.n2421 0.109875
R35219 C10_P_btm.n2466 C10_P_btm.n2421 0.109875
R35220 C10_P_btm.n2465 C10_P_btm.n2461 0.109875
R35221 C10_P_btm.n2463 C10_P_btm.n2461 0.109875
R35222 C10_P_btm.n2518 C10_P_btm.n2369 0.109875
R35223 C10_P_btm.n2520 C10_P_btm.n2369 0.109875
R35224 C10_P_btm.n2515 C10_P_btm.n2372 0.109875
R35225 C10_P_btm.n2517 C10_P_btm.n2372 0.109875
R35226 C10_P_btm.n2512 C10_P_btm.n2373 0.109875
R35227 C10_P_btm.n2514 C10_P_btm.n2373 0.109875
R35228 C10_P_btm.n2509 C10_P_btm.n2374 0.109875
R35229 C10_P_btm.n2511 C10_P_btm.n2374 0.109875
R35230 C10_P_btm.n2506 C10_P_btm.n2375 0.109875
R35231 C10_P_btm.n2508 C10_P_btm.n2375 0.109875
R35232 C10_P_btm.n2503 C10_P_btm.n2376 0.109875
R35233 C10_P_btm.n2505 C10_P_btm.n2376 0.109875
R35234 C10_P_btm.n2500 C10_P_btm.n2377 0.109875
R35235 C10_P_btm.n2502 C10_P_btm.n2377 0.109875
R35236 C10_P_btm.n2497 C10_P_btm.n2378 0.109875
R35237 C10_P_btm.n2499 C10_P_btm.n2378 0.109875
R35238 C10_P_btm.n2494 C10_P_btm.n2412 0.109875
R35239 C10_P_btm.n2496 C10_P_btm.n2412 0.109875
R35240 C10_P_btm.n2411 C10_P_btm.n2380 0.109875
R35241 C10_P_btm.n2411 C10_P_btm.n2410 0.109875
R35242 C10_P_btm.n2408 C10_P_btm.n2381 0.109875
R35243 C10_P_btm.n2406 C10_P_btm.n2381 0.109875
R35244 C10_P_btm.n2405 C10_P_btm.n2382 0.109875
R35245 C10_P_btm.n2403 C10_P_btm.n2382 0.109875
R35246 C10_P_btm.n2402 C10_P_btm.n2383 0.109875
R35247 C10_P_btm.n2400 C10_P_btm.n2383 0.109875
R35248 C10_P_btm.n2399 C10_P_btm.n2384 0.109875
R35249 C10_P_btm.n2397 C10_P_btm.n2384 0.109875
R35250 C10_P_btm.n2396 C10_P_btm.n2385 0.109875
R35251 C10_P_btm.n2394 C10_P_btm.n2385 0.109875
R35252 C10_P_btm.n2393 C10_P_btm.n2386 0.109875
R35253 C10_P_btm.n2391 C10_P_btm.n2386 0.109875
R35254 C10_P_btm.n2390 C10_P_btm.n2387 0.109875
R35255 C10_P_btm.n2388 C10_P_btm.n2387 0.109875
R35256 C10_P_btm.n2527 C10_P_btm.n2370 0.109875
R35257 C10_P_btm.n2527 C10_P_btm.n2526 0.109875
R35258 C10_P_btm.n2532 C10_P_btm.n2528 0.109875
R35259 C10_P_btm.n2530 C10_P_btm.n2528 0.109875
R35260 C10_P_btm.n2535 C10_P_btm.n2368 0.109875
R35261 C10_P_btm.n2533 C10_P_btm.n2368 0.109875
R35262 C10_P_btm.n2538 C10_P_btm.n2367 0.109875
R35263 C10_P_btm.n2536 C10_P_btm.n2367 0.109875
R35264 C10_P_btm.n2541 C10_P_btm.n2366 0.109875
R35265 C10_P_btm.n2539 C10_P_btm.n2366 0.109875
R35266 C10_P_btm.n2544 C10_P_btm.n2365 0.109875
R35267 C10_P_btm.n2542 C10_P_btm.n2365 0.109875
R35268 C10_P_btm.n2547 C10_P_btm.n2364 0.109875
R35269 C10_P_btm.n2545 C10_P_btm.n2364 0.109875
R35270 C10_P_btm.n2550 C10_P_btm.n2363 0.109875
R35271 C10_P_btm.n2548 C10_P_btm.n2363 0.109875
R35272 C10_P_btm.n2553 C10_P_btm.n2362 0.109875
R35273 C10_P_btm.n2551 C10_P_btm.n2362 0.109875
R35274 C10_P_btm.n2556 C10_P_btm.n2361 0.109875
R35275 C10_P_btm.n2554 C10_P_btm.n2361 0.109875
R35276 C10_P_btm.n2561 C10_P_btm.n2359 0.109875
R35277 C10_P_btm.n2563 C10_P_btm.n2359 0.109875
R35278 C10_P_btm.n2564 C10_P_btm.n2325 0.109875
R35279 C10_P_btm.n2566 C10_P_btm.n2325 0.109875
R35280 C10_P_btm.n2567 C10_P_btm.n2324 0.109875
R35281 C10_P_btm.n2569 C10_P_btm.n2324 0.109875
R35282 C10_P_btm.n2570 C10_P_btm.n2323 0.109875
R35283 C10_P_btm.n2572 C10_P_btm.n2323 0.109875
R35284 C10_P_btm.n2573 C10_P_btm.n2322 0.109875
R35285 C10_P_btm.n2575 C10_P_btm.n2322 0.109875
R35286 C10_P_btm.n2576 C10_P_btm.n2321 0.109875
R35287 C10_P_btm.n2578 C10_P_btm.n2321 0.109875
R35288 C10_P_btm.n2579 C10_P_btm.n2320 0.109875
R35289 C10_P_btm.n2581 C10_P_btm.n2320 0.109875
R35290 C10_P_btm.n2582 C10_P_btm.n2319 0.109875
R35291 C10_P_btm.n2584 C10_P_btm.n2319 0.109875
R35292 C10_P_btm.n2585 C10_P_btm.n2316 0.109875
R35293 C10_P_btm.n2587 C10_P_btm.n2316 0.109875
R35294 C10_P_btm.n2594 C10_P_btm.n2317 0.109875
R35295 C10_P_btm.n2594 C10_P_btm.n2593 0.109875
R35296 C10_P_btm.n2337 C10_P_btm.n2334 0.109875
R35297 C10_P_btm.n2335 C10_P_btm.n2334 0.109875
R35298 C10_P_btm.n2340 C10_P_btm.n2333 0.109875
R35299 C10_P_btm.n2338 C10_P_btm.n2333 0.109875
R35300 C10_P_btm.n2343 C10_P_btm.n2332 0.109875
R35301 C10_P_btm.n2341 C10_P_btm.n2332 0.109875
R35302 C10_P_btm.n2346 C10_P_btm.n2331 0.109875
R35303 C10_P_btm.n2344 C10_P_btm.n2331 0.109875
R35304 C10_P_btm.n2349 C10_P_btm.n2330 0.109875
R35305 C10_P_btm.n2347 C10_P_btm.n2330 0.109875
R35306 C10_P_btm.n2352 C10_P_btm.n2329 0.109875
R35307 C10_P_btm.n2350 C10_P_btm.n2329 0.109875
R35308 C10_P_btm.n2355 C10_P_btm.n2328 0.109875
R35309 C10_P_btm.n2353 C10_P_btm.n2328 0.109875
R35310 C10_P_btm.n2358 C10_P_btm.n2327 0.109875
R35311 C10_P_btm.n2358 C10_P_btm.n2357 0.109875
R35312 C10_P_btm.n2623 C10_P_btm.n2308 0.109875
R35313 C10_P_btm.n2621 C10_P_btm.n2308 0.109875
R35314 C10_P_btm.n2620 C10_P_btm.n2309 0.109875
R35315 C10_P_btm.n2618 C10_P_btm.n2309 0.109875
R35316 C10_P_btm.n2617 C10_P_btm.n2310 0.109875
R35317 C10_P_btm.n2615 C10_P_btm.n2310 0.109875
R35318 C10_P_btm.n2614 C10_P_btm.n2311 0.109875
R35319 C10_P_btm.n2612 C10_P_btm.n2311 0.109875
R35320 C10_P_btm.n2611 C10_P_btm.n2312 0.109875
R35321 C10_P_btm.n2609 C10_P_btm.n2312 0.109875
R35322 C10_P_btm.n2608 C10_P_btm.n2313 0.109875
R35323 C10_P_btm.n2606 C10_P_btm.n2313 0.109875
R35324 C10_P_btm.n2605 C10_P_btm.n2314 0.109875
R35325 C10_P_btm.n2603 C10_P_btm.n2314 0.109875
R35326 C10_P_btm.n2602 C10_P_btm.n2315 0.109875
R35327 C10_P_btm.n2600 C10_P_btm.n2315 0.109875
R35328 C10_P_btm.n2599 C10_P_btm.n2595 0.109875
R35329 C10_P_btm.n2597 C10_P_btm.n2595 0.109875
R35330 C10_P_btm.n2652 C10_P_btm.n2263 0.109875
R35331 C10_P_btm.n2654 C10_P_btm.n2263 0.109875
R35332 C10_P_btm.n2649 C10_P_btm.n2266 0.109875
R35333 C10_P_btm.n2651 C10_P_btm.n2266 0.109875
R35334 C10_P_btm.n2646 C10_P_btm.n2267 0.109875
R35335 C10_P_btm.n2648 C10_P_btm.n2267 0.109875
R35336 C10_P_btm.n2643 C10_P_btm.n2268 0.109875
R35337 C10_P_btm.n2645 C10_P_btm.n2268 0.109875
R35338 C10_P_btm.n2640 C10_P_btm.n2269 0.109875
R35339 C10_P_btm.n2642 C10_P_btm.n2269 0.109875
R35340 C10_P_btm.n2637 C10_P_btm.n2270 0.109875
R35341 C10_P_btm.n2639 C10_P_btm.n2270 0.109875
R35342 C10_P_btm.n2634 C10_P_btm.n2271 0.109875
R35343 C10_P_btm.n2636 C10_P_btm.n2271 0.109875
R35344 C10_P_btm.n2631 C10_P_btm.n2272 0.109875
R35345 C10_P_btm.n2633 C10_P_btm.n2272 0.109875
R35346 C10_P_btm.n2628 C10_P_btm.n2306 0.109875
R35347 C10_P_btm.n2630 C10_P_btm.n2306 0.109875
R35348 C10_P_btm.n2305 C10_P_btm.n2274 0.109875
R35349 C10_P_btm.n2305 C10_P_btm.n2304 0.109875
R35350 C10_P_btm.n2302 C10_P_btm.n2275 0.109875
R35351 C10_P_btm.n2300 C10_P_btm.n2275 0.109875
R35352 C10_P_btm.n2299 C10_P_btm.n2276 0.109875
R35353 C10_P_btm.n2297 C10_P_btm.n2276 0.109875
R35354 C10_P_btm.n2296 C10_P_btm.n2277 0.109875
R35355 C10_P_btm.n2294 C10_P_btm.n2277 0.109875
R35356 C10_P_btm.n2293 C10_P_btm.n2278 0.109875
R35357 C10_P_btm.n2291 C10_P_btm.n2278 0.109875
R35358 C10_P_btm.n2290 C10_P_btm.n2279 0.109875
R35359 C10_P_btm.n2288 C10_P_btm.n2279 0.109875
R35360 C10_P_btm.n2287 C10_P_btm.n2280 0.109875
R35361 C10_P_btm.n2285 C10_P_btm.n2280 0.109875
R35362 C10_P_btm.n2284 C10_P_btm.n2281 0.109875
R35363 C10_P_btm.n2282 C10_P_btm.n2281 0.109875
R35364 C10_P_btm.n2661 C10_P_btm.n2264 0.109875
R35365 C10_P_btm.n2661 C10_P_btm.n2660 0.109875
R35366 C10_P_btm.n2666 C10_P_btm.n2662 0.109875
R35367 C10_P_btm.n2664 C10_P_btm.n2662 0.109875
R35368 C10_P_btm.n2669 C10_P_btm.n2262 0.109875
R35369 C10_P_btm.n2667 C10_P_btm.n2262 0.109875
R35370 C10_P_btm.n2672 C10_P_btm.n2261 0.109875
R35371 C10_P_btm.n2670 C10_P_btm.n2261 0.109875
R35372 C10_P_btm.n2675 C10_P_btm.n2260 0.109875
R35373 C10_P_btm.n2673 C10_P_btm.n2260 0.109875
R35374 C10_P_btm.n2678 C10_P_btm.n2259 0.109875
R35375 C10_P_btm.n2676 C10_P_btm.n2259 0.109875
R35376 C10_P_btm.n2681 C10_P_btm.n2258 0.109875
R35377 C10_P_btm.n2679 C10_P_btm.n2258 0.109875
R35378 C10_P_btm.n2684 C10_P_btm.n2257 0.109875
R35379 C10_P_btm.n2682 C10_P_btm.n2257 0.109875
R35380 C10_P_btm.n2687 C10_P_btm.n2256 0.109875
R35381 C10_P_btm.n2685 C10_P_btm.n2256 0.109875
R35382 C10_P_btm.n2690 C10_P_btm.n2255 0.109875
R35383 C10_P_btm.n2688 C10_P_btm.n2255 0.109875
R35384 C10_P_btm.n2695 C10_P_btm.n2253 0.109875
R35385 C10_P_btm.n2697 C10_P_btm.n2253 0.109875
R35386 C10_P_btm.n2698 C10_P_btm.n2219 0.109875
R35387 C10_P_btm.n2700 C10_P_btm.n2219 0.109875
R35388 C10_P_btm.n2701 C10_P_btm.n2218 0.109875
R35389 C10_P_btm.n2703 C10_P_btm.n2218 0.109875
R35390 C10_P_btm.n2704 C10_P_btm.n2217 0.109875
R35391 C10_P_btm.n2706 C10_P_btm.n2217 0.109875
R35392 C10_P_btm.n2707 C10_P_btm.n2216 0.109875
R35393 C10_P_btm.n2709 C10_P_btm.n2216 0.109875
R35394 C10_P_btm.n2710 C10_P_btm.n2215 0.109875
R35395 C10_P_btm.n2712 C10_P_btm.n2215 0.109875
R35396 C10_P_btm.n2713 C10_P_btm.n2214 0.109875
R35397 C10_P_btm.n2715 C10_P_btm.n2214 0.109875
R35398 C10_P_btm.n2716 C10_P_btm.n2213 0.109875
R35399 C10_P_btm.n2718 C10_P_btm.n2213 0.109875
R35400 C10_P_btm.n2719 C10_P_btm.n2210 0.109875
R35401 C10_P_btm.n2721 C10_P_btm.n2210 0.109875
R35402 C10_P_btm.n2728 C10_P_btm.n2211 0.109875
R35403 C10_P_btm.n2728 C10_P_btm.n2727 0.109875
R35404 C10_P_btm.n2231 C10_P_btm.n2228 0.109875
R35405 C10_P_btm.n2229 C10_P_btm.n2228 0.109875
R35406 C10_P_btm.n2234 C10_P_btm.n2227 0.109875
R35407 C10_P_btm.n2232 C10_P_btm.n2227 0.109875
R35408 C10_P_btm.n2237 C10_P_btm.n2226 0.109875
R35409 C10_P_btm.n2235 C10_P_btm.n2226 0.109875
R35410 C10_P_btm.n2240 C10_P_btm.n2225 0.109875
R35411 C10_P_btm.n2238 C10_P_btm.n2225 0.109875
R35412 C10_P_btm.n2243 C10_P_btm.n2224 0.109875
R35413 C10_P_btm.n2241 C10_P_btm.n2224 0.109875
R35414 C10_P_btm.n2246 C10_P_btm.n2223 0.109875
R35415 C10_P_btm.n2244 C10_P_btm.n2223 0.109875
R35416 C10_P_btm.n2249 C10_P_btm.n2222 0.109875
R35417 C10_P_btm.n2247 C10_P_btm.n2222 0.109875
R35418 C10_P_btm.n2252 C10_P_btm.n2221 0.109875
R35419 C10_P_btm.n2252 C10_P_btm.n2251 0.109875
R35420 C10_P_btm.n2757 C10_P_btm.n2202 0.109875
R35421 C10_P_btm.n2755 C10_P_btm.n2202 0.109875
R35422 C10_P_btm.n2754 C10_P_btm.n2203 0.109875
R35423 C10_P_btm.n2752 C10_P_btm.n2203 0.109875
R35424 C10_P_btm.n2751 C10_P_btm.n2204 0.109875
R35425 C10_P_btm.n2749 C10_P_btm.n2204 0.109875
R35426 C10_P_btm.n2748 C10_P_btm.n2205 0.109875
R35427 C10_P_btm.n2746 C10_P_btm.n2205 0.109875
R35428 C10_P_btm.n2745 C10_P_btm.n2206 0.109875
R35429 C10_P_btm.n2743 C10_P_btm.n2206 0.109875
R35430 C10_P_btm.n2742 C10_P_btm.n2207 0.109875
R35431 C10_P_btm.n2740 C10_P_btm.n2207 0.109875
R35432 C10_P_btm.n2739 C10_P_btm.n2208 0.109875
R35433 C10_P_btm.n2737 C10_P_btm.n2208 0.109875
R35434 C10_P_btm.n2736 C10_P_btm.n2209 0.109875
R35435 C10_P_btm.n2734 C10_P_btm.n2209 0.109875
R35436 C10_P_btm.n2733 C10_P_btm.n2729 0.109875
R35437 C10_P_btm.n2731 C10_P_btm.n2729 0.109875
R35438 C10_P_btm.n2786 C10_P_btm.n2157 0.109875
R35439 C10_P_btm.n2788 C10_P_btm.n2157 0.109875
R35440 C10_P_btm.n2783 C10_P_btm.n2160 0.109875
R35441 C10_P_btm.n2785 C10_P_btm.n2160 0.109875
R35442 C10_P_btm.n2780 C10_P_btm.n2161 0.109875
R35443 C10_P_btm.n2782 C10_P_btm.n2161 0.109875
R35444 C10_P_btm.n2777 C10_P_btm.n2162 0.109875
R35445 C10_P_btm.n2779 C10_P_btm.n2162 0.109875
R35446 C10_P_btm.n2774 C10_P_btm.n2163 0.109875
R35447 C10_P_btm.n2776 C10_P_btm.n2163 0.109875
R35448 C10_P_btm.n2771 C10_P_btm.n2164 0.109875
R35449 C10_P_btm.n2773 C10_P_btm.n2164 0.109875
R35450 C10_P_btm.n2768 C10_P_btm.n2165 0.109875
R35451 C10_P_btm.n2770 C10_P_btm.n2165 0.109875
R35452 C10_P_btm.n2765 C10_P_btm.n2166 0.109875
R35453 C10_P_btm.n2767 C10_P_btm.n2166 0.109875
R35454 C10_P_btm.n2762 C10_P_btm.n2200 0.109875
R35455 C10_P_btm.n2764 C10_P_btm.n2200 0.109875
R35456 C10_P_btm.n2199 C10_P_btm.n2168 0.109875
R35457 C10_P_btm.n2199 C10_P_btm.n2198 0.109875
R35458 C10_P_btm.n2196 C10_P_btm.n2169 0.109875
R35459 C10_P_btm.n2194 C10_P_btm.n2169 0.109875
R35460 C10_P_btm.n2193 C10_P_btm.n2170 0.109875
R35461 C10_P_btm.n2191 C10_P_btm.n2170 0.109875
R35462 C10_P_btm.n2190 C10_P_btm.n2171 0.109875
R35463 C10_P_btm.n2188 C10_P_btm.n2171 0.109875
R35464 C10_P_btm.n2187 C10_P_btm.n2172 0.109875
R35465 C10_P_btm.n2185 C10_P_btm.n2172 0.109875
R35466 C10_P_btm.n2184 C10_P_btm.n2173 0.109875
R35467 C10_P_btm.n2182 C10_P_btm.n2173 0.109875
R35468 C10_P_btm.n2181 C10_P_btm.n2174 0.109875
R35469 C10_P_btm.n2179 C10_P_btm.n2174 0.109875
R35470 C10_P_btm.n2178 C10_P_btm.n2175 0.109875
R35471 C10_P_btm.n2176 C10_P_btm.n2175 0.109875
R35472 C10_P_btm.n2795 C10_P_btm.n2158 0.109875
R35473 C10_P_btm.n2795 C10_P_btm.n2794 0.109875
R35474 C10_P_btm.n2800 C10_P_btm.n2796 0.109875
R35475 C10_P_btm.n2798 C10_P_btm.n2796 0.109875
R35476 C10_P_btm.n2803 C10_P_btm.n2156 0.109875
R35477 C10_P_btm.n2801 C10_P_btm.n2156 0.109875
R35478 C10_P_btm.n2806 C10_P_btm.n2155 0.109875
R35479 C10_P_btm.n2804 C10_P_btm.n2155 0.109875
R35480 C10_P_btm.n2809 C10_P_btm.n2154 0.109875
R35481 C10_P_btm.n2807 C10_P_btm.n2154 0.109875
R35482 C10_P_btm.n2812 C10_P_btm.n2153 0.109875
R35483 C10_P_btm.n2810 C10_P_btm.n2153 0.109875
R35484 C10_P_btm.n2815 C10_P_btm.n2152 0.109875
R35485 C10_P_btm.n2813 C10_P_btm.n2152 0.109875
R35486 C10_P_btm.n2818 C10_P_btm.n2151 0.109875
R35487 C10_P_btm.n2816 C10_P_btm.n2151 0.109875
R35488 C10_P_btm.n2821 C10_P_btm.n2150 0.109875
R35489 C10_P_btm.n2819 C10_P_btm.n2150 0.109875
R35490 C10_P_btm.n2824 C10_P_btm.n2149 0.109875
R35491 C10_P_btm.n2822 C10_P_btm.n2149 0.109875
R35492 C10_P_btm.n2829 C10_P_btm.n2147 0.109875
R35493 C10_P_btm.n2831 C10_P_btm.n2147 0.109875
R35494 C10_P_btm.n2832 C10_P_btm.n2113 0.109875
R35495 C10_P_btm.n2834 C10_P_btm.n2113 0.109875
R35496 C10_P_btm.n2835 C10_P_btm.n2112 0.109875
R35497 C10_P_btm.n2837 C10_P_btm.n2112 0.109875
R35498 C10_P_btm.n2838 C10_P_btm.n2111 0.109875
R35499 C10_P_btm.n2840 C10_P_btm.n2111 0.109875
R35500 C10_P_btm.n2841 C10_P_btm.n2110 0.109875
R35501 C10_P_btm.n2843 C10_P_btm.n2110 0.109875
R35502 C10_P_btm.n2844 C10_P_btm.n2109 0.109875
R35503 C10_P_btm.n2846 C10_P_btm.n2109 0.109875
R35504 C10_P_btm.n2847 C10_P_btm.n2108 0.109875
R35505 C10_P_btm.n2849 C10_P_btm.n2108 0.109875
R35506 C10_P_btm.n2850 C10_P_btm.n2107 0.109875
R35507 C10_P_btm.n2852 C10_P_btm.n2107 0.109875
R35508 C10_P_btm.n2853 C10_P_btm.n2104 0.109875
R35509 C10_P_btm.n2855 C10_P_btm.n2104 0.109875
R35510 C10_P_btm.n2862 C10_P_btm.n2105 0.109875
R35511 C10_P_btm.n2862 C10_P_btm.n2861 0.109875
R35512 C10_P_btm.n2125 C10_P_btm.n2122 0.109875
R35513 C10_P_btm.n2123 C10_P_btm.n2122 0.109875
R35514 C10_P_btm.n2128 C10_P_btm.n2121 0.109875
R35515 C10_P_btm.n2126 C10_P_btm.n2121 0.109875
R35516 C10_P_btm.n2131 C10_P_btm.n2120 0.109875
R35517 C10_P_btm.n2129 C10_P_btm.n2120 0.109875
R35518 C10_P_btm.n2134 C10_P_btm.n2119 0.109875
R35519 C10_P_btm.n2132 C10_P_btm.n2119 0.109875
R35520 C10_P_btm.n2137 C10_P_btm.n2118 0.109875
R35521 C10_P_btm.n2135 C10_P_btm.n2118 0.109875
R35522 C10_P_btm.n2140 C10_P_btm.n2117 0.109875
R35523 C10_P_btm.n2138 C10_P_btm.n2117 0.109875
R35524 C10_P_btm.n2143 C10_P_btm.n2116 0.109875
R35525 C10_P_btm.n2141 C10_P_btm.n2116 0.109875
R35526 C10_P_btm.n2146 C10_P_btm.n2115 0.109875
R35527 C10_P_btm.n2146 C10_P_btm.n2145 0.109875
R35528 C10_P_btm.n2891 C10_P_btm.n2096 0.109875
R35529 C10_P_btm.n2889 C10_P_btm.n2096 0.109875
R35530 C10_P_btm.n2888 C10_P_btm.n2097 0.109875
R35531 C10_P_btm.n2886 C10_P_btm.n2097 0.109875
R35532 C10_P_btm.n2885 C10_P_btm.n2098 0.109875
R35533 C10_P_btm.n2883 C10_P_btm.n2098 0.109875
R35534 C10_P_btm.n2882 C10_P_btm.n2099 0.109875
R35535 C10_P_btm.n2880 C10_P_btm.n2099 0.109875
R35536 C10_P_btm.n2879 C10_P_btm.n2100 0.109875
R35537 C10_P_btm.n2877 C10_P_btm.n2100 0.109875
R35538 C10_P_btm.n2876 C10_P_btm.n2101 0.109875
R35539 C10_P_btm.n2874 C10_P_btm.n2101 0.109875
R35540 C10_P_btm.n2873 C10_P_btm.n2102 0.109875
R35541 C10_P_btm.n2871 C10_P_btm.n2102 0.109875
R35542 C10_P_btm.n2870 C10_P_btm.n2103 0.109875
R35543 C10_P_btm.n2868 C10_P_btm.n2103 0.109875
R35544 C10_P_btm.n2867 C10_P_btm.n2863 0.109875
R35545 C10_P_btm.n2865 C10_P_btm.n2863 0.109875
R35546 C10_P_btm.n2955 C10_P_btm.n2084 0.109875
R35547 C10_P_btm.n2957 C10_P_btm.n2084 0.109875
R35548 C10_P_btm.n2952 C10_P_btm.n2087 0.109875
R35549 C10_P_btm.n2954 C10_P_btm.n2087 0.109875
R35550 C10_P_btm.n2949 C10_P_btm.n2088 0.109875
R35551 C10_P_btm.n2951 C10_P_btm.n2088 0.109875
R35552 C10_P_btm.n2946 C10_P_btm.n2089 0.109875
R35553 C10_P_btm.n2948 C10_P_btm.n2089 0.109875
R35554 C10_P_btm.n2943 C10_P_btm.n2090 0.109875
R35555 C10_P_btm.n2945 C10_P_btm.n2090 0.109875
R35556 C10_P_btm.n2940 C10_P_btm.n2091 0.109875
R35557 C10_P_btm.n2942 C10_P_btm.n2091 0.109875
R35558 C10_P_btm.n2937 C10_P_btm.n2092 0.109875
R35559 C10_P_btm.n2939 C10_P_btm.n2092 0.109875
R35560 C10_P_btm.n2934 C10_P_btm.n2093 0.109875
R35561 C10_P_btm.n2936 C10_P_btm.n2093 0.109875
R35562 C10_P_btm.n2931 C10_P_btm.n2094 0.109875
R35563 C10_P_btm.n2933 C10_P_btm.n2094 0.109875
R35564 C10_P_btm.n2926 C10_P_btm.n2075 0.109875
R35565 C10_P_btm.n2924 C10_P_btm.n2075 0.109875
R35566 C10_P_btm.n2923 C10_P_btm.n2896 0.109875
R35567 C10_P_btm.n2921 C10_P_btm.n2896 0.109875
R35568 C10_P_btm.n2920 C10_P_btm.n2897 0.109875
R35569 C10_P_btm.n2918 C10_P_btm.n2897 0.109875
R35570 C10_P_btm.n2917 C10_P_btm.n2898 0.109875
R35571 C10_P_btm.n2915 C10_P_btm.n2898 0.109875
R35572 C10_P_btm.n2914 C10_P_btm.n2899 0.109875
R35573 C10_P_btm.n2912 C10_P_btm.n2899 0.109875
R35574 C10_P_btm.n2911 C10_P_btm.n2900 0.109875
R35575 C10_P_btm.n2909 C10_P_btm.n2900 0.109875
R35576 C10_P_btm.n2908 C10_P_btm.n2901 0.109875
R35577 C10_P_btm.n2906 C10_P_btm.n2901 0.109875
R35578 C10_P_btm.n2905 C10_P_btm.n2902 0.109875
R35579 C10_P_btm.n2903 C10_P_btm.n2902 0.109875
R35580 C10_P_btm.n2964 C10_P_btm.n2085 0.109875
R35581 C10_P_btm.n2964 C10_P_btm.n2963 0.109875
R35582 C10_P_btm.n2969 C10_P_btm.n2965 0.109875
R35583 C10_P_btm.n2967 C10_P_btm.n2965 0.109875
R35584 C10_P_btm.n2972 C10_P_btm.n2083 0.109875
R35585 C10_P_btm.n2970 C10_P_btm.n2083 0.109875
R35586 C10_P_btm.n2975 C10_P_btm.n2082 0.109875
R35587 C10_P_btm.n2973 C10_P_btm.n2082 0.109875
R35588 C10_P_btm.n2978 C10_P_btm.n2081 0.109875
R35589 C10_P_btm.n2976 C10_P_btm.n2081 0.109875
R35590 C10_P_btm.n2981 C10_P_btm.n2080 0.109875
R35591 C10_P_btm.n2979 C10_P_btm.n2080 0.109875
R35592 C10_P_btm.n2984 C10_P_btm.n2079 0.109875
R35593 C10_P_btm.n2982 C10_P_btm.n2079 0.109875
R35594 C10_P_btm.n2987 C10_P_btm.n2078 0.109875
R35595 C10_P_btm.n2985 C10_P_btm.n2078 0.109875
R35596 C10_P_btm.n2990 C10_P_btm.n2077 0.109875
R35597 C10_P_btm.n2988 C10_P_btm.n2077 0.109875
R35598 C10_P_btm.n2993 C10_P_btm.n2076 0.109875
R35599 C10_P_btm.n2993 C10_P_btm.n2992 0.109875
R35600 C10_P_btm.n2996 C10_P_btm.n2994 0.109875
R35601 C10_P_btm.n2998 C10_P_btm.n2994 0.109875
R35602 C10_P_btm.n2999 C10_P_btm.n2074 0.109875
R35603 C10_P_btm.n3001 C10_P_btm.n2074 0.109875
R35604 C10_P_btm.n3002 C10_P_btm.n2073 0.109875
R35605 C10_P_btm.n3004 C10_P_btm.n2073 0.109875
R35606 C10_P_btm.n3005 C10_P_btm.n2072 0.109875
R35607 C10_P_btm.n3007 C10_P_btm.n2072 0.109875
R35608 C10_P_btm.n3008 C10_P_btm.n2071 0.109875
R35609 C10_P_btm.n3010 C10_P_btm.n2071 0.109875
R35610 C10_P_btm.n3011 C10_P_btm.n2070 0.109875
R35611 C10_P_btm.n3013 C10_P_btm.n2070 0.109875
R35612 C10_P_btm.n3014 C10_P_btm.n2069 0.109875
R35613 C10_P_btm.n3016 C10_P_btm.n2069 0.109875
R35614 C10_P_btm.n3017 C10_P_btm.n2068 0.109875
R35615 C10_P_btm.n3019 C10_P_btm.n2068 0.109875
R35616 C10_P_btm.n3020 C10_P_btm.n2067 0.109875
R35617 C10_P_btm.n3022 C10_P_btm.n2067 0.109875
R35618 C10_P_btm.n3041 C10_P_btm.n3037 0.109875
R35619 C10_P_btm.n3039 C10_P_btm.n3037 0.109875
R35620 C10_P_btm.n3044 C10_P_btm.n3036 0.109875
R35621 C10_P_btm.n3042 C10_P_btm.n3036 0.109875
R35622 C10_P_btm.n3047 C10_P_btm.n3035 0.109875
R35623 C10_P_btm.n3045 C10_P_btm.n3035 0.109875
R35624 C10_P_btm.n3050 C10_P_btm.n3034 0.109875
R35625 C10_P_btm.n3048 C10_P_btm.n3034 0.109875
R35626 C10_P_btm.n3053 C10_P_btm.n3033 0.109875
R35627 C10_P_btm.n3051 C10_P_btm.n3033 0.109875
R35628 C10_P_btm.n3056 C10_P_btm.n3032 0.109875
R35629 C10_P_btm.n3054 C10_P_btm.n3032 0.109875
R35630 C10_P_btm.n3059 C10_P_btm.n3031 0.109875
R35631 C10_P_btm.n3057 C10_P_btm.n3031 0.109875
R35632 C10_P_btm.n3062 C10_P_btm.n3030 0.109875
R35633 C10_P_btm.n3060 C10_P_btm.n3030 0.109875
R35634 C10_P_btm.n3065 C10_P_btm.n3029 0.109875
R35635 C10_P_btm.n3063 C10_P_btm.n3029 0.109875
R35636 C10_P_btm.n3068 C10_P_btm.n3028 0.109875
R35637 C10_P_btm.n3066 C10_P_btm.n3028 0.109875
R35638 C10_P_btm.n3071 C10_P_btm.n3027 0.109875
R35639 C10_P_btm.n3069 C10_P_btm.n3027 0.109875
R35640 C10_P_btm.n3074 C10_P_btm.n3026 0.109875
R35641 C10_P_btm.n3072 C10_P_btm.n3026 0.109875
R35642 C10_P_btm.n3077 C10_P_btm.n3025 0.109875
R35643 C10_P_btm.n3075 C10_P_btm.n3025 0.109875
R35644 C10_P_btm.n3080 C10_P_btm.n2065 0.109875
R35645 C10_P_btm.n3078 C10_P_btm.n2065 0.109875
R35646 C10_P_btm.n3083 C10_P_btm.n2064 0.109875
R35647 C10_P_btm.n3081 C10_P_btm.n2064 0.109875
R35648 C10_P_btm.n3086 C10_P_btm.n2063 0.109875
R35649 C10_P_btm.n3084 C10_P_btm.n2063 0.109875
R35650 C10_P_btm.n3089 C10_P_btm.n2062 0.109875
R35651 C10_P_btm.n3087 C10_P_btm.n2062 0.109875
R35652 C10_P_btm.n3092 C10_P_btm.n2061 0.109875
R35653 C10_P_btm.n3090 C10_P_btm.n2061 0.109875
R35654 C10_P_btm.n3095 C10_P_btm.n2060 0.109875
R35655 C10_P_btm.n3093 C10_P_btm.n2060 0.109875
R35656 C10_P_btm.n3098 C10_P_btm.n2059 0.109875
R35657 C10_P_btm.n3096 C10_P_btm.n2059 0.109875
R35658 C10_P_btm.n3101 C10_P_btm.n2058 0.109875
R35659 C10_P_btm.n3099 C10_P_btm.n2058 0.109875
R35660 C10_P_btm.n3104 C10_P_btm.n2057 0.109875
R35661 C10_P_btm.n3102 C10_P_btm.n2057 0.109875
R35662 C10_P_btm.n1289 C10_P_btm.n1287 0.109875
R35663 C10_P_btm.n1291 C10_P_btm.n1287 0.109875
R35664 C10_P_btm.n1292 C10_P_btm.n1041 0.109875
R35665 C10_P_btm.n1294 C10_P_btm.n1041 0.109875
R35666 C10_P_btm.n1295 C10_P_btm.n1040 0.109875
R35667 C10_P_btm.n1297 C10_P_btm.n1040 0.109875
R35668 C10_P_btm.n1298 C10_P_btm.n1039 0.109875
R35669 C10_P_btm.n1300 C10_P_btm.n1039 0.109875
R35670 C10_P_btm.n1301 C10_P_btm.n1038 0.109875
R35671 C10_P_btm.n1303 C10_P_btm.n1038 0.109875
R35672 C10_P_btm.n1304 C10_P_btm.n1037 0.109875
R35673 C10_P_btm.n1306 C10_P_btm.n1037 0.109875
R35674 C10_P_btm.n1307 C10_P_btm.n1036 0.109875
R35675 C10_P_btm.n1309 C10_P_btm.n1036 0.109875
R35676 C10_P_btm.n1310 C10_P_btm.n1035 0.109875
R35677 C10_P_btm.n1312 C10_P_btm.n1035 0.109875
R35678 C10_P_btm.n1313 C10_P_btm.n1034 0.109875
R35679 C10_P_btm.n1315 C10_P_btm.n1034 0.109875
R35680 C10_P_btm.n1316 C10_P_btm.n1033 0.109875
R35681 C10_P_btm.n1318 C10_P_btm.n1033 0.109875
R35682 C10_P_btm.n1319 C10_P_btm.n1032 0.109875
R35683 C10_P_btm.n1321 C10_P_btm.n1032 0.109875
R35684 C10_P_btm.n1322 C10_P_btm.n1031 0.109875
R35685 C10_P_btm.n1324 C10_P_btm.n1031 0.109875
R35686 C10_P_btm.n1325 C10_P_btm.n1030 0.109875
R35687 C10_P_btm.n1327 C10_P_btm.n1030 0.109875
R35688 C10_P_btm.n1328 C10_P_btm.n1029 0.109875
R35689 C10_P_btm.n1330 C10_P_btm.n1029 0.109875
R35690 C10_P_btm.n1331 C10_P_btm.n1028 0.109875
R35691 C10_P_btm.n1333 C10_P_btm.n1028 0.109875
R35692 C10_P_btm.n1334 C10_P_btm.n1027 0.109875
R35693 C10_P_btm.n1336 C10_P_btm.n1027 0.109875
R35694 C10_P_btm.n1337 C10_P_btm.n1026 0.109875
R35695 C10_P_btm.n1339 C10_P_btm.n1026 0.109875
R35696 C10_P_btm.n1340 C10_P_btm.n1025 0.109875
R35697 C10_P_btm.n1342 C10_P_btm.n1025 0.109875
R35698 C10_P_btm.n1343 C10_P_btm.n1024 0.109875
R35699 C10_P_btm.n1345 C10_P_btm.n1024 0.109875
R35700 C10_P_btm.n1346 C10_P_btm.n1023 0.109875
R35701 C10_P_btm.n1348 C10_P_btm.n1023 0.109875
R35702 C10_P_btm.n1349 C10_P_btm.n1022 0.109875
R35703 C10_P_btm.n1351 C10_P_btm.n1022 0.109875
R35704 C10_P_btm.n1352 C10_P_btm.n1021 0.109875
R35705 C10_P_btm.n1354 C10_P_btm.n1021 0.109875
R35706 C10_P_btm.n1355 C10_P_btm.n1020 0.109875
R35707 C10_P_btm.n1357 C10_P_btm.n1020 0.109875
R35708 C10_P_btm.n1358 C10_P_btm.n1019 0.109875
R35709 C10_P_btm.n1360 C10_P_btm.n1019 0.109875
R35710 C10_P_btm.n1361 C10_P_btm.n1018 0.109875
R35711 C10_P_btm.n1363 C10_P_btm.n1018 0.109875
R35712 C10_P_btm.n1364 C10_P_btm.n1017 0.109875
R35713 C10_P_btm.n1366 C10_P_btm.n1017 0.109875
R35714 C10_P_btm.n1367 C10_P_btm.n1016 0.109875
R35715 C10_P_btm.n1369 C10_P_btm.n1016 0.109875
R35716 C10_P_btm.n1370 C10_P_btm.n1015 0.109875
R35717 C10_P_btm.n1372 C10_P_btm.n1015 0.109875
R35718 C10_P_btm.n1373 C10_P_btm.n1014 0.109875
R35719 C10_P_btm.n1375 C10_P_btm.n1014 0.109875
R35720 C10_P_btm.n1376 C10_P_btm.n1013 0.109875
R35721 C10_P_btm.n1378 C10_P_btm.n1013 0.109875
R35722 C10_P_btm.n1379 C10_P_btm.n1012 0.109875
R35723 C10_P_btm.n1381 C10_P_btm.n1012 0.109875
R35724 C10_P_btm.n1382 C10_P_btm.n1011 0.109875
R35725 C10_P_btm.n1384 C10_P_btm.n1011 0.109875
R35726 C10_P_btm.n1385 C10_P_btm.n1010 0.109875
R35727 C10_P_btm.n1387 C10_P_btm.n1010 0.109875
R35728 C10_P_btm.n1388 C10_P_btm.n1009 0.109875
R35729 C10_P_btm.n1390 C10_P_btm.n1009 0.109875
R35730 C10_P_btm.n1391 C10_P_btm.n1008 0.109875
R35731 C10_P_btm.n1393 C10_P_btm.n1008 0.109875
R35732 C10_P_btm.n1394 C10_P_btm.n1007 0.109875
R35733 C10_P_btm.n1396 C10_P_btm.n1007 0.109875
R35734 C10_P_btm.n1397 C10_P_btm.n1006 0.109875
R35735 C10_P_btm.n1399 C10_P_btm.n1006 0.109875
R35736 C10_P_btm.n1400 C10_P_btm.n1005 0.109875
R35737 C10_P_btm.n1402 C10_P_btm.n1005 0.109875
R35738 C10_P_btm.n1403 C10_P_btm.n1004 0.109875
R35739 C10_P_btm.n1405 C10_P_btm.n1004 0.109875
R35740 C10_P_btm.n1406 C10_P_btm.n1003 0.109875
R35741 C10_P_btm.n1408 C10_P_btm.n1003 0.109875
R35742 C10_P_btm.n1409 C10_P_btm.n1002 0.109875
R35743 C10_P_btm.n1411 C10_P_btm.n1002 0.109875
R35744 C10_P_btm.n1412 C10_P_btm.n1001 0.109875
R35745 C10_P_btm.n1414 C10_P_btm.n1001 0.109875
R35746 C10_P_btm.n1415 C10_P_btm.n1000 0.109875
R35747 C10_P_btm.n1417 C10_P_btm.n1000 0.109875
R35748 C10_P_btm.n1418 C10_P_btm.n999 0.109875
R35749 C10_P_btm.n1420 C10_P_btm.n999 0.109875
R35750 C10_P_btm.n1421 C10_P_btm.n998 0.109875
R35751 C10_P_btm.n1423 C10_P_btm.n998 0.109875
R35752 C10_P_btm.n1424 C10_P_btm.n997 0.109875
R35753 C10_P_btm.n1426 C10_P_btm.n997 0.109875
R35754 C10_P_btm.n1427 C10_P_btm.n996 0.109875
R35755 C10_P_btm.n1429 C10_P_btm.n996 0.109875
R35756 C10_P_btm.n1430 C10_P_btm.n995 0.109875
R35757 C10_P_btm.n1432 C10_P_btm.n995 0.109875
R35758 C10_P_btm.n1433 C10_P_btm.n994 0.109875
R35759 C10_P_btm.n1435 C10_P_btm.n994 0.109875
R35760 C10_P_btm.n1436 C10_P_btm.n993 0.109875
R35761 C10_P_btm.n1438 C10_P_btm.n993 0.109875
R35762 C10_P_btm.n1439 C10_P_btm.n992 0.109875
R35763 C10_P_btm.n1441 C10_P_btm.n992 0.109875
R35764 C10_P_btm.n1442 C10_P_btm.n991 0.109875
R35765 C10_P_btm.n1444 C10_P_btm.n991 0.109875
R35766 C10_P_btm.n1445 C10_P_btm.n990 0.109875
R35767 C10_P_btm.n1447 C10_P_btm.n990 0.109875
R35768 C10_P_btm.n1448 C10_P_btm.n989 0.109875
R35769 C10_P_btm.n1450 C10_P_btm.n989 0.109875
R35770 C10_P_btm.n1451 C10_P_btm.n988 0.109875
R35771 C10_P_btm.n1453 C10_P_btm.n988 0.109875
R35772 C10_P_btm.n1454 C10_P_btm.n987 0.109875
R35773 C10_P_btm.n1456 C10_P_btm.n987 0.109875
R35774 C10_P_btm.n1457 C10_P_btm.n986 0.109875
R35775 C10_P_btm.n1459 C10_P_btm.n986 0.109875
R35776 C10_P_btm.n1460 C10_P_btm.n985 0.109875
R35777 C10_P_btm.n1462 C10_P_btm.n985 0.109875
R35778 C10_P_btm.n1463 C10_P_btm.n984 0.109875
R35779 C10_P_btm.n1465 C10_P_btm.n984 0.109875
R35780 C10_P_btm.n1466 C10_P_btm.n983 0.109875
R35781 C10_P_btm.n1468 C10_P_btm.n983 0.109875
R35782 C10_P_btm.n1469 C10_P_btm.n982 0.109875
R35783 C10_P_btm.n1471 C10_P_btm.n982 0.109875
R35784 C10_P_btm.n1472 C10_P_btm.n980 0.109875
R35785 C10_P_btm.n1474 C10_P_btm.n980 0.109875
R35786 C10_P_btm.n1480 C10_P_btm.n981 0.109875
R35787 C10_P_btm.n1480 C10_P_btm.n1479 0.109875
R35788 C10_P_btm.n1106 C10_P_btm.n1103 0.109875
R35789 C10_P_btm.n1104 C10_P_btm.n1103 0.109875
R35790 C10_P_btm.n1109 C10_P_btm.n1102 0.109875
R35791 C10_P_btm.n1107 C10_P_btm.n1102 0.109875
R35792 C10_P_btm.n1112 C10_P_btm.n1101 0.109875
R35793 C10_P_btm.n1110 C10_P_btm.n1101 0.109875
R35794 C10_P_btm.n1115 C10_P_btm.n1100 0.109875
R35795 C10_P_btm.n1113 C10_P_btm.n1100 0.109875
R35796 C10_P_btm.n1118 C10_P_btm.n1099 0.109875
R35797 C10_P_btm.n1116 C10_P_btm.n1099 0.109875
R35798 C10_P_btm.n1121 C10_P_btm.n1098 0.109875
R35799 C10_P_btm.n1119 C10_P_btm.n1098 0.109875
R35800 C10_P_btm.n1124 C10_P_btm.n1097 0.109875
R35801 C10_P_btm.n1122 C10_P_btm.n1097 0.109875
R35802 C10_P_btm.n1127 C10_P_btm.n1096 0.109875
R35803 C10_P_btm.n1125 C10_P_btm.n1096 0.109875
R35804 C10_P_btm.n1130 C10_P_btm.n1095 0.109875
R35805 C10_P_btm.n1128 C10_P_btm.n1095 0.109875
R35806 C10_P_btm.n1133 C10_P_btm.n1094 0.109875
R35807 C10_P_btm.n1131 C10_P_btm.n1094 0.109875
R35808 C10_P_btm.n1136 C10_P_btm.n1093 0.109875
R35809 C10_P_btm.n1134 C10_P_btm.n1093 0.109875
R35810 C10_P_btm.n1139 C10_P_btm.n1092 0.109875
R35811 C10_P_btm.n1137 C10_P_btm.n1092 0.109875
R35812 C10_P_btm.n1142 C10_P_btm.n1091 0.109875
R35813 C10_P_btm.n1140 C10_P_btm.n1091 0.109875
R35814 C10_P_btm.n1145 C10_P_btm.n1090 0.109875
R35815 C10_P_btm.n1143 C10_P_btm.n1090 0.109875
R35816 C10_P_btm.n1148 C10_P_btm.n1089 0.109875
R35817 C10_P_btm.n1146 C10_P_btm.n1089 0.109875
R35818 C10_P_btm.n1151 C10_P_btm.n1088 0.109875
R35819 C10_P_btm.n1149 C10_P_btm.n1088 0.109875
R35820 C10_P_btm.n1154 C10_P_btm.n1087 0.109875
R35821 C10_P_btm.n1152 C10_P_btm.n1087 0.109875
R35822 C10_P_btm.n1157 C10_P_btm.n1086 0.109875
R35823 C10_P_btm.n1155 C10_P_btm.n1086 0.109875
R35824 C10_P_btm.n1160 C10_P_btm.n1085 0.109875
R35825 C10_P_btm.n1158 C10_P_btm.n1085 0.109875
R35826 C10_P_btm.n1163 C10_P_btm.n1084 0.109875
R35827 C10_P_btm.n1161 C10_P_btm.n1084 0.109875
R35828 C10_P_btm.n1166 C10_P_btm.n1083 0.109875
R35829 C10_P_btm.n1164 C10_P_btm.n1083 0.109875
R35830 C10_P_btm.n1169 C10_P_btm.n1082 0.109875
R35831 C10_P_btm.n1167 C10_P_btm.n1082 0.109875
R35832 C10_P_btm.n1172 C10_P_btm.n1081 0.109875
R35833 C10_P_btm.n1170 C10_P_btm.n1081 0.109875
R35834 C10_P_btm.n1175 C10_P_btm.n1080 0.109875
R35835 C10_P_btm.n1173 C10_P_btm.n1080 0.109875
R35836 C10_P_btm.n1178 C10_P_btm.n1079 0.109875
R35837 C10_P_btm.n1176 C10_P_btm.n1079 0.109875
R35838 C10_P_btm.n1181 C10_P_btm.n1078 0.109875
R35839 C10_P_btm.n1179 C10_P_btm.n1078 0.109875
R35840 C10_P_btm.n1184 C10_P_btm.n1077 0.109875
R35841 C10_P_btm.n1182 C10_P_btm.n1077 0.109875
R35842 C10_P_btm.n1187 C10_P_btm.n1076 0.109875
R35843 C10_P_btm.n1185 C10_P_btm.n1076 0.109875
R35844 C10_P_btm.n1190 C10_P_btm.n1075 0.109875
R35845 C10_P_btm.n1188 C10_P_btm.n1075 0.109875
R35846 C10_P_btm.n1193 C10_P_btm.n1074 0.109875
R35847 C10_P_btm.n1191 C10_P_btm.n1074 0.109875
R35848 C10_P_btm.n1196 C10_P_btm.n1073 0.109875
R35849 C10_P_btm.n1194 C10_P_btm.n1073 0.109875
R35850 C10_P_btm.n1199 C10_P_btm.n1072 0.109875
R35851 C10_P_btm.n1197 C10_P_btm.n1072 0.109875
R35852 C10_P_btm.n1202 C10_P_btm.n1071 0.109875
R35853 C10_P_btm.n1200 C10_P_btm.n1071 0.109875
R35854 C10_P_btm.n1205 C10_P_btm.n1070 0.109875
R35855 C10_P_btm.n1203 C10_P_btm.n1070 0.109875
R35856 C10_P_btm.n1208 C10_P_btm.n1069 0.109875
R35857 C10_P_btm.n1206 C10_P_btm.n1069 0.109875
R35858 C10_P_btm.n1211 C10_P_btm.n1068 0.109875
R35859 C10_P_btm.n1209 C10_P_btm.n1068 0.109875
R35860 C10_P_btm.n1214 C10_P_btm.n1067 0.109875
R35861 C10_P_btm.n1212 C10_P_btm.n1067 0.109875
R35862 C10_P_btm.n1217 C10_P_btm.n1066 0.109875
R35863 C10_P_btm.n1215 C10_P_btm.n1066 0.109875
R35864 C10_P_btm.n1220 C10_P_btm.n1065 0.109875
R35865 C10_P_btm.n1218 C10_P_btm.n1065 0.109875
R35866 C10_P_btm.n1223 C10_P_btm.n1064 0.109875
R35867 C10_P_btm.n1221 C10_P_btm.n1064 0.109875
R35868 C10_P_btm.n1226 C10_P_btm.n1063 0.109875
R35869 C10_P_btm.n1224 C10_P_btm.n1063 0.109875
R35870 C10_P_btm.n1229 C10_P_btm.n1062 0.109875
R35871 C10_P_btm.n1227 C10_P_btm.n1062 0.109875
R35872 C10_P_btm.n1232 C10_P_btm.n1061 0.109875
R35873 C10_P_btm.n1230 C10_P_btm.n1061 0.109875
R35874 C10_P_btm.n1235 C10_P_btm.n1060 0.109875
R35875 C10_P_btm.n1233 C10_P_btm.n1060 0.109875
R35876 C10_P_btm.n1238 C10_P_btm.n1059 0.109875
R35877 C10_P_btm.n1236 C10_P_btm.n1059 0.109875
R35878 C10_P_btm.n1241 C10_P_btm.n1058 0.109875
R35879 C10_P_btm.n1239 C10_P_btm.n1058 0.109875
R35880 C10_P_btm.n1244 C10_P_btm.n1057 0.109875
R35881 C10_P_btm.n1242 C10_P_btm.n1057 0.109875
R35882 C10_P_btm.n1247 C10_P_btm.n1056 0.109875
R35883 C10_P_btm.n1245 C10_P_btm.n1056 0.109875
R35884 C10_P_btm.n1250 C10_P_btm.n1055 0.109875
R35885 C10_P_btm.n1248 C10_P_btm.n1055 0.109875
R35886 C10_P_btm.n1253 C10_P_btm.n1054 0.109875
R35887 C10_P_btm.n1251 C10_P_btm.n1054 0.109875
R35888 C10_P_btm.n1256 C10_P_btm.n1053 0.109875
R35889 C10_P_btm.n1254 C10_P_btm.n1053 0.109875
R35890 C10_P_btm.n1259 C10_P_btm.n1052 0.109875
R35891 C10_P_btm.n1257 C10_P_btm.n1052 0.109875
R35892 C10_P_btm.n1262 C10_P_btm.n1051 0.109875
R35893 C10_P_btm.n1260 C10_P_btm.n1051 0.109875
R35894 C10_P_btm.n1265 C10_P_btm.n1050 0.109875
R35895 C10_P_btm.n1263 C10_P_btm.n1050 0.109875
R35896 C10_P_btm.n1268 C10_P_btm.n1049 0.109875
R35897 C10_P_btm.n1266 C10_P_btm.n1049 0.109875
R35898 C10_P_btm.n1271 C10_P_btm.n1048 0.109875
R35899 C10_P_btm.n1269 C10_P_btm.n1048 0.109875
R35900 C10_P_btm.n1274 C10_P_btm.n1047 0.109875
R35901 C10_P_btm.n1272 C10_P_btm.n1047 0.109875
R35902 C10_P_btm.n1277 C10_P_btm.n1046 0.109875
R35903 C10_P_btm.n1275 C10_P_btm.n1046 0.109875
R35904 C10_P_btm.n1280 C10_P_btm.n1045 0.109875
R35905 C10_P_btm.n1278 C10_P_btm.n1045 0.109875
R35906 C10_P_btm.n1283 C10_P_btm.n1044 0.109875
R35907 C10_P_btm.n1281 C10_P_btm.n1044 0.109875
R35908 C10_P_btm.n1286 C10_P_btm.n1043 0.109875
R35909 C10_P_btm.n1286 C10_P_btm.n1285 0.109875
R35910 C10_P_btm.n1668 C10_P_btm.n919 0.109875
R35911 C10_P_btm.n1666 C10_P_btm.n919 0.109875
R35912 C10_P_btm.n1665 C10_P_btm.n920 0.109875
R35913 C10_P_btm.n1663 C10_P_btm.n920 0.109875
R35914 C10_P_btm.n1662 C10_P_btm.n921 0.109875
R35915 C10_P_btm.n1660 C10_P_btm.n921 0.109875
R35916 C10_P_btm.n1659 C10_P_btm.n922 0.109875
R35917 C10_P_btm.n1657 C10_P_btm.n922 0.109875
R35918 C10_P_btm.n1656 C10_P_btm.n923 0.109875
R35919 C10_P_btm.n1654 C10_P_btm.n923 0.109875
R35920 C10_P_btm.n1653 C10_P_btm.n924 0.109875
R35921 C10_P_btm.n1651 C10_P_btm.n924 0.109875
R35922 C10_P_btm.n1650 C10_P_btm.n925 0.109875
R35923 C10_P_btm.n1648 C10_P_btm.n925 0.109875
R35924 C10_P_btm.n1647 C10_P_btm.n926 0.109875
R35925 C10_P_btm.n1645 C10_P_btm.n926 0.109875
R35926 C10_P_btm.n1644 C10_P_btm.n927 0.109875
R35927 C10_P_btm.n1642 C10_P_btm.n927 0.109875
R35928 C10_P_btm.n1641 C10_P_btm.n928 0.109875
R35929 C10_P_btm.n1639 C10_P_btm.n928 0.109875
R35930 C10_P_btm.n1638 C10_P_btm.n929 0.109875
R35931 C10_P_btm.n1636 C10_P_btm.n929 0.109875
R35932 C10_P_btm.n1635 C10_P_btm.n930 0.109875
R35933 C10_P_btm.n1633 C10_P_btm.n930 0.109875
R35934 C10_P_btm.n1632 C10_P_btm.n931 0.109875
R35935 C10_P_btm.n1630 C10_P_btm.n931 0.109875
R35936 C10_P_btm.n1629 C10_P_btm.n932 0.109875
R35937 C10_P_btm.n1627 C10_P_btm.n932 0.109875
R35938 C10_P_btm.n1626 C10_P_btm.n933 0.109875
R35939 C10_P_btm.n1624 C10_P_btm.n933 0.109875
R35940 C10_P_btm.n1623 C10_P_btm.n934 0.109875
R35941 C10_P_btm.n1621 C10_P_btm.n934 0.109875
R35942 C10_P_btm.n1620 C10_P_btm.n935 0.109875
R35943 C10_P_btm.n1618 C10_P_btm.n935 0.109875
R35944 C10_P_btm.n1617 C10_P_btm.n936 0.109875
R35945 C10_P_btm.n1615 C10_P_btm.n936 0.109875
R35946 C10_P_btm.n1614 C10_P_btm.n937 0.109875
R35947 C10_P_btm.n1612 C10_P_btm.n937 0.109875
R35948 C10_P_btm.n1611 C10_P_btm.n938 0.109875
R35949 C10_P_btm.n1609 C10_P_btm.n938 0.109875
R35950 C10_P_btm.n1608 C10_P_btm.n939 0.109875
R35951 C10_P_btm.n1606 C10_P_btm.n939 0.109875
R35952 C10_P_btm.n1605 C10_P_btm.n940 0.109875
R35953 C10_P_btm.n1603 C10_P_btm.n940 0.109875
R35954 C10_P_btm.n1602 C10_P_btm.n941 0.109875
R35955 C10_P_btm.n1600 C10_P_btm.n941 0.109875
R35956 C10_P_btm.n1599 C10_P_btm.n942 0.109875
R35957 C10_P_btm.n1597 C10_P_btm.n942 0.109875
R35958 C10_P_btm.n1596 C10_P_btm.n943 0.109875
R35959 C10_P_btm.n1594 C10_P_btm.n943 0.109875
R35960 C10_P_btm.n1593 C10_P_btm.n944 0.109875
R35961 C10_P_btm.n1591 C10_P_btm.n944 0.109875
R35962 C10_P_btm.n1590 C10_P_btm.n945 0.109875
R35963 C10_P_btm.n1588 C10_P_btm.n945 0.109875
R35964 C10_P_btm.n1587 C10_P_btm.n946 0.109875
R35965 C10_P_btm.n1585 C10_P_btm.n946 0.109875
R35966 C10_P_btm.n1584 C10_P_btm.n947 0.109875
R35967 C10_P_btm.n1582 C10_P_btm.n947 0.109875
R35968 C10_P_btm.n1581 C10_P_btm.n948 0.109875
R35969 C10_P_btm.n1579 C10_P_btm.n948 0.109875
R35970 C10_P_btm.n1578 C10_P_btm.n949 0.109875
R35971 C10_P_btm.n1576 C10_P_btm.n949 0.109875
R35972 C10_P_btm.n1575 C10_P_btm.n950 0.109875
R35973 C10_P_btm.n1573 C10_P_btm.n950 0.109875
R35974 C10_P_btm.n1572 C10_P_btm.n951 0.109875
R35975 C10_P_btm.n1570 C10_P_btm.n951 0.109875
R35976 C10_P_btm.n1569 C10_P_btm.n952 0.109875
R35977 C10_P_btm.n1567 C10_P_btm.n952 0.109875
R35978 C10_P_btm.n1566 C10_P_btm.n953 0.109875
R35979 C10_P_btm.n1564 C10_P_btm.n953 0.109875
R35980 C10_P_btm.n1563 C10_P_btm.n954 0.109875
R35981 C10_P_btm.n1561 C10_P_btm.n954 0.109875
R35982 C10_P_btm.n1560 C10_P_btm.n955 0.109875
R35983 C10_P_btm.n1558 C10_P_btm.n955 0.109875
R35984 C10_P_btm.n1557 C10_P_btm.n956 0.109875
R35985 C10_P_btm.n1555 C10_P_btm.n956 0.109875
R35986 C10_P_btm.n1554 C10_P_btm.n957 0.109875
R35987 C10_P_btm.n1552 C10_P_btm.n957 0.109875
R35988 C10_P_btm.n1551 C10_P_btm.n958 0.109875
R35989 C10_P_btm.n1549 C10_P_btm.n958 0.109875
R35990 C10_P_btm.n1548 C10_P_btm.n959 0.109875
R35991 C10_P_btm.n1546 C10_P_btm.n959 0.109875
R35992 C10_P_btm.n1545 C10_P_btm.n960 0.109875
R35993 C10_P_btm.n1543 C10_P_btm.n960 0.109875
R35994 C10_P_btm.n1542 C10_P_btm.n961 0.109875
R35995 C10_P_btm.n1540 C10_P_btm.n961 0.109875
R35996 C10_P_btm.n1539 C10_P_btm.n962 0.109875
R35997 C10_P_btm.n1537 C10_P_btm.n962 0.109875
R35998 C10_P_btm.n1536 C10_P_btm.n963 0.109875
R35999 C10_P_btm.n1534 C10_P_btm.n963 0.109875
R36000 C10_P_btm.n1533 C10_P_btm.n964 0.109875
R36001 C10_P_btm.n1531 C10_P_btm.n964 0.109875
R36002 C10_P_btm.n1530 C10_P_btm.n965 0.109875
R36003 C10_P_btm.n1528 C10_P_btm.n965 0.109875
R36004 C10_P_btm.n1527 C10_P_btm.n966 0.109875
R36005 C10_P_btm.n1525 C10_P_btm.n966 0.109875
R36006 C10_P_btm.n1524 C10_P_btm.n967 0.109875
R36007 C10_P_btm.n1522 C10_P_btm.n967 0.109875
R36008 C10_P_btm.n1521 C10_P_btm.n968 0.109875
R36009 C10_P_btm.n1519 C10_P_btm.n968 0.109875
R36010 C10_P_btm.n1518 C10_P_btm.n969 0.109875
R36011 C10_P_btm.n1516 C10_P_btm.n969 0.109875
R36012 C10_P_btm.n1515 C10_P_btm.n970 0.109875
R36013 C10_P_btm.n1513 C10_P_btm.n970 0.109875
R36014 C10_P_btm.n1512 C10_P_btm.n971 0.109875
R36015 C10_P_btm.n1510 C10_P_btm.n971 0.109875
R36016 C10_P_btm.n1509 C10_P_btm.n972 0.109875
R36017 C10_P_btm.n1507 C10_P_btm.n972 0.109875
R36018 C10_P_btm.n1506 C10_P_btm.n973 0.109875
R36019 C10_P_btm.n1504 C10_P_btm.n973 0.109875
R36020 C10_P_btm.n1503 C10_P_btm.n974 0.109875
R36021 C10_P_btm.n1501 C10_P_btm.n974 0.109875
R36022 C10_P_btm.n1500 C10_P_btm.n975 0.109875
R36023 C10_P_btm.n1498 C10_P_btm.n975 0.109875
R36024 C10_P_btm.n1497 C10_P_btm.n976 0.109875
R36025 C10_P_btm.n1495 C10_P_btm.n976 0.109875
R36026 C10_P_btm.n1494 C10_P_btm.n977 0.109875
R36027 C10_P_btm.n1492 C10_P_btm.n977 0.109875
R36028 C10_P_btm.n1491 C10_P_btm.n978 0.109875
R36029 C10_P_btm.n1489 C10_P_btm.n978 0.109875
R36030 C10_P_btm.n1488 C10_P_btm.n979 0.109875
R36031 C10_P_btm.n1486 C10_P_btm.n979 0.109875
R36032 C10_P_btm.n1485 C10_P_btm.n1481 0.109875
R36033 C10_P_btm.n1483 C10_P_btm.n1481 0.109875
R36034 C10_P_btm.n1856 C10_P_btm.n609 0.109875
R36035 C10_P_btm.n1858 C10_P_btm.n609 0.109875
R36036 C10_P_btm.n1853 C10_P_btm.n612 0.109875
R36037 C10_P_btm.n1855 C10_P_btm.n612 0.109875
R36038 C10_P_btm.n1850 C10_P_btm.n613 0.109875
R36039 C10_P_btm.n1852 C10_P_btm.n613 0.109875
R36040 C10_P_btm.n1847 C10_P_btm.n614 0.109875
R36041 C10_P_btm.n1849 C10_P_btm.n614 0.109875
R36042 C10_P_btm.n1844 C10_P_btm.n615 0.109875
R36043 C10_P_btm.n1846 C10_P_btm.n615 0.109875
R36044 C10_P_btm.n1841 C10_P_btm.n616 0.109875
R36045 C10_P_btm.n1843 C10_P_btm.n616 0.109875
R36046 C10_P_btm.n1838 C10_P_btm.n617 0.109875
R36047 C10_P_btm.n1840 C10_P_btm.n617 0.109875
R36048 C10_P_btm.n1835 C10_P_btm.n618 0.109875
R36049 C10_P_btm.n1837 C10_P_btm.n618 0.109875
R36050 C10_P_btm.n1832 C10_P_btm.n619 0.109875
R36051 C10_P_btm.n1834 C10_P_btm.n619 0.109875
R36052 C10_P_btm.n1829 C10_P_btm.n620 0.109875
R36053 C10_P_btm.n1831 C10_P_btm.n620 0.109875
R36054 C10_P_btm.n1826 C10_P_btm.n621 0.109875
R36055 C10_P_btm.n1828 C10_P_btm.n621 0.109875
R36056 C10_P_btm.n1823 C10_P_btm.n622 0.109875
R36057 C10_P_btm.n1825 C10_P_btm.n622 0.109875
R36058 C10_P_btm.n1820 C10_P_btm.n623 0.109875
R36059 C10_P_btm.n1822 C10_P_btm.n623 0.109875
R36060 C10_P_btm.n1817 C10_P_btm.n624 0.109875
R36061 C10_P_btm.n1819 C10_P_btm.n624 0.109875
R36062 C10_P_btm.n1814 C10_P_btm.n625 0.109875
R36063 C10_P_btm.n1816 C10_P_btm.n625 0.109875
R36064 C10_P_btm.n1811 C10_P_btm.n626 0.109875
R36065 C10_P_btm.n1813 C10_P_btm.n626 0.109875
R36066 C10_P_btm.n1808 C10_P_btm.n627 0.109875
R36067 C10_P_btm.n1810 C10_P_btm.n627 0.109875
R36068 C10_P_btm.n1805 C10_P_btm.n628 0.109875
R36069 C10_P_btm.n1807 C10_P_btm.n628 0.109875
R36070 C10_P_btm.n1802 C10_P_btm.n629 0.109875
R36071 C10_P_btm.n1804 C10_P_btm.n629 0.109875
R36072 C10_P_btm.n1799 C10_P_btm.n630 0.109875
R36073 C10_P_btm.n1801 C10_P_btm.n630 0.109875
R36074 C10_P_btm.n1796 C10_P_btm.n631 0.109875
R36075 C10_P_btm.n1798 C10_P_btm.n631 0.109875
R36076 C10_P_btm.n1793 C10_P_btm.n632 0.109875
R36077 C10_P_btm.n1795 C10_P_btm.n632 0.109875
R36078 C10_P_btm.n1790 C10_P_btm.n633 0.109875
R36079 C10_P_btm.n1792 C10_P_btm.n633 0.109875
R36080 C10_P_btm.n1787 C10_P_btm.n634 0.109875
R36081 C10_P_btm.n1789 C10_P_btm.n634 0.109875
R36082 C10_P_btm.n1784 C10_P_btm.n635 0.109875
R36083 C10_P_btm.n1786 C10_P_btm.n635 0.109875
R36084 C10_P_btm.n1781 C10_P_btm.n636 0.109875
R36085 C10_P_btm.n1783 C10_P_btm.n636 0.109875
R36086 C10_P_btm.n1778 C10_P_btm.n637 0.109875
R36087 C10_P_btm.n1780 C10_P_btm.n637 0.109875
R36088 C10_P_btm.n1775 C10_P_btm.n638 0.109875
R36089 C10_P_btm.n1777 C10_P_btm.n638 0.109875
R36090 C10_P_btm.n1772 C10_P_btm.n639 0.109875
R36091 C10_P_btm.n1774 C10_P_btm.n639 0.109875
R36092 C10_P_btm.n1769 C10_P_btm.n640 0.109875
R36093 C10_P_btm.n1771 C10_P_btm.n640 0.109875
R36094 C10_P_btm.n1766 C10_P_btm.n641 0.109875
R36095 C10_P_btm.n1768 C10_P_btm.n641 0.109875
R36096 C10_P_btm.n1763 C10_P_btm.n642 0.109875
R36097 C10_P_btm.n1765 C10_P_btm.n642 0.109875
R36098 C10_P_btm.n1760 C10_P_btm.n643 0.109875
R36099 C10_P_btm.n1762 C10_P_btm.n643 0.109875
R36100 C10_P_btm.n1757 C10_P_btm.n644 0.109875
R36101 C10_P_btm.n1759 C10_P_btm.n644 0.109875
R36102 C10_P_btm.n1754 C10_P_btm.n645 0.109875
R36103 C10_P_btm.n1756 C10_P_btm.n645 0.109875
R36104 C10_P_btm.n1751 C10_P_btm.n646 0.109875
R36105 C10_P_btm.n1753 C10_P_btm.n646 0.109875
R36106 C10_P_btm.n1748 C10_P_btm.n647 0.109875
R36107 C10_P_btm.n1750 C10_P_btm.n647 0.109875
R36108 C10_P_btm.n1745 C10_P_btm.n648 0.109875
R36109 C10_P_btm.n1747 C10_P_btm.n648 0.109875
R36110 C10_P_btm.n1742 C10_P_btm.n649 0.109875
R36111 C10_P_btm.n1744 C10_P_btm.n649 0.109875
R36112 C10_P_btm.n1739 C10_P_btm.n650 0.109875
R36113 C10_P_btm.n1741 C10_P_btm.n650 0.109875
R36114 C10_P_btm.n1736 C10_P_btm.n651 0.109875
R36115 C10_P_btm.n1738 C10_P_btm.n651 0.109875
R36116 C10_P_btm.n1733 C10_P_btm.n652 0.109875
R36117 C10_P_btm.n1735 C10_P_btm.n652 0.109875
R36118 C10_P_btm.n1730 C10_P_btm.n653 0.109875
R36119 C10_P_btm.n1732 C10_P_btm.n653 0.109875
R36120 C10_P_btm.n1727 C10_P_btm.n654 0.109875
R36121 C10_P_btm.n1729 C10_P_btm.n654 0.109875
R36122 C10_P_btm.n1724 C10_P_btm.n655 0.109875
R36123 C10_P_btm.n1726 C10_P_btm.n655 0.109875
R36124 C10_P_btm.n1721 C10_P_btm.n656 0.109875
R36125 C10_P_btm.n1723 C10_P_btm.n656 0.109875
R36126 C10_P_btm.n1718 C10_P_btm.n657 0.109875
R36127 C10_P_btm.n1720 C10_P_btm.n657 0.109875
R36128 C10_P_btm.n1715 C10_P_btm.n658 0.109875
R36129 C10_P_btm.n1717 C10_P_btm.n658 0.109875
R36130 C10_P_btm.n1712 C10_P_btm.n659 0.109875
R36131 C10_P_btm.n1714 C10_P_btm.n659 0.109875
R36132 C10_P_btm.n1709 C10_P_btm.n660 0.109875
R36133 C10_P_btm.n1711 C10_P_btm.n660 0.109875
R36134 C10_P_btm.n1706 C10_P_btm.n661 0.109875
R36135 C10_P_btm.n1708 C10_P_btm.n661 0.109875
R36136 C10_P_btm.n1703 C10_P_btm.n662 0.109875
R36137 C10_P_btm.n1705 C10_P_btm.n662 0.109875
R36138 C10_P_btm.n1700 C10_P_btm.n663 0.109875
R36139 C10_P_btm.n1702 C10_P_btm.n663 0.109875
R36140 C10_P_btm.n1697 C10_P_btm.n664 0.109875
R36141 C10_P_btm.n1699 C10_P_btm.n664 0.109875
R36142 C10_P_btm.n1694 C10_P_btm.n665 0.109875
R36143 C10_P_btm.n1696 C10_P_btm.n665 0.109875
R36144 C10_P_btm.n1691 C10_P_btm.n666 0.109875
R36145 C10_P_btm.n1693 C10_P_btm.n666 0.109875
R36146 C10_P_btm.n1688 C10_P_btm.n667 0.109875
R36147 C10_P_btm.n1690 C10_P_btm.n667 0.109875
R36148 C10_P_btm.n1685 C10_P_btm.n668 0.109875
R36149 C10_P_btm.n1687 C10_P_btm.n668 0.109875
R36150 C10_P_btm.n1682 C10_P_btm.n669 0.109875
R36151 C10_P_btm.n1684 C10_P_btm.n669 0.109875
R36152 C10_P_btm.n1679 C10_P_btm.n670 0.109875
R36153 C10_P_btm.n1681 C10_P_btm.n670 0.109875
R36154 C10_P_btm.n1676 C10_P_btm.n671 0.109875
R36155 C10_P_btm.n1678 C10_P_btm.n671 0.109875
R36156 C10_P_btm.n1673 C10_P_btm.n917 0.109875
R36157 C10_P_btm.n1675 C10_P_btm.n917 0.109875
R36158 C10_P_btm.n916 C10_P_btm.n673 0.109875
R36159 C10_P_btm.n916 C10_P_btm.n915 0.109875
R36160 C10_P_btm.n913 C10_P_btm.n674 0.109875
R36161 C10_P_btm.n911 C10_P_btm.n674 0.109875
R36162 C10_P_btm.n910 C10_P_btm.n675 0.109875
R36163 C10_P_btm.n908 C10_P_btm.n675 0.109875
R36164 C10_P_btm.n907 C10_P_btm.n676 0.109875
R36165 C10_P_btm.n905 C10_P_btm.n676 0.109875
R36166 C10_P_btm.n904 C10_P_btm.n677 0.109875
R36167 C10_P_btm.n902 C10_P_btm.n677 0.109875
R36168 C10_P_btm.n901 C10_P_btm.n678 0.109875
R36169 C10_P_btm.n899 C10_P_btm.n678 0.109875
R36170 C10_P_btm.n898 C10_P_btm.n679 0.109875
R36171 C10_P_btm.n896 C10_P_btm.n679 0.109875
R36172 C10_P_btm.n895 C10_P_btm.n680 0.109875
R36173 C10_P_btm.n893 C10_P_btm.n680 0.109875
R36174 C10_P_btm.n892 C10_P_btm.n681 0.109875
R36175 C10_P_btm.n890 C10_P_btm.n681 0.109875
R36176 C10_P_btm.n889 C10_P_btm.n682 0.109875
R36177 C10_P_btm.n887 C10_P_btm.n682 0.109875
R36178 C10_P_btm.n886 C10_P_btm.n683 0.109875
R36179 C10_P_btm.n884 C10_P_btm.n683 0.109875
R36180 C10_P_btm.n883 C10_P_btm.n684 0.109875
R36181 C10_P_btm.n881 C10_P_btm.n684 0.109875
R36182 C10_P_btm.n880 C10_P_btm.n685 0.109875
R36183 C10_P_btm.n878 C10_P_btm.n685 0.109875
R36184 C10_P_btm.n877 C10_P_btm.n686 0.109875
R36185 C10_P_btm.n875 C10_P_btm.n686 0.109875
R36186 C10_P_btm.n874 C10_P_btm.n687 0.109875
R36187 C10_P_btm.n872 C10_P_btm.n687 0.109875
R36188 C10_P_btm.n871 C10_P_btm.n688 0.109875
R36189 C10_P_btm.n869 C10_P_btm.n688 0.109875
R36190 C10_P_btm.n868 C10_P_btm.n689 0.109875
R36191 C10_P_btm.n866 C10_P_btm.n689 0.109875
R36192 C10_P_btm.n865 C10_P_btm.n690 0.109875
R36193 C10_P_btm.n863 C10_P_btm.n690 0.109875
R36194 C10_P_btm.n862 C10_P_btm.n691 0.109875
R36195 C10_P_btm.n860 C10_P_btm.n691 0.109875
R36196 C10_P_btm.n859 C10_P_btm.n692 0.109875
R36197 C10_P_btm.n857 C10_P_btm.n692 0.109875
R36198 C10_P_btm.n856 C10_P_btm.n693 0.109875
R36199 C10_P_btm.n854 C10_P_btm.n693 0.109875
R36200 C10_P_btm.n853 C10_P_btm.n694 0.109875
R36201 C10_P_btm.n851 C10_P_btm.n694 0.109875
R36202 C10_P_btm.n850 C10_P_btm.n695 0.109875
R36203 C10_P_btm.n848 C10_P_btm.n695 0.109875
R36204 C10_P_btm.n847 C10_P_btm.n696 0.109875
R36205 C10_P_btm.n845 C10_P_btm.n696 0.109875
R36206 C10_P_btm.n844 C10_P_btm.n697 0.109875
R36207 C10_P_btm.n842 C10_P_btm.n697 0.109875
R36208 C10_P_btm.n841 C10_P_btm.n698 0.109875
R36209 C10_P_btm.n839 C10_P_btm.n698 0.109875
R36210 C10_P_btm.n838 C10_P_btm.n699 0.109875
R36211 C10_P_btm.n836 C10_P_btm.n699 0.109875
R36212 C10_P_btm.n835 C10_P_btm.n700 0.109875
R36213 C10_P_btm.n833 C10_P_btm.n700 0.109875
R36214 C10_P_btm.n832 C10_P_btm.n701 0.109875
R36215 C10_P_btm.n830 C10_P_btm.n701 0.109875
R36216 C10_P_btm.n829 C10_P_btm.n702 0.109875
R36217 C10_P_btm.n827 C10_P_btm.n702 0.109875
R36218 C10_P_btm.n826 C10_P_btm.n703 0.109875
R36219 C10_P_btm.n824 C10_P_btm.n703 0.109875
R36220 C10_P_btm.n823 C10_P_btm.n704 0.109875
R36221 C10_P_btm.n821 C10_P_btm.n704 0.109875
R36222 C10_P_btm.n820 C10_P_btm.n705 0.109875
R36223 C10_P_btm.n818 C10_P_btm.n705 0.109875
R36224 C10_P_btm.n817 C10_P_btm.n706 0.109875
R36225 C10_P_btm.n815 C10_P_btm.n706 0.109875
R36226 C10_P_btm.n814 C10_P_btm.n707 0.109875
R36227 C10_P_btm.n812 C10_P_btm.n707 0.109875
R36228 C10_P_btm.n811 C10_P_btm.n708 0.109875
R36229 C10_P_btm.n809 C10_P_btm.n708 0.109875
R36230 C10_P_btm.n808 C10_P_btm.n709 0.109875
R36231 C10_P_btm.n806 C10_P_btm.n709 0.109875
R36232 C10_P_btm.n805 C10_P_btm.n710 0.109875
R36233 C10_P_btm.n803 C10_P_btm.n710 0.109875
R36234 C10_P_btm.n802 C10_P_btm.n711 0.109875
R36235 C10_P_btm.n800 C10_P_btm.n711 0.109875
R36236 C10_P_btm.n799 C10_P_btm.n712 0.109875
R36237 C10_P_btm.n797 C10_P_btm.n712 0.109875
R36238 C10_P_btm.n796 C10_P_btm.n713 0.109875
R36239 C10_P_btm.n794 C10_P_btm.n713 0.109875
R36240 C10_P_btm.n793 C10_P_btm.n714 0.109875
R36241 C10_P_btm.n791 C10_P_btm.n714 0.109875
R36242 C10_P_btm.n790 C10_P_btm.n715 0.109875
R36243 C10_P_btm.n788 C10_P_btm.n715 0.109875
R36244 C10_P_btm.n787 C10_P_btm.n716 0.109875
R36245 C10_P_btm.n785 C10_P_btm.n716 0.109875
R36246 C10_P_btm.n784 C10_P_btm.n717 0.109875
R36247 C10_P_btm.n782 C10_P_btm.n717 0.109875
R36248 C10_P_btm.n781 C10_P_btm.n718 0.109875
R36249 C10_P_btm.n779 C10_P_btm.n718 0.109875
R36250 C10_P_btm.n778 C10_P_btm.n719 0.109875
R36251 C10_P_btm.n776 C10_P_btm.n719 0.109875
R36252 C10_P_btm.n775 C10_P_btm.n720 0.109875
R36253 C10_P_btm.n773 C10_P_btm.n720 0.109875
R36254 C10_P_btm.n772 C10_P_btm.n721 0.109875
R36255 C10_P_btm.n770 C10_P_btm.n721 0.109875
R36256 C10_P_btm.n769 C10_P_btm.n722 0.109875
R36257 C10_P_btm.n767 C10_P_btm.n722 0.109875
R36258 C10_P_btm.n766 C10_P_btm.n723 0.109875
R36259 C10_P_btm.n764 C10_P_btm.n723 0.109875
R36260 C10_P_btm.n763 C10_P_btm.n724 0.109875
R36261 C10_P_btm.n761 C10_P_btm.n724 0.109875
R36262 C10_P_btm.n760 C10_P_btm.n725 0.109875
R36263 C10_P_btm.n758 C10_P_btm.n725 0.109875
R36264 C10_P_btm.n757 C10_P_btm.n726 0.109875
R36265 C10_P_btm.n755 C10_P_btm.n726 0.109875
R36266 C10_P_btm.n754 C10_P_btm.n727 0.109875
R36267 C10_P_btm.n752 C10_P_btm.n727 0.109875
R36268 C10_P_btm.n751 C10_P_btm.n728 0.109875
R36269 C10_P_btm.n749 C10_P_btm.n728 0.109875
R36270 C10_P_btm.n748 C10_P_btm.n729 0.109875
R36271 C10_P_btm.n746 C10_P_btm.n729 0.109875
R36272 C10_P_btm.n745 C10_P_btm.n730 0.109875
R36273 C10_P_btm.n743 C10_P_btm.n730 0.109875
R36274 C10_P_btm.n742 C10_P_btm.n731 0.109875
R36275 C10_P_btm.n740 C10_P_btm.n731 0.109875
R36276 C10_P_btm.n739 C10_P_btm.n732 0.109875
R36277 C10_P_btm.n737 C10_P_btm.n732 0.109875
R36278 C10_P_btm.n736 C10_P_btm.n733 0.109875
R36279 C10_P_btm.n734 C10_P_btm.n733 0.109875
R36280 C10_P_btm.n1865 C10_P_btm.n610 0.109875
R36281 C10_P_btm.n1865 C10_P_btm.n1864 0.109875
R36282 C10_P_btm.n1870 C10_P_btm.n1866 0.109875
R36283 C10_P_btm.n1868 C10_P_btm.n1866 0.109875
R36284 C10_P_btm.n1873 C10_P_btm.n608 0.109875
R36285 C10_P_btm.n1871 C10_P_btm.n608 0.109875
R36286 C10_P_btm.n1876 C10_P_btm.n607 0.109875
R36287 C10_P_btm.n1874 C10_P_btm.n607 0.109875
R36288 C10_P_btm.n1879 C10_P_btm.n606 0.109875
R36289 C10_P_btm.n1877 C10_P_btm.n606 0.109875
R36290 C10_P_btm.n1882 C10_P_btm.n605 0.109875
R36291 C10_P_btm.n1880 C10_P_btm.n605 0.109875
R36292 C10_P_btm.n1885 C10_P_btm.n604 0.109875
R36293 C10_P_btm.n1883 C10_P_btm.n604 0.109875
R36294 C10_P_btm.n1888 C10_P_btm.n603 0.109875
R36295 C10_P_btm.n1886 C10_P_btm.n603 0.109875
R36296 C10_P_btm.n1891 C10_P_btm.n602 0.109875
R36297 C10_P_btm.n1889 C10_P_btm.n602 0.109875
R36298 C10_P_btm.n1894 C10_P_btm.n601 0.109875
R36299 C10_P_btm.n1892 C10_P_btm.n601 0.109875
R36300 C10_P_btm.n1897 C10_P_btm.n600 0.109875
R36301 C10_P_btm.n1895 C10_P_btm.n600 0.109875
R36302 C10_P_btm.n1900 C10_P_btm.n599 0.109875
R36303 C10_P_btm.n1898 C10_P_btm.n599 0.109875
R36304 C10_P_btm.n1903 C10_P_btm.n598 0.109875
R36305 C10_P_btm.n1901 C10_P_btm.n598 0.109875
R36306 C10_P_btm.n1906 C10_P_btm.n597 0.109875
R36307 C10_P_btm.n1904 C10_P_btm.n597 0.109875
R36308 C10_P_btm.n1909 C10_P_btm.n596 0.109875
R36309 C10_P_btm.n1907 C10_P_btm.n596 0.109875
R36310 C10_P_btm.n1912 C10_P_btm.n595 0.109875
R36311 C10_P_btm.n1910 C10_P_btm.n595 0.109875
R36312 C10_P_btm.n1915 C10_P_btm.n594 0.109875
R36313 C10_P_btm.n1913 C10_P_btm.n594 0.109875
R36314 C10_P_btm.n1918 C10_P_btm.n593 0.109875
R36315 C10_P_btm.n1916 C10_P_btm.n593 0.109875
R36316 C10_P_btm.n1921 C10_P_btm.n592 0.109875
R36317 C10_P_btm.n1919 C10_P_btm.n592 0.109875
R36318 C10_P_btm.n1924 C10_P_btm.n591 0.109875
R36319 C10_P_btm.n1922 C10_P_btm.n591 0.109875
R36320 C10_P_btm.n1927 C10_P_btm.n590 0.109875
R36321 C10_P_btm.n1925 C10_P_btm.n590 0.109875
R36322 C10_P_btm.n1930 C10_P_btm.n589 0.109875
R36323 C10_P_btm.n1928 C10_P_btm.n589 0.109875
R36324 C10_P_btm.n1933 C10_P_btm.n588 0.109875
R36325 C10_P_btm.n1931 C10_P_btm.n588 0.109875
R36326 C10_P_btm.n1936 C10_P_btm.n587 0.109875
R36327 C10_P_btm.n1934 C10_P_btm.n587 0.109875
R36328 C10_P_btm.n1939 C10_P_btm.n586 0.109875
R36329 C10_P_btm.n1937 C10_P_btm.n586 0.109875
R36330 C10_P_btm.n1942 C10_P_btm.n585 0.109875
R36331 C10_P_btm.n1940 C10_P_btm.n585 0.109875
R36332 C10_P_btm.n1945 C10_P_btm.n584 0.109875
R36333 C10_P_btm.n1943 C10_P_btm.n584 0.109875
R36334 C10_P_btm.n1948 C10_P_btm.n583 0.109875
R36335 C10_P_btm.n1946 C10_P_btm.n583 0.109875
R36336 C10_P_btm.n1951 C10_P_btm.n582 0.109875
R36337 C10_P_btm.n1949 C10_P_btm.n582 0.109875
R36338 C10_P_btm.n1954 C10_P_btm.n581 0.109875
R36339 C10_P_btm.n1952 C10_P_btm.n581 0.109875
R36340 C10_P_btm.n1957 C10_P_btm.n580 0.109875
R36341 C10_P_btm.n1955 C10_P_btm.n580 0.109875
R36342 C10_P_btm.n1960 C10_P_btm.n579 0.109875
R36343 C10_P_btm.n1958 C10_P_btm.n579 0.109875
R36344 C10_P_btm.n1963 C10_P_btm.n578 0.109875
R36345 C10_P_btm.n1961 C10_P_btm.n578 0.109875
R36346 C10_P_btm.n1966 C10_P_btm.n577 0.109875
R36347 C10_P_btm.n1964 C10_P_btm.n577 0.109875
R36348 C10_P_btm.n1969 C10_P_btm.n576 0.109875
R36349 C10_P_btm.n1967 C10_P_btm.n576 0.109875
R36350 C10_P_btm.n1972 C10_P_btm.n575 0.109875
R36351 C10_P_btm.n1970 C10_P_btm.n575 0.109875
R36352 C10_P_btm.n1975 C10_P_btm.n574 0.109875
R36353 C10_P_btm.n1973 C10_P_btm.n574 0.109875
R36354 C10_P_btm.n1978 C10_P_btm.n573 0.109875
R36355 C10_P_btm.n1976 C10_P_btm.n573 0.109875
R36356 C10_P_btm.n1981 C10_P_btm.n572 0.109875
R36357 C10_P_btm.n1979 C10_P_btm.n572 0.109875
R36358 C10_P_btm.n1984 C10_P_btm.n571 0.109875
R36359 C10_P_btm.n1982 C10_P_btm.n571 0.109875
R36360 C10_P_btm.n1987 C10_P_btm.n570 0.109875
R36361 C10_P_btm.n1985 C10_P_btm.n570 0.109875
R36362 C10_P_btm.n1990 C10_P_btm.n569 0.109875
R36363 C10_P_btm.n1988 C10_P_btm.n569 0.109875
R36364 C10_P_btm.n1993 C10_P_btm.n568 0.109875
R36365 C10_P_btm.n1991 C10_P_btm.n568 0.109875
R36366 C10_P_btm.n1996 C10_P_btm.n567 0.109875
R36367 C10_P_btm.n1994 C10_P_btm.n567 0.109875
R36368 C10_P_btm.n1999 C10_P_btm.n566 0.109875
R36369 C10_P_btm.n1997 C10_P_btm.n566 0.109875
R36370 C10_P_btm.n2002 C10_P_btm.n565 0.109875
R36371 C10_P_btm.n2000 C10_P_btm.n565 0.109875
R36372 C10_P_btm.n2005 C10_P_btm.n564 0.109875
R36373 C10_P_btm.n2003 C10_P_btm.n564 0.109875
R36374 C10_P_btm.n2008 C10_P_btm.n563 0.109875
R36375 C10_P_btm.n2006 C10_P_btm.n563 0.109875
R36376 C10_P_btm.n2011 C10_P_btm.n562 0.109875
R36377 C10_P_btm.n2009 C10_P_btm.n562 0.109875
R36378 C10_P_btm.n2014 C10_P_btm.n561 0.109875
R36379 C10_P_btm.n2012 C10_P_btm.n561 0.109875
R36380 C10_P_btm.n2017 C10_P_btm.n560 0.109875
R36381 C10_P_btm.n2015 C10_P_btm.n560 0.109875
R36382 C10_P_btm.n2020 C10_P_btm.n559 0.109875
R36383 C10_P_btm.n2018 C10_P_btm.n559 0.109875
R36384 C10_P_btm.n2023 C10_P_btm.n558 0.109875
R36385 C10_P_btm.n2021 C10_P_btm.n558 0.109875
R36386 C10_P_btm.n2026 C10_P_btm.n557 0.109875
R36387 C10_P_btm.n2024 C10_P_btm.n557 0.109875
R36388 C10_P_btm.n2029 C10_P_btm.n556 0.109875
R36389 C10_P_btm.n2027 C10_P_btm.n556 0.109875
R36390 C10_P_btm.n2032 C10_P_btm.n555 0.109875
R36391 C10_P_btm.n2030 C10_P_btm.n555 0.109875
R36392 C10_P_btm.n2035 C10_P_btm.n554 0.109875
R36393 C10_P_btm.n2033 C10_P_btm.n554 0.109875
R36394 C10_P_btm.n2038 C10_P_btm.n553 0.109875
R36395 C10_P_btm.n2036 C10_P_btm.n553 0.109875
R36396 C10_P_btm.n2041 C10_P_btm.n552 0.109875
R36397 C10_P_btm.n2039 C10_P_btm.n552 0.109875
R36398 C10_P_btm.n2044 C10_P_btm.n551 0.109875
R36399 C10_P_btm.n2042 C10_P_btm.n551 0.109875
R36400 C10_P_btm.n2047 C10_P_btm.n550 0.109875
R36401 C10_P_btm.n2045 C10_P_btm.n550 0.109875
R36402 C10_P_btm.n2050 C10_P_btm.n549 0.109875
R36403 C10_P_btm.n2048 C10_P_btm.n549 0.109875
R36404 C10_P_btm.n2053 C10_P_btm.n548 0.109875
R36405 C10_P_btm.n2051 C10_P_btm.n548 0.109875
R36406 C10_P_btm.n3109 C10_P_btm.n546 0.109875
R36407 C10_P_btm.n3111 C10_P_btm.n546 0.109875
R36408 C10_P_btm.n3112 C10_P_btm.n545 0.109875
R36409 C10_P_btm.n3114 C10_P_btm.n545 0.109875
R36410 C10_P_btm.n3115 C10_P_btm.n544 0.109875
R36411 C10_P_btm.n3117 C10_P_btm.n544 0.109875
R36412 C10_P_btm.n3118 C10_P_btm.n543 0.109875
R36413 C10_P_btm.n3120 C10_P_btm.n543 0.109875
R36414 C10_P_btm.n3121 C10_P_btm.n542 0.109875
R36415 C10_P_btm.n3123 C10_P_btm.n542 0.109875
R36416 C10_P_btm.n3124 C10_P_btm.n541 0.109875
R36417 C10_P_btm.n3126 C10_P_btm.n541 0.109875
R36418 C10_P_btm.n3127 C10_P_btm.n540 0.109875
R36419 C10_P_btm.n3129 C10_P_btm.n540 0.109875
R36420 C10_P_btm.n3130 C10_P_btm.n539 0.109875
R36421 C10_P_btm.n3132 C10_P_btm.n539 0.109875
R36422 C10_P_btm.n3133 C10_P_btm.n538 0.109875
R36423 C10_P_btm.n3135 C10_P_btm.n538 0.109875
R36424 C10_P_btm.n3136 C10_P_btm.n537 0.109875
R36425 C10_P_btm.n3138 C10_P_btm.n537 0.109875
R36426 C10_P_btm.n3139 C10_P_btm.n536 0.109875
R36427 C10_P_btm.n3141 C10_P_btm.n536 0.109875
R36428 C10_P_btm.n3142 C10_P_btm.n535 0.109875
R36429 C10_P_btm.n3144 C10_P_btm.n535 0.109875
R36430 C10_P_btm.n3145 C10_P_btm.n534 0.109875
R36431 C10_P_btm.n3147 C10_P_btm.n534 0.109875
R36432 C10_P_btm.n3148 C10_P_btm.n533 0.109875
R36433 C10_P_btm.n3150 C10_P_btm.n533 0.109875
R36434 C10_P_btm.n3151 C10_P_btm.n532 0.109875
R36435 C10_P_btm.n3153 C10_P_btm.n532 0.109875
R36436 C10_P_btm.n3154 C10_P_btm.n531 0.109875
R36437 C10_P_btm.n3156 C10_P_btm.n531 0.109875
R36438 C10_P_btm.n3157 C10_P_btm.n530 0.109875
R36439 C10_P_btm.n3159 C10_P_btm.n530 0.109875
R36440 C10_P_btm.n3160 C10_P_btm.n529 0.109875
R36441 C10_P_btm.n3162 C10_P_btm.n529 0.109875
R36442 C10_P_btm.n3163 C10_P_btm.n528 0.109875
R36443 C10_P_btm.n3165 C10_P_btm.n528 0.109875
R36444 C10_P_btm.n3166 C10_P_btm.n527 0.109875
R36445 C10_P_btm.n3168 C10_P_btm.n527 0.109875
R36446 C10_P_btm.n3169 C10_P_btm.n526 0.109875
R36447 C10_P_btm.n3171 C10_P_btm.n526 0.109875
R36448 C10_P_btm.n3172 C10_P_btm.n525 0.109875
R36449 C10_P_btm.n3174 C10_P_btm.n525 0.109875
R36450 C10_P_btm.n3175 C10_P_btm.n524 0.109875
R36451 C10_P_btm.n3177 C10_P_btm.n524 0.109875
R36452 C10_P_btm.n3178 C10_P_btm.n523 0.109875
R36453 C10_P_btm.n3180 C10_P_btm.n523 0.109875
R36454 C10_P_btm.n3181 C10_P_btm.n522 0.109875
R36455 C10_P_btm.n3183 C10_P_btm.n522 0.109875
R36456 C10_P_btm.n3184 C10_P_btm.n521 0.109875
R36457 C10_P_btm.n3186 C10_P_btm.n521 0.109875
R36458 C10_P_btm.n3187 C10_P_btm.n520 0.109875
R36459 C10_P_btm.n3189 C10_P_btm.n520 0.109875
R36460 C10_P_btm.n3190 C10_P_btm.n519 0.109875
R36461 C10_P_btm.n3192 C10_P_btm.n519 0.109875
R36462 C10_P_btm.n3193 C10_P_btm.n518 0.109875
R36463 C10_P_btm.n3195 C10_P_btm.n518 0.109875
R36464 C10_P_btm.n3196 C10_P_btm.n517 0.109875
R36465 C10_P_btm.n3198 C10_P_btm.n517 0.109875
R36466 C10_P_btm.n3199 C10_P_btm.n516 0.109875
R36467 C10_P_btm.n3201 C10_P_btm.n516 0.109875
R36468 C10_P_btm.n3202 C10_P_btm.n515 0.109875
R36469 C10_P_btm.n3204 C10_P_btm.n515 0.109875
R36470 C10_P_btm.n3205 C10_P_btm.n514 0.109875
R36471 C10_P_btm.n3207 C10_P_btm.n514 0.109875
R36472 C10_P_btm.n3208 C10_P_btm.n513 0.109875
R36473 C10_P_btm.n3210 C10_P_btm.n513 0.109875
R36474 C10_P_btm.n3211 C10_P_btm.n512 0.109875
R36475 C10_P_btm.n3213 C10_P_btm.n512 0.109875
R36476 C10_P_btm.n3214 C10_P_btm.n511 0.109875
R36477 C10_P_btm.n3216 C10_P_btm.n511 0.109875
R36478 C10_P_btm.n3217 C10_P_btm.n510 0.109875
R36479 C10_P_btm.n3219 C10_P_btm.n510 0.109875
R36480 C10_P_btm.n3220 C10_P_btm.n509 0.109875
R36481 C10_P_btm.n3222 C10_P_btm.n509 0.109875
R36482 C10_P_btm.n3223 C10_P_btm.n508 0.109875
R36483 C10_P_btm.n3225 C10_P_btm.n508 0.109875
R36484 C10_P_btm.n3226 C10_P_btm.n507 0.109875
R36485 C10_P_btm.n3228 C10_P_btm.n507 0.109875
R36486 C10_P_btm.n3229 C10_P_btm.n422 0.109875
R36487 C10_P_btm.n3231 C10_P_btm.n422 0.109875
R36488 C10_P_btm.n3232 C10_P_btm.n421 0.109875
R36489 C10_P_btm.n3234 C10_P_btm.n421 0.109875
R36490 C10_P_btm.n3235 C10_P_btm.n420 0.109875
R36491 C10_P_btm.n3237 C10_P_btm.n420 0.109875
R36492 C10_P_btm.n3238 C10_P_btm.n419 0.109875
R36493 C10_P_btm.n3240 C10_P_btm.n419 0.109875
R36494 C10_P_btm.n3241 C10_P_btm.n418 0.109875
R36495 C10_P_btm.n3243 C10_P_btm.n418 0.109875
R36496 C10_P_btm.n3244 C10_P_btm.n417 0.109875
R36497 C10_P_btm.n3246 C10_P_btm.n417 0.109875
R36498 C10_P_btm.n3247 C10_P_btm.n416 0.109875
R36499 C10_P_btm.n3249 C10_P_btm.n416 0.109875
R36500 C10_P_btm.n3250 C10_P_btm.n415 0.109875
R36501 C10_P_btm.n3252 C10_P_btm.n415 0.109875
R36502 C10_P_btm.n3253 C10_P_btm.n414 0.109875
R36503 C10_P_btm.n3255 C10_P_btm.n414 0.109875
R36504 C10_P_btm.n3256 C10_P_btm.n413 0.109875
R36505 C10_P_btm.n3258 C10_P_btm.n413 0.109875
R36506 C10_P_btm.n3259 C10_P_btm.n412 0.109875
R36507 C10_P_btm.n3261 C10_P_btm.n412 0.109875
R36508 C10_P_btm.n3262 C10_P_btm.n411 0.109875
R36509 C10_P_btm.n3264 C10_P_btm.n411 0.109875
R36510 C10_P_btm.n3265 C10_P_btm.n410 0.109875
R36511 C10_P_btm.n3267 C10_P_btm.n410 0.109875
R36512 C10_P_btm.n3268 C10_P_btm.n409 0.109875
R36513 C10_P_btm.n3270 C10_P_btm.n409 0.109875
R36514 C10_P_btm.n3271 C10_P_btm.n408 0.109875
R36515 C10_P_btm.n3273 C10_P_btm.n408 0.109875
R36516 C10_P_btm.n3274 C10_P_btm.n407 0.109875
R36517 C10_P_btm.n3276 C10_P_btm.n407 0.109875
R36518 C10_P_btm.n3277 C10_P_btm.n406 0.109875
R36519 C10_P_btm.n3279 C10_P_btm.n406 0.109875
R36520 C10_P_btm.n3280 C10_P_btm.n405 0.109875
R36521 C10_P_btm.n3282 C10_P_btm.n405 0.109875
R36522 C10_P_btm.n3283 C10_P_btm.n404 0.109875
R36523 C10_P_btm.n3285 C10_P_btm.n404 0.109875
R36524 C10_P_btm.n3286 C10_P_btm.n403 0.109875
R36525 C10_P_btm.n3288 C10_P_btm.n403 0.109875
R36526 C10_P_btm.n3289 C10_P_btm.n402 0.109875
R36527 C10_P_btm.n3291 C10_P_btm.n402 0.109875
R36528 C10_P_btm.n3292 C10_P_btm.n399 0.109875
R36529 C10_P_btm.n3294 C10_P_btm.n399 0.109875
R36530 C10_P_btm.n3301 C10_P_btm.n400 0.109875
R36531 C10_P_btm.n3301 C10_P_btm.n3300 0.109875
R36532 C10_P_btm.n445 C10_P_btm.n442 0.109875
R36533 C10_P_btm.n443 C10_P_btm.n442 0.109875
R36534 C10_P_btm.n448 C10_P_btm.n441 0.109875
R36535 C10_P_btm.n446 C10_P_btm.n441 0.109875
R36536 C10_P_btm.n451 C10_P_btm.n440 0.109875
R36537 C10_P_btm.n449 C10_P_btm.n440 0.109875
R36538 C10_P_btm.n454 C10_P_btm.n439 0.109875
R36539 C10_P_btm.n452 C10_P_btm.n439 0.109875
R36540 C10_P_btm.n457 C10_P_btm.n438 0.109875
R36541 C10_P_btm.n455 C10_P_btm.n438 0.109875
R36542 C10_P_btm.n460 C10_P_btm.n437 0.109875
R36543 C10_P_btm.n458 C10_P_btm.n437 0.109875
R36544 C10_P_btm.n463 C10_P_btm.n436 0.109875
R36545 C10_P_btm.n461 C10_P_btm.n436 0.109875
R36546 C10_P_btm.n466 C10_P_btm.n435 0.109875
R36547 C10_P_btm.n464 C10_P_btm.n435 0.109875
R36548 C10_P_btm.n469 C10_P_btm.n390 0.109875
R36549 C10_P_btm.n467 C10_P_btm.n390 0.109875
R36550 C10_P_btm.n3330 C10_P_btm.n391 0.109875
R36551 C10_P_btm.n3328 C10_P_btm.n391 0.109875
R36552 C10_P_btm.n3327 C10_P_btm.n392 0.109875
R36553 C10_P_btm.n3325 C10_P_btm.n392 0.109875
R36554 C10_P_btm.n3324 C10_P_btm.n393 0.109875
R36555 C10_P_btm.n3322 C10_P_btm.n393 0.109875
R36556 C10_P_btm.n3321 C10_P_btm.n394 0.109875
R36557 C10_P_btm.n3319 C10_P_btm.n394 0.109875
R36558 C10_P_btm.n3318 C10_P_btm.n395 0.109875
R36559 C10_P_btm.n3316 C10_P_btm.n395 0.109875
R36560 C10_P_btm.n3315 C10_P_btm.n396 0.109875
R36561 C10_P_btm.n3313 C10_P_btm.n396 0.109875
R36562 C10_P_btm.n3312 C10_P_btm.n397 0.109875
R36563 C10_P_btm.n3310 C10_P_btm.n397 0.109875
R36564 C10_P_btm.n3309 C10_P_btm.n398 0.109875
R36565 C10_P_btm.n3307 C10_P_btm.n398 0.109875
R36566 C10_P_btm.n3306 C10_P_btm.n3302 0.109875
R36567 C10_P_btm.n3304 C10_P_btm.n3302 0.109875
R36568 C10_P_btm.n3359 C10_P_btm.n346 0.109875
R36569 C10_P_btm.n3361 C10_P_btm.n346 0.109875
R36570 C10_P_btm.n3356 C10_P_btm.n349 0.109875
R36571 C10_P_btm.n3358 C10_P_btm.n349 0.109875
R36572 C10_P_btm.n3353 C10_P_btm.n350 0.109875
R36573 C10_P_btm.n3355 C10_P_btm.n350 0.109875
R36574 C10_P_btm.n3350 C10_P_btm.n351 0.109875
R36575 C10_P_btm.n3352 C10_P_btm.n351 0.109875
R36576 C10_P_btm.n3347 C10_P_btm.n352 0.109875
R36577 C10_P_btm.n3349 C10_P_btm.n352 0.109875
R36578 C10_P_btm.n3344 C10_P_btm.n353 0.109875
R36579 C10_P_btm.n3346 C10_P_btm.n353 0.109875
R36580 C10_P_btm.n3341 C10_P_btm.n354 0.109875
R36581 C10_P_btm.n3343 C10_P_btm.n354 0.109875
R36582 C10_P_btm.n3338 C10_P_btm.n355 0.109875
R36583 C10_P_btm.n3340 C10_P_btm.n355 0.109875
R36584 C10_P_btm.n3335 C10_P_btm.n389 0.109875
R36585 C10_P_btm.n3337 C10_P_btm.n389 0.109875
R36586 C10_P_btm.n388 C10_P_btm.n357 0.109875
R36587 C10_P_btm.n388 C10_P_btm.n387 0.109875
R36588 C10_P_btm.n385 C10_P_btm.n358 0.109875
R36589 C10_P_btm.n383 C10_P_btm.n358 0.109875
R36590 C10_P_btm.n382 C10_P_btm.n359 0.109875
R36591 C10_P_btm.n380 C10_P_btm.n359 0.109875
R36592 C10_P_btm.n379 C10_P_btm.n360 0.109875
R36593 C10_P_btm.n377 C10_P_btm.n360 0.109875
R36594 C10_P_btm.n376 C10_P_btm.n361 0.109875
R36595 C10_P_btm.n374 C10_P_btm.n361 0.109875
R36596 C10_P_btm.n373 C10_P_btm.n362 0.109875
R36597 C10_P_btm.n371 C10_P_btm.n362 0.109875
R36598 C10_P_btm.n370 C10_P_btm.n363 0.109875
R36599 C10_P_btm.n368 C10_P_btm.n363 0.109875
R36600 C10_P_btm.n367 C10_P_btm.n364 0.109875
R36601 C10_P_btm.n365 C10_P_btm.n364 0.109875
R36602 C10_P_btm.n3368 C10_P_btm.n347 0.109875
R36603 C10_P_btm.n3368 C10_P_btm.n3367 0.109875
R36604 C10_P_btm.n3373 C10_P_btm.n3369 0.109875
R36605 C10_P_btm.n3371 C10_P_btm.n3369 0.109875
R36606 C10_P_btm.n3376 C10_P_btm.n345 0.109875
R36607 C10_P_btm.n3374 C10_P_btm.n345 0.109875
R36608 C10_P_btm.n3379 C10_P_btm.n344 0.109875
R36609 C10_P_btm.n3377 C10_P_btm.n344 0.109875
R36610 C10_P_btm.n3382 C10_P_btm.n343 0.109875
R36611 C10_P_btm.n3380 C10_P_btm.n343 0.109875
R36612 C10_P_btm.n3385 C10_P_btm.n342 0.109875
R36613 C10_P_btm.n3383 C10_P_btm.n342 0.109875
R36614 C10_P_btm.n3388 C10_P_btm.n341 0.109875
R36615 C10_P_btm.n3386 C10_P_btm.n341 0.109875
R36616 C10_P_btm.n3391 C10_P_btm.n340 0.109875
R36617 C10_P_btm.n3389 C10_P_btm.n340 0.109875
R36618 C10_P_btm.n3394 C10_P_btm.n339 0.109875
R36619 C10_P_btm.n3392 C10_P_btm.n339 0.109875
R36620 C10_P_btm.n3397 C10_P_btm.n338 0.109875
R36621 C10_P_btm.n3395 C10_P_btm.n338 0.109875
R36622 C10_P_btm.n3402 C10_P_btm.n336 0.109875
R36623 C10_P_btm.n3404 C10_P_btm.n336 0.109875
R36624 C10_P_btm.n3405 C10_P_btm.n302 0.109875
R36625 C10_P_btm.n3407 C10_P_btm.n302 0.109875
R36626 C10_P_btm.n3408 C10_P_btm.n301 0.109875
R36627 C10_P_btm.n3410 C10_P_btm.n301 0.109875
R36628 C10_P_btm.n3411 C10_P_btm.n300 0.109875
R36629 C10_P_btm.n3413 C10_P_btm.n300 0.109875
R36630 C10_P_btm.n3414 C10_P_btm.n299 0.109875
R36631 C10_P_btm.n3416 C10_P_btm.n299 0.109875
R36632 C10_P_btm.n3417 C10_P_btm.n298 0.109875
R36633 C10_P_btm.n3419 C10_P_btm.n298 0.109875
R36634 C10_P_btm.n3420 C10_P_btm.n297 0.109875
R36635 C10_P_btm.n3422 C10_P_btm.n297 0.109875
R36636 C10_P_btm.n3423 C10_P_btm.n296 0.109875
R36637 C10_P_btm.n3425 C10_P_btm.n296 0.109875
R36638 C10_P_btm.n3426 C10_P_btm.n293 0.109875
R36639 C10_P_btm.n3428 C10_P_btm.n293 0.109875
R36640 C10_P_btm.n3435 C10_P_btm.n294 0.109875
R36641 C10_P_btm.n3435 C10_P_btm.n3434 0.109875
R36642 C10_P_btm.n314 C10_P_btm.n311 0.109875
R36643 C10_P_btm.n312 C10_P_btm.n311 0.109875
R36644 C10_P_btm.n317 C10_P_btm.n310 0.109875
R36645 C10_P_btm.n315 C10_P_btm.n310 0.109875
R36646 C10_P_btm.n320 C10_P_btm.n309 0.109875
R36647 C10_P_btm.n318 C10_P_btm.n309 0.109875
R36648 C10_P_btm.n323 C10_P_btm.n308 0.109875
R36649 C10_P_btm.n321 C10_P_btm.n308 0.109875
R36650 C10_P_btm.n326 C10_P_btm.n307 0.109875
R36651 C10_P_btm.n324 C10_P_btm.n307 0.109875
R36652 C10_P_btm.n329 C10_P_btm.n306 0.109875
R36653 C10_P_btm.n327 C10_P_btm.n306 0.109875
R36654 C10_P_btm.n332 C10_P_btm.n305 0.109875
R36655 C10_P_btm.n330 C10_P_btm.n305 0.109875
R36656 C10_P_btm.n335 C10_P_btm.n304 0.109875
R36657 C10_P_btm.n335 C10_P_btm.n334 0.109875
R36658 C10_P_btm.n3464 C10_P_btm.n285 0.109875
R36659 C10_P_btm.n3462 C10_P_btm.n285 0.109875
R36660 C10_P_btm.n3461 C10_P_btm.n286 0.109875
R36661 C10_P_btm.n3459 C10_P_btm.n286 0.109875
R36662 C10_P_btm.n3458 C10_P_btm.n287 0.109875
R36663 C10_P_btm.n3456 C10_P_btm.n287 0.109875
R36664 C10_P_btm.n3455 C10_P_btm.n288 0.109875
R36665 C10_P_btm.n3453 C10_P_btm.n288 0.109875
R36666 C10_P_btm.n3452 C10_P_btm.n289 0.109875
R36667 C10_P_btm.n3450 C10_P_btm.n289 0.109875
R36668 C10_P_btm.n3449 C10_P_btm.n290 0.109875
R36669 C10_P_btm.n3447 C10_P_btm.n290 0.109875
R36670 C10_P_btm.n3446 C10_P_btm.n291 0.109875
R36671 C10_P_btm.n3444 C10_P_btm.n291 0.109875
R36672 C10_P_btm.n3443 C10_P_btm.n292 0.109875
R36673 C10_P_btm.n3441 C10_P_btm.n292 0.109875
R36674 C10_P_btm.n3440 C10_P_btm.n3436 0.109875
R36675 C10_P_btm.n3438 C10_P_btm.n3436 0.109875
R36676 C10_P_btm.n3493 C10_P_btm.n240 0.109875
R36677 C10_P_btm.n3495 C10_P_btm.n240 0.109875
R36678 C10_P_btm.n3490 C10_P_btm.n243 0.109875
R36679 C10_P_btm.n3492 C10_P_btm.n243 0.109875
R36680 C10_P_btm.n3487 C10_P_btm.n244 0.109875
R36681 C10_P_btm.n3489 C10_P_btm.n244 0.109875
R36682 C10_P_btm.n3484 C10_P_btm.n245 0.109875
R36683 C10_P_btm.n3486 C10_P_btm.n245 0.109875
R36684 C10_P_btm.n3481 C10_P_btm.n246 0.109875
R36685 C10_P_btm.n3483 C10_P_btm.n246 0.109875
R36686 C10_P_btm.n3478 C10_P_btm.n247 0.109875
R36687 C10_P_btm.n3480 C10_P_btm.n247 0.109875
R36688 C10_P_btm.n3475 C10_P_btm.n248 0.109875
R36689 C10_P_btm.n3477 C10_P_btm.n248 0.109875
R36690 C10_P_btm.n3472 C10_P_btm.n249 0.109875
R36691 C10_P_btm.n3474 C10_P_btm.n249 0.109875
R36692 C10_P_btm.n3469 C10_P_btm.n283 0.109875
R36693 C10_P_btm.n3471 C10_P_btm.n283 0.109875
R36694 C10_P_btm.n282 C10_P_btm.n251 0.109875
R36695 C10_P_btm.n282 C10_P_btm.n281 0.109875
R36696 C10_P_btm.n279 C10_P_btm.n252 0.109875
R36697 C10_P_btm.n277 C10_P_btm.n252 0.109875
R36698 C10_P_btm.n276 C10_P_btm.n253 0.109875
R36699 C10_P_btm.n274 C10_P_btm.n253 0.109875
R36700 C10_P_btm.n273 C10_P_btm.n254 0.109875
R36701 C10_P_btm.n271 C10_P_btm.n254 0.109875
R36702 C10_P_btm.n270 C10_P_btm.n255 0.109875
R36703 C10_P_btm.n268 C10_P_btm.n255 0.109875
R36704 C10_P_btm.n267 C10_P_btm.n256 0.109875
R36705 C10_P_btm.n265 C10_P_btm.n256 0.109875
R36706 C10_P_btm.n264 C10_P_btm.n257 0.109875
R36707 C10_P_btm.n262 C10_P_btm.n257 0.109875
R36708 C10_P_btm.n261 C10_P_btm.n258 0.109875
R36709 C10_P_btm.n259 C10_P_btm.n258 0.109875
R36710 C10_P_btm.n3502 C10_P_btm.n241 0.109875
R36711 C10_P_btm.n3502 C10_P_btm.n3501 0.109875
R36712 C10_P_btm.n3507 C10_P_btm.n3503 0.109875
R36713 C10_P_btm.n3505 C10_P_btm.n3503 0.109875
R36714 C10_P_btm.n3510 C10_P_btm.n239 0.109875
R36715 C10_P_btm.n3508 C10_P_btm.n239 0.109875
R36716 C10_P_btm.n3513 C10_P_btm.n238 0.109875
R36717 C10_P_btm.n3511 C10_P_btm.n238 0.109875
R36718 C10_P_btm.n3516 C10_P_btm.n237 0.109875
R36719 C10_P_btm.n3514 C10_P_btm.n237 0.109875
R36720 C10_P_btm.n3519 C10_P_btm.n236 0.109875
R36721 C10_P_btm.n3517 C10_P_btm.n236 0.109875
R36722 C10_P_btm.n3522 C10_P_btm.n235 0.109875
R36723 C10_P_btm.n3520 C10_P_btm.n235 0.109875
R36724 C10_P_btm.n3525 C10_P_btm.n234 0.109875
R36725 C10_P_btm.n3523 C10_P_btm.n234 0.109875
R36726 C10_P_btm.n3528 C10_P_btm.n233 0.109875
R36727 C10_P_btm.n3526 C10_P_btm.n233 0.109875
R36728 C10_P_btm.n3531 C10_P_btm.n232 0.109875
R36729 C10_P_btm.n3529 C10_P_btm.n232 0.109875
R36730 C10_P_btm.n3536 C10_P_btm.n230 0.109875
R36731 C10_P_btm.n3538 C10_P_btm.n230 0.109875
R36732 C10_P_btm.n3539 C10_P_btm.n196 0.109875
R36733 C10_P_btm.n3541 C10_P_btm.n196 0.109875
R36734 C10_P_btm.n3542 C10_P_btm.n195 0.109875
R36735 C10_P_btm.n3544 C10_P_btm.n195 0.109875
R36736 C10_P_btm.n3545 C10_P_btm.n194 0.109875
R36737 C10_P_btm.n3547 C10_P_btm.n194 0.109875
R36738 C10_P_btm.n3548 C10_P_btm.n193 0.109875
R36739 C10_P_btm.n3550 C10_P_btm.n193 0.109875
R36740 C10_P_btm.n3551 C10_P_btm.n192 0.109875
R36741 C10_P_btm.n3553 C10_P_btm.n192 0.109875
R36742 C10_P_btm.n3554 C10_P_btm.n191 0.109875
R36743 C10_P_btm.n3556 C10_P_btm.n191 0.109875
R36744 C10_P_btm.n3557 C10_P_btm.n190 0.109875
R36745 C10_P_btm.n3559 C10_P_btm.n190 0.109875
R36746 C10_P_btm.n3560 C10_P_btm.n187 0.109875
R36747 C10_P_btm.n3562 C10_P_btm.n187 0.109875
R36748 C10_P_btm.n3569 C10_P_btm.n188 0.109875
R36749 C10_P_btm.n3569 C10_P_btm.n3568 0.109875
R36750 C10_P_btm.n208 C10_P_btm.n205 0.109875
R36751 C10_P_btm.n206 C10_P_btm.n205 0.109875
R36752 C10_P_btm.n211 C10_P_btm.n204 0.109875
R36753 C10_P_btm.n209 C10_P_btm.n204 0.109875
R36754 C10_P_btm.n214 C10_P_btm.n203 0.109875
R36755 C10_P_btm.n212 C10_P_btm.n203 0.109875
R36756 C10_P_btm.n217 C10_P_btm.n202 0.109875
R36757 C10_P_btm.n215 C10_P_btm.n202 0.109875
R36758 C10_P_btm.n220 C10_P_btm.n201 0.109875
R36759 C10_P_btm.n218 C10_P_btm.n201 0.109875
R36760 C10_P_btm.n223 C10_P_btm.n200 0.109875
R36761 C10_P_btm.n221 C10_P_btm.n200 0.109875
R36762 C10_P_btm.n226 C10_P_btm.n199 0.109875
R36763 C10_P_btm.n224 C10_P_btm.n199 0.109875
R36764 C10_P_btm.n229 C10_P_btm.n198 0.109875
R36765 C10_P_btm.n229 C10_P_btm.n228 0.109875
R36766 C10_P_btm.n3598 C10_P_btm.n179 0.109875
R36767 C10_P_btm.n3596 C10_P_btm.n179 0.109875
R36768 C10_P_btm.n3595 C10_P_btm.n180 0.109875
R36769 C10_P_btm.n3593 C10_P_btm.n180 0.109875
R36770 C10_P_btm.n3592 C10_P_btm.n181 0.109875
R36771 C10_P_btm.n3590 C10_P_btm.n181 0.109875
R36772 C10_P_btm.n3589 C10_P_btm.n182 0.109875
R36773 C10_P_btm.n3587 C10_P_btm.n182 0.109875
R36774 C10_P_btm.n3586 C10_P_btm.n183 0.109875
R36775 C10_P_btm.n3584 C10_P_btm.n183 0.109875
R36776 C10_P_btm.n3583 C10_P_btm.n184 0.109875
R36777 C10_P_btm.n3581 C10_P_btm.n184 0.109875
R36778 C10_P_btm.n3580 C10_P_btm.n185 0.109875
R36779 C10_P_btm.n3578 C10_P_btm.n185 0.109875
R36780 C10_P_btm.n3577 C10_P_btm.n186 0.109875
R36781 C10_P_btm.n3575 C10_P_btm.n186 0.109875
R36782 C10_P_btm.n3574 C10_P_btm.n3570 0.109875
R36783 C10_P_btm.n3572 C10_P_btm.n3570 0.109875
R36784 C10_P_btm.n3627 C10_P_btm.n134 0.109875
R36785 C10_P_btm.n3629 C10_P_btm.n134 0.109875
R36786 C10_P_btm.n3624 C10_P_btm.n137 0.109875
R36787 C10_P_btm.n3626 C10_P_btm.n137 0.109875
R36788 C10_P_btm.n3621 C10_P_btm.n138 0.109875
R36789 C10_P_btm.n3623 C10_P_btm.n138 0.109875
R36790 C10_P_btm.n3618 C10_P_btm.n139 0.109875
R36791 C10_P_btm.n3620 C10_P_btm.n139 0.109875
R36792 C10_P_btm.n3615 C10_P_btm.n140 0.109875
R36793 C10_P_btm.n3617 C10_P_btm.n140 0.109875
R36794 C10_P_btm.n3612 C10_P_btm.n141 0.109875
R36795 C10_P_btm.n3614 C10_P_btm.n141 0.109875
R36796 C10_P_btm.n3609 C10_P_btm.n142 0.109875
R36797 C10_P_btm.n3611 C10_P_btm.n142 0.109875
R36798 C10_P_btm.n3606 C10_P_btm.n143 0.109875
R36799 C10_P_btm.n3608 C10_P_btm.n143 0.109875
R36800 C10_P_btm.n3603 C10_P_btm.n177 0.109875
R36801 C10_P_btm.n3605 C10_P_btm.n177 0.109875
R36802 C10_P_btm.n176 C10_P_btm.n145 0.109875
R36803 C10_P_btm.n176 C10_P_btm.n175 0.109875
R36804 C10_P_btm.n173 C10_P_btm.n146 0.109875
R36805 C10_P_btm.n171 C10_P_btm.n146 0.109875
R36806 C10_P_btm.n170 C10_P_btm.n147 0.109875
R36807 C10_P_btm.n168 C10_P_btm.n147 0.109875
R36808 C10_P_btm.n167 C10_P_btm.n148 0.109875
R36809 C10_P_btm.n165 C10_P_btm.n148 0.109875
R36810 C10_P_btm.n164 C10_P_btm.n149 0.109875
R36811 C10_P_btm.n162 C10_P_btm.n149 0.109875
R36812 C10_P_btm.n161 C10_P_btm.n150 0.109875
R36813 C10_P_btm.n159 C10_P_btm.n150 0.109875
R36814 C10_P_btm.n158 C10_P_btm.n151 0.109875
R36815 C10_P_btm.n156 C10_P_btm.n151 0.109875
R36816 C10_P_btm.n155 C10_P_btm.n152 0.109875
R36817 C10_P_btm.n153 C10_P_btm.n152 0.109875
R36818 C10_P_btm.n3636 C10_P_btm.n135 0.109875
R36819 C10_P_btm.n3636 C10_P_btm.n3635 0.109875
R36820 C10_P_btm.n3641 C10_P_btm.n3637 0.109875
R36821 C10_P_btm.n3639 C10_P_btm.n3637 0.109875
R36822 C10_P_btm.n3644 C10_P_btm.n133 0.109875
R36823 C10_P_btm.n3642 C10_P_btm.n133 0.109875
R36824 C10_P_btm.n3647 C10_P_btm.n132 0.109875
R36825 C10_P_btm.n3645 C10_P_btm.n132 0.109875
R36826 C10_P_btm.n3650 C10_P_btm.n131 0.109875
R36827 C10_P_btm.n3648 C10_P_btm.n131 0.109875
R36828 C10_P_btm.n3653 C10_P_btm.n130 0.109875
R36829 C10_P_btm.n3651 C10_P_btm.n130 0.109875
R36830 C10_P_btm.n3656 C10_P_btm.n129 0.109875
R36831 C10_P_btm.n3654 C10_P_btm.n129 0.109875
R36832 C10_P_btm.n3659 C10_P_btm.n128 0.109875
R36833 C10_P_btm.n3657 C10_P_btm.n128 0.109875
R36834 C10_P_btm.n3662 C10_P_btm.n127 0.109875
R36835 C10_P_btm.n3660 C10_P_btm.n127 0.109875
R36836 C10_P_btm.n3665 C10_P_btm.n126 0.109875
R36837 C10_P_btm.n3663 C10_P_btm.n126 0.109875
R36838 C10_P_btm.n3670 C10_P_btm.n124 0.109875
R36839 C10_P_btm.n3672 C10_P_btm.n124 0.109875
R36840 C10_P_btm.n3673 C10_P_btm.n90 0.109875
R36841 C10_P_btm.n3675 C10_P_btm.n90 0.109875
R36842 C10_P_btm.n3676 C10_P_btm.n89 0.109875
R36843 C10_P_btm.n3678 C10_P_btm.n89 0.109875
R36844 C10_P_btm.n3679 C10_P_btm.n88 0.109875
R36845 C10_P_btm.n3681 C10_P_btm.n88 0.109875
R36846 C10_P_btm.n3682 C10_P_btm.n87 0.109875
R36847 C10_P_btm.n3684 C10_P_btm.n87 0.109875
R36848 C10_P_btm.n3685 C10_P_btm.n86 0.109875
R36849 C10_P_btm.n3687 C10_P_btm.n86 0.109875
R36850 C10_P_btm.n3688 C10_P_btm.n85 0.109875
R36851 C10_P_btm.n3690 C10_P_btm.n85 0.109875
R36852 C10_P_btm.n3691 C10_P_btm.n84 0.109875
R36853 C10_P_btm.n3693 C10_P_btm.n84 0.109875
R36854 C10_P_btm.n3694 C10_P_btm.n81 0.109875
R36855 C10_P_btm.n3696 C10_P_btm.n81 0.109875
R36856 C10_P_btm.n3703 C10_P_btm.n82 0.109875
R36857 C10_P_btm.n3703 C10_P_btm.n3702 0.109875
R36858 C10_P_btm.n102 C10_P_btm.n99 0.109875
R36859 C10_P_btm.n100 C10_P_btm.n99 0.109875
R36860 C10_P_btm.n105 C10_P_btm.n98 0.109875
R36861 C10_P_btm.n103 C10_P_btm.n98 0.109875
R36862 C10_P_btm.n108 C10_P_btm.n97 0.109875
R36863 C10_P_btm.n106 C10_P_btm.n97 0.109875
R36864 C10_P_btm.n111 C10_P_btm.n96 0.109875
R36865 C10_P_btm.n109 C10_P_btm.n96 0.109875
R36866 C10_P_btm.n114 C10_P_btm.n95 0.109875
R36867 C10_P_btm.n112 C10_P_btm.n95 0.109875
R36868 C10_P_btm.n117 C10_P_btm.n94 0.109875
R36869 C10_P_btm.n115 C10_P_btm.n94 0.109875
R36870 C10_P_btm.n120 C10_P_btm.n93 0.109875
R36871 C10_P_btm.n118 C10_P_btm.n93 0.109875
R36872 C10_P_btm.n123 C10_P_btm.n92 0.109875
R36873 C10_P_btm.n123 C10_P_btm.n122 0.109875
R36874 C10_P_btm.n3732 C10_P_btm.n73 0.109875
R36875 C10_P_btm.n3730 C10_P_btm.n73 0.109875
R36876 C10_P_btm.n3729 C10_P_btm.n74 0.109875
R36877 C10_P_btm.n3727 C10_P_btm.n74 0.109875
R36878 C10_P_btm.n3726 C10_P_btm.n75 0.109875
R36879 C10_P_btm.n3724 C10_P_btm.n75 0.109875
R36880 C10_P_btm.n3723 C10_P_btm.n76 0.109875
R36881 C10_P_btm.n3721 C10_P_btm.n76 0.109875
R36882 C10_P_btm.n3720 C10_P_btm.n77 0.109875
R36883 C10_P_btm.n3718 C10_P_btm.n77 0.109875
R36884 C10_P_btm.n3717 C10_P_btm.n78 0.109875
R36885 C10_P_btm.n3715 C10_P_btm.n78 0.109875
R36886 C10_P_btm.n3714 C10_P_btm.n79 0.109875
R36887 C10_P_btm.n3712 C10_P_btm.n79 0.109875
R36888 C10_P_btm.n3711 C10_P_btm.n80 0.109875
R36889 C10_P_btm.n3709 C10_P_btm.n80 0.109875
R36890 C10_P_btm.n3708 C10_P_btm.n3704 0.109875
R36891 C10_P_btm.n3706 C10_P_btm.n3704 0.109875
R36892 C10_P_btm.n3796 C10_P_btm.n61 0.109875
R36893 C10_P_btm.n3798 C10_P_btm.n61 0.109875
R36894 C10_P_btm.n3793 C10_P_btm.n64 0.109875
R36895 C10_P_btm.n3795 C10_P_btm.n64 0.109875
R36896 C10_P_btm.n3790 C10_P_btm.n65 0.109875
R36897 C10_P_btm.n3792 C10_P_btm.n65 0.109875
R36898 C10_P_btm.n3787 C10_P_btm.n66 0.109875
R36899 C10_P_btm.n3789 C10_P_btm.n66 0.109875
R36900 C10_P_btm.n3784 C10_P_btm.n67 0.109875
R36901 C10_P_btm.n3786 C10_P_btm.n67 0.109875
R36902 C10_P_btm.n3781 C10_P_btm.n68 0.109875
R36903 C10_P_btm.n3783 C10_P_btm.n68 0.109875
R36904 C10_P_btm.n3778 C10_P_btm.n69 0.109875
R36905 C10_P_btm.n3780 C10_P_btm.n69 0.109875
R36906 C10_P_btm.n3775 C10_P_btm.n70 0.109875
R36907 C10_P_btm.n3777 C10_P_btm.n70 0.109875
R36908 C10_P_btm.n3772 C10_P_btm.n71 0.109875
R36909 C10_P_btm.n3774 C10_P_btm.n71 0.109875
R36910 C10_P_btm.n3767 C10_P_btm.n52 0.109875
R36911 C10_P_btm.n3765 C10_P_btm.n52 0.109875
R36912 C10_P_btm.n3764 C10_P_btm.n3737 0.109875
R36913 C10_P_btm.n3762 C10_P_btm.n3737 0.109875
R36914 C10_P_btm.n3761 C10_P_btm.n3738 0.109875
R36915 C10_P_btm.n3759 C10_P_btm.n3738 0.109875
R36916 C10_P_btm.n3758 C10_P_btm.n3739 0.109875
R36917 C10_P_btm.n3756 C10_P_btm.n3739 0.109875
R36918 C10_P_btm.n3755 C10_P_btm.n3740 0.109875
R36919 C10_P_btm.n3753 C10_P_btm.n3740 0.109875
R36920 C10_P_btm.n3752 C10_P_btm.n3741 0.109875
R36921 C10_P_btm.n3750 C10_P_btm.n3741 0.109875
R36922 C10_P_btm.n3749 C10_P_btm.n3742 0.109875
R36923 C10_P_btm.n3747 C10_P_btm.n3742 0.109875
R36924 C10_P_btm.n3746 C10_P_btm.n3743 0.109875
R36925 C10_P_btm.n3744 C10_P_btm.n3743 0.109875
R36926 C10_P_btm.n3805 C10_P_btm.n62 0.109875
R36927 C10_P_btm.n3805 C10_P_btm.n3804 0.109875
R36928 C10_P_btm.n3810 C10_P_btm.n3806 0.109875
R36929 C10_P_btm.n3808 C10_P_btm.n3806 0.109875
R36930 C10_P_btm.n3813 C10_P_btm.n60 0.109875
R36931 C10_P_btm.n3811 C10_P_btm.n60 0.109875
R36932 C10_P_btm.n3816 C10_P_btm.n59 0.109875
R36933 C10_P_btm.n3814 C10_P_btm.n59 0.109875
R36934 C10_P_btm.n3819 C10_P_btm.n58 0.109875
R36935 C10_P_btm.n3817 C10_P_btm.n58 0.109875
R36936 C10_P_btm.n3822 C10_P_btm.n57 0.109875
R36937 C10_P_btm.n3820 C10_P_btm.n57 0.109875
R36938 C10_P_btm.n3825 C10_P_btm.n56 0.109875
R36939 C10_P_btm.n3823 C10_P_btm.n56 0.109875
R36940 C10_P_btm.n3828 C10_P_btm.n55 0.109875
R36941 C10_P_btm.n3826 C10_P_btm.n55 0.109875
R36942 C10_P_btm.n3831 C10_P_btm.n54 0.109875
R36943 C10_P_btm.n3829 C10_P_btm.n54 0.109875
R36944 C10_P_btm.n3834 C10_P_btm.n53 0.109875
R36945 C10_P_btm.n3834 C10_P_btm.n3833 0.109875
R36946 C10_P_btm.n3837 C10_P_btm.n3835 0.109875
R36947 C10_P_btm.n3839 C10_P_btm.n3835 0.109875
R36948 C10_P_btm.n3840 C10_P_btm.n51 0.109875
R36949 C10_P_btm.n3842 C10_P_btm.n51 0.109875
R36950 C10_P_btm.n3843 C10_P_btm.n50 0.109875
R36951 C10_P_btm.n3845 C10_P_btm.n50 0.109875
R36952 C10_P_btm.n3846 C10_P_btm.n49 0.109875
R36953 C10_P_btm.n3848 C10_P_btm.n49 0.109875
R36954 C10_P_btm.n3849 C10_P_btm.n48 0.109875
R36955 C10_P_btm.n3851 C10_P_btm.n48 0.109875
R36956 C10_P_btm.n3852 C10_P_btm.n47 0.109875
R36957 C10_P_btm.n3854 C10_P_btm.n47 0.109875
R36958 C10_P_btm.n3855 C10_P_btm.n46 0.109875
R36959 C10_P_btm.n3857 C10_P_btm.n46 0.109875
R36960 C10_P_btm.n3858 C10_P_btm.n45 0.109875
R36961 C10_P_btm.n3860 C10_P_btm.n45 0.109875
R36962 C10_P_btm.n3861 C10_P_btm.n44 0.109875
R36963 C10_P_btm.n3863 C10_P_btm.n44 0.109875
R36964 C10_P_btm.n3870 C10_P_btm.n42 0.109875
R36965 C10_P_btm.n3868 C10_P_btm.n42 0.109875
R36966 C10_P_btm.n3873 C10_P_btm.n41 0.109875
R36967 C10_P_btm.n3871 C10_P_btm.n41 0.109875
R36968 C10_P_btm.n3876 C10_P_btm.n40 0.109875
R36969 C10_P_btm.n3874 C10_P_btm.n40 0.109875
R36970 C10_P_btm.n3879 C10_P_btm.n39 0.109875
R36971 C10_P_btm.n3877 C10_P_btm.n39 0.109875
R36972 C10_P_btm.n3882 C10_P_btm.n38 0.109875
R36973 C10_P_btm.n3880 C10_P_btm.n38 0.109875
R36974 C10_P_btm.n3885 C10_P_btm.n37 0.109875
R36975 C10_P_btm.n3883 C10_P_btm.n37 0.109875
R36976 C10_P_btm.n3888 C10_P_btm.n36 0.109875
R36977 C10_P_btm.n3886 C10_P_btm.n36 0.109875
R36978 C10_P_btm.n3891 C10_P_btm.n35 0.109875
R36979 C10_P_btm.n3889 C10_P_btm.n35 0.109875
R36980 C10_P_btm.n3894 C10_P_btm.n34 0.109875
R36981 C10_P_btm.n3892 C10_P_btm.n34 0.109875
R36982 C10_P_btm.n2457 C10_P_btm.n2456 0.0556875
R36983 C10_P_btm.n2430 C10_P_btm.n2413 0.0556875
R36984 C10_P_btm.n2491 C10_P_btm.n2490 0.0556875
R36985 C10_P_btm.n2462 C10_P_btm.n2371 0.0556875
R36986 C10_P_btm.n2522 C10_P_btm.n2521 0.0556875
R36987 C10_P_btm.n2493 C10_P_btm.n2492 0.0556875
R36988 C10_P_btm.n2379 C10_P_btm.n2360 0.0556875
R36989 C10_P_btm.n2524 C10_P_btm.n2523 0.0556875
R36990 C10_P_btm.n2529 C10_P_btm.n2318 0.0556875
R36991 C10_P_btm.n2558 C10_P_btm.n2557 0.0556875
R36992 C10_P_btm.n2560 C10_P_btm.n2559 0.0556875
R36993 C10_P_btm.n2589 C10_P_btm.n2588 0.0556875
R36994 C10_P_btm.n2591 C10_P_btm.n2590 0.0556875
R36995 C10_P_btm.n2326 C10_P_btm.n2307 0.0556875
R36996 C10_P_btm.n2625 C10_P_btm.n2624 0.0556875
R36997 C10_P_btm.n2596 C10_P_btm.n2265 0.0556875
R36998 C10_P_btm.n2656 C10_P_btm.n2655 0.0556875
R36999 C10_P_btm.n2627 C10_P_btm.n2626 0.0556875
R37000 C10_P_btm.n2273 C10_P_btm.n2254 0.0556875
R37001 C10_P_btm.n2658 C10_P_btm.n2657 0.0556875
R37002 C10_P_btm.n2663 C10_P_btm.n2212 0.0556875
R37003 C10_P_btm.n2692 C10_P_btm.n2691 0.0556875
R37004 C10_P_btm.n2694 C10_P_btm.n2693 0.0556875
R37005 C10_P_btm.n2723 C10_P_btm.n2722 0.0556875
R37006 C10_P_btm.n2725 C10_P_btm.n2724 0.0556875
R37007 C10_P_btm.n2220 C10_P_btm.n2201 0.0556875
R37008 C10_P_btm.n2759 C10_P_btm.n2758 0.0556875
R37009 C10_P_btm.n2730 C10_P_btm.n2159 0.0556875
R37010 C10_P_btm.n2790 C10_P_btm.n2789 0.0556875
R37011 C10_P_btm.n2761 C10_P_btm.n2760 0.0556875
R37012 C10_P_btm.n2167 C10_P_btm.n2148 0.0556875
R37013 C10_P_btm.n2792 C10_P_btm.n2791 0.0556875
R37014 C10_P_btm.n2797 C10_P_btm.n2106 0.0556875
R37015 C10_P_btm.n2826 C10_P_btm.n2825 0.0556875
R37016 C10_P_btm.n2828 C10_P_btm.n2827 0.0556875
R37017 C10_P_btm.n2857 C10_P_btm.n2856 0.0556875
R37018 C10_P_btm.n2859 C10_P_btm.n2858 0.0556875
R37019 C10_P_btm.n2114 C10_P_btm.n2095 0.0556875
R37020 C10_P_btm.n2893 C10_P_btm.n2892 0.0556875
R37021 C10_P_btm.n2864 C10_P_btm.n2086 0.0556875
R37022 C10_P_btm.n2959 C10_P_btm.n2958 0.0556875
R37023 C10_P_btm.n2930 C10_P_btm.n2929 0.0556875
R37024 C10_P_btm.n2928 C10_P_btm.n2927 0.0556875
R37025 C10_P_btm.n2961 C10_P_btm.n2960 0.0556875
R37026 C10_P_btm.n2966 C10_P_btm.n2066 0.0556875
R37027 C10_P_btm.n2895 C10_P_btm.n2894 0.0556875
R37028 C10_P_btm.n2995 C10_P_btm.n2056 0.0556875
R37029 C10_P_btm.n3024 C10_P_btm.n3023 0.0556875
R37030 C10_P_btm.n3106 C10_P_btm.n3105 0.0556875
R37031 C10_P_btm.n1477 C10_P_btm.n1476 0.0556875
R37032 C10_P_btm.n1042 C10_P_btm.n918 0.0556875
R37033 C10_P_btm.n1670 C10_P_btm.n1669 0.0556875
R37034 C10_P_btm.n1482 C10_P_btm.n611 0.0556875
R37035 C10_P_btm.n1860 C10_P_btm.n1859 0.0556875
R37036 C10_P_btm.n1672 C10_P_btm.n1671 0.0556875
R37037 C10_P_btm.n672 C10_P_btm.n547 0.0556875
R37038 C10_P_btm.n1862 C10_P_btm.n1861 0.0556875
R37039 C10_P_btm.n1867 C10_P_btm.n401 0.0556875
R37040 C10_P_btm.n2055 C10_P_btm.n2054 0.0556875
R37041 C10_P_btm.n3108 C10_P_btm.n3107 0.0556875
R37042 C10_P_btm.n3296 C10_P_btm.n3295 0.0556875
R37043 C10_P_btm.n3298 C10_P_btm.n3297 0.0556875
R37044 C10_P_btm.n3332 C10_P_btm.n3331 0.0556875
R37045 C10_P_btm.n3303 C10_P_btm.n348 0.0556875
R37046 C10_P_btm.n3363 C10_P_btm.n3362 0.0556875
R37047 C10_P_btm.n3334 C10_P_btm.n3333 0.0556875
R37048 C10_P_btm.n356 C10_P_btm.n337 0.0556875
R37049 C10_P_btm.n3365 C10_P_btm.n3364 0.0556875
R37050 C10_P_btm.n3370 C10_P_btm.n295 0.0556875
R37051 C10_P_btm.n3399 C10_P_btm.n3398 0.0556875
R37052 C10_P_btm.n3401 C10_P_btm.n3400 0.0556875
R37053 C10_P_btm.n3430 C10_P_btm.n3429 0.0556875
R37054 C10_P_btm.n3432 C10_P_btm.n3431 0.0556875
R37055 C10_P_btm.n303 C10_P_btm.n284 0.0556875
R37056 C10_P_btm.n3466 C10_P_btm.n3465 0.0556875
R37057 C10_P_btm.n3437 C10_P_btm.n242 0.0556875
R37058 C10_P_btm.n3497 C10_P_btm.n3496 0.0556875
R37059 C10_P_btm.n3468 C10_P_btm.n3467 0.0556875
R37060 C10_P_btm.n250 C10_P_btm.n231 0.0556875
R37061 C10_P_btm.n3499 C10_P_btm.n3498 0.0556875
R37062 C10_P_btm.n3504 C10_P_btm.n189 0.0556875
R37063 C10_P_btm.n3533 C10_P_btm.n3532 0.0556875
R37064 C10_P_btm.n3535 C10_P_btm.n3534 0.0556875
R37065 C10_P_btm.n3564 C10_P_btm.n3563 0.0556875
R37066 C10_P_btm.n3566 C10_P_btm.n3565 0.0556875
R37067 C10_P_btm.n197 C10_P_btm.n178 0.0556875
R37068 C10_P_btm.n3600 C10_P_btm.n3599 0.0556875
R37069 C10_P_btm.n3571 C10_P_btm.n136 0.0556875
R37070 C10_P_btm.n3631 C10_P_btm.n3630 0.0556875
R37071 C10_P_btm.n3602 C10_P_btm.n3601 0.0556875
R37072 C10_P_btm.n144 C10_P_btm.n125 0.0556875
R37073 C10_P_btm.n3633 C10_P_btm.n3632 0.0556875
R37074 C10_P_btm.n3638 C10_P_btm.n83 0.0556875
R37075 C10_P_btm.n3667 C10_P_btm.n3666 0.0556875
R37076 C10_P_btm.n3669 C10_P_btm.n3668 0.0556875
R37077 C10_P_btm.n3698 C10_P_btm.n3697 0.0556875
R37078 C10_P_btm.n3700 C10_P_btm.n3699 0.0556875
R37079 C10_P_btm.n91 C10_P_btm.n72 0.0556875
R37080 C10_P_btm.n3734 C10_P_btm.n3733 0.0556875
R37081 C10_P_btm.n3705 C10_P_btm.n63 0.0556875
R37082 C10_P_btm.n3800 C10_P_btm.n3799 0.0556875
R37083 C10_P_btm.n3771 C10_P_btm.n3770 0.0556875
R37084 C10_P_btm.n3769 C10_P_btm.n3768 0.0556875
R37085 C10_P_btm.n3802 C10_P_btm.n3801 0.0556875
R37086 C10_P_btm.n3807 C10_P_btm.n43 0.0556875
R37087 C10_P_btm.n3736 C10_P_btm.n3735 0.0556875
R37088 C10_P_btm.n3836 C10_P_btm.n33 0.0556875
R37089 C10_P_btm.n3865 C10_P_btm.n3864 0.0556875
R37090 C10_P_btm.n3867 C10_P_btm.n3866 0.0556875
R37091 C10_P_btm.n3896 C10_P_btm.n3895 0.0556875
R37092 a_n1522_42718.n1 a_n1522_42718.t4 685.552
R37093 a_n1522_42718.n1 a_n1522_42718.n0 296.139
R37094 a_n1522_42718.n2 a_n1522_42718.n1 269.182
R37095 a_n1522_42718.n0 a_n1522_42718.t2 26.5955
R37096 a_n1522_42718.n0 a_n1522_42718.t3 26.5955
R37097 a_n1522_42718.n2 a_n1522_42718.t0 24.9236
R37098 a_n1522_42718.t1 a_n1522_42718.n2 24.9236
R37099 C10_N_btm C10_N_btm.n32 92.1672
R37100 C10_N_btm.n2 C10_N_btm.n0 33.0802
R37101 C10_N_btm.n14 C10_N_btm.n13 32.3614
R37102 C10_N_btm.n12 C10_N_btm.n11 32.3614
R37103 C10_N_btm.n10 C10_N_btm.n9 32.3614
R37104 C10_N_btm.n8 C10_N_btm.n7 32.3614
R37105 C10_N_btm.n6 C10_N_btm.n5 32.3614
R37106 C10_N_btm.n4 C10_N_btm.n3 32.3614
R37107 C10_N_btm.n2 C10_N_btm.n1 32.3614
R37108 C10_N_btm.n22 C10_N_btm.n14 29.1203
R37109 C10_N_btm.n24 C10_N_btm.n23 20.3263
R37110 C10_N_btm.n27 C10_N_btm.n25 15.4755
R37111 C10_N_btm.n17 C10_N_btm.n15 15.394
R37112 C10_N_btm.n31 C10_N_btm.n30 14.9755
R37113 C10_N_btm.n29 C10_N_btm.n28 14.9755
R37114 C10_N_btm.n27 C10_N_btm.n26 14.9755
R37115 C10_N_btm.n21 C10_N_btm.n20 14.894
R37116 C10_N_btm.n19 C10_N_btm.n18 14.894
R37117 C10_N_btm.n17 C10_N_btm.n16 14.894
R37118 C10_N_btm.n24 C10_N_btm.n22 6.29217
R37119 C10_N_btm C10_N_btm.n3897 6.2755
R37120 C10_N_btm.n22 C10_N_btm.n21 5.43279
R37121 C10_N_btm.n32 C10_N_btm.n31 5.33904
R37122 C10_N_btm.n34 C10_N_btm.t1061 5.03712
R37123 C10_N_btm.n35 C10_N_btm.t1074 5.03712
R37124 C10_N_btm.n36 C10_N_btm.t1069 5.03712
R37125 C10_N_btm.n37 C10_N_btm.t1067 5.03712
R37126 C10_N_btm.n38 C10_N_btm.t1079 5.03712
R37127 C10_N_btm.n39 C10_N_btm.t1065 5.03712
R37128 C10_N_btm.n40 C10_N_btm.t1071 5.03712
R37129 C10_N_btm.n41 C10_N_btm.t1062 5.03712
R37130 C10_N_btm.n42 C10_N_btm.t1070 5.03712
R37131 C10_N_btm.n904 C10_N_btm.t1078 5.03712
R37132 C10_N_btm.n920 C10_N_btm.t1072 5.03712
R37133 C10_N_btm.n919 C10_N_btm.t1076 5.03712
R37134 C10_N_btm.n918 C10_N_btm.t1063 5.03712
R37135 C10_N_btm.n917 C10_N_btm.t1073 5.03712
R37136 C10_N_btm.n916 C10_N_btm.t1060 5.03712
R37137 C10_N_btm.n915 C10_N_btm.t1068 5.03712
R37138 C10_N_btm.n914 C10_N_btm.t1058 5.03712
R37139 C10_N_btm.n913 C10_N_btm.t1066 5.03712
R37140 C10_N_btm.n951 C10_N_btm.t1077 5.03712
R37141 C10_N_btm.n947 C10_N_btm.t1064 5.03712
R37142 C10_N_btm.n3866 C10_N_btm.t1059 5.03712
R37143 C10_N_btm.n32 C10_N_btm.n24 4.7505
R37144 C10_N_btm.n3893 C10_N_btm.n3892 4.60698
R37145 C10_N_btm.n3894 C10_N_btm.n3893 4.60698
R37146 C10_N_btm.n3890 C10_N_btm.n3889 4.60698
R37147 C10_N_btm.n3891 C10_N_btm.n3890 4.60698
R37148 C10_N_btm.n3887 C10_N_btm.n3886 4.60698
R37149 C10_N_btm.n3888 C10_N_btm.n3887 4.60698
R37150 C10_N_btm.n3884 C10_N_btm.n3883 4.60698
R37151 C10_N_btm.n3885 C10_N_btm.n3884 4.60698
R37152 C10_N_btm.n3881 C10_N_btm.n3880 4.60698
R37153 C10_N_btm.n3882 C10_N_btm.n3881 4.60698
R37154 C10_N_btm.n3878 C10_N_btm.n3877 4.60698
R37155 C10_N_btm.n3879 C10_N_btm.n3878 4.60698
R37156 C10_N_btm.n3875 C10_N_btm.n3874 4.60698
R37157 C10_N_btm.n3876 C10_N_btm.n3875 4.60698
R37158 C10_N_btm.n3872 C10_N_btm.n3871 4.60698
R37159 C10_N_btm.n3873 C10_N_btm.n3872 4.60698
R37160 C10_N_btm.n3869 C10_N_btm.n3868 4.60698
R37161 C10_N_btm.n3870 C10_N_btm.n3869 4.60698
R37162 C10_N_btm.n3863 C10_N_btm.n3862 4.60698
R37163 C10_N_btm.n3862 C10_N_btm.n3861 4.60698
R37164 C10_N_btm.n3860 C10_N_btm.n3859 4.60698
R37165 C10_N_btm.n3859 C10_N_btm.n3858 4.60698
R37166 C10_N_btm.n3857 C10_N_btm.n3856 4.60698
R37167 C10_N_btm.n3856 C10_N_btm.n3855 4.60698
R37168 C10_N_btm.n3854 C10_N_btm.n3853 4.60698
R37169 C10_N_btm.n3853 C10_N_btm.n3852 4.60698
R37170 C10_N_btm.n3851 C10_N_btm.n3850 4.60698
R37171 C10_N_btm.n3850 C10_N_btm.n3849 4.60698
R37172 C10_N_btm.n3848 C10_N_btm.n3847 4.60698
R37173 C10_N_btm.n3847 C10_N_btm.n3846 4.60698
R37174 C10_N_btm.n3845 C10_N_btm.n3844 4.60698
R37175 C10_N_btm.n3844 C10_N_btm.n3843 4.60698
R37176 C10_N_btm.n3842 C10_N_btm.n3841 4.60698
R37177 C10_N_btm.n3841 C10_N_btm.n3840 4.60698
R37178 C10_N_btm.n3839 C10_N_btm.n3838 4.60698
R37179 C10_N_btm.n3838 C10_N_btm.n3837 4.60698
R37180 C10_N_btm.n3833 C10_N_btm.n3832 4.60698
R37181 C10_N_btm.n3832 C10_N_btm.n53 4.60698
R37182 C10_N_btm.n3830 C10_N_btm.n3829 4.60698
R37183 C10_N_btm.n3831 C10_N_btm.n3830 4.60698
R37184 C10_N_btm.n3827 C10_N_btm.n3826 4.60698
R37185 C10_N_btm.n3828 C10_N_btm.n3827 4.60698
R37186 C10_N_btm.n3824 C10_N_btm.n3823 4.60698
R37187 C10_N_btm.n3825 C10_N_btm.n3824 4.60698
R37188 C10_N_btm.n3821 C10_N_btm.n3820 4.60698
R37189 C10_N_btm.n3822 C10_N_btm.n3821 4.60698
R37190 C10_N_btm.n3818 C10_N_btm.n3817 4.60698
R37191 C10_N_btm.n3819 C10_N_btm.n3818 4.60698
R37192 C10_N_btm.n3815 C10_N_btm.n3814 4.60698
R37193 C10_N_btm.n3816 C10_N_btm.n3815 4.60698
R37194 C10_N_btm.n3812 C10_N_btm.n3811 4.60698
R37195 C10_N_btm.n3813 C10_N_btm.n3812 4.60698
R37196 C10_N_btm.n3809 C10_N_btm.n3808 4.60698
R37197 C10_N_btm.n3810 C10_N_btm.n3809 4.60698
R37198 C10_N_btm.n3804 C10_N_btm.n3803 4.60698
R37199 C10_N_btm.n3803 C10_N_btm.n62 4.60698
R37200 C10_N_btm.n3745 C10_N_btm.n3744 4.60698
R37201 C10_N_btm.n3746 C10_N_btm.n3745 4.60698
R37202 C10_N_btm.n3748 C10_N_btm.n3747 4.60698
R37203 C10_N_btm.n3749 C10_N_btm.n3748 4.60698
R37204 C10_N_btm.n3751 C10_N_btm.n3750 4.60698
R37205 C10_N_btm.n3752 C10_N_btm.n3751 4.60698
R37206 C10_N_btm.n3754 C10_N_btm.n3753 4.60698
R37207 C10_N_btm.n3755 C10_N_btm.n3754 4.60698
R37208 C10_N_btm.n3757 C10_N_btm.n3756 4.60698
R37209 C10_N_btm.n3758 C10_N_btm.n3757 4.60698
R37210 C10_N_btm.n3760 C10_N_btm.n3759 4.60698
R37211 C10_N_btm.n3761 C10_N_btm.n3760 4.60698
R37212 C10_N_btm.n3763 C10_N_btm.n3762 4.60698
R37213 C10_N_btm.n3764 C10_N_btm.n3763 4.60698
R37214 C10_N_btm.n3766 C10_N_btm.n3765 4.60698
R37215 C10_N_btm.n3767 C10_N_btm.n3766 4.60698
R37216 C10_N_btm.n3774 C10_N_btm.n3773 4.60698
R37217 C10_N_btm.n3773 C10_N_btm.n3772 4.60698
R37218 C10_N_btm.n3777 C10_N_btm.n3776 4.60698
R37219 C10_N_btm.n3776 C10_N_btm.n3775 4.60698
R37220 C10_N_btm.n3780 C10_N_btm.n3779 4.60698
R37221 C10_N_btm.n3779 C10_N_btm.n3778 4.60698
R37222 C10_N_btm.n3783 C10_N_btm.n3782 4.60698
R37223 C10_N_btm.n3782 C10_N_btm.n3781 4.60698
R37224 C10_N_btm.n3786 C10_N_btm.n3785 4.60698
R37225 C10_N_btm.n3785 C10_N_btm.n3784 4.60698
R37226 C10_N_btm.n3789 C10_N_btm.n3788 4.60698
R37227 C10_N_btm.n3788 C10_N_btm.n3787 4.60698
R37228 C10_N_btm.n3792 C10_N_btm.n3791 4.60698
R37229 C10_N_btm.n3791 C10_N_btm.n3790 4.60698
R37230 C10_N_btm.n3795 C10_N_btm.n3794 4.60698
R37231 C10_N_btm.n3794 C10_N_btm.n3793 4.60698
R37232 C10_N_btm.n3798 C10_N_btm.n3797 4.60698
R37233 C10_N_btm.n3797 C10_N_btm.n3796 4.60698
R37234 C10_N_btm.n3707 C10_N_btm.n3706 4.60698
R37235 C10_N_btm.n3708 C10_N_btm.n3707 4.60698
R37236 C10_N_btm.n3710 C10_N_btm.n3709 4.60698
R37237 C10_N_btm.n3711 C10_N_btm.n3710 4.60698
R37238 C10_N_btm.n3713 C10_N_btm.n3712 4.60698
R37239 C10_N_btm.n3714 C10_N_btm.n3713 4.60698
R37240 C10_N_btm.n3716 C10_N_btm.n3715 4.60698
R37241 C10_N_btm.n3717 C10_N_btm.n3716 4.60698
R37242 C10_N_btm.n3719 C10_N_btm.n3718 4.60698
R37243 C10_N_btm.n3720 C10_N_btm.n3719 4.60698
R37244 C10_N_btm.n3722 C10_N_btm.n3721 4.60698
R37245 C10_N_btm.n3723 C10_N_btm.n3722 4.60698
R37246 C10_N_btm.n3725 C10_N_btm.n3724 4.60698
R37247 C10_N_btm.n3726 C10_N_btm.n3725 4.60698
R37248 C10_N_btm.n3728 C10_N_btm.n3727 4.60698
R37249 C10_N_btm.n3729 C10_N_btm.n3728 4.60698
R37250 C10_N_btm.n3731 C10_N_btm.n3730 4.60698
R37251 C10_N_btm.n3732 C10_N_btm.n3731 4.60698
R37252 C10_N_btm.n122 C10_N_btm.n121 4.60698
R37253 C10_N_btm.n121 C10_N_btm.n92 4.60698
R37254 C10_N_btm.n119 C10_N_btm.n118 4.60698
R37255 C10_N_btm.n120 C10_N_btm.n119 4.60698
R37256 C10_N_btm.n116 C10_N_btm.n115 4.60698
R37257 C10_N_btm.n117 C10_N_btm.n116 4.60698
R37258 C10_N_btm.n113 C10_N_btm.n112 4.60698
R37259 C10_N_btm.n114 C10_N_btm.n113 4.60698
R37260 C10_N_btm.n110 C10_N_btm.n109 4.60698
R37261 C10_N_btm.n111 C10_N_btm.n110 4.60698
R37262 C10_N_btm.n107 C10_N_btm.n106 4.60698
R37263 C10_N_btm.n108 C10_N_btm.n107 4.60698
R37264 C10_N_btm.n104 C10_N_btm.n103 4.60698
R37265 C10_N_btm.n105 C10_N_btm.n104 4.60698
R37266 C10_N_btm.n101 C10_N_btm.n100 4.60698
R37267 C10_N_btm.n102 C10_N_btm.n101 4.60698
R37268 C10_N_btm.n3702 C10_N_btm.n3701 4.60698
R37269 C10_N_btm.n3701 C10_N_btm.n82 4.60698
R37270 C10_N_btm.n3696 C10_N_btm.n3695 4.60698
R37271 C10_N_btm.n3695 C10_N_btm.n3694 4.60698
R37272 C10_N_btm.n3693 C10_N_btm.n3692 4.60698
R37273 C10_N_btm.n3692 C10_N_btm.n3691 4.60698
R37274 C10_N_btm.n3690 C10_N_btm.n3689 4.60698
R37275 C10_N_btm.n3689 C10_N_btm.n3688 4.60698
R37276 C10_N_btm.n3687 C10_N_btm.n3686 4.60698
R37277 C10_N_btm.n3686 C10_N_btm.n3685 4.60698
R37278 C10_N_btm.n3684 C10_N_btm.n3683 4.60698
R37279 C10_N_btm.n3683 C10_N_btm.n3682 4.60698
R37280 C10_N_btm.n3681 C10_N_btm.n3680 4.60698
R37281 C10_N_btm.n3680 C10_N_btm.n3679 4.60698
R37282 C10_N_btm.n3678 C10_N_btm.n3677 4.60698
R37283 C10_N_btm.n3677 C10_N_btm.n3676 4.60698
R37284 C10_N_btm.n3675 C10_N_btm.n3674 4.60698
R37285 C10_N_btm.n3674 C10_N_btm.n3673 4.60698
R37286 C10_N_btm.n3672 C10_N_btm.n3671 4.60698
R37287 C10_N_btm.n3671 C10_N_btm.n3670 4.60698
R37288 C10_N_btm.n3664 C10_N_btm.n3663 4.60698
R37289 C10_N_btm.n3665 C10_N_btm.n3664 4.60698
R37290 C10_N_btm.n3661 C10_N_btm.n3660 4.60698
R37291 C10_N_btm.n3662 C10_N_btm.n3661 4.60698
R37292 C10_N_btm.n3658 C10_N_btm.n3657 4.60698
R37293 C10_N_btm.n3659 C10_N_btm.n3658 4.60698
R37294 C10_N_btm.n3655 C10_N_btm.n3654 4.60698
R37295 C10_N_btm.n3656 C10_N_btm.n3655 4.60698
R37296 C10_N_btm.n3652 C10_N_btm.n3651 4.60698
R37297 C10_N_btm.n3653 C10_N_btm.n3652 4.60698
R37298 C10_N_btm.n3649 C10_N_btm.n3648 4.60698
R37299 C10_N_btm.n3650 C10_N_btm.n3649 4.60698
R37300 C10_N_btm.n3646 C10_N_btm.n3645 4.60698
R37301 C10_N_btm.n3647 C10_N_btm.n3646 4.60698
R37302 C10_N_btm.n3643 C10_N_btm.n3642 4.60698
R37303 C10_N_btm.n3644 C10_N_btm.n3643 4.60698
R37304 C10_N_btm.n3640 C10_N_btm.n3639 4.60698
R37305 C10_N_btm.n3641 C10_N_btm.n3640 4.60698
R37306 C10_N_btm.n3635 C10_N_btm.n3634 4.60698
R37307 C10_N_btm.n3634 C10_N_btm.n135 4.60698
R37308 C10_N_btm.n154 C10_N_btm.n153 4.60698
R37309 C10_N_btm.n155 C10_N_btm.n154 4.60698
R37310 C10_N_btm.n157 C10_N_btm.n156 4.60698
R37311 C10_N_btm.n158 C10_N_btm.n157 4.60698
R37312 C10_N_btm.n160 C10_N_btm.n159 4.60698
R37313 C10_N_btm.n161 C10_N_btm.n160 4.60698
R37314 C10_N_btm.n163 C10_N_btm.n162 4.60698
R37315 C10_N_btm.n164 C10_N_btm.n163 4.60698
R37316 C10_N_btm.n166 C10_N_btm.n165 4.60698
R37317 C10_N_btm.n167 C10_N_btm.n166 4.60698
R37318 C10_N_btm.n169 C10_N_btm.n168 4.60698
R37319 C10_N_btm.n170 C10_N_btm.n169 4.60698
R37320 C10_N_btm.n172 C10_N_btm.n171 4.60698
R37321 C10_N_btm.n173 C10_N_btm.n172 4.60698
R37322 C10_N_btm.n175 C10_N_btm.n174 4.60698
R37323 C10_N_btm.n174 C10_N_btm.n145 4.60698
R37324 C10_N_btm.n3605 C10_N_btm.n3604 4.60698
R37325 C10_N_btm.n3604 C10_N_btm.n3603 4.60698
R37326 C10_N_btm.n3608 C10_N_btm.n3607 4.60698
R37327 C10_N_btm.n3607 C10_N_btm.n3606 4.60698
R37328 C10_N_btm.n3611 C10_N_btm.n3610 4.60698
R37329 C10_N_btm.n3610 C10_N_btm.n3609 4.60698
R37330 C10_N_btm.n3614 C10_N_btm.n3613 4.60698
R37331 C10_N_btm.n3613 C10_N_btm.n3612 4.60698
R37332 C10_N_btm.n3617 C10_N_btm.n3616 4.60698
R37333 C10_N_btm.n3616 C10_N_btm.n3615 4.60698
R37334 C10_N_btm.n3620 C10_N_btm.n3619 4.60698
R37335 C10_N_btm.n3619 C10_N_btm.n3618 4.60698
R37336 C10_N_btm.n3623 C10_N_btm.n3622 4.60698
R37337 C10_N_btm.n3622 C10_N_btm.n3621 4.60698
R37338 C10_N_btm.n3626 C10_N_btm.n3625 4.60698
R37339 C10_N_btm.n3625 C10_N_btm.n3624 4.60698
R37340 C10_N_btm.n3629 C10_N_btm.n3628 4.60698
R37341 C10_N_btm.n3628 C10_N_btm.n3627 4.60698
R37342 C10_N_btm.n3573 C10_N_btm.n3572 4.60698
R37343 C10_N_btm.n3574 C10_N_btm.n3573 4.60698
R37344 C10_N_btm.n3576 C10_N_btm.n3575 4.60698
R37345 C10_N_btm.n3577 C10_N_btm.n3576 4.60698
R37346 C10_N_btm.n3579 C10_N_btm.n3578 4.60698
R37347 C10_N_btm.n3580 C10_N_btm.n3579 4.60698
R37348 C10_N_btm.n3582 C10_N_btm.n3581 4.60698
R37349 C10_N_btm.n3583 C10_N_btm.n3582 4.60698
R37350 C10_N_btm.n3585 C10_N_btm.n3584 4.60698
R37351 C10_N_btm.n3586 C10_N_btm.n3585 4.60698
R37352 C10_N_btm.n3588 C10_N_btm.n3587 4.60698
R37353 C10_N_btm.n3589 C10_N_btm.n3588 4.60698
R37354 C10_N_btm.n3591 C10_N_btm.n3590 4.60698
R37355 C10_N_btm.n3592 C10_N_btm.n3591 4.60698
R37356 C10_N_btm.n3594 C10_N_btm.n3593 4.60698
R37357 C10_N_btm.n3595 C10_N_btm.n3594 4.60698
R37358 C10_N_btm.n3597 C10_N_btm.n3596 4.60698
R37359 C10_N_btm.n3598 C10_N_btm.n3597 4.60698
R37360 C10_N_btm.n228 C10_N_btm.n227 4.60698
R37361 C10_N_btm.n227 C10_N_btm.n198 4.60698
R37362 C10_N_btm.n225 C10_N_btm.n224 4.60698
R37363 C10_N_btm.n226 C10_N_btm.n225 4.60698
R37364 C10_N_btm.n222 C10_N_btm.n221 4.60698
R37365 C10_N_btm.n223 C10_N_btm.n222 4.60698
R37366 C10_N_btm.n219 C10_N_btm.n218 4.60698
R37367 C10_N_btm.n220 C10_N_btm.n219 4.60698
R37368 C10_N_btm.n216 C10_N_btm.n215 4.60698
R37369 C10_N_btm.n217 C10_N_btm.n216 4.60698
R37370 C10_N_btm.n213 C10_N_btm.n212 4.60698
R37371 C10_N_btm.n214 C10_N_btm.n213 4.60698
R37372 C10_N_btm.n210 C10_N_btm.n209 4.60698
R37373 C10_N_btm.n211 C10_N_btm.n210 4.60698
R37374 C10_N_btm.n207 C10_N_btm.n206 4.60698
R37375 C10_N_btm.n208 C10_N_btm.n207 4.60698
R37376 C10_N_btm.n3568 C10_N_btm.n3567 4.60698
R37377 C10_N_btm.n3567 C10_N_btm.n188 4.60698
R37378 C10_N_btm.n3562 C10_N_btm.n3561 4.60698
R37379 C10_N_btm.n3561 C10_N_btm.n3560 4.60698
R37380 C10_N_btm.n3559 C10_N_btm.n3558 4.60698
R37381 C10_N_btm.n3558 C10_N_btm.n3557 4.60698
R37382 C10_N_btm.n3556 C10_N_btm.n3555 4.60698
R37383 C10_N_btm.n3555 C10_N_btm.n3554 4.60698
R37384 C10_N_btm.n3553 C10_N_btm.n3552 4.60698
R37385 C10_N_btm.n3552 C10_N_btm.n3551 4.60698
R37386 C10_N_btm.n3550 C10_N_btm.n3549 4.60698
R37387 C10_N_btm.n3549 C10_N_btm.n3548 4.60698
R37388 C10_N_btm.n3547 C10_N_btm.n3546 4.60698
R37389 C10_N_btm.n3546 C10_N_btm.n3545 4.60698
R37390 C10_N_btm.n3544 C10_N_btm.n3543 4.60698
R37391 C10_N_btm.n3543 C10_N_btm.n3542 4.60698
R37392 C10_N_btm.n3541 C10_N_btm.n3540 4.60698
R37393 C10_N_btm.n3540 C10_N_btm.n3539 4.60698
R37394 C10_N_btm.n3538 C10_N_btm.n3537 4.60698
R37395 C10_N_btm.n3537 C10_N_btm.n3536 4.60698
R37396 C10_N_btm.n3530 C10_N_btm.n3529 4.60698
R37397 C10_N_btm.n3531 C10_N_btm.n3530 4.60698
R37398 C10_N_btm.n3527 C10_N_btm.n3526 4.60698
R37399 C10_N_btm.n3528 C10_N_btm.n3527 4.60698
R37400 C10_N_btm.n3524 C10_N_btm.n3523 4.60698
R37401 C10_N_btm.n3525 C10_N_btm.n3524 4.60698
R37402 C10_N_btm.n3521 C10_N_btm.n3520 4.60698
R37403 C10_N_btm.n3522 C10_N_btm.n3521 4.60698
R37404 C10_N_btm.n3518 C10_N_btm.n3517 4.60698
R37405 C10_N_btm.n3519 C10_N_btm.n3518 4.60698
R37406 C10_N_btm.n3515 C10_N_btm.n3514 4.60698
R37407 C10_N_btm.n3516 C10_N_btm.n3515 4.60698
R37408 C10_N_btm.n3512 C10_N_btm.n3511 4.60698
R37409 C10_N_btm.n3513 C10_N_btm.n3512 4.60698
R37410 C10_N_btm.n3509 C10_N_btm.n3508 4.60698
R37411 C10_N_btm.n3510 C10_N_btm.n3509 4.60698
R37412 C10_N_btm.n3506 C10_N_btm.n3505 4.60698
R37413 C10_N_btm.n3507 C10_N_btm.n3506 4.60698
R37414 C10_N_btm.n3501 C10_N_btm.n3500 4.60698
R37415 C10_N_btm.n3500 C10_N_btm.n241 4.60698
R37416 C10_N_btm.n260 C10_N_btm.n259 4.60698
R37417 C10_N_btm.n261 C10_N_btm.n260 4.60698
R37418 C10_N_btm.n263 C10_N_btm.n262 4.60698
R37419 C10_N_btm.n264 C10_N_btm.n263 4.60698
R37420 C10_N_btm.n266 C10_N_btm.n265 4.60698
R37421 C10_N_btm.n267 C10_N_btm.n266 4.60698
R37422 C10_N_btm.n269 C10_N_btm.n268 4.60698
R37423 C10_N_btm.n270 C10_N_btm.n269 4.60698
R37424 C10_N_btm.n272 C10_N_btm.n271 4.60698
R37425 C10_N_btm.n273 C10_N_btm.n272 4.60698
R37426 C10_N_btm.n275 C10_N_btm.n274 4.60698
R37427 C10_N_btm.n276 C10_N_btm.n275 4.60698
R37428 C10_N_btm.n278 C10_N_btm.n277 4.60698
R37429 C10_N_btm.n279 C10_N_btm.n278 4.60698
R37430 C10_N_btm.n281 C10_N_btm.n280 4.60698
R37431 C10_N_btm.n280 C10_N_btm.n251 4.60698
R37432 C10_N_btm.n3471 C10_N_btm.n3470 4.60698
R37433 C10_N_btm.n3470 C10_N_btm.n3469 4.60698
R37434 C10_N_btm.n3474 C10_N_btm.n3473 4.60698
R37435 C10_N_btm.n3473 C10_N_btm.n3472 4.60698
R37436 C10_N_btm.n3477 C10_N_btm.n3476 4.60698
R37437 C10_N_btm.n3476 C10_N_btm.n3475 4.60698
R37438 C10_N_btm.n3480 C10_N_btm.n3479 4.60698
R37439 C10_N_btm.n3479 C10_N_btm.n3478 4.60698
R37440 C10_N_btm.n3483 C10_N_btm.n3482 4.60698
R37441 C10_N_btm.n3482 C10_N_btm.n3481 4.60698
R37442 C10_N_btm.n3486 C10_N_btm.n3485 4.60698
R37443 C10_N_btm.n3485 C10_N_btm.n3484 4.60698
R37444 C10_N_btm.n3489 C10_N_btm.n3488 4.60698
R37445 C10_N_btm.n3488 C10_N_btm.n3487 4.60698
R37446 C10_N_btm.n3492 C10_N_btm.n3491 4.60698
R37447 C10_N_btm.n3491 C10_N_btm.n3490 4.60698
R37448 C10_N_btm.n3495 C10_N_btm.n3494 4.60698
R37449 C10_N_btm.n3494 C10_N_btm.n3493 4.60698
R37450 C10_N_btm.n3439 C10_N_btm.n3438 4.60698
R37451 C10_N_btm.n3440 C10_N_btm.n3439 4.60698
R37452 C10_N_btm.n3442 C10_N_btm.n3441 4.60698
R37453 C10_N_btm.n3443 C10_N_btm.n3442 4.60698
R37454 C10_N_btm.n3445 C10_N_btm.n3444 4.60698
R37455 C10_N_btm.n3446 C10_N_btm.n3445 4.60698
R37456 C10_N_btm.n3448 C10_N_btm.n3447 4.60698
R37457 C10_N_btm.n3449 C10_N_btm.n3448 4.60698
R37458 C10_N_btm.n3451 C10_N_btm.n3450 4.60698
R37459 C10_N_btm.n3452 C10_N_btm.n3451 4.60698
R37460 C10_N_btm.n3454 C10_N_btm.n3453 4.60698
R37461 C10_N_btm.n3455 C10_N_btm.n3454 4.60698
R37462 C10_N_btm.n3457 C10_N_btm.n3456 4.60698
R37463 C10_N_btm.n3458 C10_N_btm.n3457 4.60698
R37464 C10_N_btm.n3460 C10_N_btm.n3459 4.60698
R37465 C10_N_btm.n3461 C10_N_btm.n3460 4.60698
R37466 C10_N_btm.n3463 C10_N_btm.n3462 4.60698
R37467 C10_N_btm.n3464 C10_N_btm.n3463 4.60698
R37468 C10_N_btm.n334 C10_N_btm.n333 4.60698
R37469 C10_N_btm.n333 C10_N_btm.n304 4.60698
R37470 C10_N_btm.n331 C10_N_btm.n330 4.60698
R37471 C10_N_btm.n332 C10_N_btm.n331 4.60698
R37472 C10_N_btm.n328 C10_N_btm.n327 4.60698
R37473 C10_N_btm.n329 C10_N_btm.n328 4.60698
R37474 C10_N_btm.n325 C10_N_btm.n324 4.60698
R37475 C10_N_btm.n326 C10_N_btm.n325 4.60698
R37476 C10_N_btm.n322 C10_N_btm.n321 4.60698
R37477 C10_N_btm.n323 C10_N_btm.n322 4.60698
R37478 C10_N_btm.n319 C10_N_btm.n318 4.60698
R37479 C10_N_btm.n320 C10_N_btm.n319 4.60698
R37480 C10_N_btm.n316 C10_N_btm.n315 4.60698
R37481 C10_N_btm.n317 C10_N_btm.n316 4.60698
R37482 C10_N_btm.n313 C10_N_btm.n312 4.60698
R37483 C10_N_btm.n314 C10_N_btm.n313 4.60698
R37484 C10_N_btm.n3434 C10_N_btm.n3433 4.60698
R37485 C10_N_btm.n3433 C10_N_btm.n294 4.60698
R37486 C10_N_btm.n3428 C10_N_btm.n3427 4.60698
R37487 C10_N_btm.n3427 C10_N_btm.n3426 4.60698
R37488 C10_N_btm.n3425 C10_N_btm.n3424 4.60698
R37489 C10_N_btm.n3424 C10_N_btm.n3423 4.60698
R37490 C10_N_btm.n3422 C10_N_btm.n3421 4.60698
R37491 C10_N_btm.n3421 C10_N_btm.n3420 4.60698
R37492 C10_N_btm.n3419 C10_N_btm.n3418 4.60698
R37493 C10_N_btm.n3418 C10_N_btm.n3417 4.60698
R37494 C10_N_btm.n3416 C10_N_btm.n3415 4.60698
R37495 C10_N_btm.n3415 C10_N_btm.n3414 4.60698
R37496 C10_N_btm.n3413 C10_N_btm.n3412 4.60698
R37497 C10_N_btm.n3412 C10_N_btm.n3411 4.60698
R37498 C10_N_btm.n3410 C10_N_btm.n3409 4.60698
R37499 C10_N_btm.n3409 C10_N_btm.n3408 4.60698
R37500 C10_N_btm.n3407 C10_N_btm.n3406 4.60698
R37501 C10_N_btm.n3406 C10_N_btm.n3405 4.60698
R37502 C10_N_btm.n3404 C10_N_btm.n3403 4.60698
R37503 C10_N_btm.n3403 C10_N_btm.n3402 4.60698
R37504 C10_N_btm.n3396 C10_N_btm.n3395 4.60698
R37505 C10_N_btm.n3397 C10_N_btm.n3396 4.60698
R37506 C10_N_btm.n3393 C10_N_btm.n3392 4.60698
R37507 C10_N_btm.n3394 C10_N_btm.n3393 4.60698
R37508 C10_N_btm.n3390 C10_N_btm.n3389 4.60698
R37509 C10_N_btm.n3391 C10_N_btm.n3390 4.60698
R37510 C10_N_btm.n3387 C10_N_btm.n3386 4.60698
R37511 C10_N_btm.n3388 C10_N_btm.n3387 4.60698
R37512 C10_N_btm.n3384 C10_N_btm.n3383 4.60698
R37513 C10_N_btm.n3385 C10_N_btm.n3384 4.60698
R37514 C10_N_btm.n3381 C10_N_btm.n3380 4.60698
R37515 C10_N_btm.n3382 C10_N_btm.n3381 4.60698
R37516 C10_N_btm.n3378 C10_N_btm.n3377 4.60698
R37517 C10_N_btm.n3379 C10_N_btm.n3378 4.60698
R37518 C10_N_btm.n3375 C10_N_btm.n3374 4.60698
R37519 C10_N_btm.n3376 C10_N_btm.n3375 4.60698
R37520 C10_N_btm.n3372 C10_N_btm.n3371 4.60698
R37521 C10_N_btm.n3373 C10_N_btm.n3372 4.60698
R37522 C10_N_btm.n3367 C10_N_btm.n3366 4.60698
R37523 C10_N_btm.n3366 C10_N_btm.n347 4.60698
R37524 C10_N_btm.n366 C10_N_btm.n365 4.60698
R37525 C10_N_btm.n367 C10_N_btm.n366 4.60698
R37526 C10_N_btm.n369 C10_N_btm.n368 4.60698
R37527 C10_N_btm.n370 C10_N_btm.n369 4.60698
R37528 C10_N_btm.n372 C10_N_btm.n371 4.60698
R37529 C10_N_btm.n373 C10_N_btm.n372 4.60698
R37530 C10_N_btm.n375 C10_N_btm.n374 4.60698
R37531 C10_N_btm.n376 C10_N_btm.n375 4.60698
R37532 C10_N_btm.n378 C10_N_btm.n377 4.60698
R37533 C10_N_btm.n379 C10_N_btm.n378 4.60698
R37534 C10_N_btm.n381 C10_N_btm.n380 4.60698
R37535 C10_N_btm.n382 C10_N_btm.n381 4.60698
R37536 C10_N_btm.n384 C10_N_btm.n383 4.60698
R37537 C10_N_btm.n385 C10_N_btm.n384 4.60698
R37538 C10_N_btm.n387 C10_N_btm.n386 4.60698
R37539 C10_N_btm.n386 C10_N_btm.n357 4.60698
R37540 C10_N_btm.n3337 C10_N_btm.n3336 4.60698
R37541 C10_N_btm.n3336 C10_N_btm.n3335 4.60698
R37542 C10_N_btm.n3340 C10_N_btm.n3339 4.60698
R37543 C10_N_btm.n3339 C10_N_btm.n3338 4.60698
R37544 C10_N_btm.n3343 C10_N_btm.n3342 4.60698
R37545 C10_N_btm.n3342 C10_N_btm.n3341 4.60698
R37546 C10_N_btm.n3346 C10_N_btm.n3345 4.60698
R37547 C10_N_btm.n3345 C10_N_btm.n3344 4.60698
R37548 C10_N_btm.n3349 C10_N_btm.n3348 4.60698
R37549 C10_N_btm.n3348 C10_N_btm.n3347 4.60698
R37550 C10_N_btm.n3352 C10_N_btm.n3351 4.60698
R37551 C10_N_btm.n3351 C10_N_btm.n3350 4.60698
R37552 C10_N_btm.n3355 C10_N_btm.n3354 4.60698
R37553 C10_N_btm.n3354 C10_N_btm.n3353 4.60698
R37554 C10_N_btm.n3358 C10_N_btm.n3357 4.60698
R37555 C10_N_btm.n3357 C10_N_btm.n3356 4.60698
R37556 C10_N_btm.n3361 C10_N_btm.n3360 4.60698
R37557 C10_N_btm.n3360 C10_N_btm.n3359 4.60698
R37558 C10_N_btm.n3305 C10_N_btm.n3304 4.60698
R37559 C10_N_btm.n3306 C10_N_btm.n3305 4.60698
R37560 C10_N_btm.n3308 C10_N_btm.n3307 4.60698
R37561 C10_N_btm.n3309 C10_N_btm.n3308 4.60698
R37562 C10_N_btm.n3311 C10_N_btm.n3310 4.60698
R37563 C10_N_btm.n3312 C10_N_btm.n3311 4.60698
R37564 C10_N_btm.n3314 C10_N_btm.n3313 4.60698
R37565 C10_N_btm.n3315 C10_N_btm.n3314 4.60698
R37566 C10_N_btm.n3317 C10_N_btm.n3316 4.60698
R37567 C10_N_btm.n3318 C10_N_btm.n3317 4.60698
R37568 C10_N_btm.n3320 C10_N_btm.n3319 4.60698
R37569 C10_N_btm.n3321 C10_N_btm.n3320 4.60698
R37570 C10_N_btm.n3323 C10_N_btm.n3322 4.60698
R37571 C10_N_btm.n3324 C10_N_btm.n3323 4.60698
R37572 C10_N_btm.n3326 C10_N_btm.n3325 4.60698
R37573 C10_N_btm.n3327 C10_N_btm.n3326 4.60698
R37574 C10_N_btm.n3329 C10_N_btm.n3328 4.60698
R37575 C10_N_btm.n3330 C10_N_btm.n3329 4.60698
R37576 C10_N_btm.n468 C10_N_btm.n467 4.60698
R37577 C10_N_btm.n469 C10_N_btm.n468 4.60698
R37578 C10_N_btm.n465 C10_N_btm.n464 4.60698
R37579 C10_N_btm.n466 C10_N_btm.n465 4.60698
R37580 C10_N_btm.n462 C10_N_btm.n461 4.60698
R37581 C10_N_btm.n463 C10_N_btm.n462 4.60698
R37582 C10_N_btm.n459 C10_N_btm.n458 4.60698
R37583 C10_N_btm.n460 C10_N_btm.n459 4.60698
R37584 C10_N_btm.n456 C10_N_btm.n455 4.60698
R37585 C10_N_btm.n457 C10_N_btm.n456 4.60698
R37586 C10_N_btm.n453 C10_N_btm.n452 4.60698
R37587 C10_N_btm.n454 C10_N_btm.n453 4.60698
R37588 C10_N_btm.n450 C10_N_btm.n449 4.60698
R37589 C10_N_btm.n451 C10_N_btm.n450 4.60698
R37590 C10_N_btm.n447 C10_N_btm.n446 4.60698
R37591 C10_N_btm.n448 C10_N_btm.n447 4.60698
R37592 C10_N_btm.n444 C10_N_btm.n443 4.60698
R37593 C10_N_btm.n445 C10_N_btm.n444 4.60698
R37594 C10_N_btm.n3300 C10_N_btm.n3299 4.60698
R37595 C10_N_btm.n3299 C10_N_btm.n400 4.60698
R37596 C10_N_btm.n3294 C10_N_btm.n3293 4.60698
R37597 C10_N_btm.n3293 C10_N_btm.n3292 4.60698
R37598 C10_N_btm.n3291 C10_N_btm.n3290 4.60698
R37599 C10_N_btm.n3290 C10_N_btm.n3289 4.60698
R37600 C10_N_btm.n3288 C10_N_btm.n3287 4.60698
R37601 C10_N_btm.n3287 C10_N_btm.n3286 4.60698
R37602 C10_N_btm.n3285 C10_N_btm.n3284 4.60698
R37603 C10_N_btm.n3284 C10_N_btm.n3283 4.60698
R37604 C10_N_btm.n3282 C10_N_btm.n3281 4.60698
R37605 C10_N_btm.n3281 C10_N_btm.n3280 4.60698
R37606 C10_N_btm.n3279 C10_N_btm.n3278 4.60698
R37607 C10_N_btm.n3278 C10_N_btm.n3277 4.60698
R37608 C10_N_btm.n3276 C10_N_btm.n3275 4.60698
R37609 C10_N_btm.n3275 C10_N_btm.n3274 4.60698
R37610 C10_N_btm.n3273 C10_N_btm.n3272 4.60698
R37611 C10_N_btm.n3272 C10_N_btm.n3271 4.60698
R37612 C10_N_btm.n3270 C10_N_btm.n3269 4.60698
R37613 C10_N_btm.n3269 C10_N_btm.n3268 4.60698
R37614 C10_N_btm.n3267 C10_N_btm.n3266 4.60698
R37615 C10_N_btm.n3266 C10_N_btm.n3265 4.60698
R37616 C10_N_btm.n3264 C10_N_btm.n3263 4.60698
R37617 C10_N_btm.n3263 C10_N_btm.n3262 4.60698
R37618 C10_N_btm.n3261 C10_N_btm.n3260 4.60698
R37619 C10_N_btm.n3260 C10_N_btm.n3259 4.60698
R37620 C10_N_btm.n3258 C10_N_btm.n3257 4.60698
R37621 C10_N_btm.n3257 C10_N_btm.n3256 4.60698
R37622 C10_N_btm.n3255 C10_N_btm.n3254 4.60698
R37623 C10_N_btm.n3254 C10_N_btm.n3253 4.60698
R37624 C10_N_btm.n3252 C10_N_btm.n3251 4.60698
R37625 C10_N_btm.n3251 C10_N_btm.n3250 4.60698
R37626 C10_N_btm.n3249 C10_N_btm.n3248 4.60698
R37627 C10_N_btm.n3248 C10_N_btm.n3247 4.60698
R37628 C10_N_btm.n3246 C10_N_btm.n3245 4.60698
R37629 C10_N_btm.n3245 C10_N_btm.n3244 4.60698
R37630 C10_N_btm.n3243 C10_N_btm.n3242 4.60698
R37631 C10_N_btm.n3242 C10_N_btm.n3241 4.60698
R37632 C10_N_btm.n3240 C10_N_btm.n3239 4.60698
R37633 C10_N_btm.n3239 C10_N_btm.n3238 4.60698
R37634 C10_N_btm.n3237 C10_N_btm.n3236 4.60698
R37635 C10_N_btm.n3236 C10_N_btm.n3235 4.60698
R37636 C10_N_btm.n3234 C10_N_btm.n3233 4.60698
R37637 C10_N_btm.n3233 C10_N_btm.n3232 4.60698
R37638 C10_N_btm.n3231 C10_N_btm.n3230 4.60698
R37639 C10_N_btm.n3230 C10_N_btm.n3229 4.60698
R37640 C10_N_btm.n3228 C10_N_btm.n3227 4.60698
R37641 C10_N_btm.n3227 C10_N_btm.n3226 4.60698
R37642 C10_N_btm.n504 C10_N_btm.n503 4.60698
R37643 C10_N_btm.n505 C10_N_btm.n504 4.60698
R37644 C10_N_btm.n501 C10_N_btm.n500 4.60698
R37645 C10_N_btm.n502 C10_N_btm.n501 4.60698
R37646 C10_N_btm.n498 C10_N_btm.n497 4.60698
R37647 C10_N_btm.n499 C10_N_btm.n498 4.60698
R37648 C10_N_btm.n495 C10_N_btm.n494 4.60698
R37649 C10_N_btm.n496 C10_N_btm.n495 4.60698
R37650 C10_N_btm.n492 C10_N_btm.n491 4.60698
R37651 C10_N_btm.n493 C10_N_btm.n492 4.60698
R37652 C10_N_btm.n489 C10_N_btm.n488 4.60698
R37653 C10_N_btm.n490 C10_N_btm.n489 4.60698
R37654 C10_N_btm.n486 C10_N_btm.n485 4.60698
R37655 C10_N_btm.n487 C10_N_btm.n486 4.60698
R37656 C10_N_btm.n483 C10_N_btm.n482 4.60698
R37657 C10_N_btm.n484 C10_N_btm.n483 4.60698
R37658 C10_N_btm.n480 C10_N_btm.n479 4.60698
R37659 C10_N_btm.n481 C10_N_btm.n480 4.60698
R37660 C10_N_btm.n477 C10_N_btm.n476 4.60698
R37661 C10_N_btm.n478 C10_N_btm.n477 4.60698
R37662 C10_N_btm.n474 C10_N_btm.n473 4.60698
R37663 C10_N_btm.n475 C10_N_btm.n474 4.60698
R37664 C10_N_btm.n471 C10_N_btm.n470 4.60698
R37665 C10_N_btm.n472 C10_N_btm.n471 4.60698
R37666 C10_N_btm.n3225 C10_N_btm.n3224 4.60698
R37667 C10_N_btm.n3224 C10_N_btm.n3223 4.60698
R37668 C10_N_btm.n3222 C10_N_btm.n3221 4.60698
R37669 C10_N_btm.n3221 C10_N_btm.n3220 4.60698
R37670 C10_N_btm.n3219 C10_N_btm.n3218 4.60698
R37671 C10_N_btm.n3218 C10_N_btm.n3217 4.60698
R37672 C10_N_btm.n3216 C10_N_btm.n3215 4.60698
R37673 C10_N_btm.n3215 C10_N_btm.n3214 4.60698
R37674 C10_N_btm.n3213 C10_N_btm.n3212 4.60698
R37675 C10_N_btm.n3212 C10_N_btm.n3211 4.60698
R37676 C10_N_btm.n3210 C10_N_btm.n3209 4.60698
R37677 C10_N_btm.n3209 C10_N_btm.n3208 4.60698
R37678 C10_N_btm.n3207 C10_N_btm.n3206 4.60698
R37679 C10_N_btm.n3206 C10_N_btm.n3205 4.60698
R37680 C10_N_btm.n3204 C10_N_btm.n3203 4.60698
R37681 C10_N_btm.n3203 C10_N_btm.n3202 4.60698
R37682 C10_N_btm.n3201 C10_N_btm.n3200 4.60698
R37683 C10_N_btm.n3200 C10_N_btm.n3199 4.60698
R37684 C10_N_btm.n3198 C10_N_btm.n3197 4.60698
R37685 C10_N_btm.n3197 C10_N_btm.n3196 4.60698
R37686 C10_N_btm.n3195 C10_N_btm.n3194 4.60698
R37687 C10_N_btm.n3194 C10_N_btm.n3193 4.60698
R37688 C10_N_btm.n3192 C10_N_btm.n3191 4.60698
R37689 C10_N_btm.n3191 C10_N_btm.n3190 4.60698
R37690 C10_N_btm.n3189 C10_N_btm.n3188 4.60698
R37691 C10_N_btm.n3188 C10_N_btm.n3187 4.60698
R37692 C10_N_btm.n3186 C10_N_btm.n3185 4.60698
R37693 C10_N_btm.n3185 C10_N_btm.n3184 4.60698
R37694 C10_N_btm.n3183 C10_N_btm.n3182 4.60698
R37695 C10_N_btm.n3182 C10_N_btm.n3181 4.60698
R37696 C10_N_btm.n3180 C10_N_btm.n3179 4.60698
R37697 C10_N_btm.n3179 C10_N_btm.n3178 4.60698
R37698 C10_N_btm.n3177 C10_N_btm.n3176 4.60698
R37699 C10_N_btm.n3176 C10_N_btm.n3175 4.60698
R37700 C10_N_btm.n3174 C10_N_btm.n3173 4.60698
R37701 C10_N_btm.n3173 C10_N_btm.n3172 4.60698
R37702 C10_N_btm.n3171 C10_N_btm.n3170 4.60698
R37703 C10_N_btm.n3170 C10_N_btm.n3169 4.60698
R37704 C10_N_btm.n3168 C10_N_btm.n3167 4.60698
R37705 C10_N_btm.n3167 C10_N_btm.n3166 4.60698
R37706 C10_N_btm.n3165 C10_N_btm.n3164 4.60698
R37707 C10_N_btm.n3164 C10_N_btm.n3163 4.60698
R37708 C10_N_btm.n3162 C10_N_btm.n3161 4.60698
R37709 C10_N_btm.n3161 C10_N_btm.n3160 4.60698
R37710 C10_N_btm.n3159 C10_N_btm.n3158 4.60698
R37711 C10_N_btm.n3158 C10_N_btm.n3157 4.60698
R37712 C10_N_btm.n3156 C10_N_btm.n3155 4.60698
R37713 C10_N_btm.n3155 C10_N_btm.n3154 4.60698
R37714 C10_N_btm.n3153 C10_N_btm.n3152 4.60698
R37715 C10_N_btm.n3152 C10_N_btm.n3151 4.60698
R37716 C10_N_btm.n3150 C10_N_btm.n3149 4.60698
R37717 C10_N_btm.n3149 C10_N_btm.n3148 4.60698
R37718 C10_N_btm.n3147 C10_N_btm.n3146 4.60698
R37719 C10_N_btm.n3146 C10_N_btm.n3145 4.60698
R37720 C10_N_btm.n3144 C10_N_btm.n3143 4.60698
R37721 C10_N_btm.n3143 C10_N_btm.n3142 4.60698
R37722 C10_N_btm.n3141 C10_N_btm.n3140 4.60698
R37723 C10_N_btm.n3140 C10_N_btm.n3139 4.60698
R37724 C10_N_btm.n3138 C10_N_btm.n3137 4.60698
R37725 C10_N_btm.n3137 C10_N_btm.n3136 4.60698
R37726 C10_N_btm.n3135 C10_N_btm.n3134 4.60698
R37727 C10_N_btm.n3134 C10_N_btm.n3133 4.60698
R37728 C10_N_btm.n3132 C10_N_btm.n3131 4.60698
R37729 C10_N_btm.n3131 C10_N_btm.n3130 4.60698
R37730 C10_N_btm.n3129 C10_N_btm.n3128 4.60698
R37731 C10_N_btm.n3128 C10_N_btm.n3127 4.60698
R37732 C10_N_btm.n3126 C10_N_btm.n3125 4.60698
R37733 C10_N_btm.n3125 C10_N_btm.n3124 4.60698
R37734 C10_N_btm.n3123 C10_N_btm.n3122 4.60698
R37735 C10_N_btm.n3122 C10_N_btm.n3121 4.60698
R37736 C10_N_btm.n3120 C10_N_btm.n3119 4.60698
R37737 C10_N_btm.n3119 C10_N_btm.n3118 4.60698
R37738 C10_N_btm.n3117 C10_N_btm.n3116 4.60698
R37739 C10_N_btm.n3116 C10_N_btm.n3115 4.60698
R37740 C10_N_btm.n3114 C10_N_btm.n3113 4.60698
R37741 C10_N_btm.n3113 C10_N_btm.n3112 4.60698
R37742 C10_N_btm.n3111 C10_N_btm.n3110 4.60698
R37743 C10_N_btm.n3110 C10_N_btm.n3109 4.60698
R37744 C10_N_btm.n3103 C10_N_btm.n3102 4.60698
R37745 C10_N_btm.n3104 C10_N_btm.n3103 4.60698
R37746 C10_N_btm.n3100 C10_N_btm.n3099 4.60698
R37747 C10_N_btm.n3101 C10_N_btm.n3100 4.60698
R37748 C10_N_btm.n3097 C10_N_btm.n3096 4.60698
R37749 C10_N_btm.n3098 C10_N_btm.n3097 4.60698
R37750 C10_N_btm.n3094 C10_N_btm.n3093 4.60698
R37751 C10_N_btm.n3095 C10_N_btm.n3094 4.60698
R37752 C10_N_btm.n3091 C10_N_btm.n3090 4.60698
R37753 C10_N_btm.n3092 C10_N_btm.n3091 4.60698
R37754 C10_N_btm.n3088 C10_N_btm.n3087 4.60698
R37755 C10_N_btm.n3089 C10_N_btm.n3088 4.60698
R37756 C10_N_btm.n3085 C10_N_btm.n3084 4.60698
R37757 C10_N_btm.n3086 C10_N_btm.n3085 4.60698
R37758 C10_N_btm.n3082 C10_N_btm.n3081 4.60698
R37759 C10_N_btm.n3083 C10_N_btm.n3082 4.60698
R37760 C10_N_btm.n3079 C10_N_btm.n3078 4.60698
R37761 C10_N_btm.n3080 C10_N_btm.n3079 4.60698
R37762 C10_N_btm.n3076 C10_N_btm.n3075 4.60698
R37763 C10_N_btm.n3077 C10_N_btm.n3076 4.60698
R37764 C10_N_btm.n3073 C10_N_btm.n3072 4.60698
R37765 C10_N_btm.n3074 C10_N_btm.n3073 4.60698
R37766 C10_N_btm.n3070 C10_N_btm.n3069 4.60698
R37767 C10_N_btm.n3071 C10_N_btm.n3070 4.60698
R37768 C10_N_btm.n3067 C10_N_btm.n3066 4.60698
R37769 C10_N_btm.n3068 C10_N_btm.n3067 4.60698
R37770 C10_N_btm.n3064 C10_N_btm.n3063 4.60698
R37771 C10_N_btm.n3065 C10_N_btm.n3064 4.60698
R37772 C10_N_btm.n3061 C10_N_btm.n3060 4.60698
R37773 C10_N_btm.n3062 C10_N_btm.n3061 4.60698
R37774 C10_N_btm.n3058 C10_N_btm.n3057 4.60698
R37775 C10_N_btm.n3059 C10_N_btm.n3058 4.60698
R37776 C10_N_btm.n3055 C10_N_btm.n3054 4.60698
R37777 C10_N_btm.n3056 C10_N_btm.n3055 4.60698
R37778 C10_N_btm.n3052 C10_N_btm.n3051 4.60698
R37779 C10_N_btm.n3053 C10_N_btm.n3052 4.60698
R37780 C10_N_btm.n3049 C10_N_btm.n3048 4.60698
R37781 C10_N_btm.n3050 C10_N_btm.n3049 4.60698
R37782 C10_N_btm.n3046 C10_N_btm.n3045 4.60698
R37783 C10_N_btm.n3047 C10_N_btm.n3046 4.60698
R37784 C10_N_btm.n3043 C10_N_btm.n3042 4.60698
R37785 C10_N_btm.n3044 C10_N_btm.n3043 4.60698
R37786 C10_N_btm.n3040 C10_N_btm.n3039 4.60698
R37787 C10_N_btm.n3041 C10_N_btm.n3040 4.60698
R37788 C10_N_btm.n3037 C10_N_btm.n3036 4.60698
R37789 C10_N_btm.n3038 C10_N_btm.n3037 4.60698
R37790 C10_N_btm.n3034 C10_N_btm.n3033 4.60698
R37791 C10_N_btm.n3035 C10_N_btm.n3034 4.60698
R37792 C10_N_btm.n3031 C10_N_btm.n3030 4.60698
R37793 C10_N_btm.n3032 C10_N_btm.n3031 4.60698
R37794 C10_N_btm.n3028 C10_N_btm.n3027 4.60698
R37795 C10_N_btm.n3029 C10_N_btm.n3028 4.60698
R37796 C10_N_btm.n3025 C10_N_btm.n3024 4.60698
R37797 C10_N_btm.n3026 C10_N_btm.n3025 4.60698
R37798 C10_N_btm.n3022 C10_N_btm.n3021 4.60698
R37799 C10_N_btm.n3023 C10_N_btm.n3022 4.60698
R37800 C10_N_btm.n3019 C10_N_btm.n3018 4.60698
R37801 C10_N_btm.n3020 C10_N_btm.n3019 4.60698
R37802 C10_N_btm.n3016 C10_N_btm.n3015 4.60698
R37803 C10_N_btm.n3017 C10_N_btm.n3016 4.60698
R37804 C10_N_btm.n3013 C10_N_btm.n3012 4.60698
R37805 C10_N_btm.n3014 C10_N_btm.n3013 4.60698
R37806 C10_N_btm.n3010 C10_N_btm.n3009 4.60698
R37807 C10_N_btm.n3011 C10_N_btm.n3010 4.60698
R37808 C10_N_btm.n3007 C10_N_btm.n3006 4.60698
R37809 C10_N_btm.n3008 C10_N_btm.n3007 4.60698
R37810 C10_N_btm.n3004 C10_N_btm.n3003 4.60698
R37811 C10_N_btm.n3005 C10_N_btm.n3004 4.60698
R37812 C10_N_btm.n3001 C10_N_btm.n3000 4.60698
R37813 C10_N_btm.n3002 C10_N_btm.n3001 4.60698
R37814 C10_N_btm.n2998 C10_N_btm.n2997 4.60698
R37815 C10_N_btm.n2999 C10_N_btm.n2998 4.60698
R37816 C10_N_btm.n2995 C10_N_btm.n2994 4.60698
R37817 C10_N_btm.n2996 C10_N_btm.n2995 4.60698
R37818 C10_N_btm.n2992 C10_N_btm.n2991 4.60698
R37819 C10_N_btm.n2993 C10_N_btm.n2992 4.60698
R37820 C10_N_btm.n2989 C10_N_btm.n2988 4.60698
R37821 C10_N_btm.n2990 C10_N_btm.n2989 4.60698
R37822 C10_N_btm.n2986 C10_N_btm.n2985 4.60698
R37823 C10_N_btm.n2987 C10_N_btm.n2986 4.60698
R37824 C10_N_btm.n2983 C10_N_btm.n2982 4.60698
R37825 C10_N_btm.n2984 C10_N_btm.n2983 4.60698
R37826 C10_N_btm.n2980 C10_N_btm.n2979 4.60698
R37827 C10_N_btm.n2981 C10_N_btm.n2980 4.60698
R37828 C10_N_btm.n2977 C10_N_btm.n2976 4.60698
R37829 C10_N_btm.n2978 C10_N_btm.n2977 4.60698
R37830 C10_N_btm.n2974 C10_N_btm.n2973 4.60698
R37831 C10_N_btm.n2975 C10_N_btm.n2974 4.60698
R37832 C10_N_btm.n2971 C10_N_btm.n2970 4.60698
R37833 C10_N_btm.n2972 C10_N_btm.n2971 4.60698
R37834 C10_N_btm.n2968 C10_N_btm.n2967 4.60698
R37835 C10_N_btm.n2969 C10_N_btm.n2968 4.60698
R37836 C10_N_btm.n2965 C10_N_btm.n2964 4.60698
R37837 C10_N_btm.n2966 C10_N_btm.n2965 4.60698
R37838 C10_N_btm.n2962 C10_N_btm.n2961 4.60698
R37839 C10_N_btm.n2963 C10_N_btm.n2962 4.60698
R37840 C10_N_btm.n2959 C10_N_btm.n2958 4.60698
R37841 C10_N_btm.n2960 C10_N_btm.n2959 4.60698
R37842 C10_N_btm.n2956 C10_N_btm.n2955 4.60698
R37843 C10_N_btm.n2957 C10_N_btm.n2956 4.60698
R37844 C10_N_btm.n2953 C10_N_btm.n2952 4.60698
R37845 C10_N_btm.n2954 C10_N_btm.n2953 4.60698
R37846 C10_N_btm.n2950 C10_N_btm.n2949 4.60698
R37847 C10_N_btm.n2951 C10_N_btm.n2950 4.60698
R37848 C10_N_btm.n2947 C10_N_btm.n2946 4.60698
R37849 C10_N_btm.n2948 C10_N_btm.n2947 4.60698
R37850 C10_N_btm.n2944 C10_N_btm.n2943 4.60698
R37851 C10_N_btm.n2945 C10_N_btm.n2944 4.60698
R37852 C10_N_btm.n2941 C10_N_btm.n2940 4.60698
R37853 C10_N_btm.n2942 C10_N_btm.n2941 4.60698
R37854 C10_N_btm.n2938 C10_N_btm.n2937 4.60698
R37855 C10_N_btm.n2939 C10_N_btm.n2938 4.60698
R37856 C10_N_btm.n2935 C10_N_btm.n2934 4.60698
R37857 C10_N_btm.n2936 C10_N_btm.n2935 4.60698
R37858 C10_N_btm.n2932 C10_N_btm.n2931 4.60698
R37859 C10_N_btm.n2933 C10_N_btm.n2932 4.60698
R37860 C10_N_btm.n2929 C10_N_btm.n2928 4.60698
R37861 C10_N_btm.n2930 C10_N_btm.n2929 4.60698
R37862 C10_N_btm.n2926 C10_N_btm.n2925 4.60698
R37863 C10_N_btm.n2927 C10_N_btm.n2926 4.60698
R37864 C10_N_btm.n2923 C10_N_btm.n2922 4.60698
R37865 C10_N_btm.n2924 C10_N_btm.n2923 4.60698
R37866 C10_N_btm.n2920 C10_N_btm.n2919 4.60698
R37867 C10_N_btm.n2921 C10_N_btm.n2920 4.60698
R37868 C10_N_btm.n2915 C10_N_btm.n2914 4.60698
R37869 C10_N_btm.n2914 C10_N_btm.n1661 4.60698
R37870 C10_N_btm.n1786 C10_N_btm.n1785 4.60698
R37871 C10_N_btm.n1787 C10_N_btm.n1786 4.60698
R37872 C10_N_btm.n1789 C10_N_btm.n1788 4.60698
R37873 C10_N_btm.n1790 C10_N_btm.n1789 4.60698
R37874 C10_N_btm.n1792 C10_N_btm.n1791 4.60698
R37875 C10_N_btm.n1793 C10_N_btm.n1792 4.60698
R37876 C10_N_btm.n1795 C10_N_btm.n1794 4.60698
R37877 C10_N_btm.n1796 C10_N_btm.n1795 4.60698
R37878 C10_N_btm.n1798 C10_N_btm.n1797 4.60698
R37879 C10_N_btm.n1799 C10_N_btm.n1798 4.60698
R37880 C10_N_btm.n1801 C10_N_btm.n1800 4.60698
R37881 C10_N_btm.n1802 C10_N_btm.n1801 4.60698
R37882 C10_N_btm.n1804 C10_N_btm.n1803 4.60698
R37883 C10_N_btm.n1805 C10_N_btm.n1804 4.60698
R37884 C10_N_btm.n1807 C10_N_btm.n1806 4.60698
R37885 C10_N_btm.n1808 C10_N_btm.n1807 4.60698
R37886 C10_N_btm.n1810 C10_N_btm.n1809 4.60698
R37887 C10_N_btm.n1811 C10_N_btm.n1810 4.60698
R37888 C10_N_btm.n1813 C10_N_btm.n1812 4.60698
R37889 C10_N_btm.n1814 C10_N_btm.n1813 4.60698
R37890 C10_N_btm.n1816 C10_N_btm.n1815 4.60698
R37891 C10_N_btm.n1817 C10_N_btm.n1816 4.60698
R37892 C10_N_btm.n1819 C10_N_btm.n1818 4.60698
R37893 C10_N_btm.n1820 C10_N_btm.n1819 4.60698
R37894 C10_N_btm.n1822 C10_N_btm.n1821 4.60698
R37895 C10_N_btm.n1823 C10_N_btm.n1822 4.60698
R37896 C10_N_btm.n1825 C10_N_btm.n1824 4.60698
R37897 C10_N_btm.n1826 C10_N_btm.n1825 4.60698
R37898 C10_N_btm.n1828 C10_N_btm.n1827 4.60698
R37899 C10_N_btm.n1829 C10_N_btm.n1828 4.60698
R37900 C10_N_btm.n1831 C10_N_btm.n1830 4.60698
R37901 C10_N_btm.n1832 C10_N_btm.n1831 4.60698
R37902 C10_N_btm.n1834 C10_N_btm.n1833 4.60698
R37903 C10_N_btm.n1835 C10_N_btm.n1834 4.60698
R37904 C10_N_btm.n1837 C10_N_btm.n1836 4.60698
R37905 C10_N_btm.n1838 C10_N_btm.n1837 4.60698
R37906 C10_N_btm.n1840 C10_N_btm.n1839 4.60698
R37907 C10_N_btm.n1841 C10_N_btm.n1840 4.60698
R37908 C10_N_btm.n1843 C10_N_btm.n1842 4.60698
R37909 C10_N_btm.n1844 C10_N_btm.n1843 4.60698
R37910 C10_N_btm.n1846 C10_N_btm.n1845 4.60698
R37911 C10_N_btm.n1847 C10_N_btm.n1846 4.60698
R37912 C10_N_btm.n1849 C10_N_btm.n1848 4.60698
R37913 C10_N_btm.n1850 C10_N_btm.n1849 4.60698
R37914 C10_N_btm.n1852 C10_N_btm.n1851 4.60698
R37915 C10_N_btm.n1853 C10_N_btm.n1852 4.60698
R37916 C10_N_btm.n1855 C10_N_btm.n1854 4.60698
R37917 C10_N_btm.n1856 C10_N_btm.n1855 4.60698
R37918 C10_N_btm.n1858 C10_N_btm.n1857 4.60698
R37919 C10_N_btm.n1859 C10_N_btm.n1858 4.60698
R37920 C10_N_btm.n1861 C10_N_btm.n1860 4.60698
R37921 C10_N_btm.n1862 C10_N_btm.n1861 4.60698
R37922 C10_N_btm.n1864 C10_N_btm.n1863 4.60698
R37923 C10_N_btm.n1865 C10_N_btm.n1864 4.60698
R37924 C10_N_btm.n1867 C10_N_btm.n1866 4.60698
R37925 C10_N_btm.n1868 C10_N_btm.n1867 4.60698
R37926 C10_N_btm.n1870 C10_N_btm.n1869 4.60698
R37927 C10_N_btm.n1871 C10_N_btm.n1870 4.60698
R37928 C10_N_btm.n1873 C10_N_btm.n1872 4.60698
R37929 C10_N_btm.n1874 C10_N_btm.n1873 4.60698
R37930 C10_N_btm.n1876 C10_N_btm.n1875 4.60698
R37931 C10_N_btm.n1877 C10_N_btm.n1876 4.60698
R37932 C10_N_btm.n1879 C10_N_btm.n1878 4.60698
R37933 C10_N_btm.n1880 C10_N_btm.n1879 4.60698
R37934 C10_N_btm.n1882 C10_N_btm.n1881 4.60698
R37935 C10_N_btm.n1883 C10_N_btm.n1882 4.60698
R37936 C10_N_btm.n1885 C10_N_btm.n1884 4.60698
R37937 C10_N_btm.n1886 C10_N_btm.n1885 4.60698
R37938 C10_N_btm.n1888 C10_N_btm.n1887 4.60698
R37939 C10_N_btm.n1889 C10_N_btm.n1888 4.60698
R37940 C10_N_btm.n1891 C10_N_btm.n1890 4.60698
R37941 C10_N_btm.n1892 C10_N_btm.n1891 4.60698
R37942 C10_N_btm.n1894 C10_N_btm.n1893 4.60698
R37943 C10_N_btm.n1895 C10_N_btm.n1894 4.60698
R37944 C10_N_btm.n1897 C10_N_btm.n1896 4.60698
R37945 C10_N_btm.n1898 C10_N_btm.n1897 4.60698
R37946 C10_N_btm.n1900 C10_N_btm.n1899 4.60698
R37947 C10_N_btm.n1901 C10_N_btm.n1900 4.60698
R37948 C10_N_btm.n1903 C10_N_btm.n1902 4.60698
R37949 C10_N_btm.n1904 C10_N_btm.n1903 4.60698
R37950 C10_N_btm.n1906 C10_N_btm.n1905 4.60698
R37951 C10_N_btm.n1907 C10_N_btm.n1906 4.60698
R37952 C10_N_btm.n1909 C10_N_btm.n1908 4.60698
R37953 C10_N_btm.n1910 C10_N_btm.n1909 4.60698
R37954 C10_N_btm.n1912 C10_N_btm.n1911 4.60698
R37955 C10_N_btm.n1913 C10_N_btm.n1912 4.60698
R37956 C10_N_btm.n1915 C10_N_btm.n1914 4.60698
R37957 C10_N_btm.n1916 C10_N_btm.n1915 4.60698
R37958 C10_N_btm.n1918 C10_N_btm.n1917 4.60698
R37959 C10_N_btm.n1919 C10_N_btm.n1918 4.60698
R37960 C10_N_btm.n1921 C10_N_btm.n1920 4.60698
R37961 C10_N_btm.n1922 C10_N_btm.n1921 4.60698
R37962 C10_N_btm.n1924 C10_N_btm.n1923 4.60698
R37963 C10_N_btm.n1925 C10_N_btm.n1924 4.60698
R37964 C10_N_btm.n1927 C10_N_btm.n1926 4.60698
R37965 C10_N_btm.n1928 C10_N_btm.n1927 4.60698
R37966 C10_N_btm.n1930 C10_N_btm.n1929 4.60698
R37967 C10_N_btm.n1931 C10_N_btm.n1930 4.60698
R37968 C10_N_btm.n1933 C10_N_btm.n1932 4.60698
R37969 C10_N_btm.n1934 C10_N_btm.n1933 4.60698
R37970 C10_N_btm.n1936 C10_N_btm.n1935 4.60698
R37971 C10_N_btm.n1937 C10_N_btm.n1936 4.60698
R37972 C10_N_btm.n1939 C10_N_btm.n1938 4.60698
R37973 C10_N_btm.n1940 C10_N_btm.n1939 4.60698
R37974 C10_N_btm.n1942 C10_N_btm.n1941 4.60698
R37975 C10_N_btm.n1943 C10_N_btm.n1942 4.60698
R37976 C10_N_btm.n1945 C10_N_btm.n1944 4.60698
R37977 C10_N_btm.n1946 C10_N_btm.n1945 4.60698
R37978 C10_N_btm.n1948 C10_N_btm.n1947 4.60698
R37979 C10_N_btm.n1949 C10_N_btm.n1948 4.60698
R37980 C10_N_btm.n1951 C10_N_btm.n1950 4.60698
R37981 C10_N_btm.n1952 C10_N_btm.n1951 4.60698
R37982 C10_N_btm.n1954 C10_N_btm.n1953 4.60698
R37983 C10_N_btm.n1955 C10_N_btm.n1954 4.60698
R37984 C10_N_btm.n1957 C10_N_btm.n1956 4.60698
R37985 C10_N_btm.n1958 C10_N_btm.n1957 4.60698
R37986 C10_N_btm.n1960 C10_N_btm.n1959 4.60698
R37987 C10_N_btm.n1961 C10_N_btm.n1960 4.60698
R37988 C10_N_btm.n1963 C10_N_btm.n1962 4.60698
R37989 C10_N_btm.n1964 C10_N_btm.n1963 4.60698
R37990 C10_N_btm.n1966 C10_N_btm.n1965 4.60698
R37991 C10_N_btm.n1965 C10_N_btm.n1724 4.60698
R37992 C10_N_btm.n2726 C10_N_btm.n2725 4.60698
R37993 C10_N_btm.n2725 C10_N_btm.n2724 4.60698
R37994 C10_N_btm.n2729 C10_N_btm.n2728 4.60698
R37995 C10_N_btm.n2728 C10_N_btm.n2727 4.60698
R37996 C10_N_btm.n2732 C10_N_btm.n2731 4.60698
R37997 C10_N_btm.n2731 C10_N_btm.n2730 4.60698
R37998 C10_N_btm.n2735 C10_N_btm.n2734 4.60698
R37999 C10_N_btm.n2734 C10_N_btm.n2733 4.60698
R38000 C10_N_btm.n2738 C10_N_btm.n2737 4.60698
R38001 C10_N_btm.n2737 C10_N_btm.n2736 4.60698
R38002 C10_N_btm.n2741 C10_N_btm.n2740 4.60698
R38003 C10_N_btm.n2740 C10_N_btm.n2739 4.60698
R38004 C10_N_btm.n2744 C10_N_btm.n2743 4.60698
R38005 C10_N_btm.n2743 C10_N_btm.n2742 4.60698
R38006 C10_N_btm.n2747 C10_N_btm.n2746 4.60698
R38007 C10_N_btm.n2746 C10_N_btm.n2745 4.60698
R38008 C10_N_btm.n2750 C10_N_btm.n2749 4.60698
R38009 C10_N_btm.n2749 C10_N_btm.n2748 4.60698
R38010 C10_N_btm.n2753 C10_N_btm.n2752 4.60698
R38011 C10_N_btm.n2752 C10_N_btm.n2751 4.60698
R38012 C10_N_btm.n2756 C10_N_btm.n2755 4.60698
R38013 C10_N_btm.n2755 C10_N_btm.n2754 4.60698
R38014 C10_N_btm.n2759 C10_N_btm.n2758 4.60698
R38015 C10_N_btm.n2758 C10_N_btm.n2757 4.60698
R38016 C10_N_btm.n2762 C10_N_btm.n2761 4.60698
R38017 C10_N_btm.n2761 C10_N_btm.n2760 4.60698
R38018 C10_N_btm.n2765 C10_N_btm.n2764 4.60698
R38019 C10_N_btm.n2764 C10_N_btm.n2763 4.60698
R38020 C10_N_btm.n2768 C10_N_btm.n2767 4.60698
R38021 C10_N_btm.n2767 C10_N_btm.n2766 4.60698
R38022 C10_N_btm.n2771 C10_N_btm.n2770 4.60698
R38023 C10_N_btm.n2770 C10_N_btm.n2769 4.60698
R38024 C10_N_btm.n2774 C10_N_btm.n2773 4.60698
R38025 C10_N_btm.n2773 C10_N_btm.n2772 4.60698
R38026 C10_N_btm.n2777 C10_N_btm.n2776 4.60698
R38027 C10_N_btm.n2776 C10_N_btm.n2775 4.60698
R38028 C10_N_btm.n2780 C10_N_btm.n2779 4.60698
R38029 C10_N_btm.n2779 C10_N_btm.n2778 4.60698
R38030 C10_N_btm.n2783 C10_N_btm.n2782 4.60698
R38031 C10_N_btm.n2782 C10_N_btm.n2781 4.60698
R38032 C10_N_btm.n2786 C10_N_btm.n2785 4.60698
R38033 C10_N_btm.n2785 C10_N_btm.n2784 4.60698
R38034 C10_N_btm.n2789 C10_N_btm.n2788 4.60698
R38035 C10_N_btm.n2788 C10_N_btm.n2787 4.60698
R38036 C10_N_btm.n2792 C10_N_btm.n2791 4.60698
R38037 C10_N_btm.n2791 C10_N_btm.n2790 4.60698
R38038 C10_N_btm.n2795 C10_N_btm.n2794 4.60698
R38039 C10_N_btm.n2794 C10_N_btm.n2793 4.60698
R38040 C10_N_btm.n2798 C10_N_btm.n2797 4.60698
R38041 C10_N_btm.n2797 C10_N_btm.n2796 4.60698
R38042 C10_N_btm.n2801 C10_N_btm.n2800 4.60698
R38043 C10_N_btm.n2800 C10_N_btm.n2799 4.60698
R38044 C10_N_btm.n2804 C10_N_btm.n2803 4.60698
R38045 C10_N_btm.n2803 C10_N_btm.n2802 4.60698
R38046 C10_N_btm.n2807 C10_N_btm.n2806 4.60698
R38047 C10_N_btm.n2806 C10_N_btm.n2805 4.60698
R38048 C10_N_btm.n2810 C10_N_btm.n2809 4.60698
R38049 C10_N_btm.n2809 C10_N_btm.n2808 4.60698
R38050 C10_N_btm.n2813 C10_N_btm.n2812 4.60698
R38051 C10_N_btm.n2812 C10_N_btm.n2811 4.60698
R38052 C10_N_btm.n2816 C10_N_btm.n2815 4.60698
R38053 C10_N_btm.n2815 C10_N_btm.n2814 4.60698
R38054 C10_N_btm.n2819 C10_N_btm.n2818 4.60698
R38055 C10_N_btm.n2818 C10_N_btm.n2817 4.60698
R38056 C10_N_btm.n2822 C10_N_btm.n2821 4.60698
R38057 C10_N_btm.n2821 C10_N_btm.n2820 4.60698
R38058 C10_N_btm.n2825 C10_N_btm.n2824 4.60698
R38059 C10_N_btm.n2824 C10_N_btm.n2823 4.60698
R38060 C10_N_btm.n2828 C10_N_btm.n2827 4.60698
R38061 C10_N_btm.n2827 C10_N_btm.n2826 4.60698
R38062 C10_N_btm.n2831 C10_N_btm.n2830 4.60698
R38063 C10_N_btm.n2830 C10_N_btm.n2829 4.60698
R38064 C10_N_btm.n2834 C10_N_btm.n2833 4.60698
R38065 C10_N_btm.n2833 C10_N_btm.n2832 4.60698
R38066 C10_N_btm.n2837 C10_N_btm.n2836 4.60698
R38067 C10_N_btm.n2836 C10_N_btm.n2835 4.60698
R38068 C10_N_btm.n2840 C10_N_btm.n2839 4.60698
R38069 C10_N_btm.n2839 C10_N_btm.n2838 4.60698
R38070 C10_N_btm.n2843 C10_N_btm.n2842 4.60698
R38071 C10_N_btm.n2842 C10_N_btm.n2841 4.60698
R38072 C10_N_btm.n2846 C10_N_btm.n2845 4.60698
R38073 C10_N_btm.n2845 C10_N_btm.n2844 4.60698
R38074 C10_N_btm.n2849 C10_N_btm.n2848 4.60698
R38075 C10_N_btm.n2848 C10_N_btm.n2847 4.60698
R38076 C10_N_btm.n2852 C10_N_btm.n2851 4.60698
R38077 C10_N_btm.n2851 C10_N_btm.n2850 4.60698
R38078 C10_N_btm.n2855 C10_N_btm.n2854 4.60698
R38079 C10_N_btm.n2854 C10_N_btm.n2853 4.60698
R38080 C10_N_btm.n2858 C10_N_btm.n2857 4.60698
R38081 C10_N_btm.n2857 C10_N_btm.n2856 4.60698
R38082 C10_N_btm.n2861 C10_N_btm.n2860 4.60698
R38083 C10_N_btm.n2860 C10_N_btm.n2859 4.60698
R38084 C10_N_btm.n2864 C10_N_btm.n2863 4.60698
R38085 C10_N_btm.n2863 C10_N_btm.n2862 4.60698
R38086 C10_N_btm.n2867 C10_N_btm.n2866 4.60698
R38087 C10_N_btm.n2866 C10_N_btm.n2865 4.60698
R38088 C10_N_btm.n2870 C10_N_btm.n2869 4.60698
R38089 C10_N_btm.n2869 C10_N_btm.n2868 4.60698
R38090 C10_N_btm.n2873 C10_N_btm.n2872 4.60698
R38091 C10_N_btm.n2872 C10_N_btm.n2871 4.60698
R38092 C10_N_btm.n2876 C10_N_btm.n2875 4.60698
R38093 C10_N_btm.n2875 C10_N_btm.n2874 4.60698
R38094 C10_N_btm.n2879 C10_N_btm.n2878 4.60698
R38095 C10_N_btm.n2878 C10_N_btm.n2877 4.60698
R38096 C10_N_btm.n2882 C10_N_btm.n2881 4.60698
R38097 C10_N_btm.n2881 C10_N_btm.n2880 4.60698
R38098 C10_N_btm.n2885 C10_N_btm.n2884 4.60698
R38099 C10_N_btm.n2884 C10_N_btm.n2883 4.60698
R38100 C10_N_btm.n2888 C10_N_btm.n2887 4.60698
R38101 C10_N_btm.n2887 C10_N_btm.n2886 4.60698
R38102 C10_N_btm.n2891 C10_N_btm.n2890 4.60698
R38103 C10_N_btm.n2890 C10_N_btm.n2889 4.60698
R38104 C10_N_btm.n2894 C10_N_btm.n2893 4.60698
R38105 C10_N_btm.n2893 C10_N_btm.n2892 4.60698
R38106 C10_N_btm.n2897 C10_N_btm.n2896 4.60698
R38107 C10_N_btm.n2896 C10_N_btm.n2895 4.60698
R38108 C10_N_btm.n2900 C10_N_btm.n2899 4.60698
R38109 C10_N_btm.n2899 C10_N_btm.n2898 4.60698
R38110 C10_N_btm.n2903 C10_N_btm.n2902 4.60698
R38111 C10_N_btm.n2902 C10_N_btm.n2901 4.60698
R38112 C10_N_btm.n2906 C10_N_btm.n2905 4.60698
R38113 C10_N_btm.n2905 C10_N_btm.n2904 4.60698
R38114 C10_N_btm.n2909 C10_N_btm.n2908 4.60698
R38115 C10_N_btm.n2908 C10_N_btm.n2907 4.60698
R38116 C10_N_btm.n2535 C10_N_btm.n2534 4.60698
R38117 C10_N_btm.n2536 C10_N_btm.n2535 4.60698
R38118 C10_N_btm.n2538 C10_N_btm.n2537 4.60698
R38119 C10_N_btm.n2539 C10_N_btm.n2538 4.60698
R38120 C10_N_btm.n2541 C10_N_btm.n2540 4.60698
R38121 C10_N_btm.n2542 C10_N_btm.n2541 4.60698
R38122 C10_N_btm.n2544 C10_N_btm.n2543 4.60698
R38123 C10_N_btm.n2545 C10_N_btm.n2544 4.60698
R38124 C10_N_btm.n2547 C10_N_btm.n2546 4.60698
R38125 C10_N_btm.n2548 C10_N_btm.n2547 4.60698
R38126 C10_N_btm.n2550 C10_N_btm.n2549 4.60698
R38127 C10_N_btm.n2551 C10_N_btm.n2550 4.60698
R38128 C10_N_btm.n2553 C10_N_btm.n2552 4.60698
R38129 C10_N_btm.n2554 C10_N_btm.n2553 4.60698
R38130 C10_N_btm.n2556 C10_N_btm.n2555 4.60698
R38131 C10_N_btm.n2557 C10_N_btm.n2556 4.60698
R38132 C10_N_btm.n2559 C10_N_btm.n2558 4.60698
R38133 C10_N_btm.n2560 C10_N_btm.n2559 4.60698
R38134 C10_N_btm.n2562 C10_N_btm.n2561 4.60698
R38135 C10_N_btm.n2563 C10_N_btm.n2562 4.60698
R38136 C10_N_btm.n2565 C10_N_btm.n2564 4.60698
R38137 C10_N_btm.n2566 C10_N_btm.n2565 4.60698
R38138 C10_N_btm.n2568 C10_N_btm.n2567 4.60698
R38139 C10_N_btm.n2569 C10_N_btm.n2568 4.60698
R38140 C10_N_btm.n2571 C10_N_btm.n2570 4.60698
R38141 C10_N_btm.n2572 C10_N_btm.n2571 4.60698
R38142 C10_N_btm.n2574 C10_N_btm.n2573 4.60698
R38143 C10_N_btm.n2575 C10_N_btm.n2574 4.60698
R38144 C10_N_btm.n2577 C10_N_btm.n2576 4.60698
R38145 C10_N_btm.n2578 C10_N_btm.n2577 4.60698
R38146 C10_N_btm.n2580 C10_N_btm.n2579 4.60698
R38147 C10_N_btm.n2581 C10_N_btm.n2580 4.60698
R38148 C10_N_btm.n2583 C10_N_btm.n2582 4.60698
R38149 C10_N_btm.n2584 C10_N_btm.n2583 4.60698
R38150 C10_N_btm.n2586 C10_N_btm.n2585 4.60698
R38151 C10_N_btm.n2587 C10_N_btm.n2586 4.60698
R38152 C10_N_btm.n2589 C10_N_btm.n2588 4.60698
R38153 C10_N_btm.n2590 C10_N_btm.n2589 4.60698
R38154 C10_N_btm.n2592 C10_N_btm.n2591 4.60698
R38155 C10_N_btm.n2593 C10_N_btm.n2592 4.60698
R38156 C10_N_btm.n2595 C10_N_btm.n2594 4.60698
R38157 C10_N_btm.n2596 C10_N_btm.n2595 4.60698
R38158 C10_N_btm.n2598 C10_N_btm.n2597 4.60698
R38159 C10_N_btm.n2599 C10_N_btm.n2598 4.60698
R38160 C10_N_btm.n2601 C10_N_btm.n2600 4.60698
R38161 C10_N_btm.n2602 C10_N_btm.n2601 4.60698
R38162 C10_N_btm.n2604 C10_N_btm.n2603 4.60698
R38163 C10_N_btm.n2605 C10_N_btm.n2604 4.60698
R38164 C10_N_btm.n2607 C10_N_btm.n2606 4.60698
R38165 C10_N_btm.n2608 C10_N_btm.n2607 4.60698
R38166 C10_N_btm.n2610 C10_N_btm.n2609 4.60698
R38167 C10_N_btm.n2611 C10_N_btm.n2610 4.60698
R38168 C10_N_btm.n2613 C10_N_btm.n2612 4.60698
R38169 C10_N_btm.n2614 C10_N_btm.n2613 4.60698
R38170 C10_N_btm.n2616 C10_N_btm.n2615 4.60698
R38171 C10_N_btm.n2617 C10_N_btm.n2616 4.60698
R38172 C10_N_btm.n2619 C10_N_btm.n2618 4.60698
R38173 C10_N_btm.n2620 C10_N_btm.n2619 4.60698
R38174 C10_N_btm.n2622 C10_N_btm.n2621 4.60698
R38175 C10_N_btm.n2623 C10_N_btm.n2622 4.60698
R38176 C10_N_btm.n2625 C10_N_btm.n2624 4.60698
R38177 C10_N_btm.n2626 C10_N_btm.n2625 4.60698
R38178 C10_N_btm.n2628 C10_N_btm.n2627 4.60698
R38179 C10_N_btm.n2629 C10_N_btm.n2628 4.60698
R38180 C10_N_btm.n2631 C10_N_btm.n2630 4.60698
R38181 C10_N_btm.n2632 C10_N_btm.n2631 4.60698
R38182 C10_N_btm.n2634 C10_N_btm.n2633 4.60698
R38183 C10_N_btm.n2635 C10_N_btm.n2634 4.60698
R38184 C10_N_btm.n2637 C10_N_btm.n2636 4.60698
R38185 C10_N_btm.n2638 C10_N_btm.n2637 4.60698
R38186 C10_N_btm.n2640 C10_N_btm.n2639 4.60698
R38187 C10_N_btm.n2641 C10_N_btm.n2640 4.60698
R38188 C10_N_btm.n2643 C10_N_btm.n2642 4.60698
R38189 C10_N_btm.n2644 C10_N_btm.n2643 4.60698
R38190 C10_N_btm.n2646 C10_N_btm.n2645 4.60698
R38191 C10_N_btm.n2647 C10_N_btm.n2646 4.60698
R38192 C10_N_btm.n2649 C10_N_btm.n2648 4.60698
R38193 C10_N_btm.n2650 C10_N_btm.n2649 4.60698
R38194 C10_N_btm.n2652 C10_N_btm.n2651 4.60698
R38195 C10_N_btm.n2653 C10_N_btm.n2652 4.60698
R38196 C10_N_btm.n2655 C10_N_btm.n2654 4.60698
R38197 C10_N_btm.n2656 C10_N_btm.n2655 4.60698
R38198 C10_N_btm.n2658 C10_N_btm.n2657 4.60698
R38199 C10_N_btm.n2659 C10_N_btm.n2658 4.60698
R38200 C10_N_btm.n2661 C10_N_btm.n2660 4.60698
R38201 C10_N_btm.n2662 C10_N_btm.n2661 4.60698
R38202 C10_N_btm.n2664 C10_N_btm.n2663 4.60698
R38203 C10_N_btm.n2665 C10_N_btm.n2664 4.60698
R38204 C10_N_btm.n2667 C10_N_btm.n2666 4.60698
R38205 C10_N_btm.n2668 C10_N_btm.n2667 4.60698
R38206 C10_N_btm.n2670 C10_N_btm.n2669 4.60698
R38207 C10_N_btm.n2671 C10_N_btm.n2670 4.60698
R38208 C10_N_btm.n2673 C10_N_btm.n2672 4.60698
R38209 C10_N_btm.n2674 C10_N_btm.n2673 4.60698
R38210 C10_N_btm.n2676 C10_N_btm.n2675 4.60698
R38211 C10_N_btm.n2677 C10_N_btm.n2676 4.60698
R38212 C10_N_btm.n2679 C10_N_btm.n2678 4.60698
R38213 C10_N_btm.n2680 C10_N_btm.n2679 4.60698
R38214 C10_N_btm.n2682 C10_N_btm.n2681 4.60698
R38215 C10_N_btm.n2683 C10_N_btm.n2682 4.60698
R38216 C10_N_btm.n2685 C10_N_btm.n2684 4.60698
R38217 C10_N_btm.n2686 C10_N_btm.n2685 4.60698
R38218 C10_N_btm.n2688 C10_N_btm.n2687 4.60698
R38219 C10_N_btm.n2689 C10_N_btm.n2688 4.60698
R38220 C10_N_btm.n2691 C10_N_btm.n2690 4.60698
R38221 C10_N_btm.n2692 C10_N_btm.n2691 4.60698
R38222 C10_N_btm.n2694 C10_N_btm.n2693 4.60698
R38223 C10_N_btm.n2695 C10_N_btm.n2694 4.60698
R38224 C10_N_btm.n2697 C10_N_btm.n2696 4.60698
R38225 C10_N_btm.n2698 C10_N_btm.n2697 4.60698
R38226 C10_N_btm.n2700 C10_N_btm.n2699 4.60698
R38227 C10_N_btm.n2701 C10_N_btm.n2700 4.60698
R38228 C10_N_btm.n2703 C10_N_btm.n2702 4.60698
R38229 C10_N_btm.n2704 C10_N_btm.n2703 4.60698
R38230 C10_N_btm.n2706 C10_N_btm.n2705 4.60698
R38231 C10_N_btm.n2707 C10_N_btm.n2706 4.60698
R38232 C10_N_btm.n2709 C10_N_btm.n2708 4.60698
R38233 C10_N_btm.n2710 C10_N_btm.n2709 4.60698
R38234 C10_N_btm.n2712 C10_N_btm.n2711 4.60698
R38235 C10_N_btm.n2713 C10_N_btm.n2712 4.60698
R38236 C10_N_btm.n2715 C10_N_btm.n2714 4.60698
R38237 C10_N_btm.n2716 C10_N_btm.n2715 4.60698
R38238 C10_N_btm.n2718 C10_N_btm.n2717 4.60698
R38239 C10_N_btm.n2719 C10_N_btm.n2718 4.60698
R38240 C10_N_btm.n2336 C10_N_btm.n2335 4.60698
R38241 C10_N_btm.n2335 C10_N_btm.n2094 4.60698
R38242 C10_N_btm.n2333 C10_N_btm.n2332 4.60698
R38243 C10_N_btm.n2334 C10_N_btm.n2333 4.60698
R38244 C10_N_btm.n2330 C10_N_btm.n2329 4.60698
R38245 C10_N_btm.n2331 C10_N_btm.n2330 4.60698
R38246 C10_N_btm.n2327 C10_N_btm.n2326 4.60698
R38247 C10_N_btm.n2328 C10_N_btm.n2327 4.60698
R38248 C10_N_btm.n2324 C10_N_btm.n2323 4.60698
R38249 C10_N_btm.n2325 C10_N_btm.n2324 4.60698
R38250 C10_N_btm.n2321 C10_N_btm.n2320 4.60698
R38251 C10_N_btm.n2322 C10_N_btm.n2321 4.60698
R38252 C10_N_btm.n2318 C10_N_btm.n2317 4.60698
R38253 C10_N_btm.n2319 C10_N_btm.n2318 4.60698
R38254 C10_N_btm.n2315 C10_N_btm.n2314 4.60698
R38255 C10_N_btm.n2316 C10_N_btm.n2315 4.60698
R38256 C10_N_btm.n2312 C10_N_btm.n2311 4.60698
R38257 C10_N_btm.n2313 C10_N_btm.n2312 4.60698
R38258 C10_N_btm.n2309 C10_N_btm.n2308 4.60698
R38259 C10_N_btm.n2310 C10_N_btm.n2309 4.60698
R38260 C10_N_btm.n2306 C10_N_btm.n2305 4.60698
R38261 C10_N_btm.n2307 C10_N_btm.n2306 4.60698
R38262 C10_N_btm.n2303 C10_N_btm.n2302 4.60698
R38263 C10_N_btm.n2304 C10_N_btm.n2303 4.60698
R38264 C10_N_btm.n2300 C10_N_btm.n2299 4.60698
R38265 C10_N_btm.n2301 C10_N_btm.n2300 4.60698
R38266 C10_N_btm.n2297 C10_N_btm.n2296 4.60698
R38267 C10_N_btm.n2298 C10_N_btm.n2297 4.60698
R38268 C10_N_btm.n2294 C10_N_btm.n2293 4.60698
R38269 C10_N_btm.n2295 C10_N_btm.n2294 4.60698
R38270 C10_N_btm.n2291 C10_N_btm.n2290 4.60698
R38271 C10_N_btm.n2292 C10_N_btm.n2291 4.60698
R38272 C10_N_btm.n2288 C10_N_btm.n2287 4.60698
R38273 C10_N_btm.n2289 C10_N_btm.n2288 4.60698
R38274 C10_N_btm.n2285 C10_N_btm.n2284 4.60698
R38275 C10_N_btm.n2286 C10_N_btm.n2285 4.60698
R38276 C10_N_btm.n2282 C10_N_btm.n2281 4.60698
R38277 C10_N_btm.n2283 C10_N_btm.n2282 4.60698
R38278 C10_N_btm.n2279 C10_N_btm.n2278 4.60698
R38279 C10_N_btm.n2280 C10_N_btm.n2279 4.60698
R38280 C10_N_btm.n2276 C10_N_btm.n2275 4.60698
R38281 C10_N_btm.n2277 C10_N_btm.n2276 4.60698
R38282 C10_N_btm.n2273 C10_N_btm.n2272 4.60698
R38283 C10_N_btm.n2274 C10_N_btm.n2273 4.60698
R38284 C10_N_btm.n2270 C10_N_btm.n2269 4.60698
R38285 C10_N_btm.n2271 C10_N_btm.n2270 4.60698
R38286 C10_N_btm.n2267 C10_N_btm.n2266 4.60698
R38287 C10_N_btm.n2268 C10_N_btm.n2267 4.60698
R38288 C10_N_btm.n2264 C10_N_btm.n2263 4.60698
R38289 C10_N_btm.n2265 C10_N_btm.n2264 4.60698
R38290 C10_N_btm.n2261 C10_N_btm.n2260 4.60698
R38291 C10_N_btm.n2262 C10_N_btm.n2261 4.60698
R38292 C10_N_btm.n2258 C10_N_btm.n2257 4.60698
R38293 C10_N_btm.n2259 C10_N_btm.n2258 4.60698
R38294 C10_N_btm.n2255 C10_N_btm.n2254 4.60698
R38295 C10_N_btm.n2256 C10_N_btm.n2255 4.60698
R38296 C10_N_btm.n2252 C10_N_btm.n2251 4.60698
R38297 C10_N_btm.n2253 C10_N_btm.n2252 4.60698
R38298 C10_N_btm.n2249 C10_N_btm.n2248 4.60698
R38299 C10_N_btm.n2250 C10_N_btm.n2249 4.60698
R38300 C10_N_btm.n2246 C10_N_btm.n2245 4.60698
R38301 C10_N_btm.n2247 C10_N_btm.n2246 4.60698
R38302 C10_N_btm.n2243 C10_N_btm.n2242 4.60698
R38303 C10_N_btm.n2244 C10_N_btm.n2243 4.60698
R38304 C10_N_btm.n2240 C10_N_btm.n2239 4.60698
R38305 C10_N_btm.n2241 C10_N_btm.n2240 4.60698
R38306 C10_N_btm.n2237 C10_N_btm.n2236 4.60698
R38307 C10_N_btm.n2238 C10_N_btm.n2237 4.60698
R38308 C10_N_btm.n2234 C10_N_btm.n2233 4.60698
R38309 C10_N_btm.n2235 C10_N_btm.n2234 4.60698
R38310 C10_N_btm.n2231 C10_N_btm.n2230 4.60698
R38311 C10_N_btm.n2232 C10_N_btm.n2231 4.60698
R38312 C10_N_btm.n2228 C10_N_btm.n2227 4.60698
R38313 C10_N_btm.n2229 C10_N_btm.n2228 4.60698
R38314 C10_N_btm.n2225 C10_N_btm.n2224 4.60698
R38315 C10_N_btm.n2226 C10_N_btm.n2225 4.60698
R38316 C10_N_btm.n2222 C10_N_btm.n2221 4.60698
R38317 C10_N_btm.n2223 C10_N_btm.n2222 4.60698
R38318 C10_N_btm.n2219 C10_N_btm.n2218 4.60698
R38319 C10_N_btm.n2220 C10_N_btm.n2219 4.60698
R38320 C10_N_btm.n2216 C10_N_btm.n2215 4.60698
R38321 C10_N_btm.n2217 C10_N_btm.n2216 4.60698
R38322 C10_N_btm.n2213 C10_N_btm.n2212 4.60698
R38323 C10_N_btm.n2214 C10_N_btm.n2213 4.60698
R38324 C10_N_btm.n2210 C10_N_btm.n2209 4.60698
R38325 C10_N_btm.n2211 C10_N_btm.n2210 4.60698
R38326 C10_N_btm.n2207 C10_N_btm.n2206 4.60698
R38327 C10_N_btm.n2208 C10_N_btm.n2207 4.60698
R38328 C10_N_btm.n2204 C10_N_btm.n2203 4.60698
R38329 C10_N_btm.n2205 C10_N_btm.n2204 4.60698
R38330 C10_N_btm.n2201 C10_N_btm.n2200 4.60698
R38331 C10_N_btm.n2202 C10_N_btm.n2201 4.60698
R38332 C10_N_btm.n2198 C10_N_btm.n2197 4.60698
R38333 C10_N_btm.n2199 C10_N_btm.n2198 4.60698
R38334 C10_N_btm.n2195 C10_N_btm.n2194 4.60698
R38335 C10_N_btm.n2196 C10_N_btm.n2195 4.60698
R38336 C10_N_btm.n2192 C10_N_btm.n2191 4.60698
R38337 C10_N_btm.n2193 C10_N_btm.n2192 4.60698
R38338 C10_N_btm.n2189 C10_N_btm.n2188 4.60698
R38339 C10_N_btm.n2190 C10_N_btm.n2189 4.60698
R38340 C10_N_btm.n2186 C10_N_btm.n2185 4.60698
R38341 C10_N_btm.n2187 C10_N_btm.n2186 4.60698
R38342 C10_N_btm.n2183 C10_N_btm.n2182 4.60698
R38343 C10_N_btm.n2184 C10_N_btm.n2183 4.60698
R38344 C10_N_btm.n2180 C10_N_btm.n2179 4.60698
R38345 C10_N_btm.n2181 C10_N_btm.n2180 4.60698
R38346 C10_N_btm.n2177 C10_N_btm.n2176 4.60698
R38347 C10_N_btm.n2178 C10_N_btm.n2177 4.60698
R38348 C10_N_btm.n2174 C10_N_btm.n2173 4.60698
R38349 C10_N_btm.n2175 C10_N_btm.n2174 4.60698
R38350 C10_N_btm.n2171 C10_N_btm.n2170 4.60698
R38351 C10_N_btm.n2172 C10_N_btm.n2171 4.60698
R38352 C10_N_btm.n2168 C10_N_btm.n2167 4.60698
R38353 C10_N_btm.n2169 C10_N_btm.n2168 4.60698
R38354 C10_N_btm.n2165 C10_N_btm.n2164 4.60698
R38355 C10_N_btm.n2166 C10_N_btm.n2165 4.60698
R38356 C10_N_btm.n2162 C10_N_btm.n2161 4.60698
R38357 C10_N_btm.n2163 C10_N_btm.n2162 4.60698
R38358 C10_N_btm.n2159 C10_N_btm.n2158 4.60698
R38359 C10_N_btm.n2160 C10_N_btm.n2159 4.60698
R38360 C10_N_btm.n2156 C10_N_btm.n2155 4.60698
R38361 C10_N_btm.n2157 C10_N_btm.n2156 4.60698
R38362 C10_N_btm.n2530 C10_N_btm.n2529 4.60698
R38363 C10_N_btm.n2529 C10_N_btm.n2032 4.60698
R38364 C10_N_btm.n2524 C10_N_btm.n2523 4.60698
R38365 C10_N_btm.n2525 C10_N_btm.n2524 4.60698
R38366 C10_N_btm.n2521 C10_N_btm.n2520 4.60698
R38367 C10_N_btm.n2522 C10_N_btm.n2521 4.60698
R38368 C10_N_btm.n2518 C10_N_btm.n2517 4.60698
R38369 C10_N_btm.n2519 C10_N_btm.n2518 4.60698
R38370 C10_N_btm.n2515 C10_N_btm.n2514 4.60698
R38371 C10_N_btm.n2516 C10_N_btm.n2515 4.60698
R38372 C10_N_btm.n2512 C10_N_btm.n2511 4.60698
R38373 C10_N_btm.n2513 C10_N_btm.n2512 4.60698
R38374 C10_N_btm.n2509 C10_N_btm.n2508 4.60698
R38375 C10_N_btm.n2510 C10_N_btm.n2509 4.60698
R38376 C10_N_btm.n2506 C10_N_btm.n2505 4.60698
R38377 C10_N_btm.n2507 C10_N_btm.n2506 4.60698
R38378 C10_N_btm.n2503 C10_N_btm.n2502 4.60698
R38379 C10_N_btm.n2504 C10_N_btm.n2503 4.60698
R38380 C10_N_btm.n2500 C10_N_btm.n2499 4.60698
R38381 C10_N_btm.n2501 C10_N_btm.n2500 4.60698
R38382 C10_N_btm.n2497 C10_N_btm.n2496 4.60698
R38383 C10_N_btm.n2498 C10_N_btm.n2497 4.60698
R38384 C10_N_btm.n2494 C10_N_btm.n2493 4.60698
R38385 C10_N_btm.n2495 C10_N_btm.n2494 4.60698
R38386 C10_N_btm.n2491 C10_N_btm.n2490 4.60698
R38387 C10_N_btm.n2492 C10_N_btm.n2491 4.60698
R38388 C10_N_btm.n2488 C10_N_btm.n2487 4.60698
R38389 C10_N_btm.n2489 C10_N_btm.n2488 4.60698
R38390 C10_N_btm.n2485 C10_N_btm.n2484 4.60698
R38391 C10_N_btm.n2486 C10_N_btm.n2485 4.60698
R38392 C10_N_btm.n2482 C10_N_btm.n2481 4.60698
R38393 C10_N_btm.n2483 C10_N_btm.n2482 4.60698
R38394 C10_N_btm.n2479 C10_N_btm.n2478 4.60698
R38395 C10_N_btm.n2480 C10_N_btm.n2479 4.60698
R38396 C10_N_btm.n2476 C10_N_btm.n2475 4.60698
R38397 C10_N_btm.n2477 C10_N_btm.n2476 4.60698
R38398 C10_N_btm.n2473 C10_N_btm.n2472 4.60698
R38399 C10_N_btm.n2474 C10_N_btm.n2473 4.60698
R38400 C10_N_btm.n2470 C10_N_btm.n2469 4.60698
R38401 C10_N_btm.n2471 C10_N_btm.n2470 4.60698
R38402 C10_N_btm.n2467 C10_N_btm.n2466 4.60698
R38403 C10_N_btm.n2468 C10_N_btm.n2467 4.60698
R38404 C10_N_btm.n2464 C10_N_btm.n2463 4.60698
R38405 C10_N_btm.n2465 C10_N_btm.n2464 4.60698
R38406 C10_N_btm.n2461 C10_N_btm.n2460 4.60698
R38407 C10_N_btm.n2462 C10_N_btm.n2461 4.60698
R38408 C10_N_btm.n2458 C10_N_btm.n2457 4.60698
R38409 C10_N_btm.n2459 C10_N_btm.n2458 4.60698
R38410 C10_N_btm.n2455 C10_N_btm.n2454 4.60698
R38411 C10_N_btm.n2456 C10_N_btm.n2455 4.60698
R38412 C10_N_btm.n2452 C10_N_btm.n2451 4.60698
R38413 C10_N_btm.n2453 C10_N_btm.n2452 4.60698
R38414 C10_N_btm.n2449 C10_N_btm.n2448 4.60698
R38415 C10_N_btm.n2450 C10_N_btm.n2449 4.60698
R38416 C10_N_btm.n2446 C10_N_btm.n2445 4.60698
R38417 C10_N_btm.n2447 C10_N_btm.n2446 4.60698
R38418 C10_N_btm.n2443 C10_N_btm.n2442 4.60698
R38419 C10_N_btm.n2444 C10_N_btm.n2443 4.60698
R38420 C10_N_btm.n2440 C10_N_btm.n2439 4.60698
R38421 C10_N_btm.n2441 C10_N_btm.n2440 4.60698
R38422 C10_N_btm.n2437 C10_N_btm.n2436 4.60698
R38423 C10_N_btm.n2438 C10_N_btm.n2437 4.60698
R38424 C10_N_btm.n2434 C10_N_btm.n2433 4.60698
R38425 C10_N_btm.n2435 C10_N_btm.n2434 4.60698
R38426 C10_N_btm.n2431 C10_N_btm.n2430 4.60698
R38427 C10_N_btm.n2432 C10_N_btm.n2431 4.60698
R38428 C10_N_btm.n2428 C10_N_btm.n2427 4.60698
R38429 C10_N_btm.n2429 C10_N_btm.n2428 4.60698
R38430 C10_N_btm.n2425 C10_N_btm.n2424 4.60698
R38431 C10_N_btm.n2426 C10_N_btm.n2425 4.60698
R38432 C10_N_btm.n2422 C10_N_btm.n2421 4.60698
R38433 C10_N_btm.n2423 C10_N_btm.n2422 4.60698
R38434 C10_N_btm.n2419 C10_N_btm.n2418 4.60698
R38435 C10_N_btm.n2420 C10_N_btm.n2419 4.60698
R38436 C10_N_btm.n2416 C10_N_btm.n2415 4.60698
R38437 C10_N_btm.n2417 C10_N_btm.n2416 4.60698
R38438 C10_N_btm.n2413 C10_N_btm.n2412 4.60698
R38439 C10_N_btm.n2414 C10_N_btm.n2413 4.60698
R38440 C10_N_btm.n2410 C10_N_btm.n2409 4.60698
R38441 C10_N_btm.n2411 C10_N_btm.n2410 4.60698
R38442 C10_N_btm.n2407 C10_N_btm.n2406 4.60698
R38443 C10_N_btm.n2408 C10_N_btm.n2407 4.60698
R38444 C10_N_btm.n2404 C10_N_btm.n2403 4.60698
R38445 C10_N_btm.n2405 C10_N_btm.n2404 4.60698
R38446 C10_N_btm.n2401 C10_N_btm.n2400 4.60698
R38447 C10_N_btm.n2402 C10_N_btm.n2401 4.60698
R38448 C10_N_btm.n2398 C10_N_btm.n2397 4.60698
R38449 C10_N_btm.n2399 C10_N_btm.n2398 4.60698
R38450 C10_N_btm.n2395 C10_N_btm.n2394 4.60698
R38451 C10_N_btm.n2396 C10_N_btm.n2395 4.60698
R38452 C10_N_btm.n2392 C10_N_btm.n2391 4.60698
R38453 C10_N_btm.n2393 C10_N_btm.n2392 4.60698
R38454 C10_N_btm.n2389 C10_N_btm.n2388 4.60698
R38455 C10_N_btm.n2390 C10_N_btm.n2389 4.60698
R38456 C10_N_btm.n2386 C10_N_btm.n2385 4.60698
R38457 C10_N_btm.n2387 C10_N_btm.n2386 4.60698
R38458 C10_N_btm.n2383 C10_N_btm.n2382 4.60698
R38459 C10_N_btm.n2384 C10_N_btm.n2383 4.60698
R38460 C10_N_btm.n2380 C10_N_btm.n2379 4.60698
R38461 C10_N_btm.n2381 C10_N_btm.n2380 4.60698
R38462 C10_N_btm.n2377 C10_N_btm.n2376 4.60698
R38463 C10_N_btm.n2378 C10_N_btm.n2377 4.60698
R38464 C10_N_btm.n2374 C10_N_btm.n2373 4.60698
R38465 C10_N_btm.n2375 C10_N_btm.n2374 4.60698
R38466 C10_N_btm.n2371 C10_N_btm.n2370 4.60698
R38467 C10_N_btm.n2372 C10_N_btm.n2371 4.60698
R38468 C10_N_btm.n2368 C10_N_btm.n2367 4.60698
R38469 C10_N_btm.n2369 C10_N_btm.n2368 4.60698
R38470 C10_N_btm.n2365 C10_N_btm.n2364 4.60698
R38471 C10_N_btm.n2366 C10_N_btm.n2365 4.60698
R38472 C10_N_btm.n2362 C10_N_btm.n2361 4.60698
R38473 C10_N_btm.n2363 C10_N_btm.n2362 4.60698
R38474 C10_N_btm.n2359 C10_N_btm.n2358 4.60698
R38475 C10_N_btm.n2360 C10_N_btm.n2359 4.60698
R38476 C10_N_btm.n2356 C10_N_btm.n2355 4.60698
R38477 C10_N_btm.n2357 C10_N_btm.n2356 4.60698
R38478 C10_N_btm.n2353 C10_N_btm.n2352 4.60698
R38479 C10_N_btm.n2354 C10_N_btm.n2353 4.60698
R38480 C10_N_btm.n2350 C10_N_btm.n2349 4.60698
R38481 C10_N_btm.n2351 C10_N_btm.n2350 4.60698
R38482 C10_N_btm.n2347 C10_N_btm.n2346 4.60698
R38483 C10_N_btm.n2348 C10_N_btm.n2347 4.60698
R38484 C10_N_btm.n2344 C10_N_btm.n2343 4.60698
R38485 C10_N_btm.n2345 C10_N_btm.n2344 4.60698
R38486 C10_N_btm.n2341 C10_N_btm.n2340 4.60698
R38487 C10_N_btm.n2342 C10_N_btm.n2341 4.60698
R38488 C10_N_btm.n1594 C10_N_btm.n1593 4.60698
R38489 C10_N_btm.n1595 C10_N_btm.n1594 4.60698
R38490 C10_N_btm.n1591 C10_N_btm.n1590 4.60698
R38491 C10_N_btm.n1592 C10_N_btm.n1591 4.60698
R38492 C10_N_btm.n1588 C10_N_btm.n1587 4.60698
R38493 C10_N_btm.n1589 C10_N_btm.n1588 4.60698
R38494 C10_N_btm.n1585 C10_N_btm.n1584 4.60698
R38495 C10_N_btm.n1586 C10_N_btm.n1585 4.60698
R38496 C10_N_btm.n1582 C10_N_btm.n1581 4.60698
R38497 C10_N_btm.n1583 C10_N_btm.n1582 4.60698
R38498 C10_N_btm.n1579 C10_N_btm.n1578 4.60698
R38499 C10_N_btm.n1580 C10_N_btm.n1579 4.60698
R38500 C10_N_btm.n1576 C10_N_btm.n1575 4.60698
R38501 C10_N_btm.n1577 C10_N_btm.n1576 4.60698
R38502 C10_N_btm.n1573 C10_N_btm.n1572 4.60698
R38503 C10_N_btm.n1574 C10_N_btm.n1573 4.60698
R38504 C10_N_btm.n1570 C10_N_btm.n1569 4.60698
R38505 C10_N_btm.n1571 C10_N_btm.n1570 4.60698
R38506 C10_N_btm.n1567 C10_N_btm.n1566 4.60698
R38507 C10_N_btm.n1568 C10_N_btm.n1567 4.60698
R38508 C10_N_btm.n1513 C10_N_btm.n1512 4.60698
R38509 C10_N_btm.n1512 C10_N_btm.n1511 4.60698
R38510 C10_N_btm.n1510 C10_N_btm.n1509 4.60698
R38511 C10_N_btm.n1509 C10_N_btm.n1508 4.60698
R38512 C10_N_btm.n1507 C10_N_btm.n1506 4.60698
R38513 C10_N_btm.n1506 C10_N_btm.n1505 4.60698
R38514 C10_N_btm.n1504 C10_N_btm.n1503 4.60698
R38515 C10_N_btm.n1503 C10_N_btm.n1502 4.60698
R38516 C10_N_btm.n1501 C10_N_btm.n1500 4.60698
R38517 C10_N_btm.n1500 C10_N_btm.n1499 4.60698
R38518 C10_N_btm.n1498 C10_N_btm.n1497 4.60698
R38519 C10_N_btm.n1497 C10_N_btm.n1496 4.60698
R38520 C10_N_btm.n1495 C10_N_btm.n1494 4.60698
R38521 C10_N_btm.n1494 C10_N_btm.n1493 4.60698
R38522 C10_N_btm.n1492 C10_N_btm.n1491 4.60698
R38523 C10_N_btm.n1491 C10_N_btm.n1490 4.60698
R38524 C10_N_btm.n1489 C10_N_btm.n1488 4.60698
R38525 C10_N_btm.n1488 C10_N_btm.n1487 4.60698
R38526 C10_N_btm.n1483 C10_N_btm.n1482 4.60698
R38527 C10_N_btm.n1482 C10_N_btm.n567 4.60698
R38528 C10_N_btm.n1480 C10_N_btm.n1479 4.60698
R38529 C10_N_btm.n1481 C10_N_btm.n1480 4.60698
R38530 C10_N_btm.n1477 C10_N_btm.n1476 4.60698
R38531 C10_N_btm.n1478 C10_N_btm.n1477 4.60698
R38532 C10_N_btm.n1474 C10_N_btm.n1473 4.60698
R38533 C10_N_btm.n1475 C10_N_btm.n1474 4.60698
R38534 C10_N_btm.n1471 C10_N_btm.n1470 4.60698
R38535 C10_N_btm.n1472 C10_N_btm.n1471 4.60698
R38536 C10_N_btm.n1468 C10_N_btm.n1467 4.60698
R38537 C10_N_btm.n1469 C10_N_btm.n1468 4.60698
R38538 C10_N_btm.n1465 C10_N_btm.n1464 4.60698
R38539 C10_N_btm.n1466 C10_N_btm.n1465 4.60698
R38540 C10_N_btm.n1462 C10_N_btm.n1461 4.60698
R38541 C10_N_btm.n1463 C10_N_btm.n1462 4.60698
R38542 C10_N_btm.n1459 C10_N_btm.n1458 4.60698
R38543 C10_N_btm.n1460 C10_N_btm.n1459 4.60698
R38544 C10_N_btm.n1454 C10_N_btm.n1453 4.60698
R38545 C10_N_btm.n1453 C10_N_btm.n576 4.60698
R38546 C10_N_btm.n1395 C10_N_btm.n1394 4.60698
R38547 C10_N_btm.n1396 C10_N_btm.n1395 4.60698
R38548 C10_N_btm.n1398 C10_N_btm.n1397 4.60698
R38549 C10_N_btm.n1399 C10_N_btm.n1398 4.60698
R38550 C10_N_btm.n1401 C10_N_btm.n1400 4.60698
R38551 C10_N_btm.n1402 C10_N_btm.n1401 4.60698
R38552 C10_N_btm.n1404 C10_N_btm.n1403 4.60698
R38553 C10_N_btm.n1405 C10_N_btm.n1404 4.60698
R38554 C10_N_btm.n1407 C10_N_btm.n1406 4.60698
R38555 C10_N_btm.n1408 C10_N_btm.n1407 4.60698
R38556 C10_N_btm.n1410 C10_N_btm.n1409 4.60698
R38557 C10_N_btm.n1411 C10_N_btm.n1410 4.60698
R38558 C10_N_btm.n1413 C10_N_btm.n1412 4.60698
R38559 C10_N_btm.n1414 C10_N_btm.n1413 4.60698
R38560 C10_N_btm.n1416 C10_N_btm.n1415 4.60698
R38561 C10_N_btm.n1417 C10_N_btm.n1416 4.60698
R38562 C10_N_btm.n1424 C10_N_btm.n1423 4.60698
R38563 C10_N_btm.n1423 C10_N_btm.n1422 4.60698
R38564 C10_N_btm.n1427 C10_N_btm.n1426 4.60698
R38565 C10_N_btm.n1426 C10_N_btm.n1425 4.60698
R38566 C10_N_btm.n1430 C10_N_btm.n1429 4.60698
R38567 C10_N_btm.n1429 C10_N_btm.n1428 4.60698
R38568 C10_N_btm.n1433 C10_N_btm.n1432 4.60698
R38569 C10_N_btm.n1432 C10_N_btm.n1431 4.60698
R38570 C10_N_btm.n1436 C10_N_btm.n1435 4.60698
R38571 C10_N_btm.n1435 C10_N_btm.n1434 4.60698
R38572 C10_N_btm.n1439 C10_N_btm.n1438 4.60698
R38573 C10_N_btm.n1438 C10_N_btm.n1437 4.60698
R38574 C10_N_btm.n1442 C10_N_btm.n1441 4.60698
R38575 C10_N_btm.n1441 C10_N_btm.n1440 4.60698
R38576 C10_N_btm.n1445 C10_N_btm.n1444 4.60698
R38577 C10_N_btm.n1444 C10_N_btm.n1443 4.60698
R38578 C10_N_btm.n1448 C10_N_btm.n1447 4.60698
R38579 C10_N_btm.n1447 C10_N_btm.n1446 4.60698
R38580 C10_N_btm.n1357 C10_N_btm.n1356 4.60698
R38581 C10_N_btm.n1358 C10_N_btm.n1357 4.60698
R38582 C10_N_btm.n1360 C10_N_btm.n1359 4.60698
R38583 C10_N_btm.n1361 C10_N_btm.n1360 4.60698
R38584 C10_N_btm.n1363 C10_N_btm.n1362 4.60698
R38585 C10_N_btm.n1364 C10_N_btm.n1363 4.60698
R38586 C10_N_btm.n1366 C10_N_btm.n1365 4.60698
R38587 C10_N_btm.n1367 C10_N_btm.n1366 4.60698
R38588 C10_N_btm.n1369 C10_N_btm.n1368 4.60698
R38589 C10_N_btm.n1370 C10_N_btm.n1369 4.60698
R38590 C10_N_btm.n1372 C10_N_btm.n1371 4.60698
R38591 C10_N_btm.n1373 C10_N_btm.n1372 4.60698
R38592 C10_N_btm.n1375 C10_N_btm.n1374 4.60698
R38593 C10_N_btm.n1376 C10_N_btm.n1375 4.60698
R38594 C10_N_btm.n1378 C10_N_btm.n1377 4.60698
R38595 C10_N_btm.n1379 C10_N_btm.n1378 4.60698
R38596 C10_N_btm.n1381 C10_N_btm.n1380 4.60698
R38597 C10_N_btm.n1382 C10_N_btm.n1381 4.60698
R38598 C10_N_btm.n636 C10_N_btm.n635 4.60698
R38599 C10_N_btm.n635 C10_N_btm.n606 4.60698
R38600 C10_N_btm.n633 C10_N_btm.n632 4.60698
R38601 C10_N_btm.n634 C10_N_btm.n633 4.60698
R38602 C10_N_btm.n630 C10_N_btm.n629 4.60698
R38603 C10_N_btm.n631 C10_N_btm.n630 4.60698
R38604 C10_N_btm.n627 C10_N_btm.n626 4.60698
R38605 C10_N_btm.n628 C10_N_btm.n627 4.60698
R38606 C10_N_btm.n624 C10_N_btm.n623 4.60698
R38607 C10_N_btm.n625 C10_N_btm.n624 4.60698
R38608 C10_N_btm.n621 C10_N_btm.n620 4.60698
R38609 C10_N_btm.n622 C10_N_btm.n621 4.60698
R38610 C10_N_btm.n618 C10_N_btm.n617 4.60698
R38611 C10_N_btm.n619 C10_N_btm.n618 4.60698
R38612 C10_N_btm.n615 C10_N_btm.n614 4.60698
R38613 C10_N_btm.n616 C10_N_btm.n615 4.60698
R38614 C10_N_btm.n1352 C10_N_btm.n1351 4.60698
R38615 C10_N_btm.n1351 C10_N_btm.n596 4.60698
R38616 C10_N_btm.n1346 C10_N_btm.n1345 4.60698
R38617 C10_N_btm.n1345 C10_N_btm.n1344 4.60698
R38618 C10_N_btm.n1343 C10_N_btm.n1342 4.60698
R38619 C10_N_btm.n1342 C10_N_btm.n1341 4.60698
R38620 C10_N_btm.n1340 C10_N_btm.n1339 4.60698
R38621 C10_N_btm.n1339 C10_N_btm.n1338 4.60698
R38622 C10_N_btm.n1337 C10_N_btm.n1336 4.60698
R38623 C10_N_btm.n1336 C10_N_btm.n1335 4.60698
R38624 C10_N_btm.n1334 C10_N_btm.n1333 4.60698
R38625 C10_N_btm.n1333 C10_N_btm.n1332 4.60698
R38626 C10_N_btm.n1331 C10_N_btm.n1330 4.60698
R38627 C10_N_btm.n1330 C10_N_btm.n1329 4.60698
R38628 C10_N_btm.n1328 C10_N_btm.n1327 4.60698
R38629 C10_N_btm.n1327 C10_N_btm.n1326 4.60698
R38630 C10_N_btm.n1325 C10_N_btm.n1324 4.60698
R38631 C10_N_btm.n1324 C10_N_btm.n1323 4.60698
R38632 C10_N_btm.n1322 C10_N_btm.n1321 4.60698
R38633 C10_N_btm.n1321 C10_N_btm.n1320 4.60698
R38634 C10_N_btm.n1314 C10_N_btm.n1313 4.60698
R38635 C10_N_btm.n1315 C10_N_btm.n1314 4.60698
R38636 C10_N_btm.n1311 C10_N_btm.n1310 4.60698
R38637 C10_N_btm.n1312 C10_N_btm.n1311 4.60698
R38638 C10_N_btm.n1308 C10_N_btm.n1307 4.60698
R38639 C10_N_btm.n1309 C10_N_btm.n1308 4.60698
R38640 C10_N_btm.n1305 C10_N_btm.n1304 4.60698
R38641 C10_N_btm.n1306 C10_N_btm.n1305 4.60698
R38642 C10_N_btm.n1302 C10_N_btm.n1301 4.60698
R38643 C10_N_btm.n1303 C10_N_btm.n1302 4.60698
R38644 C10_N_btm.n1299 C10_N_btm.n1298 4.60698
R38645 C10_N_btm.n1300 C10_N_btm.n1299 4.60698
R38646 C10_N_btm.n1296 C10_N_btm.n1295 4.60698
R38647 C10_N_btm.n1297 C10_N_btm.n1296 4.60698
R38648 C10_N_btm.n1293 C10_N_btm.n1292 4.60698
R38649 C10_N_btm.n1294 C10_N_btm.n1293 4.60698
R38650 C10_N_btm.n1290 C10_N_btm.n1289 4.60698
R38651 C10_N_btm.n1291 C10_N_btm.n1290 4.60698
R38652 C10_N_btm.n1285 C10_N_btm.n1284 4.60698
R38653 C10_N_btm.n1284 C10_N_btm.n649 4.60698
R38654 C10_N_btm.n668 C10_N_btm.n667 4.60698
R38655 C10_N_btm.n669 C10_N_btm.n668 4.60698
R38656 C10_N_btm.n671 C10_N_btm.n670 4.60698
R38657 C10_N_btm.n672 C10_N_btm.n671 4.60698
R38658 C10_N_btm.n674 C10_N_btm.n673 4.60698
R38659 C10_N_btm.n675 C10_N_btm.n674 4.60698
R38660 C10_N_btm.n677 C10_N_btm.n676 4.60698
R38661 C10_N_btm.n678 C10_N_btm.n677 4.60698
R38662 C10_N_btm.n680 C10_N_btm.n679 4.60698
R38663 C10_N_btm.n681 C10_N_btm.n680 4.60698
R38664 C10_N_btm.n683 C10_N_btm.n682 4.60698
R38665 C10_N_btm.n684 C10_N_btm.n683 4.60698
R38666 C10_N_btm.n686 C10_N_btm.n685 4.60698
R38667 C10_N_btm.n687 C10_N_btm.n686 4.60698
R38668 C10_N_btm.n689 C10_N_btm.n688 4.60698
R38669 C10_N_btm.n688 C10_N_btm.n659 4.60698
R38670 C10_N_btm.n1255 C10_N_btm.n1254 4.60698
R38671 C10_N_btm.n1254 C10_N_btm.n1253 4.60698
R38672 C10_N_btm.n1258 C10_N_btm.n1257 4.60698
R38673 C10_N_btm.n1257 C10_N_btm.n1256 4.60698
R38674 C10_N_btm.n1261 C10_N_btm.n1260 4.60698
R38675 C10_N_btm.n1260 C10_N_btm.n1259 4.60698
R38676 C10_N_btm.n1264 C10_N_btm.n1263 4.60698
R38677 C10_N_btm.n1263 C10_N_btm.n1262 4.60698
R38678 C10_N_btm.n1267 C10_N_btm.n1266 4.60698
R38679 C10_N_btm.n1266 C10_N_btm.n1265 4.60698
R38680 C10_N_btm.n1270 C10_N_btm.n1269 4.60698
R38681 C10_N_btm.n1269 C10_N_btm.n1268 4.60698
R38682 C10_N_btm.n1273 C10_N_btm.n1272 4.60698
R38683 C10_N_btm.n1272 C10_N_btm.n1271 4.60698
R38684 C10_N_btm.n1276 C10_N_btm.n1275 4.60698
R38685 C10_N_btm.n1275 C10_N_btm.n1274 4.60698
R38686 C10_N_btm.n1279 C10_N_btm.n1278 4.60698
R38687 C10_N_btm.n1278 C10_N_btm.n1277 4.60698
R38688 C10_N_btm.n1223 C10_N_btm.n1222 4.60698
R38689 C10_N_btm.n1224 C10_N_btm.n1223 4.60698
R38690 C10_N_btm.n1226 C10_N_btm.n1225 4.60698
R38691 C10_N_btm.n1227 C10_N_btm.n1226 4.60698
R38692 C10_N_btm.n1229 C10_N_btm.n1228 4.60698
R38693 C10_N_btm.n1230 C10_N_btm.n1229 4.60698
R38694 C10_N_btm.n1232 C10_N_btm.n1231 4.60698
R38695 C10_N_btm.n1233 C10_N_btm.n1232 4.60698
R38696 C10_N_btm.n1235 C10_N_btm.n1234 4.60698
R38697 C10_N_btm.n1236 C10_N_btm.n1235 4.60698
R38698 C10_N_btm.n1238 C10_N_btm.n1237 4.60698
R38699 C10_N_btm.n1239 C10_N_btm.n1238 4.60698
R38700 C10_N_btm.n1241 C10_N_btm.n1240 4.60698
R38701 C10_N_btm.n1242 C10_N_btm.n1241 4.60698
R38702 C10_N_btm.n1244 C10_N_btm.n1243 4.60698
R38703 C10_N_btm.n1245 C10_N_btm.n1244 4.60698
R38704 C10_N_btm.n1247 C10_N_btm.n1246 4.60698
R38705 C10_N_btm.n1248 C10_N_btm.n1247 4.60698
R38706 C10_N_btm.n742 C10_N_btm.n741 4.60698
R38707 C10_N_btm.n741 C10_N_btm.n712 4.60698
R38708 C10_N_btm.n739 C10_N_btm.n738 4.60698
R38709 C10_N_btm.n740 C10_N_btm.n739 4.60698
R38710 C10_N_btm.n736 C10_N_btm.n735 4.60698
R38711 C10_N_btm.n737 C10_N_btm.n736 4.60698
R38712 C10_N_btm.n733 C10_N_btm.n732 4.60698
R38713 C10_N_btm.n734 C10_N_btm.n733 4.60698
R38714 C10_N_btm.n730 C10_N_btm.n729 4.60698
R38715 C10_N_btm.n731 C10_N_btm.n730 4.60698
R38716 C10_N_btm.n727 C10_N_btm.n726 4.60698
R38717 C10_N_btm.n728 C10_N_btm.n727 4.60698
R38718 C10_N_btm.n724 C10_N_btm.n723 4.60698
R38719 C10_N_btm.n725 C10_N_btm.n724 4.60698
R38720 C10_N_btm.n721 C10_N_btm.n720 4.60698
R38721 C10_N_btm.n722 C10_N_btm.n721 4.60698
R38722 C10_N_btm.n1218 C10_N_btm.n1217 4.60698
R38723 C10_N_btm.n1217 C10_N_btm.n702 4.60698
R38724 C10_N_btm.n1212 C10_N_btm.n1211 4.60698
R38725 C10_N_btm.n1211 C10_N_btm.n1210 4.60698
R38726 C10_N_btm.n1209 C10_N_btm.n1208 4.60698
R38727 C10_N_btm.n1208 C10_N_btm.n1207 4.60698
R38728 C10_N_btm.n1206 C10_N_btm.n1205 4.60698
R38729 C10_N_btm.n1205 C10_N_btm.n1204 4.60698
R38730 C10_N_btm.n1203 C10_N_btm.n1202 4.60698
R38731 C10_N_btm.n1202 C10_N_btm.n1201 4.60698
R38732 C10_N_btm.n1200 C10_N_btm.n1199 4.60698
R38733 C10_N_btm.n1199 C10_N_btm.n1198 4.60698
R38734 C10_N_btm.n1197 C10_N_btm.n1196 4.60698
R38735 C10_N_btm.n1196 C10_N_btm.n1195 4.60698
R38736 C10_N_btm.n1194 C10_N_btm.n1193 4.60698
R38737 C10_N_btm.n1193 C10_N_btm.n1192 4.60698
R38738 C10_N_btm.n1191 C10_N_btm.n1190 4.60698
R38739 C10_N_btm.n1190 C10_N_btm.n1189 4.60698
R38740 C10_N_btm.n1188 C10_N_btm.n1187 4.60698
R38741 C10_N_btm.n1187 C10_N_btm.n1186 4.60698
R38742 C10_N_btm.n1180 C10_N_btm.n1179 4.60698
R38743 C10_N_btm.n1181 C10_N_btm.n1180 4.60698
R38744 C10_N_btm.n1177 C10_N_btm.n1176 4.60698
R38745 C10_N_btm.n1178 C10_N_btm.n1177 4.60698
R38746 C10_N_btm.n1174 C10_N_btm.n1173 4.60698
R38747 C10_N_btm.n1175 C10_N_btm.n1174 4.60698
R38748 C10_N_btm.n1171 C10_N_btm.n1170 4.60698
R38749 C10_N_btm.n1172 C10_N_btm.n1171 4.60698
R38750 C10_N_btm.n1168 C10_N_btm.n1167 4.60698
R38751 C10_N_btm.n1169 C10_N_btm.n1168 4.60698
R38752 C10_N_btm.n1165 C10_N_btm.n1164 4.60698
R38753 C10_N_btm.n1166 C10_N_btm.n1165 4.60698
R38754 C10_N_btm.n1162 C10_N_btm.n1161 4.60698
R38755 C10_N_btm.n1163 C10_N_btm.n1162 4.60698
R38756 C10_N_btm.n1159 C10_N_btm.n1158 4.60698
R38757 C10_N_btm.n1160 C10_N_btm.n1159 4.60698
R38758 C10_N_btm.n1156 C10_N_btm.n1155 4.60698
R38759 C10_N_btm.n1157 C10_N_btm.n1156 4.60698
R38760 C10_N_btm.n1151 C10_N_btm.n1150 4.60698
R38761 C10_N_btm.n1150 C10_N_btm.n755 4.60698
R38762 C10_N_btm.n774 C10_N_btm.n773 4.60698
R38763 C10_N_btm.n775 C10_N_btm.n774 4.60698
R38764 C10_N_btm.n777 C10_N_btm.n776 4.60698
R38765 C10_N_btm.n778 C10_N_btm.n777 4.60698
R38766 C10_N_btm.n780 C10_N_btm.n779 4.60698
R38767 C10_N_btm.n781 C10_N_btm.n780 4.60698
R38768 C10_N_btm.n783 C10_N_btm.n782 4.60698
R38769 C10_N_btm.n784 C10_N_btm.n783 4.60698
R38770 C10_N_btm.n786 C10_N_btm.n785 4.60698
R38771 C10_N_btm.n787 C10_N_btm.n786 4.60698
R38772 C10_N_btm.n789 C10_N_btm.n788 4.60698
R38773 C10_N_btm.n790 C10_N_btm.n789 4.60698
R38774 C10_N_btm.n792 C10_N_btm.n791 4.60698
R38775 C10_N_btm.n793 C10_N_btm.n792 4.60698
R38776 C10_N_btm.n795 C10_N_btm.n794 4.60698
R38777 C10_N_btm.n794 C10_N_btm.n765 4.60698
R38778 C10_N_btm.n1121 C10_N_btm.n1120 4.60698
R38779 C10_N_btm.n1120 C10_N_btm.n1119 4.60698
R38780 C10_N_btm.n1124 C10_N_btm.n1123 4.60698
R38781 C10_N_btm.n1123 C10_N_btm.n1122 4.60698
R38782 C10_N_btm.n1127 C10_N_btm.n1126 4.60698
R38783 C10_N_btm.n1126 C10_N_btm.n1125 4.60698
R38784 C10_N_btm.n1130 C10_N_btm.n1129 4.60698
R38785 C10_N_btm.n1129 C10_N_btm.n1128 4.60698
R38786 C10_N_btm.n1133 C10_N_btm.n1132 4.60698
R38787 C10_N_btm.n1132 C10_N_btm.n1131 4.60698
R38788 C10_N_btm.n1136 C10_N_btm.n1135 4.60698
R38789 C10_N_btm.n1135 C10_N_btm.n1134 4.60698
R38790 C10_N_btm.n1139 C10_N_btm.n1138 4.60698
R38791 C10_N_btm.n1138 C10_N_btm.n1137 4.60698
R38792 C10_N_btm.n1142 C10_N_btm.n1141 4.60698
R38793 C10_N_btm.n1141 C10_N_btm.n1140 4.60698
R38794 C10_N_btm.n1145 C10_N_btm.n1144 4.60698
R38795 C10_N_btm.n1144 C10_N_btm.n1143 4.60698
R38796 C10_N_btm.n1089 C10_N_btm.n1088 4.60698
R38797 C10_N_btm.n1090 C10_N_btm.n1089 4.60698
R38798 C10_N_btm.n1092 C10_N_btm.n1091 4.60698
R38799 C10_N_btm.n1093 C10_N_btm.n1092 4.60698
R38800 C10_N_btm.n1095 C10_N_btm.n1094 4.60698
R38801 C10_N_btm.n1096 C10_N_btm.n1095 4.60698
R38802 C10_N_btm.n1098 C10_N_btm.n1097 4.60698
R38803 C10_N_btm.n1099 C10_N_btm.n1098 4.60698
R38804 C10_N_btm.n1101 C10_N_btm.n1100 4.60698
R38805 C10_N_btm.n1102 C10_N_btm.n1101 4.60698
R38806 C10_N_btm.n1104 C10_N_btm.n1103 4.60698
R38807 C10_N_btm.n1105 C10_N_btm.n1104 4.60698
R38808 C10_N_btm.n1107 C10_N_btm.n1106 4.60698
R38809 C10_N_btm.n1108 C10_N_btm.n1107 4.60698
R38810 C10_N_btm.n1110 C10_N_btm.n1109 4.60698
R38811 C10_N_btm.n1111 C10_N_btm.n1110 4.60698
R38812 C10_N_btm.n1113 C10_N_btm.n1112 4.60698
R38813 C10_N_btm.n1114 C10_N_btm.n1113 4.60698
R38814 C10_N_btm.n848 C10_N_btm.n847 4.60698
R38815 C10_N_btm.n847 C10_N_btm.n818 4.60698
R38816 C10_N_btm.n845 C10_N_btm.n844 4.60698
R38817 C10_N_btm.n846 C10_N_btm.n845 4.60698
R38818 C10_N_btm.n842 C10_N_btm.n841 4.60698
R38819 C10_N_btm.n843 C10_N_btm.n842 4.60698
R38820 C10_N_btm.n839 C10_N_btm.n838 4.60698
R38821 C10_N_btm.n840 C10_N_btm.n839 4.60698
R38822 C10_N_btm.n836 C10_N_btm.n835 4.60698
R38823 C10_N_btm.n837 C10_N_btm.n836 4.60698
R38824 C10_N_btm.n833 C10_N_btm.n832 4.60698
R38825 C10_N_btm.n834 C10_N_btm.n833 4.60698
R38826 C10_N_btm.n830 C10_N_btm.n829 4.60698
R38827 C10_N_btm.n831 C10_N_btm.n830 4.60698
R38828 C10_N_btm.n827 C10_N_btm.n826 4.60698
R38829 C10_N_btm.n828 C10_N_btm.n827 4.60698
R38830 C10_N_btm.n1084 C10_N_btm.n1083 4.60698
R38831 C10_N_btm.n1083 C10_N_btm.n808 4.60698
R38832 C10_N_btm.n1078 C10_N_btm.n1077 4.60698
R38833 C10_N_btm.n1077 C10_N_btm.n1076 4.60698
R38834 C10_N_btm.n1075 C10_N_btm.n1074 4.60698
R38835 C10_N_btm.n1074 C10_N_btm.n1073 4.60698
R38836 C10_N_btm.n1072 C10_N_btm.n1071 4.60698
R38837 C10_N_btm.n1071 C10_N_btm.n1070 4.60698
R38838 C10_N_btm.n1069 C10_N_btm.n1068 4.60698
R38839 C10_N_btm.n1068 C10_N_btm.n1067 4.60698
R38840 C10_N_btm.n1066 C10_N_btm.n1065 4.60698
R38841 C10_N_btm.n1065 C10_N_btm.n1064 4.60698
R38842 C10_N_btm.n1063 C10_N_btm.n1062 4.60698
R38843 C10_N_btm.n1062 C10_N_btm.n1061 4.60698
R38844 C10_N_btm.n1060 C10_N_btm.n1059 4.60698
R38845 C10_N_btm.n1059 C10_N_btm.n1058 4.60698
R38846 C10_N_btm.n1057 C10_N_btm.n1056 4.60698
R38847 C10_N_btm.n1056 C10_N_btm.n1055 4.60698
R38848 C10_N_btm.n1054 C10_N_btm.n1053 4.60698
R38849 C10_N_btm.n1053 C10_N_btm.n1052 4.60698
R38850 C10_N_btm.n1046 C10_N_btm.n1045 4.60698
R38851 C10_N_btm.n1047 C10_N_btm.n1046 4.60698
R38852 C10_N_btm.n1043 C10_N_btm.n1042 4.60698
R38853 C10_N_btm.n1044 C10_N_btm.n1043 4.60698
R38854 C10_N_btm.n1040 C10_N_btm.n1039 4.60698
R38855 C10_N_btm.n1041 C10_N_btm.n1040 4.60698
R38856 C10_N_btm.n1037 C10_N_btm.n1036 4.60698
R38857 C10_N_btm.n1038 C10_N_btm.n1037 4.60698
R38858 C10_N_btm.n1034 C10_N_btm.n1033 4.60698
R38859 C10_N_btm.n1035 C10_N_btm.n1034 4.60698
R38860 C10_N_btm.n1031 C10_N_btm.n1030 4.60698
R38861 C10_N_btm.n1032 C10_N_btm.n1031 4.60698
R38862 C10_N_btm.n1028 C10_N_btm.n1027 4.60698
R38863 C10_N_btm.n1029 C10_N_btm.n1028 4.60698
R38864 C10_N_btm.n1025 C10_N_btm.n1024 4.60698
R38865 C10_N_btm.n1026 C10_N_btm.n1025 4.60698
R38866 C10_N_btm.n1022 C10_N_btm.n1021 4.60698
R38867 C10_N_btm.n1023 C10_N_btm.n1022 4.60698
R38868 C10_N_btm.n1017 C10_N_btm.n1016 4.60698
R38869 C10_N_btm.n1016 C10_N_btm.n861 4.60698
R38870 C10_N_btm.n880 C10_N_btm.n879 4.60698
R38871 C10_N_btm.n881 C10_N_btm.n880 4.60698
R38872 C10_N_btm.n883 C10_N_btm.n882 4.60698
R38873 C10_N_btm.n884 C10_N_btm.n883 4.60698
R38874 C10_N_btm.n886 C10_N_btm.n885 4.60698
R38875 C10_N_btm.n887 C10_N_btm.n886 4.60698
R38876 C10_N_btm.n889 C10_N_btm.n888 4.60698
R38877 C10_N_btm.n890 C10_N_btm.n889 4.60698
R38878 C10_N_btm.n892 C10_N_btm.n891 4.60698
R38879 C10_N_btm.n893 C10_N_btm.n892 4.60698
R38880 C10_N_btm.n895 C10_N_btm.n894 4.60698
R38881 C10_N_btm.n896 C10_N_btm.n895 4.60698
R38882 C10_N_btm.n898 C10_N_btm.n897 4.60698
R38883 C10_N_btm.n899 C10_N_btm.n898 4.60698
R38884 C10_N_btm.n901 C10_N_btm.n900 4.60698
R38885 C10_N_btm.n900 C10_N_btm.n871 4.60698
R38886 C10_N_btm.n987 C10_N_btm.n986 4.60698
R38887 C10_N_btm.n986 C10_N_btm.n985 4.60698
R38888 C10_N_btm.n990 C10_N_btm.n989 4.60698
R38889 C10_N_btm.n989 C10_N_btm.n988 4.60698
R38890 C10_N_btm.n993 C10_N_btm.n992 4.60698
R38891 C10_N_btm.n992 C10_N_btm.n991 4.60698
R38892 C10_N_btm.n996 C10_N_btm.n995 4.60698
R38893 C10_N_btm.n995 C10_N_btm.n994 4.60698
R38894 C10_N_btm.n999 C10_N_btm.n998 4.60698
R38895 C10_N_btm.n998 C10_N_btm.n997 4.60698
R38896 C10_N_btm.n1002 C10_N_btm.n1001 4.60698
R38897 C10_N_btm.n1001 C10_N_btm.n1000 4.60698
R38898 C10_N_btm.n1005 C10_N_btm.n1004 4.60698
R38899 C10_N_btm.n1004 C10_N_btm.n1003 4.60698
R38900 C10_N_btm.n1008 C10_N_btm.n1007 4.60698
R38901 C10_N_btm.n1007 C10_N_btm.n1006 4.60698
R38902 C10_N_btm.n1011 C10_N_btm.n1010 4.60698
R38903 C10_N_btm.n1010 C10_N_btm.n1009 4.60698
R38904 C10_N_btm.n955 C10_N_btm.n954 4.60698
R38905 C10_N_btm.n956 C10_N_btm.n955 4.60698
R38906 C10_N_btm.n958 C10_N_btm.n957 4.60698
R38907 C10_N_btm.n959 C10_N_btm.n958 4.60698
R38908 C10_N_btm.n961 C10_N_btm.n960 4.60698
R38909 C10_N_btm.n962 C10_N_btm.n961 4.60698
R38910 C10_N_btm.n964 C10_N_btm.n963 4.60698
R38911 C10_N_btm.n965 C10_N_btm.n964 4.60698
R38912 C10_N_btm.n967 C10_N_btm.n966 4.60698
R38913 C10_N_btm.n968 C10_N_btm.n967 4.60698
R38914 C10_N_btm.n970 C10_N_btm.n969 4.60698
R38915 C10_N_btm.n971 C10_N_btm.n970 4.60698
R38916 C10_N_btm.n973 C10_N_btm.n972 4.60698
R38917 C10_N_btm.n974 C10_N_btm.n973 4.60698
R38918 C10_N_btm.n976 C10_N_btm.n975 4.60698
R38919 C10_N_btm.n977 C10_N_btm.n976 4.60698
R38920 C10_N_btm.n979 C10_N_btm.n978 4.60698
R38921 C10_N_btm.n980 C10_N_btm.n979 4.60698
R38922 C10_N_btm.n924 C10_N_btm.n923 4.60698
R38923 C10_N_btm.n923 C10_N_btm.n922 4.60698
R38924 C10_N_btm.n927 C10_N_btm.n926 4.60698
R38925 C10_N_btm.n926 C10_N_btm.n925 4.60698
R38926 C10_N_btm.n930 C10_N_btm.n929 4.60698
R38927 C10_N_btm.n929 C10_N_btm.n928 4.60698
R38928 C10_N_btm.n933 C10_N_btm.n932 4.60698
R38929 C10_N_btm.n932 C10_N_btm.n931 4.60698
R38930 C10_N_btm.n936 C10_N_btm.n935 4.60698
R38931 C10_N_btm.n935 C10_N_btm.n934 4.60698
R38932 C10_N_btm.n939 C10_N_btm.n938 4.60698
R38933 C10_N_btm.n938 C10_N_btm.n937 4.60698
R38934 C10_N_btm.n942 C10_N_btm.n941 4.60698
R38935 C10_N_btm.n941 C10_N_btm.n940 4.60698
R38936 C10_N_btm.n945 C10_N_btm.n944 4.60698
R38937 C10_N_btm.n944 C10_N_btm.n943 4.60698
R38938 C10_N_btm.n950 C10_N_btm.n949 4.60698
R38939 C10_N_btm.n949 C10_N_btm.n946 4.60698
R38940 C10_N_btm.n1564 C10_N_btm.n1563 4.60698
R38941 C10_N_btm.n1565 C10_N_btm.n1564 4.60698
R38942 C10_N_btm.n1561 C10_N_btm.n1560 4.60698
R38943 C10_N_btm.n1562 C10_N_btm.n1561 4.60698
R38944 C10_N_btm.n1558 C10_N_btm.n1557 4.60698
R38945 C10_N_btm.n1559 C10_N_btm.n1558 4.60698
R38946 C10_N_btm.n1555 C10_N_btm.n1554 4.60698
R38947 C10_N_btm.n1556 C10_N_btm.n1555 4.60698
R38948 C10_N_btm.n1552 C10_N_btm.n1551 4.60698
R38949 C10_N_btm.n1553 C10_N_btm.n1552 4.60698
R38950 C10_N_btm.n1549 C10_N_btm.n1548 4.60698
R38951 C10_N_btm.n1550 C10_N_btm.n1549 4.60698
R38952 C10_N_btm.n1546 C10_N_btm.n1545 4.60698
R38953 C10_N_btm.n1547 C10_N_btm.n1546 4.60698
R38954 C10_N_btm.n1543 C10_N_btm.n1542 4.60698
R38955 C10_N_btm.n1544 C10_N_btm.n1543 4.60698
R38956 C10_N_btm.n1540 C10_N_btm.n1539 4.60698
R38957 C10_N_btm.n1541 C10_N_btm.n1540 4.60698
R38958 C10_N_btm.n1537 C10_N_btm.n1536 4.60698
R38959 C10_N_btm.n1538 C10_N_btm.n1537 4.60698
R38960 C10_N_btm.n1534 C10_N_btm.n1533 4.60698
R38961 C10_N_btm.n1535 C10_N_btm.n1534 4.60698
R38962 C10_N_btm.n1531 C10_N_btm.n1530 4.60698
R38963 C10_N_btm.n1532 C10_N_btm.n1531 4.60698
R38964 C10_N_btm.n3897 C10_N_btm.t1075 4.03712
R38965 C10_N_btm.n3895 C10_N_btm.t513 3.98193
R38966 C10_N_btm.n3836 C10_N_btm.t1001 3.98193
R38967 C10_N_btm.n3735 C10_N_btm.t322 3.98193
R38968 C10_N_btm.n3768 C10_N_btm.t825 3.98193
R38969 C10_N_btm.n3771 C10_N_btm.t168 3.98193
R38970 C10_N_btm.n3733 C10_N_btm.t526 3.98193
R38971 C10_N_btm.n91 C10_N_btm.t634 3.98193
R38972 C10_N_btm.n3669 C10_N_btm.t364 3.98193
R38973 C10_N_btm.n3666 C10_N_btm.t876 3.98193
R38974 C10_N_btm.n144 C10_N_btm.t207 3.98193
R38975 C10_N_btm.n3602 C10_N_btm.t576 3.98193
R38976 C10_N_btm.n3599 C10_N_btm.t106 3.98193
R38977 C10_N_btm.n197 C10_N_btm.t410 3.98193
R38978 C10_N_btm.n3535 C10_N_btm.t927 3.98193
R38979 C10_N_btm.n3532 C10_N_btm.t256 3.98193
R38980 C10_N_btm.n250 C10_N_btm.t628 3.98193
R38981 C10_N_btm.n3468 C10_N_btm.t104 3.98193
R38982 C10_N_btm.n3465 C10_N_btm.t454 3.98193
R38983 C10_N_btm.n303 C10_N_btm.t972 3.98193
R38984 C10_N_btm.n3401 C10_N_btm.t293 3.98193
R38985 C10_N_btm.n3398 C10_N_btm.t681 3.98193
R38986 C10_N_btm.n356 C10_N_btm.t725 3.98193
R38987 C10_N_btm.n3334 C10_N_btm.t73 3.98193
R38988 C10_N_btm.n3331 C10_N_btm.t550 3.98193
R38989 C10_N_btm.n506 C10_N_btm.t127 3.98193
R38990 C10_N_btm.n3108 C10_N_btm.t1044 3.98193
R38991 C10_N_btm.n3105 C10_N_btm.t177 3.98193
R38992 C10_N_btm.n1723 C10_N_btm.t264 3.98193
R38993 C10_N_btm.n2723 C10_N_btm.t964 3.98193
R38994 C10_N_btm.n2720 C10_N_btm.t117 3.98193
R38995 C10_N_btm.n2093 C10_N_btm.t212 3.98193
R38996 C10_N_btm.n2526 C10_N_btm.t633 3.98193
R38997 C10_N_btm.n2339 C10_N_btm.t791 3.98193
R38998 C10_N_btm.n2528 C10_N_btm.t146 3.98193
R38999 C10_N_btm.n2533 C10_N_btm.t806 3.98193
R39000 C10_N_btm.n2910 C10_N_btm.t414 3.98193
R39001 C10_N_btm.n2913 C10_N_btm.t980 3.98193
R39002 C10_N_btm.n2918 C10_N_btm.t579 3.98193
R39003 C10_N_btm.n1596 C10_N_btm.t421 3.98193
R39004 C10_N_btm.n1486 C10_N_btm.t328 3.98193
R39005 C10_N_btm.n1385 C10_N_btm.t689 3.98193
R39006 C10_N_btm.n1418 C10_N_btm.t585 3.98193
R39007 C10_N_btm.n1421 C10_N_btm.t1046 3.98193
R39008 C10_N_btm.n1383 C10_N_btm.t423 3.98193
R39009 C10_N_btm.n605 C10_N_btm.t333 3.98193
R39010 C10_N_btm.n1319 C10_N_btm.t691 3.98193
R39011 C10_N_btm.n1316 C10_N_btm.t588 3.98193
R39012 C10_N_btm.n658 C10_N_btm.t959 3.98193
R39013 C10_N_btm.n1252 C10_N_btm.t863 3.98193
R39014 C10_N_btm.n1249 C10_N_btm.t763 3.98193
R39015 C10_N_btm.n711 C10_N_btm.t76 3.98193
R39016 C10_N_btm.n1185 C10_N_btm.t46 3.98193
R39017 C10_N_btm.n1182 C10_N_btm.t324 3.98193
R39018 C10_N_btm.n764 C10_N_btm.t514 3.98193
R39019 C10_N_btm.n1118 C10_N_btm.t151 3.98193
R39020 C10_N_btm.n1115 C10_N_btm.t597 3.98193
R39021 C10_N_btm.n817 C10_N_btm.t390 3.98193
R39022 C10_N_btm.n1051 C10_N_btm.t756 3.98193
R39023 C10_N_btm.n1048 C10_N_btm.t662 3.98193
R39024 C10_N_btm.n870 C10_N_btm.t556 3.98193
R39025 C10_N_btm.n984 C10_N_btm.t930 3.98193
R39026 C10_N_btm.n981 C10_N_btm.t831 3.98193
R39027 C10_N_btm.n921 C10_N_btm.t139 3.98193
R39028 C10_N_btm.n948 C10_N_btm.t1003 3.98193
R39029 C10_N_btm.n953 C10_N_btm.t636 3.98193
R39030 C10_N_btm.n1012 C10_N_btm.t728 3.98193
R39031 C10_N_btm.n1015 C10_N_btm.t372 3.98193
R39032 C10_N_btm.n1020 C10_N_btm.t463 3.98193
R39033 C10_N_btm.n1079 C10_N_btm.t555 3.98193
R39034 C10_N_btm.n1082 C10_N_btm.t227 3.98193
R39035 C10_N_btm.n1087 C10_N_btm.t303 3.98193
R39036 C10_N_btm.n1146 C10_N_btm.t1016 3.98193
R39037 C10_N_btm.n1149 C10_N_btm.t775 3.98193
R39038 C10_N_btm.n1154 C10_N_btm.t150 3.98193
R39039 C10_N_btm.n1213 C10_N_btm.t838 3.98193
R39040 C10_N_btm.n1216 C10_N_btm.t937 3.98193
R39041 C10_N_btm.n1221 C10_N_btm.t561 3.98193
R39042 C10_N_btm.n1280 C10_N_btm.t669 3.98193
R39043 C10_N_btm.n1283 C10_N_btm.t762 3.98193
R39044 C10_N_btm.n1288 C10_N_btm.t397 3.98193
R39045 C10_N_btm.n1347 C10_N_btm.t892 3.98193
R39046 C10_N_btm.n1350 C10_N_btm.t158 3.98193
R39047 C10_N_btm.n1355 C10_N_btm.t992 3.98193
R39048 C10_N_btm.n1449 C10_N_btm.t332 3.98193
R39049 C10_N_btm.n1452 C10_N_btm.t395 3.98193
R39050 C10_N_btm.n1457 C10_N_btm.t619 3.98193
R39051 C10_N_btm.n1514 C10_N_btm.t155 3.98193
R39052 C10_N_btm.n1529 C10_N_btm.t886 3.98193
R39053 C10_N_btm.n3295 C10_N_btm.t112 3.98193
R39054 C10_N_btm.n3298 C10_N_btm.t758 3.98193
R39055 C10_N_btm.n3303 C10_N_btm.t370 3.98193
R39056 C10_N_btm.n3362 C10_N_btm.t932 3.98193
R39057 C10_N_btm.n3365 C10_N_btm.t531 3.98193
R39058 C10_N_btm.n3370 C10_N_btm.t512 3.98193
R39059 C10_N_btm.n3429 C10_N_btm.t500 3.98193
R39060 C10_N_btm.n3432 C10_N_btm.t783 3.98193
R39061 C10_N_btm.n3437 C10_N_btm.t273 3.98193
R39062 C10_N_btm.n3496 C10_N_btm.t953 3.98193
R39063 C10_N_btm.n3499 C10_N_btm.t435 3.98193
R39064 C10_N_btm.n3504 C10_N_btm.t70 3.98193
R39065 C10_N_btm.n3563 C10_N_btm.t723 3.98193
R39066 C10_N_btm.n3566 C10_N_btm.t499 3.98193
R39067 C10_N_btm.n3571 C10_N_btm.t902 3.98193
R39068 C10_N_btm.n3630 C10_N_btm.t1053 3.98193
R39069 C10_N_btm.n3633 C10_N_btm.t477 3.98193
R39070 C10_N_btm.n3638 C10_N_btm.t684 3.98193
R39071 C10_N_btm.n3697 C10_N_btm.t187 3.98193
R39072 C10_N_btm.n3700 C10_N_btm.t857 3.98193
R39073 C10_N_btm.n3705 C10_N_btm.t346 3.98193
R39074 C10_N_btm.n3799 C10_N_btm.t222 3.98193
R39075 C10_N_btm.n3802 C10_N_btm.t632 3.98193
R39076 C10_N_btm.n3807 C10_N_btm.t145 3.98193
R39077 C10_N_btm.n3864 C10_N_btm.t805 3.98193
R39078 C10_N_btm.n3867 C10_N_btm.t298 3.98193
R39079 C10_N_btm.n13 C10_N_btm.t19 3.57113
R39080 C10_N_btm.n13 C10_N_btm.t27 3.57113
R39081 C10_N_btm.n11 C10_N_btm.t21 3.57113
R39082 C10_N_btm.n11 C10_N_btm.t25 3.57113
R39083 C10_N_btm.n9 C10_N_btm.t29 3.57113
R39084 C10_N_btm.n9 C10_N_btm.t33 3.57113
R39085 C10_N_btm.n7 C10_N_btm.t28 3.57113
R39086 C10_N_btm.n7 C10_N_btm.t32 3.57113
R39087 C10_N_btm.n5 C10_N_btm.t26 3.57113
R39088 C10_N_btm.n5 C10_N_btm.t18 3.57113
R39089 C10_N_btm.n3 C10_N_btm.t22 3.57113
R39090 C10_N_btm.n3 C10_N_btm.t20 3.57113
R39091 C10_N_btm.n1 C10_N_btm.t30 3.57113
R39092 C10_N_btm.n1 C10_N_btm.t24 3.57113
R39093 C10_N_btm.n0 C10_N_btm.t31 3.57113
R39094 C10_N_btm.n0 C10_N_btm.t23 3.57113
R39095 C10_N_btm.n18 C10_N_btm.t2 2.4755
R39096 C10_N_btm.n18 C10_N_btm.t6 2.4755
R39097 C10_N_btm.n16 C10_N_btm.t3 2.4755
R39098 C10_N_btm.n16 C10_N_btm.t4 2.4755
R39099 C10_N_btm.n15 C10_N_btm.t5 2.4755
R39100 C10_N_btm.n15 C10_N_btm.t1 2.4755
R39101 C10_N_btm.n23 C10_N_btm.t17 2.4755
R39102 C10_N_btm.n23 C10_N_btm.t16 2.4755
R39103 C10_N_btm.n30 C10_N_btm.t11 2.4755
R39104 C10_N_btm.n30 C10_N_btm.t10 2.4755
R39105 C10_N_btm.n28 C10_N_btm.t13 2.4755
R39106 C10_N_btm.n28 C10_N_btm.t14 2.4755
R39107 C10_N_btm.n26 C10_N_btm.t15 2.4755
R39108 C10_N_btm.n26 C10_N_btm.t12 2.4755
R39109 C10_N_btm.n25 C10_N_btm.t9 2.4755
R39110 C10_N_btm.n25 C10_N_btm.t8 2.4755
R39111 C10_N_btm.n20 C10_N_btm.t0 2.4755
R39112 C10_N_btm.n20 C10_N_btm.t7 2.4755
R39113 C10_N_btm.n3893 C10_N_btm.t267 1.67819
R39114 C10_N_btm.n3890 C10_N_btm.t533 1.67819
R39115 C10_N_btm.n3887 C10_N_btm.t316 1.67819
R39116 C10_N_btm.n3884 C10_N_btm.t115 1.67819
R39117 C10_N_btm.n3881 C10_N_btm.t363 1.67819
R39118 C10_N_btm.n3878 C10_N_btm.t156 1.67819
R39119 C10_N_btm.n3875 C10_N_btm.t973 1.67819
R39120 C10_N_btm.n3872 C10_N_btm.t252 1.67819
R39121 C10_N_btm.n3869 C10_N_btm.t36 1.67819
R39122 C10_N_btm.n3862 C10_N_btm.t458 1.67819
R39123 C10_N_btm.n3859 C10_N_btm.t748 1.67819
R39124 C10_N_btm.n3856 C10_N_btm.t404 1.67819
R39125 C10_N_btm.n3853 C10_N_btm.t641 1.67819
R39126 C10_N_btm.n3850 C10_N_btm.t875 1.67819
R39127 C10_N_btm.n3847 C10_N_btm.t581 1.67819
R39128 C10_N_btm.n3844 C10_N_btm.t817 1.67819
R39129 C10_N_btm.n3841 C10_N_btm.t515 1.67819
R39130 C10_N_btm.n3838 C10_N_btm.t766 1.67819
R39131 C10_N_btm.n3832 C10_N_btm.t219 1.67819
R39132 C10_N_btm.n3830 C10_N_btm.t373 1.67819
R39133 C10_N_btm.n3827 C10_N_btm.t163 1.67819
R39134 C10_N_btm.n3824 C10_N_btm.t982 1.67819
R39135 C10_N_btm.n3821 C10_N_btm.t206 1.67819
R39136 C10_N_btm.n3818 C10_N_btm.t994 1.67819
R39137 C10_N_btm.n3815 C10_N_btm.t799 1.67819
R39138 C10_N_btm.n3812 C10_N_btm.t98 1.67819
R39139 C10_N_btm.n3809 C10_N_btm.t859 1.67819
R39140 C10_N_btm.n3803 C10_N_btm.t297 1.67819
R39141 C10_N_btm.n3745 C10_N_btm.t570 1.67819
R39142 C10_N_btm.n3748 C10_N_btm.t251 1.67819
R39143 C10_N_btm.n3751 C10_N_btm.t472 1.67819
R39144 C10_N_btm.n3754 C10_N_btm.t700 1.67819
R39145 C10_N_btm.n3757 C10_N_btm.t415 1.67819
R39146 C10_N_btm.n3760 C10_N_btm.t650 1.67819
R39147 C10_N_btm.n3763 C10_N_btm.t881 1.67819
R39148 C10_N_btm.n3766 C10_N_btm.t590 1.67819
R39149 C10_N_btm.n3773 C10_N_btm.t988 1.67819
R39150 C10_N_btm.n3776 C10_N_btm.t218 1.67819
R39151 C10_N_btm.n3779 C10_N_btm.t920 1.67819
R39152 C10_N_btm.n3782 C10_N_btm.t807 1.67819
R39153 C10_N_btm.n3785 C10_N_btm.t99 1.67819
R39154 C10_N_btm.n3788 C10_N_btm.t866 1.67819
R39155 C10_N_btm.n3791 C10_N_btm.t625 1.67819
R39156 C10_N_btm.n3794 C10_N_btm.t970 1.67819
R39157 C10_N_btm.n3797 C10_N_btm.t685 1.67819
R39158 C10_N_btm.n3707 C10_N_btm.t517 1.67819
R39159 C10_N_btm.n3710 C10_N_btm.t288 1.67819
R39160 C10_N_btm.n3713 C10_N_btm.t1036 1.67819
R39161 C10_N_btm.n3716 C10_N_btm.t193 1.67819
R39162 C10_N_btm.n3719 C10_N_btm.t409 1.67819
R39163 C10_N_btm.n3722 C10_N_btm.t148 1.67819
R39164 C10_N_btm.n3725 C10_N_btm.t354 1.67819
R39165 C10_N_btm.n3728 C10_N_btm.t587 1.67819
R39166 C10_N_btm.n3731 C10_N_btm.t308 1.67819
R39167 C10_N_btm.n121 C10_N_btm.t813 1.67819
R39168 C10_N_btm.n119 C10_N_btm.t493 1.67819
R39169 C10_N_btm.n116 C10_N_btm.t870 1.67819
R39170 C10_N_btm.n113 C10_N_btm.t635 1.67819
R39171 C10_N_btm.n110 C10_N_btm.t926 1.67819
R39172 C10_N_btm.n107 C10_N_btm.t692 1.67819
R39173 C10_N_btm.n104 C10_N_btm.t449 1.67819
R39174 C10_N_btm.n101 C10_N_btm.t797 1.67819
R39175 C10_N_btm.n3701 C10_N_btm.t1038 1.67819
R39176 C10_N_btm.n3695 C10_N_btm.t904 1.67819
R39177 C10_N_btm.n3692 C10_N_btm.t134 1.67819
R39178 C10_N_btm.n3689 C10_N_btm.t852 1.67819
R39179 C10_N_btm.n3686 C10_N_btm.t42 1.67819
R39180 C10_N_btm.n3683 C10_N_btm.t255 1.67819
R39181 C10_N_btm.n3680 C10_N_btm.t39 1.67819
R39182 C10_N_btm.n3677 C10_N_btm.t200 1.67819
R39183 C10_N_btm.n3674 C10_N_btm.t420 1.67819
R39184 C10_N_btm.n3671 C10_N_btm.t157 1.67819
R39185 C10_N_btm.n3664 C10_N_btm.t642 1.67819
R39186 C10_N_btm.n3661 C10_N_btm.t933 1.67819
R39187 C10_N_btm.n3658 C10_N_btm.t694 1.67819
R39188 C10_N_btm.n3655 C10_N_btm.t459 1.67819
R39189 C10_N_btm.n3652 C10_N_btm.t751 1.67819
R39190 C10_N_btm.n3649 C10_N_btm.t1048 1.67819
R39191 C10_N_btm.n3646 C10_N_btm.t287 1.67819
R39192 C10_N_btm.n3643 C10_N_btm.t623 1.67819
R39193 C10_N_btm.n3640 C10_N_btm.t345 1.67819
R39194 C10_N_btm.n3634 C10_N_btm.t726 1.67819
R39195 C10_N_btm.n154 C10_N_btm.t96 1.67819
R39196 C10_N_btm.n157 C10_N_btm.t678 1.67819
R39197 C10_N_btm.n160 C10_N_btm.t913 1.67819
R39198 C10_N_btm.n163 C10_N_btm.t101 1.67819
R39199 C10_N_btm.n166 C10_N_btm.t860 1.67819
R39200 C10_N_btm.n169 C10_N_btm.t52 1.67819
R39201 C10_N_btm.n172 C10_N_btm.t262 1.67819
R39202 C10_N_btm.n174 C10_N_btm.t979 1.67819
R39203 C10_N_btm.n3604 C10_N_btm.t350 1.67819
R39204 C10_N_btm.n3607 C10_N_btm.t638 1.67819
R39205 C10_N_btm.n3610 C10_N_btm.t401 1.67819
R39206 C10_N_btm.n3613 C10_N_btm.t188 1.67819
R39207 C10_N_btm.n3616 C10_N_btm.t452 1.67819
R39208 C10_N_btm.n3619 C10_N_btm.t773 1.67819
R39209 C10_N_btm.n3622 C10_N_btm.t103 1.67819
R39210 C10_N_btm.n3625 C10_N_btm.t340 1.67819
R39211 C10_N_btm.n3628 C10_N_btm.t74 1.67819
R39212 C10_N_btm.n3573 C10_N_btm.t551 1.67819
R39213 C10_N_btm.n3576 C10_N_btm.t848 1.67819
R39214 C10_N_btm.n3579 C10_N_btm.t503 1.67819
R39215 C10_N_btm.n3582 C10_N_btm.t735 1.67819
R39216 C10_N_btm.n3585 C10_N_btm.t971 1.67819
R39217 C10_N_btm.n3588 C10_N_btm.t687 1.67819
R39218 C10_N_btm.n3591 C10_N_btm.t918 1.67819
R39219 C10_N_btm.n3594 C10_N_btm.t113 1.67819
R39220 C10_N_btm.n3597 C10_N_btm.t868 1.67819
R39221 C10_N_btm.n227 C10_N_btm.t194 1.67819
R39222 C10_N_btm.n225 C10_N_btm.t464 1.67819
R39223 C10_N_btm.n222 C10_N_btm.t249 1.67819
R39224 C10_N_btm.n219 C10_N_btm.t34 1.67819
R39225 C10_N_btm.n216 C10_N_btm.t292 1.67819
R39226 C10_N_btm.n213 C10_N_btm.t80 1.67819
R39227 C10_N_btm.n210 C10_N_btm.t897 1.67819
R39228 C10_N_btm.n207 C10_N_btm.t182 1.67819
R39229 C10_N_btm.n3567 C10_N_btm.t956 1.67819
R39230 C10_N_btm.n3561 C10_N_btm.t1052 1.67819
R39231 C10_N_btm.n3558 C10_N_btm.t676 1.67819
R39232 C10_N_btm.n3555 C10_N_btm.t339 1.67819
R39233 C10_N_btm.n3552 C10_N_btm.t560 1.67819
R39234 C10_N_btm.n3549 C10_N_btm.t798 1.67819
R39235 C10_N_btm.n3546 C10_N_btm.t1040 1.67819
R39236 C10_N_btm.n3543 C10_N_btm.t744 1.67819
R39237 C10_N_btm.n3540 C10_N_btm.t981 1.67819
R39238 C10_N_btm.n3537 C10_N_btm.t693 1.67819
R39239 C10_N_btm.n3530 C10_N_btm.t44 1.67819
R39240 C10_N_btm.n3527 C10_N_btm.t301 1.67819
R39241 C10_N_btm.n3524 C10_N_btm.t88 1.67819
R39242 C10_N_btm.n3521 C10_N_btm.t907 1.67819
R39243 C10_N_btm.n3518 C10_N_btm.t135 1.67819
R39244 C10_N_btm.n3515 C10_N_btm.t962 1.67819
R39245 C10_N_btm.n3512 C10_N_btm.t717 1.67819
R39246 C10_N_btm.n3509 C10_N_btm.t86 1.67819
R39247 C10_N_btm.n3506 C10_N_btm.t785 1.67819
R39248 C10_N_btm.n3500 C10_N_btm.t993 1.67819
R39249 C10_N_btm.n260 C10_N_btm.t385 1.67819
R39250 C10_N_btm.n263 C10_N_btm.t67 1.67819
R39251 C10_N_btm.n266 C10_N_btm.t282 1.67819
R39252 C10_N_btm.n269 C10_N_btm.t506 1.67819
R39253 C10_N_btm.n272 C10_N_btm.t511 1.67819
R39254 C10_N_btm.n275 C10_N_btm.t446 1.67819
R39255 C10_N_btm.n278 C10_N_btm.t690 1.67819
R39256 C10_N_btm.n280 C10_N_btm.t396 1.67819
R39257 C10_N_btm.n3470 C10_N_btm.t914 1.67819
R39258 C10_N_btm.n3473 C10_N_btm.t147 1.67819
R39259 C10_N_btm.n3476 C10_N_btm.t965 1.67819
R39260 C10_N_btm.n3479 C10_N_btm.t727 1.67819
R39261 C10_N_btm.n3482 C10_N_btm.t223 1.67819
R39262 C10_N_btm.n3485 C10_N_btm.t789 1.67819
R39263 C10_N_btm.n3488 C10_N_btm.t542 1.67819
R39264 C10_N_btm.n3491 C10_N_btm.t893 1.67819
R39265 C10_N_btm.n3494 C10_N_btm.t607 1.67819
R39266 C10_N_btm.n3439 C10_N_btm.t1006 1.67819
R39267 C10_N_btm.n3442 C10_N_btm.t467 1.67819
R39268 C10_N_btm.n3445 C10_N_btm.t950 1.67819
R39269 C10_N_btm.n3448 C10_N_btm.t126 1.67819
R39270 C10_N_btm.n3451 C10_N_btm.t341 1.67819
R39271 C10_N_btm.n3454 C10_N_btm.t75 1.67819
R39272 C10_N_btm.n3457 C10_N_btm.t286 1.67819
R39273 C10_N_btm.n3460 C10_N_btm.t1042 1.67819
R39274 C10_N_btm.n3463 C10_N_btm.t906 1.67819
R39275 C10_N_btm.n333 C10_N_btm.t736 1.67819
R39276 C10_N_btm.n331 C10_N_btm.t478 1.67819
R39277 C10_N_btm.n328 C10_N_btm.t792 1.67819
R39278 C10_N_btm.n325 C10_N_btm.t552 1.67819
R39279 C10_N_btm.n322 C10_N_btm.t851 1.67819
R39280 C10_N_btm.n319 C10_N_btm.t614 1.67819
R39281 C10_N_btm.n316 C10_N_btm.t1041 1.67819
R39282 C10_N_btm.n313 C10_N_btm.t713 1.67819
R39283 C10_N_btm.n3433 C10_N_btm.t434 1.67819
R39284 C10_N_btm.n3427 C10_N_btm.t829 1.67819
R39285 C10_N_btm.n3424 C10_N_btm.t65 1.67819
R39286 C10_N_btm.n3421 C10_N_btm.t779 1.67819
R39287 C10_N_btm.n3418 C10_N_btm.t1017 1.67819
R39288 C10_N_btm.n3415 C10_N_btm.t184 1.67819
R39289 C10_N_btm.n3412 C10_N_btm.t957 1.67819
R39290 C10_N_btm.n3409 C10_N_btm.t132 1.67819
R39291 C10_N_btm.n3406 C10_N_btm.t347 1.67819
R39292 C10_N_btm.n3403 C10_N_btm.t81 1.67819
R39293 C10_N_btm.n3396 C10_N_btm.t441 1.67819
R39294 C10_N_btm.n3393 C10_N_btm.t731 1.67819
R39295 C10_N_btm.n3390 C10_N_btm.t1027 1.67819
R39296 C10_N_btm.n3387 C10_N_btm.t277 1.67819
R39297 C10_N_btm.n3384 C10_N_btm.t546 1.67819
R39298 C10_N_btm.n3381 C10_N_btm.t331 1.67819
R39299 C10_N_btm.n3378 C10_N_btm.t244 1.67819
R39300 C10_N_btm.n3375 C10_N_btm.t428 1.67819
R39301 C10_N_btm.n3372 C10_N_btm.t172 1.67819
R39302 C10_N_btm.n3366 C10_N_btm.t215 1.67819
R39303 C10_N_btm.n366 C10_N_btm.t498 1.67819
R39304 C10_N_btm.n369 C10_N_btm.t166 1.67819
R39305 C10_N_btm.n372 C10_N_btm.t377 1.67819
R39306 C10_N_btm.n375 C10_N_btm.t605 1.67819
R39307 C10_N_btm.n378 C10_N_btm.t326 1.67819
R39308 C10_N_btm.n381 C10_N_btm.t540 1.67819
R39309 C10_N_btm.n384 C10_N_btm.t388 1.67819
R39310 C10_N_btm.n386 C10_N_btm.t991 1.67819
R39311 C10_N_btm.n3336 C10_N_btm.t888 1.67819
R39312 C10_N_btm.n3339 C10_N_btm.t124 1.67819
R39313 C10_N_btm.n3342 C10_N_btm.t948 1.67819
R39314 C10_N_btm.n3345 C10_N_btm.t705 1.67819
R39315 C10_N_btm.n3348 C10_N_btm.t1004 1.67819
R39316 C10_N_btm.n3351 C10_N_btm.t769 1.67819
R39317 C10_N_btm.n3354 C10_N_btm.t525 1.67819
R39318 C10_N_btm.n3357 C10_N_btm.t874 1.67819
R39319 C10_N_btm.n3360 C10_N_btm.t583 1.67819
R39320 C10_N_btm.n3305 C10_N_btm.t476 1.67819
R39321 C10_N_btm.n3308 C10_N_btm.t320 1.67819
R39322 C10_N_btm.n3311 C10_N_btm.t738 1.67819
R39323 C10_N_btm.n3314 C10_N_btm.t234 1.67819
R39324 C10_N_btm.n3317 C10_N_btm.t433 1.67819
R39325 C10_N_btm.n3320 C10_N_btm.t174 1.67819
R39326 C10_N_btm.n3323 C10_N_btm.t384 1.67819
R39327 C10_N_btm.n3326 C10_N_btm.t613 1.67819
R39328 C10_N_btm.n3329 C10_N_btm.t335 1.67819
R39329 C10_N_btm.n468 C10_N_btm.t954 1.67819
R39330 C10_N_btm.n465 C10_N_btm.t710 1.67819
R39331 C10_N_btm.n462 C10_N_btm.t1014 1.67819
R39332 C10_N_btm.n459 C10_N_btm.t776 1.67819
R39333 C10_N_btm.n456 C10_N_btm.t1057 1.67819
R39334 C10_N_btm.n453 C10_N_btm.t827 1.67819
R39335 C10_N_btm.n450 C10_N_btm.t592 1.67819
R39336 C10_N_btm.n447 C10_N_btm.t360 1.67819
R39337 C10_N_btm.n444 C10_N_btm.t698 1.67819
R39338 C10_N_btm.n3299 C10_N_btm.t417 1.67819
R39339 C10_N_btm.n3293 C10_N_btm.t808 1.67819
R39340 C10_N_btm.n3290 C10_N_btm.t93 1.67819
R39341 C10_N_btm.n3287 C10_N_btm.t753 1.67819
R39342 C10_N_btm.n3284 C10_N_btm.t989 1.67819
R39343 C10_N_btm.n3281 C10_N_btm.t171 1.67819
R39344 C10_N_btm.n3278 C10_N_btm.t935 1.67819
R39345 C10_N_btm.n3275 C10_N_btm.t241 1.67819
R39346 C10_N_btm.n3272 C10_N_btm.t330 1.67819
R39347 C10_N_btm.n3269 C10_N_btm.t59 1.67819
R39348 C10_N_btm.n3266 C10_N_btm.t276 1.67819
R39349 C10_N_btm.n3263 C10_N_btm.t1011 1.67819
R39350 C10_N_btm.n3260 C10_N_btm.t471 1.67819
R39351 C10_N_btm.n3257 C10_N_btm.t440 1.67819
R39352 C10_N_btm.n3254 C10_N_btm.t741 1.67819
R39353 C10_N_btm.n3251 C10_N_btm.t976 1.67819
R39354 C10_N_btm.n3248 C10_N_btm.t201 1.67819
R39355 C10_N_btm.n3245 C10_N_btm.t922 1.67819
R39356 C10_N_btm.n3242 C10_N_btm.t119 1.67819
R39357 C10_N_btm.n3239 C10_N_btm.t365 1.67819
R39358 C10_N_btm.n3236 C10_N_btm.t220 1.67819
R39359 C10_N_btm.n3233 C10_N_btm.t268 1.67819
R39360 C10_N_btm.n3230 C10_N_btm.t793 1.67819
R39361 C10_N_btm.n3227 C10_N_btm.t228 1.67819
R39362 C10_N_btm.n504 C10_N_btm.t951 1.67819
R39363 C10_N_btm.n501 C10_N_btm.t180 1.67819
R39364 C10_N_btm.n498 C10_N_btm.t1008 1.67819
R39365 C10_N_btm.n495 C10_N_btm.t274 1.67819
R39366 C10_N_btm.n492 C10_N_btm.t83 1.67819
R39367 C10_N_btm.n489 C10_N_btm.t821 1.67819
R39368 C10_N_btm.n486 C10_N_btm.t236 1.67819
R39369 C10_N_btm.n483 C10_N_btm.t878 1.67819
R39370 C10_N_btm.n480 C10_N_btm.t647 1.67819
R39371 C10_N_btm.n477 C10_N_btm.t78 1.67819
R39372 C10_N_btm.n474 C10_N_btm.t895 1.67819
R39373 C10_N_btm.n471 C10_N_btm.t608 1.67819
R39374 C10_N_btm.n3224 C10_N_btm.t431 1.67819
R39375 C10_N_btm.n3221 C10_N_btm.t485 1.67819
R39376 C10_N_btm.n3218 C10_N_btm.t1039 1.67819
R39377 C10_N_btm.n3215 C10_N_btm.t611 1.67819
R39378 C10_N_btm.n3212 C10_N_btm.t279 1.67819
R39379 C10_N_btm.n3209 C10_N_btm.t547 1.67819
R39380 C10_N_btm.n3206 C10_N_btm.t488 1.67819
R39381 C10_N_btm.n3203 C10_N_btm.t443 1.67819
R39382 C10_N_btm.n3200 C10_N_btm.t732 1.67819
R39383 C10_N_btm.n3197 C10_N_btm.t392 1.67819
R39384 C10_N_btm.n3194 C10_N_btm.t622 1.67819
R39385 C10_N_btm.n3191 C10_N_btm.t865 1.67819
R39386 C10_N_btm.n3188 C10_N_btm.t564 1.67819
R39387 C10_N_btm.n3185 C10_N_btm.t804 1.67819
R39388 C10_N_btm.n3182 C10_N_btm.t457 1.67819
R39389 C10_N_btm.n3179 C10_N_btm.t747 1.67819
R39390 C10_N_btm.n3176 C10_N_btm.t986 1.67819
R39391 C10_N_btm.n3173 C10_N_btm.t686 1.67819
R39392 C10_N_btm.n3170 C10_N_btm.t969 1.67819
R39393 C10_N_btm.n3167 C10_N_btm.t154 1.67819
R39394 C10_N_btm.n3164 C10_N_btm.t867 1.67819
R39395 C10_N_btm.n3161 C10_N_btm.t102 1.67819
R39396 C10_N_btm.n3158 C10_N_btm.t314 1.67819
R39397 C10_N_btm.n3155 C10_N_btm.t924 1.67819
R39398 C10_N_btm.n3152 C10_N_btm.t224 1.67819
R39399 C10_N_btm.n3149 C10_N_btm.t987 1.67819
R39400 C10_N_btm.n3146 C10_N_btm.t167 1.67819
R39401 C10_N_btm.n3143 C10_N_btm.t379 1.67819
R39402 C10_N_btm.n3140 C10_N_btm.t233 1.67819
R39403 C10_N_btm.n3137 C10_N_btm.t327 1.67819
R39404 C10_N_btm.n3134 C10_N_btm.t543 1.67819
R39405 C10_N_btm.n3131 C10_N_btm.t474 1.67819
R39406 C10_N_btm.n3128 C10_N_btm.t1012 1.67819
R39407 C10_N_btm.n3125 C10_N_btm.t179 1.67819
R39408 C10_N_btm.n3122 C10_N_btm.t389 1.67819
R39409 C10_N_btm.n3119 C10_N_btm.t679 1.67819
R39410 C10_N_btm.n3116 C10_N_btm.t342 1.67819
R39411 C10_N_btm.n3113 C10_N_btm.t563 1.67819
R39412 C10_N_btm.n3110 C10_N_btm.t861 1.67819
R39413 C10_N_btm.n3103 C10_N_btm.t757 1.67819
R39414 C10_N_btm.n3100 C10_N_btm.t239 1.67819
R39415 C10_N_btm.n3097 C10_N_btm.t361 1.67819
R39416 C10_N_btm.n3094 C10_N_btm.t321 1.67819
R39417 C10_N_btm.n3091 C10_N_btm.t516 1.67819
R39418 C10_N_btm.n3088 C10_N_btm.t872 1.67819
R39419 C10_N_btm.n3085 C10_N_btm.t162 1.67819
R39420 C10_N_btm.n3082 C10_N_btm.t928 1.67819
R39421 C10_N_btm.n3079 C10_N_btm.t205 1.67819
R39422 C10_N_btm.n3076 C10_N_btm.t1055 1.67819
R39423 C10_N_btm.n3073 C10_N_btm.t394 1.67819
R39424 C10_N_btm.n3070 C10_N_btm.t50 1.67819
R39425 C10_N_btm.n3067 C10_N_btm.t858 1.67819
R39426 C10_N_btm.n3064 C10_N_btm.t618 1.67819
R39427 C10_N_btm.n3061 C10_N_btm.t912 1.67819
R39428 C10_N_btm.n3058 C10_N_btm.t677 1.67819
R39429 C10_N_btm.n3055 C10_N_btm.t48 1.67819
R39430 C10_N_btm.n3052 C10_N_btm.t724 1.67819
R39431 C10_N_btm.n3049 C10_N_btm.t974 1.67819
R39432 C10_N_btm.n3046 C10_N_btm.t843 1.67819
R39433 C10_N_btm.n3043 C10_N_btm.t604 1.67819
R39434 C10_N_btm.n3040 C10_N_btm.t325 1.67819
R39435 C10_N_btm.n3037 C10_N_btm.t617 1.67819
R39436 C10_N_btm.n3034 C10_N_btm.t387 1.67819
R39437 C10_N_btm.n3031 C10_N_btm.t121 1.67819
R39438 C10_N_btm.n3028 C10_N_btm.t439 1.67819
R39439 C10_N_btm.n3025 C10_N_btm.t243 1.67819
R39440 C10_N_btm.n3022 C10_N_btm.t905 1.67819
R39441 C10_N_btm.n3019 C10_N_btm.t272 1.67819
R39442 C10_N_btm.n3016 C10_N_btm.t57 1.67819
R39443 C10_N_btm.n3013 C10_N_btm.t375 1.67819
R39444 C10_N_btm.n3010 C10_N_btm.t229 1.67819
R39445 C10_N_btm.n3007 C10_N_btm.t931 1.67819
R39446 C10_N_btm.n3004 C10_N_btm.t211 1.67819
R39447 C10_N_btm.n3001 C10_N_btm.t985 1.67819
R39448 C10_N_btm.n2998 C10_N_btm.t265 1.67819
R39449 C10_N_btm.n2995 C10_N_btm.t56 1.67819
R39450 C10_N_btm.n2992 C10_N_btm.t803 1.67819
R39451 C10_N_btm.n2989 C10_N_btm.t107 1.67819
R39452 C10_N_btm.n2986 C10_N_btm.t916 1.67819
R39453 C10_N_btm.n2983 C10_N_btm.t680 1.67819
R39454 C10_N_btm.n2980 C10_N_btm.t968 1.67819
R39455 C10_N_btm.n2977 C10_N_btm.t730 1.67819
R39456 C10_N_btm.n2974 C10_N_btm.t1034 1.67819
R39457 C10_N_btm.n2971 C10_N_btm.t790 1.67819
R39458 C10_N_btm.n2968 C10_N_btm.t545 1.67819
R39459 C10_N_btm.n2965 C10_N_btm.t896 1.67819
R39460 C10_N_btm.n2962 C10_N_btm.t609 1.67819
R39461 C10_N_btm.n2959 C10_N_btm.t382 1.67819
R39462 C10_N_btm.n2956 C10_N_btm.t961 1.67819
R39463 C10_N_btm.n2953 C10_N_btm.t715 1.67819
R39464 C10_N_btm.n2950 C10_N_btm.t436 1.67819
R39465 C10_N_btm.n2947 C10_N_btm.t784 1.67819
R39466 C10_N_btm.n2944 C10_N_btm.t537 1.67819
R39467 C10_N_btm.n2941 C10_N_btm.t836 1.67819
R39468 C10_N_btm.n2938 C10_N_btm.t294 1.67819
R39469 C10_N_btm.n2935 C10_N_btm.t371 1.67819
R39470 C10_N_btm.n2932 C10_N_btm.t658 1.67819
R39471 C10_N_btm.n2929 C10_N_btm.t425 1.67819
R39472 C10_N_btm.n2926 C10_N_btm.t204 1.67819
R39473 C10_N_btm.n2923 C10_N_btm.t522 1.67819
R39474 C10_N_btm.n2920 C10_N_btm.t261 1.67819
R39475 C10_N_btm.n2914 C10_N_btm.t637 1.67819
R39476 C10_N_btm.n1786 C10_N_btm.t925 1.67819
R39477 C10_N_btm.n1789 C10_N_btm.t575 1.67819
R39478 C10_N_btm.n1792 C10_N_btm.t815 1.67819
R39479 C10_N_btm.n1795 C10_N_btm.t573 1.67819
R39480 C10_N_btm.n1798 C10_N_btm.t761 1.67819
R39481 C10_N_btm.n1801 C10_N_btm.t996 1.67819
R39482 C10_N_btm.n1804 C10_N_btm.t176 1.67819
R39483 C10_N_btm.n1807 C10_N_btm.t942 1.67819
R39484 C10_N_btm.n1810 C10_N_btm.t774 1.67819
R39485 C10_N_btm.n1813 C10_N_btm.t833 1.67819
R39486 C10_N_btm.n1816 C10_N_btm.t66 1.67819
R39487 C10_N_btm.n1819 C10_N_btm.t281 1.67819
R39488 C10_N_btm.n1822 C10_N_btm.t486 1.67819
R39489 C10_N_btm.n1825 C10_N_btm.t703 1.67819
R39490 C10_N_btm.n1828 C10_N_btm.t997 1.67819
R39491 C10_N_btm.n1831 C10_N_btm.t655 1.67819
R39492 C10_N_btm.n1834 C10_N_btm.t884 1.67819
R39493 C10_N_btm.n1837 C10_N_btm.t1032 1.67819
R39494 C10_N_btm.n1840 C10_N_btm.t412 1.67819
R39495 C10_N_btm.n1843 C10_N_btm.t532 1.67819
R39496 C10_N_btm.n1846 C10_N_btm.t781 1.67819
R39497 C10_N_btm.n1849 C10_N_btm.t1018 1.67819
R39498 C10_N_btm.n1852 C10_N_btm.t185 1.67819
R39499 C10_N_btm.n1855 C10_N_btm.t900 1.67819
R39500 C10_N_btm.n1858 C10_N_btm.t1051 1.67819
R39501 C10_N_btm.n1861 C10_N_btm.t349 1.67819
R39502 C10_N_btm.n1864 C10_N_btm.t37 1.67819
R39503 C10_N_btm.n1867 C10_N_btm.t295 1.67819
R39504 C10_N_btm.n1870 C10_N_btm.t95 1.67819
R39505 C10_N_btm.n1873 C10_N_btm.t196 1.67819
R39506 C10_N_btm.n1876 C10_N_btm.t469 1.67819
R39507 C10_N_btm.n1879 C10_N_btm.t153 1.67819
R39508 C10_N_btm.n1882 C10_N_btm.t357 1.67819
R39509 C10_N_btm.n1885 C10_N_btm.t589 1.67819
R39510 C10_N_btm.n1888 C10_N_btm.t313 1.67819
R39511 C10_N_btm.n1891 C10_N_btm.t530 1.67819
R39512 C10_N_btm.n1894 C10_N_btm.t214 1.67819
R39513 C10_N_btm.n1897 C10_N_btm.t497 1.67819
R39514 C10_N_btm.n1900 C10_N_btm.t709 1.67819
R39515 C10_N_btm.n1903 C10_N_btm.t416 1.67819
R39516 C10_N_btm.n1906 C10_N_btm.t699 1.67819
R39517 C10_N_btm.n1909 C10_N_btm.t940 1.67819
R39518 C10_N_btm.n1912 C10_N_btm.t591 1.67819
R39519 C10_N_btm.n1915 C10_N_btm.t826 1.67819
R39520 C10_N_btm.n1918 C10_N_btm.t64 1.67819
R39521 C10_N_btm.n1921 C10_N_btm.t777 1.67819
R39522 C10_N_btm.n1924 C10_N_btm.t1029 1.67819
R39523 C10_N_btm.n1927 C10_N_btm.t711 1.67819
R39524 C10_N_btm.n1930 C10_N_btm.t955 1.67819
R39525 C10_N_btm.n1933 C10_N_btm.t130 1.67819
R39526 C10_N_btm.n1936 C10_N_btm.t894 1.67819
R39527 C10_N_btm.n1939 C10_N_btm.t79 1.67819
R39528 C10_N_btm.n1942 C10_N_btm.t290 1.67819
R39529 C10_N_btm.n1945 C10_N_btm.t40 1.67819
R39530 C10_N_btm.n1948 C10_N_btm.t248 1.67819
R39531 C10_N_btm.n1951 C10_N_btm.t967 1.67819
R39532 C10_N_btm.n1954 C10_N_btm.t149 1.67819
R39533 C10_N_btm.n1957 C10_N_btm.t408 1.67819
R39534 C10_N_btm.n1960 C10_N_btm.t105 1.67819
R39535 C10_N_btm.n1963 C10_N_btm.t311 1.67819
R39536 C10_N_btm.n1965 C10_N_btm.t586 1.67819
R39537 C10_N_btm.n2725 C10_N_btm.t620 1.67819
R39538 C10_N_btm.n2728 C10_N_btm.t1023 1.67819
R39539 C10_N_btm.n2731 C10_N_btm.t787 1.67819
R39540 C10_N_btm.n2734 C10_N_btm.t72 1.67819
R39541 C10_N_btm.n2737 C10_N_btm.t839 1.67819
R39542 C10_N_btm.n2740 C10_N_btm.t602 1.67819
R39543 C10_N_btm.n2743 C10_N_btm.t947 1.67819
R39544 C10_N_btm.n2746 C10_N_btm.t660 1.67819
R39545 C10_N_btm.n2749 C10_N_btm.t1002 1.67819
R39546 C10_N_btm.n2752 C10_N_btm.t768 1.67819
R39547 C10_N_btm.n2755 C10_N_btm.t524 1.67819
R39548 C10_N_btm.n2758 C10_N_btm.t818 1.67819
R39549 C10_N_btm.n2761 C10_N_btm.t582 1.67819
R39550 C10_N_btm.n2764 C10_N_btm.t353 1.67819
R39551 C10_N_btm.n2767 C10_N_btm.t643 1.67819
R39552 C10_N_btm.n2770 C10_N_btm.t405 1.67819
R39553 C10_N_btm.n2773 C10_N_btm.t749 1.67819
R39554 C10_N_btm.n2776 C10_N_btm.t460 1.67819
R39555 C10_N_btm.n2779 C10_N_btm.t1031 1.67819
R39556 C10_N_btm.n2782 C10_N_btm.t566 1.67819
R39557 C10_N_btm.n2785 C10_N_btm.t344 1.67819
R39558 C10_N_btm.n2788 C10_N_btm.t77 1.67819
R39559 C10_N_btm.n2791 C10_N_btm.t352 1.67819
R39560 C10_N_btm.n2794 C10_N_btm.t142 1.67819
R39561 C10_N_btm.n2797 C10_N_btm.t911 1.67819
R39562 C10_N_btm.n2800 C10_N_btm.t192 1.67819
R39563 C10_N_btm.n2803 C10_N_btm.t1037 1.67819
R39564 C10_N_btm.n2806 C10_N_btm.t1013 1.67819
R39565 C10_N_btm.n2809 C10_N_btm.t238 1.67819
R39566 C10_N_btm.n2812 C10_N_btm.t842 1.67819
R39567 C10_N_btm.n2815 C10_N_btm.t128 1.67819
R39568 C10_N_btm.n2818 C10_N_btm.t891 1.67819
R39569 C10_N_btm.n2821 C10_N_btm.t665 1.67819
R39570 C10_N_btm.n2824 C10_N_btm.t1010 1.67819
R39571 C10_N_btm.n2827 C10_N_btm.t708 1.67819
R39572 C10_N_btm.n2830 C10_N_btm.t41 1.67819
R39573 C10_N_btm.n2833 C10_N_btm.t823 1.67819
R39574 C10_N_btm.n2836 C10_N_btm.t529 1.67819
R39575 C10_N_btm.n2839 C10_N_btm.t880 1.67819
R39576 C10_N_btm.n2842 C10_N_btm.t648 1.67819
R39577 C10_N_btm.n2845 C10_N_btm.t411 1.67819
R39578 C10_N_btm.n2848 C10_N_btm.t697 1.67819
R39579 C10_N_btm.n2851 C10_N_btm.t465 1.67819
R39580 C10_N_btm.n2854 C10_N_btm.t809 1.67819
R39581 C10_N_btm.n2857 C10_N_btm.t1050 1.67819
R39582 C10_N_btm.n2860 C10_N_btm.t143 1.67819
R39583 C10_N_btm.n2863 C10_N_btm.t627 1.67819
R39584 C10_N_btm.n2866 C10_N_btm.t348 1.67819
R39585 C10_N_btm.n2869 C10_N_btm.t133 1.67819
R39586 C10_N_btm.n2872 C10_N_btm.t788 1.67819
R39587 C10_N_btm.n2875 C10_N_btm.t541 1.67819
R39588 C10_N_btm.n2878 C10_N_btm.t275 1.67819
R39589 C10_N_btm.n2881 C10_N_btm.t606 1.67819
R39590 C10_N_btm.n2884 C10_N_btm.t378 1.67819
R39591 C10_N_btm.n2887 C10_N_btm.t666 1.67819
R39592 C10_N_btm.n2890 C10_N_btm.t427 1.67819
R39593 C10_N_btm.n2893 C10_N_btm.t217 1.67819
R39594 C10_N_btm.n2896 C10_N_btm.t510 1.67819
R39595 C10_N_btm.n2899 C10_N_btm.t266 1.67819
R39596 C10_N_btm.n2902 C10_N_btm.t89 1.67819
R39597 C10_N_btm.n2905 C10_N_btm.t358 1.67819
R39598 C10_N_btm.n2908 C10_N_btm.t108 1.67819
R39599 C10_N_btm.n2535 C10_N_btm.t461 1.67819
R39600 C10_N_btm.n2538 C10_N_btm.t750 1.67819
R39601 C10_N_btm.n2541 C10_N_btm.t406 1.67819
R39602 C10_N_btm.n2544 C10_N_btm.t644 1.67819
R39603 C10_N_btm.n2547 C10_N_btm.t877 1.67819
R39604 C10_N_btm.n2550 C10_N_btm.t584 1.67819
R39605 C10_N_btm.n2553 C10_N_btm.t819 1.67819
R39606 C10_N_btm.n2556 C10_N_btm.t116 1.67819
R39607 C10_N_btm.n2559 C10_N_btm.t770 1.67819
R39608 C10_N_btm.n2562 C10_N_btm.t1005 1.67819
R39609 C10_N_btm.n2565 C10_N_btm.t661 1.67819
R39610 C10_N_btm.n2568 C10_N_btm.t949 1.67819
R39611 C10_N_btm.n2571 C10_N_btm.t125 1.67819
R39612 C10_N_btm.n2574 C10_N_btm.t242 1.67819
R39613 C10_N_btm.n2577 C10_N_btm.t438 1.67819
R39614 C10_N_btm.n2580 C10_N_btm.t719 1.67819
R39615 C10_N_btm.n2583 C10_N_btm.t1047 1.67819
R39616 C10_N_btm.n2586 C10_N_btm.t616 1.67819
R39617 C10_N_btm.n2589 C10_N_btm.t908 1.67819
R39618 C10_N_btm.n2592 C10_N_btm.t558 1.67819
R39619 C10_N_btm.n2595 C10_N_btm.t796 1.67819
R39620 C10_N_btm.n2598 C10_N_btm.t507 1.67819
R39621 C10_N_btm.n2601 C10_N_btm.t742 1.67819
R39622 C10_N_btm.n2604 C10_N_btm.t978 1.67819
R39623 C10_N_btm.n2607 C10_N_btm.t631 1.67819
R39624 C10_N_btm.n2610 C10_N_btm.t923 1.67819
R39625 C10_N_btm.n2613 C10_N_btm.t216 1.67819
R39626 C10_N_btm.n2616 C10_N_btm.t811 1.67819
R39627 C10_N_btm.n2619 C10_N_btm.t230 1.67819
R39628 C10_N_btm.n2622 C10_N_btm.t374 1.67819
R39629 C10_N_btm.n2625 C10_N_btm.t990 1.67819
R39630 C10_N_btm.n2628 C10_N_btm.t231 1.67819
R39631 C10_N_btm.n2631 C10_N_btm.t939 1.67819
R39632 C10_N_btm.n2634 C10_N_btm.t492 1.67819
R39633 C10_N_btm.n2637 C10_N_btm.t334 1.67819
R39634 C10_N_btm.n2640 C10_N_btm.t63 1.67819
R39635 C10_N_btm.n2643 C10_N_btm.t280 1.67819
R39636 C10_N_btm.n2646 C10_N_btm.t1026 1.67819
R39637 C10_N_btm.n2649 C10_N_btm.t491 1.67819
R39638 C10_N_btm.n2652 C10_N_btm.t444 1.67819
R39639 C10_N_btm.n2655 C10_N_btm.t175 1.67819
R39640 C10_N_btm.n2658 C10_N_btm.t432 1.67819
R39641 C10_N_btm.n2661 C10_N_btm.t672 1.67819
R39642 C10_N_btm.n2664 C10_N_btm.t336 1.67819
R39643 C10_N_btm.n2667 C10_N_btm.t553 1.67819
R39644 C10_N_btm.n2670 C10_N_btm.t849 1.67819
R39645 C10_N_btm.n2673 C10_N_btm.t504 1.67819
R39646 C10_N_btm.n2676 C10_N_btm.t737 1.67819
R39647 C10_N_btm.n2679 C10_N_btm.t445 1.67819
R39648 C10_N_btm.n2682 C10_N_btm.t688 1.67819
R39649 C10_N_btm.n2685 C10_N_btm.t919 1.67819
R39650 C10_N_btm.n2688 C10_N_btm.t626 1.67819
R39651 C10_N_btm.n2691 C10_N_btm.t869 1.67819
R39652 C10_N_btm.n2694 C10_N_btm.t114 1.67819
R39653 C10_N_btm.n2697 C10_N_btm.t754 1.67819
R39654 C10_N_btm.n2700 C10_N_btm.t812 1.67819
R39655 C10_N_btm.n2703 C10_N_btm.t696 1.67819
R39656 C10_N_btm.n2706 C10_N_btm.t936 1.67819
R39657 C10_N_btm.n2709 C10_N_btm.t170 1.67819
R39658 C10_N_btm.n2712 C10_N_btm.t879 1.67819
R39659 C10_N_btm.n2715 C10_N_btm.t61 1.67819
R39660 C10_N_btm.n2718 C10_N_btm.t329 1.67819
R39661 C10_N_btm.n2335 C10_N_btm.t422 1.67819
R39662 C10_N_btm.n2333 C10_N_btm.t160 1.67819
R39663 C10_N_btm.n2330 C10_N_btm.t977 1.67819
R39664 C10_N_btm.n2327 C10_N_btm.t258 1.67819
R39665 C10_N_btm.n2324 C10_N_btm.t43 1.67819
R39666 C10_N_btm.n2321 C10_N_btm.t795 1.67819
R39667 C10_N_btm.n2318 C10_N_btm.t92 1.67819
R39668 C10_N_btm.n2315 C10_N_btm.t853 1.67819
R39669 C10_N_btm.n2312 C10_N_btm.t137 1.67819
R39670 C10_N_btm.n2309 C10_N_btm.t963 1.67819
R39671 C10_N_btm.n2306 C10_N_btm.t718 1.67819
R39672 C10_N_btm.n2303 C10_N_btm.t1022 1.67819
R39673 C10_N_btm.n2300 C10_N_btm.t786 1.67819
R39674 C10_N_btm.n2297 C10_N_btm.t539 1.67819
R39675 C10_N_btm.n2294 C10_N_btm.t837 1.67819
R39676 C10_N_btm.n2291 C10_N_btm.t601 1.67819
R39677 C10_N_btm.n2288 C10_N_btm.t946 1.67819
R39678 C10_N_btm.n2285 C10_N_btm.t659 1.67819
R39679 C10_N_btm.n2282 C10_N_btm.t426 1.67819
R39680 C10_N_btm.n2279 C10_N_btm.t767 1.67819
R39681 C10_N_btm.n2276 C10_N_btm.t523 1.67819
R39682 C10_N_btm.n2273 C10_N_btm.t263 1.67819
R39683 C10_N_btm.n2270 C10_N_btm.t536 1.67819
R39684 C10_N_btm.n2267 C10_N_btm.t319 1.67819
R39685 C10_N_btm.n2264 C10_N_btm.t245 1.67819
R39686 C10_N_btm.n2261 C10_N_btm.t369 1.67819
R39687 C10_N_btm.n2258 C10_N_btm.t161 1.67819
R39688 C10_N_btm.n2255 C10_N_btm.t424 1.67819
R39689 C10_N_btm.n2252 C10_N_btm.t203 1.67819
R39690 C10_N_btm.n2249 C10_N_btm.t54 1.67819
R39691 C10_N_btm.n2246 C10_N_btm.t306 1.67819
R39692 C10_N_btm.n2243 C10_N_btm.t49 1.67819
R39693 C10_N_btm.n2240 C10_N_btm.t856 1.67819
R39694 C10_N_btm.n2237 C10_N_btm.t141 1.67819
R39695 C10_N_btm.n2234 C10_N_btm.t910 1.67819
R39696 C10_N_btm.n2231 C10_N_btm.t191 1.67819
R39697 C10_N_btm.n2228 C10_N_btm.t1028 1.67819
R39698 C10_N_btm.n2225 C10_N_btm.t722 1.67819
R39699 C10_N_btm.n2222 C10_N_btm.t221 1.67819
R39700 C10_N_btm.n2219 C10_N_btm.t841 1.67819
R39701 C10_N_btm.n2216 C10_N_btm.t603 1.67819
R39702 C10_N_btm.n2213 C10_N_btm.t890 1.67819
R39703 C10_N_btm.n2210 C10_N_btm.t664 1.67819
R39704 C10_N_btm.n2207 C10_N_btm.t1009 1.67819
R39705 C10_N_btm.n2204 C10_N_btm.t707 1.67819
R39706 C10_N_btm.n2201 C10_N_btm.t495 1.67819
R39707 C10_N_btm.n2198 C10_N_btm.t822 1.67819
R39708 C10_N_btm.n2195 C10_N_btm.t528 1.67819
R39709 C10_N_btm.n2192 C10_N_btm.t312 1.67819
R39710 C10_N_btm.n2189 C10_N_btm.t772 1.67819
R39711 C10_N_btm.n2186 C10_N_btm.t271 1.67819
R39712 C10_N_btm.n2183 C10_N_btm.t198 1.67819
R39713 C10_N_btm.n2180 C10_N_btm.t323 1.67819
R39714 C10_N_btm.n2177 C10_N_btm.t226 1.67819
R39715 C10_N_btm.n2174 C10_N_btm.t183 1.67819
R39716 C10_N_btm.n2171 C10_N_btm.t164 1.67819
R39717 C10_N_btm.n2168 C10_N_btm.t983 1.67819
R39718 C10_N_btm.n2165 C10_N_btm.t209 1.67819
R39719 C10_N_btm.n2162 C10_N_btm.t975 1.67819
R39720 C10_N_btm.n2159 C10_N_btm.t800 1.67819
R39721 C10_N_btm.n2156 C10_N_btm.t100 1.67819
R39722 C10_N_btm.n2529 C10_N_btm.t862 1.67819
R39723 C10_N_btm.n2524 C10_N_btm.t299 1.67819
R39724 C10_N_btm.n2521 C10_N_btm.t571 1.67819
R39725 C10_N_btm.n2518 C10_N_btm.t253 1.67819
R39726 C10_N_btm.n2515 C10_N_btm.t473 1.67819
R39727 C10_N_btm.n2512 C10_N_btm.t701 1.67819
R39728 C10_N_btm.n2509 C10_N_btm.t418 1.67819
R39729 C10_N_btm.n2506 C10_N_btm.t651 1.67819
R39730 C10_N_btm.n2503 C10_N_btm.t882 1.67819
R39731 C10_N_btm.n2500 C10_N_btm.t593 1.67819
R39732 C10_N_btm.n2497 C10_N_btm.t828 1.67819
R39733 C10_N_btm.n2494 C10_N_btm.t518 1.67819
R39734 C10_N_btm.n2491 C10_N_btm.t778 1.67819
R39735 C10_N_btm.n2488 C10_N_btm.t1015 1.67819
R39736 C10_N_btm.n2485 C10_N_btm.t508 1.67819
R39737 C10_N_btm.n2482 C10_N_btm.t190 1.67819
R39738 C10_N_btm.n2479 C10_N_btm.t453 1.67819
R39739 C10_N_btm.n2476 C10_N_btm.t140 1.67819
R39740 C10_N_btm.n2473 C10_N_btm.t351 1.67819
R39741 C10_N_btm.n2470 C10_N_btm.t639 1.67819
R39742 C10_N_btm.n2467 C10_N_btm.t305 1.67819
R39743 C10_N_btm.n2464 C10_N_btm.t521 1.67819
R39744 C10_N_btm.n2461 C10_N_btm.t259 1.67819
R39745 C10_N_btm.n2458 C10_N_btm.t487 1.67819
R39746 C10_N_btm.n2455 C10_N_btm.t704 1.67819
R39747 C10_N_btm.n2452 C10_N_btm.t368 1.67819
R39748 C10_N_btm.n2449 C10_N_btm.t656 1.67819
R39749 C10_N_btm.n2446 C10_N_btm.t885 1.67819
R39750 C10_N_btm.n2443 C10_N_btm.t535 1.67819
R39751 C10_N_btm.n2440 C10_N_btm.t834 1.67819
R39752 C10_N_btm.n2437 C10_N_btm.t612 1.67819
R39753 C10_N_btm.n2434 C10_N_btm.t712 1.67819
R39754 C10_N_btm.n2431 C10_N_btm.t1019 1.67819
R39755 C10_N_btm.n2428 C10_N_btm.t671 1.67819
R39756 C10_N_btm.n2425 C10_N_btm.t901 1.67819
R39757 C10_N_btm.n2422 C10_N_btm.t84 1.67819
R39758 C10_N_btm.n2419 C10_N_btm.t847 1.67819
R39759 C10_N_btm.n2416 C10_N_btm.t38 1.67819
R39760 C10_N_btm.n2413 C10_N_btm.t734 1.67819
R39761 C10_N_btm.n2410 C10_N_btm.t111 1.67819
R39762 C10_N_btm.n2407 C10_N_btm.t197 1.67819
R39763 C10_N_btm.n2404 C10_N_btm.t960 1.67819
R39764 C10_N_btm.n2401 C10_N_btm.t186 1.67819
R39765 C10_N_btm.n2398 C10_N_btm.t399 1.67819
R39766 C10_N_btm.n2395 C10_N_btm.t87 1.67819
R39767 C10_N_btm.n2392 C10_N_btm.t300 1.67819
R39768 C10_N_btm.n2389 C10_N_btm.t572 1.67819
R39769 C10_N_btm.n2386 C10_N_btm.t254 1.67819
R39770 C10_N_btm.n2383 C10_N_btm.t479 1.67819
R39771 C10_N_btm.n2380 C10_N_btm.t199 1.67819
R39772 C10_N_btm.n2377 C10_N_btm.t419 1.67819
R39773 C10_N_btm.n2374 C10_N_btm.t652 1.67819
R39774 C10_N_btm.n2371 C10_N_btm.t362 1.67819
R39775 C10_N_btm.n2368 C10_N_btm.t594 1.67819
R39776 C10_N_btm.n2365 C10_N_btm.t830 1.67819
R39777 C10_N_btm.n2362 C10_N_btm.t519 1.67819
R39778 C10_N_btm.n2359 C10_N_btm.t780 1.67819
R39779 C10_N_btm.n2356 C10_N_btm.t430 1.67819
R39780 C10_N_btm.n2353 C10_N_btm.t668 1.67819
R39781 C10_N_btm.n2350 C10_N_btm.t958 1.67819
R39782 C10_N_btm.n2347 C10_N_btm.t610 1.67819
R39783 C10_N_btm.n2344 C10_N_btm.t846 1.67819
R39784 C10_N_btm.n2341 C10_N_btm.t82 1.67819
R39785 C10_N_btm.n1594 C10_N_btm.t760 1.67819
R39786 C10_N_btm.n1591 C10_N_btm.t482 1.67819
R39787 C10_N_btm.n1588 C10_N_btm.t257 1.67819
R39788 C10_N_btm.n1585 C10_N_btm.t574 1.67819
R39789 C10_N_btm.n1582 C10_N_btm.t302 1.67819
R39790 C10_N_btm.n1579 C10_N_btm.t90 1.67819
R39791 C10_N_btm.n1576 C10_N_btm.t400 1.67819
R39792 C10_N_btm.n1573 C10_N_btm.t136 1.67819
R39793 C10_N_btm.n1570 C10_N_btm.t450 1.67819
R39794 C10_N_btm.n1567 C10_N_btm.t598 1.67819
R39795 C10_N_btm.n1512 C10_N_btm.t359 1.67819
R39796 C10_N_btm.n1509 C10_N_btm.t109 1.67819
R39797 C10_N_btm.n1506 C10_N_btm.t315 1.67819
R39798 C10_N_btm.n1503 C10_N_btm.t903 1.67819
R39799 C10_N_btm.n1500 C10_N_btm.t225 1.67819
R39800 C10_N_btm.n1497 C10_N_btm.t501 1.67819
R39801 C10_N_btm.n1494 C10_N_btm.t169 1.67819
R39802 C10_N_btm.n1491 C10_N_btm.t381 1.67819
R39803 C10_N_btm.n1488 C10_N_btm.t667 1.67819
R39804 C10_N_btm.n1482 C10_N_btm.t1035 1.67819
R39805 C10_N_btm.n1480 C10_N_btm.t739 1.67819
R39806 C10_N_btm.n1477 C10_N_btm.t505 1.67819
R39807 C10_N_btm.n1474 C10_N_btm.t850 1.67819
R39808 C10_N_btm.n1471 C10_N_btm.t554 1.67819
R39809 C10_N_btm.n1468 C10_N_btm.t337 1.67819
R39810 C10_N_btm.n1465 C10_N_btm.t673 1.67819
R39811 C10_N_btm.n1462 C10_N_btm.t1043 1.67819
R39812 C10_N_btm.n1459 C10_N_btm.t714 1.67819
R39813 C10_N_btm.n1453 C10_N_btm.t624 1.67819
R39814 C10_N_btm.n1395 C10_N_btm.t289 1.67819
R39815 C10_N_btm.n1398 C10_N_btm.t567 1.67819
R39816 C10_N_btm.n1401 C10_N_btm.t247 1.67819
R39817 C10_N_btm.n1404 C10_N_btm.t462 1.67819
R39818 C10_N_btm.n1407 C10_N_btm.t752 1.67819
R39819 C10_N_btm.n1410 C10_N_btm.t407 1.67819
R39820 C10_N_btm.n1413 C10_N_btm.t645 1.67819
R39821 C10_N_btm.n1416 C10_N_btm.t934 1.67819
R39822 C10_N_btm.n1423 C10_N_btm.t864 1.67819
R39823 C10_N_btm.n1426 C10_N_btm.t565 1.67819
R39824 C10_N_btm.n1429 C10_N_btm.t343 1.67819
R39825 C10_N_btm.n1432 C10_N_btm.t683 1.67819
R39826 C10_N_btm.n1435 C10_N_btm.t393 1.67819
R39827 C10_N_btm.n1438 C10_N_btm.t181 1.67819
R39828 C10_N_btm.n1441 C10_N_btm.t502 1.67819
R39829 C10_N_btm.n1444 C10_N_btm.t496 1.67819
R39830 C10_N_btm.n1447 C10_N_btm.t549 1.67819
R39831 C10_N_btm.n1357 C10_N_btm.t456 1.67819
R39832 C10_N_btm.n1360 C10_N_btm.t144 1.67819
R39833 C10_N_btm.n1363 C10_N_btm.t403 1.67819
R39834 C10_N_btm.n1366 C10_N_btm.t97 1.67819
R39835 C10_N_btm.n1369 C10_N_btm.t307 1.67819
R39836 C10_N_btm.n1372 C10_N_btm.t578 1.67819
R39837 C10_N_btm.n1375 C10_N_btm.t260 1.67819
R39838 C10_N_btm.n1378 C10_N_btm.t489 1.67819
R39839 C10_N_btm.n1381 C10_N_btm.t764 1.67819
R39840 C10_N_btm.n635 C10_N_btm.t670 1.67819
R39841 C10_N_btm.n633 C10_N_btm.t383 1.67819
R39842 C10_N_btm.n630 C10_N_btm.t173 1.67819
R39843 C10_N_btm.n627 C10_N_btm.t595 1.67819
R39844 C10_N_btm.n624 C10_N_btm.t232 1.67819
R39845 C10_N_btm.n621 C10_N_btm.t759 1.67819
R39846 C10_N_btm.n618 C10_N_btm.t317 1.67819
R39847 C10_N_btm.n615 C10_N_btm.t237 1.67819
R39848 C10_N_btm.n1351 C10_N_btm.t366 1.67819
R39849 C10_N_btm.n1345 C10_N_btm.t721 1.67819
R39850 C10_N_btm.n1342 C10_N_btm.t1049 1.67819
R39851 C10_N_btm.n1339 C10_N_btm.t675 1.67819
R39852 C10_N_btm.n1336 C10_N_btm.t338 1.67819
R39853 C10_N_btm.n1333 C10_N_btm.t559 1.67819
R39854 C10_N_btm.n1330 C10_N_btm.t855 1.67819
R39855 C10_N_btm.n1327 C10_N_btm.t509 1.67819
R39856 C10_N_btm.n1324 C10_N_btm.t743 1.67819
R39857 C10_N_btm.n1321 C10_N_btm.t51 1.67819
R39858 C10_N_btm.n1314 C10_N_btm.t938 1.67819
R39859 C10_N_btm.n1311 C10_N_btm.t649 1.67819
R39860 C10_N_btm.n1308 C10_N_btm.t413 1.67819
R39861 C10_N_btm.n1305 C10_N_btm.t755 1.67819
R39862 C10_N_btm.n1302 C10_N_btm.t470 1.67819
R39863 C10_N_btm.n1299 C10_N_btm.t250 1.67819
R39864 C10_N_btm.n1296 C10_N_btm.t568 1.67819
R39865 C10_N_btm.n1293 C10_N_btm.t296 1.67819
R39866 C10_N_btm.n1290 C10_N_btm.t629 1.67819
R39867 C10_N_btm.n1284 C10_N_btm.t999 1.67819
R39868 C10_N_btm.n668 C10_N_btm.t657 1.67819
R39869 C10_N_btm.n671 C10_N_btm.t944 1.67819
R39870 C10_N_btm.n674 C10_N_btm.t596 1.67819
R39871 C10_N_btm.n677 C10_N_btm.t835 1.67819
R39872 C10_N_btm.n680 C10_N_btm.t69 1.67819
R39873 C10_N_btm.n683 C10_N_btm.t782 1.67819
R39874 C10_N_btm.n686 C10_N_btm.t1020 1.67819
R39875 C10_N_btm.n688 C10_N_btm.t520 1.67819
R39876 C10_N_btm.n1254 C10_N_btm.t152 1.67819
R39877 C10_N_btm.n1257 C10_N_btm.t917 1.67819
R39878 C10_N_btm.n1260 C10_N_btm.t682 1.67819
R39879 C10_N_btm.n1263 C10_N_btm.t55 1.67819
R39880 C10_N_btm.n1266 C10_N_btm.t733 1.67819
R39881 C10_N_btm.n1269 C10_N_btm.t1030 1.67819
R39882 C10_N_btm.n1272 C10_N_btm.t845 1.67819
R39883 C10_N_btm.n1275 C10_N_btm.t548 1.67819
R39884 C10_N_btm.n1278 C10_N_btm.t899 1.67819
R39885 C10_N_btm.n1223 C10_N_btm.t801 1.67819
R39886 C10_N_btm.n1226 C10_N_btm.t455 1.67819
R39887 C10_N_btm.n1229 C10_N_btm.t745 1.67819
R39888 C10_N_btm.n1232 C10_N_btm.t402 1.67819
R39889 C10_N_btm.n1235 C10_N_btm.t640 1.67819
R39890 C10_N_btm.n1238 C10_N_btm.t929 1.67819
R39891 C10_N_btm.n1241 C10_N_btm.t577 1.67819
R39892 C10_N_btm.n1244 C10_N_btm.t816 1.67819
R39893 C10_N_btm.n1247 C10_N_btm.t1033 1.67819
R39894 C10_N_btm.n741 C10_N_btm.t391 1.67819
R39895 C10_N_btm.n739 C10_N_btm.t129 1.67819
R39896 C10_N_btm.n736 C10_N_btm.t952 1.67819
R39897 C10_N_btm.n733 C10_N_btm.t484 1.67819
R39898 C10_N_btm.n730 C10_N_btm.t1021 1.67819
R39899 C10_N_btm.n727 C10_N_btm.t771 1.67819
R39900 C10_N_btm.n724 C10_N_btm.t62 1.67819
R39901 C10_N_btm.n721 C10_N_btm.t824 1.67819
R39902 C10_N_btm.n1217 C10_N_btm.t475 1.67819
R39903 C10_N_btm.n1211 C10_N_btm.t110 1.67819
R39904 C10_N_btm.n1208 C10_N_btm.t720 1.67819
R39905 C10_N_btm.n1205 C10_N_btm.t1024 1.67819
R39906 C10_N_btm.n1202 C10_N_btm.t674 1.67819
R39907 C10_N_btm.n1199 C10_N_btm.t909 1.67819
R39908 C10_N_btm.n1196 C10_N_btm.t138 1.67819
R39909 C10_N_btm.n1193 C10_N_btm.t854 1.67819
R39910 C10_N_btm.n1190 C10_N_btm.t45 1.67819
R39911 C10_N_btm.n1187 C10_N_btm.t304 1.67819
R39912 C10_N_btm.n1180 C10_N_btm.t663 1.67819
R39913 C10_N_btm.n1177 C10_N_btm.t376 1.67819
R39914 C10_N_btm.n1174 C10_N_btm.t165 1.67819
R39915 C10_N_btm.n1171 C10_N_btm.t494 1.67819
R39916 C10_N_btm.n1168 C10_N_btm.t210 1.67819
R39917 C10_N_btm.n1165 C10_N_btm.t941 1.67819
R39918 C10_N_btm.n1162 C10_N_btm.t310 1.67819
R39919 C10_N_btm.n1159 C10_N_btm.t85 1.67819
R39920 C10_N_btm.n1156 C10_N_btm.t356 1.67819
R39921 C10_N_btm.n1150 C10_N_btm.t270 1.67819
R39922 C10_N_btm.n774 C10_N_btm.t998 1.67819
R39923 C10_N_btm.n777 C10_N_btm.t240 1.67819
R39924 C10_N_btm.n780 C10_N_btm.t943 1.67819
R39925 C10_N_btm.n783 C10_N_btm.t120 1.67819
R39926 C10_N_btm.n786 C10_N_btm.t1045 1.67819
R39927 C10_N_btm.n789 C10_N_btm.t68 1.67819
R39928 C10_N_btm.n792 C10_N_btm.t283 1.67819
R39929 C10_N_btm.n794 C10_N_btm.t557 1.67819
R39930 C10_N_btm.n1120 C10_N_btm.t466 1.67819
R39931 C10_N_btm.n1123 C10_N_btm.t195 1.67819
R39932 C10_N_btm.n1126 C10_N_btm.t47 1.67819
R39933 C10_N_btm.n1129 C10_N_btm.t291 1.67819
R39934 C10_N_btm.n1132 C10_N_btm.t35 1.67819
R39935 C10_N_btm.n1135 C10_N_btm.t844 1.67819
R39936 C10_N_btm.n1138 C10_N_btm.t131 1.67819
R39937 C10_N_btm.n1141 C10_N_btm.t898 1.67819
R39938 C10_N_btm.n1144 C10_N_btm.t91 1.67819
R39939 C10_N_btm.n1089 C10_N_btm.t1056 1.67819
R39940 C10_N_btm.n1092 C10_N_btm.t202 1.67819
R39941 C10_N_btm.n1095 C10_N_btm.t483 1.67819
R39942 C10_N_btm.n1098 C10_N_btm.t159 1.67819
R39943 C10_N_btm.n1101 C10_N_btm.t367 1.67819
R39944 C10_N_btm.n1104 C10_N_btm.t654 1.67819
R39945 C10_N_btm.n1107 C10_N_btm.t318 1.67819
R39946 C10_N_btm.n1110 C10_N_btm.t534 1.67819
R39947 C10_N_btm.n1113 C10_N_btm.t832 1.67819
R39948 C10_N_btm.n847 C10_N_btm.t729 1.67819
R39949 C10_N_btm.n845 C10_N_btm.t442 1.67819
R39950 C10_N_btm.n842 C10_N_btm.t481 1.67819
R39951 C10_N_btm.n839 C10_N_btm.t544 1.67819
R39952 C10_N_btm.n836 C10_N_btm.t278 1.67819
R39953 C10_N_btm.n833 C10_N_btm.t60 1.67819
R39954 C10_N_btm.n830 C10_N_btm.t380 1.67819
R39955 C10_N_btm.n827 C10_N_btm.t468 1.67819
R39956 C10_N_btm.n1083 C10_N_btm.t429 1.67819
R39957 C10_N_btm.n1077 C10_N_btm.t794 1.67819
R39958 C10_N_btm.n1074 C10_N_btm.t447 1.67819
R39959 C10_N_btm.n1071 C10_N_btm.t740 1.67819
R39960 C10_N_btm.n1068 C10_N_btm.t398 1.67819
R39961 C10_N_btm.n1065 C10_N_btm.t630 1.67819
R39962 C10_N_btm.n1062 C10_N_btm.t921 1.67819
R39963 C10_N_btm.n1059 C10_N_btm.t569 1.67819
R39964 C10_N_btm.n1056 C10_N_btm.t810 1.67819
R39965 C10_N_btm.n1053 C10_N_btm.t213 1.67819
R39966 C10_N_btm.n1046 C10_N_btm.t1007 1.67819
R39967 C10_N_btm.n1043 C10_N_btm.t706 1.67819
R39968 C10_N_btm.n1040 C10_N_btm.t490 1.67819
R39969 C10_N_btm.n1037 C10_N_btm.t820 1.67819
R39970 C10_N_btm.n1034 C10_N_btm.t527 1.67819
R39971 C10_N_btm.n1031 C10_N_btm.t309 1.67819
R39972 C10_N_btm.n1028 C10_N_btm.t646 1.67819
R39973 C10_N_btm.n1025 C10_N_btm.t355 1.67819
R39974 C10_N_btm.n1022 C10_N_btm.t695 1.67819
R39975 C10_N_btm.n1016 C10_N_btm.t600 1.67819
R39976 C10_N_btm.n880 C10_N_btm.t269 1.67819
R39977 C10_N_btm.n883 C10_N_btm.t538 1.67819
R39978 C10_N_btm.n886 C10_N_btm.t235 1.67819
R39979 C10_N_btm.n889 C10_N_btm.t437 1.67819
R39980 C10_N_btm.n892 C10_N_btm.t716 1.67819
R39981 C10_N_btm.n895 C10_N_btm.t386 1.67819
R39982 C10_N_btm.n898 C10_N_btm.t615 1.67819
R39983 C10_N_btm.n900 C10_N_btm.t448 1.67819
R39984 C10_N_btm.n986 C10_N_btm.t208 1.67819
R39985 C10_N_btm.n989 C10_N_btm.t984 1.67819
R39986 C10_N_btm.n992 C10_N_btm.t746 1.67819
R39987 C10_N_btm.n995 C10_N_btm.t53 1.67819
R39988 C10_N_btm.n998 C10_N_btm.t802 1.67819
R39989 C10_N_btm.n1001 C10_N_btm.t562 1.67819
R39990 C10_N_btm.n1004 C10_N_btm.t915 1.67819
R39991 C10_N_btm.n1007 C10_N_btm.t621 1.67819
R39992 C10_N_btm.n1010 C10_N_btm.t966 1.67819
R39993 C10_N_btm.n955 C10_N_btm.t871 1.67819
R39994 C10_N_btm.n958 C10_N_btm.t1054 1.67819
R39995 C10_N_btm.n961 C10_N_btm.t814 1.67819
R39996 C10_N_btm.n964 C10_N_btm.t480 1.67819
R39997 C10_N_btm.n967 C10_N_btm.t702 1.67819
R39998 C10_N_btm.n970 C10_N_btm.t995 1.67819
R39999 C10_N_btm.n973 C10_N_btm.t653 1.67819
R40000 C10_N_btm.n976 C10_N_btm.t883 1.67819
R40001 C10_N_btm.n979 C10_N_btm.t599 1.67819
R40002 C10_N_btm.n923 C10_N_btm.t451 1.67819
R40003 C10_N_btm.n926 C10_N_btm.t189 1.67819
R40004 C10_N_btm.n929 C10_N_btm.t1025 1.67819
R40005 C10_N_btm.n932 C10_N_btm.t285 1.67819
R40006 C10_N_btm.n935 C10_N_btm.t118 1.67819
R40007 C10_N_btm.n938 C10_N_btm.t840 1.67819
R40008 C10_N_btm.n941 C10_N_btm.t123 1.67819
R40009 C10_N_btm.n944 C10_N_btm.t889 1.67819
R40010 C10_N_btm.n949 C10_N_btm.t178 1.67819
R40011 C10_N_btm.n1564 C10_N_btm.t94 1.67819
R40012 C10_N_btm.n1561 C10_N_btm.t284 1.67819
R40013 C10_N_btm.n1558 C10_N_btm.t71 1.67819
R40014 C10_N_btm.n1555 C10_N_btm.t887 1.67819
R40015 C10_N_btm.n1552 C10_N_btm.t122 1.67819
R40016 C10_N_btm.n1549 C10_N_btm.t945 1.67819
R40017 C10_N_btm.n1546 C10_N_btm.t246 1.67819
R40018 C10_N_btm.n1543 C10_N_btm.t1000 1.67819
R40019 C10_N_btm.n1540 C10_N_btm.t765 1.67819
R40020 C10_N_btm.n1537 C10_N_btm.t58 1.67819
R40021 C10_N_btm.n1534 C10_N_btm.t873 1.67819
R40022 C10_N_btm.n1531 C10_N_btm.t580 1.67819
R40023 C10_N_btm.n507 C10_N_btm.n506 1.05569
R40024 C10_N_btm.n2339 C10_N_btm.n1969 1.05569
R40025 C10_N_btm.n2527 C10_N_btm.n2526 1.05569
R40026 C10_N_btm.n1529 C10_N_btm.n524 1.05569
R40027 C10_N_btm.n44 C10_N_btm.n42 1.0005
R40028 C10_N_btm.n45 C10_N_btm.n41 1.0005
R40029 C10_N_btm.n46 C10_N_btm.n40 1.0005
R40030 C10_N_btm.n47 C10_N_btm.n39 1.0005
R40031 C10_N_btm.n48 C10_N_btm.n38 1.0005
R40032 C10_N_btm.n49 C10_N_btm.n37 1.0005
R40033 C10_N_btm.n50 C10_N_btm.n36 1.0005
R40034 C10_N_btm.n51 C10_N_btm.n35 1.0005
R40035 C10_N_btm.n3835 C10_N_btm.n34 1.0005
R40036 C10_N_btm.n3835 C10_N_btm.n3834 1.0005
R40037 C10_N_btm.n54 C10_N_btm.n51 1.0005
R40038 C10_N_btm.n55 C10_N_btm.n50 1.0005
R40039 C10_N_btm.n56 C10_N_btm.n49 1.0005
R40040 C10_N_btm.n57 C10_N_btm.n48 1.0005
R40041 C10_N_btm.n58 C10_N_btm.n47 1.0005
R40042 C10_N_btm.n59 C10_N_btm.n46 1.0005
R40043 C10_N_btm.n60 C10_N_btm.n45 1.0005
R40044 C10_N_btm.n3806 C10_N_btm.n44 1.0005
R40045 C10_N_btm.n3806 C10_N_btm.n3805 1.0005
R40046 C10_N_btm.n3743 C10_N_btm.n60 1.0005
R40047 C10_N_btm.n3742 C10_N_btm.n59 1.0005
R40048 C10_N_btm.n3741 C10_N_btm.n58 1.0005
R40049 C10_N_btm.n3740 C10_N_btm.n57 1.0005
R40050 C10_N_btm.n3739 C10_N_btm.n56 1.0005
R40051 C10_N_btm.n3738 C10_N_btm.n55 1.0005
R40052 C10_N_btm.n3737 C10_N_btm.n54 1.0005
R40053 C10_N_btm.n3834 C10_N_btm.n52 1.0005
R40054 C10_N_btm.n71 C10_N_btm.n52 1.0005
R40055 C10_N_btm.n3737 C10_N_btm.n70 1.0005
R40056 C10_N_btm.n3738 C10_N_btm.n69 1.0005
R40057 C10_N_btm.n3739 C10_N_btm.n68 1.0005
R40058 C10_N_btm.n3740 C10_N_btm.n67 1.0005
R40059 C10_N_btm.n3741 C10_N_btm.n66 1.0005
R40060 C10_N_btm.n3742 C10_N_btm.n65 1.0005
R40061 C10_N_btm.n3743 C10_N_btm.n64 1.0005
R40062 C10_N_btm.n3805 C10_N_btm.n61 1.0005
R40063 C10_N_btm.n3704 C10_N_btm.n61 1.0005
R40064 C10_N_btm.n80 C10_N_btm.n64 1.0005
R40065 C10_N_btm.n79 C10_N_btm.n65 1.0005
R40066 C10_N_btm.n78 C10_N_btm.n66 1.0005
R40067 C10_N_btm.n77 C10_N_btm.n67 1.0005
R40068 C10_N_btm.n76 C10_N_btm.n68 1.0005
R40069 C10_N_btm.n75 C10_N_btm.n69 1.0005
R40070 C10_N_btm.n74 C10_N_btm.n70 1.0005
R40071 C10_N_btm.n73 C10_N_btm.n71 1.0005
R40072 C10_N_btm.n123 C10_N_btm.n73 1.0005
R40073 C10_N_btm.n93 C10_N_btm.n74 1.0005
R40074 C10_N_btm.n94 C10_N_btm.n75 1.0005
R40075 C10_N_btm.n95 C10_N_btm.n76 1.0005
R40076 C10_N_btm.n96 C10_N_btm.n77 1.0005
R40077 C10_N_btm.n97 C10_N_btm.n78 1.0005
R40078 C10_N_btm.n98 C10_N_btm.n79 1.0005
R40079 C10_N_btm.n99 C10_N_btm.n80 1.0005
R40080 C10_N_btm.n3704 C10_N_btm.n3703 1.0005
R40081 C10_N_btm.n3703 C10_N_btm.n81 1.0005
R40082 C10_N_btm.n99 C10_N_btm.n84 1.0005
R40083 C10_N_btm.n98 C10_N_btm.n85 1.0005
R40084 C10_N_btm.n97 C10_N_btm.n86 1.0005
R40085 C10_N_btm.n96 C10_N_btm.n87 1.0005
R40086 C10_N_btm.n95 C10_N_btm.n88 1.0005
R40087 C10_N_btm.n94 C10_N_btm.n89 1.0005
R40088 C10_N_btm.n93 C10_N_btm.n90 1.0005
R40089 C10_N_btm.n124 C10_N_btm.n123 1.0005
R40090 C10_N_btm.n126 C10_N_btm.n124 1.0005
R40091 C10_N_btm.n127 C10_N_btm.n90 1.0005
R40092 C10_N_btm.n128 C10_N_btm.n89 1.0005
R40093 C10_N_btm.n129 C10_N_btm.n88 1.0005
R40094 C10_N_btm.n130 C10_N_btm.n87 1.0005
R40095 C10_N_btm.n131 C10_N_btm.n86 1.0005
R40096 C10_N_btm.n132 C10_N_btm.n85 1.0005
R40097 C10_N_btm.n133 C10_N_btm.n84 1.0005
R40098 C10_N_btm.n3637 C10_N_btm.n81 1.0005
R40099 C10_N_btm.n3637 C10_N_btm.n3636 1.0005
R40100 C10_N_btm.n152 C10_N_btm.n133 1.0005
R40101 C10_N_btm.n151 C10_N_btm.n132 1.0005
R40102 C10_N_btm.n150 C10_N_btm.n131 1.0005
R40103 C10_N_btm.n149 C10_N_btm.n130 1.0005
R40104 C10_N_btm.n148 C10_N_btm.n129 1.0005
R40105 C10_N_btm.n147 C10_N_btm.n128 1.0005
R40106 C10_N_btm.n146 C10_N_btm.n127 1.0005
R40107 C10_N_btm.n176 C10_N_btm.n126 1.0005
R40108 C10_N_btm.n177 C10_N_btm.n176 1.0005
R40109 C10_N_btm.n146 C10_N_btm.n143 1.0005
R40110 C10_N_btm.n147 C10_N_btm.n142 1.0005
R40111 C10_N_btm.n148 C10_N_btm.n141 1.0005
R40112 C10_N_btm.n149 C10_N_btm.n140 1.0005
R40113 C10_N_btm.n150 C10_N_btm.n139 1.0005
R40114 C10_N_btm.n151 C10_N_btm.n138 1.0005
R40115 C10_N_btm.n152 C10_N_btm.n137 1.0005
R40116 C10_N_btm.n3636 C10_N_btm.n134 1.0005
R40117 C10_N_btm.n3570 C10_N_btm.n134 1.0005
R40118 C10_N_btm.n186 C10_N_btm.n137 1.0005
R40119 C10_N_btm.n185 C10_N_btm.n138 1.0005
R40120 C10_N_btm.n184 C10_N_btm.n139 1.0005
R40121 C10_N_btm.n183 C10_N_btm.n140 1.0005
R40122 C10_N_btm.n182 C10_N_btm.n141 1.0005
R40123 C10_N_btm.n181 C10_N_btm.n142 1.0005
R40124 C10_N_btm.n180 C10_N_btm.n143 1.0005
R40125 C10_N_btm.n179 C10_N_btm.n177 1.0005
R40126 C10_N_btm.n229 C10_N_btm.n179 1.0005
R40127 C10_N_btm.n199 C10_N_btm.n180 1.0005
R40128 C10_N_btm.n200 C10_N_btm.n181 1.0005
R40129 C10_N_btm.n201 C10_N_btm.n182 1.0005
R40130 C10_N_btm.n202 C10_N_btm.n183 1.0005
R40131 C10_N_btm.n203 C10_N_btm.n184 1.0005
R40132 C10_N_btm.n204 C10_N_btm.n185 1.0005
R40133 C10_N_btm.n205 C10_N_btm.n186 1.0005
R40134 C10_N_btm.n3570 C10_N_btm.n3569 1.0005
R40135 C10_N_btm.n3569 C10_N_btm.n187 1.0005
R40136 C10_N_btm.n205 C10_N_btm.n190 1.0005
R40137 C10_N_btm.n204 C10_N_btm.n191 1.0005
R40138 C10_N_btm.n203 C10_N_btm.n192 1.0005
R40139 C10_N_btm.n202 C10_N_btm.n193 1.0005
R40140 C10_N_btm.n201 C10_N_btm.n194 1.0005
R40141 C10_N_btm.n200 C10_N_btm.n195 1.0005
R40142 C10_N_btm.n199 C10_N_btm.n196 1.0005
R40143 C10_N_btm.n230 C10_N_btm.n229 1.0005
R40144 C10_N_btm.n232 C10_N_btm.n230 1.0005
R40145 C10_N_btm.n233 C10_N_btm.n196 1.0005
R40146 C10_N_btm.n234 C10_N_btm.n195 1.0005
R40147 C10_N_btm.n235 C10_N_btm.n194 1.0005
R40148 C10_N_btm.n236 C10_N_btm.n193 1.0005
R40149 C10_N_btm.n237 C10_N_btm.n192 1.0005
R40150 C10_N_btm.n238 C10_N_btm.n191 1.0005
R40151 C10_N_btm.n239 C10_N_btm.n190 1.0005
R40152 C10_N_btm.n3503 C10_N_btm.n187 1.0005
R40153 C10_N_btm.n3503 C10_N_btm.n3502 1.0005
R40154 C10_N_btm.n258 C10_N_btm.n239 1.0005
R40155 C10_N_btm.n257 C10_N_btm.n238 1.0005
R40156 C10_N_btm.n256 C10_N_btm.n237 1.0005
R40157 C10_N_btm.n255 C10_N_btm.n236 1.0005
R40158 C10_N_btm.n254 C10_N_btm.n235 1.0005
R40159 C10_N_btm.n253 C10_N_btm.n234 1.0005
R40160 C10_N_btm.n252 C10_N_btm.n233 1.0005
R40161 C10_N_btm.n282 C10_N_btm.n232 1.0005
R40162 C10_N_btm.n283 C10_N_btm.n282 1.0005
R40163 C10_N_btm.n252 C10_N_btm.n249 1.0005
R40164 C10_N_btm.n253 C10_N_btm.n248 1.0005
R40165 C10_N_btm.n254 C10_N_btm.n247 1.0005
R40166 C10_N_btm.n255 C10_N_btm.n246 1.0005
R40167 C10_N_btm.n256 C10_N_btm.n245 1.0005
R40168 C10_N_btm.n257 C10_N_btm.n244 1.0005
R40169 C10_N_btm.n258 C10_N_btm.n243 1.0005
R40170 C10_N_btm.n3502 C10_N_btm.n240 1.0005
R40171 C10_N_btm.n3436 C10_N_btm.n240 1.0005
R40172 C10_N_btm.n292 C10_N_btm.n243 1.0005
R40173 C10_N_btm.n291 C10_N_btm.n244 1.0005
R40174 C10_N_btm.n290 C10_N_btm.n245 1.0005
R40175 C10_N_btm.n289 C10_N_btm.n246 1.0005
R40176 C10_N_btm.n288 C10_N_btm.n247 1.0005
R40177 C10_N_btm.n287 C10_N_btm.n248 1.0005
R40178 C10_N_btm.n286 C10_N_btm.n249 1.0005
R40179 C10_N_btm.n285 C10_N_btm.n283 1.0005
R40180 C10_N_btm.n335 C10_N_btm.n285 1.0005
R40181 C10_N_btm.n305 C10_N_btm.n286 1.0005
R40182 C10_N_btm.n306 C10_N_btm.n287 1.0005
R40183 C10_N_btm.n307 C10_N_btm.n288 1.0005
R40184 C10_N_btm.n308 C10_N_btm.n289 1.0005
R40185 C10_N_btm.n309 C10_N_btm.n290 1.0005
R40186 C10_N_btm.n310 C10_N_btm.n291 1.0005
R40187 C10_N_btm.n311 C10_N_btm.n292 1.0005
R40188 C10_N_btm.n3436 C10_N_btm.n3435 1.0005
R40189 C10_N_btm.n3435 C10_N_btm.n293 1.0005
R40190 C10_N_btm.n311 C10_N_btm.n296 1.0005
R40191 C10_N_btm.n310 C10_N_btm.n297 1.0005
R40192 C10_N_btm.n309 C10_N_btm.n298 1.0005
R40193 C10_N_btm.n308 C10_N_btm.n299 1.0005
R40194 C10_N_btm.n307 C10_N_btm.n300 1.0005
R40195 C10_N_btm.n306 C10_N_btm.n301 1.0005
R40196 C10_N_btm.n305 C10_N_btm.n302 1.0005
R40197 C10_N_btm.n336 C10_N_btm.n335 1.0005
R40198 C10_N_btm.n338 C10_N_btm.n336 1.0005
R40199 C10_N_btm.n339 C10_N_btm.n302 1.0005
R40200 C10_N_btm.n340 C10_N_btm.n301 1.0005
R40201 C10_N_btm.n341 C10_N_btm.n300 1.0005
R40202 C10_N_btm.n342 C10_N_btm.n299 1.0005
R40203 C10_N_btm.n343 C10_N_btm.n298 1.0005
R40204 C10_N_btm.n344 C10_N_btm.n297 1.0005
R40205 C10_N_btm.n345 C10_N_btm.n296 1.0005
R40206 C10_N_btm.n3369 C10_N_btm.n293 1.0005
R40207 C10_N_btm.n3369 C10_N_btm.n3368 1.0005
R40208 C10_N_btm.n364 C10_N_btm.n345 1.0005
R40209 C10_N_btm.n363 C10_N_btm.n344 1.0005
R40210 C10_N_btm.n362 C10_N_btm.n343 1.0005
R40211 C10_N_btm.n361 C10_N_btm.n342 1.0005
R40212 C10_N_btm.n360 C10_N_btm.n341 1.0005
R40213 C10_N_btm.n359 C10_N_btm.n340 1.0005
R40214 C10_N_btm.n358 C10_N_btm.n339 1.0005
R40215 C10_N_btm.n388 C10_N_btm.n338 1.0005
R40216 C10_N_btm.n389 C10_N_btm.n388 1.0005
R40217 C10_N_btm.n358 C10_N_btm.n355 1.0005
R40218 C10_N_btm.n359 C10_N_btm.n354 1.0005
R40219 C10_N_btm.n360 C10_N_btm.n353 1.0005
R40220 C10_N_btm.n361 C10_N_btm.n352 1.0005
R40221 C10_N_btm.n362 C10_N_btm.n351 1.0005
R40222 C10_N_btm.n363 C10_N_btm.n350 1.0005
R40223 C10_N_btm.n364 C10_N_btm.n349 1.0005
R40224 C10_N_btm.n3368 C10_N_btm.n346 1.0005
R40225 C10_N_btm.n3302 C10_N_btm.n346 1.0005
R40226 C10_N_btm.n398 C10_N_btm.n349 1.0005
R40227 C10_N_btm.n397 C10_N_btm.n350 1.0005
R40228 C10_N_btm.n396 C10_N_btm.n351 1.0005
R40229 C10_N_btm.n395 C10_N_btm.n352 1.0005
R40230 C10_N_btm.n394 C10_N_btm.n353 1.0005
R40231 C10_N_btm.n393 C10_N_btm.n354 1.0005
R40232 C10_N_btm.n392 C10_N_btm.n355 1.0005
R40233 C10_N_btm.n391 C10_N_btm.n389 1.0005
R40234 C10_N_btm.n435 C10_N_btm.n391 1.0005
R40235 C10_N_btm.n436 C10_N_btm.n392 1.0005
R40236 C10_N_btm.n437 C10_N_btm.n393 1.0005
R40237 C10_N_btm.n438 C10_N_btm.n394 1.0005
R40238 C10_N_btm.n439 C10_N_btm.n395 1.0005
R40239 C10_N_btm.n440 C10_N_btm.n396 1.0005
R40240 C10_N_btm.n441 C10_N_btm.n397 1.0005
R40241 C10_N_btm.n442 C10_N_btm.n398 1.0005
R40242 C10_N_btm.n3302 C10_N_btm.n3301 1.0005
R40243 C10_N_btm.n3301 C10_N_btm.n399 1.0005
R40244 C10_N_btm.n442 C10_N_btm.n402 1.0005
R40245 C10_N_btm.n441 C10_N_btm.n403 1.0005
R40246 C10_N_btm.n440 C10_N_btm.n404 1.0005
R40247 C10_N_btm.n439 C10_N_btm.n405 1.0005
R40248 C10_N_btm.n438 C10_N_btm.n406 1.0005
R40249 C10_N_btm.n437 C10_N_btm.n407 1.0005
R40250 C10_N_btm.n436 C10_N_btm.n408 1.0005
R40251 C10_N_btm.n435 C10_N_btm.n409 1.0005
R40252 C10_N_btm.n410 C10_N_btm.n390 1.0005
R40253 C10_N_btm.n423 C10_N_btm.n422 1.0005
R40254 C10_N_btm.n424 C10_N_btm.n421 1.0005
R40255 C10_N_btm.n425 C10_N_btm.n420 1.0005
R40256 C10_N_btm.n426 C10_N_btm.n419 1.0005
R40257 C10_N_btm.n427 C10_N_btm.n418 1.0005
R40258 C10_N_btm.n428 C10_N_btm.n417 1.0005
R40259 C10_N_btm.n429 C10_N_btm.n416 1.0005
R40260 C10_N_btm.n430 C10_N_btm.n415 1.0005
R40261 C10_N_btm.n431 C10_N_btm.n414 1.0005
R40262 C10_N_btm.n432 C10_N_btm.n413 1.0005
R40263 C10_N_btm.n433 C10_N_btm.n412 1.0005
R40264 C10_N_btm.n434 C10_N_btm.n411 1.0005
R40265 C10_N_btm.n1599 C10_N_btm.n546 1.0005
R40266 C10_N_btm.n1600 C10_N_btm.n545 1.0005
R40267 C10_N_btm.n1601 C10_N_btm.n544 1.0005
R40268 C10_N_btm.n1602 C10_N_btm.n543 1.0005
R40269 C10_N_btm.n1603 C10_N_btm.n542 1.0005
R40270 C10_N_btm.n1604 C10_N_btm.n541 1.0005
R40271 C10_N_btm.n1605 C10_N_btm.n540 1.0005
R40272 C10_N_btm.n1606 C10_N_btm.n539 1.0005
R40273 C10_N_btm.n1607 C10_N_btm.n538 1.0005
R40274 C10_N_btm.n1608 C10_N_btm.n537 1.0005
R40275 C10_N_btm.n1609 C10_N_btm.n536 1.0005
R40276 C10_N_btm.n1610 C10_N_btm.n535 1.0005
R40277 C10_N_btm.n1611 C10_N_btm.n534 1.0005
R40278 C10_N_btm.n1612 C10_N_btm.n533 1.0005
R40279 C10_N_btm.n1613 C10_N_btm.n532 1.0005
R40280 C10_N_btm.n1614 C10_N_btm.n531 1.0005
R40281 C10_N_btm.n1615 C10_N_btm.n530 1.0005
R40282 C10_N_btm.n1616 C10_N_btm.n529 1.0005
R40283 C10_N_btm.n1617 C10_N_btm.n528 1.0005
R40284 C10_N_btm.n1618 C10_N_btm.n527 1.0005
R40285 C10_N_btm.n1619 C10_N_btm.n526 1.0005
R40286 C10_N_btm.n1620 C10_N_btm.n525 1.0005
R40287 C10_N_btm.n1621 C10_N_btm.n524 1.0005
R40288 C10_N_btm.n1622 C10_N_btm.n523 1.0005
R40289 C10_N_btm.n1623 C10_N_btm.n522 1.0005
R40290 C10_N_btm.n1624 C10_N_btm.n521 1.0005
R40291 C10_N_btm.n1625 C10_N_btm.n520 1.0005
R40292 C10_N_btm.n1626 C10_N_btm.n519 1.0005
R40293 C10_N_btm.n1627 C10_N_btm.n518 1.0005
R40294 C10_N_btm.n1628 C10_N_btm.n517 1.0005
R40295 C10_N_btm.n1629 C10_N_btm.n516 1.0005
R40296 C10_N_btm.n1630 C10_N_btm.n515 1.0005
R40297 C10_N_btm.n1631 C10_N_btm.n514 1.0005
R40298 C10_N_btm.n1632 C10_N_btm.n513 1.0005
R40299 C10_N_btm.n1633 C10_N_btm.n512 1.0005
R40300 C10_N_btm.n1634 C10_N_btm.n511 1.0005
R40301 C10_N_btm.n1635 C10_N_btm.n510 1.0005
R40302 C10_N_btm.n1636 C10_N_btm.n509 1.0005
R40303 C10_N_btm.n1637 C10_N_btm.n508 1.0005
R40304 C10_N_btm.n1638 C10_N_btm.n507 1.0005
R40305 C10_N_btm.n1639 C10_N_btm.n422 1.0005
R40306 C10_N_btm.n1640 C10_N_btm.n421 1.0005
R40307 C10_N_btm.n1641 C10_N_btm.n420 1.0005
R40308 C10_N_btm.n1642 C10_N_btm.n419 1.0005
R40309 C10_N_btm.n1643 C10_N_btm.n418 1.0005
R40310 C10_N_btm.n1644 C10_N_btm.n417 1.0005
R40311 C10_N_btm.n1645 C10_N_btm.n416 1.0005
R40312 C10_N_btm.n1646 C10_N_btm.n415 1.0005
R40313 C10_N_btm.n1647 C10_N_btm.n414 1.0005
R40314 C10_N_btm.n1648 C10_N_btm.n413 1.0005
R40315 C10_N_btm.n1649 C10_N_btm.n412 1.0005
R40316 C10_N_btm.n1650 C10_N_btm.n411 1.0005
R40317 C10_N_btm.n1651 C10_N_btm.n410 1.0005
R40318 C10_N_btm.n1652 C10_N_btm.n409 1.0005
R40319 C10_N_btm.n1653 C10_N_btm.n408 1.0005
R40320 C10_N_btm.n1654 C10_N_btm.n407 1.0005
R40321 C10_N_btm.n1655 C10_N_btm.n406 1.0005
R40322 C10_N_btm.n1656 C10_N_btm.n405 1.0005
R40323 C10_N_btm.n1657 C10_N_btm.n404 1.0005
R40324 C10_N_btm.n1658 C10_N_btm.n403 1.0005
R40325 C10_N_btm.n1659 C10_N_btm.n402 1.0005
R40326 C10_N_btm.n2917 C10_N_btm.n399 1.0005
R40327 C10_N_btm.n2917 C10_N_btm.n2916 1.0005
R40328 C10_N_btm.n1784 C10_N_btm.n1659 1.0005
R40329 C10_N_btm.n1783 C10_N_btm.n1658 1.0005
R40330 C10_N_btm.n1782 C10_N_btm.n1657 1.0005
R40331 C10_N_btm.n1781 C10_N_btm.n1656 1.0005
R40332 C10_N_btm.n1780 C10_N_btm.n1655 1.0005
R40333 C10_N_btm.n1779 C10_N_btm.n1654 1.0005
R40334 C10_N_btm.n1778 C10_N_btm.n1653 1.0005
R40335 C10_N_btm.n1777 C10_N_btm.n1652 1.0005
R40336 C10_N_btm.n1776 C10_N_btm.n1651 1.0005
R40337 C10_N_btm.n1775 C10_N_btm.n1650 1.0005
R40338 C10_N_btm.n1774 C10_N_btm.n1649 1.0005
R40339 C10_N_btm.n1773 C10_N_btm.n1648 1.0005
R40340 C10_N_btm.n1772 C10_N_btm.n1647 1.0005
R40341 C10_N_btm.n1771 C10_N_btm.n1646 1.0005
R40342 C10_N_btm.n1770 C10_N_btm.n1645 1.0005
R40343 C10_N_btm.n1769 C10_N_btm.n1644 1.0005
R40344 C10_N_btm.n1768 C10_N_btm.n1643 1.0005
R40345 C10_N_btm.n1767 C10_N_btm.n1642 1.0005
R40346 C10_N_btm.n1766 C10_N_btm.n1641 1.0005
R40347 C10_N_btm.n1765 C10_N_btm.n1640 1.0005
R40348 C10_N_btm.n1764 C10_N_btm.n1639 1.0005
R40349 C10_N_btm.n1763 C10_N_btm.n1638 1.0005
R40350 C10_N_btm.n1762 C10_N_btm.n1637 1.0005
R40351 C10_N_btm.n1761 C10_N_btm.n1636 1.0005
R40352 C10_N_btm.n1760 C10_N_btm.n1635 1.0005
R40353 C10_N_btm.n1759 C10_N_btm.n1634 1.0005
R40354 C10_N_btm.n1758 C10_N_btm.n1633 1.0005
R40355 C10_N_btm.n1757 C10_N_btm.n1632 1.0005
R40356 C10_N_btm.n1756 C10_N_btm.n1631 1.0005
R40357 C10_N_btm.n1755 C10_N_btm.n1630 1.0005
R40358 C10_N_btm.n1754 C10_N_btm.n1629 1.0005
R40359 C10_N_btm.n1753 C10_N_btm.n1628 1.0005
R40360 C10_N_btm.n1752 C10_N_btm.n1627 1.0005
R40361 C10_N_btm.n1751 C10_N_btm.n1626 1.0005
R40362 C10_N_btm.n1750 C10_N_btm.n1625 1.0005
R40363 C10_N_btm.n1749 C10_N_btm.n1624 1.0005
R40364 C10_N_btm.n1748 C10_N_btm.n1623 1.0005
R40365 C10_N_btm.n1747 C10_N_btm.n1622 1.0005
R40366 C10_N_btm.n1746 C10_N_btm.n1621 1.0005
R40367 C10_N_btm.n1745 C10_N_btm.n1620 1.0005
R40368 C10_N_btm.n1744 C10_N_btm.n1619 1.0005
R40369 C10_N_btm.n1743 C10_N_btm.n1618 1.0005
R40370 C10_N_btm.n1742 C10_N_btm.n1617 1.0005
R40371 C10_N_btm.n1741 C10_N_btm.n1616 1.0005
R40372 C10_N_btm.n1740 C10_N_btm.n1615 1.0005
R40373 C10_N_btm.n1739 C10_N_btm.n1614 1.0005
R40374 C10_N_btm.n1738 C10_N_btm.n1613 1.0005
R40375 C10_N_btm.n1737 C10_N_btm.n1612 1.0005
R40376 C10_N_btm.n1736 C10_N_btm.n1611 1.0005
R40377 C10_N_btm.n1735 C10_N_btm.n1610 1.0005
R40378 C10_N_btm.n1734 C10_N_btm.n1609 1.0005
R40379 C10_N_btm.n1733 C10_N_btm.n1608 1.0005
R40380 C10_N_btm.n1732 C10_N_btm.n1607 1.0005
R40381 C10_N_btm.n1731 C10_N_btm.n1606 1.0005
R40382 C10_N_btm.n1730 C10_N_btm.n1605 1.0005
R40383 C10_N_btm.n1729 C10_N_btm.n1604 1.0005
R40384 C10_N_btm.n1728 C10_N_btm.n1603 1.0005
R40385 C10_N_btm.n1727 C10_N_btm.n1602 1.0005
R40386 C10_N_btm.n1726 C10_N_btm.n1601 1.0005
R40387 C10_N_btm.n1725 C10_N_btm.n1600 1.0005
R40388 C10_N_btm.n1967 C10_N_btm.n1599 1.0005
R40389 C10_N_btm.n1968 C10_N_btm.n1967 1.0005
R40390 C10_N_btm.n1725 C10_N_btm.n1722 1.0005
R40391 C10_N_btm.n1726 C10_N_btm.n1721 1.0005
R40392 C10_N_btm.n1727 C10_N_btm.n1720 1.0005
R40393 C10_N_btm.n1728 C10_N_btm.n1719 1.0005
R40394 C10_N_btm.n1729 C10_N_btm.n1718 1.0005
R40395 C10_N_btm.n1730 C10_N_btm.n1717 1.0005
R40396 C10_N_btm.n1731 C10_N_btm.n1716 1.0005
R40397 C10_N_btm.n1732 C10_N_btm.n1715 1.0005
R40398 C10_N_btm.n1733 C10_N_btm.n1714 1.0005
R40399 C10_N_btm.n1734 C10_N_btm.n1713 1.0005
R40400 C10_N_btm.n1735 C10_N_btm.n1712 1.0005
R40401 C10_N_btm.n1736 C10_N_btm.n1711 1.0005
R40402 C10_N_btm.n1737 C10_N_btm.n1710 1.0005
R40403 C10_N_btm.n1738 C10_N_btm.n1709 1.0005
R40404 C10_N_btm.n1739 C10_N_btm.n1708 1.0005
R40405 C10_N_btm.n1740 C10_N_btm.n1707 1.0005
R40406 C10_N_btm.n1741 C10_N_btm.n1706 1.0005
R40407 C10_N_btm.n1742 C10_N_btm.n1705 1.0005
R40408 C10_N_btm.n1743 C10_N_btm.n1704 1.0005
R40409 C10_N_btm.n1744 C10_N_btm.n1703 1.0005
R40410 C10_N_btm.n1745 C10_N_btm.n1702 1.0005
R40411 C10_N_btm.n1746 C10_N_btm.n1701 1.0005
R40412 C10_N_btm.n1747 C10_N_btm.n1700 1.0005
R40413 C10_N_btm.n1748 C10_N_btm.n1699 1.0005
R40414 C10_N_btm.n1749 C10_N_btm.n1698 1.0005
R40415 C10_N_btm.n1750 C10_N_btm.n1697 1.0005
R40416 C10_N_btm.n1751 C10_N_btm.n1696 1.0005
R40417 C10_N_btm.n1752 C10_N_btm.n1695 1.0005
R40418 C10_N_btm.n1753 C10_N_btm.n1694 1.0005
R40419 C10_N_btm.n1754 C10_N_btm.n1693 1.0005
R40420 C10_N_btm.n1755 C10_N_btm.n1692 1.0005
R40421 C10_N_btm.n1756 C10_N_btm.n1691 1.0005
R40422 C10_N_btm.n1757 C10_N_btm.n1690 1.0005
R40423 C10_N_btm.n1758 C10_N_btm.n1689 1.0005
R40424 C10_N_btm.n1759 C10_N_btm.n1688 1.0005
R40425 C10_N_btm.n1760 C10_N_btm.n1687 1.0005
R40426 C10_N_btm.n1761 C10_N_btm.n1686 1.0005
R40427 C10_N_btm.n1762 C10_N_btm.n1685 1.0005
R40428 C10_N_btm.n1763 C10_N_btm.n1684 1.0005
R40429 C10_N_btm.n1764 C10_N_btm.n1683 1.0005
R40430 C10_N_btm.n1765 C10_N_btm.n1682 1.0005
R40431 C10_N_btm.n1766 C10_N_btm.n1681 1.0005
R40432 C10_N_btm.n1767 C10_N_btm.n1680 1.0005
R40433 C10_N_btm.n1768 C10_N_btm.n1679 1.0005
R40434 C10_N_btm.n1769 C10_N_btm.n1678 1.0005
R40435 C10_N_btm.n1770 C10_N_btm.n1677 1.0005
R40436 C10_N_btm.n1771 C10_N_btm.n1676 1.0005
R40437 C10_N_btm.n1772 C10_N_btm.n1675 1.0005
R40438 C10_N_btm.n1773 C10_N_btm.n1674 1.0005
R40439 C10_N_btm.n1774 C10_N_btm.n1673 1.0005
R40440 C10_N_btm.n1775 C10_N_btm.n1672 1.0005
R40441 C10_N_btm.n1776 C10_N_btm.n1671 1.0005
R40442 C10_N_btm.n1777 C10_N_btm.n1670 1.0005
R40443 C10_N_btm.n1778 C10_N_btm.n1669 1.0005
R40444 C10_N_btm.n1779 C10_N_btm.n1668 1.0005
R40445 C10_N_btm.n1780 C10_N_btm.n1667 1.0005
R40446 C10_N_btm.n1781 C10_N_btm.n1666 1.0005
R40447 C10_N_btm.n1782 C10_N_btm.n1665 1.0005
R40448 C10_N_btm.n1783 C10_N_btm.n1664 1.0005
R40449 C10_N_btm.n1784 C10_N_btm.n1663 1.0005
R40450 C10_N_btm.n2916 C10_N_btm.n1660 1.0005
R40451 C10_N_btm.n2532 C10_N_btm.n1660 1.0005
R40452 C10_N_btm.n2030 C10_N_btm.n1663 1.0005
R40453 C10_N_btm.n2029 C10_N_btm.n1664 1.0005
R40454 C10_N_btm.n2028 C10_N_btm.n1665 1.0005
R40455 C10_N_btm.n2027 C10_N_btm.n1666 1.0005
R40456 C10_N_btm.n2026 C10_N_btm.n1667 1.0005
R40457 C10_N_btm.n2025 C10_N_btm.n1668 1.0005
R40458 C10_N_btm.n2024 C10_N_btm.n1669 1.0005
R40459 C10_N_btm.n2023 C10_N_btm.n1670 1.0005
R40460 C10_N_btm.n2022 C10_N_btm.n1671 1.0005
R40461 C10_N_btm.n2021 C10_N_btm.n1672 1.0005
R40462 C10_N_btm.n2020 C10_N_btm.n1673 1.0005
R40463 C10_N_btm.n2019 C10_N_btm.n1674 1.0005
R40464 C10_N_btm.n2018 C10_N_btm.n1675 1.0005
R40465 C10_N_btm.n2017 C10_N_btm.n1676 1.0005
R40466 C10_N_btm.n2016 C10_N_btm.n1677 1.0005
R40467 C10_N_btm.n2015 C10_N_btm.n1678 1.0005
R40468 C10_N_btm.n2014 C10_N_btm.n1679 1.0005
R40469 C10_N_btm.n2013 C10_N_btm.n1680 1.0005
R40470 C10_N_btm.n2012 C10_N_btm.n1681 1.0005
R40471 C10_N_btm.n2011 C10_N_btm.n1682 1.0005
R40472 C10_N_btm.n2010 C10_N_btm.n1683 1.0005
R40473 C10_N_btm.n2009 C10_N_btm.n1684 1.0005
R40474 C10_N_btm.n2008 C10_N_btm.n1685 1.0005
R40475 C10_N_btm.n2007 C10_N_btm.n1686 1.0005
R40476 C10_N_btm.n2006 C10_N_btm.n1687 1.0005
R40477 C10_N_btm.n2005 C10_N_btm.n1688 1.0005
R40478 C10_N_btm.n2004 C10_N_btm.n1689 1.0005
R40479 C10_N_btm.n2003 C10_N_btm.n1690 1.0005
R40480 C10_N_btm.n2002 C10_N_btm.n1691 1.0005
R40481 C10_N_btm.n2001 C10_N_btm.n1692 1.0005
R40482 C10_N_btm.n2000 C10_N_btm.n1693 1.0005
R40483 C10_N_btm.n1999 C10_N_btm.n1694 1.0005
R40484 C10_N_btm.n1998 C10_N_btm.n1695 1.0005
R40485 C10_N_btm.n1997 C10_N_btm.n1696 1.0005
R40486 C10_N_btm.n1996 C10_N_btm.n1697 1.0005
R40487 C10_N_btm.n1995 C10_N_btm.n1698 1.0005
R40488 C10_N_btm.n1994 C10_N_btm.n1699 1.0005
R40489 C10_N_btm.n1993 C10_N_btm.n1700 1.0005
R40490 C10_N_btm.n1992 C10_N_btm.n1701 1.0005
R40491 C10_N_btm.n1991 C10_N_btm.n1702 1.0005
R40492 C10_N_btm.n1990 C10_N_btm.n1703 1.0005
R40493 C10_N_btm.n1989 C10_N_btm.n1704 1.0005
R40494 C10_N_btm.n1988 C10_N_btm.n1705 1.0005
R40495 C10_N_btm.n1987 C10_N_btm.n1706 1.0005
R40496 C10_N_btm.n1986 C10_N_btm.n1707 1.0005
R40497 C10_N_btm.n1985 C10_N_btm.n1708 1.0005
R40498 C10_N_btm.n1984 C10_N_btm.n1709 1.0005
R40499 C10_N_btm.n1983 C10_N_btm.n1710 1.0005
R40500 C10_N_btm.n1982 C10_N_btm.n1711 1.0005
R40501 C10_N_btm.n1981 C10_N_btm.n1712 1.0005
R40502 C10_N_btm.n1980 C10_N_btm.n1713 1.0005
R40503 C10_N_btm.n1979 C10_N_btm.n1714 1.0005
R40504 C10_N_btm.n1978 C10_N_btm.n1715 1.0005
R40505 C10_N_btm.n1977 C10_N_btm.n1716 1.0005
R40506 C10_N_btm.n1976 C10_N_btm.n1717 1.0005
R40507 C10_N_btm.n1975 C10_N_btm.n1718 1.0005
R40508 C10_N_btm.n1974 C10_N_btm.n1719 1.0005
R40509 C10_N_btm.n1973 C10_N_btm.n1720 1.0005
R40510 C10_N_btm.n1972 C10_N_btm.n1721 1.0005
R40511 C10_N_btm.n1971 C10_N_btm.n1722 1.0005
R40512 C10_N_btm.n1970 C10_N_btm.n1968 1.0005
R40513 C10_N_btm.n2337 C10_N_btm.n1970 1.0005
R40514 C10_N_btm.n2095 C10_N_btm.n1971 1.0005
R40515 C10_N_btm.n2096 C10_N_btm.n1972 1.0005
R40516 C10_N_btm.n2097 C10_N_btm.n1973 1.0005
R40517 C10_N_btm.n2098 C10_N_btm.n1974 1.0005
R40518 C10_N_btm.n2099 C10_N_btm.n1975 1.0005
R40519 C10_N_btm.n2100 C10_N_btm.n1976 1.0005
R40520 C10_N_btm.n2101 C10_N_btm.n1977 1.0005
R40521 C10_N_btm.n2102 C10_N_btm.n1978 1.0005
R40522 C10_N_btm.n2103 C10_N_btm.n1979 1.0005
R40523 C10_N_btm.n2104 C10_N_btm.n1980 1.0005
R40524 C10_N_btm.n2105 C10_N_btm.n1981 1.0005
R40525 C10_N_btm.n2106 C10_N_btm.n1982 1.0005
R40526 C10_N_btm.n2107 C10_N_btm.n1983 1.0005
R40527 C10_N_btm.n2108 C10_N_btm.n1984 1.0005
R40528 C10_N_btm.n2109 C10_N_btm.n1985 1.0005
R40529 C10_N_btm.n2110 C10_N_btm.n1986 1.0005
R40530 C10_N_btm.n2111 C10_N_btm.n1987 1.0005
R40531 C10_N_btm.n2112 C10_N_btm.n1988 1.0005
R40532 C10_N_btm.n2113 C10_N_btm.n1989 1.0005
R40533 C10_N_btm.n2114 C10_N_btm.n1990 1.0005
R40534 C10_N_btm.n2115 C10_N_btm.n1991 1.0005
R40535 C10_N_btm.n2116 C10_N_btm.n1992 1.0005
R40536 C10_N_btm.n2117 C10_N_btm.n1993 1.0005
R40537 C10_N_btm.n2118 C10_N_btm.n1994 1.0005
R40538 C10_N_btm.n2119 C10_N_btm.n1995 1.0005
R40539 C10_N_btm.n2120 C10_N_btm.n1996 1.0005
R40540 C10_N_btm.n2121 C10_N_btm.n1997 1.0005
R40541 C10_N_btm.n2122 C10_N_btm.n1998 1.0005
R40542 C10_N_btm.n2123 C10_N_btm.n1999 1.0005
R40543 C10_N_btm.n2124 C10_N_btm.n2000 1.0005
R40544 C10_N_btm.n2125 C10_N_btm.n2001 1.0005
R40545 C10_N_btm.n2126 C10_N_btm.n2002 1.0005
R40546 C10_N_btm.n2127 C10_N_btm.n2003 1.0005
R40547 C10_N_btm.n2128 C10_N_btm.n2004 1.0005
R40548 C10_N_btm.n2129 C10_N_btm.n2005 1.0005
R40549 C10_N_btm.n2130 C10_N_btm.n2006 1.0005
R40550 C10_N_btm.n2131 C10_N_btm.n2007 1.0005
R40551 C10_N_btm.n2132 C10_N_btm.n2008 1.0005
R40552 C10_N_btm.n2133 C10_N_btm.n2009 1.0005
R40553 C10_N_btm.n2134 C10_N_btm.n2010 1.0005
R40554 C10_N_btm.n2135 C10_N_btm.n2011 1.0005
R40555 C10_N_btm.n2136 C10_N_btm.n2012 1.0005
R40556 C10_N_btm.n2137 C10_N_btm.n2013 1.0005
R40557 C10_N_btm.n2138 C10_N_btm.n2014 1.0005
R40558 C10_N_btm.n2139 C10_N_btm.n2015 1.0005
R40559 C10_N_btm.n2140 C10_N_btm.n2016 1.0005
R40560 C10_N_btm.n2141 C10_N_btm.n2017 1.0005
R40561 C10_N_btm.n2142 C10_N_btm.n2018 1.0005
R40562 C10_N_btm.n2143 C10_N_btm.n2019 1.0005
R40563 C10_N_btm.n2144 C10_N_btm.n2020 1.0005
R40564 C10_N_btm.n2145 C10_N_btm.n2021 1.0005
R40565 C10_N_btm.n2146 C10_N_btm.n2022 1.0005
R40566 C10_N_btm.n2147 C10_N_btm.n2023 1.0005
R40567 C10_N_btm.n2148 C10_N_btm.n2024 1.0005
R40568 C10_N_btm.n2149 C10_N_btm.n2025 1.0005
R40569 C10_N_btm.n2150 C10_N_btm.n2026 1.0005
R40570 C10_N_btm.n2151 C10_N_btm.n2027 1.0005
R40571 C10_N_btm.n2152 C10_N_btm.n2028 1.0005
R40572 C10_N_btm.n2153 C10_N_btm.n2029 1.0005
R40573 C10_N_btm.n2154 C10_N_btm.n2030 1.0005
R40574 C10_N_btm.n2532 C10_N_btm.n2531 1.0005
R40575 C10_N_btm.n2531 C10_N_btm.n2031 1.0005
R40576 C10_N_btm.n2154 C10_N_btm.n2033 1.0005
R40577 C10_N_btm.n2153 C10_N_btm.n2034 1.0005
R40578 C10_N_btm.n2152 C10_N_btm.n2035 1.0005
R40579 C10_N_btm.n2151 C10_N_btm.n2036 1.0005
R40580 C10_N_btm.n2150 C10_N_btm.n2037 1.0005
R40581 C10_N_btm.n2149 C10_N_btm.n2038 1.0005
R40582 C10_N_btm.n2148 C10_N_btm.n2039 1.0005
R40583 C10_N_btm.n2147 C10_N_btm.n2040 1.0005
R40584 C10_N_btm.n2146 C10_N_btm.n2041 1.0005
R40585 C10_N_btm.n2145 C10_N_btm.n2042 1.0005
R40586 C10_N_btm.n2144 C10_N_btm.n2043 1.0005
R40587 C10_N_btm.n2143 C10_N_btm.n2044 1.0005
R40588 C10_N_btm.n2142 C10_N_btm.n2045 1.0005
R40589 C10_N_btm.n2141 C10_N_btm.n2046 1.0005
R40590 C10_N_btm.n2140 C10_N_btm.n2047 1.0005
R40591 C10_N_btm.n2139 C10_N_btm.n2048 1.0005
R40592 C10_N_btm.n2138 C10_N_btm.n2049 1.0005
R40593 C10_N_btm.n2137 C10_N_btm.n2050 1.0005
R40594 C10_N_btm.n2136 C10_N_btm.n2051 1.0005
R40595 C10_N_btm.n2135 C10_N_btm.n2052 1.0005
R40596 C10_N_btm.n2134 C10_N_btm.n2053 1.0005
R40597 C10_N_btm.n2133 C10_N_btm.n2054 1.0005
R40598 C10_N_btm.n2132 C10_N_btm.n2055 1.0005
R40599 C10_N_btm.n2131 C10_N_btm.n2056 1.0005
R40600 C10_N_btm.n2130 C10_N_btm.n2057 1.0005
R40601 C10_N_btm.n2129 C10_N_btm.n2058 1.0005
R40602 C10_N_btm.n2128 C10_N_btm.n2059 1.0005
R40603 C10_N_btm.n2127 C10_N_btm.n2060 1.0005
R40604 C10_N_btm.n2126 C10_N_btm.n2061 1.0005
R40605 C10_N_btm.n2125 C10_N_btm.n2062 1.0005
R40606 C10_N_btm.n2124 C10_N_btm.n2063 1.0005
R40607 C10_N_btm.n2123 C10_N_btm.n2064 1.0005
R40608 C10_N_btm.n2122 C10_N_btm.n2065 1.0005
R40609 C10_N_btm.n2121 C10_N_btm.n2066 1.0005
R40610 C10_N_btm.n2120 C10_N_btm.n2067 1.0005
R40611 C10_N_btm.n2119 C10_N_btm.n2068 1.0005
R40612 C10_N_btm.n2118 C10_N_btm.n2069 1.0005
R40613 C10_N_btm.n2117 C10_N_btm.n2070 1.0005
R40614 C10_N_btm.n2116 C10_N_btm.n2071 1.0005
R40615 C10_N_btm.n2115 C10_N_btm.n2072 1.0005
R40616 C10_N_btm.n2114 C10_N_btm.n2073 1.0005
R40617 C10_N_btm.n2113 C10_N_btm.n2074 1.0005
R40618 C10_N_btm.n2112 C10_N_btm.n2075 1.0005
R40619 C10_N_btm.n2111 C10_N_btm.n2076 1.0005
R40620 C10_N_btm.n2110 C10_N_btm.n2077 1.0005
R40621 C10_N_btm.n2109 C10_N_btm.n2078 1.0005
R40622 C10_N_btm.n2108 C10_N_btm.n2079 1.0005
R40623 C10_N_btm.n2107 C10_N_btm.n2080 1.0005
R40624 C10_N_btm.n2106 C10_N_btm.n2081 1.0005
R40625 C10_N_btm.n2105 C10_N_btm.n2082 1.0005
R40626 C10_N_btm.n2104 C10_N_btm.n2083 1.0005
R40627 C10_N_btm.n2103 C10_N_btm.n2084 1.0005
R40628 C10_N_btm.n2102 C10_N_btm.n2085 1.0005
R40629 C10_N_btm.n2101 C10_N_btm.n2086 1.0005
R40630 C10_N_btm.n2100 C10_N_btm.n2087 1.0005
R40631 C10_N_btm.n2099 C10_N_btm.n2088 1.0005
R40632 C10_N_btm.n2098 C10_N_btm.n2089 1.0005
R40633 C10_N_btm.n2097 C10_N_btm.n2090 1.0005
R40634 C10_N_btm.n2096 C10_N_btm.n2091 1.0005
R40635 C10_N_btm.n2095 C10_N_btm.n2092 1.0005
R40636 C10_N_btm.n2338 C10_N_btm.n2337 1.0005
R40637 C10_N_btm.n2527 C10_N_btm.n1662 1.0005
R40638 C10_N_btm.n2722 C10_N_btm.n2721 1.0005
R40639 C10_N_btm.n2721 C10_N_btm.n1969 1.0005
R40640 C10_N_btm.n2912 C10_N_btm.n2911 1.0005
R40641 C10_N_btm.n2911 C10_N_btm.n1662 1.0005
R40642 C10_N_btm.n3106 C10_N_btm.n1598 1.0005
R40643 C10_N_btm.n2722 C10_N_btm.n1598 1.0005
R40644 C10_N_btm.n3296 C10_N_btm.n401 1.0005
R40645 C10_N_btm.n2912 C10_N_btm.n401 1.0005
R40646 C10_N_btm.n548 C10_N_btm.n546 1.0005
R40647 C10_N_btm.n549 C10_N_btm.n545 1.0005
R40648 C10_N_btm.n550 C10_N_btm.n544 1.0005
R40649 C10_N_btm.n551 C10_N_btm.n543 1.0005
R40650 C10_N_btm.n552 C10_N_btm.n542 1.0005
R40651 C10_N_btm.n553 C10_N_btm.n541 1.0005
R40652 C10_N_btm.n554 C10_N_btm.n540 1.0005
R40653 C10_N_btm.n555 C10_N_btm.n539 1.0005
R40654 C10_N_btm.n556 C10_N_btm.n538 1.0005
R40655 C10_N_btm.n558 C10_N_btm.n556 1.0005
R40656 C10_N_btm.n559 C10_N_btm.n555 1.0005
R40657 C10_N_btm.n560 C10_N_btm.n554 1.0005
R40658 C10_N_btm.n561 C10_N_btm.n553 1.0005
R40659 C10_N_btm.n562 C10_N_btm.n552 1.0005
R40660 C10_N_btm.n563 C10_N_btm.n551 1.0005
R40661 C10_N_btm.n564 C10_N_btm.n550 1.0005
R40662 C10_N_btm.n565 C10_N_btm.n549 1.0005
R40663 C10_N_btm.n1485 C10_N_btm.n548 1.0005
R40664 C10_N_btm.n1485 C10_N_btm.n1484 1.0005
R40665 C10_N_btm.n568 C10_N_btm.n565 1.0005
R40666 C10_N_btm.n569 C10_N_btm.n564 1.0005
R40667 C10_N_btm.n570 C10_N_btm.n563 1.0005
R40668 C10_N_btm.n571 C10_N_btm.n562 1.0005
R40669 C10_N_btm.n572 C10_N_btm.n561 1.0005
R40670 C10_N_btm.n573 C10_N_btm.n560 1.0005
R40671 C10_N_btm.n574 C10_N_btm.n559 1.0005
R40672 C10_N_btm.n1456 C10_N_btm.n558 1.0005
R40673 C10_N_btm.n1456 C10_N_btm.n1455 1.0005
R40674 C10_N_btm.n1393 C10_N_btm.n574 1.0005
R40675 C10_N_btm.n1392 C10_N_btm.n573 1.0005
R40676 C10_N_btm.n1391 C10_N_btm.n572 1.0005
R40677 C10_N_btm.n1390 C10_N_btm.n571 1.0005
R40678 C10_N_btm.n1389 C10_N_btm.n570 1.0005
R40679 C10_N_btm.n1388 C10_N_btm.n569 1.0005
R40680 C10_N_btm.n1387 C10_N_btm.n568 1.0005
R40681 C10_N_btm.n1484 C10_N_btm.n566 1.0005
R40682 C10_N_btm.n585 C10_N_btm.n566 1.0005
R40683 C10_N_btm.n1387 C10_N_btm.n584 1.0005
R40684 C10_N_btm.n1388 C10_N_btm.n583 1.0005
R40685 C10_N_btm.n1389 C10_N_btm.n582 1.0005
R40686 C10_N_btm.n1390 C10_N_btm.n581 1.0005
R40687 C10_N_btm.n1391 C10_N_btm.n580 1.0005
R40688 C10_N_btm.n1392 C10_N_btm.n579 1.0005
R40689 C10_N_btm.n1393 C10_N_btm.n578 1.0005
R40690 C10_N_btm.n1455 C10_N_btm.n575 1.0005
R40691 C10_N_btm.n1354 C10_N_btm.n575 1.0005
R40692 C10_N_btm.n594 C10_N_btm.n578 1.0005
R40693 C10_N_btm.n593 C10_N_btm.n579 1.0005
R40694 C10_N_btm.n592 C10_N_btm.n580 1.0005
R40695 C10_N_btm.n591 C10_N_btm.n581 1.0005
R40696 C10_N_btm.n590 C10_N_btm.n582 1.0005
R40697 C10_N_btm.n589 C10_N_btm.n583 1.0005
R40698 C10_N_btm.n588 C10_N_btm.n584 1.0005
R40699 C10_N_btm.n587 C10_N_btm.n585 1.0005
R40700 C10_N_btm.n637 C10_N_btm.n587 1.0005
R40701 C10_N_btm.n607 C10_N_btm.n588 1.0005
R40702 C10_N_btm.n608 C10_N_btm.n589 1.0005
R40703 C10_N_btm.n609 C10_N_btm.n590 1.0005
R40704 C10_N_btm.n610 C10_N_btm.n591 1.0005
R40705 C10_N_btm.n611 C10_N_btm.n592 1.0005
R40706 C10_N_btm.n612 C10_N_btm.n593 1.0005
R40707 C10_N_btm.n613 C10_N_btm.n594 1.0005
R40708 C10_N_btm.n1354 C10_N_btm.n1353 1.0005
R40709 C10_N_btm.n1353 C10_N_btm.n595 1.0005
R40710 C10_N_btm.n613 C10_N_btm.n598 1.0005
R40711 C10_N_btm.n612 C10_N_btm.n599 1.0005
R40712 C10_N_btm.n611 C10_N_btm.n600 1.0005
R40713 C10_N_btm.n610 C10_N_btm.n601 1.0005
R40714 C10_N_btm.n609 C10_N_btm.n602 1.0005
R40715 C10_N_btm.n608 C10_N_btm.n603 1.0005
R40716 C10_N_btm.n607 C10_N_btm.n604 1.0005
R40717 C10_N_btm.n638 C10_N_btm.n637 1.0005
R40718 C10_N_btm.n640 C10_N_btm.n638 1.0005
R40719 C10_N_btm.n641 C10_N_btm.n604 1.0005
R40720 C10_N_btm.n642 C10_N_btm.n603 1.0005
R40721 C10_N_btm.n643 C10_N_btm.n602 1.0005
R40722 C10_N_btm.n644 C10_N_btm.n601 1.0005
R40723 C10_N_btm.n645 C10_N_btm.n600 1.0005
R40724 C10_N_btm.n646 C10_N_btm.n599 1.0005
R40725 C10_N_btm.n647 C10_N_btm.n598 1.0005
R40726 C10_N_btm.n1287 C10_N_btm.n595 1.0005
R40727 C10_N_btm.n1287 C10_N_btm.n1286 1.0005
R40728 C10_N_btm.n666 C10_N_btm.n647 1.0005
R40729 C10_N_btm.n665 C10_N_btm.n646 1.0005
R40730 C10_N_btm.n664 C10_N_btm.n645 1.0005
R40731 C10_N_btm.n663 C10_N_btm.n644 1.0005
R40732 C10_N_btm.n662 C10_N_btm.n643 1.0005
R40733 C10_N_btm.n661 C10_N_btm.n642 1.0005
R40734 C10_N_btm.n660 C10_N_btm.n641 1.0005
R40735 C10_N_btm.n690 C10_N_btm.n640 1.0005
R40736 C10_N_btm.n691 C10_N_btm.n690 1.0005
R40737 C10_N_btm.n660 C10_N_btm.n657 1.0005
R40738 C10_N_btm.n661 C10_N_btm.n656 1.0005
R40739 C10_N_btm.n662 C10_N_btm.n655 1.0005
R40740 C10_N_btm.n663 C10_N_btm.n654 1.0005
R40741 C10_N_btm.n664 C10_N_btm.n653 1.0005
R40742 C10_N_btm.n665 C10_N_btm.n652 1.0005
R40743 C10_N_btm.n666 C10_N_btm.n651 1.0005
R40744 C10_N_btm.n1286 C10_N_btm.n648 1.0005
R40745 C10_N_btm.n1220 C10_N_btm.n648 1.0005
R40746 C10_N_btm.n700 C10_N_btm.n651 1.0005
R40747 C10_N_btm.n699 C10_N_btm.n652 1.0005
R40748 C10_N_btm.n698 C10_N_btm.n653 1.0005
R40749 C10_N_btm.n697 C10_N_btm.n654 1.0005
R40750 C10_N_btm.n696 C10_N_btm.n655 1.0005
R40751 C10_N_btm.n695 C10_N_btm.n656 1.0005
R40752 C10_N_btm.n694 C10_N_btm.n657 1.0005
R40753 C10_N_btm.n693 C10_N_btm.n691 1.0005
R40754 C10_N_btm.n743 C10_N_btm.n693 1.0005
R40755 C10_N_btm.n713 C10_N_btm.n694 1.0005
R40756 C10_N_btm.n714 C10_N_btm.n695 1.0005
R40757 C10_N_btm.n715 C10_N_btm.n696 1.0005
R40758 C10_N_btm.n716 C10_N_btm.n697 1.0005
R40759 C10_N_btm.n717 C10_N_btm.n698 1.0005
R40760 C10_N_btm.n718 C10_N_btm.n699 1.0005
R40761 C10_N_btm.n719 C10_N_btm.n700 1.0005
R40762 C10_N_btm.n1220 C10_N_btm.n1219 1.0005
R40763 C10_N_btm.n1219 C10_N_btm.n701 1.0005
R40764 C10_N_btm.n719 C10_N_btm.n704 1.0005
R40765 C10_N_btm.n718 C10_N_btm.n705 1.0005
R40766 C10_N_btm.n717 C10_N_btm.n706 1.0005
R40767 C10_N_btm.n716 C10_N_btm.n707 1.0005
R40768 C10_N_btm.n715 C10_N_btm.n708 1.0005
R40769 C10_N_btm.n714 C10_N_btm.n709 1.0005
R40770 C10_N_btm.n713 C10_N_btm.n710 1.0005
R40771 C10_N_btm.n744 C10_N_btm.n743 1.0005
R40772 C10_N_btm.n746 C10_N_btm.n744 1.0005
R40773 C10_N_btm.n747 C10_N_btm.n710 1.0005
R40774 C10_N_btm.n748 C10_N_btm.n709 1.0005
R40775 C10_N_btm.n749 C10_N_btm.n708 1.0005
R40776 C10_N_btm.n750 C10_N_btm.n707 1.0005
R40777 C10_N_btm.n751 C10_N_btm.n706 1.0005
R40778 C10_N_btm.n752 C10_N_btm.n705 1.0005
R40779 C10_N_btm.n753 C10_N_btm.n704 1.0005
R40780 C10_N_btm.n1153 C10_N_btm.n701 1.0005
R40781 C10_N_btm.n1153 C10_N_btm.n1152 1.0005
R40782 C10_N_btm.n772 C10_N_btm.n753 1.0005
R40783 C10_N_btm.n771 C10_N_btm.n752 1.0005
R40784 C10_N_btm.n770 C10_N_btm.n751 1.0005
R40785 C10_N_btm.n769 C10_N_btm.n750 1.0005
R40786 C10_N_btm.n768 C10_N_btm.n749 1.0005
R40787 C10_N_btm.n767 C10_N_btm.n748 1.0005
R40788 C10_N_btm.n766 C10_N_btm.n747 1.0005
R40789 C10_N_btm.n796 C10_N_btm.n746 1.0005
R40790 C10_N_btm.n797 C10_N_btm.n796 1.0005
R40791 C10_N_btm.n766 C10_N_btm.n763 1.0005
R40792 C10_N_btm.n767 C10_N_btm.n762 1.0005
R40793 C10_N_btm.n768 C10_N_btm.n761 1.0005
R40794 C10_N_btm.n769 C10_N_btm.n760 1.0005
R40795 C10_N_btm.n770 C10_N_btm.n759 1.0005
R40796 C10_N_btm.n771 C10_N_btm.n758 1.0005
R40797 C10_N_btm.n772 C10_N_btm.n757 1.0005
R40798 C10_N_btm.n1152 C10_N_btm.n754 1.0005
R40799 C10_N_btm.n1086 C10_N_btm.n754 1.0005
R40800 C10_N_btm.n806 C10_N_btm.n757 1.0005
R40801 C10_N_btm.n805 C10_N_btm.n758 1.0005
R40802 C10_N_btm.n804 C10_N_btm.n759 1.0005
R40803 C10_N_btm.n803 C10_N_btm.n760 1.0005
R40804 C10_N_btm.n802 C10_N_btm.n761 1.0005
R40805 C10_N_btm.n801 C10_N_btm.n762 1.0005
R40806 C10_N_btm.n800 C10_N_btm.n763 1.0005
R40807 C10_N_btm.n799 C10_N_btm.n797 1.0005
R40808 C10_N_btm.n849 C10_N_btm.n799 1.0005
R40809 C10_N_btm.n819 C10_N_btm.n800 1.0005
R40810 C10_N_btm.n820 C10_N_btm.n801 1.0005
R40811 C10_N_btm.n821 C10_N_btm.n802 1.0005
R40812 C10_N_btm.n822 C10_N_btm.n803 1.0005
R40813 C10_N_btm.n823 C10_N_btm.n804 1.0005
R40814 C10_N_btm.n824 C10_N_btm.n805 1.0005
R40815 C10_N_btm.n825 C10_N_btm.n806 1.0005
R40816 C10_N_btm.n1086 C10_N_btm.n1085 1.0005
R40817 C10_N_btm.n1085 C10_N_btm.n807 1.0005
R40818 C10_N_btm.n825 C10_N_btm.n810 1.0005
R40819 C10_N_btm.n824 C10_N_btm.n811 1.0005
R40820 C10_N_btm.n823 C10_N_btm.n812 1.0005
R40821 C10_N_btm.n822 C10_N_btm.n813 1.0005
R40822 C10_N_btm.n821 C10_N_btm.n814 1.0005
R40823 C10_N_btm.n820 C10_N_btm.n815 1.0005
R40824 C10_N_btm.n819 C10_N_btm.n816 1.0005
R40825 C10_N_btm.n850 C10_N_btm.n849 1.0005
R40826 C10_N_btm.n852 C10_N_btm.n850 1.0005
R40827 C10_N_btm.n853 C10_N_btm.n816 1.0005
R40828 C10_N_btm.n854 C10_N_btm.n815 1.0005
R40829 C10_N_btm.n855 C10_N_btm.n814 1.0005
R40830 C10_N_btm.n856 C10_N_btm.n813 1.0005
R40831 C10_N_btm.n857 C10_N_btm.n812 1.0005
R40832 C10_N_btm.n858 C10_N_btm.n811 1.0005
R40833 C10_N_btm.n859 C10_N_btm.n810 1.0005
R40834 C10_N_btm.n1019 C10_N_btm.n807 1.0005
R40835 C10_N_btm.n1019 C10_N_btm.n1018 1.0005
R40836 C10_N_btm.n878 C10_N_btm.n859 1.0005
R40837 C10_N_btm.n877 C10_N_btm.n858 1.0005
R40838 C10_N_btm.n876 C10_N_btm.n857 1.0005
R40839 C10_N_btm.n875 C10_N_btm.n856 1.0005
R40840 C10_N_btm.n874 C10_N_btm.n855 1.0005
R40841 C10_N_btm.n873 C10_N_btm.n854 1.0005
R40842 C10_N_btm.n872 C10_N_btm.n853 1.0005
R40843 C10_N_btm.n902 C10_N_btm.n852 1.0005
R40844 C10_N_btm.n903 C10_N_btm.n902 1.0005
R40845 C10_N_btm.n872 C10_N_btm.n869 1.0005
R40846 C10_N_btm.n873 C10_N_btm.n868 1.0005
R40847 C10_N_btm.n874 C10_N_btm.n867 1.0005
R40848 C10_N_btm.n875 C10_N_btm.n866 1.0005
R40849 C10_N_btm.n876 C10_N_btm.n865 1.0005
R40850 C10_N_btm.n877 C10_N_btm.n864 1.0005
R40851 C10_N_btm.n878 C10_N_btm.n863 1.0005
R40852 C10_N_btm.n1018 C10_N_btm.n860 1.0005
R40853 C10_N_btm.n952 C10_N_btm.n860 1.0005
R40854 C10_N_btm.n912 C10_N_btm.n863 1.0005
R40855 C10_N_btm.n911 C10_N_btm.n864 1.0005
R40856 C10_N_btm.n910 C10_N_btm.n865 1.0005
R40857 C10_N_btm.n909 C10_N_btm.n866 1.0005
R40858 C10_N_btm.n908 C10_N_btm.n867 1.0005
R40859 C10_N_btm.n907 C10_N_btm.n868 1.0005
R40860 C10_N_btm.n906 C10_N_btm.n869 1.0005
R40861 C10_N_btm.n905 C10_N_btm.n903 1.0005
R40862 C10_N_btm.n920 C10_N_btm.n905 1.0005
R40863 C10_N_btm.n919 C10_N_btm.n906 1.0005
R40864 C10_N_btm.n918 C10_N_btm.n907 1.0005
R40865 C10_N_btm.n917 C10_N_btm.n908 1.0005
R40866 C10_N_btm.n916 C10_N_btm.n909 1.0005
R40867 C10_N_btm.n915 C10_N_btm.n910 1.0005
R40868 C10_N_btm.n914 C10_N_btm.n911 1.0005
R40869 C10_N_btm.n913 C10_N_btm.n912 1.0005
R40870 C10_N_btm.n952 C10_N_btm.n951 1.0005
R40871 C10_N_btm.n947 C10_N_btm.n862 1.0005
R40872 C10_N_btm.n982 C10_N_btm.n904 1.0005
R40873 C10_N_btm.n983 C10_N_btm.n982 1.0005
R40874 C10_N_btm.n1013 C10_N_btm.n862 1.0005
R40875 C10_N_btm.n1014 C10_N_btm.n1013 1.0005
R40876 C10_N_btm.n983 C10_N_btm.n851 1.0005
R40877 C10_N_btm.n1049 C10_N_btm.n851 1.0005
R40878 C10_N_btm.n1014 C10_N_btm.n809 1.0005
R40879 C10_N_btm.n1080 C10_N_btm.n809 1.0005
R40880 C10_N_btm.n1050 C10_N_btm.n1049 1.0005
R40881 C10_N_btm.n1050 C10_N_btm.n798 1.0005
R40882 C10_N_btm.n1081 C10_N_btm.n1080 1.0005
R40883 C10_N_btm.n1081 C10_N_btm.n756 1.0005
R40884 C10_N_btm.n1116 C10_N_btm.n798 1.0005
R40885 C10_N_btm.n1117 C10_N_btm.n1116 1.0005
R40886 C10_N_btm.n1147 C10_N_btm.n756 1.0005
R40887 C10_N_btm.n1148 C10_N_btm.n1147 1.0005
R40888 C10_N_btm.n1117 C10_N_btm.n745 1.0005
R40889 C10_N_btm.n1183 C10_N_btm.n745 1.0005
R40890 C10_N_btm.n1148 C10_N_btm.n703 1.0005
R40891 C10_N_btm.n1214 C10_N_btm.n703 1.0005
R40892 C10_N_btm.n1184 C10_N_btm.n1183 1.0005
R40893 C10_N_btm.n1184 C10_N_btm.n692 1.0005
R40894 C10_N_btm.n1215 C10_N_btm.n1214 1.0005
R40895 C10_N_btm.n1215 C10_N_btm.n650 1.0005
R40896 C10_N_btm.n1250 C10_N_btm.n692 1.0005
R40897 C10_N_btm.n1251 C10_N_btm.n1250 1.0005
R40898 C10_N_btm.n1281 C10_N_btm.n650 1.0005
R40899 C10_N_btm.n1282 C10_N_btm.n1281 1.0005
R40900 C10_N_btm.n1251 C10_N_btm.n639 1.0005
R40901 C10_N_btm.n1317 C10_N_btm.n639 1.0005
R40902 C10_N_btm.n1282 C10_N_btm.n597 1.0005
R40903 C10_N_btm.n1348 C10_N_btm.n597 1.0005
R40904 C10_N_btm.n1318 C10_N_btm.n1317 1.0005
R40905 C10_N_btm.n1318 C10_N_btm.n586 1.0005
R40906 C10_N_btm.n1349 C10_N_btm.n1348 1.0005
R40907 C10_N_btm.n1349 C10_N_btm.n577 1.0005
R40908 C10_N_btm.n1384 C10_N_btm.n586 1.0005
R40909 C10_N_btm.n1420 C10_N_btm.n1384 1.0005
R40910 C10_N_btm.n1450 C10_N_btm.n577 1.0005
R40911 C10_N_btm.n1451 C10_N_btm.n1450 1.0005
R40912 C10_N_btm.n1420 C10_N_btm.n1419 1.0005
R40913 C10_N_btm.n1419 C10_N_btm.n1386 1.0005
R40914 C10_N_btm.n1451 C10_N_btm.n557 1.0005
R40915 C10_N_btm.n1515 C10_N_btm.n557 1.0005
R40916 C10_N_btm.n1386 C10_N_btm.n547 1.0005
R40917 C10_N_btm.n1597 C10_N_btm.n547 1.0005
R40918 C10_N_btm.n1516 C10_N_btm.n1515 1.0005
R40919 C10_N_btm.n1516 C10_N_btm.n537 1.0005
R40920 C10_N_btm.n1517 C10_N_btm.n536 1.0005
R40921 C10_N_btm.n1518 C10_N_btm.n535 1.0005
R40922 C10_N_btm.n1519 C10_N_btm.n534 1.0005
R40923 C10_N_btm.n1520 C10_N_btm.n533 1.0005
R40924 C10_N_btm.n1521 C10_N_btm.n532 1.0005
R40925 C10_N_btm.n1522 C10_N_btm.n531 1.0005
R40926 C10_N_btm.n1523 C10_N_btm.n530 1.0005
R40927 C10_N_btm.n1524 C10_N_btm.n529 1.0005
R40928 C10_N_btm.n1525 C10_N_btm.n528 1.0005
R40929 C10_N_btm.n1526 C10_N_btm.n527 1.0005
R40930 C10_N_btm.n1527 C10_N_btm.n526 1.0005
R40931 C10_N_btm.n1528 C10_N_btm.n525 1.0005
R40932 C10_N_btm.n3107 C10_N_btm.n1597 1.0005
R40933 C10_N_btm.n3107 C10_N_btm.n3106 1.0005
R40934 C10_N_btm.n3297 C10_N_btm.n348 1.0005
R40935 C10_N_btm.n3297 C10_N_btm.n3296 1.0005
R40936 C10_N_btm.n3333 C10_N_btm.n3332 1.0005
R40937 C10_N_btm.n3332 C10_N_btm.n390 1.0005
R40938 C10_N_btm.n3364 C10_N_btm.n3363 1.0005
R40939 C10_N_btm.n3363 C10_N_btm.n348 1.0005
R40940 C10_N_btm.n3399 C10_N_btm.n337 1.0005
R40941 C10_N_btm.n3333 C10_N_btm.n337 1.0005
R40942 C10_N_btm.n3430 C10_N_btm.n295 1.0005
R40943 C10_N_btm.n3364 C10_N_btm.n295 1.0005
R40944 C10_N_btm.n3400 C10_N_btm.n284 1.0005
R40945 C10_N_btm.n3400 C10_N_btm.n3399 1.0005
R40946 C10_N_btm.n3431 C10_N_btm.n242 1.0005
R40947 C10_N_btm.n3431 C10_N_btm.n3430 1.0005
R40948 C10_N_btm.n3467 C10_N_btm.n3466 1.0005
R40949 C10_N_btm.n3466 C10_N_btm.n284 1.0005
R40950 C10_N_btm.n3498 C10_N_btm.n3497 1.0005
R40951 C10_N_btm.n3497 C10_N_btm.n242 1.0005
R40952 C10_N_btm.n3533 C10_N_btm.n231 1.0005
R40953 C10_N_btm.n3467 C10_N_btm.n231 1.0005
R40954 C10_N_btm.n3564 C10_N_btm.n189 1.0005
R40955 C10_N_btm.n3498 C10_N_btm.n189 1.0005
R40956 C10_N_btm.n3534 C10_N_btm.n178 1.0005
R40957 C10_N_btm.n3534 C10_N_btm.n3533 1.0005
R40958 C10_N_btm.n3565 C10_N_btm.n136 1.0005
R40959 C10_N_btm.n3565 C10_N_btm.n3564 1.0005
R40960 C10_N_btm.n3601 C10_N_btm.n3600 1.0005
R40961 C10_N_btm.n3600 C10_N_btm.n178 1.0005
R40962 C10_N_btm.n3632 C10_N_btm.n3631 1.0005
R40963 C10_N_btm.n3631 C10_N_btm.n136 1.0005
R40964 C10_N_btm.n3667 C10_N_btm.n125 1.0005
R40965 C10_N_btm.n3601 C10_N_btm.n125 1.0005
R40966 C10_N_btm.n3698 C10_N_btm.n83 1.0005
R40967 C10_N_btm.n3632 C10_N_btm.n83 1.0005
R40968 C10_N_btm.n3668 C10_N_btm.n72 1.0005
R40969 C10_N_btm.n3668 C10_N_btm.n3667 1.0005
R40970 C10_N_btm.n3699 C10_N_btm.n63 1.0005
R40971 C10_N_btm.n3699 C10_N_btm.n3698 1.0005
R40972 C10_N_btm.n3770 C10_N_btm.n3734 1.0005
R40973 C10_N_btm.n3734 C10_N_btm.n72 1.0005
R40974 C10_N_btm.n3801 C10_N_btm.n3800 1.0005
R40975 C10_N_btm.n3800 C10_N_btm.n63 1.0005
R40976 C10_N_btm.n3769 C10_N_btm.n3736 1.0005
R40977 C10_N_btm.n3770 C10_N_btm.n3769 1.0005
R40978 C10_N_btm.n3865 C10_N_btm.n43 1.0005
R40979 C10_N_btm.n3801 C10_N_btm.n43 1.0005
R40980 C10_N_btm.n3896 C10_N_btm.n33 1.0005
R40981 C10_N_btm.n3736 C10_N_btm.n33 1.0005
R40982 C10_N_btm.n3866 C10_N_btm.n3865 1.0005
R40983 C10_N_btm.n3897 C10_N_btm.n3896 1.0005
R40984 C10_N_btm.n4 C10_N_btm.n2 0.71925
R40985 C10_N_btm.n8 C10_N_btm.n6 0.71925
R40986 C10_N_btm.n12 C10_N_btm.n10 0.71925
R40987 C10_N_btm.n6 C10_N_btm.n4 0.688
R40988 C10_N_btm.n10 C10_N_btm.n8 0.688
R40989 C10_N_btm.n506 C10_N_btm.n505 0.679419
R40990 C10_N_btm.n2340 C10_N_btm.n2339 0.679419
R40991 C10_N_btm.n2526 C10_N_btm.n2525 0.679419
R40992 C10_N_btm.n2530 C10_N_btm.n2528 0.679419
R40993 C10_N_btm.n2094 C10_N_btm.n2093 0.679419
R40994 C10_N_btm.n2720 C10_N_btm.n2719 0.679419
R40995 C10_N_btm.n2534 C10_N_btm.n2533 0.679419
R40996 C10_N_btm.n2910 C10_N_btm.n2909 0.679419
R40997 C10_N_btm.n2724 C10_N_btm.n2723 0.679419
R40998 C10_N_btm.n1724 C10_N_btm.n1723 0.679419
R40999 C10_N_btm.n2915 C10_N_btm.n2913 0.679419
R41000 C10_N_btm.n2919 C10_N_btm.n2918 0.679419
R41001 C10_N_btm.n3105 C10_N_btm.n3104 0.679419
R41002 C10_N_btm.n950 C10_N_btm.n948 0.679419
R41003 C10_N_btm.n922 C10_N_btm.n921 0.679419
R41004 C10_N_btm.n981 C10_N_btm.n980 0.679419
R41005 C10_N_btm.n954 C10_N_btm.n953 0.679419
R41006 C10_N_btm.n1012 C10_N_btm.n1011 0.679419
R41007 C10_N_btm.n985 C10_N_btm.n984 0.679419
R41008 C10_N_btm.n871 C10_N_btm.n870 0.679419
R41009 C10_N_btm.n1017 C10_N_btm.n1015 0.679419
R41010 C10_N_btm.n1021 C10_N_btm.n1020 0.679419
R41011 C10_N_btm.n1048 C10_N_btm.n1047 0.679419
R41012 C10_N_btm.n1052 C10_N_btm.n1051 0.679419
R41013 C10_N_btm.n1079 C10_N_btm.n1078 0.679419
R41014 C10_N_btm.n1084 C10_N_btm.n1082 0.679419
R41015 C10_N_btm.n818 C10_N_btm.n817 0.679419
R41016 C10_N_btm.n1115 C10_N_btm.n1114 0.679419
R41017 C10_N_btm.n1088 C10_N_btm.n1087 0.679419
R41018 C10_N_btm.n1146 C10_N_btm.n1145 0.679419
R41019 C10_N_btm.n1119 C10_N_btm.n1118 0.679419
R41020 C10_N_btm.n765 C10_N_btm.n764 0.679419
R41021 C10_N_btm.n1151 C10_N_btm.n1149 0.679419
R41022 C10_N_btm.n1155 C10_N_btm.n1154 0.679419
R41023 C10_N_btm.n1182 C10_N_btm.n1181 0.679419
R41024 C10_N_btm.n1186 C10_N_btm.n1185 0.679419
R41025 C10_N_btm.n1213 C10_N_btm.n1212 0.679419
R41026 C10_N_btm.n1218 C10_N_btm.n1216 0.679419
R41027 C10_N_btm.n712 C10_N_btm.n711 0.679419
R41028 C10_N_btm.n1249 C10_N_btm.n1248 0.679419
R41029 C10_N_btm.n1222 C10_N_btm.n1221 0.679419
R41030 C10_N_btm.n1280 C10_N_btm.n1279 0.679419
R41031 C10_N_btm.n1253 C10_N_btm.n1252 0.679419
R41032 C10_N_btm.n659 C10_N_btm.n658 0.679419
R41033 C10_N_btm.n1285 C10_N_btm.n1283 0.679419
R41034 C10_N_btm.n1289 C10_N_btm.n1288 0.679419
R41035 C10_N_btm.n1316 C10_N_btm.n1315 0.679419
R41036 C10_N_btm.n1320 C10_N_btm.n1319 0.679419
R41037 C10_N_btm.n1347 C10_N_btm.n1346 0.679419
R41038 C10_N_btm.n1352 C10_N_btm.n1350 0.679419
R41039 C10_N_btm.n606 C10_N_btm.n605 0.679419
R41040 C10_N_btm.n1383 C10_N_btm.n1382 0.679419
R41041 C10_N_btm.n1356 C10_N_btm.n1355 0.679419
R41042 C10_N_btm.n1449 C10_N_btm.n1448 0.679419
R41043 C10_N_btm.n1422 C10_N_btm.n1421 0.679419
R41044 C10_N_btm.n1418 C10_N_btm.n1417 0.679419
R41045 C10_N_btm.n1454 C10_N_btm.n1452 0.679419
R41046 C10_N_btm.n1458 C10_N_btm.n1457 0.679419
R41047 C10_N_btm.n1385 C10_N_btm.n567 0.679419
R41048 C10_N_btm.n1487 C10_N_btm.n1486 0.679419
R41049 C10_N_btm.n1514 C10_N_btm.n1513 0.679419
R41050 C10_N_btm.n1530 C10_N_btm.n1529 0.679419
R41051 C10_N_btm.n1596 C10_N_btm.n1595 0.679419
R41052 C10_N_btm.n3109 C10_N_btm.n3108 0.679419
R41053 C10_N_btm.n3295 C10_N_btm.n3294 0.679419
R41054 C10_N_btm.n3300 C10_N_btm.n3298 0.679419
R41055 C10_N_btm.n3331 C10_N_btm.n3330 0.679419
R41056 C10_N_btm.n3304 C10_N_btm.n3303 0.679419
R41057 C10_N_btm.n3362 C10_N_btm.n3361 0.679419
R41058 C10_N_btm.n3335 C10_N_btm.n3334 0.679419
R41059 C10_N_btm.n357 C10_N_btm.n356 0.679419
R41060 C10_N_btm.n3367 C10_N_btm.n3365 0.679419
R41061 C10_N_btm.n3371 C10_N_btm.n3370 0.679419
R41062 C10_N_btm.n3398 C10_N_btm.n3397 0.679419
R41063 C10_N_btm.n3402 C10_N_btm.n3401 0.679419
R41064 C10_N_btm.n3429 C10_N_btm.n3428 0.679419
R41065 C10_N_btm.n3434 C10_N_btm.n3432 0.679419
R41066 C10_N_btm.n304 C10_N_btm.n303 0.679419
R41067 C10_N_btm.n3465 C10_N_btm.n3464 0.679419
R41068 C10_N_btm.n3438 C10_N_btm.n3437 0.679419
R41069 C10_N_btm.n3496 C10_N_btm.n3495 0.679419
R41070 C10_N_btm.n3469 C10_N_btm.n3468 0.679419
R41071 C10_N_btm.n251 C10_N_btm.n250 0.679419
R41072 C10_N_btm.n3501 C10_N_btm.n3499 0.679419
R41073 C10_N_btm.n3505 C10_N_btm.n3504 0.679419
R41074 C10_N_btm.n3532 C10_N_btm.n3531 0.679419
R41075 C10_N_btm.n3536 C10_N_btm.n3535 0.679419
R41076 C10_N_btm.n3563 C10_N_btm.n3562 0.679419
R41077 C10_N_btm.n3568 C10_N_btm.n3566 0.679419
R41078 C10_N_btm.n198 C10_N_btm.n197 0.679419
R41079 C10_N_btm.n3599 C10_N_btm.n3598 0.679419
R41080 C10_N_btm.n3572 C10_N_btm.n3571 0.679419
R41081 C10_N_btm.n3630 C10_N_btm.n3629 0.679419
R41082 C10_N_btm.n3603 C10_N_btm.n3602 0.679419
R41083 C10_N_btm.n145 C10_N_btm.n144 0.679419
R41084 C10_N_btm.n3635 C10_N_btm.n3633 0.679419
R41085 C10_N_btm.n3639 C10_N_btm.n3638 0.679419
R41086 C10_N_btm.n3666 C10_N_btm.n3665 0.679419
R41087 C10_N_btm.n3670 C10_N_btm.n3669 0.679419
R41088 C10_N_btm.n3697 C10_N_btm.n3696 0.679419
R41089 C10_N_btm.n3702 C10_N_btm.n3700 0.679419
R41090 C10_N_btm.n92 C10_N_btm.n91 0.679419
R41091 C10_N_btm.n3733 C10_N_btm.n3732 0.679419
R41092 C10_N_btm.n3706 C10_N_btm.n3705 0.679419
R41093 C10_N_btm.n3799 C10_N_btm.n3798 0.679419
R41094 C10_N_btm.n3772 C10_N_btm.n3771 0.679419
R41095 C10_N_btm.n3768 C10_N_btm.n3767 0.679419
R41096 C10_N_btm.n3804 C10_N_btm.n3802 0.679419
R41097 C10_N_btm.n3808 C10_N_btm.n3807 0.679419
R41098 C10_N_btm.n3735 C10_N_btm.n53 0.679419
R41099 C10_N_btm.n3837 C10_N_btm.n3836 0.679419
R41100 C10_N_btm.n3864 C10_N_btm.n3863 0.679419
R41101 C10_N_btm.n3868 C10_N_btm.n3867 0.679419
R41102 C10_N_btm.n3895 C10_N_btm.n3894 0.679419
R41103 C10_N_btm.n14 C10_N_btm.n12 0.672375
R41104 C10_N_btm.n470 C10_N_btm.n469 0.6255
R41105 C10_N_btm.n473 C10_N_btm.n472 0.6255
R41106 C10_N_btm.n476 C10_N_btm.n475 0.6255
R41107 C10_N_btm.n479 C10_N_btm.n478 0.6255
R41108 C10_N_btm.n482 C10_N_btm.n481 0.6255
R41109 C10_N_btm.n485 C10_N_btm.n484 0.6255
R41110 C10_N_btm.n488 C10_N_btm.n487 0.6255
R41111 C10_N_btm.n491 C10_N_btm.n490 0.6255
R41112 C10_N_btm.n494 C10_N_btm.n493 0.6255
R41113 C10_N_btm.n497 C10_N_btm.n496 0.6255
R41114 C10_N_btm.n500 C10_N_btm.n499 0.6255
R41115 C10_N_btm.n503 C10_N_btm.n502 0.6255
R41116 C10_N_btm.n2343 C10_N_btm.n2342 0.6255
R41117 C10_N_btm.n2346 C10_N_btm.n2345 0.6255
R41118 C10_N_btm.n2349 C10_N_btm.n2348 0.6255
R41119 C10_N_btm.n2352 C10_N_btm.n2351 0.6255
R41120 C10_N_btm.n2355 C10_N_btm.n2354 0.6255
R41121 C10_N_btm.n2358 C10_N_btm.n2357 0.6255
R41122 C10_N_btm.n2361 C10_N_btm.n2360 0.6255
R41123 C10_N_btm.n2364 C10_N_btm.n2363 0.6255
R41124 C10_N_btm.n2367 C10_N_btm.n2366 0.6255
R41125 C10_N_btm.n2370 C10_N_btm.n2369 0.6255
R41126 C10_N_btm.n2373 C10_N_btm.n2372 0.6255
R41127 C10_N_btm.n2376 C10_N_btm.n2375 0.6255
R41128 C10_N_btm.n2379 C10_N_btm.n2378 0.6255
R41129 C10_N_btm.n2382 C10_N_btm.n2381 0.6255
R41130 C10_N_btm.n2385 C10_N_btm.n2384 0.6255
R41131 C10_N_btm.n2388 C10_N_btm.n2387 0.6255
R41132 C10_N_btm.n2391 C10_N_btm.n2390 0.6255
R41133 C10_N_btm.n2394 C10_N_btm.n2393 0.6255
R41134 C10_N_btm.n2397 C10_N_btm.n2396 0.6255
R41135 C10_N_btm.n2400 C10_N_btm.n2399 0.6255
R41136 C10_N_btm.n2403 C10_N_btm.n2402 0.6255
R41137 C10_N_btm.n2406 C10_N_btm.n2405 0.6255
R41138 C10_N_btm.n2409 C10_N_btm.n2408 0.6255
R41139 C10_N_btm.n2412 C10_N_btm.n2411 0.6255
R41140 C10_N_btm.n2415 C10_N_btm.n2414 0.6255
R41141 C10_N_btm.n2418 C10_N_btm.n2417 0.6255
R41142 C10_N_btm.n2421 C10_N_btm.n2420 0.6255
R41143 C10_N_btm.n2424 C10_N_btm.n2423 0.6255
R41144 C10_N_btm.n2427 C10_N_btm.n2426 0.6255
R41145 C10_N_btm.n2430 C10_N_btm.n2429 0.6255
R41146 C10_N_btm.n2433 C10_N_btm.n2432 0.6255
R41147 C10_N_btm.n2436 C10_N_btm.n2435 0.6255
R41148 C10_N_btm.n2439 C10_N_btm.n2438 0.6255
R41149 C10_N_btm.n2442 C10_N_btm.n2441 0.6255
R41150 C10_N_btm.n2445 C10_N_btm.n2444 0.6255
R41151 C10_N_btm.n2448 C10_N_btm.n2447 0.6255
R41152 C10_N_btm.n2451 C10_N_btm.n2450 0.6255
R41153 C10_N_btm.n2454 C10_N_btm.n2453 0.6255
R41154 C10_N_btm.n2457 C10_N_btm.n2456 0.6255
R41155 C10_N_btm.n2460 C10_N_btm.n2459 0.6255
R41156 C10_N_btm.n2463 C10_N_btm.n2462 0.6255
R41157 C10_N_btm.n2466 C10_N_btm.n2465 0.6255
R41158 C10_N_btm.n2469 C10_N_btm.n2468 0.6255
R41159 C10_N_btm.n2472 C10_N_btm.n2471 0.6255
R41160 C10_N_btm.n2475 C10_N_btm.n2474 0.6255
R41161 C10_N_btm.n2478 C10_N_btm.n2477 0.6255
R41162 C10_N_btm.n2481 C10_N_btm.n2480 0.6255
R41163 C10_N_btm.n2484 C10_N_btm.n2483 0.6255
R41164 C10_N_btm.n2487 C10_N_btm.n2486 0.6255
R41165 C10_N_btm.n2490 C10_N_btm.n2489 0.6255
R41166 C10_N_btm.n2493 C10_N_btm.n2492 0.6255
R41167 C10_N_btm.n2496 C10_N_btm.n2495 0.6255
R41168 C10_N_btm.n2499 C10_N_btm.n2498 0.6255
R41169 C10_N_btm.n2502 C10_N_btm.n2501 0.6255
R41170 C10_N_btm.n2505 C10_N_btm.n2504 0.6255
R41171 C10_N_btm.n2508 C10_N_btm.n2507 0.6255
R41172 C10_N_btm.n2511 C10_N_btm.n2510 0.6255
R41173 C10_N_btm.n2514 C10_N_btm.n2513 0.6255
R41174 C10_N_btm.n2517 C10_N_btm.n2516 0.6255
R41175 C10_N_btm.n2520 C10_N_btm.n2519 0.6255
R41176 C10_N_btm.n2523 C10_N_btm.n2522 0.6255
R41177 C10_N_btm.n2155 C10_N_btm.n2032 0.6255
R41178 C10_N_btm.n2158 C10_N_btm.n2157 0.6255
R41179 C10_N_btm.n2161 C10_N_btm.n2160 0.6255
R41180 C10_N_btm.n2164 C10_N_btm.n2163 0.6255
R41181 C10_N_btm.n2167 C10_N_btm.n2166 0.6255
R41182 C10_N_btm.n2170 C10_N_btm.n2169 0.6255
R41183 C10_N_btm.n2173 C10_N_btm.n2172 0.6255
R41184 C10_N_btm.n2176 C10_N_btm.n2175 0.6255
R41185 C10_N_btm.n2179 C10_N_btm.n2178 0.6255
R41186 C10_N_btm.n2182 C10_N_btm.n2181 0.6255
R41187 C10_N_btm.n2185 C10_N_btm.n2184 0.6255
R41188 C10_N_btm.n2188 C10_N_btm.n2187 0.6255
R41189 C10_N_btm.n2191 C10_N_btm.n2190 0.6255
R41190 C10_N_btm.n2194 C10_N_btm.n2193 0.6255
R41191 C10_N_btm.n2197 C10_N_btm.n2196 0.6255
R41192 C10_N_btm.n2200 C10_N_btm.n2199 0.6255
R41193 C10_N_btm.n2203 C10_N_btm.n2202 0.6255
R41194 C10_N_btm.n2206 C10_N_btm.n2205 0.6255
R41195 C10_N_btm.n2209 C10_N_btm.n2208 0.6255
R41196 C10_N_btm.n2212 C10_N_btm.n2211 0.6255
R41197 C10_N_btm.n2215 C10_N_btm.n2214 0.6255
R41198 C10_N_btm.n2218 C10_N_btm.n2217 0.6255
R41199 C10_N_btm.n2221 C10_N_btm.n2220 0.6255
R41200 C10_N_btm.n2224 C10_N_btm.n2223 0.6255
R41201 C10_N_btm.n2227 C10_N_btm.n2226 0.6255
R41202 C10_N_btm.n2230 C10_N_btm.n2229 0.6255
R41203 C10_N_btm.n2233 C10_N_btm.n2232 0.6255
R41204 C10_N_btm.n2236 C10_N_btm.n2235 0.6255
R41205 C10_N_btm.n2239 C10_N_btm.n2238 0.6255
R41206 C10_N_btm.n2242 C10_N_btm.n2241 0.6255
R41207 C10_N_btm.n2245 C10_N_btm.n2244 0.6255
R41208 C10_N_btm.n2248 C10_N_btm.n2247 0.6255
R41209 C10_N_btm.n2251 C10_N_btm.n2250 0.6255
R41210 C10_N_btm.n2254 C10_N_btm.n2253 0.6255
R41211 C10_N_btm.n2257 C10_N_btm.n2256 0.6255
R41212 C10_N_btm.n2260 C10_N_btm.n2259 0.6255
R41213 C10_N_btm.n2263 C10_N_btm.n2262 0.6255
R41214 C10_N_btm.n2266 C10_N_btm.n2265 0.6255
R41215 C10_N_btm.n2269 C10_N_btm.n2268 0.6255
R41216 C10_N_btm.n2272 C10_N_btm.n2271 0.6255
R41217 C10_N_btm.n2275 C10_N_btm.n2274 0.6255
R41218 C10_N_btm.n2278 C10_N_btm.n2277 0.6255
R41219 C10_N_btm.n2281 C10_N_btm.n2280 0.6255
R41220 C10_N_btm.n2284 C10_N_btm.n2283 0.6255
R41221 C10_N_btm.n2287 C10_N_btm.n2286 0.6255
R41222 C10_N_btm.n2290 C10_N_btm.n2289 0.6255
R41223 C10_N_btm.n2293 C10_N_btm.n2292 0.6255
R41224 C10_N_btm.n2296 C10_N_btm.n2295 0.6255
R41225 C10_N_btm.n2299 C10_N_btm.n2298 0.6255
R41226 C10_N_btm.n2302 C10_N_btm.n2301 0.6255
R41227 C10_N_btm.n2305 C10_N_btm.n2304 0.6255
R41228 C10_N_btm.n2308 C10_N_btm.n2307 0.6255
R41229 C10_N_btm.n2311 C10_N_btm.n2310 0.6255
R41230 C10_N_btm.n2314 C10_N_btm.n2313 0.6255
R41231 C10_N_btm.n2317 C10_N_btm.n2316 0.6255
R41232 C10_N_btm.n2320 C10_N_btm.n2319 0.6255
R41233 C10_N_btm.n2323 C10_N_btm.n2322 0.6255
R41234 C10_N_btm.n2326 C10_N_btm.n2325 0.6255
R41235 C10_N_btm.n2329 C10_N_btm.n2328 0.6255
R41236 C10_N_btm.n2332 C10_N_btm.n2331 0.6255
R41237 C10_N_btm.n2336 C10_N_btm.n2334 0.6255
R41238 C10_N_btm.n2717 C10_N_btm.n2716 0.6255
R41239 C10_N_btm.n2714 C10_N_btm.n2713 0.6255
R41240 C10_N_btm.n2711 C10_N_btm.n2710 0.6255
R41241 C10_N_btm.n2708 C10_N_btm.n2707 0.6255
R41242 C10_N_btm.n2705 C10_N_btm.n2704 0.6255
R41243 C10_N_btm.n2702 C10_N_btm.n2701 0.6255
R41244 C10_N_btm.n2699 C10_N_btm.n2698 0.6255
R41245 C10_N_btm.n2696 C10_N_btm.n2695 0.6255
R41246 C10_N_btm.n2693 C10_N_btm.n2692 0.6255
R41247 C10_N_btm.n2690 C10_N_btm.n2689 0.6255
R41248 C10_N_btm.n2687 C10_N_btm.n2686 0.6255
R41249 C10_N_btm.n2684 C10_N_btm.n2683 0.6255
R41250 C10_N_btm.n2681 C10_N_btm.n2680 0.6255
R41251 C10_N_btm.n2678 C10_N_btm.n2677 0.6255
R41252 C10_N_btm.n2675 C10_N_btm.n2674 0.6255
R41253 C10_N_btm.n2672 C10_N_btm.n2671 0.6255
R41254 C10_N_btm.n2669 C10_N_btm.n2668 0.6255
R41255 C10_N_btm.n2666 C10_N_btm.n2665 0.6255
R41256 C10_N_btm.n2663 C10_N_btm.n2662 0.6255
R41257 C10_N_btm.n2660 C10_N_btm.n2659 0.6255
R41258 C10_N_btm.n2657 C10_N_btm.n2656 0.6255
R41259 C10_N_btm.n2654 C10_N_btm.n2653 0.6255
R41260 C10_N_btm.n2651 C10_N_btm.n2650 0.6255
R41261 C10_N_btm.n2648 C10_N_btm.n2647 0.6255
R41262 C10_N_btm.n2645 C10_N_btm.n2644 0.6255
R41263 C10_N_btm.n2642 C10_N_btm.n2641 0.6255
R41264 C10_N_btm.n2639 C10_N_btm.n2638 0.6255
R41265 C10_N_btm.n2636 C10_N_btm.n2635 0.6255
R41266 C10_N_btm.n2633 C10_N_btm.n2632 0.6255
R41267 C10_N_btm.n2630 C10_N_btm.n2629 0.6255
R41268 C10_N_btm.n2627 C10_N_btm.n2626 0.6255
R41269 C10_N_btm.n2624 C10_N_btm.n2623 0.6255
R41270 C10_N_btm.n2621 C10_N_btm.n2620 0.6255
R41271 C10_N_btm.n2618 C10_N_btm.n2617 0.6255
R41272 C10_N_btm.n2615 C10_N_btm.n2614 0.6255
R41273 C10_N_btm.n2612 C10_N_btm.n2611 0.6255
R41274 C10_N_btm.n2609 C10_N_btm.n2608 0.6255
R41275 C10_N_btm.n2606 C10_N_btm.n2605 0.6255
R41276 C10_N_btm.n2603 C10_N_btm.n2602 0.6255
R41277 C10_N_btm.n2600 C10_N_btm.n2599 0.6255
R41278 C10_N_btm.n2597 C10_N_btm.n2596 0.6255
R41279 C10_N_btm.n2594 C10_N_btm.n2593 0.6255
R41280 C10_N_btm.n2591 C10_N_btm.n2590 0.6255
R41281 C10_N_btm.n2588 C10_N_btm.n2587 0.6255
R41282 C10_N_btm.n2585 C10_N_btm.n2584 0.6255
R41283 C10_N_btm.n2582 C10_N_btm.n2581 0.6255
R41284 C10_N_btm.n2579 C10_N_btm.n2578 0.6255
R41285 C10_N_btm.n2576 C10_N_btm.n2575 0.6255
R41286 C10_N_btm.n2573 C10_N_btm.n2572 0.6255
R41287 C10_N_btm.n2570 C10_N_btm.n2569 0.6255
R41288 C10_N_btm.n2567 C10_N_btm.n2566 0.6255
R41289 C10_N_btm.n2564 C10_N_btm.n2563 0.6255
R41290 C10_N_btm.n2561 C10_N_btm.n2560 0.6255
R41291 C10_N_btm.n2558 C10_N_btm.n2557 0.6255
R41292 C10_N_btm.n2555 C10_N_btm.n2554 0.6255
R41293 C10_N_btm.n2552 C10_N_btm.n2551 0.6255
R41294 C10_N_btm.n2549 C10_N_btm.n2548 0.6255
R41295 C10_N_btm.n2546 C10_N_btm.n2545 0.6255
R41296 C10_N_btm.n2543 C10_N_btm.n2542 0.6255
R41297 C10_N_btm.n2540 C10_N_btm.n2539 0.6255
R41298 C10_N_btm.n2537 C10_N_btm.n2536 0.6255
R41299 C10_N_btm.n2907 C10_N_btm.n2906 0.6255
R41300 C10_N_btm.n2904 C10_N_btm.n2903 0.6255
R41301 C10_N_btm.n2901 C10_N_btm.n2900 0.6255
R41302 C10_N_btm.n2898 C10_N_btm.n2897 0.6255
R41303 C10_N_btm.n2895 C10_N_btm.n2894 0.6255
R41304 C10_N_btm.n2892 C10_N_btm.n2891 0.6255
R41305 C10_N_btm.n2889 C10_N_btm.n2888 0.6255
R41306 C10_N_btm.n2886 C10_N_btm.n2885 0.6255
R41307 C10_N_btm.n2883 C10_N_btm.n2882 0.6255
R41308 C10_N_btm.n2880 C10_N_btm.n2879 0.6255
R41309 C10_N_btm.n2877 C10_N_btm.n2876 0.6255
R41310 C10_N_btm.n2874 C10_N_btm.n2873 0.6255
R41311 C10_N_btm.n2871 C10_N_btm.n2870 0.6255
R41312 C10_N_btm.n2868 C10_N_btm.n2867 0.6255
R41313 C10_N_btm.n2865 C10_N_btm.n2864 0.6255
R41314 C10_N_btm.n2862 C10_N_btm.n2861 0.6255
R41315 C10_N_btm.n2859 C10_N_btm.n2858 0.6255
R41316 C10_N_btm.n2856 C10_N_btm.n2855 0.6255
R41317 C10_N_btm.n2853 C10_N_btm.n2852 0.6255
R41318 C10_N_btm.n2850 C10_N_btm.n2849 0.6255
R41319 C10_N_btm.n2847 C10_N_btm.n2846 0.6255
R41320 C10_N_btm.n2844 C10_N_btm.n2843 0.6255
R41321 C10_N_btm.n2841 C10_N_btm.n2840 0.6255
R41322 C10_N_btm.n2838 C10_N_btm.n2837 0.6255
R41323 C10_N_btm.n2835 C10_N_btm.n2834 0.6255
R41324 C10_N_btm.n2832 C10_N_btm.n2831 0.6255
R41325 C10_N_btm.n2829 C10_N_btm.n2828 0.6255
R41326 C10_N_btm.n2826 C10_N_btm.n2825 0.6255
R41327 C10_N_btm.n2823 C10_N_btm.n2822 0.6255
R41328 C10_N_btm.n2820 C10_N_btm.n2819 0.6255
R41329 C10_N_btm.n2817 C10_N_btm.n2816 0.6255
R41330 C10_N_btm.n2814 C10_N_btm.n2813 0.6255
R41331 C10_N_btm.n2811 C10_N_btm.n2810 0.6255
R41332 C10_N_btm.n2808 C10_N_btm.n2807 0.6255
R41333 C10_N_btm.n2805 C10_N_btm.n2804 0.6255
R41334 C10_N_btm.n2802 C10_N_btm.n2801 0.6255
R41335 C10_N_btm.n2799 C10_N_btm.n2798 0.6255
R41336 C10_N_btm.n2796 C10_N_btm.n2795 0.6255
R41337 C10_N_btm.n2793 C10_N_btm.n2792 0.6255
R41338 C10_N_btm.n2790 C10_N_btm.n2789 0.6255
R41339 C10_N_btm.n2787 C10_N_btm.n2786 0.6255
R41340 C10_N_btm.n2784 C10_N_btm.n2783 0.6255
R41341 C10_N_btm.n2781 C10_N_btm.n2780 0.6255
R41342 C10_N_btm.n2778 C10_N_btm.n2777 0.6255
R41343 C10_N_btm.n2775 C10_N_btm.n2774 0.6255
R41344 C10_N_btm.n2772 C10_N_btm.n2771 0.6255
R41345 C10_N_btm.n2769 C10_N_btm.n2768 0.6255
R41346 C10_N_btm.n2766 C10_N_btm.n2765 0.6255
R41347 C10_N_btm.n2763 C10_N_btm.n2762 0.6255
R41348 C10_N_btm.n2760 C10_N_btm.n2759 0.6255
R41349 C10_N_btm.n2757 C10_N_btm.n2756 0.6255
R41350 C10_N_btm.n2754 C10_N_btm.n2753 0.6255
R41351 C10_N_btm.n2751 C10_N_btm.n2750 0.6255
R41352 C10_N_btm.n2748 C10_N_btm.n2747 0.6255
R41353 C10_N_btm.n2745 C10_N_btm.n2744 0.6255
R41354 C10_N_btm.n2742 C10_N_btm.n2741 0.6255
R41355 C10_N_btm.n2739 C10_N_btm.n2738 0.6255
R41356 C10_N_btm.n2736 C10_N_btm.n2735 0.6255
R41357 C10_N_btm.n2733 C10_N_btm.n2732 0.6255
R41358 C10_N_btm.n2730 C10_N_btm.n2729 0.6255
R41359 C10_N_btm.n2727 C10_N_btm.n2726 0.6255
R41360 C10_N_btm.n1966 C10_N_btm.n1964 0.6255
R41361 C10_N_btm.n1962 C10_N_btm.n1961 0.6255
R41362 C10_N_btm.n1959 C10_N_btm.n1958 0.6255
R41363 C10_N_btm.n1956 C10_N_btm.n1955 0.6255
R41364 C10_N_btm.n1953 C10_N_btm.n1952 0.6255
R41365 C10_N_btm.n1950 C10_N_btm.n1949 0.6255
R41366 C10_N_btm.n1947 C10_N_btm.n1946 0.6255
R41367 C10_N_btm.n1944 C10_N_btm.n1943 0.6255
R41368 C10_N_btm.n1941 C10_N_btm.n1940 0.6255
R41369 C10_N_btm.n1938 C10_N_btm.n1937 0.6255
R41370 C10_N_btm.n1935 C10_N_btm.n1934 0.6255
R41371 C10_N_btm.n1932 C10_N_btm.n1931 0.6255
R41372 C10_N_btm.n1929 C10_N_btm.n1928 0.6255
R41373 C10_N_btm.n1926 C10_N_btm.n1925 0.6255
R41374 C10_N_btm.n1923 C10_N_btm.n1922 0.6255
R41375 C10_N_btm.n1920 C10_N_btm.n1919 0.6255
R41376 C10_N_btm.n1917 C10_N_btm.n1916 0.6255
R41377 C10_N_btm.n1914 C10_N_btm.n1913 0.6255
R41378 C10_N_btm.n1911 C10_N_btm.n1910 0.6255
R41379 C10_N_btm.n1908 C10_N_btm.n1907 0.6255
R41380 C10_N_btm.n1905 C10_N_btm.n1904 0.6255
R41381 C10_N_btm.n1902 C10_N_btm.n1901 0.6255
R41382 C10_N_btm.n1899 C10_N_btm.n1898 0.6255
R41383 C10_N_btm.n1896 C10_N_btm.n1895 0.6255
R41384 C10_N_btm.n1893 C10_N_btm.n1892 0.6255
R41385 C10_N_btm.n1890 C10_N_btm.n1889 0.6255
R41386 C10_N_btm.n1887 C10_N_btm.n1886 0.6255
R41387 C10_N_btm.n1884 C10_N_btm.n1883 0.6255
R41388 C10_N_btm.n1881 C10_N_btm.n1880 0.6255
R41389 C10_N_btm.n1878 C10_N_btm.n1877 0.6255
R41390 C10_N_btm.n1875 C10_N_btm.n1874 0.6255
R41391 C10_N_btm.n1872 C10_N_btm.n1871 0.6255
R41392 C10_N_btm.n1869 C10_N_btm.n1868 0.6255
R41393 C10_N_btm.n1866 C10_N_btm.n1865 0.6255
R41394 C10_N_btm.n1863 C10_N_btm.n1862 0.6255
R41395 C10_N_btm.n1860 C10_N_btm.n1859 0.6255
R41396 C10_N_btm.n1857 C10_N_btm.n1856 0.6255
R41397 C10_N_btm.n1854 C10_N_btm.n1853 0.6255
R41398 C10_N_btm.n1851 C10_N_btm.n1850 0.6255
R41399 C10_N_btm.n1848 C10_N_btm.n1847 0.6255
R41400 C10_N_btm.n1845 C10_N_btm.n1844 0.6255
R41401 C10_N_btm.n1842 C10_N_btm.n1841 0.6255
R41402 C10_N_btm.n1839 C10_N_btm.n1838 0.6255
R41403 C10_N_btm.n1836 C10_N_btm.n1835 0.6255
R41404 C10_N_btm.n1833 C10_N_btm.n1832 0.6255
R41405 C10_N_btm.n1830 C10_N_btm.n1829 0.6255
R41406 C10_N_btm.n1827 C10_N_btm.n1826 0.6255
R41407 C10_N_btm.n1824 C10_N_btm.n1823 0.6255
R41408 C10_N_btm.n1821 C10_N_btm.n1820 0.6255
R41409 C10_N_btm.n1818 C10_N_btm.n1817 0.6255
R41410 C10_N_btm.n1815 C10_N_btm.n1814 0.6255
R41411 C10_N_btm.n1812 C10_N_btm.n1811 0.6255
R41412 C10_N_btm.n1809 C10_N_btm.n1808 0.6255
R41413 C10_N_btm.n1806 C10_N_btm.n1805 0.6255
R41414 C10_N_btm.n1803 C10_N_btm.n1802 0.6255
R41415 C10_N_btm.n1800 C10_N_btm.n1799 0.6255
R41416 C10_N_btm.n1797 C10_N_btm.n1796 0.6255
R41417 C10_N_btm.n1794 C10_N_btm.n1793 0.6255
R41418 C10_N_btm.n1791 C10_N_btm.n1790 0.6255
R41419 C10_N_btm.n1788 C10_N_btm.n1787 0.6255
R41420 C10_N_btm.n1785 C10_N_btm.n1661 0.6255
R41421 C10_N_btm.n2922 C10_N_btm.n2921 0.6255
R41422 C10_N_btm.n2925 C10_N_btm.n2924 0.6255
R41423 C10_N_btm.n2928 C10_N_btm.n2927 0.6255
R41424 C10_N_btm.n2931 C10_N_btm.n2930 0.6255
R41425 C10_N_btm.n2934 C10_N_btm.n2933 0.6255
R41426 C10_N_btm.n2937 C10_N_btm.n2936 0.6255
R41427 C10_N_btm.n2940 C10_N_btm.n2939 0.6255
R41428 C10_N_btm.n2943 C10_N_btm.n2942 0.6255
R41429 C10_N_btm.n2946 C10_N_btm.n2945 0.6255
R41430 C10_N_btm.n2949 C10_N_btm.n2948 0.6255
R41431 C10_N_btm.n2952 C10_N_btm.n2951 0.6255
R41432 C10_N_btm.n2955 C10_N_btm.n2954 0.6255
R41433 C10_N_btm.n2958 C10_N_btm.n2957 0.6255
R41434 C10_N_btm.n2961 C10_N_btm.n2960 0.6255
R41435 C10_N_btm.n2964 C10_N_btm.n2963 0.6255
R41436 C10_N_btm.n2967 C10_N_btm.n2966 0.6255
R41437 C10_N_btm.n2970 C10_N_btm.n2969 0.6255
R41438 C10_N_btm.n2973 C10_N_btm.n2972 0.6255
R41439 C10_N_btm.n2976 C10_N_btm.n2975 0.6255
R41440 C10_N_btm.n2979 C10_N_btm.n2978 0.6255
R41441 C10_N_btm.n2982 C10_N_btm.n2981 0.6255
R41442 C10_N_btm.n2985 C10_N_btm.n2984 0.6255
R41443 C10_N_btm.n2988 C10_N_btm.n2987 0.6255
R41444 C10_N_btm.n2991 C10_N_btm.n2990 0.6255
R41445 C10_N_btm.n2994 C10_N_btm.n2993 0.6255
R41446 C10_N_btm.n2997 C10_N_btm.n2996 0.6255
R41447 C10_N_btm.n3000 C10_N_btm.n2999 0.6255
R41448 C10_N_btm.n3003 C10_N_btm.n3002 0.6255
R41449 C10_N_btm.n3006 C10_N_btm.n3005 0.6255
R41450 C10_N_btm.n3009 C10_N_btm.n3008 0.6255
R41451 C10_N_btm.n3012 C10_N_btm.n3011 0.6255
R41452 C10_N_btm.n3015 C10_N_btm.n3014 0.6255
R41453 C10_N_btm.n3018 C10_N_btm.n3017 0.6255
R41454 C10_N_btm.n3021 C10_N_btm.n3020 0.6255
R41455 C10_N_btm.n3024 C10_N_btm.n3023 0.6255
R41456 C10_N_btm.n3027 C10_N_btm.n3026 0.6255
R41457 C10_N_btm.n3030 C10_N_btm.n3029 0.6255
R41458 C10_N_btm.n3033 C10_N_btm.n3032 0.6255
R41459 C10_N_btm.n3036 C10_N_btm.n3035 0.6255
R41460 C10_N_btm.n3039 C10_N_btm.n3038 0.6255
R41461 C10_N_btm.n3042 C10_N_btm.n3041 0.6255
R41462 C10_N_btm.n3045 C10_N_btm.n3044 0.6255
R41463 C10_N_btm.n3048 C10_N_btm.n3047 0.6255
R41464 C10_N_btm.n3051 C10_N_btm.n3050 0.6255
R41465 C10_N_btm.n3054 C10_N_btm.n3053 0.6255
R41466 C10_N_btm.n3057 C10_N_btm.n3056 0.6255
R41467 C10_N_btm.n3060 C10_N_btm.n3059 0.6255
R41468 C10_N_btm.n3063 C10_N_btm.n3062 0.6255
R41469 C10_N_btm.n3066 C10_N_btm.n3065 0.6255
R41470 C10_N_btm.n3069 C10_N_btm.n3068 0.6255
R41471 C10_N_btm.n3072 C10_N_btm.n3071 0.6255
R41472 C10_N_btm.n3075 C10_N_btm.n3074 0.6255
R41473 C10_N_btm.n3078 C10_N_btm.n3077 0.6255
R41474 C10_N_btm.n3081 C10_N_btm.n3080 0.6255
R41475 C10_N_btm.n3084 C10_N_btm.n3083 0.6255
R41476 C10_N_btm.n3087 C10_N_btm.n3086 0.6255
R41477 C10_N_btm.n3090 C10_N_btm.n3089 0.6255
R41478 C10_N_btm.n3093 C10_N_btm.n3092 0.6255
R41479 C10_N_btm.n3096 C10_N_btm.n3095 0.6255
R41480 C10_N_btm.n3099 C10_N_btm.n3098 0.6255
R41481 C10_N_btm.n3102 C10_N_btm.n3101 0.6255
R41482 C10_N_btm.n946 C10_N_btm.n945 0.6255
R41483 C10_N_btm.n943 C10_N_btm.n942 0.6255
R41484 C10_N_btm.n940 C10_N_btm.n939 0.6255
R41485 C10_N_btm.n937 C10_N_btm.n936 0.6255
R41486 C10_N_btm.n934 C10_N_btm.n933 0.6255
R41487 C10_N_btm.n931 C10_N_btm.n930 0.6255
R41488 C10_N_btm.n928 C10_N_btm.n927 0.6255
R41489 C10_N_btm.n925 C10_N_btm.n924 0.6255
R41490 C10_N_btm.n978 C10_N_btm.n977 0.6255
R41491 C10_N_btm.n975 C10_N_btm.n974 0.6255
R41492 C10_N_btm.n972 C10_N_btm.n971 0.6255
R41493 C10_N_btm.n969 C10_N_btm.n968 0.6255
R41494 C10_N_btm.n966 C10_N_btm.n965 0.6255
R41495 C10_N_btm.n963 C10_N_btm.n962 0.6255
R41496 C10_N_btm.n960 C10_N_btm.n959 0.6255
R41497 C10_N_btm.n957 C10_N_btm.n956 0.6255
R41498 C10_N_btm.n1009 C10_N_btm.n1008 0.6255
R41499 C10_N_btm.n1006 C10_N_btm.n1005 0.6255
R41500 C10_N_btm.n1003 C10_N_btm.n1002 0.6255
R41501 C10_N_btm.n1000 C10_N_btm.n999 0.6255
R41502 C10_N_btm.n997 C10_N_btm.n996 0.6255
R41503 C10_N_btm.n994 C10_N_btm.n993 0.6255
R41504 C10_N_btm.n991 C10_N_btm.n990 0.6255
R41505 C10_N_btm.n988 C10_N_btm.n987 0.6255
R41506 C10_N_btm.n901 C10_N_btm.n899 0.6255
R41507 C10_N_btm.n897 C10_N_btm.n896 0.6255
R41508 C10_N_btm.n894 C10_N_btm.n893 0.6255
R41509 C10_N_btm.n891 C10_N_btm.n890 0.6255
R41510 C10_N_btm.n888 C10_N_btm.n887 0.6255
R41511 C10_N_btm.n885 C10_N_btm.n884 0.6255
R41512 C10_N_btm.n882 C10_N_btm.n881 0.6255
R41513 C10_N_btm.n879 C10_N_btm.n861 0.6255
R41514 C10_N_btm.n1024 C10_N_btm.n1023 0.6255
R41515 C10_N_btm.n1027 C10_N_btm.n1026 0.6255
R41516 C10_N_btm.n1030 C10_N_btm.n1029 0.6255
R41517 C10_N_btm.n1033 C10_N_btm.n1032 0.6255
R41518 C10_N_btm.n1036 C10_N_btm.n1035 0.6255
R41519 C10_N_btm.n1039 C10_N_btm.n1038 0.6255
R41520 C10_N_btm.n1042 C10_N_btm.n1041 0.6255
R41521 C10_N_btm.n1045 C10_N_btm.n1044 0.6255
R41522 C10_N_btm.n1055 C10_N_btm.n1054 0.6255
R41523 C10_N_btm.n1058 C10_N_btm.n1057 0.6255
R41524 C10_N_btm.n1061 C10_N_btm.n1060 0.6255
R41525 C10_N_btm.n1064 C10_N_btm.n1063 0.6255
R41526 C10_N_btm.n1067 C10_N_btm.n1066 0.6255
R41527 C10_N_btm.n1070 C10_N_btm.n1069 0.6255
R41528 C10_N_btm.n1073 C10_N_btm.n1072 0.6255
R41529 C10_N_btm.n1076 C10_N_btm.n1075 0.6255
R41530 C10_N_btm.n826 C10_N_btm.n808 0.6255
R41531 C10_N_btm.n829 C10_N_btm.n828 0.6255
R41532 C10_N_btm.n832 C10_N_btm.n831 0.6255
R41533 C10_N_btm.n835 C10_N_btm.n834 0.6255
R41534 C10_N_btm.n838 C10_N_btm.n837 0.6255
R41535 C10_N_btm.n841 C10_N_btm.n840 0.6255
R41536 C10_N_btm.n844 C10_N_btm.n843 0.6255
R41537 C10_N_btm.n848 C10_N_btm.n846 0.6255
R41538 C10_N_btm.n1112 C10_N_btm.n1111 0.6255
R41539 C10_N_btm.n1109 C10_N_btm.n1108 0.6255
R41540 C10_N_btm.n1106 C10_N_btm.n1105 0.6255
R41541 C10_N_btm.n1103 C10_N_btm.n1102 0.6255
R41542 C10_N_btm.n1100 C10_N_btm.n1099 0.6255
R41543 C10_N_btm.n1097 C10_N_btm.n1096 0.6255
R41544 C10_N_btm.n1094 C10_N_btm.n1093 0.6255
R41545 C10_N_btm.n1091 C10_N_btm.n1090 0.6255
R41546 C10_N_btm.n1143 C10_N_btm.n1142 0.6255
R41547 C10_N_btm.n1140 C10_N_btm.n1139 0.6255
R41548 C10_N_btm.n1137 C10_N_btm.n1136 0.6255
R41549 C10_N_btm.n1134 C10_N_btm.n1133 0.6255
R41550 C10_N_btm.n1131 C10_N_btm.n1130 0.6255
R41551 C10_N_btm.n1128 C10_N_btm.n1127 0.6255
R41552 C10_N_btm.n1125 C10_N_btm.n1124 0.6255
R41553 C10_N_btm.n1122 C10_N_btm.n1121 0.6255
R41554 C10_N_btm.n795 C10_N_btm.n793 0.6255
R41555 C10_N_btm.n791 C10_N_btm.n790 0.6255
R41556 C10_N_btm.n788 C10_N_btm.n787 0.6255
R41557 C10_N_btm.n785 C10_N_btm.n784 0.6255
R41558 C10_N_btm.n782 C10_N_btm.n781 0.6255
R41559 C10_N_btm.n779 C10_N_btm.n778 0.6255
R41560 C10_N_btm.n776 C10_N_btm.n775 0.6255
R41561 C10_N_btm.n773 C10_N_btm.n755 0.6255
R41562 C10_N_btm.n1158 C10_N_btm.n1157 0.6255
R41563 C10_N_btm.n1161 C10_N_btm.n1160 0.6255
R41564 C10_N_btm.n1164 C10_N_btm.n1163 0.6255
R41565 C10_N_btm.n1167 C10_N_btm.n1166 0.6255
R41566 C10_N_btm.n1170 C10_N_btm.n1169 0.6255
R41567 C10_N_btm.n1173 C10_N_btm.n1172 0.6255
R41568 C10_N_btm.n1176 C10_N_btm.n1175 0.6255
R41569 C10_N_btm.n1179 C10_N_btm.n1178 0.6255
R41570 C10_N_btm.n1189 C10_N_btm.n1188 0.6255
R41571 C10_N_btm.n1192 C10_N_btm.n1191 0.6255
R41572 C10_N_btm.n1195 C10_N_btm.n1194 0.6255
R41573 C10_N_btm.n1198 C10_N_btm.n1197 0.6255
R41574 C10_N_btm.n1201 C10_N_btm.n1200 0.6255
R41575 C10_N_btm.n1204 C10_N_btm.n1203 0.6255
R41576 C10_N_btm.n1207 C10_N_btm.n1206 0.6255
R41577 C10_N_btm.n1210 C10_N_btm.n1209 0.6255
R41578 C10_N_btm.n720 C10_N_btm.n702 0.6255
R41579 C10_N_btm.n723 C10_N_btm.n722 0.6255
R41580 C10_N_btm.n726 C10_N_btm.n725 0.6255
R41581 C10_N_btm.n729 C10_N_btm.n728 0.6255
R41582 C10_N_btm.n732 C10_N_btm.n731 0.6255
R41583 C10_N_btm.n735 C10_N_btm.n734 0.6255
R41584 C10_N_btm.n738 C10_N_btm.n737 0.6255
R41585 C10_N_btm.n742 C10_N_btm.n740 0.6255
R41586 C10_N_btm.n1246 C10_N_btm.n1245 0.6255
R41587 C10_N_btm.n1243 C10_N_btm.n1242 0.6255
R41588 C10_N_btm.n1240 C10_N_btm.n1239 0.6255
R41589 C10_N_btm.n1237 C10_N_btm.n1236 0.6255
R41590 C10_N_btm.n1234 C10_N_btm.n1233 0.6255
R41591 C10_N_btm.n1231 C10_N_btm.n1230 0.6255
R41592 C10_N_btm.n1228 C10_N_btm.n1227 0.6255
R41593 C10_N_btm.n1225 C10_N_btm.n1224 0.6255
R41594 C10_N_btm.n1277 C10_N_btm.n1276 0.6255
R41595 C10_N_btm.n1274 C10_N_btm.n1273 0.6255
R41596 C10_N_btm.n1271 C10_N_btm.n1270 0.6255
R41597 C10_N_btm.n1268 C10_N_btm.n1267 0.6255
R41598 C10_N_btm.n1265 C10_N_btm.n1264 0.6255
R41599 C10_N_btm.n1262 C10_N_btm.n1261 0.6255
R41600 C10_N_btm.n1259 C10_N_btm.n1258 0.6255
R41601 C10_N_btm.n1256 C10_N_btm.n1255 0.6255
R41602 C10_N_btm.n689 C10_N_btm.n687 0.6255
R41603 C10_N_btm.n685 C10_N_btm.n684 0.6255
R41604 C10_N_btm.n682 C10_N_btm.n681 0.6255
R41605 C10_N_btm.n679 C10_N_btm.n678 0.6255
R41606 C10_N_btm.n676 C10_N_btm.n675 0.6255
R41607 C10_N_btm.n673 C10_N_btm.n672 0.6255
R41608 C10_N_btm.n670 C10_N_btm.n669 0.6255
R41609 C10_N_btm.n667 C10_N_btm.n649 0.6255
R41610 C10_N_btm.n1292 C10_N_btm.n1291 0.6255
R41611 C10_N_btm.n1295 C10_N_btm.n1294 0.6255
R41612 C10_N_btm.n1298 C10_N_btm.n1297 0.6255
R41613 C10_N_btm.n1301 C10_N_btm.n1300 0.6255
R41614 C10_N_btm.n1304 C10_N_btm.n1303 0.6255
R41615 C10_N_btm.n1307 C10_N_btm.n1306 0.6255
R41616 C10_N_btm.n1310 C10_N_btm.n1309 0.6255
R41617 C10_N_btm.n1313 C10_N_btm.n1312 0.6255
R41618 C10_N_btm.n1323 C10_N_btm.n1322 0.6255
R41619 C10_N_btm.n1326 C10_N_btm.n1325 0.6255
R41620 C10_N_btm.n1329 C10_N_btm.n1328 0.6255
R41621 C10_N_btm.n1332 C10_N_btm.n1331 0.6255
R41622 C10_N_btm.n1335 C10_N_btm.n1334 0.6255
R41623 C10_N_btm.n1338 C10_N_btm.n1337 0.6255
R41624 C10_N_btm.n1341 C10_N_btm.n1340 0.6255
R41625 C10_N_btm.n1344 C10_N_btm.n1343 0.6255
R41626 C10_N_btm.n614 C10_N_btm.n596 0.6255
R41627 C10_N_btm.n617 C10_N_btm.n616 0.6255
R41628 C10_N_btm.n620 C10_N_btm.n619 0.6255
R41629 C10_N_btm.n623 C10_N_btm.n622 0.6255
R41630 C10_N_btm.n626 C10_N_btm.n625 0.6255
R41631 C10_N_btm.n629 C10_N_btm.n628 0.6255
R41632 C10_N_btm.n632 C10_N_btm.n631 0.6255
R41633 C10_N_btm.n636 C10_N_btm.n634 0.6255
R41634 C10_N_btm.n1380 C10_N_btm.n1379 0.6255
R41635 C10_N_btm.n1377 C10_N_btm.n1376 0.6255
R41636 C10_N_btm.n1374 C10_N_btm.n1373 0.6255
R41637 C10_N_btm.n1371 C10_N_btm.n1370 0.6255
R41638 C10_N_btm.n1368 C10_N_btm.n1367 0.6255
R41639 C10_N_btm.n1365 C10_N_btm.n1364 0.6255
R41640 C10_N_btm.n1362 C10_N_btm.n1361 0.6255
R41641 C10_N_btm.n1359 C10_N_btm.n1358 0.6255
R41642 C10_N_btm.n1446 C10_N_btm.n1445 0.6255
R41643 C10_N_btm.n1443 C10_N_btm.n1442 0.6255
R41644 C10_N_btm.n1440 C10_N_btm.n1439 0.6255
R41645 C10_N_btm.n1437 C10_N_btm.n1436 0.6255
R41646 C10_N_btm.n1434 C10_N_btm.n1433 0.6255
R41647 C10_N_btm.n1431 C10_N_btm.n1430 0.6255
R41648 C10_N_btm.n1428 C10_N_btm.n1427 0.6255
R41649 C10_N_btm.n1425 C10_N_btm.n1424 0.6255
R41650 C10_N_btm.n1415 C10_N_btm.n1414 0.6255
R41651 C10_N_btm.n1412 C10_N_btm.n1411 0.6255
R41652 C10_N_btm.n1409 C10_N_btm.n1408 0.6255
R41653 C10_N_btm.n1406 C10_N_btm.n1405 0.6255
R41654 C10_N_btm.n1403 C10_N_btm.n1402 0.6255
R41655 C10_N_btm.n1400 C10_N_btm.n1399 0.6255
R41656 C10_N_btm.n1397 C10_N_btm.n1396 0.6255
R41657 C10_N_btm.n1394 C10_N_btm.n576 0.6255
R41658 C10_N_btm.n1461 C10_N_btm.n1460 0.6255
R41659 C10_N_btm.n1464 C10_N_btm.n1463 0.6255
R41660 C10_N_btm.n1467 C10_N_btm.n1466 0.6255
R41661 C10_N_btm.n1470 C10_N_btm.n1469 0.6255
R41662 C10_N_btm.n1473 C10_N_btm.n1472 0.6255
R41663 C10_N_btm.n1476 C10_N_btm.n1475 0.6255
R41664 C10_N_btm.n1479 C10_N_btm.n1478 0.6255
R41665 C10_N_btm.n1483 C10_N_btm.n1481 0.6255
R41666 C10_N_btm.n1490 C10_N_btm.n1489 0.6255
R41667 C10_N_btm.n1493 C10_N_btm.n1492 0.6255
R41668 C10_N_btm.n1496 C10_N_btm.n1495 0.6255
R41669 C10_N_btm.n1499 C10_N_btm.n1498 0.6255
R41670 C10_N_btm.n1502 C10_N_btm.n1501 0.6255
R41671 C10_N_btm.n1505 C10_N_btm.n1504 0.6255
R41672 C10_N_btm.n1508 C10_N_btm.n1507 0.6255
R41673 C10_N_btm.n1511 C10_N_btm.n1510 0.6255
R41674 C10_N_btm.n1533 C10_N_btm.n1532 0.6255
R41675 C10_N_btm.n1536 C10_N_btm.n1535 0.6255
R41676 C10_N_btm.n1539 C10_N_btm.n1538 0.6255
R41677 C10_N_btm.n1542 C10_N_btm.n1541 0.6255
R41678 C10_N_btm.n1545 C10_N_btm.n1544 0.6255
R41679 C10_N_btm.n1548 C10_N_btm.n1547 0.6255
R41680 C10_N_btm.n1551 C10_N_btm.n1550 0.6255
R41681 C10_N_btm.n1554 C10_N_btm.n1553 0.6255
R41682 C10_N_btm.n1557 C10_N_btm.n1556 0.6255
R41683 C10_N_btm.n1560 C10_N_btm.n1559 0.6255
R41684 C10_N_btm.n1563 C10_N_btm.n1562 0.6255
R41685 C10_N_btm.n1566 C10_N_btm.n1565 0.6255
R41686 C10_N_btm.n1569 C10_N_btm.n1568 0.6255
R41687 C10_N_btm.n1572 C10_N_btm.n1571 0.6255
R41688 C10_N_btm.n1575 C10_N_btm.n1574 0.6255
R41689 C10_N_btm.n1578 C10_N_btm.n1577 0.6255
R41690 C10_N_btm.n1581 C10_N_btm.n1580 0.6255
R41691 C10_N_btm.n1584 C10_N_btm.n1583 0.6255
R41692 C10_N_btm.n1587 C10_N_btm.n1586 0.6255
R41693 C10_N_btm.n1590 C10_N_btm.n1589 0.6255
R41694 C10_N_btm.n1593 C10_N_btm.n1592 0.6255
R41695 C10_N_btm.n3112 C10_N_btm.n3111 0.6255
R41696 C10_N_btm.n3115 C10_N_btm.n3114 0.6255
R41697 C10_N_btm.n3118 C10_N_btm.n3117 0.6255
R41698 C10_N_btm.n3121 C10_N_btm.n3120 0.6255
R41699 C10_N_btm.n3124 C10_N_btm.n3123 0.6255
R41700 C10_N_btm.n3127 C10_N_btm.n3126 0.6255
R41701 C10_N_btm.n3130 C10_N_btm.n3129 0.6255
R41702 C10_N_btm.n3133 C10_N_btm.n3132 0.6255
R41703 C10_N_btm.n3136 C10_N_btm.n3135 0.6255
R41704 C10_N_btm.n3139 C10_N_btm.n3138 0.6255
R41705 C10_N_btm.n3142 C10_N_btm.n3141 0.6255
R41706 C10_N_btm.n3145 C10_N_btm.n3144 0.6255
R41707 C10_N_btm.n3148 C10_N_btm.n3147 0.6255
R41708 C10_N_btm.n3151 C10_N_btm.n3150 0.6255
R41709 C10_N_btm.n3154 C10_N_btm.n3153 0.6255
R41710 C10_N_btm.n3157 C10_N_btm.n3156 0.6255
R41711 C10_N_btm.n3160 C10_N_btm.n3159 0.6255
R41712 C10_N_btm.n3163 C10_N_btm.n3162 0.6255
R41713 C10_N_btm.n3166 C10_N_btm.n3165 0.6255
R41714 C10_N_btm.n3169 C10_N_btm.n3168 0.6255
R41715 C10_N_btm.n3172 C10_N_btm.n3171 0.6255
R41716 C10_N_btm.n3175 C10_N_btm.n3174 0.6255
R41717 C10_N_btm.n3178 C10_N_btm.n3177 0.6255
R41718 C10_N_btm.n3181 C10_N_btm.n3180 0.6255
R41719 C10_N_btm.n3184 C10_N_btm.n3183 0.6255
R41720 C10_N_btm.n3187 C10_N_btm.n3186 0.6255
R41721 C10_N_btm.n3190 C10_N_btm.n3189 0.6255
R41722 C10_N_btm.n3193 C10_N_btm.n3192 0.6255
R41723 C10_N_btm.n3196 C10_N_btm.n3195 0.6255
R41724 C10_N_btm.n3199 C10_N_btm.n3198 0.6255
R41725 C10_N_btm.n3202 C10_N_btm.n3201 0.6255
R41726 C10_N_btm.n3205 C10_N_btm.n3204 0.6255
R41727 C10_N_btm.n3208 C10_N_btm.n3207 0.6255
R41728 C10_N_btm.n3211 C10_N_btm.n3210 0.6255
R41729 C10_N_btm.n3214 C10_N_btm.n3213 0.6255
R41730 C10_N_btm.n3217 C10_N_btm.n3216 0.6255
R41731 C10_N_btm.n3220 C10_N_btm.n3219 0.6255
R41732 C10_N_btm.n3223 C10_N_btm.n3222 0.6255
R41733 C10_N_btm.n3226 C10_N_btm.n3225 0.6255
R41734 C10_N_btm.n3229 C10_N_btm.n3228 0.6255
R41735 C10_N_btm.n3232 C10_N_btm.n3231 0.6255
R41736 C10_N_btm.n3235 C10_N_btm.n3234 0.6255
R41737 C10_N_btm.n3238 C10_N_btm.n3237 0.6255
R41738 C10_N_btm.n3241 C10_N_btm.n3240 0.6255
R41739 C10_N_btm.n3244 C10_N_btm.n3243 0.6255
R41740 C10_N_btm.n3247 C10_N_btm.n3246 0.6255
R41741 C10_N_btm.n3250 C10_N_btm.n3249 0.6255
R41742 C10_N_btm.n3253 C10_N_btm.n3252 0.6255
R41743 C10_N_btm.n3256 C10_N_btm.n3255 0.6255
R41744 C10_N_btm.n3259 C10_N_btm.n3258 0.6255
R41745 C10_N_btm.n3262 C10_N_btm.n3261 0.6255
R41746 C10_N_btm.n3265 C10_N_btm.n3264 0.6255
R41747 C10_N_btm.n3268 C10_N_btm.n3267 0.6255
R41748 C10_N_btm.n3271 C10_N_btm.n3270 0.6255
R41749 C10_N_btm.n3274 C10_N_btm.n3273 0.6255
R41750 C10_N_btm.n3277 C10_N_btm.n3276 0.6255
R41751 C10_N_btm.n3280 C10_N_btm.n3279 0.6255
R41752 C10_N_btm.n3283 C10_N_btm.n3282 0.6255
R41753 C10_N_btm.n3286 C10_N_btm.n3285 0.6255
R41754 C10_N_btm.n3289 C10_N_btm.n3288 0.6255
R41755 C10_N_btm.n3292 C10_N_btm.n3291 0.6255
R41756 C10_N_btm.n443 C10_N_btm.n400 0.6255
R41757 C10_N_btm.n446 C10_N_btm.n445 0.6255
R41758 C10_N_btm.n449 C10_N_btm.n448 0.6255
R41759 C10_N_btm.n452 C10_N_btm.n451 0.6255
R41760 C10_N_btm.n455 C10_N_btm.n454 0.6255
R41761 C10_N_btm.n458 C10_N_btm.n457 0.6255
R41762 C10_N_btm.n461 C10_N_btm.n460 0.6255
R41763 C10_N_btm.n464 C10_N_btm.n463 0.6255
R41764 C10_N_btm.n467 C10_N_btm.n466 0.6255
R41765 C10_N_btm.n3328 C10_N_btm.n3327 0.6255
R41766 C10_N_btm.n3325 C10_N_btm.n3324 0.6255
R41767 C10_N_btm.n3322 C10_N_btm.n3321 0.6255
R41768 C10_N_btm.n3319 C10_N_btm.n3318 0.6255
R41769 C10_N_btm.n3316 C10_N_btm.n3315 0.6255
R41770 C10_N_btm.n3313 C10_N_btm.n3312 0.6255
R41771 C10_N_btm.n3310 C10_N_btm.n3309 0.6255
R41772 C10_N_btm.n3307 C10_N_btm.n3306 0.6255
R41773 C10_N_btm.n3359 C10_N_btm.n3358 0.6255
R41774 C10_N_btm.n3356 C10_N_btm.n3355 0.6255
R41775 C10_N_btm.n3353 C10_N_btm.n3352 0.6255
R41776 C10_N_btm.n3350 C10_N_btm.n3349 0.6255
R41777 C10_N_btm.n3347 C10_N_btm.n3346 0.6255
R41778 C10_N_btm.n3344 C10_N_btm.n3343 0.6255
R41779 C10_N_btm.n3341 C10_N_btm.n3340 0.6255
R41780 C10_N_btm.n3338 C10_N_btm.n3337 0.6255
R41781 C10_N_btm.n387 C10_N_btm.n385 0.6255
R41782 C10_N_btm.n383 C10_N_btm.n382 0.6255
R41783 C10_N_btm.n380 C10_N_btm.n379 0.6255
R41784 C10_N_btm.n377 C10_N_btm.n376 0.6255
R41785 C10_N_btm.n374 C10_N_btm.n373 0.6255
R41786 C10_N_btm.n371 C10_N_btm.n370 0.6255
R41787 C10_N_btm.n368 C10_N_btm.n367 0.6255
R41788 C10_N_btm.n365 C10_N_btm.n347 0.6255
R41789 C10_N_btm.n3374 C10_N_btm.n3373 0.6255
R41790 C10_N_btm.n3377 C10_N_btm.n3376 0.6255
R41791 C10_N_btm.n3380 C10_N_btm.n3379 0.6255
R41792 C10_N_btm.n3383 C10_N_btm.n3382 0.6255
R41793 C10_N_btm.n3386 C10_N_btm.n3385 0.6255
R41794 C10_N_btm.n3389 C10_N_btm.n3388 0.6255
R41795 C10_N_btm.n3392 C10_N_btm.n3391 0.6255
R41796 C10_N_btm.n3395 C10_N_btm.n3394 0.6255
R41797 C10_N_btm.n3405 C10_N_btm.n3404 0.6255
R41798 C10_N_btm.n3408 C10_N_btm.n3407 0.6255
R41799 C10_N_btm.n3411 C10_N_btm.n3410 0.6255
R41800 C10_N_btm.n3414 C10_N_btm.n3413 0.6255
R41801 C10_N_btm.n3417 C10_N_btm.n3416 0.6255
R41802 C10_N_btm.n3420 C10_N_btm.n3419 0.6255
R41803 C10_N_btm.n3423 C10_N_btm.n3422 0.6255
R41804 C10_N_btm.n3426 C10_N_btm.n3425 0.6255
R41805 C10_N_btm.n312 C10_N_btm.n294 0.6255
R41806 C10_N_btm.n315 C10_N_btm.n314 0.6255
R41807 C10_N_btm.n318 C10_N_btm.n317 0.6255
R41808 C10_N_btm.n321 C10_N_btm.n320 0.6255
R41809 C10_N_btm.n324 C10_N_btm.n323 0.6255
R41810 C10_N_btm.n327 C10_N_btm.n326 0.6255
R41811 C10_N_btm.n330 C10_N_btm.n329 0.6255
R41812 C10_N_btm.n334 C10_N_btm.n332 0.6255
R41813 C10_N_btm.n3462 C10_N_btm.n3461 0.6255
R41814 C10_N_btm.n3459 C10_N_btm.n3458 0.6255
R41815 C10_N_btm.n3456 C10_N_btm.n3455 0.6255
R41816 C10_N_btm.n3453 C10_N_btm.n3452 0.6255
R41817 C10_N_btm.n3450 C10_N_btm.n3449 0.6255
R41818 C10_N_btm.n3447 C10_N_btm.n3446 0.6255
R41819 C10_N_btm.n3444 C10_N_btm.n3443 0.6255
R41820 C10_N_btm.n3441 C10_N_btm.n3440 0.6255
R41821 C10_N_btm.n3493 C10_N_btm.n3492 0.6255
R41822 C10_N_btm.n3490 C10_N_btm.n3489 0.6255
R41823 C10_N_btm.n3487 C10_N_btm.n3486 0.6255
R41824 C10_N_btm.n3484 C10_N_btm.n3483 0.6255
R41825 C10_N_btm.n3481 C10_N_btm.n3480 0.6255
R41826 C10_N_btm.n3478 C10_N_btm.n3477 0.6255
R41827 C10_N_btm.n3475 C10_N_btm.n3474 0.6255
R41828 C10_N_btm.n3472 C10_N_btm.n3471 0.6255
R41829 C10_N_btm.n281 C10_N_btm.n279 0.6255
R41830 C10_N_btm.n277 C10_N_btm.n276 0.6255
R41831 C10_N_btm.n274 C10_N_btm.n273 0.6255
R41832 C10_N_btm.n271 C10_N_btm.n270 0.6255
R41833 C10_N_btm.n268 C10_N_btm.n267 0.6255
R41834 C10_N_btm.n265 C10_N_btm.n264 0.6255
R41835 C10_N_btm.n262 C10_N_btm.n261 0.6255
R41836 C10_N_btm.n259 C10_N_btm.n241 0.6255
R41837 C10_N_btm.n3508 C10_N_btm.n3507 0.6255
R41838 C10_N_btm.n3511 C10_N_btm.n3510 0.6255
R41839 C10_N_btm.n3514 C10_N_btm.n3513 0.6255
R41840 C10_N_btm.n3517 C10_N_btm.n3516 0.6255
R41841 C10_N_btm.n3520 C10_N_btm.n3519 0.6255
R41842 C10_N_btm.n3523 C10_N_btm.n3522 0.6255
R41843 C10_N_btm.n3526 C10_N_btm.n3525 0.6255
R41844 C10_N_btm.n3529 C10_N_btm.n3528 0.6255
R41845 C10_N_btm.n3539 C10_N_btm.n3538 0.6255
R41846 C10_N_btm.n3542 C10_N_btm.n3541 0.6255
R41847 C10_N_btm.n3545 C10_N_btm.n3544 0.6255
R41848 C10_N_btm.n3548 C10_N_btm.n3547 0.6255
R41849 C10_N_btm.n3551 C10_N_btm.n3550 0.6255
R41850 C10_N_btm.n3554 C10_N_btm.n3553 0.6255
R41851 C10_N_btm.n3557 C10_N_btm.n3556 0.6255
R41852 C10_N_btm.n3560 C10_N_btm.n3559 0.6255
R41853 C10_N_btm.n206 C10_N_btm.n188 0.6255
R41854 C10_N_btm.n209 C10_N_btm.n208 0.6255
R41855 C10_N_btm.n212 C10_N_btm.n211 0.6255
R41856 C10_N_btm.n215 C10_N_btm.n214 0.6255
R41857 C10_N_btm.n218 C10_N_btm.n217 0.6255
R41858 C10_N_btm.n221 C10_N_btm.n220 0.6255
R41859 C10_N_btm.n224 C10_N_btm.n223 0.6255
R41860 C10_N_btm.n228 C10_N_btm.n226 0.6255
R41861 C10_N_btm.n3596 C10_N_btm.n3595 0.6255
R41862 C10_N_btm.n3593 C10_N_btm.n3592 0.6255
R41863 C10_N_btm.n3590 C10_N_btm.n3589 0.6255
R41864 C10_N_btm.n3587 C10_N_btm.n3586 0.6255
R41865 C10_N_btm.n3584 C10_N_btm.n3583 0.6255
R41866 C10_N_btm.n3581 C10_N_btm.n3580 0.6255
R41867 C10_N_btm.n3578 C10_N_btm.n3577 0.6255
R41868 C10_N_btm.n3575 C10_N_btm.n3574 0.6255
R41869 C10_N_btm.n3627 C10_N_btm.n3626 0.6255
R41870 C10_N_btm.n3624 C10_N_btm.n3623 0.6255
R41871 C10_N_btm.n3621 C10_N_btm.n3620 0.6255
R41872 C10_N_btm.n3618 C10_N_btm.n3617 0.6255
R41873 C10_N_btm.n3615 C10_N_btm.n3614 0.6255
R41874 C10_N_btm.n3612 C10_N_btm.n3611 0.6255
R41875 C10_N_btm.n3609 C10_N_btm.n3608 0.6255
R41876 C10_N_btm.n3606 C10_N_btm.n3605 0.6255
R41877 C10_N_btm.n175 C10_N_btm.n173 0.6255
R41878 C10_N_btm.n171 C10_N_btm.n170 0.6255
R41879 C10_N_btm.n168 C10_N_btm.n167 0.6255
R41880 C10_N_btm.n165 C10_N_btm.n164 0.6255
R41881 C10_N_btm.n162 C10_N_btm.n161 0.6255
R41882 C10_N_btm.n159 C10_N_btm.n158 0.6255
R41883 C10_N_btm.n156 C10_N_btm.n155 0.6255
R41884 C10_N_btm.n153 C10_N_btm.n135 0.6255
R41885 C10_N_btm.n3642 C10_N_btm.n3641 0.6255
R41886 C10_N_btm.n3645 C10_N_btm.n3644 0.6255
R41887 C10_N_btm.n3648 C10_N_btm.n3647 0.6255
R41888 C10_N_btm.n3651 C10_N_btm.n3650 0.6255
R41889 C10_N_btm.n3654 C10_N_btm.n3653 0.6255
R41890 C10_N_btm.n3657 C10_N_btm.n3656 0.6255
R41891 C10_N_btm.n3660 C10_N_btm.n3659 0.6255
R41892 C10_N_btm.n3663 C10_N_btm.n3662 0.6255
R41893 C10_N_btm.n3673 C10_N_btm.n3672 0.6255
R41894 C10_N_btm.n3676 C10_N_btm.n3675 0.6255
R41895 C10_N_btm.n3679 C10_N_btm.n3678 0.6255
R41896 C10_N_btm.n3682 C10_N_btm.n3681 0.6255
R41897 C10_N_btm.n3685 C10_N_btm.n3684 0.6255
R41898 C10_N_btm.n3688 C10_N_btm.n3687 0.6255
R41899 C10_N_btm.n3691 C10_N_btm.n3690 0.6255
R41900 C10_N_btm.n3694 C10_N_btm.n3693 0.6255
R41901 C10_N_btm.n100 C10_N_btm.n82 0.6255
R41902 C10_N_btm.n103 C10_N_btm.n102 0.6255
R41903 C10_N_btm.n106 C10_N_btm.n105 0.6255
R41904 C10_N_btm.n109 C10_N_btm.n108 0.6255
R41905 C10_N_btm.n112 C10_N_btm.n111 0.6255
R41906 C10_N_btm.n115 C10_N_btm.n114 0.6255
R41907 C10_N_btm.n118 C10_N_btm.n117 0.6255
R41908 C10_N_btm.n122 C10_N_btm.n120 0.6255
R41909 C10_N_btm.n3730 C10_N_btm.n3729 0.6255
R41910 C10_N_btm.n3727 C10_N_btm.n3726 0.6255
R41911 C10_N_btm.n3724 C10_N_btm.n3723 0.6255
R41912 C10_N_btm.n3721 C10_N_btm.n3720 0.6255
R41913 C10_N_btm.n3718 C10_N_btm.n3717 0.6255
R41914 C10_N_btm.n3715 C10_N_btm.n3714 0.6255
R41915 C10_N_btm.n3712 C10_N_btm.n3711 0.6255
R41916 C10_N_btm.n3709 C10_N_btm.n3708 0.6255
R41917 C10_N_btm.n3796 C10_N_btm.n3795 0.6255
R41918 C10_N_btm.n3793 C10_N_btm.n3792 0.6255
R41919 C10_N_btm.n3790 C10_N_btm.n3789 0.6255
R41920 C10_N_btm.n3787 C10_N_btm.n3786 0.6255
R41921 C10_N_btm.n3784 C10_N_btm.n3783 0.6255
R41922 C10_N_btm.n3781 C10_N_btm.n3780 0.6255
R41923 C10_N_btm.n3778 C10_N_btm.n3777 0.6255
R41924 C10_N_btm.n3775 C10_N_btm.n3774 0.6255
R41925 C10_N_btm.n3765 C10_N_btm.n3764 0.6255
R41926 C10_N_btm.n3762 C10_N_btm.n3761 0.6255
R41927 C10_N_btm.n3759 C10_N_btm.n3758 0.6255
R41928 C10_N_btm.n3756 C10_N_btm.n3755 0.6255
R41929 C10_N_btm.n3753 C10_N_btm.n3752 0.6255
R41930 C10_N_btm.n3750 C10_N_btm.n3749 0.6255
R41931 C10_N_btm.n3747 C10_N_btm.n3746 0.6255
R41932 C10_N_btm.n3744 C10_N_btm.n62 0.6255
R41933 C10_N_btm.n3811 C10_N_btm.n3810 0.6255
R41934 C10_N_btm.n3814 C10_N_btm.n3813 0.6255
R41935 C10_N_btm.n3817 C10_N_btm.n3816 0.6255
R41936 C10_N_btm.n3820 C10_N_btm.n3819 0.6255
R41937 C10_N_btm.n3823 C10_N_btm.n3822 0.6255
R41938 C10_N_btm.n3826 C10_N_btm.n3825 0.6255
R41939 C10_N_btm.n3829 C10_N_btm.n3828 0.6255
R41940 C10_N_btm.n3833 C10_N_btm.n3831 0.6255
R41941 C10_N_btm.n3840 C10_N_btm.n3839 0.6255
R41942 C10_N_btm.n3843 C10_N_btm.n3842 0.6255
R41943 C10_N_btm.n3846 C10_N_btm.n3845 0.6255
R41944 C10_N_btm.n3849 C10_N_btm.n3848 0.6255
R41945 C10_N_btm.n3852 C10_N_btm.n3851 0.6255
R41946 C10_N_btm.n3855 C10_N_btm.n3854 0.6255
R41947 C10_N_btm.n3858 C10_N_btm.n3857 0.6255
R41948 C10_N_btm.n3861 C10_N_btm.n3860 0.6255
R41949 C10_N_btm.n3871 C10_N_btm.n3870 0.6255
R41950 C10_N_btm.n3874 C10_N_btm.n3873 0.6255
R41951 C10_N_btm.n3877 C10_N_btm.n3876 0.6255
R41952 C10_N_btm.n3880 C10_N_btm.n3879 0.6255
R41953 C10_N_btm.n3883 C10_N_btm.n3882 0.6255
R41954 C10_N_btm.n3886 C10_N_btm.n3885 0.6255
R41955 C10_N_btm.n3889 C10_N_btm.n3888 0.6255
R41956 C10_N_btm.n3892 C10_N_btm.n3891 0.6255
R41957 C10_N_btm.n19 C10_N_btm.n17 0.5005
R41958 C10_N_btm.n29 C10_N_btm.n27 0.5005
R41959 C10_N_btm.n31 C10_N_btm.n29 0.484875
R41960 C10_N_btm.n21 C10_N_btm.n19 0.453625
R41961 C10_N_btm.n472 C10_N_btm.n434 0.109875
R41962 C10_N_btm.n470 C10_N_btm.n434 0.109875
R41963 C10_N_btm.n475 C10_N_btm.n433 0.109875
R41964 C10_N_btm.n473 C10_N_btm.n433 0.109875
R41965 C10_N_btm.n478 C10_N_btm.n432 0.109875
R41966 C10_N_btm.n476 C10_N_btm.n432 0.109875
R41967 C10_N_btm.n481 C10_N_btm.n431 0.109875
R41968 C10_N_btm.n479 C10_N_btm.n431 0.109875
R41969 C10_N_btm.n484 C10_N_btm.n430 0.109875
R41970 C10_N_btm.n482 C10_N_btm.n430 0.109875
R41971 C10_N_btm.n487 C10_N_btm.n429 0.109875
R41972 C10_N_btm.n485 C10_N_btm.n429 0.109875
R41973 C10_N_btm.n490 C10_N_btm.n428 0.109875
R41974 C10_N_btm.n488 C10_N_btm.n428 0.109875
R41975 C10_N_btm.n493 C10_N_btm.n427 0.109875
R41976 C10_N_btm.n491 C10_N_btm.n427 0.109875
R41977 C10_N_btm.n496 C10_N_btm.n426 0.109875
R41978 C10_N_btm.n494 C10_N_btm.n426 0.109875
R41979 C10_N_btm.n499 C10_N_btm.n425 0.109875
R41980 C10_N_btm.n497 C10_N_btm.n425 0.109875
R41981 C10_N_btm.n502 C10_N_btm.n424 0.109875
R41982 C10_N_btm.n500 C10_N_btm.n424 0.109875
R41983 C10_N_btm.n505 C10_N_btm.n423 0.109875
R41984 C10_N_btm.n503 C10_N_btm.n423 0.109875
R41985 C10_N_btm.n2340 C10_N_btm.n2338 0.109875
R41986 C10_N_btm.n2342 C10_N_btm.n2338 0.109875
R41987 C10_N_btm.n2343 C10_N_btm.n2092 0.109875
R41988 C10_N_btm.n2345 C10_N_btm.n2092 0.109875
R41989 C10_N_btm.n2346 C10_N_btm.n2091 0.109875
R41990 C10_N_btm.n2348 C10_N_btm.n2091 0.109875
R41991 C10_N_btm.n2349 C10_N_btm.n2090 0.109875
R41992 C10_N_btm.n2351 C10_N_btm.n2090 0.109875
R41993 C10_N_btm.n2352 C10_N_btm.n2089 0.109875
R41994 C10_N_btm.n2354 C10_N_btm.n2089 0.109875
R41995 C10_N_btm.n2355 C10_N_btm.n2088 0.109875
R41996 C10_N_btm.n2357 C10_N_btm.n2088 0.109875
R41997 C10_N_btm.n2358 C10_N_btm.n2087 0.109875
R41998 C10_N_btm.n2360 C10_N_btm.n2087 0.109875
R41999 C10_N_btm.n2361 C10_N_btm.n2086 0.109875
R42000 C10_N_btm.n2363 C10_N_btm.n2086 0.109875
R42001 C10_N_btm.n2364 C10_N_btm.n2085 0.109875
R42002 C10_N_btm.n2366 C10_N_btm.n2085 0.109875
R42003 C10_N_btm.n2367 C10_N_btm.n2084 0.109875
R42004 C10_N_btm.n2369 C10_N_btm.n2084 0.109875
R42005 C10_N_btm.n2370 C10_N_btm.n2083 0.109875
R42006 C10_N_btm.n2372 C10_N_btm.n2083 0.109875
R42007 C10_N_btm.n2373 C10_N_btm.n2082 0.109875
R42008 C10_N_btm.n2375 C10_N_btm.n2082 0.109875
R42009 C10_N_btm.n2376 C10_N_btm.n2081 0.109875
R42010 C10_N_btm.n2378 C10_N_btm.n2081 0.109875
R42011 C10_N_btm.n2379 C10_N_btm.n2080 0.109875
R42012 C10_N_btm.n2381 C10_N_btm.n2080 0.109875
R42013 C10_N_btm.n2382 C10_N_btm.n2079 0.109875
R42014 C10_N_btm.n2384 C10_N_btm.n2079 0.109875
R42015 C10_N_btm.n2385 C10_N_btm.n2078 0.109875
R42016 C10_N_btm.n2387 C10_N_btm.n2078 0.109875
R42017 C10_N_btm.n2388 C10_N_btm.n2077 0.109875
R42018 C10_N_btm.n2390 C10_N_btm.n2077 0.109875
R42019 C10_N_btm.n2391 C10_N_btm.n2076 0.109875
R42020 C10_N_btm.n2393 C10_N_btm.n2076 0.109875
R42021 C10_N_btm.n2394 C10_N_btm.n2075 0.109875
R42022 C10_N_btm.n2396 C10_N_btm.n2075 0.109875
R42023 C10_N_btm.n2397 C10_N_btm.n2074 0.109875
R42024 C10_N_btm.n2399 C10_N_btm.n2074 0.109875
R42025 C10_N_btm.n2400 C10_N_btm.n2073 0.109875
R42026 C10_N_btm.n2402 C10_N_btm.n2073 0.109875
R42027 C10_N_btm.n2403 C10_N_btm.n2072 0.109875
R42028 C10_N_btm.n2405 C10_N_btm.n2072 0.109875
R42029 C10_N_btm.n2406 C10_N_btm.n2071 0.109875
R42030 C10_N_btm.n2408 C10_N_btm.n2071 0.109875
R42031 C10_N_btm.n2409 C10_N_btm.n2070 0.109875
R42032 C10_N_btm.n2411 C10_N_btm.n2070 0.109875
R42033 C10_N_btm.n2412 C10_N_btm.n2069 0.109875
R42034 C10_N_btm.n2414 C10_N_btm.n2069 0.109875
R42035 C10_N_btm.n2415 C10_N_btm.n2068 0.109875
R42036 C10_N_btm.n2417 C10_N_btm.n2068 0.109875
R42037 C10_N_btm.n2418 C10_N_btm.n2067 0.109875
R42038 C10_N_btm.n2420 C10_N_btm.n2067 0.109875
R42039 C10_N_btm.n2421 C10_N_btm.n2066 0.109875
R42040 C10_N_btm.n2423 C10_N_btm.n2066 0.109875
R42041 C10_N_btm.n2424 C10_N_btm.n2065 0.109875
R42042 C10_N_btm.n2426 C10_N_btm.n2065 0.109875
R42043 C10_N_btm.n2427 C10_N_btm.n2064 0.109875
R42044 C10_N_btm.n2429 C10_N_btm.n2064 0.109875
R42045 C10_N_btm.n2430 C10_N_btm.n2063 0.109875
R42046 C10_N_btm.n2432 C10_N_btm.n2063 0.109875
R42047 C10_N_btm.n2433 C10_N_btm.n2062 0.109875
R42048 C10_N_btm.n2435 C10_N_btm.n2062 0.109875
R42049 C10_N_btm.n2436 C10_N_btm.n2061 0.109875
R42050 C10_N_btm.n2438 C10_N_btm.n2061 0.109875
R42051 C10_N_btm.n2439 C10_N_btm.n2060 0.109875
R42052 C10_N_btm.n2441 C10_N_btm.n2060 0.109875
R42053 C10_N_btm.n2442 C10_N_btm.n2059 0.109875
R42054 C10_N_btm.n2444 C10_N_btm.n2059 0.109875
R42055 C10_N_btm.n2445 C10_N_btm.n2058 0.109875
R42056 C10_N_btm.n2447 C10_N_btm.n2058 0.109875
R42057 C10_N_btm.n2448 C10_N_btm.n2057 0.109875
R42058 C10_N_btm.n2450 C10_N_btm.n2057 0.109875
R42059 C10_N_btm.n2451 C10_N_btm.n2056 0.109875
R42060 C10_N_btm.n2453 C10_N_btm.n2056 0.109875
R42061 C10_N_btm.n2454 C10_N_btm.n2055 0.109875
R42062 C10_N_btm.n2456 C10_N_btm.n2055 0.109875
R42063 C10_N_btm.n2457 C10_N_btm.n2054 0.109875
R42064 C10_N_btm.n2459 C10_N_btm.n2054 0.109875
R42065 C10_N_btm.n2460 C10_N_btm.n2053 0.109875
R42066 C10_N_btm.n2462 C10_N_btm.n2053 0.109875
R42067 C10_N_btm.n2463 C10_N_btm.n2052 0.109875
R42068 C10_N_btm.n2465 C10_N_btm.n2052 0.109875
R42069 C10_N_btm.n2466 C10_N_btm.n2051 0.109875
R42070 C10_N_btm.n2468 C10_N_btm.n2051 0.109875
R42071 C10_N_btm.n2469 C10_N_btm.n2050 0.109875
R42072 C10_N_btm.n2471 C10_N_btm.n2050 0.109875
R42073 C10_N_btm.n2472 C10_N_btm.n2049 0.109875
R42074 C10_N_btm.n2474 C10_N_btm.n2049 0.109875
R42075 C10_N_btm.n2475 C10_N_btm.n2048 0.109875
R42076 C10_N_btm.n2477 C10_N_btm.n2048 0.109875
R42077 C10_N_btm.n2478 C10_N_btm.n2047 0.109875
R42078 C10_N_btm.n2480 C10_N_btm.n2047 0.109875
R42079 C10_N_btm.n2481 C10_N_btm.n2046 0.109875
R42080 C10_N_btm.n2483 C10_N_btm.n2046 0.109875
R42081 C10_N_btm.n2484 C10_N_btm.n2045 0.109875
R42082 C10_N_btm.n2486 C10_N_btm.n2045 0.109875
R42083 C10_N_btm.n2487 C10_N_btm.n2044 0.109875
R42084 C10_N_btm.n2489 C10_N_btm.n2044 0.109875
R42085 C10_N_btm.n2490 C10_N_btm.n2043 0.109875
R42086 C10_N_btm.n2492 C10_N_btm.n2043 0.109875
R42087 C10_N_btm.n2493 C10_N_btm.n2042 0.109875
R42088 C10_N_btm.n2495 C10_N_btm.n2042 0.109875
R42089 C10_N_btm.n2496 C10_N_btm.n2041 0.109875
R42090 C10_N_btm.n2498 C10_N_btm.n2041 0.109875
R42091 C10_N_btm.n2499 C10_N_btm.n2040 0.109875
R42092 C10_N_btm.n2501 C10_N_btm.n2040 0.109875
R42093 C10_N_btm.n2502 C10_N_btm.n2039 0.109875
R42094 C10_N_btm.n2504 C10_N_btm.n2039 0.109875
R42095 C10_N_btm.n2505 C10_N_btm.n2038 0.109875
R42096 C10_N_btm.n2507 C10_N_btm.n2038 0.109875
R42097 C10_N_btm.n2508 C10_N_btm.n2037 0.109875
R42098 C10_N_btm.n2510 C10_N_btm.n2037 0.109875
R42099 C10_N_btm.n2511 C10_N_btm.n2036 0.109875
R42100 C10_N_btm.n2513 C10_N_btm.n2036 0.109875
R42101 C10_N_btm.n2514 C10_N_btm.n2035 0.109875
R42102 C10_N_btm.n2516 C10_N_btm.n2035 0.109875
R42103 C10_N_btm.n2517 C10_N_btm.n2034 0.109875
R42104 C10_N_btm.n2519 C10_N_btm.n2034 0.109875
R42105 C10_N_btm.n2520 C10_N_btm.n2033 0.109875
R42106 C10_N_btm.n2522 C10_N_btm.n2033 0.109875
R42107 C10_N_btm.n2523 C10_N_btm.n2031 0.109875
R42108 C10_N_btm.n2525 C10_N_btm.n2031 0.109875
R42109 C10_N_btm.n2531 C10_N_btm.n2032 0.109875
R42110 C10_N_btm.n2531 C10_N_btm.n2530 0.109875
R42111 C10_N_btm.n2157 C10_N_btm.n2154 0.109875
R42112 C10_N_btm.n2155 C10_N_btm.n2154 0.109875
R42113 C10_N_btm.n2160 C10_N_btm.n2153 0.109875
R42114 C10_N_btm.n2158 C10_N_btm.n2153 0.109875
R42115 C10_N_btm.n2163 C10_N_btm.n2152 0.109875
R42116 C10_N_btm.n2161 C10_N_btm.n2152 0.109875
R42117 C10_N_btm.n2166 C10_N_btm.n2151 0.109875
R42118 C10_N_btm.n2164 C10_N_btm.n2151 0.109875
R42119 C10_N_btm.n2169 C10_N_btm.n2150 0.109875
R42120 C10_N_btm.n2167 C10_N_btm.n2150 0.109875
R42121 C10_N_btm.n2172 C10_N_btm.n2149 0.109875
R42122 C10_N_btm.n2170 C10_N_btm.n2149 0.109875
R42123 C10_N_btm.n2175 C10_N_btm.n2148 0.109875
R42124 C10_N_btm.n2173 C10_N_btm.n2148 0.109875
R42125 C10_N_btm.n2178 C10_N_btm.n2147 0.109875
R42126 C10_N_btm.n2176 C10_N_btm.n2147 0.109875
R42127 C10_N_btm.n2181 C10_N_btm.n2146 0.109875
R42128 C10_N_btm.n2179 C10_N_btm.n2146 0.109875
R42129 C10_N_btm.n2184 C10_N_btm.n2145 0.109875
R42130 C10_N_btm.n2182 C10_N_btm.n2145 0.109875
R42131 C10_N_btm.n2187 C10_N_btm.n2144 0.109875
R42132 C10_N_btm.n2185 C10_N_btm.n2144 0.109875
R42133 C10_N_btm.n2190 C10_N_btm.n2143 0.109875
R42134 C10_N_btm.n2188 C10_N_btm.n2143 0.109875
R42135 C10_N_btm.n2193 C10_N_btm.n2142 0.109875
R42136 C10_N_btm.n2191 C10_N_btm.n2142 0.109875
R42137 C10_N_btm.n2196 C10_N_btm.n2141 0.109875
R42138 C10_N_btm.n2194 C10_N_btm.n2141 0.109875
R42139 C10_N_btm.n2199 C10_N_btm.n2140 0.109875
R42140 C10_N_btm.n2197 C10_N_btm.n2140 0.109875
R42141 C10_N_btm.n2202 C10_N_btm.n2139 0.109875
R42142 C10_N_btm.n2200 C10_N_btm.n2139 0.109875
R42143 C10_N_btm.n2205 C10_N_btm.n2138 0.109875
R42144 C10_N_btm.n2203 C10_N_btm.n2138 0.109875
R42145 C10_N_btm.n2208 C10_N_btm.n2137 0.109875
R42146 C10_N_btm.n2206 C10_N_btm.n2137 0.109875
R42147 C10_N_btm.n2211 C10_N_btm.n2136 0.109875
R42148 C10_N_btm.n2209 C10_N_btm.n2136 0.109875
R42149 C10_N_btm.n2214 C10_N_btm.n2135 0.109875
R42150 C10_N_btm.n2212 C10_N_btm.n2135 0.109875
R42151 C10_N_btm.n2217 C10_N_btm.n2134 0.109875
R42152 C10_N_btm.n2215 C10_N_btm.n2134 0.109875
R42153 C10_N_btm.n2220 C10_N_btm.n2133 0.109875
R42154 C10_N_btm.n2218 C10_N_btm.n2133 0.109875
R42155 C10_N_btm.n2223 C10_N_btm.n2132 0.109875
R42156 C10_N_btm.n2221 C10_N_btm.n2132 0.109875
R42157 C10_N_btm.n2226 C10_N_btm.n2131 0.109875
R42158 C10_N_btm.n2224 C10_N_btm.n2131 0.109875
R42159 C10_N_btm.n2229 C10_N_btm.n2130 0.109875
R42160 C10_N_btm.n2227 C10_N_btm.n2130 0.109875
R42161 C10_N_btm.n2232 C10_N_btm.n2129 0.109875
R42162 C10_N_btm.n2230 C10_N_btm.n2129 0.109875
R42163 C10_N_btm.n2235 C10_N_btm.n2128 0.109875
R42164 C10_N_btm.n2233 C10_N_btm.n2128 0.109875
R42165 C10_N_btm.n2238 C10_N_btm.n2127 0.109875
R42166 C10_N_btm.n2236 C10_N_btm.n2127 0.109875
R42167 C10_N_btm.n2241 C10_N_btm.n2126 0.109875
R42168 C10_N_btm.n2239 C10_N_btm.n2126 0.109875
R42169 C10_N_btm.n2244 C10_N_btm.n2125 0.109875
R42170 C10_N_btm.n2242 C10_N_btm.n2125 0.109875
R42171 C10_N_btm.n2247 C10_N_btm.n2124 0.109875
R42172 C10_N_btm.n2245 C10_N_btm.n2124 0.109875
R42173 C10_N_btm.n2250 C10_N_btm.n2123 0.109875
R42174 C10_N_btm.n2248 C10_N_btm.n2123 0.109875
R42175 C10_N_btm.n2253 C10_N_btm.n2122 0.109875
R42176 C10_N_btm.n2251 C10_N_btm.n2122 0.109875
R42177 C10_N_btm.n2256 C10_N_btm.n2121 0.109875
R42178 C10_N_btm.n2254 C10_N_btm.n2121 0.109875
R42179 C10_N_btm.n2259 C10_N_btm.n2120 0.109875
R42180 C10_N_btm.n2257 C10_N_btm.n2120 0.109875
R42181 C10_N_btm.n2262 C10_N_btm.n2119 0.109875
R42182 C10_N_btm.n2260 C10_N_btm.n2119 0.109875
R42183 C10_N_btm.n2265 C10_N_btm.n2118 0.109875
R42184 C10_N_btm.n2263 C10_N_btm.n2118 0.109875
R42185 C10_N_btm.n2268 C10_N_btm.n2117 0.109875
R42186 C10_N_btm.n2266 C10_N_btm.n2117 0.109875
R42187 C10_N_btm.n2271 C10_N_btm.n2116 0.109875
R42188 C10_N_btm.n2269 C10_N_btm.n2116 0.109875
R42189 C10_N_btm.n2274 C10_N_btm.n2115 0.109875
R42190 C10_N_btm.n2272 C10_N_btm.n2115 0.109875
R42191 C10_N_btm.n2277 C10_N_btm.n2114 0.109875
R42192 C10_N_btm.n2275 C10_N_btm.n2114 0.109875
R42193 C10_N_btm.n2280 C10_N_btm.n2113 0.109875
R42194 C10_N_btm.n2278 C10_N_btm.n2113 0.109875
R42195 C10_N_btm.n2283 C10_N_btm.n2112 0.109875
R42196 C10_N_btm.n2281 C10_N_btm.n2112 0.109875
R42197 C10_N_btm.n2286 C10_N_btm.n2111 0.109875
R42198 C10_N_btm.n2284 C10_N_btm.n2111 0.109875
R42199 C10_N_btm.n2289 C10_N_btm.n2110 0.109875
R42200 C10_N_btm.n2287 C10_N_btm.n2110 0.109875
R42201 C10_N_btm.n2292 C10_N_btm.n2109 0.109875
R42202 C10_N_btm.n2290 C10_N_btm.n2109 0.109875
R42203 C10_N_btm.n2295 C10_N_btm.n2108 0.109875
R42204 C10_N_btm.n2293 C10_N_btm.n2108 0.109875
R42205 C10_N_btm.n2298 C10_N_btm.n2107 0.109875
R42206 C10_N_btm.n2296 C10_N_btm.n2107 0.109875
R42207 C10_N_btm.n2301 C10_N_btm.n2106 0.109875
R42208 C10_N_btm.n2299 C10_N_btm.n2106 0.109875
R42209 C10_N_btm.n2304 C10_N_btm.n2105 0.109875
R42210 C10_N_btm.n2302 C10_N_btm.n2105 0.109875
R42211 C10_N_btm.n2307 C10_N_btm.n2104 0.109875
R42212 C10_N_btm.n2305 C10_N_btm.n2104 0.109875
R42213 C10_N_btm.n2310 C10_N_btm.n2103 0.109875
R42214 C10_N_btm.n2308 C10_N_btm.n2103 0.109875
R42215 C10_N_btm.n2313 C10_N_btm.n2102 0.109875
R42216 C10_N_btm.n2311 C10_N_btm.n2102 0.109875
R42217 C10_N_btm.n2316 C10_N_btm.n2101 0.109875
R42218 C10_N_btm.n2314 C10_N_btm.n2101 0.109875
R42219 C10_N_btm.n2319 C10_N_btm.n2100 0.109875
R42220 C10_N_btm.n2317 C10_N_btm.n2100 0.109875
R42221 C10_N_btm.n2322 C10_N_btm.n2099 0.109875
R42222 C10_N_btm.n2320 C10_N_btm.n2099 0.109875
R42223 C10_N_btm.n2325 C10_N_btm.n2098 0.109875
R42224 C10_N_btm.n2323 C10_N_btm.n2098 0.109875
R42225 C10_N_btm.n2328 C10_N_btm.n2097 0.109875
R42226 C10_N_btm.n2326 C10_N_btm.n2097 0.109875
R42227 C10_N_btm.n2331 C10_N_btm.n2096 0.109875
R42228 C10_N_btm.n2329 C10_N_btm.n2096 0.109875
R42229 C10_N_btm.n2334 C10_N_btm.n2095 0.109875
R42230 C10_N_btm.n2332 C10_N_btm.n2095 0.109875
R42231 C10_N_btm.n2337 C10_N_btm.n2094 0.109875
R42232 C10_N_btm.n2337 C10_N_btm.n2336 0.109875
R42233 C10_N_btm.n2719 C10_N_btm.n1970 0.109875
R42234 C10_N_btm.n2717 C10_N_btm.n1970 0.109875
R42235 C10_N_btm.n2716 C10_N_btm.n1971 0.109875
R42236 C10_N_btm.n2714 C10_N_btm.n1971 0.109875
R42237 C10_N_btm.n2713 C10_N_btm.n1972 0.109875
R42238 C10_N_btm.n2711 C10_N_btm.n1972 0.109875
R42239 C10_N_btm.n2710 C10_N_btm.n1973 0.109875
R42240 C10_N_btm.n2708 C10_N_btm.n1973 0.109875
R42241 C10_N_btm.n2707 C10_N_btm.n1974 0.109875
R42242 C10_N_btm.n2705 C10_N_btm.n1974 0.109875
R42243 C10_N_btm.n2704 C10_N_btm.n1975 0.109875
R42244 C10_N_btm.n2702 C10_N_btm.n1975 0.109875
R42245 C10_N_btm.n2701 C10_N_btm.n1976 0.109875
R42246 C10_N_btm.n2699 C10_N_btm.n1976 0.109875
R42247 C10_N_btm.n2698 C10_N_btm.n1977 0.109875
R42248 C10_N_btm.n2696 C10_N_btm.n1977 0.109875
R42249 C10_N_btm.n2695 C10_N_btm.n1978 0.109875
R42250 C10_N_btm.n2693 C10_N_btm.n1978 0.109875
R42251 C10_N_btm.n2692 C10_N_btm.n1979 0.109875
R42252 C10_N_btm.n2690 C10_N_btm.n1979 0.109875
R42253 C10_N_btm.n2689 C10_N_btm.n1980 0.109875
R42254 C10_N_btm.n2687 C10_N_btm.n1980 0.109875
R42255 C10_N_btm.n2686 C10_N_btm.n1981 0.109875
R42256 C10_N_btm.n2684 C10_N_btm.n1981 0.109875
R42257 C10_N_btm.n2683 C10_N_btm.n1982 0.109875
R42258 C10_N_btm.n2681 C10_N_btm.n1982 0.109875
R42259 C10_N_btm.n2680 C10_N_btm.n1983 0.109875
R42260 C10_N_btm.n2678 C10_N_btm.n1983 0.109875
R42261 C10_N_btm.n2677 C10_N_btm.n1984 0.109875
R42262 C10_N_btm.n2675 C10_N_btm.n1984 0.109875
R42263 C10_N_btm.n2674 C10_N_btm.n1985 0.109875
R42264 C10_N_btm.n2672 C10_N_btm.n1985 0.109875
R42265 C10_N_btm.n2671 C10_N_btm.n1986 0.109875
R42266 C10_N_btm.n2669 C10_N_btm.n1986 0.109875
R42267 C10_N_btm.n2668 C10_N_btm.n1987 0.109875
R42268 C10_N_btm.n2666 C10_N_btm.n1987 0.109875
R42269 C10_N_btm.n2665 C10_N_btm.n1988 0.109875
R42270 C10_N_btm.n2663 C10_N_btm.n1988 0.109875
R42271 C10_N_btm.n2662 C10_N_btm.n1989 0.109875
R42272 C10_N_btm.n2660 C10_N_btm.n1989 0.109875
R42273 C10_N_btm.n2659 C10_N_btm.n1990 0.109875
R42274 C10_N_btm.n2657 C10_N_btm.n1990 0.109875
R42275 C10_N_btm.n2656 C10_N_btm.n1991 0.109875
R42276 C10_N_btm.n2654 C10_N_btm.n1991 0.109875
R42277 C10_N_btm.n2653 C10_N_btm.n1992 0.109875
R42278 C10_N_btm.n2651 C10_N_btm.n1992 0.109875
R42279 C10_N_btm.n2650 C10_N_btm.n1993 0.109875
R42280 C10_N_btm.n2648 C10_N_btm.n1993 0.109875
R42281 C10_N_btm.n2647 C10_N_btm.n1994 0.109875
R42282 C10_N_btm.n2645 C10_N_btm.n1994 0.109875
R42283 C10_N_btm.n2644 C10_N_btm.n1995 0.109875
R42284 C10_N_btm.n2642 C10_N_btm.n1995 0.109875
R42285 C10_N_btm.n2641 C10_N_btm.n1996 0.109875
R42286 C10_N_btm.n2639 C10_N_btm.n1996 0.109875
R42287 C10_N_btm.n2638 C10_N_btm.n1997 0.109875
R42288 C10_N_btm.n2636 C10_N_btm.n1997 0.109875
R42289 C10_N_btm.n2635 C10_N_btm.n1998 0.109875
R42290 C10_N_btm.n2633 C10_N_btm.n1998 0.109875
R42291 C10_N_btm.n2632 C10_N_btm.n1999 0.109875
R42292 C10_N_btm.n2630 C10_N_btm.n1999 0.109875
R42293 C10_N_btm.n2629 C10_N_btm.n2000 0.109875
R42294 C10_N_btm.n2627 C10_N_btm.n2000 0.109875
R42295 C10_N_btm.n2626 C10_N_btm.n2001 0.109875
R42296 C10_N_btm.n2624 C10_N_btm.n2001 0.109875
R42297 C10_N_btm.n2623 C10_N_btm.n2002 0.109875
R42298 C10_N_btm.n2621 C10_N_btm.n2002 0.109875
R42299 C10_N_btm.n2620 C10_N_btm.n2003 0.109875
R42300 C10_N_btm.n2618 C10_N_btm.n2003 0.109875
R42301 C10_N_btm.n2617 C10_N_btm.n2004 0.109875
R42302 C10_N_btm.n2615 C10_N_btm.n2004 0.109875
R42303 C10_N_btm.n2614 C10_N_btm.n2005 0.109875
R42304 C10_N_btm.n2612 C10_N_btm.n2005 0.109875
R42305 C10_N_btm.n2611 C10_N_btm.n2006 0.109875
R42306 C10_N_btm.n2609 C10_N_btm.n2006 0.109875
R42307 C10_N_btm.n2608 C10_N_btm.n2007 0.109875
R42308 C10_N_btm.n2606 C10_N_btm.n2007 0.109875
R42309 C10_N_btm.n2605 C10_N_btm.n2008 0.109875
R42310 C10_N_btm.n2603 C10_N_btm.n2008 0.109875
R42311 C10_N_btm.n2602 C10_N_btm.n2009 0.109875
R42312 C10_N_btm.n2600 C10_N_btm.n2009 0.109875
R42313 C10_N_btm.n2599 C10_N_btm.n2010 0.109875
R42314 C10_N_btm.n2597 C10_N_btm.n2010 0.109875
R42315 C10_N_btm.n2596 C10_N_btm.n2011 0.109875
R42316 C10_N_btm.n2594 C10_N_btm.n2011 0.109875
R42317 C10_N_btm.n2593 C10_N_btm.n2012 0.109875
R42318 C10_N_btm.n2591 C10_N_btm.n2012 0.109875
R42319 C10_N_btm.n2590 C10_N_btm.n2013 0.109875
R42320 C10_N_btm.n2588 C10_N_btm.n2013 0.109875
R42321 C10_N_btm.n2587 C10_N_btm.n2014 0.109875
R42322 C10_N_btm.n2585 C10_N_btm.n2014 0.109875
R42323 C10_N_btm.n2584 C10_N_btm.n2015 0.109875
R42324 C10_N_btm.n2582 C10_N_btm.n2015 0.109875
R42325 C10_N_btm.n2581 C10_N_btm.n2016 0.109875
R42326 C10_N_btm.n2579 C10_N_btm.n2016 0.109875
R42327 C10_N_btm.n2578 C10_N_btm.n2017 0.109875
R42328 C10_N_btm.n2576 C10_N_btm.n2017 0.109875
R42329 C10_N_btm.n2575 C10_N_btm.n2018 0.109875
R42330 C10_N_btm.n2573 C10_N_btm.n2018 0.109875
R42331 C10_N_btm.n2572 C10_N_btm.n2019 0.109875
R42332 C10_N_btm.n2570 C10_N_btm.n2019 0.109875
R42333 C10_N_btm.n2569 C10_N_btm.n2020 0.109875
R42334 C10_N_btm.n2567 C10_N_btm.n2020 0.109875
R42335 C10_N_btm.n2566 C10_N_btm.n2021 0.109875
R42336 C10_N_btm.n2564 C10_N_btm.n2021 0.109875
R42337 C10_N_btm.n2563 C10_N_btm.n2022 0.109875
R42338 C10_N_btm.n2561 C10_N_btm.n2022 0.109875
R42339 C10_N_btm.n2560 C10_N_btm.n2023 0.109875
R42340 C10_N_btm.n2558 C10_N_btm.n2023 0.109875
R42341 C10_N_btm.n2557 C10_N_btm.n2024 0.109875
R42342 C10_N_btm.n2555 C10_N_btm.n2024 0.109875
R42343 C10_N_btm.n2554 C10_N_btm.n2025 0.109875
R42344 C10_N_btm.n2552 C10_N_btm.n2025 0.109875
R42345 C10_N_btm.n2551 C10_N_btm.n2026 0.109875
R42346 C10_N_btm.n2549 C10_N_btm.n2026 0.109875
R42347 C10_N_btm.n2548 C10_N_btm.n2027 0.109875
R42348 C10_N_btm.n2546 C10_N_btm.n2027 0.109875
R42349 C10_N_btm.n2545 C10_N_btm.n2028 0.109875
R42350 C10_N_btm.n2543 C10_N_btm.n2028 0.109875
R42351 C10_N_btm.n2542 C10_N_btm.n2029 0.109875
R42352 C10_N_btm.n2540 C10_N_btm.n2029 0.109875
R42353 C10_N_btm.n2539 C10_N_btm.n2030 0.109875
R42354 C10_N_btm.n2537 C10_N_btm.n2030 0.109875
R42355 C10_N_btm.n2536 C10_N_btm.n2532 0.109875
R42356 C10_N_btm.n2534 C10_N_btm.n2532 0.109875
R42357 C10_N_btm.n2907 C10_N_btm.n1660 0.109875
R42358 C10_N_btm.n2909 C10_N_btm.n1660 0.109875
R42359 C10_N_btm.n2904 C10_N_btm.n1663 0.109875
R42360 C10_N_btm.n2906 C10_N_btm.n1663 0.109875
R42361 C10_N_btm.n2901 C10_N_btm.n1664 0.109875
R42362 C10_N_btm.n2903 C10_N_btm.n1664 0.109875
R42363 C10_N_btm.n2898 C10_N_btm.n1665 0.109875
R42364 C10_N_btm.n2900 C10_N_btm.n1665 0.109875
R42365 C10_N_btm.n2895 C10_N_btm.n1666 0.109875
R42366 C10_N_btm.n2897 C10_N_btm.n1666 0.109875
R42367 C10_N_btm.n2892 C10_N_btm.n1667 0.109875
R42368 C10_N_btm.n2894 C10_N_btm.n1667 0.109875
R42369 C10_N_btm.n2889 C10_N_btm.n1668 0.109875
R42370 C10_N_btm.n2891 C10_N_btm.n1668 0.109875
R42371 C10_N_btm.n2886 C10_N_btm.n1669 0.109875
R42372 C10_N_btm.n2888 C10_N_btm.n1669 0.109875
R42373 C10_N_btm.n2883 C10_N_btm.n1670 0.109875
R42374 C10_N_btm.n2885 C10_N_btm.n1670 0.109875
R42375 C10_N_btm.n2880 C10_N_btm.n1671 0.109875
R42376 C10_N_btm.n2882 C10_N_btm.n1671 0.109875
R42377 C10_N_btm.n2877 C10_N_btm.n1672 0.109875
R42378 C10_N_btm.n2879 C10_N_btm.n1672 0.109875
R42379 C10_N_btm.n2874 C10_N_btm.n1673 0.109875
R42380 C10_N_btm.n2876 C10_N_btm.n1673 0.109875
R42381 C10_N_btm.n2871 C10_N_btm.n1674 0.109875
R42382 C10_N_btm.n2873 C10_N_btm.n1674 0.109875
R42383 C10_N_btm.n2868 C10_N_btm.n1675 0.109875
R42384 C10_N_btm.n2870 C10_N_btm.n1675 0.109875
R42385 C10_N_btm.n2865 C10_N_btm.n1676 0.109875
R42386 C10_N_btm.n2867 C10_N_btm.n1676 0.109875
R42387 C10_N_btm.n2862 C10_N_btm.n1677 0.109875
R42388 C10_N_btm.n2864 C10_N_btm.n1677 0.109875
R42389 C10_N_btm.n2859 C10_N_btm.n1678 0.109875
R42390 C10_N_btm.n2861 C10_N_btm.n1678 0.109875
R42391 C10_N_btm.n2856 C10_N_btm.n1679 0.109875
R42392 C10_N_btm.n2858 C10_N_btm.n1679 0.109875
R42393 C10_N_btm.n2853 C10_N_btm.n1680 0.109875
R42394 C10_N_btm.n2855 C10_N_btm.n1680 0.109875
R42395 C10_N_btm.n2850 C10_N_btm.n1681 0.109875
R42396 C10_N_btm.n2852 C10_N_btm.n1681 0.109875
R42397 C10_N_btm.n2847 C10_N_btm.n1682 0.109875
R42398 C10_N_btm.n2849 C10_N_btm.n1682 0.109875
R42399 C10_N_btm.n2844 C10_N_btm.n1683 0.109875
R42400 C10_N_btm.n2846 C10_N_btm.n1683 0.109875
R42401 C10_N_btm.n2841 C10_N_btm.n1684 0.109875
R42402 C10_N_btm.n2843 C10_N_btm.n1684 0.109875
R42403 C10_N_btm.n2838 C10_N_btm.n1685 0.109875
R42404 C10_N_btm.n2840 C10_N_btm.n1685 0.109875
R42405 C10_N_btm.n2835 C10_N_btm.n1686 0.109875
R42406 C10_N_btm.n2837 C10_N_btm.n1686 0.109875
R42407 C10_N_btm.n2832 C10_N_btm.n1687 0.109875
R42408 C10_N_btm.n2834 C10_N_btm.n1687 0.109875
R42409 C10_N_btm.n2829 C10_N_btm.n1688 0.109875
R42410 C10_N_btm.n2831 C10_N_btm.n1688 0.109875
R42411 C10_N_btm.n2826 C10_N_btm.n1689 0.109875
R42412 C10_N_btm.n2828 C10_N_btm.n1689 0.109875
R42413 C10_N_btm.n2823 C10_N_btm.n1690 0.109875
R42414 C10_N_btm.n2825 C10_N_btm.n1690 0.109875
R42415 C10_N_btm.n2820 C10_N_btm.n1691 0.109875
R42416 C10_N_btm.n2822 C10_N_btm.n1691 0.109875
R42417 C10_N_btm.n2817 C10_N_btm.n1692 0.109875
R42418 C10_N_btm.n2819 C10_N_btm.n1692 0.109875
R42419 C10_N_btm.n2814 C10_N_btm.n1693 0.109875
R42420 C10_N_btm.n2816 C10_N_btm.n1693 0.109875
R42421 C10_N_btm.n2811 C10_N_btm.n1694 0.109875
R42422 C10_N_btm.n2813 C10_N_btm.n1694 0.109875
R42423 C10_N_btm.n2808 C10_N_btm.n1695 0.109875
R42424 C10_N_btm.n2810 C10_N_btm.n1695 0.109875
R42425 C10_N_btm.n2805 C10_N_btm.n1696 0.109875
R42426 C10_N_btm.n2807 C10_N_btm.n1696 0.109875
R42427 C10_N_btm.n2802 C10_N_btm.n1697 0.109875
R42428 C10_N_btm.n2804 C10_N_btm.n1697 0.109875
R42429 C10_N_btm.n2799 C10_N_btm.n1698 0.109875
R42430 C10_N_btm.n2801 C10_N_btm.n1698 0.109875
R42431 C10_N_btm.n2796 C10_N_btm.n1699 0.109875
R42432 C10_N_btm.n2798 C10_N_btm.n1699 0.109875
R42433 C10_N_btm.n2793 C10_N_btm.n1700 0.109875
R42434 C10_N_btm.n2795 C10_N_btm.n1700 0.109875
R42435 C10_N_btm.n2790 C10_N_btm.n1701 0.109875
R42436 C10_N_btm.n2792 C10_N_btm.n1701 0.109875
R42437 C10_N_btm.n2787 C10_N_btm.n1702 0.109875
R42438 C10_N_btm.n2789 C10_N_btm.n1702 0.109875
R42439 C10_N_btm.n2784 C10_N_btm.n1703 0.109875
R42440 C10_N_btm.n2786 C10_N_btm.n1703 0.109875
R42441 C10_N_btm.n2781 C10_N_btm.n1704 0.109875
R42442 C10_N_btm.n2783 C10_N_btm.n1704 0.109875
R42443 C10_N_btm.n2778 C10_N_btm.n1705 0.109875
R42444 C10_N_btm.n2780 C10_N_btm.n1705 0.109875
R42445 C10_N_btm.n2775 C10_N_btm.n1706 0.109875
R42446 C10_N_btm.n2777 C10_N_btm.n1706 0.109875
R42447 C10_N_btm.n2772 C10_N_btm.n1707 0.109875
R42448 C10_N_btm.n2774 C10_N_btm.n1707 0.109875
R42449 C10_N_btm.n2769 C10_N_btm.n1708 0.109875
R42450 C10_N_btm.n2771 C10_N_btm.n1708 0.109875
R42451 C10_N_btm.n2766 C10_N_btm.n1709 0.109875
R42452 C10_N_btm.n2768 C10_N_btm.n1709 0.109875
R42453 C10_N_btm.n2763 C10_N_btm.n1710 0.109875
R42454 C10_N_btm.n2765 C10_N_btm.n1710 0.109875
R42455 C10_N_btm.n2760 C10_N_btm.n1711 0.109875
R42456 C10_N_btm.n2762 C10_N_btm.n1711 0.109875
R42457 C10_N_btm.n2757 C10_N_btm.n1712 0.109875
R42458 C10_N_btm.n2759 C10_N_btm.n1712 0.109875
R42459 C10_N_btm.n2754 C10_N_btm.n1713 0.109875
R42460 C10_N_btm.n2756 C10_N_btm.n1713 0.109875
R42461 C10_N_btm.n2751 C10_N_btm.n1714 0.109875
R42462 C10_N_btm.n2753 C10_N_btm.n1714 0.109875
R42463 C10_N_btm.n2748 C10_N_btm.n1715 0.109875
R42464 C10_N_btm.n2750 C10_N_btm.n1715 0.109875
R42465 C10_N_btm.n2745 C10_N_btm.n1716 0.109875
R42466 C10_N_btm.n2747 C10_N_btm.n1716 0.109875
R42467 C10_N_btm.n2742 C10_N_btm.n1717 0.109875
R42468 C10_N_btm.n2744 C10_N_btm.n1717 0.109875
R42469 C10_N_btm.n2739 C10_N_btm.n1718 0.109875
R42470 C10_N_btm.n2741 C10_N_btm.n1718 0.109875
R42471 C10_N_btm.n2736 C10_N_btm.n1719 0.109875
R42472 C10_N_btm.n2738 C10_N_btm.n1719 0.109875
R42473 C10_N_btm.n2733 C10_N_btm.n1720 0.109875
R42474 C10_N_btm.n2735 C10_N_btm.n1720 0.109875
R42475 C10_N_btm.n2730 C10_N_btm.n1721 0.109875
R42476 C10_N_btm.n2732 C10_N_btm.n1721 0.109875
R42477 C10_N_btm.n2727 C10_N_btm.n1722 0.109875
R42478 C10_N_btm.n2729 C10_N_btm.n1722 0.109875
R42479 C10_N_btm.n2724 C10_N_btm.n1968 0.109875
R42480 C10_N_btm.n2726 C10_N_btm.n1968 0.109875
R42481 C10_N_btm.n1967 C10_N_btm.n1724 0.109875
R42482 C10_N_btm.n1967 C10_N_btm.n1966 0.109875
R42483 C10_N_btm.n1964 C10_N_btm.n1725 0.109875
R42484 C10_N_btm.n1962 C10_N_btm.n1725 0.109875
R42485 C10_N_btm.n1961 C10_N_btm.n1726 0.109875
R42486 C10_N_btm.n1959 C10_N_btm.n1726 0.109875
R42487 C10_N_btm.n1958 C10_N_btm.n1727 0.109875
R42488 C10_N_btm.n1956 C10_N_btm.n1727 0.109875
R42489 C10_N_btm.n1955 C10_N_btm.n1728 0.109875
R42490 C10_N_btm.n1953 C10_N_btm.n1728 0.109875
R42491 C10_N_btm.n1952 C10_N_btm.n1729 0.109875
R42492 C10_N_btm.n1950 C10_N_btm.n1729 0.109875
R42493 C10_N_btm.n1949 C10_N_btm.n1730 0.109875
R42494 C10_N_btm.n1947 C10_N_btm.n1730 0.109875
R42495 C10_N_btm.n1946 C10_N_btm.n1731 0.109875
R42496 C10_N_btm.n1944 C10_N_btm.n1731 0.109875
R42497 C10_N_btm.n1943 C10_N_btm.n1732 0.109875
R42498 C10_N_btm.n1941 C10_N_btm.n1732 0.109875
R42499 C10_N_btm.n1940 C10_N_btm.n1733 0.109875
R42500 C10_N_btm.n1938 C10_N_btm.n1733 0.109875
R42501 C10_N_btm.n1937 C10_N_btm.n1734 0.109875
R42502 C10_N_btm.n1935 C10_N_btm.n1734 0.109875
R42503 C10_N_btm.n1934 C10_N_btm.n1735 0.109875
R42504 C10_N_btm.n1932 C10_N_btm.n1735 0.109875
R42505 C10_N_btm.n1931 C10_N_btm.n1736 0.109875
R42506 C10_N_btm.n1929 C10_N_btm.n1736 0.109875
R42507 C10_N_btm.n1928 C10_N_btm.n1737 0.109875
R42508 C10_N_btm.n1926 C10_N_btm.n1737 0.109875
R42509 C10_N_btm.n1925 C10_N_btm.n1738 0.109875
R42510 C10_N_btm.n1923 C10_N_btm.n1738 0.109875
R42511 C10_N_btm.n1922 C10_N_btm.n1739 0.109875
R42512 C10_N_btm.n1920 C10_N_btm.n1739 0.109875
R42513 C10_N_btm.n1919 C10_N_btm.n1740 0.109875
R42514 C10_N_btm.n1917 C10_N_btm.n1740 0.109875
R42515 C10_N_btm.n1916 C10_N_btm.n1741 0.109875
R42516 C10_N_btm.n1914 C10_N_btm.n1741 0.109875
R42517 C10_N_btm.n1913 C10_N_btm.n1742 0.109875
R42518 C10_N_btm.n1911 C10_N_btm.n1742 0.109875
R42519 C10_N_btm.n1910 C10_N_btm.n1743 0.109875
R42520 C10_N_btm.n1908 C10_N_btm.n1743 0.109875
R42521 C10_N_btm.n1907 C10_N_btm.n1744 0.109875
R42522 C10_N_btm.n1905 C10_N_btm.n1744 0.109875
R42523 C10_N_btm.n1904 C10_N_btm.n1745 0.109875
R42524 C10_N_btm.n1902 C10_N_btm.n1745 0.109875
R42525 C10_N_btm.n1901 C10_N_btm.n1746 0.109875
R42526 C10_N_btm.n1899 C10_N_btm.n1746 0.109875
R42527 C10_N_btm.n1898 C10_N_btm.n1747 0.109875
R42528 C10_N_btm.n1896 C10_N_btm.n1747 0.109875
R42529 C10_N_btm.n1895 C10_N_btm.n1748 0.109875
R42530 C10_N_btm.n1893 C10_N_btm.n1748 0.109875
R42531 C10_N_btm.n1892 C10_N_btm.n1749 0.109875
R42532 C10_N_btm.n1890 C10_N_btm.n1749 0.109875
R42533 C10_N_btm.n1889 C10_N_btm.n1750 0.109875
R42534 C10_N_btm.n1887 C10_N_btm.n1750 0.109875
R42535 C10_N_btm.n1886 C10_N_btm.n1751 0.109875
R42536 C10_N_btm.n1884 C10_N_btm.n1751 0.109875
R42537 C10_N_btm.n1883 C10_N_btm.n1752 0.109875
R42538 C10_N_btm.n1881 C10_N_btm.n1752 0.109875
R42539 C10_N_btm.n1880 C10_N_btm.n1753 0.109875
R42540 C10_N_btm.n1878 C10_N_btm.n1753 0.109875
R42541 C10_N_btm.n1877 C10_N_btm.n1754 0.109875
R42542 C10_N_btm.n1875 C10_N_btm.n1754 0.109875
R42543 C10_N_btm.n1874 C10_N_btm.n1755 0.109875
R42544 C10_N_btm.n1872 C10_N_btm.n1755 0.109875
R42545 C10_N_btm.n1871 C10_N_btm.n1756 0.109875
R42546 C10_N_btm.n1869 C10_N_btm.n1756 0.109875
R42547 C10_N_btm.n1868 C10_N_btm.n1757 0.109875
R42548 C10_N_btm.n1866 C10_N_btm.n1757 0.109875
R42549 C10_N_btm.n1865 C10_N_btm.n1758 0.109875
R42550 C10_N_btm.n1863 C10_N_btm.n1758 0.109875
R42551 C10_N_btm.n1862 C10_N_btm.n1759 0.109875
R42552 C10_N_btm.n1860 C10_N_btm.n1759 0.109875
R42553 C10_N_btm.n1859 C10_N_btm.n1760 0.109875
R42554 C10_N_btm.n1857 C10_N_btm.n1760 0.109875
R42555 C10_N_btm.n1856 C10_N_btm.n1761 0.109875
R42556 C10_N_btm.n1854 C10_N_btm.n1761 0.109875
R42557 C10_N_btm.n1853 C10_N_btm.n1762 0.109875
R42558 C10_N_btm.n1851 C10_N_btm.n1762 0.109875
R42559 C10_N_btm.n1850 C10_N_btm.n1763 0.109875
R42560 C10_N_btm.n1848 C10_N_btm.n1763 0.109875
R42561 C10_N_btm.n1847 C10_N_btm.n1764 0.109875
R42562 C10_N_btm.n1845 C10_N_btm.n1764 0.109875
R42563 C10_N_btm.n1844 C10_N_btm.n1765 0.109875
R42564 C10_N_btm.n1842 C10_N_btm.n1765 0.109875
R42565 C10_N_btm.n1841 C10_N_btm.n1766 0.109875
R42566 C10_N_btm.n1839 C10_N_btm.n1766 0.109875
R42567 C10_N_btm.n1838 C10_N_btm.n1767 0.109875
R42568 C10_N_btm.n1836 C10_N_btm.n1767 0.109875
R42569 C10_N_btm.n1835 C10_N_btm.n1768 0.109875
R42570 C10_N_btm.n1833 C10_N_btm.n1768 0.109875
R42571 C10_N_btm.n1832 C10_N_btm.n1769 0.109875
R42572 C10_N_btm.n1830 C10_N_btm.n1769 0.109875
R42573 C10_N_btm.n1829 C10_N_btm.n1770 0.109875
R42574 C10_N_btm.n1827 C10_N_btm.n1770 0.109875
R42575 C10_N_btm.n1826 C10_N_btm.n1771 0.109875
R42576 C10_N_btm.n1824 C10_N_btm.n1771 0.109875
R42577 C10_N_btm.n1823 C10_N_btm.n1772 0.109875
R42578 C10_N_btm.n1821 C10_N_btm.n1772 0.109875
R42579 C10_N_btm.n1820 C10_N_btm.n1773 0.109875
R42580 C10_N_btm.n1818 C10_N_btm.n1773 0.109875
R42581 C10_N_btm.n1817 C10_N_btm.n1774 0.109875
R42582 C10_N_btm.n1815 C10_N_btm.n1774 0.109875
R42583 C10_N_btm.n1814 C10_N_btm.n1775 0.109875
R42584 C10_N_btm.n1812 C10_N_btm.n1775 0.109875
R42585 C10_N_btm.n1811 C10_N_btm.n1776 0.109875
R42586 C10_N_btm.n1809 C10_N_btm.n1776 0.109875
R42587 C10_N_btm.n1808 C10_N_btm.n1777 0.109875
R42588 C10_N_btm.n1806 C10_N_btm.n1777 0.109875
R42589 C10_N_btm.n1805 C10_N_btm.n1778 0.109875
R42590 C10_N_btm.n1803 C10_N_btm.n1778 0.109875
R42591 C10_N_btm.n1802 C10_N_btm.n1779 0.109875
R42592 C10_N_btm.n1800 C10_N_btm.n1779 0.109875
R42593 C10_N_btm.n1799 C10_N_btm.n1780 0.109875
R42594 C10_N_btm.n1797 C10_N_btm.n1780 0.109875
R42595 C10_N_btm.n1796 C10_N_btm.n1781 0.109875
R42596 C10_N_btm.n1794 C10_N_btm.n1781 0.109875
R42597 C10_N_btm.n1793 C10_N_btm.n1782 0.109875
R42598 C10_N_btm.n1791 C10_N_btm.n1782 0.109875
R42599 C10_N_btm.n1790 C10_N_btm.n1783 0.109875
R42600 C10_N_btm.n1788 C10_N_btm.n1783 0.109875
R42601 C10_N_btm.n1787 C10_N_btm.n1784 0.109875
R42602 C10_N_btm.n1785 C10_N_btm.n1784 0.109875
R42603 C10_N_btm.n2916 C10_N_btm.n1661 0.109875
R42604 C10_N_btm.n2916 C10_N_btm.n2915 0.109875
R42605 C10_N_btm.n2921 C10_N_btm.n2917 0.109875
R42606 C10_N_btm.n2919 C10_N_btm.n2917 0.109875
R42607 C10_N_btm.n2924 C10_N_btm.n1659 0.109875
R42608 C10_N_btm.n2922 C10_N_btm.n1659 0.109875
R42609 C10_N_btm.n2927 C10_N_btm.n1658 0.109875
R42610 C10_N_btm.n2925 C10_N_btm.n1658 0.109875
R42611 C10_N_btm.n2930 C10_N_btm.n1657 0.109875
R42612 C10_N_btm.n2928 C10_N_btm.n1657 0.109875
R42613 C10_N_btm.n2933 C10_N_btm.n1656 0.109875
R42614 C10_N_btm.n2931 C10_N_btm.n1656 0.109875
R42615 C10_N_btm.n2936 C10_N_btm.n1655 0.109875
R42616 C10_N_btm.n2934 C10_N_btm.n1655 0.109875
R42617 C10_N_btm.n2939 C10_N_btm.n1654 0.109875
R42618 C10_N_btm.n2937 C10_N_btm.n1654 0.109875
R42619 C10_N_btm.n2942 C10_N_btm.n1653 0.109875
R42620 C10_N_btm.n2940 C10_N_btm.n1653 0.109875
R42621 C10_N_btm.n2945 C10_N_btm.n1652 0.109875
R42622 C10_N_btm.n2943 C10_N_btm.n1652 0.109875
R42623 C10_N_btm.n2948 C10_N_btm.n1651 0.109875
R42624 C10_N_btm.n2946 C10_N_btm.n1651 0.109875
R42625 C10_N_btm.n2951 C10_N_btm.n1650 0.109875
R42626 C10_N_btm.n2949 C10_N_btm.n1650 0.109875
R42627 C10_N_btm.n2954 C10_N_btm.n1649 0.109875
R42628 C10_N_btm.n2952 C10_N_btm.n1649 0.109875
R42629 C10_N_btm.n2957 C10_N_btm.n1648 0.109875
R42630 C10_N_btm.n2955 C10_N_btm.n1648 0.109875
R42631 C10_N_btm.n2960 C10_N_btm.n1647 0.109875
R42632 C10_N_btm.n2958 C10_N_btm.n1647 0.109875
R42633 C10_N_btm.n2963 C10_N_btm.n1646 0.109875
R42634 C10_N_btm.n2961 C10_N_btm.n1646 0.109875
R42635 C10_N_btm.n2966 C10_N_btm.n1645 0.109875
R42636 C10_N_btm.n2964 C10_N_btm.n1645 0.109875
R42637 C10_N_btm.n2969 C10_N_btm.n1644 0.109875
R42638 C10_N_btm.n2967 C10_N_btm.n1644 0.109875
R42639 C10_N_btm.n2972 C10_N_btm.n1643 0.109875
R42640 C10_N_btm.n2970 C10_N_btm.n1643 0.109875
R42641 C10_N_btm.n2975 C10_N_btm.n1642 0.109875
R42642 C10_N_btm.n2973 C10_N_btm.n1642 0.109875
R42643 C10_N_btm.n2978 C10_N_btm.n1641 0.109875
R42644 C10_N_btm.n2976 C10_N_btm.n1641 0.109875
R42645 C10_N_btm.n2981 C10_N_btm.n1640 0.109875
R42646 C10_N_btm.n2979 C10_N_btm.n1640 0.109875
R42647 C10_N_btm.n2984 C10_N_btm.n1639 0.109875
R42648 C10_N_btm.n2982 C10_N_btm.n1639 0.109875
R42649 C10_N_btm.n2987 C10_N_btm.n1638 0.109875
R42650 C10_N_btm.n2985 C10_N_btm.n1638 0.109875
R42651 C10_N_btm.n2990 C10_N_btm.n1637 0.109875
R42652 C10_N_btm.n2988 C10_N_btm.n1637 0.109875
R42653 C10_N_btm.n2993 C10_N_btm.n1636 0.109875
R42654 C10_N_btm.n2991 C10_N_btm.n1636 0.109875
R42655 C10_N_btm.n2996 C10_N_btm.n1635 0.109875
R42656 C10_N_btm.n2994 C10_N_btm.n1635 0.109875
R42657 C10_N_btm.n2999 C10_N_btm.n1634 0.109875
R42658 C10_N_btm.n2997 C10_N_btm.n1634 0.109875
R42659 C10_N_btm.n3002 C10_N_btm.n1633 0.109875
R42660 C10_N_btm.n3000 C10_N_btm.n1633 0.109875
R42661 C10_N_btm.n3005 C10_N_btm.n1632 0.109875
R42662 C10_N_btm.n3003 C10_N_btm.n1632 0.109875
R42663 C10_N_btm.n3008 C10_N_btm.n1631 0.109875
R42664 C10_N_btm.n3006 C10_N_btm.n1631 0.109875
R42665 C10_N_btm.n3011 C10_N_btm.n1630 0.109875
R42666 C10_N_btm.n3009 C10_N_btm.n1630 0.109875
R42667 C10_N_btm.n3014 C10_N_btm.n1629 0.109875
R42668 C10_N_btm.n3012 C10_N_btm.n1629 0.109875
R42669 C10_N_btm.n3017 C10_N_btm.n1628 0.109875
R42670 C10_N_btm.n3015 C10_N_btm.n1628 0.109875
R42671 C10_N_btm.n3020 C10_N_btm.n1627 0.109875
R42672 C10_N_btm.n3018 C10_N_btm.n1627 0.109875
R42673 C10_N_btm.n3023 C10_N_btm.n1626 0.109875
R42674 C10_N_btm.n3021 C10_N_btm.n1626 0.109875
R42675 C10_N_btm.n3026 C10_N_btm.n1625 0.109875
R42676 C10_N_btm.n3024 C10_N_btm.n1625 0.109875
R42677 C10_N_btm.n3029 C10_N_btm.n1624 0.109875
R42678 C10_N_btm.n3027 C10_N_btm.n1624 0.109875
R42679 C10_N_btm.n3032 C10_N_btm.n1623 0.109875
R42680 C10_N_btm.n3030 C10_N_btm.n1623 0.109875
R42681 C10_N_btm.n3035 C10_N_btm.n1622 0.109875
R42682 C10_N_btm.n3033 C10_N_btm.n1622 0.109875
R42683 C10_N_btm.n3038 C10_N_btm.n1621 0.109875
R42684 C10_N_btm.n3036 C10_N_btm.n1621 0.109875
R42685 C10_N_btm.n3041 C10_N_btm.n1620 0.109875
R42686 C10_N_btm.n3039 C10_N_btm.n1620 0.109875
R42687 C10_N_btm.n3044 C10_N_btm.n1619 0.109875
R42688 C10_N_btm.n3042 C10_N_btm.n1619 0.109875
R42689 C10_N_btm.n3047 C10_N_btm.n1618 0.109875
R42690 C10_N_btm.n3045 C10_N_btm.n1618 0.109875
R42691 C10_N_btm.n3050 C10_N_btm.n1617 0.109875
R42692 C10_N_btm.n3048 C10_N_btm.n1617 0.109875
R42693 C10_N_btm.n3053 C10_N_btm.n1616 0.109875
R42694 C10_N_btm.n3051 C10_N_btm.n1616 0.109875
R42695 C10_N_btm.n3056 C10_N_btm.n1615 0.109875
R42696 C10_N_btm.n3054 C10_N_btm.n1615 0.109875
R42697 C10_N_btm.n3059 C10_N_btm.n1614 0.109875
R42698 C10_N_btm.n3057 C10_N_btm.n1614 0.109875
R42699 C10_N_btm.n3062 C10_N_btm.n1613 0.109875
R42700 C10_N_btm.n3060 C10_N_btm.n1613 0.109875
R42701 C10_N_btm.n3065 C10_N_btm.n1612 0.109875
R42702 C10_N_btm.n3063 C10_N_btm.n1612 0.109875
R42703 C10_N_btm.n3068 C10_N_btm.n1611 0.109875
R42704 C10_N_btm.n3066 C10_N_btm.n1611 0.109875
R42705 C10_N_btm.n3071 C10_N_btm.n1610 0.109875
R42706 C10_N_btm.n3069 C10_N_btm.n1610 0.109875
R42707 C10_N_btm.n3074 C10_N_btm.n1609 0.109875
R42708 C10_N_btm.n3072 C10_N_btm.n1609 0.109875
R42709 C10_N_btm.n3077 C10_N_btm.n1608 0.109875
R42710 C10_N_btm.n3075 C10_N_btm.n1608 0.109875
R42711 C10_N_btm.n3080 C10_N_btm.n1607 0.109875
R42712 C10_N_btm.n3078 C10_N_btm.n1607 0.109875
R42713 C10_N_btm.n3083 C10_N_btm.n1606 0.109875
R42714 C10_N_btm.n3081 C10_N_btm.n1606 0.109875
R42715 C10_N_btm.n3086 C10_N_btm.n1605 0.109875
R42716 C10_N_btm.n3084 C10_N_btm.n1605 0.109875
R42717 C10_N_btm.n3089 C10_N_btm.n1604 0.109875
R42718 C10_N_btm.n3087 C10_N_btm.n1604 0.109875
R42719 C10_N_btm.n3092 C10_N_btm.n1603 0.109875
R42720 C10_N_btm.n3090 C10_N_btm.n1603 0.109875
R42721 C10_N_btm.n3095 C10_N_btm.n1602 0.109875
R42722 C10_N_btm.n3093 C10_N_btm.n1602 0.109875
R42723 C10_N_btm.n3098 C10_N_btm.n1601 0.109875
R42724 C10_N_btm.n3096 C10_N_btm.n1601 0.109875
R42725 C10_N_btm.n3101 C10_N_btm.n1600 0.109875
R42726 C10_N_btm.n3099 C10_N_btm.n1600 0.109875
R42727 C10_N_btm.n3104 C10_N_btm.n1599 0.109875
R42728 C10_N_btm.n3102 C10_N_btm.n1599 0.109875
R42729 C10_N_btm.n951 C10_N_btm.n946 0.109875
R42730 C10_N_btm.n951 C10_N_btm.n950 0.109875
R42731 C10_N_btm.n943 C10_N_btm.n913 0.109875
R42732 C10_N_btm.n945 C10_N_btm.n913 0.109875
R42733 C10_N_btm.n940 C10_N_btm.n914 0.109875
R42734 C10_N_btm.n942 C10_N_btm.n914 0.109875
R42735 C10_N_btm.n937 C10_N_btm.n915 0.109875
R42736 C10_N_btm.n939 C10_N_btm.n915 0.109875
R42737 C10_N_btm.n934 C10_N_btm.n916 0.109875
R42738 C10_N_btm.n936 C10_N_btm.n916 0.109875
R42739 C10_N_btm.n931 C10_N_btm.n917 0.109875
R42740 C10_N_btm.n933 C10_N_btm.n917 0.109875
R42741 C10_N_btm.n928 C10_N_btm.n918 0.109875
R42742 C10_N_btm.n930 C10_N_btm.n918 0.109875
R42743 C10_N_btm.n925 C10_N_btm.n919 0.109875
R42744 C10_N_btm.n927 C10_N_btm.n919 0.109875
R42745 C10_N_btm.n922 C10_N_btm.n920 0.109875
R42746 C10_N_btm.n924 C10_N_btm.n920 0.109875
R42747 C10_N_btm.n980 C10_N_btm.n905 0.109875
R42748 C10_N_btm.n978 C10_N_btm.n905 0.109875
R42749 C10_N_btm.n977 C10_N_btm.n906 0.109875
R42750 C10_N_btm.n975 C10_N_btm.n906 0.109875
R42751 C10_N_btm.n974 C10_N_btm.n907 0.109875
R42752 C10_N_btm.n972 C10_N_btm.n907 0.109875
R42753 C10_N_btm.n971 C10_N_btm.n908 0.109875
R42754 C10_N_btm.n969 C10_N_btm.n908 0.109875
R42755 C10_N_btm.n968 C10_N_btm.n909 0.109875
R42756 C10_N_btm.n966 C10_N_btm.n909 0.109875
R42757 C10_N_btm.n965 C10_N_btm.n910 0.109875
R42758 C10_N_btm.n963 C10_N_btm.n910 0.109875
R42759 C10_N_btm.n962 C10_N_btm.n911 0.109875
R42760 C10_N_btm.n960 C10_N_btm.n911 0.109875
R42761 C10_N_btm.n959 C10_N_btm.n912 0.109875
R42762 C10_N_btm.n957 C10_N_btm.n912 0.109875
R42763 C10_N_btm.n956 C10_N_btm.n952 0.109875
R42764 C10_N_btm.n954 C10_N_btm.n952 0.109875
R42765 C10_N_btm.n1009 C10_N_btm.n860 0.109875
R42766 C10_N_btm.n1011 C10_N_btm.n860 0.109875
R42767 C10_N_btm.n1006 C10_N_btm.n863 0.109875
R42768 C10_N_btm.n1008 C10_N_btm.n863 0.109875
R42769 C10_N_btm.n1003 C10_N_btm.n864 0.109875
R42770 C10_N_btm.n1005 C10_N_btm.n864 0.109875
R42771 C10_N_btm.n1000 C10_N_btm.n865 0.109875
R42772 C10_N_btm.n1002 C10_N_btm.n865 0.109875
R42773 C10_N_btm.n997 C10_N_btm.n866 0.109875
R42774 C10_N_btm.n999 C10_N_btm.n866 0.109875
R42775 C10_N_btm.n994 C10_N_btm.n867 0.109875
R42776 C10_N_btm.n996 C10_N_btm.n867 0.109875
R42777 C10_N_btm.n991 C10_N_btm.n868 0.109875
R42778 C10_N_btm.n993 C10_N_btm.n868 0.109875
R42779 C10_N_btm.n988 C10_N_btm.n869 0.109875
R42780 C10_N_btm.n990 C10_N_btm.n869 0.109875
R42781 C10_N_btm.n985 C10_N_btm.n903 0.109875
R42782 C10_N_btm.n987 C10_N_btm.n903 0.109875
R42783 C10_N_btm.n902 C10_N_btm.n871 0.109875
R42784 C10_N_btm.n902 C10_N_btm.n901 0.109875
R42785 C10_N_btm.n899 C10_N_btm.n872 0.109875
R42786 C10_N_btm.n897 C10_N_btm.n872 0.109875
R42787 C10_N_btm.n896 C10_N_btm.n873 0.109875
R42788 C10_N_btm.n894 C10_N_btm.n873 0.109875
R42789 C10_N_btm.n893 C10_N_btm.n874 0.109875
R42790 C10_N_btm.n891 C10_N_btm.n874 0.109875
R42791 C10_N_btm.n890 C10_N_btm.n875 0.109875
R42792 C10_N_btm.n888 C10_N_btm.n875 0.109875
R42793 C10_N_btm.n887 C10_N_btm.n876 0.109875
R42794 C10_N_btm.n885 C10_N_btm.n876 0.109875
R42795 C10_N_btm.n884 C10_N_btm.n877 0.109875
R42796 C10_N_btm.n882 C10_N_btm.n877 0.109875
R42797 C10_N_btm.n881 C10_N_btm.n878 0.109875
R42798 C10_N_btm.n879 C10_N_btm.n878 0.109875
R42799 C10_N_btm.n1018 C10_N_btm.n861 0.109875
R42800 C10_N_btm.n1018 C10_N_btm.n1017 0.109875
R42801 C10_N_btm.n1023 C10_N_btm.n1019 0.109875
R42802 C10_N_btm.n1021 C10_N_btm.n1019 0.109875
R42803 C10_N_btm.n1026 C10_N_btm.n859 0.109875
R42804 C10_N_btm.n1024 C10_N_btm.n859 0.109875
R42805 C10_N_btm.n1029 C10_N_btm.n858 0.109875
R42806 C10_N_btm.n1027 C10_N_btm.n858 0.109875
R42807 C10_N_btm.n1032 C10_N_btm.n857 0.109875
R42808 C10_N_btm.n1030 C10_N_btm.n857 0.109875
R42809 C10_N_btm.n1035 C10_N_btm.n856 0.109875
R42810 C10_N_btm.n1033 C10_N_btm.n856 0.109875
R42811 C10_N_btm.n1038 C10_N_btm.n855 0.109875
R42812 C10_N_btm.n1036 C10_N_btm.n855 0.109875
R42813 C10_N_btm.n1041 C10_N_btm.n854 0.109875
R42814 C10_N_btm.n1039 C10_N_btm.n854 0.109875
R42815 C10_N_btm.n1044 C10_N_btm.n853 0.109875
R42816 C10_N_btm.n1042 C10_N_btm.n853 0.109875
R42817 C10_N_btm.n1047 C10_N_btm.n852 0.109875
R42818 C10_N_btm.n1045 C10_N_btm.n852 0.109875
R42819 C10_N_btm.n1052 C10_N_btm.n850 0.109875
R42820 C10_N_btm.n1054 C10_N_btm.n850 0.109875
R42821 C10_N_btm.n1055 C10_N_btm.n816 0.109875
R42822 C10_N_btm.n1057 C10_N_btm.n816 0.109875
R42823 C10_N_btm.n1058 C10_N_btm.n815 0.109875
R42824 C10_N_btm.n1060 C10_N_btm.n815 0.109875
R42825 C10_N_btm.n1061 C10_N_btm.n814 0.109875
R42826 C10_N_btm.n1063 C10_N_btm.n814 0.109875
R42827 C10_N_btm.n1064 C10_N_btm.n813 0.109875
R42828 C10_N_btm.n1066 C10_N_btm.n813 0.109875
R42829 C10_N_btm.n1067 C10_N_btm.n812 0.109875
R42830 C10_N_btm.n1069 C10_N_btm.n812 0.109875
R42831 C10_N_btm.n1070 C10_N_btm.n811 0.109875
R42832 C10_N_btm.n1072 C10_N_btm.n811 0.109875
R42833 C10_N_btm.n1073 C10_N_btm.n810 0.109875
R42834 C10_N_btm.n1075 C10_N_btm.n810 0.109875
R42835 C10_N_btm.n1076 C10_N_btm.n807 0.109875
R42836 C10_N_btm.n1078 C10_N_btm.n807 0.109875
R42837 C10_N_btm.n1085 C10_N_btm.n808 0.109875
R42838 C10_N_btm.n1085 C10_N_btm.n1084 0.109875
R42839 C10_N_btm.n828 C10_N_btm.n825 0.109875
R42840 C10_N_btm.n826 C10_N_btm.n825 0.109875
R42841 C10_N_btm.n831 C10_N_btm.n824 0.109875
R42842 C10_N_btm.n829 C10_N_btm.n824 0.109875
R42843 C10_N_btm.n834 C10_N_btm.n823 0.109875
R42844 C10_N_btm.n832 C10_N_btm.n823 0.109875
R42845 C10_N_btm.n837 C10_N_btm.n822 0.109875
R42846 C10_N_btm.n835 C10_N_btm.n822 0.109875
R42847 C10_N_btm.n840 C10_N_btm.n821 0.109875
R42848 C10_N_btm.n838 C10_N_btm.n821 0.109875
R42849 C10_N_btm.n843 C10_N_btm.n820 0.109875
R42850 C10_N_btm.n841 C10_N_btm.n820 0.109875
R42851 C10_N_btm.n846 C10_N_btm.n819 0.109875
R42852 C10_N_btm.n844 C10_N_btm.n819 0.109875
R42853 C10_N_btm.n849 C10_N_btm.n818 0.109875
R42854 C10_N_btm.n849 C10_N_btm.n848 0.109875
R42855 C10_N_btm.n1114 C10_N_btm.n799 0.109875
R42856 C10_N_btm.n1112 C10_N_btm.n799 0.109875
R42857 C10_N_btm.n1111 C10_N_btm.n800 0.109875
R42858 C10_N_btm.n1109 C10_N_btm.n800 0.109875
R42859 C10_N_btm.n1108 C10_N_btm.n801 0.109875
R42860 C10_N_btm.n1106 C10_N_btm.n801 0.109875
R42861 C10_N_btm.n1105 C10_N_btm.n802 0.109875
R42862 C10_N_btm.n1103 C10_N_btm.n802 0.109875
R42863 C10_N_btm.n1102 C10_N_btm.n803 0.109875
R42864 C10_N_btm.n1100 C10_N_btm.n803 0.109875
R42865 C10_N_btm.n1099 C10_N_btm.n804 0.109875
R42866 C10_N_btm.n1097 C10_N_btm.n804 0.109875
R42867 C10_N_btm.n1096 C10_N_btm.n805 0.109875
R42868 C10_N_btm.n1094 C10_N_btm.n805 0.109875
R42869 C10_N_btm.n1093 C10_N_btm.n806 0.109875
R42870 C10_N_btm.n1091 C10_N_btm.n806 0.109875
R42871 C10_N_btm.n1090 C10_N_btm.n1086 0.109875
R42872 C10_N_btm.n1088 C10_N_btm.n1086 0.109875
R42873 C10_N_btm.n1143 C10_N_btm.n754 0.109875
R42874 C10_N_btm.n1145 C10_N_btm.n754 0.109875
R42875 C10_N_btm.n1140 C10_N_btm.n757 0.109875
R42876 C10_N_btm.n1142 C10_N_btm.n757 0.109875
R42877 C10_N_btm.n1137 C10_N_btm.n758 0.109875
R42878 C10_N_btm.n1139 C10_N_btm.n758 0.109875
R42879 C10_N_btm.n1134 C10_N_btm.n759 0.109875
R42880 C10_N_btm.n1136 C10_N_btm.n759 0.109875
R42881 C10_N_btm.n1131 C10_N_btm.n760 0.109875
R42882 C10_N_btm.n1133 C10_N_btm.n760 0.109875
R42883 C10_N_btm.n1128 C10_N_btm.n761 0.109875
R42884 C10_N_btm.n1130 C10_N_btm.n761 0.109875
R42885 C10_N_btm.n1125 C10_N_btm.n762 0.109875
R42886 C10_N_btm.n1127 C10_N_btm.n762 0.109875
R42887 C10_N_btm.n1122 C10_N_btm.n763 0.109875
R42888 C10_N_btm.n1124 C10_N_btm.n763 0.109875
R42889 C10_N_btm.n1119 C10_N_btm.n797 0.109875
R42890 C10_N_btm.n1121 C10_N_btm.n797 0.109875
R42891 C10_N_btm.n796 C10_N_btm.n765 0.109875
R42892 C10_N_btm.n796 C10_N_btm.n795 0.109875
R42893 C10_N_btm.n793 C10_N_btm.n766 0.109875
R42894 C10_N_btm.n791 C10_N_btm.n766 0.109875
R42895 C10_N_btm.n790 C10_N_btm.n767 0.109875
R42896 C10_N_btm.n788 C10_N_btm.n767 0.109875
R42897 C10_N_btm.n787 C10_N_btm.n768 0.109875
R42898 C10_N_btm.n785 C10_N_btm.n768 0.109875
R42899 C10_N_btm.n784 C10_N_btm.n769 0.109875
R42900 C10_N_btm.n782 C10_N_btm.n769 0.109875
R42901 C10_N_btm.n781 C10_N_btm.n770 0.109875
R42902 C10_N_btm.n779 C10_N_btm.n770 0.109875
R42903 C10_N_btm.n778 C10_N_btm.n771 0.109875
R42904 C10_N_btm.n776 C10_N_btm.n771 0.109875
R42905 C10_N_btm.n775 C10_N_btm.n772 0.109875
R42906 C10_N_btm.n773 C10_N_btm.n772 0.109875
R42907 C10_N_btm.n1152 C10_N_btm.n755 0.109875
R42908 C10_N_btm.n1152 C10_N_btm.n1151 0.109875
R42909 C10_N_btm.n1157 C10_N_btm.n1153 0.109875
R42910 C10_N_btm.n1155 C10_N_btm.n1153 0.109875
R42911 C10_N_btm.n1160 C10_N_btm.n753 0.109875
R42912 C10_N_btm.n1158 C10_N_btm.n753 0.109875
R42913 C10_N_btm.n1163 C10_N_btm.n752 0.109875
R42914 C10_N_btm.n1161 C10_N_btm.n752 0.109875
R42915 C10_N_btm.n1166 C10_N_btm.n751 0.109875
R42916 C10_N_btm.n1164 C10_N_btm.n751 0.109875
R42917 C10_N_btm.n1169 C10_N_btm.n750 0.109875
R42918 C10_N_btm.n1167 C10_N_btm.n750 0.109875
R42919 C10_N_btm.n1172 C10_N_btm.n749 0.109875
R42920 C10_N_btm.n1170 C10_N_btm.n749 0.109875
R42921 C10_N_btm.n1175 C10_N_btm.n748 0.109875
R42922 C10_N_btm.n1173 C10_N_btm.n748 0.109875
R42923 C10_N_btm.n1178 C10_N_btm.n747 0.109875
R42924 C10_N_btm.n1176 C10_N_btm.n747 0.109875
R42925 C10_N_btm.n1181 C10_N_btm.n746 0.109875
R42926 C10_N_btm.n1179 C10_N_btm.n746 0.109875
R42927 C10_N_btm.n1186 C10_N_btm.n744 0.109875
R42928 C10_N_btm.n1188 C10_N_btm.n744 0.109875
R42929 C10_N_btm.n1189 C10_N_btm.n710 0.109875
R42930 C10_N_btm.n1191 C10_N_btm.n710 0.109875
R42931 C10_N_btm.n1192 C10_N_btm.n709 0.109875
R42932 C10_N_btm.n1194 C10_N_btm.n709 0.109875
R42933 C10_N_btm.n1195 C10_N_btm.n708 0.109875
R42934 C10_N_btm.n1197 C10_N_btm.n708 0.109875
R42935 C10_N_btm.n1198 C10_N_btm.n707 0.109875
R42936 C10_N_btm.n1200 C10_N_btm.n707 0.109875
R42937 C10_N_btm.n1201 C10_N_btm.n706 0.109875
R42938 C10_N_btm.n1203 C10_N_btm.n706 0.109875
R42939 C10_N_btm.n1204 C10_N_btm.n705 0.109875
R42940 C10_N_btm.n1206 C10_N_btm.n705 0.109875
R42941 C10_N_btm.n1207 C10_N_btm.n704 0.109875
R42942 C10_N_btm.n1209 C10_N_btm.n704 0.109875
R42943 C10_N_btm.n1210 C10_N_btm.n701 0.109875
R42944 C10_N_btm.n1212 C10_N_btm.n701 0.109875
R42945 C10_N_btm.n1219 C10_N_btm.n702 0.109875
R42946 C10_N_btm.n1219 C10_N_btm.n1218 0.109875
R42947 C10_N_btm.n722 C10_N_btm.n719 0.109875
R42948 C10_N_btm.n720 C10_N_btm.n719 0.109875
R42949 C10_N_btm.n725 C10_N_btm.n718 0.109875
R42950 C10_N_btm.n723 C10_N_btm.n718 0.109875
R42951 C10_N_btm.n728 C10_N_btm.n717 0.109875
R42952 C10_N_btm.n726 C10_N_btm.n717 0.109875
R42953 C10_N_btm.n731 C10_N_btm.n716 0.109875
R42954 C10_N_btm.n729 C10_N_btm.n716 0.109875
R42955 C10_N_btm.n734 C10_N_btm.n715 0.109875
R42956 C10_N_btm.n732 C10_N_btm.n715 0.109875
R42957 C10_N_btm.n737 C10_N_btm.n714 0.109875
R42958 C10_N_btm.n735 C10_N_btm.n714 0.109875
R42959 C10_N_btm.n740 C10_N_btm.n713 0.109875
R42960 C10_N_btm.n738 C10_N_btm.n713 0.109875
R42961 C10_N_btm.n743 C10_N_btm.n712 0.109875
R42962 C10_N_btm.n743 C10_N_btm.n742 0.109875
R42963 C10_N_btm.n1248 C10_N_btm.n693 0.109875
R42964 C10_N_btm.n1246 C10_N_btm.n693 0.109875
R42965 C10_N_btm.n1245 C10_N_btm.n694 0.109875
R42966 C10_N_btm.n1243 C10_N_btm.n694 0.109875
R42967 C10_N_btm.n1242 C10_N_btm.n695 0.109875
R42968 C10_N_btm.n1240 C10_N_btm.n695 0.109875
R42969 C10_N_btm.n1239 C10_N_btm.n696 0.109875
R42970 C10_N_btm.n1237 C10_N_btm.n696 0.109875
R42971 C10_N_btm.n1236 C10_N_btm.n697 0.109875
R42972 C10_N_btm.n1234 C10_N_btm.n697 0.109875
R42973 C10_N_btm.n1233 C10_N_btm.n698 0.109875
R42974 C10_N_btm.n1231 C10_N_btm.n698 0.109875
R42975 C10_N_btm.n1230 C10_N_btm.n699 0.109875
R42976 C10_N_btm.n1228 C10_N_btm.n699 0.109875
R42977 C10_N_btm.n1227 C10_N_btm.n700 0.109875
R42978 C10_N_btm.n1225 C10_N_btm.n700 0.109875
R42979 C10_N_btm.n1224 C10_N_btm.n1220 0.109875
R42980 C10_N_btm.n1222 C10_N_btm.n1220 0.109875
R42981 C10_N_btm.n1277 C10_N_btm.n648 0.109875
R42982 C10_N_btm.n1279 C10_N_btm.n648 0.109875
R42983 C10_N_btm.n1274 C10_N_btm.n651 0.109875
R42984 C10_N_btm.n1276 C10_N_btm.n651 0.109875
R42985 C10_N_btm.n1271 C10_N_btm.n652 0.109875
R42986 C10_N_btm.n1273 C10_N_btm.n652 0.109875
R42987 C10_N_btm.n1268 C10_N_btm.n653 0.109875
R42988 C10_N_btm.n1270 C10_N_btm.n653 0.109875
R42989 C10_N_btm.n1265 C10_N_btm.n654 0.109875
R42990 C10_N_btm.n1267 C10_N_btm.n654 0.109875
R42991 C10_N_btm.n1262 C10_N_btm.n655 0.109875
R42992 C10_N_btm.n1264 C10_N_btm.n655 0.109875
R42993 C10_N_btm.n1259 C10_N_btm.n656 0.109875
R42994 C10_N_btm.n1261 C10_N_btm.n656 0.109875
R42995 C10_N_btm.n1256 C10_N_btm.n657 0.109875
R42996 C10_N_btm.n1258 C10_N_btm.n657 0.109875
R42997 C10_N_btm.n1253 C10_N_btm.n691 0.109875
R42998 C10_N_btm.n1255 C10_N_btm.n691 0.109875
R42999 C10_N_btm.n690 C10_N_btm.n659 0.109875
R43000 C10_N_btm.n690 C10_N_btm.n689 0.109875
R43001 C10_N_btm.n687 C10_N_btm.n660 0.109875
R43002 C10_N_btm.n685 C10_N_btm.n660 0.109875
R43003 C10_N_btm.n684 C10_N_btm.n661 0.109875
R43004 C10_N_btm.n682 C10_N_btm.n661 0.109875
R43005 C10_N_btm.n681 C10_N_btm.n662 0.109875
R43006 C10_N_btm.n679 C10_N_btm.n662 0.109875
R43007 C10_N_btm.n678 C10_N_btm.n663 0.109875
R43008 C10_N_btm.n676 C10_N_btm.n663 0.109875
R43009 C10_N_btm.n675 C10_N_btm.n664 0.109875
R43010 C10_N_btm.n673 C10_N_btm.n664 0.109875
R43011 C10_N_btm.n672 C10_N_btm.n665 0.109875
R43012 C10_N_btm.n670 C10_N_btm.n665 0.109875
R43013 C10_N_btm.n669 C10_N_btm.n666 0.109875
R43014 C10_N_btm.n667 C10_N_btm.n666 0.109875
R43015 C10_N_btm.n1286 C10_N_btm.n649 0.109875
R43016 C10_N_btm.n1286 C10_N_btm.n1285 0.109875
R43017 C10_N_btm.n1291 C10_N_btm.n1287 0.109875
R43018 C10_N_btm.n1289 C10_N_btm.n1287 0.109875
R43019 C10_N_btm.n1294 C10_N_btm.n647 0.109875
R43020 C10_N_btm.n1292 C10_N_btm.n647 0.109875
R43021 C10_N_btm.n1297 C10_N_btm.n646 0.109875
R43022 C10_N_btm.n1295 C10_N_btm.n646 0.109875
R43023 C10_N_btm.n1300 C10_N_btm.n645 0.109875
R43024 C10_N_btm.n1298 C10_N_btm.n645 0.109875
R43025 C10_N_btm.n1303 C10_N_btm.n644 0.109875
R43026 C10_N_btm.n1301 C10_N_btm.n644 0.109875
R43027 C10_N_btm.n1306 C10_N_btm.n643 0.109875
R43028 C10_N_btm.n1304 C10_N_btm.n643 0.109875
R43029 C10_N_btm.n1309 C10_N_btm.n642 0.109875
R43030 C10_N_btm.n1307 C10_N_btm.n642 0.109875
R43031 C10_N_btm.n1312 C10_N_btm.n641 0.109875
R43032 C10_N_btm.n1310 C10_N_btm.n641 0.109875
R43033 C10_N_btm.n1315 C10_N_btm.n640 0.109875
R43034 C10_N_btm.n1313 C10_N_btm.n640 0.109875
R43035 C10_N_btm.n1320 C10_N_btm.n638 0.109875
R43036 C10_N_btm.n1322 C10_N_btm.n638 0.109875
R43037 C10_N_btm.n1323 C10_N_btm.n604 0.109875
R43038 C10_N_btm.n1325 C10_N_btm.n604 0.109875
R43039 C10_N_btm.n1326 C10_N_btm.n603 0.109875
R43040 C10_N_btm.n1328 C10_N_btm.n603 0.109875
R43041 C10_N_btm.n1329 C10_N_btm.n602 0.109875
R43042 C10_N_btm.n1331 C10_N_btm.n602 0.109875
R43043 C10_N_btm.n1332 C10_N_btm.n601 0.109875
R43044 C10_N_btm.n1334 C10_N_btm.n601 0.109875
R43045 C10_N_btm.n1335 C10_N_btm.n600 0.109875
R43046 C10_N_btm.n1337 C10_N_btm.n600 0.109875
R43047 C10_N_btm.n1338 C10_N_btm.n599 0.109875
R43048 C10_N_btm.n1340 C10_N_btm.n599 0.109875
R43049 C10_N_btm.n1341 C10_N_btm.n598 0.109875
R43050 C10_N_btm.n1343 C10_N_btm.n598 0.109875
R43051 C10_N_btm.n1344 C10_N_btm.n595 0.109875
R43052 C10_N_btm.n1346 C10_N_btm.n595 0.109875
R43053 C10_N_btm.n1353 C10_N_btm.n596 0.109875
R43054 C10_N_btm.n1353 C10_N_btm.n1352 0.109875
R43055 C10_N_btm.n616 C10_N_btm.n613 0.109875
R43056 C10_N_btm.n614 C10_N_btm.n613 0.109875
R43057 C10_N_btm.n619 C10_N_btm.n612 0.109875
R43058 C10_N_btm.n617 C10_N_btm.n612 0.109875
R43059 C10_N_btm.n622 C10_N_btm.n611 0.109875
R43060 C10_N_btm.n620 C10_N_btm.n611 0.109875
R43061 C10_N_btm.n625 C10_N_btm.n610 0.109875
R43062 C10_N_btm.n623 C10_N_btm.n610 0.109875
R43063 C10_N_btm.n628 C10_N_btm.n609 0.109875
R43064 C10_N_btm.n626 C10_N_btm.n609 0.109875
R43065 C10_N_btm.n631 C10_N_btm.n608 0.109875
R43066 C10_N_btm.n629 C10_N_btm.n608 0.109875
R43067 C10_N_btm.n634 C10_N_btm.n607 0.109875
R43068 C10_N_btm.n632 C10_N_btm.n607 0.109875
R43069 C10_N_btm.n637 C10_N_btm.n606 0.109875
R43070 C10_N_btm.n637 C10_N_btm.n636 0.109875
R43071 C10_N_btm.n1382 C10_N_btm.n587 0.109875
R43072 C10_N_btm.n1380 C10_N_btm.n587 0.109875
R43073 C10_N_btm.n1379 C10_N_btm.n588 0.109875
R43074 C10_N_btm.n1377 C10_N_btm.n588 0.109875
R43075 C10_N_btm.n1376 C10_N_btm.n589 0.109875
R43076 C10_N_btm.n1374 C10_N_btm.n589 0.109875
R43077 C10_N_btm.n1373 C10_N_btm.n590 0.109875
R43078 C10_N_btm.n1371 C10_N_btm.n590 0.109875
R43079 C10_N_btm.n1370 C10_N_btm.n591 0.109875
R43080 C10_N_btm.n1368 C10_N_btm.n591 0.109875
R43081 C10_N_btm.n1367 C10_N_btm.n592 0.109875
R43082 C10_N_btm.n1365 C10_N_btm.n592 0.109875
R43083 C10_N_btm.n1364 C10_N_btm.n593 0.109875
R43084 C10_N_btm.n1362 C10_N_btm.n593 0.109875
R43085 C10_N_btm.n1361 C10_N_btm.n594 0.109875
R43086 C10_N_btm.n1359 C10_N_btm.n594 0.109875
R43087 C10_N_btm.n1358 C10_N_btm.n1354 0.109875
R43088 C10_N_btm.n1356 C10_N_btm.n1354 0.109875
R43089 C10_N_btm.n1446 C10_N_btm.n575 0.109875
R43090 C10_N_btm.n1448 C10_N_btm.n575 0.109875
R43091 C10_N_btm.n1443 C10_N_btm.n578 0.109875
R43092 C10_N_btm.n1445 C10_N_btm.n578 0.109875
R43093 C10_N_btm.n1440 C10_N_btm.n579 0.109875
R43094 C10_N_btm.n1442 C10_N_btm.n579 0.109875
R43095 C10_N_btm.n1437 C10_N_btm.n580 0.109875
R43096 C10_N_btm.n1439 C10_N_btm.n580 0.109875
R43097 C10_N_btm.n1434 C10_N_btm.n581 0.109875
R43098 C10_N_btm.n1436 C10_N_btm.n581 0.109875
R43099 C10_N_btm.n1431 C10_N_btm.n582 0.109875
R43100 C10_N_btm.n1433 C10_N_btm.n582 0.109875
R43101 C10_N_btm.n1428 C10_N_btm.n583 0.109875
R43102 C10_N_btm.n1430 C10_N_btm.n583 0.109875
R43103 C10_N_btm.n1425 C10_N_btm.n584 0.109875
R43104 C10_N_btm.n1427 C10_N_btm.n584 0.109875
R43105 C10_N_btm.n1422 C10_N_btm.n585 0.109875
R43106 C10_N_btm.n1424 C10_N_btm.n585 0.109875
R43107 C10_N_btm.n1417 C10_N_btm.n566 0.109875
R43108 C10_N_btm.n1415 C10_N_btm.n566 0.109875
R43109 C10_N_btm.n1414 C10_N_btm.n1387 0.109875
R43110 C10_N_btm.n1412 C10_N_btm.n1387 0.109875
R43111 C10_N_btm.n1411 C10_N_btm.n1388 0.109875
R43112 C10_N_btm.n1409 C10_N_btm.n1388 0.109875
R43113 C10_N_btm.n1408 C10_N_btm.n1389 0.109875
R43114 C10_N_btm.n1406 C10_N_btm.n1389 0.109875
R43115 C10_N_btm.n1405 C10_N_btm.n1390 0.109875
R43116 C10_N_btm.n1403 C10_N_btm.n1390 0.109875
R43117 C10_N_btm.n1402 C10_N_btm.n1391 0.109875
R43118 C10_N_btm.n1400 C10_N_btm.n1391 0.109875
R43119 C10_N_btm.n1399 C10_N_btm.n1392 0.109875
R43120 C10_N_btm.n1397 C10_N_btm.n1392 0.109875
R43121 C10_N_btm.n1396 C10_N_btm.n1393 0.109875
R43122 C10_N_btm.n1394 C10_N_btm.n1393 0.109875
R43123 C10_N_btm.n1455 C10_N_btm.n576 0.109875
R43124 C10_N_btm.n1455 C10_N_btm.n1454 0.109875
R43125 C10_N_btm.n1460 C10_N_btm.n1456 0.109875
R43126 C10_N_btm.n1458 C10_N_btm.n1456 0.109875
R43127 C10_N_btm.n1463 C10_N_btm.n574 0.109875
R43128 C10_N_btm.n1461 C10_N_btm.n574 0.109875
R43129 C10_N_btm.n1466 C10_N_btm.n573 0.109875
R43130 C10_N_btm.n1464 C10_N_btm.n573 0.109875
R43131 C10_N_btm.n1469 C10_N_btm.n572 0.109875
R43132 C10_N_btm.n1467 C10_N_btm.n572 0.109875
R43133 C10_N_btm.n1472 C10_N_btm.n571 0.109875
R43134 C10_N_btm.n1470 C10_N_btm.n571 0.109875
R43135 C10_N_btm.n1475 C10_N_btm.n570 0.109875
R43136 C10_N_btm.n1473 C10_N_btm.n570 0.109875
R43137 C10_N_btm.n1478 C10_N_btm.n569 0.109875
R43138 C10_N_btm.n1476 C10_N_btm.n569 0.109875
R43139 C10_N_btm.n1481 C10_N_btm.n568 0.109875
R43140 C10_N_btm.n1479 C10_N_btm.n568 0.109875
R43141 C10_N_btm.n1484 C10_N_btm.n567 0.109875
R43142 C10_N_btm.n1484 C10_N_btm.n1483 0.109875
R43143 C10_N_btm.n1487 C10_N_btm.n1485 0.109875
R43144 C10_N_btm.n1489 C10_N_btm.n1485 0.109875
R43145 C10_N_btm.n1490 C10_N_btm.n565 0.109875
R43146 C10_N_btm.n1492 C10_N_btm.n565 0.109875
R43147 C10_N_btm.n1493 C10_N_btm.n564 0.109875
R43148 C10_N_btm.n1495 C10_N_btm.n564 0.109875
R43149 C10_N_btm.n1496 C10_N_btm.n563 0.109875
R43150 C10_N_btm.n1498 C10_N_btm.n563 0.109875
R43151 C10_N_btm.n1499 C10_N_btm.n562 0.109875
R43152 C10_N_btm.n1501 C10_N_btm.n562 0.109875
R43153 C10_N_btm.n1502 C10_N_btm.n561 0.109875
R43154 C10_N_btm.n1504 C10_N_btm.n561 0.109875
R43155 C10_N_btm.n1505 C10_N_btm.n560 0.109875
R43156 C10_N_btm.n1507 C10_N_btm.n560 0.109875
R43157 C10_N_btm.n1508 C10_N_btm.n559 0.109875
R43158 C10_N_btm.n1510 C10_N_btm.n559 0.109875
R43159 C10_N_btm.n1511 C10_N_btm.n558 0.109875
R43160 C10_N_btm.n1513 C10_N_btm.n558 0.109875
R43161 C10_N_btm.n1532 C10_N_btm.n1528 0.109875
R43162 C10_N_btm.n1530 C10_N_btm.n1528 0.109875
R43163 C10_N_btm.n1535 C10_N_btm.n1527 0.109875
R43164 C10_N_btm.n1533 C10_N_btm.n1527 0.109875
R43165 C10_N_btm.n1538 C10_N_btm.n1526 0.109875
R43166 C10_N_btm.n1536 C10_N_btm.n1526 0.109875
R43167 C10_N_btm.n1541 C10_N_btm.n1525 0.109875
R43168 C10_N_btm.n1539 C10_N_btm.n1525 0.109875
R43169 C10_N_btm.n1544 C10_N_btm.n1524 0.109875
R43170 C10_N_btm.n1542 C10_N_btm.n1524 0.109875
R43171 C10_N_btm.n1547 C10_N_btm.n1523 0.109875
R43172 C10_N_btm.n1545 C10_N_btm.n1523 0.109875
R43173 C10_N_btm.n1550 C10_N_btm.n1522 0.109875
R43174 C10_N_btm.n1548 C10_N_btm.n1522 0.109875
R43175 C10_N_btm.n1553 C10_N_btm.n1521 0.109875
R43176 C10_N_btm.n1551 C10_N_btm.n1521 0.109875
R43177 C10_N_btm.n1556 C10_N_btm.n1520 0.109875
R43178 C10_N_btm.n1554 C10_N_btm.n1520 0.109875
R43179 C10_N_btm.n1559 C10_N_btm.n1519 0.109875
R43180 C10_N_btm.n1557 C10_N_btm.n1519 0.109875
R43181 C10_N_btm.n1562 C10_N_btm.n1518 0.109875
R43182 C10_N_btm.n1560 C10_N_btm.n1518 0.109875
R43183 C10_N_btm.n1565 C10_N_btm.n1517 0.109875
R43184 C10_N_btm.n1563 C10_N_btm.n1517 0.109875
R43185 C10_N_btm.n1568 C10_N_btm.n1516 0.109875
R43186 C10_N_btm.n1566 C10_N_btm.n1516 0.109875
R43187 C10_N_btm.n1571 C10_N_btm.n556 0.109875
R43188 C10_N_btm.n1569 C10_N_btm.n556 0.109875
R43189 C10_N_btm.n1574 C10_N_btm.n555 0.109875
R43190 C10_N_btm.n1572 C10_N_btm.n555 0.109875
R43191 C10_N_btm.n1577 C10_N_btm.n554 0.109875
R43192 C10_N_btm.n1575 C10_N_btm.n554 0.109875
R43193 C10_N_btm.n1580 C10_N_btm.n553 0.109875
R43194 C10_N_btm.n1578 C10_N_btm.n553 0.109875
R43195 C10_N_btm.n1583 C10_N_btm.n552 0.109875
R43196 C10_N_btm.n1581 C10_N_btm.n552 0.109875
R43197 C10_N_btm.n1586 C10_N_btm.n551 0.109875
R43198 C10_N_btm.n1584 C10_N_btm.n551 0.109875
R43199 C10_N_btm.n1589 C10_N_btm.n550 0.109875
R43200 C10_N_btm.n1587 C10_N_btm.n550 0.109875
R43201 C10_N_btm.n1592 C10_N_btm.n549 0.109875
R43202 C10_N_btm.n1590 C10_N_btm.n549 0.109875
R43203 C10_N_btm.n1595 C10_N_btm.n548 0.109875
R43204 C10_N_btm.n1593 C10_N_btm.n548 0.109875
R43205 C10_N_btm.n3109 C10_N_btm.n546 0.109875
R43206 C10_N_btm.n3111 C10_N_btm.n546 0.109875
R43207 C10_N_btm.n3112 C10_N_btm.n545 0.109875
R43208 C10_N_btm.n3114 C10_N_btm.n545 0.109875
R43209 C10_N_btm.n3115 C10_N_btm.n544 0.109875
R43210 C10_N_btm.n3117 C10_N_btm.n544 0.109875
R43211 C10_N_btm.n3118 C10_N_btm.n543 0.109875
R43212 C10_N_btm.n3120 C10_N_btm.n543 0.109875
R43213 C10_N_btm.n3121 C10_N_btm.n542 0.109875
R43214 C10_N_btm.n3123 C10_N_btm.n542 0.109875
R43215 C10_N_btm.n3124 C10_N_btm.n541 0.109875
R43216 C10_N_btm.n3126 C10_N_btm.n541 0.109875
R43217 C10_N_btm.n3127 C10_N_btm.n540 0.109875
R43218 C10_N_btm.n3129 C10_N_btm.n540 0.109875
R43219 C10_N_btm.n3130 C10_N_btm.n539 0.109875
R43220 C10_N_btm.n3132 C10_N_btm.n539 0.109875
R43221 C10_N_btm.n3133 C10_N_btm.n538 0.109875
R43222 C10_N_btm.n3135 C10_N_btm.n538 0.109875
R43223 C10_N_btm.n3136 C10_N_btm.n537 0.109875
R43224 C10_N_btm.n3138 C10_N_btm.n537 0.109875
R43225 C10_N_btm.n3139 C10_N_btm.n536 0.109875
R43226 C10_N_btm.n3141 C10_N_btm.n536 0.109875
R43227 C10_N_btm.n3142 C10_N_btm.n535 0.109875
R43228 C10_N_btm.n3144 C10_N_btm.n535 0.109875
R43229 C10_N_btm.n3145 C10_N_btm.n534 0.109875
R43230 C10_N_btm.n3147 C10_N_btm.n534 0.109875
R43231 C10_N_btm.n3148 C10_N_btm.n533 0.109875
R43232 C10_N_btm.n3150 C10_N_btm.n533 0.109875
R43233 C10_N_btm.n3151 C10_N_btm.n532 0.109875
R43234 C10_N_btm.n3153 C10_N_btm.n532 0.109875
R43235 C10_N_btm.n3154 C10_N_btm.n531 0.109875
R43236 C10_N_btm.n3156 C10_N_btm.n531 0.109875
R43237 C10_N_btm.n3157 C10_N_btm.n530 0.109875
R43238 C10_N_btm.n3159 C10_N_btm.n530 0.109875
R43239 C10_N_btm.n3160 C10_N_btm.n529 0.109875
R43240 C10_N_btm.n3162 C10_N_btm.n529 0.109875
R43241 C10_N_btm.n3163 C10_N_btm.n528 0.109875
R43242 C10_N_btm.n3165 C10_N_btm.n528 0.109875
R43243 C10_N_btm.n3166 C10_N_btm.n527 0.109875
R43244 C10_N_btm.n3168 C10_N_btm.n527 0.109875
R43245 C10_N_btm.n3169 C10_N_btm.n526 0.109875
R43246 C10_N_btm.n3171 C10_N_btm.n526 0.109875
R43247 C10_N_btm.n3172 C10_N_btm.n525 0.109875
R43248 C10_N_btm.n3174 C10_N_btm.n525 0.109875
R43249 C10_N_btm.n3175 C10_N_btm.n524 0.109875
R43250 C10_N_btm.n3177 C10_N_btm.n524 0.109875
R43251 C10_N_btm.n3178 C10_N_btm.n523 0.109875
R43252 C10_N_btm.n3180 C10_N_btm.n523 0.109875
R43253 C10_N_btm.n3181 C10_N_btm.n522 0.109875
R43254 C10_N_btm.n3183 C10_N_btm.n522 0.109875
R43255 C10_N_btm.n3184 C10_N_btm.n521 0.109875
R43256 C10_N_btm.n3186 C10_N_btm.n521 0.109875
R43257 C10_N_btm.n3187 C10_N_btm.n520 0.109875
R43258 C10_N_btm.n3189 C10_N_btm.n520 0.109875
R43259 C10_N_btm.n3190 C10_N_btm.n519 0.109875
R43260 C10_N_btm.n3192 C10_N_btm.n519 0.109875
R43261 C10_N_btm.n3193 C10_N_btm.n518 0.109875
R43262 C10_N_btm.n3195 C10_N_btm.n518 0.109875
R43263 C10_N_btm.n3196 C10_N_btm.n517 0.109875
R43264 C10_N_btm.n3198 C10_N_btm.n517 0.109875
R43265 C10_N_btm.n3199 C10_N_btm.n516 0.109875
R43266 C10_N_btm.n3201 C10_N_btm.n516 0.109875
R43267 C10_N_btm.n3202 C10_N_btm.n515 0.109875
R43268 C10_N_btm.n3204 C10_N_btm.n515 0.109875
R43269 C10_N_btm.n3205 C10_N_btm.n514 0.109875
R43270 C10_N_btm.n3207 C10_N_btm.n514 0.109875
R43271 C10_N_btm.n3208 C10_N_btm.n513 0.109875
R43272 C10_N_btm.n3210 C10_N_btm.n513 0.109875
R43273 C10_N_btm.n3211 C10_N_btm.n512 0.109875
R43274 C10_N_btm.n3213 C10_N_btm.n512 0.109875
R43275 C10_N_btm.n3214 C10_N_btm.n511 0.109875
R43276 C10_N_btm.n3216 C10_N_btm.n511 0.109875
R43277 C10_N_btm.n3217 C10_N_btm.n510 0.109875
R43278 C10_N_btm.n3219 C10_N_btm.n510 0.109875
R43279 C10_N_btm.n3220 C10_N_btm.n509 0.109875
R43280 C10_N_btm.n3222 C10_N_btm.n509 0.109875
R43281 C10_N_btm.n3223 C10_N_btm.n508 0.109875
R43282 C10_N_btm.n3225 C10_N_btm.n508 0.109875
R43283 C10_N_btm.n3226 C10_N_btm.n507 0.109875
R43284 C10_N_btm.n3228 C10_N_btm.n507 0.109875
R43285 C10_N_btm.n3229 C10_N_btm.n422 0.109875
R43286 C10_N_btm.n3231 C10_N_btm.n422 0.109875
R43287 C10_N_btm.n3232 C10_N_btm.n421 0.109875
R43288 C10_N_btm.n3234 C10_N_btm.n421 0.109875
R43289 C10_N_btm.n3235 C10_N_btm.n420 0.109875
R43290 C10_N_btm.n3237 C10_N_btm.n420 0.109875
R43291 C10_N_btm.n3238 C10_N_btm.n419 0.109875
R43292 C10_N_btm.n3240 C10_N_btm.n419 0.109875
R43293 C10_N_btm.n3241 C10_N_btm.n418 0.109875
R43294 C10_N_btm.n3243 C10_N_btm.n418 0.109875
R43295 C10_N_btm.n3244 C10_N_btm.n417 0.109875
R43296 C10_N_btm.n3246 C10_N_btm.n417 0.109875
R43297 C10_N_btm.n3247 C10_N_btm.n416 0.109875
R43298 C10_N_btm.n3249 C10_N_btm.n416 0.109875
R43299 C10_N_btm.n3250 C10_N_btm.n415 0.109875
R43300 C10_N_btm.n3252 C10_N_btm.n415 0.109875
R43301 C10_N_btm.n3253 C10_N_btm.n414 0.109875
R43302 C10_N_btm.n3255 C10_N_btm.n414 0.109875
R43303 C10_N_btm.n3256 C10_N_btm.n413 0.109875
R43304 C10_N_btm.n3258 C10_N_btm.n413 0.109875
R43305 C10_N_btm.n3259 C10_N_btm.n412 0.109875
R43306 C10_N_btm.n3261 C10_N_btm.n412 0.109875
R43307 C10_N_btm.n3262 C10_N_btm.n411 0.109875
R43308 C10_N_btm.n3264 C10_N_btm.n411 0.109875
R43309 C10_N_btm.n3265 C10_N_btm.n410 0.109875
R43310 C10_N_btm.n3267 C10_N_btm.n410 0.109875
R43311 C10_N_btm.n3268 C10_N_btm.n409 0.109875
R43312 C10_N_btm.n3270 C10_N_btm.n409 0.109875
R43313 C10_N_btm.n3271 C10_N_btm.n408 0.109875
R43314 C10_N_btm.n3273 C10_N_btm.n408 0.109875
R43315 C10_N_btm.n3274 C10_N_btm.n407 0.109875
R43316 C10_N_btm.n3276 C10_N_btm.n407 0.109875
R43317 C10_N_btm.n3277 C10_N_btm.n406 0.109875
R43318 C10_N_btm.n3279 C10_N_btm.n406 0.109875
R43319 C10_N_btm.n3280 C10_N_btm.n405 0.109875
R43320 C10_N_btm.n3282 C10_N_btm.n405 0.109875
R43321 C10_N_btm.n3283 C10_N_btm.n404 0.109875
R43322 C10_N_btm.n3285 C10_N_btm.n404 0.109875
R43323 C10_N_btm.n3286 C10_N_btm.n403 0.109875
R43324 C10_N_btm.n3288 C10_N_btm.n403 0.109875
R43325 C10_N_btm.n3289 C10_N_btm.n402 0.109875
R43326 C10_N_btm.n3291 C10_N_btm.n402 0.109875
R43327 C10_N_btm.n3292 C10_N_btm.n399 0.109875
R43328 C10_N_btm.n3294 C10_N_btm.n399 0.109875
R43329 C10_N_btm.n3301 C10_N_btm.n400 0.109875
R43330 C10_N_btm.n3301 C10_N_btm.n3300 0.109875
R43331 C10_N_btm.n445 C10_N_btm.n442 0.109875
R43332 C10_N_btm.n443 C10_N_btm.n442 0.109875
R43333 C10_N_btm.n448 C10_N_btm.n441 0.109875
R43334 C10_N_btm.n446 C10_N_btm.n441 0.109875
R43335 C10_N_btm.n451 C10_N_btm.n440 0.109875
R43336 C10_N_btm.n449 C10_N_btm.n440 0.109875
R43337 C10_N_btm.n454 C10_N_btm.n439 0.109875
R43338 C10_N_btm.n452 C10_N_btm.n439 0.109875
R43339 C10_N_btm.n457 C10_N_btm.n438 0.109875
R43340 C10_N_btm.n455 C10_N_btm.n438 0.109875
R43341 C10_N_btm.n460 C10_N_btm.n437 0.109875
R43342 C10_N_btm.n458 C10_N_btm.n437 0.109875
R43343 C10_N_btm.n463 C10_N_btm.n436 0.109875
R43344 C10_N_btm.n461 C10_N_btm.n436 0.109875
R43345 C10_N_btm.n466 C10_N_btm.n435 0.109875
R43346 C10_N_btm.n464 C10_N_btm.n435 0.109875
R43347 C10_N_btm.n469 C10_N_btm.n390 0.109875
R43348 C10_N_btm.n467 C10_N_btm.n390 0.109875
R43349 C10_N_btm.n3330 C10_N_btm.n391 0.109875
R43350 C10_N_btm.n3328 C10_N_btm.n391 0.109875
R43351 C10_N_btm.n3327 C10_N_btm.n392 0.109875
R43352 C10_N_btm.n3325 C10_N_btm.n392 0.109875
R43353 C10_N_btm.n3324 C10_N_btm.n393 0.109875
R43354 C10_N_btm.n3322 C10_N_btm.n393 0.109875
R43355 C10_N_btm.n3321 C10_N_btm.n394 0.109875
R43356 C10_N_btm.n3319 C10_N_btm.n394 0.109875
R43357 C10_N_btm.n3318 C10_N_btm.n395 0.109875
R43358 C10_N_btm.n3316 C10_N_btm.n395 0.109875
R43359 C10_N_btm.n3315 C10_N_btm.n396 0.109875
R43360 C10_N_btm.n3313 C10_N_btm.n396 0.109875
R43361 C10_N_btm.n3312 C10_N_btm.n397 0.109875
R43362 C10_N_btm.n3310 C10_N_btm.n397 0.109875
R43363 C10_N_btm.n3309 C10_N_btm.n398 0.109875
R43364 C10_N_btm.n3307 C10_N_btm.n398 0.109875
R43365 C10_N_btm.n3306 C10_N_btm.n3302 0.109875
R43366 C10_N_btm.n3304 C10_N_btm.n3302 0.109875
R43367 C10_N_btm.n3359 C10_N_btm.n346 0.109875
R43368 C10_N_btm.n3361 C10_N_btm.n346 0.109875
R43369 C10_N_btm.n3356 C10_N_btm.n349 0.109875
R43370 C10_N_btm.n3358 C10_N_btm.n349 0.109875
R43371 C10_N_btm.n3353 C10_N_btm.n350 0.109875
R43372 C10_N_btm.n3355 C10_N_btm.n350 0.109875
R43373 C10_N_btm.n3350 C10_N_btm.n351 0.109875
R43374 C10_N_btm.n3352 C10_N_btm.n351 0.109875
R43375 C10_N_btm.n3347 C10_N_btm.n352 0.109875
R43376 C10_N_btm.n3349 C10_N_btm.n352 0.109875
R43377 C10_N_btm.n3344 C10_N_btm.n353 0.109875
R43378 C10_N_btm.n3346 C10_N_btm.n353 0.109875
R43379 C10_N_btm.n3341 C10_N_btm.n354 0.109875
R43380 C10_N_btm.n3343 C10_N_btm.n354 0.109875
R43381 C10_N_btm.n3338 C10_N_btm.n355 0.109875
R43382 C10_N_btm.n3340 C10_N_btm.n355 0.109875
R43383 C10_N_btm.n3335 C10_N_btm.n389 0.109875
R43384 C10_N_btm.n3337 C10_N_btm.n389 0.109875
R43385 C10_N_btm.n388 C10_N_btm.n357 0.109875
R43386 C10_N_btm.n388 C10_N_btm.n387 0.109875
R43387 C10_N_btm.n385 C10_N_btm.n358 0.109875
R43388 C10_N_btm.n383 C10_N_btm.n358 0.109875
R43389 C10_N_btm.n382 C10_N_btm.n359 0.109875
R43390 C10_N_btm.n380 C10_N_btm.n359 0.109875
R43391 C10_N_btm.n379 C10_N_btm.n360 0.109875
R43392 C10_N_btm.n377 C10_N_btm.n360 0.109875
R43393 C10_N_btm.n376 C10_N_btm.n361 0.109875
R43394 C10_N_btm.n374 C10_N_btm.n361 0.109875
R43395 C10_N_btm.n373 C10_N_btm.n362 0.109875
R43396 C10_N_btm.n371 C10_N_btm.n362 0.109875
R43397 C10_N_btm.n370 C10_N_btm.n363 0.109875
R43398 C10_N_btm.n368 C10_N_btm.n363 0.109875
R43399 C10_N_btm.n367 C10_N_btm.n364 0.109875
R43400 C10_N_btm.n365 C10_N_btm.n364 0.109875
R43401 C10_N_btm.n3368 C10_N_btm.n347 0.109875
R43402 C10_N_btm.n3368 C10_N_btm.n3367 0.109875
R43403 C10_N_btm.n3373 C10_N_btm.n3369 0.109875
R43404 C10_N_btm.n3371 C10_N_btm.n3369 0.109875
R43405 C10_N_btm.n3376 C10_N_btm.n345 0.109875
R43406 C10_N_btm.n3374 C10_N_btm.n345 0.109875
R43407 C10_N_btm.n3379 C10_N_btm.n344 0.109875
R43408 C10_N_btm.n3377 C10_N_btm.n344 0.109875
R43409 C10_N_btm.n3382 C10_N_btm.n343 0.109875
R43410 C10_N_btm.n3380 C10_N_btm.n343 0.109875
R43411 C10_N_btm.n3385 C10_N_btm.n342 0.109875
R43412 C10_N_btm.n3383 C10_N_btm.n342 0.109875
R43413 C10_N_btm.n3388 C10_N_btm.n341 0.109875
R43414 C10_N_btm.n3386 C10_N_btm.n341 0.109875
R43415 C10_N_btm.n3391 C10_N_btm.n340 0.109875
R43416 C10_N_btm.n3389 C10_N_btm.n340 0.109875
R43417 C10_N_btm.n3394 C10_N_btm.n339 0.109875
R43418 C10_N_btm.n3392 C10_N_btm.n339 0.109875
R43419 C10_N_btm.n3397 C10_N_btm.n338 0.109875
R43420 C10_N_btm.n3395 C10_N_btm.n338 0.109875
R43421 C10_N_btm.n3402 C10_N_btm.n336 0.109875
R43422 C10_N_btm.n3404 C10_N_btm.n336 0.109875
R43423 C10_N_btm.n3405 C10_N_btm.n302 0.109875
R43424 C10_N_btm.n3407 C10_N_btm.n302 0.109875
R43425 C10_N_btm.n3408 C10_N_btm.n301 0.109875
R43426 C10_N_btm.n3410 C10_N_btm.n301 0.109875
R43427 C10_N_btm.n3411 C10_N_btm.n300 0.109875
R43428 C10_N_btm.n3413 C10_N_btm.n300 0.109875
R43429 C10_N_btm.n3414 C10_N_btm.n299 0.109875
R43430 C10_N_btm.n3416 C10_N_btm.n299 0.109875
R43431 C10_N_btm.n3417 C10_N_btm.n298 0.109875
R43432 C10_N_btm.n3419 C10_N_btm.n298 0.109875
R43433 C10_N_btm.n3420 C10_N_btm.n297 0.109875
R43434 C10_N_btm.n3422 C10_N_btm.n297 0.109875
R43435 C10_N_btm.n3423 C10_N_btm.n296 0.109875
R43436 C10_N_btm.n3425 C10_N_btm.n296 0.109875
R43437 C10_N_btm.n3426 C10_N_btm.n293 0.109875
R43438 C10_N_btm.n3428 C10_N_btm.n293 0.109875
R43439 C10_N_btm.n3435 C10_N_btm.n294 0.109875
R43440 C10_N_btm.n3435 C10_N_btm.n3434 0.109875
R43441 C10_N_btm.n314 C10_N_btm.n311 0.109875
R43442 C10_N_btm.n312 C10_N_btm.n311 0.109875
R43443 C10_N_btm.n317 C10_N_btm.n310 0.109875
R43444 C10_N_btm.n315 C10_N_btm.n310 0.109875
R43445 C10_N_btm.n320 C10_N_btm.n309 0.109875
R43446 C10_N_btm.n318 C10_N_btm.n309 0.109875
R43447 C10_N_btm.n323 C10_N_btm.n308 0.109875
R43448 C10_N_btm.n321 C10_N_btm.n308 0.109875
R43449 C10_N_btm.n326 C10_N_btm.n307 0.109875
R43450 C10_N_btm.n324 C10_N_btm.n307 0.109875
R43451 C10_N_btm.n329 C10_N_btm.n306 0.109875
R43452 C10_N_btm.n327 C10_N_btm.n306 0.109875
R43453 C10_N_btm.n332 C10_N_btm.n305 0.109875
R43454 C10_N_btm.n330 C10_N_btm.n305 0.109875
R43455 C10_N_btm.n335 C10_N_btm.n304 0.109875
R43456 C10_N_btm.n335 C10_N_btm.n334 0.109875
R43457 C10_N_btm.n3464 C10_N_btm.n285 0.109875
R43458 C10_N_btm.n3462 C10_N_btm.n285 0.109875
R43459 C10_N_btm.n3461 C10_N_btm.n286 0.109875
R43460 C10_N_btm.n3459 C10_N_btm.n286 0.109875
R43461 C10_N_btm.n3458 C10_N_btm.n287 0.109875
R43462 C10_N_btm.n3456 C10_N_btm.n287 0.109875
R43463 C10_N_btm.n3455 C10_N_btm.n288 0.109875
R43464 C10_N_btm.n3453 C10_N_btm.n288 0.109875
R43465 C10_N_btm.n3452 C10_N_btm.n289 0.109875
R43466 C10_N_btm.n3450 C10_N_btm.n289 0.109875
R43467 C10_N_btm.n3449 C10_N_btm.n290 0.109875
R43468 C10_N_btm.n3447 C10_N_btm.n290 0.109875
R43469 C10_N_btm.n3446 C10_N_btm.n291 0.109875
R43470 C10_N_btm.n3444 C10_N_btm.n291 0.109875
R43471 C10_N_btm.n3443 C10_N_btm.n292 0.109875
R43472 C10_N_btm.n3441 C10_N_btm.n292 0.109875
R43473 C10_N_btm.n3440 C10_N_btm.n3436 0.109875
R43474 C10_N_btm.n3438 C10_N_btm.n3436 0.109875
R43475 C10_N_btm.n3493 C10_N_btm.n240 0.109875
R43476 C10_N_btm.n3495 C10_N_btm.n240 0.109875
R43477 C10_N_btm.n3490 C10_N_btm.n243 0.109875
R43478 C10_N_btm.n3492 C10_N_btm.n243 0.109875
R43479 C10_N_btm.n3487 C10_N_btm.n244 0.109875
R43480 C10_N_btm.n3489 C10_N_btm.n244 0.109875
R43481 C10_N_btm.n3484 C10_N_btm.n245 0.109875
R43482 C10_N_btm.n3486 C10_N_btm.n245 0.109875
R43483 C10_N_btm.n3481 C10_N_btm.n246 0.109875
R43484 C10_N_btm.n3483 C10_N_btm.n246 0.109875
R43485 C10_N_btm.n3478 C10_N_btm.n247 0.109875
R43486 C10_N_btm.n3480 C10_N_btm.n247 0.109875
R43487 C10_N_btm.n3475 C10_N_btm.n248 0.109875
R43488 C10_N_btm.n3477 C10_N_btm.n248 0.109875
R43489 C10_N_btm.n3472 C10_N_btm.n249 0.109875
R43490 C10_N_btm.n3474 C10_N_btm.n249 0.109875
R43491 C10_N_btm.n3469 C10_N_btm.n283 0.109875
R43492 C10_N_btm.n3471 C10_N_btm.n283 0.109875
R43493 C10_N_btm.n282 C10_N_btm.n251 0.109875
R43494 C10_N_btm.n282 C10_N_btm.n281 0.109875
R43495 C10_N_btm.n279 C10_N_btm.n252 0.109875
R43496 C10_N_btm.n277 C10_N_btm.n252 0.109875
R43497 C10_N_btm.n276 C10_N_btm.n253 0.109875
R43498 C10_N_btm.n274 C10_N_btm.n253 0.109875
R43499 C10_N_btm.n273 C10_N_btm.n254 0.109875
R43500 C10_N_btm.n271 C10_N_btm.n254 0.109875
R43501 C10_N_btm.n270 C10_N_btm.n255 0.109875
R43502 C10_N_btm.n268 C10_N_btm.n255 0.109875
R43503 C10_N_btm.n267 C10_N_btm.n256 0.109875
R43504 C10_N_btm.n265 C10_N_btm.n256 0.109875
R43505 C10_N_btm.n264 C10_N_btm.n257 0.109875
R43506 C10_N_btm.n262 C10_N_btm.n257 0.109875
R43507 C10_N_btm.n261 C10_N_btm.n258 0.109875
R43508 C10_N_btm.n259 C10_N_btm.n258 0.109875
R43509 C10_N_btm.n3502 C10_N_btm.n241 0.109875
R43510 C10_N_btm.n3502 C10_N_btm.n3501 0.109875
R43511 C10_N_btm.n3507 C10_N_btm.n3503 0.109875
R43512 C10_N_btm.n3505 C10_N_btm.n3503 0.109875
R43513 C10_N_btm.n3510 C10_N_btm.n239 0.109875
R43514 C10_N_btm.n3508 C10_N_btm.n239 0.109875
R43515 C10_N_btm.n3513 C10_N_btm.n238 0.109875
R43516 C10_N_btm.n3511 C10_N_btm.n238 0.109875
R43517 C10_N_btm.n3516 C10_N_btm.n237 0.109875
R43518 C10_N_btm.n3514 C10_N_btm.n237 0.109875
R43519 C10_N_btm.n3519 C10_N_btm.n236 0.109875
R43520 C10_N_btm.n3517 C10_N_btm.n236 0.109875
R43521 C10_N_btm.n3522 C10_N_btm.n235 0.109875
R43522 C10_N_btm.n3520 C10_N_btm.n235 0.109875
R43523 C10_N_btm.n3525 C10_N_btm.n234 0.109875
R43524 C10_N_btm.n3523 C10_N_btm.n234 0.109875
R43525 C10_N_btm.n3528 C10_N_btm.n233 0.109875
R43526 C10_N_btm.n3526 C10_N_btm.n233 0.109875
R43527 C10_N_btm.n3531 C10_N_btm.n232 0.109875
R43528 C10_N_btm.n3529 C10_N_btm.n232 0.109875
R43529 C10_N_btm.n3536 C10_N_btm.n230 0.109875
R43530 C10_N_btm.n3538 C10_N_btm.n230 0.109875
R43531 C10_N_btm.n3539 C10_N_btm.n196 0.109875
R43532 C10_N_btm.n3541 C10_N_btm.n196 0.109875
R43533 C10_N_btm.n3542 C10_N_btm.n195 0.109875
R43534 C10_N_btm.n3544 C10_N_btm.n195 0.109875
R43535 C10_N_btm.n3545 C10_N_btm.n194 0.109875
R43536 C10_N_btm.n3547 C10_N_btm.n194 0.109875
R43537 C10_N_btm.n3548 C10_N_btm.n193 0.109875
R43538 C10_N_btm.n3550 C10_N_btm.n193 0.109875
R43539 C10_N_btm.n3551 C10_N_btm.n192 0.109875
R43540 C10_N_btm.n3553 C10_N_btm.n192 0.109875
R43541 C10_N_btm.n3554 C10_N_btm.n191 0.109875
R43542 C10_N_btm.n3556 C10_N_btm.n191 0.109875
R43543 C10_N_btm.n3557 C10_N_btm.n190 0.109875
R43544 C10_N_btm.n3559 C10_N_btm.n190 0.109875
R43545 C10_N_btm.n3560 C10_N_btm.n187 0.109875
R43546 C10_N_btm.n3562 C10_N_btm.n187 0.109875
R43547 C10_N_btm.n3569 C10_N_btm.n188 0.109875
R43548 C10_N_btm.n3569 C10_N_btm.n3568 0.109875
R43549 C10_N_btm.n208 C10_N_btm.n205 0.109875
R43550 C10_N_btm.n206 C10_N_btm.n205 0.109875
R43551 C10_N_btm.n211 C10_N_btm.n204 0.109875
R43552 C10_N_btm.n209 C10_N_btm.n204 0.109875
R43553 C10_N_btm.n214 C10_N_btm.n203 0.109875
R43554 C10_N_btm.n212 C10_N_btm.n203 0.109875
R43555 C10_N_btm.n217 C10_N_btm.n202 0.109875
R43556 C10_N_btm.n215 C10_N_btm.n202 0.109875
R43557 C10_N_btm.n220 C10_N_btm.n201 0.109875
R43558 C10_N_btm.n218 C10_N_btm.n201 0.109875
R43559 C10_N_btm.n223 C10_N_btm.n200 0.109875
R43560 C10_N_btm.n221 C10_N_btm.n200 0.109875
R43561 C10_N_btm.n226 C10_N_btm.n199 0.109875
R43562 C10_N_btm.n224 C10_N_btm.n199 0.109875
R43563 C10_N_btm.n229 C10_N_btm.n198 0.109875
R43564 C10_N_btm.n229 C10_N_btm.n228 0.109875
R43565 C10_N_btm.n3598 C10_N_btm.n179 0.109875
R43566 C10_N_btm.n3596 C10_N_btm.n179 0.109875
R43567 C10_N_btm.n3595 C10_N_btm.n180 0.109875
R43568 C10_N_btm.n3593 C10_N_btm.n180 0.109875
R43569 C10_N_btm.n3592 C10_N_btm.n181 0.109875
R43570 C10_N_btm.n3590 C10_N_btm.n181 0.109875
R43571 C10_N_btm.n3589 C10_N_btm.n182 0.109875
R43572 C10_N_btm.n3587 C10_N_btm.n182 0.109875
R43573 C10_N_btm.n3586 C10_N_btm.n183 0.109875
R43574 C10_N_btm.n3584 C10_N_btm.n183 0.109875
R43575 C10_N_btm.n3583 C10_N_btm.n184 0.109875
R43576 C10_N_btm.n3581 C10_N_btm.n184 0.109875
R43577 C10_N_btm.n3580 C10_N_btm.n185 0.109875
R43578 C10_N_btm.n3578 C10_N_btm.n185 0.109875
R43579 C10_N_btm.n3577 C10_N_btm.n186 0.109875
R43580 C10_N_btm.n3575 C10_N_btm.n186 0.109875
R43581 C10_N_btm.n3574 C10_N_btm.n3570 0.109875
R43582 C10_N_btm.n3572 C10_N_btm.n3570 0.109875
R43583 C10_N_btm.n3627 C10_N_btm.n134 0.109875
R43584 C10_N_btm.n3629 C10_N_btm.n134 0.109875
R43585 C10_N_btm.n3624 C10_N_btm.n137 0.109875
R43586 C10_N_btm.n3626 C10_N_btm.n137 0.109875
R43587 C10_N_btm.n3621 C10_N_btm.n138 0.109875
R43588 C10_N_btm.n3623 C10_N_btm.n138 0.109875
R43589 C10_N_btm.n3618 C10_N_btm.n139 0.109875
R43590 C10_N_btm.n3620 C10_N_btm.n139 0.109875
R43591 C10_N_btm.n3615 C10_N_btm.n140 0.109875
R43592 C10_N_btm.n3617 C10_N_btm.n140 0.109875
R43593 C10_N_btm.n3612 C10_N_btm.n141 0.109875
R43594 C10_N_btm.n3614 C10_N_btm.n141 0.109875
R43595 C10_N_btm.n3609 C10_N_btm.n142 0.109875
R43596 C10_N_btm.n3611 C10_N_btm.n142 0.109875
R43597 C10_N_btm.n3606 C10_N_btm.n143 0.109875
R43598 C10_N_btm.n3608 C10_N_btm.n143 0.109875
R43599 C10_N_btm.n3603 C10_N_btm.n177 0.109875
R43600 C10_N_btm.n3605 C10_N_btm.n177 0.109875
R43601 C10_N_btm.n176 C10_N_btm.n145 0.109875
R43602 C10_N_btm.n176 C10_N_btm.n175 0.109875
R43603 C10_N_btm.n173 C10_N_btm.n146 0.109875
R43604 C10_N_btm.n171 C10_N_btm.n146 0.109875
R43605 C10_N_btm.n170 C10_N_btm.n147 0.109875
R43606 C10_N_btm.n168 C10_N_btm.n147 0.109875
R43607 C10_N_btm.n167 C10_N_btm.n148 0.109875
R43608 C10_N_btm.n165 C10_N_btm.n148 0.109875
R43609 C10_N_btm.n164 C10_N_btm.n149 0.109875
R43610 C10_N_btm.n162 C10_N_btm.n149 0.109875
R43611 C10_N_btm.n161 C10_N_btm.n150 0.109875
R43612 C10_N_btm.n159 C10_N_btm.n150 0.109875
R43613 C10_N_btm.n158 C10_N_btm.n151 0.109875
R43614 C10_N_btm.n156 C10_N_btm.n151 0.109875
R43615 C10_N_btm.n155 C10_N_btm.n152 0.109875
R43616 C10_N_btm.n153 C10_N_btm.n152 0.109875
R43617 C10_N_btm.n3636 C10_N_btm.n135 0.109875
R43618 C10_N_btm.n3636 C10_N_btm.n3635 0.109875
R43619 C10_N_btm.n3641 C10_N_btm.n3637 0.109875
R43620 C10_N_btm.n3639 C10_N_btm.n3637 0.109875
R43621 C10_N_btm.n3644 C10_N_btm.n133 0.109875
R43622 C10_N_btm.n3642 C10_N_btm.n133 0.109875
R43623 C10_N_btm.n3647 C10_N_btm.n132 0.109875
R43624 C10_N_btm.n3645 C10_N_btm.n132 0.109875
R43625 C10_N_btm.n3650 C10_N_btm.n131 0.109875
R43626 C10_N_btm.n3648 C10_N_btm.n131 0.109875
R43627 C10_N_btm.n3653 C10_N_btm.n130 0.109875
R43628 C10_N_btm.n3651 C10_N_btm.n130 0.109875
R43629 C10_N_btm.n3656 C10_N_btm.n129 0.109875
R43630 C10_N_btm.n3654 C10_N_btm.n129 0.109875
R43631 C10_N_btm.n3659 C10_N_btm.n128 0.109875
R43632 C10_N_btm.n3657 C10_N_btm.n128 0.109875
R43633 C10_N_btm.n3662 C10_N_btm.n127 0.109875
R43634 C10_N_btm.n3660 C10_N_btm.n127 0.109875
R43635 C10_N_btm.n3665 C10_N_btm.n126 0.109875
R43636 C10_N_btm.n3663 C10_N_btm.n126 0.109875
R43637 C10_N_btm.n3670 C10_N_btm.n124 0.109875
R43638 C10_N_btm.n3672 C10_N_btm.n124 0.109875
R43639 C10_N_btm.n3673 C10_N_btm.n90 0.109875
R43640 C10_N_btm.n3675 C10_N_btm.n90 0.109875
R43641 C10_N_btm.n3676 C10_N_btm.n89 0.109875
R43642 C10_N_btm.n3678 C10_N_btm.n89 0.109875
R43643 C10_N_btm.n3679 C10_N_btm.n88 0.109875
R43644 C10_N_btm.n3681 C10_N_btm.n88 0.109875
R43645 C10_N_btm.n3682 C10_N_btm.n87 0.109875
R43646 C10_N_btm.n3684 C10_N_btm.n87 0.109875
R43647 C10_N_btm.n3685 C10_N_btm.n86 0.109875
R43648 C10_N_btm.n3687 C10_N_btm.n86 0.109875
R43649 C10_N_btm.n3688 C10_N_btm.n85 0.109875
R43650 C10_N_btm.n3690 C10_N_btm.n85 0.109875
R43651 C10_N_btm.n3691 C10_N_btm.n84 0.109875
R43652 C10_N_btm.n3693 C10_N_btm.n84 0.109875
R43653 C10_N_btm.n3694 C10_N_btm.n81 0.109875
R43654 C10_N_btm.n3696 C10_N_btm.n81 0.109875
R43655 C10_N_btm.n3703 C10_N_btm.n82 0.109875
R43656 C10_N_btm.n3703 C10_N_btm.n3702 0.109875
R43657 C10_N_btm.n102 C10_N_btm.n99 0.109875
R43658 C10_N_btm.n100 C10_N_btm.n99 0.109875
R43659 C10_N_btm.n105 C10_N_btm.n98 0.109875
R43660 C10_N_btm.n103 C10_N_btm.n98 0.109875
R43661 C10_N_btm.n108 C10_N_btm.n97 0.109875
R43662 C10_N_btm.n106 C10_N_btm.n97 0.109875
R43663 C10_N_btm.n111 C10_N_btm.n96 0.109875
R43664 C10_N_btm.n109 C10_N_btm.n96 0.109875
R43665 C10_N_btm.n114 C10_N_btm.n95 0.109875
R43666 C10_N_btm.n112 C10_N_btm.n95 0.109875
R43667 C10_N_btm.n117 C10_N_btm.n94 0.109875
R43668 C10_N_btm.n115 C10_N_btm.n94 0.109875
R43669 C10_N_btm.n120 C10_N_btm.n93 0.109875
R43670 C10_N_btm.n118 C10_N_btm.n93 0.109875
R43671 C10_N_btm.n123 C10_N_btm.n92 0.109875
R43672 C10_N_btm.n123 C10_N_btm.n122 0.109875
R43673 C10_N_btm.n3732 C10_N_btm.n73 0.109875
R43674 C10_N_btm.n3730 C10_N_btm.n73 0.109875
R43675 C10_N_btm.n3729 C10_N_btm.n74 0.109875
R43676 C10_N_btm.n3727 C10_N_btm.n74 0.109875
R43677 C10_N_btm.n3726 C10_N_btm.n75 0.109875
R43678 C10_N_btm.n3724 C10_N_btm.n75 0.109875
R43679 C10_N_btm.n3723 C10_N_btm.n76 0.109875
R43680 C10_N_btm.n3721 C10_N_btm.n76 0.109875
R43681 C10_N_btm.n3720 C10_N_btm.n77 0.109875
R43682 C10_N_btm.n3718 C10_N_btm.n77 0.109875
R43683 C10_N_btm.n3717 C10_N_btm.n78 0.109875
R43684 C10_N_btm.n3715 C10_N_btm.n78 0.109875
R43685 C10_N_btm.n3714 C10_N_btm.n79 0.109875
R43686 C10_N_btm.n3712 C10_N_btm.n79 0.109875
R43687 C10_N_btm.n3711 C10_N_btm.n80 0.109875
R43688 C10_N_btm.n3709 C10_N_btm.n80 0.109875
R43689 C10_N_btm.n3708 C10_N_btm.n3704 0.109875
R43690 C10_N_btm.n3706 C10_N_btm.n3704 0.109875
R43691 C10_N_btm.n3796 C10_N_btm.n61 0.109875
R43692 C10_N_btm.n3798 C10_N_btm.n61 0.109875
R43693 C10_N_btm.n3793 C10_N_btm.n64 0.109875
R43694 C10_N_btm.n3795 C10_N_btm.n64 0.109875
R43695 C10_N_btm.n3790 C10_N_btm.n65 0.109875
R43696 C10_N_btm.n3792 C10_N_btm.n65 0.109875
R43697 C10_N_btm.n3787 C10_N_btm.n66 0.109875
R43698 C10_N_btm.n3789 C10_N_btm.n66 0.109875
R43699 C10_N_btm.n3784 C10_N_btm.n67 0.109875
R43700 C10_N_btm.n3786 C10_N_btm.n67 0.109875
R43701 C10_N_btm.n3781 C10_N_btm.n68 0.109875
R43702 C10_N_btm.n3783 C10_N_btm.n68 0.109875
R43703 C10_N_btm.n3778 C10_N_btm.n69 0.109875
R43704 C10_N_btm.n3780 C10_N_btm.n69 0.109875
R43705 C10_N_btm.n3775 C10_N_btm.n70 0.109875
R43706 C10_N_btm.n3777 C10_N_btm.n70 0.109875
R43707 C10_N_btm.n3772 C10_N_btm.n71 0.109875
R43708 C10_N_btm.n3774 C10_N_btm.n71 0.109875
R43709 C10_N_btm.n3767 C10_N_btm.n52 0.109875
R43710 C10_N_btm.n3765 C10_N_btm.n52 0.109875
R43711 C10_N_btm.n3764 C10_N_btm.n3737 0.109875
R43712 C10_N_btm.n3762 C10_N_btm.n3737 0.109875
R43713 C10_N_btm.n3761 C10_N_btm.n3738 0.109875
R43714 C10_N_btm.n3759 C10_N_btm.n3738 0.109875
R43715 C10_N_btm.n3758 C10_N_btm.n3739 0.109875
R43716 C10_N_btm.n3756 C10_N_btm.n3739 0.109875
R43717 C10_N_btm.n3755 C10_N_btm.n3740 0.109875
R43718 C10_N_btm.n3753 C10_N_btm.n3740 0.109875
R43719 C10_N_btm.n3752 C10_N_btm.n3741 0.109875
R43720 C10_N_btm.n3750 C10_N_btm.n3741 0.109875
R43721 C10_N_btm.n3749 C10_N_btm.n3742 0.109875
R43722 C10_N_btm.n3747 C10_N_btm.n3742 0.109875
R43723 C10_N_btm.n3746 C10_N_btm.n3743 0.109875
R43724 C10_N_btm.n3744 C10_N_btm.n3743 0.109875
R43725 C10_N_btm.n3805 C10_N_btm.n62 0.109875
R43726 C10_N_btm.n3805 C10_N_btm.n3804 0.109875
R43727 C10_N_btm.n3810 C10_N_btm.n3806 0.109875
R43728 C10_N_btm.n3808 C10_N_btm.n3806 0.109875
R43729 C10_N_btm.n3813 C10_N_btm.n60 0.109875
R43730 C10_N_btm.n3811 C10_N_btm.n60 0.109875
R43731 C10_N_btm.n3816 C10_N_btm.n59 0.109875
R43732 C10_N_btm.n3814 C10_N_btm.n59 0.109875
R43733 C10_N_btm.n3819 C10_N_btm.n58 0.109875
R43734 C10_N_btm.n3817 C10_N_btm.n58 0.109875
R43735 C10_N_btm.n3822 C10_N_btm.n57 0.109875
R43736 C10_N_btm.n3820 C10_N_btm.n57 0.109875
R43737 C10_N_btm.n3825 C10_N_btm.n56 0.109875
R43738 C10_N_btm.n3823 C10_N_btm.n56 0.109875
R43739 C10_N_btm.n3828 C10_N_btm.n55 0.109875
R43740 C10_N_btm.n3826 C10_N_btm.n55 0.109875
R43741 C10_N_btm.n3831 C10_N_btm.n54 0.109875
R43742 C10_N_btm.n3829 C10_N_btm.n54 0.109875
R43743 C10_N_btm.n3834 C10_N_btm.n53 0.109875
R43744 C10_N_btm.n3834 C10_N_btm.n3833 0.109875
R43745 C10_N_btm.n3837 C10_N_btm.n3835 0.109875
R43746 C10_N_btm.n3839 C10_N_btm.n3835 0.109875
R43747 C10_N_btm.n3840 C10_N_btm.n51 0.109875
R43748 C10_N_btm.n3842 C10_N_btm.n51 0.109875
R43749 C10_N_btm.n3843 C10_N_btm.n50 0.109875
R43750 C10_N_btm.n3845 C10_N_btm.n50 0.109875
R43751 C10_N_btm.n3846 C10_N_btm.n49 0.109875
R43752 C10_N_btm.n3848 C10_N_btm.n49 0.109875
R43753 C10_N_btm.n3849 C10_N_btm.n48 0.109875
R43754 C10_N_btm.n3851 C10_N_btm.n48 0.109875
R43755 C10_N_btm.n3852 C10_N_btm.n47 0.109875
R43756 C10_N_btm.n3854 C10_N_btm.n47 0.109875
R43757 C10_N_btm.n3855 C10_N_btm.n46 0.109875
R43758 C10_N_btm.n3857 C10_N_btm.n46 0.109875
R43759 C10_N_btm.n3858 C10_N_btm.n45 0.109875
R43760 C10_N_btm.n3860 C10_N_btm.n45 0.109875
R43761 C10_N_btm.n3861 C10_N_btm.n44 0.109875
R43762 C10_N_btm.n3863 C10_N_btm.n44 0.109875
R43763 C10_N_btm.n3870 C10_N_btm.n42 0.109875
R43764 C10_N_btm.n3868 C10_N_btm.n42 0.109875
R43765 C10_N_btm.n3873 C10_N_btm.n41 0.109875
R43766 C10_N_btm.n3871 C10_N_btm.n41 0.109875
R43767 C10_N_btm.n3876 C10_N_btm.n40 0.109875
R43768 C10_N_btm.n3874 C10_N_btm.n40 0.109875
R43769 C10_N_btm.n3879 C10_N_btm.n39 0.109875
R43770 C10_N_btm.n3877 C10_N_btm.n39 0.109875
R43771 C10_N_btm.n3882 C10_N_btm.n38 0.109875
R43772 C10_N_btm.n3880 C10_N_btm.n38 0.109875
R43773 C10_N_btm.n3885 C10_N_btm.n37 0.109875
R43774 C10_N_btm.n3883 C10_N_btm.n37 0.109875
R43775 C10_N_btm.n3888 C10_N_btm.n36 0.109875
R43776 C10_N_btm.n3886 C10_N_btm.n36 0.109875
R43777 C10_N_btm.n3891 C10_N_btm.n35 0.109875
R43778 C10_N_btm.n3889 C10_N_btm.n35 0.109875
R43779 C10_N_btm.n3894 C10_N_btm.n34 0.109875
R43780 C10_N_btm.n3892 C10_N_btm.n34 0.109875
R43781 C10_N_btm.n2528 C10_N_btm.n2527 0.0556875
R43782 C10_N_btm.n2093 C10_N_btm.n1969 0.0556875
R43783 C10_N_btm.n2721 C10_N_btm.n2720 0.0556875
R43784 C10_N_btm.n2533 C10_N_btm.n1662 0.0556875
R43785 C10_N_btm.n2911 C10_N_btm.n2910 0.0556875
R43786 C10_N_btm.n2723 C10_N_btm.n2722 0.0556875
R43787 C10_N_btm.n1723 C10_N_btm.n1598 0.0556875
R43788 C10_N_btm.n2913 C10_N_btm.n2912 0.0556875
R43789 C10_N_btm.n2918 C10_N_btm.n401 0.0556875
R43790 C10_N_btm.n3106 C10_N_btm.n3105 0.0556875
R43791 C10_N_btm.n948 C10_N_btm.n947 0.0556875
R43792 C10_N_btm.n921 C10_N_btm.n904 0.0556875
R43793 C10_N_btm.n982 C10_N_btm.n981 0.0556875
R43794 C10_N_btm.n953 C10_N_btm.n862 0.0556875
R43795 C10_N_btm.n1013 C10_N_btm.n1012 0.0556875
R43796 C10_N_btm.n984 C10_N_btm.n983 0.0556875
R43797 C10_N_btm.n870 C10_N_btm.n851 0.0556875
R43798 C10_N_btm.n1015 C10_N_btm.n1014 0.0556875
R43799 C10_N_btm.n1020 C10_N_btm.n809 0.0556875
R43800 C10_N_btm.n1049 C10_N_btm.n1048 0.0556875
R43801 C10_N_btm.n1051 C10_N_btm.n1050 0.0556875
R43802 C10_N_btm.n1080 C10_N_btm.n1079 0.0556875
R43803 C10_N_btm.n1082 C10_N_btm.n1081 0.0556875
R43804 C10_N_btm.n817 C10_N_btm.n798 0.0556875
R43805 C10_N_btm.n1116 C10_N_btm.n1115 0.0556875
R43806 C10_N_btm.n1087 C10_N_btm.n756 0.0556875
R43807 C10_N_btm.n1147 C10_N_btm.n1146 0.0556875
R43808 C10_N_btm.n1118 C10_N_btm.n1117 0.0556875
R43809 C10_N_btm.n764 C10_N_btm.n745 0.0556875
R43810 C10_N_btm.n1149 C10_N_btm.n1148 0.0556875
R43811 C10_N_btm.n1154 C10_N_btm.n703 0.0556875
R43812 C10_N_btm.n1183 C10_N_btm.n1182 0.0556875
R43813 C10_N_btm.n1185 C10_N_btm.n1184 0.0556875
R43814 C10_N_btm.n1214 C10_N_btm.n1213 0.0556875
R43815 C10_N_btm.n1216 C10_N_btm.n1215 0.0556875
R43816 C10_N_btm.n711 C10_N_btm.n692 0.0556875
R43817 C10_N_btm.n1250 C10_N_btm.n1249 0.0556875
R43818 C10_N_btm.n1221 C10_N_btm.n650 0.0556875
R43819 C10_N_btm.n1281 C10_N_btm.n1280 0.0556875
R43820 C10_N_btm.n1252 C10_N_btm.n1251 0.0556875
R43821 C10_N_btm.n658 C10_N_btm.n639 0.0556875
R43822 C10_N_btm.n1283 C10_N_btm.n1282 0.0556875
R43823 C10_N_btm.n1288 C10_N_btm.n597 0.0556875
R43824 C10_N_btm.n1317 C10_N_btm.n1316 0.0556875
R43825 C10_N_btm.n1319 C10_N_btm.n1318 0.0556875
R43826 C10_N_btm.n1348 C10_N_btm.n1347 0.0556875
R43827 C10_N_btm.n1350 C10_N_btm.n1349 0.0556875
R43828 C10_N_btm.n605 C10_N_btm.n586 0.0556875
R43829 C10_N_btm.n1384 C10_N_btm.n1383 0.0556875
R43830 C10_N_btm.n1355 C10_N_btm.n577 0.0556875
R43831 C10_N_btm.n1450 C10_N_btm.n1449 0.0556875
R43832 C10_N_btm.n1421 C10_N_btm.n1420 0.0556875
R43833 C10_N_btm.n1419 C10_N_btm.n1418 0.0556875
R43834 C10_N_btm.n1452 C10_N_btm.n1451 0.0556875
R43835 C10_N_btm.n1457 C10_N_btm.n557 0.0556875
R43836 C10_N_btm.n1386 C10_N_btm.n1385 0.0556875
R43837 C10_N_btm.n1486 C10_N_btm.n547 0.0556875
R43838 C10_N_btm.n1515 C10_N_btm.n1514 0.0556875
R43839 C10_N_btm.n1597 C10_N_btm.n1596 0.0556875
R43840 C10_N_btm.n3108 C10_N_btm.n3107 0.0556875
R43841 C10_N_btm.n3296 C10_N_btm.n3295 0.0556875
R43842 C10_N_btm.n3298 C10_N_btm.n3297 0.0556875
R43843 C10_N_btm.n3332 C10_N_btm.n3331 0.0556875
R43844 C10_N_btm.n3303 C10_N_btm.n348 0.0556875
R43845 C10_N_btm.n3363 C10_N_btm.n3362 0.0556875
R43846 C10_N_btm.n3334 C10_N_btm.n3333 0.0556875
R43847 C10_N_btm.n356 C10_N_btm.n337 0.0556875
R43848 C10_N_btm.n3365 C10_N_btm.n3364 0.0556875
R43849 C10_N_btm.n3370 C10_N_btm.n295 0.0556875
R43850 C10_N_btm.n3399 C10_N_btm.n3398 0.0556875
R43851 C10_N_btm.n3401 C10_N_btm.n3400 0.0556875
R43852 C10_N_btm.n3430 C10_N_btm.n3429 0.0556875
R43853 C10_N_btm.n3432 C10_N_btm.n3431 0.0556875
R43854 C10_N_btm.n303 C10_N_btm.n284 0.0556875
R43855 C10_N_btm.n3466 C10_N_btm.n3465 0.0556875
R43856 C10_N_btm.n3437 C10_N_btm.n242 0.0556875
R43857 C10_N_btm.n3497 C10_N_btm.n3496 0.0556875
R43858 C10_N_btm.n3468 C10_N_btm.n3467 0.0556875
R43859 C10_N_btm.n250 C10_N_btm.n231 0.0556875
R43860 C10_N_btm.n3499 C10_N_btm.n3498 0.0556875
R43861 C10_N_btm.n3504 C10_N_btm.n189 0.0556875
R43862 C10_N_btm.n3533 C10_N_btm.n3532 0.0556875
R43863 C10_N_btm.n3535 C10_N_btm.n3534 0.0556875
R43864 C10_N_btm.n3564 C10_N_btm.n3563 0.0556875
R43865 C10_N_btm.n3566 C10_N_btm.n3565 0.0556875
R43866 C10_N_btm.n197 C10_N_btm.n178 0.0556875
R43867 C10_N_btm.n3600 C10_N_btm.n3599 0.0556875
R43868 C10_N_btm.n3571 C10_N_btm.n136 0.0556875
R43869 C10_N_btm.n3631 C10_N_btm.n3630 0.0556875
R43870 C10_N_btm.n3602 C10_N_btm.n3601 0.0556875
R43871 C10_N_btm.n144 C10_N_btm.n125 0.0556875
R43872 C10_N_btm.n3633 C10_N_btm.n3632 0.0556875
R43873 C10_N_btm.n3638 C10_N_btm.n83 0.0556875
R43874 C10_N_btm.n3667 C10_N_btm.n3666 0.0556875
R43875 C10_N_btm.n3669 C10_N_btm.n3668 0.0556875
R43876 C10_N_btm.n3698 C10_N_btm.n3697 0.0556875
R43877 C10_N_btm.n3700 C10_N_btm.n3699 0.0556875
R43878 C10_N_btm.n91 C10_N_btm.n72 0.0556875
R43879 C10_N_btm.n3734 C10_N_btm.n3733 0.0556875
R43880 C10_N_btm.n3705 C10_N_btm.n63 0.0556875
R43881 C10_N_btm.n3800 C10_N_btm.n3799 0.0556875
R43882 C10_N_btm.n3771 C10_N_btm.n3770 0.0556875
R43883 C10_N_btm.n3769 C10_N_btm.n3768 0.0556875
R43884 C10_N_btm.n3802 C10_N_btm.n3801 0.0556875
R43885 C10_N_btm.n3807 C10_N_btm.n43 0.0556875
R43886 C10_N_btm.n3736 C10_N_btm.n3735 0.0556875
R43887 C10_N_btm.n3836 C10_N_btm.n33 0.0556875
R43888 C10_N_btm.n3865 C10_N_btm.n3864 0.0556875
R43889 C10_N_btm.n3867 C10_N_btm.n3866 0.0556875
R43890 C10_N_btm.n3896 C10_N_btm.n3895 0.0556875
R43891 a_n2810_44894.n9 a_n2810_44894.t11 1415.15
R43892 a_n2810_44894.n8 a_n2810_44894.t4 1330.32
R43893 a_n2810_44894.n2 a_n2810_44894.t5 1330.32
R43894 a_n2810_44894.n6 a_n2810_44894.t10 1330.32
R43895 a_n2810_44894.n7 a_n2810_44894.t7 1320.68
R43896 a_n2810_44894.n9 a_n2810_44894.t8 1320.68
R43897 a_n2810_44894.n5 a_n2810_44894.t9 1320.68
R43898 a_n2810_44894.n3 a_n2810_44894.t6 1320.68
R43899 a_n2810_44894.n11 a_n2810_44894.n0 296.139
R43900 a_n2810_44894.n12 a_n2810_44894.n11 269.182
R43901 a_n2810_44894.n4 a_n2810_44894.n3 161.78
R43902 a_n2810_44894.n7 a_n2810_44894.n1 161.3
R43903 a_n2810_44894.n5 a_n2810_44894.n4 161.3
R43904 a_n2810_44894.n10 a_n2810_44894.n9 161.3
R43905 a_n2810_44894.n11 a_n2810_44894.n10 119.445
R43906 a_n2810_44894.n9 a_n2810_44894.n8 84.8325
R43907 a_n2810_44894.n8 a_n2810_44894.n7 84.8325
R43908 a_n2810_44894.n3 a_n2810_44894.n2 84.8325
R43909 a_n2810_44894.n5 a_n2810_44894.n2 84.8325
R43910 a_n2810_44894.n6 a_n2810_44894.n5 84.8325
R43911 a_n2810_44894.n7 a_n2810_44894.n6 84.8325
R43912 a_n2810_44894.n0 a_n2810_44894.t2 26.5955
R43913 a_n2810_44894.n0 a_n2810_44894.t3 26.5955
R43914 a_n2810_44894.n12 a_n2810_44894.t0 24.9236
R43915 a_n2810_44894.t1 a_n2810_44894.n12 24.9236
R43916 a_n2810_44894.n4 a_n2810_44894.n1 0.4805
R43917 a_n2810_44894.n10 a_n2810_44894.n1 0.4655
R43918 a_9521_45982.n20 a_9521_45982.n0 659.109
R43919 a_9521_45982.n3 a_9521_45982.t4 294.557
R43920 a_9521_45982.n2 a_9521_45982.t7 294.557
R43921 a_9521_45982.n16 a_9521_45982.t23 294.557
R43922 a_9521_45982.n13 a_9521_45982.t5 294.557
R43923 a_9521_45982.n7 a_9521_45982.t20 294.557
R43924 a_9521_45982.n6 a_9521_45982.t17 294.557
R43925 a_9521_45982.n5 a_9521_45982.t15 294.557
R43926 a_9521_45982.n1 a_9521_45982.t13 294.557
R43927 a_9521_45982.n10 a_9521_45982.t19 229.001
R43928 a_9521_45982.n21 a_9521_45982.n20 219.663
R43929 a_9521_45982.n3 a_9521_45982.t14 211.01
R43930 a_9521_45982.n2 a_9521_45982.t21 211.01
R43931 a_9521_45982.n16 a_9521_45982.t9 211.01
R43932 a_9521_45982.n13 a_9521_45982.t18 211.01
R43933 a_9521_45982.n7 a_9521_45982.t22 211.01
R43934 a_9521_45982.n6 a_9521_45982.t12 211.01
R43935 a_9521_45982.n5 a_9521_45982.t11 211.01
R43936 a_9521_45982.n1 a_9521_45982.t10 211.01
R43937 a_9521_45982.n8 a_9521_45982.t16 196.549
R43938 a_9521_45982.n4 a_9521_45982.n3 180.172
R43939 a_9521_45982.n17 a_9521_45982.n16 179.678
R43940 a_9521_45982.n4 a_9521_45982.n2 178.101
R43941 a_9521_45982.n11 a_9521_45982.n10 176.357
R43942 a_9521_45982.n14 a_9521_45982.n13 174.832
R43943 a_9521_45982.n15 a_9521_45982.n5 169.666
R43944 a_9521_45982.n12 a_9521_45982.n6 168.923
R43945 a_9521_45982.n9 a_9521_45982.n8 167.506
R43946 a_9521_45982.n9 a_9521_45982.n7 165.95
R43947 a_9521_45982.n19 a_9521_45982.n1 162.585
R43948 a_9521_45982.n10 a_9521_45982.t6 156.702
R43949 a_9521_45982.n8 a_9521_45982.t8 148.35
R43950 a_9521_45982.t1 a_9521_45982.n21 38.5719
R43951 a_9521_45982.n21 a_9521_45982.t0 38.5719
R43952 a_9521_45982.n12 a_9521_45982.n11 28.5375
R43953 a_9521_45982.n0 a_9521_45982.t2 26.5955
R43954 a_9521_45982.n0 a_9521_45982.t3 26.5955
R43955 a_9521_45982.n11 a_9521_45982.n9 23.2599
R43956 a_9521_45982.n14 a_9521_45982.n12 10.4402
R43957 a_9521_45982.n20 a_9521_45982.n19 10.0713
R43958 a_9521_45982.n15 a_9521_45982.n14 9.50153
R43959 a_9521_45982.n18 a_9521_45982.n17 7.26492
R43960 a_9521_45982.n19 a_9521_45982.n18 6.07742
R43961 a_9521_45982.n18 a_9521_45982.n4 1.99363
R43962 a_9521_45982.n17 a_9521_45982.n15 1.69349
R43963 C8_P_btm C8_P_btm.n8 66.3755
R43964 C8_P_btm.n8 C8_P_btm.n7 43.4801
R43965 C8_P_btm.n2 C8_P_btm.n1 33.0333
R43966 C8_P_btm.n2 C8_P_btm.n0 32.3614
R43967 C8_P_btm.n4 C8_P_btm.n2 21.6828
R43968 C8_P_btm.n4 C8_P_btm.n3 20.8888
R43969 C8_P_btm.n6 C8_P_btm.n5 20.8766
R43970 C8_P_btm.n6 C8_P_btm.n4 11.2088
R43971 C8_P_btm.n7 C8_P_btm.t6 9.9005
R43972 C8_P_btm.n7 C8_P_btm.t7 9.9005
R43973 C8_P_btm.n8 C8_P_btm.n6 8.45883
R43974 C8_P_btm C8_P_btm.n903 6.68175
R43975 C8_P_btm.n10 C8_P_btm.t12 5.03712
R43976 C8_P_btm.n11 C8_P_btm.t17 5.03712
R43977 C8_P_btm.n12 C8_P_btm.t8 5.03712
R43978 C8_P_btm.n890 C8_P_btm.t9 5.03712
R43979 C8_P_btm.n503 C8_P_btm.t16 5.03712
R43980 C8_P_btm.n507 C8_P_btm.t11 5.03712
R43981 C8_P_btm.n506 C8_P_btm.t13 5.03712
R43982 C8_P_btm.n520 C8_P_btm.t10 5.03712
R43983 C8_P_btm.n516 C8_P_btm.t14 5.03712
R43984 C8_P_btm.n900 C8_P_btm.n899 4.60698
R43985 C8_P_btm.n899 C8_P_btm.n898 4.60698
R43986 C8_P_btm.n897 C8_P_btm.n896 4.60698
R43987 C8_P_btm.n896 C8_P_btm.n895 4.60698
R43988 C8_P_btm.n894 C8_P_btm.n893 4.60698
R43989 C8_P_btm.n893 C8_P_btm.n892 4.60698
R43990 C8_P_btm.n887 C8_P_btm.n886 4.60698
R43991 C8_P_btm.n886 C8_P_btm.n885 4.60698
R43992 C8_P_btm.n884 C8_P_btm.n883 4.60698
R43993 C8_P_btm.n883 C8_P_btm.n882 4.60698
R43994 C8_P_btm.n881 C8_P_btm.n880 4.60698
R43995 C8_P_btm.n880 C8_P_btm.n879 4.60698
R43996 C8_P_btm.n875 C8_P_btm.n874 4.60698
R43997 C8_P_btm.n874 C8_P_btm.n17 4.60698
R43998 C8_P_btm.n872 C8_P_btm.n871 4.60698
R43999 C8_P_btm.n873 C8_P_btm.n872 4.60698
R44000 C8_P_btm.n869 C8_P_btm.n868 4.60698
R44001 C8_P_btm.n870 C8_P_btm.n869 4.60698
R44002 C8_P_btm.n864 C8_P_btm.n863 4.60698
R44003 C8_P_btm.n863 C8_P_btm.n20 4.60698
R44004 C8_P_btm.n841 C8_P_btm.n840 4.60698
R44005 C8_P_btm.n842 C8_P_btm.n841 4.60698
R44006 C8_P_btm.n844 C8_P_btm.n843 4.60698
R44007 C8_P_btm.n845 C8_P_btm.n844 4.60698
R44008 C8_P_btm.n852 C8_P_btm.n851 4.60698
R44009 C8_P_btm.n851 C8_P_btm.n850 4.60698
R44010 C8_P_btm.n855 C8_P_btm.n854 4.60698
R44011 C8_P_btm.n854 C8_P_btm.n853 4.60698
R44012 C8_P_btm.n858 C8_P_btm.n857 4.60698
R44013 C8_P_btm.n857 C8_P_btm.n856 4.60698
R44014 C8_P_btm.n827 C8_P_btm.n826 4.60698
R44015 C8_P_btm.n828 C8_P_btm.n827 4.60698
R44016 C8_P_btm.n830 C8_P_btm.n829 4.60698
R44017 C8_P_btm.n831 C8_P_btm.n830 4.60698
R44018 C8_P_btm.n833 C8_P_btm.n832 4.60698
R44019 C8_P_btm.n834 C8_P_btm.n833 4.60698
R44020 C8_P_btm.n38 C8_P_btm.n37 4.60698
R44021 C8_P_btm.n37 C8_P_btm.n32 4.60698
R44022 C8_P_btm.n35 C8_P_btm.n34 4.60698
R44023 C8_P_btm.n36 C8_P_btm.n35 4.60698
R44024 C8_P_btm.n822 C8_P_btm.n821 4.60698
R44025 C8_P_btm.n821 C8_P_btm.n28 4.60698
R44026 C8_P_btm.n816 C8_P_btm.n815 4.60698
R44027 C8_P_btm.n815 C8_P_btm.n814 4.60698
R44028 C8_P_btm.n813 C8_P_btm.n812 4.60698
R44029 C8_P_btm.n812 C8_P_btm.n811 4.60698
R44030 C8_P_btm.n810 C8_P_btm.n809 4.60698
R44031 C8_P_btm.n809 C8_P_btm.n808 4.60698
R44032 C8_P_btm.n802 C8_P_btm.n801 4.60698
R44033 C8_P_btm.n803 C8_P_btm.n802 4.60698
R44034 C8_P_btm.n799 C8_P_btm.n798 4.60698
R44035 C8_P_btm.n800 C8_P_btm.n799 4.60698
R44036 C8_P_btm.n796 C8_P_btm.n795 4.60698
R44037 C8_P_btm.n797 C8_P_btm.n796 4.60698
R44038 C8_P_btm.n791 C8_P_btm.n790 4.60698
R44039 C8_P_btm.n790 C8_P_btm.n45 4.60698
R44040 C8_P_btm.n52 C8_P_btm.n51 4.60698
R44041 C8_P_btm.n53 C8_P_btm.n52 4.60698
R44042 C8_P_btm.n55 C8_P_btm.n54 4.60698
R44043 C8_P_btm.n54 C8_P_btm.n49 4.60698
R44044 C8_P_btm.n779 C8_P_btm.n778 4.60698
R44045 C8_P_btm.n778 C8_P_btm.n777 4.60698
R44046 C8_P_btm.n782 C8_P_btm.n781 4.60698
R44047 C8_P_btm.n781 C8_P_btm.n780 4.60698
R44048 C8_P_btm.n785 C8_P_btm.n784 4.60698
R44049 C8_P_btm.n784 C8_P_btm.n783 4.60698
R44050 C8_P_btm.n765 C8_P_btm.n764 4.60698
R44051 C8_P_btm.n766 C8_P_btm.n765 4.60698
R44052 C8_P_btm.n768 C8_P_btm.n767 4.60698
R44053 C8_P_btm.n769 C8_P_btm.n768 4.60698
R44054 C8_P_btm.n771 C8_P_btm.n770 4.60698
R44055 C8_P_btm.n772 C8_P_btm.n771 4.60698
R44056 C8_P_btm.n79 C8_P_btm.n78 4.60698
R44057 C8_P_btm.n78 C8_P_btm.n77 4.60698
R44058 C8_P_btm.n75 C8_P_btm.n74 4.60698
R44059 C8_P_btm.n76 C8_P_btm.n75 4.60698
R44060 C8_P_btm.n72 C8_P_btm.n71 4.60698
R44061 C8_P_btm.n73 C8_P_btm.n72 4.60698
R44062 C8_P_btm.n760 C8_P_btm.n759 4.60698
R44063 C8_P_btm.n759 C8_P_btm.n62 4.60698
R44064 C8_P_btm.n754 C8_P_btm.n753 4.60698
R44065 C8_P_btm.n753 C8_P_btm.n752 4.60698
R44066 C8_P_btm.n751 C8_P_btm.n750 4.60698
R44067 C8_P_btm.n750 C8_P_btm.n749 4.60698
R44068 C8_P_btm.n748 C8_P_btm.n747 4.60698
R44069 C8_P_btm.n747 C8_P_btm.n746 4.60698
R44070 C8_P_btm.n745 C8_P_btm.n744 4.60698
R44071 C8_P_btm.n744 C8_P_btm.n743 4.60698
R44072 C8_P_btm.n742 C8_P_btm.n741 4.60698
R44073 C8_P_btm.n741 C8_P_btm.n740 4.60698
R44074 C8_P_btm.n738 C8_P_btm.n737 4.60698
R44075 C8_P_btm.n739 C8_P_btm.n738 4.60698
R44076 C8_P_btm.n82 C8_P_btm.n81 4.60698
R44077 C8_P_btm.n81 C8_P_btm.n80 4.60698
R44078 C8_P_btm.n735 C8_P_btm.n734 4.60698
R44079 C8_P_btm.n736 C8_P_btm.n735 4.60698
R44080 C8_P_btm.n732 C8_P_btm.n731 4.60698
R44081 C8_P_btm.n733 C8_P_btm.n732 4.60698
R44082 C8_P_btm.n729 C8_P_btm.n728 4.60698
R44083 C8_P_btm.n730 C8_P_btm.n729 4.60698
R44084 C8_P_btm.n726 C8_P_btm.n725 4.60698
R44085 C8_P_btm.n727 C8_P_btm.n726 4.60698
R44086 C8_P_btm.n723 C8_P_btm.n722 4.60698
R44087 C8_P_btm.n724 C8_P_btm.n723 4.60698
R44088 C8_P_btm.n720 C8_P_btm.n719 4.60698
R44089 C8_P_btm.n721 C8_P_btm.n720 4.60698
R44090 C8_P_btm.n717 C8_P_btm.n716 4.60698
R44091 C8_P_btm.n718 C8_P_btm.n717 4.60698
R44092 C8_P_btm.n714 C8_P_btm.n713 4.60698
R44093 C8_P_btm.n715 C8_P_btm.n714 4.60698
R44094 C8_P_btm.n711 C8_P_btm.n710 4.60698
R44095 C8_P_btm.n712 C8_P_btm.n711 4.60698
R44096 C8_P_btm.n708 C8_P_btm.n707 4.60698
R44097 C8_P_btm.n709 C8_P_btm.n708 4.60698
R44098 C8_P_btm.n705 C8_P_btm.n704 4.60698
R44099 C8_P_btm.n706 C8_P_btm.n705 4.60698
R44100 C8_P_btm.n702 C8_P_btm.n701 4.60698
R44101 C8_P_btm.n703 C8_P_btm.n702 4.60698
R44102 C8_P_btm.n699 C8_P_btm.n698 4.60698
R44103 C8_P_btm.n700 C8_P_btm.n699 4.60698
R44104 C8_P_btm.n696 C8_P_btm.n695 4.60698
R44105 C8_P_btm.n697 C8_P_btm.n696 4.60698
R44106 C8_P_btm.n693 C8_P_btm.n692 4.60698
R44107 C8_P_btm.n694 C8_P_btm.n693 4.60698
R44108 C8_P_btm.n690 C8_P_btm.n689 4.60698
R44109 C8_P_btm.n691 C8_P_btm.n690 4.60698
R44110 C8_P_btm.n688 C8_P_btm.n687 4.60698
R44111 C8_P_btm.n687 C8_P_btm.n686 4.60698
R44112 C8_P_btm.n685 C8_P_btm.n684 4.60698
R44113 C8_P_btm.n684 C8_P_btm.n683 4.60698
R44114 C8_P_btm.n682 C8_P_btm.n681 4.60698
R44115 C8_P_btm.n681 C8_P_btm.n680 4.60698
R44116 C8_P_btm.n679 C8_P_btm.n678 4.60698
R44117 C8_P_btm.n678 C8_P_btm.n677 4.60698
R44118 C8_P_btm.n676 C8_P_btm.n675 4.60698
R44119 C8_P_btm.n675 C8_P_btm.n674 4.60698
R44120 C8_P_btm.n673 C8_P_btm.n672 4.60698
R44121 C8_P_btm.n672 C8_P_btm.n671 4.60698
R44122 C8_P_btm.n665 C8_P_btm.n664 4.60698
R44123 C8_P_btm.n666 C8_P_btm.n665 4.60698
R44124 C8_P_btm.n662 C8_P_btm.n661 4.60698
R44125 C8_P_btm.n663 C8_P_btm.n662 4.60698
R44126 C8_P_btm.n659 C8_P_btm.n658 4.60698
R44127 C8_P_btm.n660 C8_P_btm.n659 4.60698
R44128 C8_P_btm.n656 C8_P_btm.n655 4.60698
R44129 C8_P_btm.n657 C8_P_btm.n656 4.60698
R44130 C8_P_btm.n646 C8_P_btm.n645 4.60698
R44131 C8_P_btm.n645 C8_P_btm.n644 4.60698
R44132 C8_P_btm.n643 C8_P_btm.n642 4.60698
R44133 C8_P_btm.n642 C8_P_btm.n641 4.60698
R44134 C8_P_btm.n640 C8_P_btm.n639 4.60698
R44135 C8_P_btm.n639 C8_P_btm.n638 4.60698
R44136 C8_P_btm.n634 C8_P_btm.n633 4.60698
R44137 C8_P_btm.n633 C8_P_btm.n462 4.60698
R44138 C8_P_btm.n631 C8_P_btm.n630 4.60698
R44139 C8_P_btm.n632 C8_P_btm.n631 4.60698
R44140 C8_P_btm.n628 C8_P_btm.n627 4.60698
R44141 C8_P_btm.n629 C8_P_btm.n628 4.60698
R44142 C8_P_btm.n623 C8_P_btm.n622 4.60698
R44143 C8_P_btm.n622 C8_P_btm.n465 4.60698
R44144 C8_P_btm.n600 C8_P_btm.n599 4.60698
R44145 C8_P_btm.n601 C8_P_btm.n600 4.60698
R44146 C8_P_btm.n603 C8_P_btm.n602 4.60698
R44147 C8_P_btm.n604 C8_P_btm.n603 4.60698
R44148 C8_P_btm.n611 C8_P_btm.n610 4.60698
R44149 C8_P_btm.n610 C8_P_btm.n609 4.60698
R44150 C8_P_btm.n614 C8_P_btm.n613 4.60698
R44151 C8_P_btm.n613 C8_P_btm.n612 4.60698
R44152 C8_P_btm.n617 C8_P_btm.n616 4.60698
R44153 C8_P_btm.n616 C8_P_btm.n615 4.60698
R44154 C8_P_btm.n586 C8_P_btm.n585 4.60698
R44155 C8_P_btm.n587 C8_P_btm.n586 4.60698
R44156 C8_P_btm.n589 C8_P_btm.n588 4.60698
R44157 C8_P_btm.n590 C8_P_btm.n589 4.60698
R44158 C8_P_btm.n592 C8_P_btm.n591 4.60698
R44159 C8_P_btm.n593 C8_P_btm.n592 4.60698
R44160 C8_P_btm.n483 C8_P_btm.n482 4.60698
R44161 C8_P_btm.n482 C8_P_btm.n477 4.60698
R44162 C8_P_btm.n480 C8_P_btm.n479 4.60698
R44163 C8_P_btm.n481 C8_P_btm.n480 4.60698
R44164 C8_P_btm.n581 C8_P_btm.n580 4.60698
R44165 C8_P_btm.n580 C8_P_btm.n473 4.60698
R44166 C8_P_btm.n575 C8_P_btm.n574 4.60698
R44167 C8_P_btm.n574 C8_P_btm.n573 4.60698
R44168 C8_P_btm.n572 C8_P_btm.n571 4.60698
R44169 C8_P_btm.n571 C8_P_btm.n570 4.60698
R44170 C8_P_btm.n569 C8_P_btm.n568 4.60698
R44171 C8_P_btm.n568 C8_P_btm.n567 4.60698
R44172 C8_P_btm.n561 C8_P_btm.n560 4.60698
R44173 C8_P_btm.n562 C8_P_btm.n561 4.60698
R44174 C8_P_btm.n558 C8_P_btm.n557 4.60698
R44175 C8_P_btm.n559 C8_P_btm.n558 4.60698
R44176 C8_P_btm.n555 C8_P_btm.n554 4.60698
R44177 C8_P_btm.n556 C8_P_btm.n555 4.60698
R44178 C8_P_btm.n550 C8_P_btm.n549 4.60698
R44179 C8_P_btm.n549 C8_P_btm.n490 4.60698
R44180 C8_P_btm.n497 C8_P_btm.n496 4.60698
R44181 C8_P_btm.n498 C8_P_btm.n497 4.60698
R44182 C8_P_btm.n500 C8_P_btm.n499 4.60698
R44183 C8_P_btm.n499 C8_P_btm.n494 4.60698
R44184 C8_P_btm.n538 C8_P_btm.n537 4.60698
R44185 C8_P_btm.n537 C8_P_btm.n536 4.60698
R44186 C8_P_btm.n541 C8_P_btm.n540 4.60698
R44187 C8_P_btm.n540 C8_P_btm.n539 4.60698
R44188 C8_P_btm.n544 C8_P_btm.n543 4.60698
R44189 C8_P_btm.n543 C8_P_btm.n542 4.60698
R44190 C8_P_btm.n524 C8_P_btm.n523 4.60698
R44191 C8_P_btm.n525 C8_P_btm.n524 4.60698
R44192 C8_P_btm.n527 C8_P_btm.n526 4.60698
R44193 C8_P_btm.n528 C8_P_btm.n527 4.60698
R44194 C8_P_btm.n530 C8_P_btm.n529 4.60698
R44195 C8_P_btm.n531 C8_P_btm.n530 4.60698
R44196 C8_P_btm.n510 C8_P_btm.n509 4.60698
R44197 C8_P_btm.n511 C8_P_btm.n510 4.60698
R44198 C8_P_btm.n513 C8_P_btm.n512 4.60698
R44199 C8_P_btm.n514 C8_P_btm.n513 4.60698
R44200 C8_P_btm.n518 C8_P_btm.n515 4.60698
R44201 C8_P_btm.n519 C8_P_btm.n518 4.60698
R44202 C8_P_btm.n654 C8_P_btm.n653 4.60698
R44203 C8_P_btm.n653 C8_P_btm.n652 4.60698
R44204 C8_P_btm.n450 C8_P_btm.n449 4.60698
R44205 C8_P_btm.n451 C8_P_btm.n450 4.60698
R44206 C8_P_btm.n447 C8_P_btm.n446 4.60698
R44207 C8_P_btm.n448 C8_P_btm.n447 4.60698
R44208 C8_P_btm.n444 C8_P_btm.n443 4.60698
R44209 C8_P_btm.n445 C8_P_btm.n444 4.60698
R44210 C8_P_btm.n441 C8_P_btm.n440 4.60698
R44211 C8_P_btm.n442 C8_P_btm.n441 4.60698
R44212 C8_P_btm.n438 C8_P_btm.n437 4.60698
R44213 C8_P_btm.n439 C8_P_btm.n438 4.60698
R44214 C8_P_btm.n435 C8_P_btm.n434 4.60698
R44215 C8_P_btm.n436 C8_P_btm.n435 4.60698
R44216 C8_P_btm.n432 C8_P_btm.n431 4.60698
R44217 C8_P_btm.n433 C8_P_btm.n432 4.60698
R44218 C8_P_btm.n429 C8_P_btm.n428 4.60698
R44219 C8_P_btm.n430 C8_P_btm.n429 4.60698
R44220 C8_P_btm.n426 C8_P_btm.n425 4.60698
R44221 C8_P_btm.n427 C8_P_btm.n426 4.60698
R44222 C8_P_btm.n423 C8_P_btm.n422 4.60698
R44223 C8_P_btm.n424 C8_P_btm.n423 4.60698
R44224 C8_P_btm.n420 C8_P_btm.n419 4.60698
R44225 C8_P_btm.n421 C8_P_btm.n420 4.60698
R44226 C8_P_btm.n417 C8_P_btm.n416 4.60698
R44227 C8_P_btm.n418 C8_P_btm.n417 4.60698
R44228 C8_P_btm.n414 C8_P_btm.n413 4.60698
R44229 C8_P_btm.n415 C8_P_btm.n414 4.60698
R44230 C8_P_btm.n411 C8_P_btm.n410 4.60698
R44231 C8_P_btm.n412 C8_P_btm.n411 4.60698
R44232 C8_P_btm.n408 C8_P_btm.n407 4.60698
R44233 C8_P_btm.n409 C8_P_btm.n408 4.60698
R44234 C8_P_btm.n405 C8_P_btm.n404 4.60698
R44235 C8_P_btm.n406 C8_P_btm.n405 4.60698
R44236 C8_P_btm.n402 C8_P_btm.n401 4.60698
R44237 C8_P_btm.n403 C8_P_btm.n402 4.60698
R44238 C8_P_btm.n399 C8_P_btm.n398 4.60698
R44239 C8_P_btm.n400 C8_P_btm.n399 4.60698
R44240 C8_P_btm.n396 C8_P_btm.n395 4.60698
R44241 C8_P_btm.n397 C8_P_btm.n396 4.60698
R44242 C8_P_btm.n393 C8_P_btm.n392 4.60698
R44243 C8_P_btm.n394 C8_P_btm.n393 4.60698
R44244 C8_P_btm.n390 C8_P_btm.n389 4.60698
R44245 C8_P_btm.n391 C8_P_btm.n390 4.60698
R44246 C8_P_btm.n387 C8_P_btm.n386 4.60698
R44247 C8_P_btm.n388 C8_P_btm.n387 4.60698
R44248 C8_P_btm.n384 C8_P_btm.n383 4.60698
R44249 C8_P_btm.n385 C8_P_btm.n384 4.60698
R44250 C8_P_btm.n381 C8_P_btm.n380 4.60698
R44251 C8_P_btm.n382 C8_P_btm.n381 4.60698
R44252 C8_P_btm.n378 C8_P_btm.n377 4.60698
R44253 C8_P_btm.n379 C8_P_btm.n378 4.60698
R44254 C8_P_btm.n375 C8_P_btm.n374 4.60698
R44255 C8_P_btm.n376 C8_P_btm.n375 4.60698
R44256 C8_P_btm.n372 C8_P_btm.n371 4.60698
R44257 C8_P_btm.n373 C8_P_btm.n372 4.60698
R44258 C8_P_btm.n369 C8_P_btm.n368 4.60698
R44259 C8_P_btm.n370 C8_P_btm.n369 4.60698
R44260 C8_P_btm.n364 C8_P_btm.n363 4.60698
R44261 C8_P_btm.n363 C8_P_btm.n136 4.60698
R44262 C8_P_btm.n194 C8_P_btm.n193 4.60698
R44263 C8_P_btm.n195 C8_P_btm.n194 4.60698
R44264 C8_P_btm.n197 C8_P_btm.n196 4.60698
R44265 C8_P_btm.n198 C8_P_btm.n197 4.60698
R44266 C8_P_btm.n200 C8_P_btm.n199 4.60698
R44267 C8_P_btm.n201 C8_P_btm.n200 4.60698
R44268 C8_P_btm.n203 C8_P_btm.n202 4.60698
R44269 C8_P_btm.n204 C8_P_btm.n203 4.60698
R44270 C8_P_btm.n206 C8_P_btm.n205 4.60698
R44271 C8_P_btm.n207 C8_P_btm.n206 4.60698
R44272 C8_P_btm.n209 C8_P_btm.n208 4.60698
R44273 C8_P_btm.n210 C8_P_btm.n209 4.60698
R44274 C8_P_btm.n212 C8_P_btm.n211 4.60698
R44275 C8_P_btm.n213 C8_P_btm.n212 4.60698
R44276 C8_P_btm.n215 C8_P_btm.n214 4.60698
R44277 C8_P_btm.n216 C8_P_btm.n215 4.60698
R44278 C8_P_btm.n218 C8_P_btm.n217 4.60698
R44279 C8_P_btm.n219 C8_P_btm.n218 4.60698
R44280 C8_P_btm.n221 C8_P_btm.n220 4.60698
R44281 C8_P_btm.n222 C8_P_btm.n221 4.60698
R44282 C8_P_btm.n224 C8_P_btm.n223 4.60698
R44283 C8_P_btm.n225 C8_P_btm.n224 4.60698
R44284 C8_P_btm.n227 C8_P_btm.n226 4.60698
R44285 C8_P_btm.n228 C8_P_btm.n227 4.60698
R44286 C8_P_btm.n230 C8_P_btm.n229 4.60698
R44287 C8_P_btm.n231 C8_P_btm.n230 4.60698
R44288 C8_P_btm.n233 C8_P_btm.n232 4.60698
R44289 C8_P_btm.n234 C8_P_btm.n233 4.60698
R44290 C8_P_btm.n236 C8_P_btm.n235 4.60698
R44291 C8_P_btm.n237 C8_P_btm.n236 4.60698
R44292 C8_P_btm.n239 C8_P_btm.n238 4.60698
R44293 C8_P_btm.n240 C8_P_btm.n239 4.60698
R44294 C8_P_btm.n242 C8_P_btm.n241 4.60698
R44295 C8_P_btm.n243 C8_P_btm.n242 4.60698
R44296 C8_P_btm.n245 C8_P_btm.n244 4.60698
R44297 C8_P_btm.n246 C8_P_btm.n245 4.60698
R44298 C8_P_btm.n248 C8_P_btm.n247 4.60698
R44299 C8_P_btm.n249 C8_P_btm.n248 4.60698
R44300 C8_P_btm.n251 C8_P_btm.n250 4.60698
R44301 C8_P_btm.n252 C8_P_btm.n251 4.60698
R44302 C8_P_btm.n254 C8_P_btm.n253 4.60698
R44303 C8_P_btm.n255 C8_P_btm.n254 4.60698
R44304 C8_P_btm.n257 C8_P_btm.n256 4.60698
R44305 C8_P_btm.n258 C8_P_btm.n257 4.60698
R44306 C8_P_btm.n260 C8_P_btm.n259 4.60698
R44307 C8_P_btm.n261 C8_P_btm.n260 4.60698
R44308 C8_P_btm.n263 C8_P_btm.n262 4.60698
R44309 C8_P_btm.n264 C8_P_btm.n263 4.60698
R44310 C8_P_btm.n266 C8_P_btm.n265 4.60698
R44311 C8_P_btm.n267 C8_P_btm.n266 4.60698
R44312 C8_P_btm.n269 C8_P_btm.n268 4.60698
R44313 C8_P_btm.n270 C8_P_btm.n269 4.60698
R44314 C8_P_btm.n272 C8_P_btm.n271 4.60698
R44315 C8_P_btm.n271 C8_P_btm.n166 4.60698
R44316 C8_P_btm.n278 C8_P_btm.n277 4.60698
R44317 C8_P_btm.n277 C8_P_btm.n276 4.60698
R44318 C8_P_btm.n281 C8_P_btm.n280 4.60698
R44319 C8_P_btm.n280 C8_P_btm.n279 4.60698
R44320 C8_P_btm.n284 C8_P_btm.n283 4.60698
R44321 C8_P_btm.n283 C8_P_btm.n282 4.60698
R44322 C8_P_btm.n287 C8_P_btm.n286 4.60698
R44323 C8_P_btm.n286 C8_P_btm.n285 4.60698
R44324 C8_P_btm.n290 C8_P_btm.n289 4.60698
R44325 C8_P_btm.n289 C8_P_btm.n288 4.60698
R44326 C8_P_btm.n293 C8_P_btm.n292 4.60698
R44327 C8_P_btm.n292 C8_P_btm.n291 4.60698
R44328 C8_P_btm.n296 C8_P_btm.n295 4.60698
R44329 C8_P_btm.n295 C8_P_btm.n294 4.60698
R44330 C8_P_btm.n299 C8_P_btm.n298 4.60698
R44331 C8_P_btm.n298 C8_P_btm.n297 4.60698
R44332 C8_P_btm.n302 C8_P_btm.n301 4.60698
R44333 C8_P_btm.n301 C8_P_btm.n300 4.60698
R44334 C8_P_btm.n305 C8_P_btm.n304 4.60698
R44335 C8_P_btm.n304 C8_P_btm.n303 4.60698
R44336 C8_P_btm.n308 C8_P_btm.n307 4.60698
R44337 C8_P_btm.n307 C8_P_btm.n306 4.60698
R44338 C8_P_btm.n311 C8_P_btm.n310 4.60698
R44339 C8_P_btm.n310 C8_P_btm.n309 4.60698
R44340 C8_P_btm.n314 C8_P_btm.n313 4.60698
R44341 C8_P_btm.n313 C8_P_btm.n312 4.60698
R44342 C8_P_btm.n317 C8_P_btm.n316 4.60698
R44343 C8_P_btm.n316 C8_P_btm.n315 4.60698
R44344 C8_P_btm.n320 C8_P_btm.n319 4.60698
R44345 C8_P_btm.n319 C8_P_btm.n318 4.60698
R44346 C8_P_btm.n323 C8_P_btm.n322 4.60698
R44347 C8_P_btm.n322 C8_P_btm.n321 4.60698
R44348 C8_P_btm.n326 C8_P_btm.n325 4.60698
R44349 C8_P_btm.n325 C8_P_btm.n324 4.60698
R44350 C8_P_btm.n329 C8_P_btm.n328 4.60698
R44351 C8_P_btm.n328 C8_P_btm.n327 4.60698
R44352 C8_P_btm.n332 C8_P_btm.n331 4.60698
R44353 C8_P_btm.n331 C8_P_btm.n330 4.60698
R44354 C8_P_btm.n335 C8_P_btm.n334 4.60698
R44355 C8_P_btm.n334 C8_P_btm.n333 4.60698
R44356 C8_P_btm.n338 C8_P_btm.n337 4.60698
R44357 C8_P_btm.n337 C8_P_btm.n336 4.60698
R44358 C8_P_btm.n341 C8_P_btm.n340 4.60698
R44359 C8_P_btm.n340 C8_P_btm.n339 4.60698
R44360 C8_P_btm.n344 C8_P_btm.n343 4.60698
R44361 C8_P_btm.n343 C8_P_btm.n342 4.60698
R44362 C8_P_btm.n347 C8_P_btm.n346 4.60698
R44363 C8_P_btm.n346 C8_P_btm.n345 4.60698
R44364 C8_P_btm.n350 C8_P_btm.n349 4.60698
R44365 C8_P_btm.n349 C8_P_btm.n348 4.60698
R44366 C8_P_btm.n353 C8_P_btm.n352 4.60698
R44367 C8_P_btm.n352 C8_P_btm.n351 4.60698
R44368 C8_P_btm.n356 C8_P_btm.n355 4.60698
R44369 C8_P_btm.n355 C8_P_btm.n354 4.60698
R44370 C8_P_btm.n359 C8_P_btm.n358 4.60698
R44371 C8_P_btm.n358 C8_P_btm.n357 4.60698
R44372 C8_P_btm.n903 C8_P_btm.t15 4.03712
R44373 C8_P_btm.n901 C8_P_btm.t196 3.98193
R44374 C8_P_btm.n891 C8_P_btm.t264 3.98193
R44375 C8_P_btm.n878 C8_P_btm.t254 3.98193
R44376 C8_P_btm.n837 C8_P_btm.t46 3.98193
R44377 C8_P_btm.n846 C8_P_btm.t88 3.98193
R44378 C8_P_btm.n849 C8_P_btm.t63 3.98193
R44379 C8_P_btm.n835 C8_P_btm.t44 3.98193
R44380 C8_P_btm.n31 C8_P_btm.t127 3.98193
R44381 C8_P_btm.n807 C8_P_btm.t106 3.98193
R44382 C8_P_btm.n804 C8_P_btm.t195 3.98193
R44383 C8_P_btm.n48 C8_P_btm.t170 3.98193
R44384 C8_P_btm.n776 C8_P_btm.t145 3.98193
R44385 C8_P_btm.n773 C8_P_btm.t239 3.98193
R44386 C8_P_btm.n83 C8_P_btm.t202 3.98193
R44387 C8_P_btm.n670 C8_P_btm.t191 3.98193
R44388 C8_P_btm.n667 C8_P_btm.t227 3.98193
R44389 C8_P_btm.n637 C8_P_btm.t257 3.98193
R44390 C8_P_btm.n596 C8_P_btm.t158 3.98193
R44391 C8_P_btm.n605 C8_P_btm.t181 3.98193
R44392 C8_P_btm.n608 C8_P_btm.t209 3.98193
R44393 C8_P_btm.n594 C8_P_btm.t246 3.98193
R44394 C8_P_btm.n476 C8_P_btm.t141 3.98193
R44395 C8_P_btm.n566 C8_P_btm.t234 3.98193
R44396 C8_P_btm.n563 C8_P_btm.t77 3.98193
R44397 C8_P_btm.n493 C8_P_btm.t99 3.98193
R44398 C8_P_btm.n535 C8_P_btm.t38 3.98193
R44399 C8_P_btm.n532 C8_P_btm.t37 3.98193
R44400 C8_P_btm.n508 C8_P_btm.t211 3.98193
R44401 C8_P_btm.n517 C8_P_btm.t115 3.98193
R44402 C8_P_btm.n522 C8_P_btm.t198 3.98193
R44403 C8_P_btm.n545 C8_P_btm.t173 3.98193
R44404 C8_P_btm.n548 C8_P_btm.t93 3.98193
R44405 C8_P_btm.n553 C8_P_btm.t241 3.98193
R44406 C8_P_btm.n576 C8_P_btm.t218 3.98193
R44407 C8_P_btm.n579 C8_P_btm.t50 3.98193
R44408 C8_P_btm.n584 C8_P_btm.t102 3.98193
R44409 C8_P_btm.n618 C8_P_btm.t112 3.98193
R44410 C8_P_btm.n621 C8_P_btm.t41 3.98193
R44411 C8_P_btm.n626 C8_P_btm.t60 3.98193
R44412 C8_P_btm.n647 C8_P_btm.t146 3.98193
R44413 C8_P_btm.n651 C8_P_btm.t126 3.98193
R44414 C8_P_btm.n452 C8_P_btm.t31 3.98193
R44415 C8_P_btm.n165 C8_P_btm.t110 3.98193
R44416 C8_P_btm.n275 C8_P_btm.t261 3.98193
R44417 C8_P_btm.n151 C8_P_btm.t84 3.98193
R44418 C8_P_btm.n150 C8_P_btm.t104 3.98193
R44419 C8_P_btm.n360 C8_P_btm.t244 3.98193
R44420 C8_P_btm.n362 C8_P_btm.t150 3.98193
R44421 C8_P_btm.n367 C8_P_btm.t177 3.98193
R44422 C8_P_btm.n755 C8_P_btm.t203 3.98193
R44423 C8_P_btm.n758 C8_P_btm.t122 3.98193
R44424 C8_P_btm.n763 C8_P_btm.t133 3.98193
R44425 C8_P_btm.n786 C8_P_btm.t108 3.98193
R44426 C8_P_btm.n789 C8_P_btm.t71 3.98193
R44427 C8_P_btm.n794 C8_P_btm.t263 3.98193
R44428 C8_P_btm.n817 C8_P_btm.t132 3.98193
R44429 C8_P_btm.n820 C8_P_btm.t32 3.98193
R44430 C8_P_btm.n825 C8_P_btm.t205 3.98193
R44431 C8_P_btm.n859 C8_P_btm.t228 3.98193
R44432 C8_P_btm.n862 C8_P_btm.t95 3.98193
R44433 C8_P_btm.n867 C8_P_btm.t159 3.98193
R44434 C8_P_btm.n888 C8_P_btm.t183 3.98193
R44435 C8_P_btm.n0 C8_P_btm.t3 3.57113
R44436 C8_P_btm.n0 C8_P_btm.t1 3.57113
R44437 C8_P_btm.n1 C8_P_btm.t2 3.57113
R44438 C8_P_btm.n1 C8_P_btm.t0 3.57113
R44439 C8_P_btm.n3 C8_P_btm.t274 2.4755
R44440 C8_P_btm.n3 C8_P_btm.t275 2.4755
R44441 C8_P_btm.n5 C8_P_btm.t5 2.4755
R44442 C8_P_btm.n5 C8_P_btm.t4 2.4755
R44443 C8_P_btm.n899 C8_P_btm.t138 1.67819
R44444 C8_P_btm.n896 C8_P_btm.t225 1.67819
R44445 C8_P_btm.n893 C8_P_btm.t149 1.67819
R44446 C8_P_btm.n886 C8_P_btm.t245 1.67819
R44447 C8_P_btm.n883 C8_P_btm.t123 1.67819
R44448 C8_P_btm.n880 C8_P_btm.t231 1.67819
R44449 C8_P_btm.n874 C8_P_btm.t207 1.67819
R44450 C8_P_btm.n872 C8_P_btm.t28 1.67819
R44451 C8_P_btm.n869 C8_P_btm.t220 1.67819
R44452 C8_P_btm.n863 C8_P_btm.t101 1.67819
R44453 C8_P_btm.n841 C8_P_btm.t188 1.67819
R44454 C8_P_btm.n844 C8_P_btm.t267 1.67819
R44455 C8_P_btm.n851 C8_P_btm.t19 1.67819
R44456 C8_P_btm.n854 C8_P_btm.t259 1.67819
R44457 C8_P_btm.n857 C8_P_btm.t131 1.67819
R44458 C8_P_btm.n827 C8_P_btm.t39 1.67819
R44459 C8_P_btm.n830 C8_P_btm.t67 1.67819
R44460 C8_P_btm.n833 C8_P_btm.t249 1.67819
R44461 C8_P_btm.n37 C8_P_btm.t74 1.67819
R44462 C8_P_btm.n35 C8_P_btm.t154 1.67819
R44463 C8_P_btm.n821 C8_P_btm.t86 1.67819
R44464 C8_P_btm.n815 C8_P_btm.t61 1.67819
R44465 C8_P_btm.n812 C8_P_btm.t270 1.67819
R44466 C8_P_btm.n809 C8_P_btm.t117 1.67819
R44467 C8_P_btm.n802 C8_P_btm.t135 1.67819
R44468 C8_P_btm.n799 C8_P_btm.t224 1.67819
R44469 C8_P_btm.n796 C8_P_btm.t148 1.67819
R44470 C8_P_btm.n790 C8_P_btm.t125 1.67819
R44471 C8_P_btm.n52 C8_P_btm.t200 1.67819
R44472 C8_P_btm.n54 C8_P_btm.t175 1.67819
R44473 C8_P_btm.n778 C8_P_btm.t92 1.67819
R44474 C8_P_btm.n781 C8_P_btm.t174 1.67819
R44475 C8_P_btm.n784 C8_P_btm.t103 1.67819
R44476 C8_P_btm.n765 C8_P_btm.t193 1.67819
R44477 C8_P_btm.n768 C8_P_btm.t45 1.67819
R44478 C8_P_btm.n771 C8_P_btm.t179 1.67819
R44479 C8_P_btm.n78 C8_P_btm.t214 1.67819
R44480 C8_P_btm.n75 C8_P_btm.t153 1.67819
R44481 C8_P_btm.n72 C8_P_btm.t242 1.67819
R44482 C8_P_btm.n759 C8_P_btm.t166 1.67819
R44483 C8_P_btm.n753 C8_P_btm.t256 1.67819
R44484 C8_P_btm.n750 C8_P_btm.t64 1.67819
R44485 C8_P_btm.n747 C8_P_btm.t251 1.67819
R44486 C8_P_btm.n744 C8_P_btm.t42 1.67819
R44487 C8_P_btm.n741 C8_P_btm.t236 1.67819
R44488 C8_P_btm.n738 C8_P_btm.t29 1.67819
R44489 C8_P_btm.n81 C8_P_btm.t142 1.67819
R44490 C8_P_btm.n735 C8_P_btm.t82 1.67819
R44491 C8_P_btm.n732 C8_P_btm.t271 1.67819
R44492 C8_P_btm.n729 C8_P_btm.t69 1.67819
R44493 C8_P_btm.n726 C8_P_btm.t124 1.67819
R44494 C8_P_btm.n723 C8_P_btm.t53 1.67819
R44495 C8_P_btm.n720 C8_P_btm.t128 1.67819
R44496 C8_P_btm.n717 C8_P_btm.t33 1.67819
R44497 C8_P_btm.n714 C8_P_btm.t87 1.67819
R44498 C8_P_btm.n711 C8_P_btm.t155 1.67819
R44499 C8_P_btm.n708 C8_P_btm.t75 1.67819
R44500 C8_P_btm.n705 C8_P_btm.t265 1.67819
R44501 C8_P_btm.n702 C8_P_btm.t185 1.67819
R44502 C8_P_btm.n699 C8_P_btm.t221 1.67819
R44503 C8_P_btm.n696 C8_P_btm.t172 1.67819
R44504 C8_P_btm.n693 C8_P_btm.t90 1.67819
R44505 C8_P_btm.n690 C8_P_btm.t157 1.67819
R44506 C8_P_btm.n687 C8_P_btm.t219 1.67819
R44507 C8_P_btm.n684 C8_P_btm.t143 1.67819
R44508 C8_P_btm.n681 C8_P_btm.t215 1.67819
R44509 C8_P_btm.n678 C8_P_btm.t21 1.67819
R44510 C8_P_btm.n675 C8_P_btm.t186 1.67819
R44511 C8_P_btm.n672 C8_P_btm.t250 1.67819
R44512 C8_P_btm.n665 C8_P_btm.t152 1.67819
R44513 C8_P_btm.n662 C8_P_btm.t98 1.67819
R44514 C8_P_btm.n659 C8_P_btm.t180 1.67819
R44515 C8_P_btm.n656 C8_P_btm.t258 1.67819
R44516 C8_P_btm.n645 C8_P_btm.t208 1.67819
R44517 C8_P_btm.n642 C8_P_btm.t120 1.67819
R44518 C8_P_btm.n639 C8_P_btm.t178 1.67819
R44519 C8_P_btm.n633 C8_P_btm.t91 1.67819
R44520 C8_P_btm.n631 C8_P_btm.t268 1.67819
R44521 C8_P_btm.n628 C8_P_btm.t233 1.67819
R44522 C8_P_btm.n622 C8_P_btm.t140 1.67819
R44523 C8_P_btm.n600 C8_P_btm.t57 1.67819
R44524 C8_P_btm.n603 C8_P_btm.t168 1.67819
R44525 C8_P_btm.n610 C8_P_btm.t134 1.67819
R44526 C8_P_btm.n613 C8_P_btm.t79 1.67819
R44527 C8_P_btm.n616 C8_P_btm.t162 1.67819
R44528 C8_P_btm.n586 C8_P_btm.t76 1.67819
R44529 C8_P_btm.n589 C8_P_btm.t24 1.67819
R44530 C8_P_btm.n592 C8_P_btm.t114 1.67819
R44531 C8_P_btm.n482 C8_P_btm.t73 1.67819
R44532 C8_P_btm.n480 C8_P_btm.t51 1.67819
R44533 C8_P_btm.n580 C8_P_btm.t100 1.67819
R44534 C8_P_btm.n574 C8_P_btm.t22 1.67819
R44535 C8_P_btm.n571 C8_P_btm.t187 1.67819
R44536 C8_P_btm.n568 C8_P_btm.t248 1.67819
R44537 C8_P_btm.n561 C8_P_btm.t18 1.67819
R44538 C8_P_btm.n558 C8_P_btm.t213 1.67819
R44539 C8_P_btm.n555 C8_P_btm.t35 1.67819
R44540 C8_P_btm.n549 C8_P_btm.t58 1.67819
R44541 C8_P_btm.n497 C8_P_btm.t238 1.67819
R44542 C8_P_btm.n499 C8_P_btm.t34 1.67819
R44543 C8_P_btm.n537 C8_P_btm.t206 1.67819
R44544 C8_P_btm.n540 C8_P_btm.t144 1.67819
R44545 C8_P_btm.n543 C8_P_btm.t235 1.67819
R44546 C8_P_btm.n524 C8_P_btm.t96 1.67819
R44547 C8_P_btm.n527 C8_P_btm.t169 1.67819
R44548 C8_P_btm.n530 C8_P_btm.t229 1.67819
R44549 C8_P_btm.n510 C8_P_btm.t136 1.67819
R44550 C8_P_btm.n513 C8_P_btm.t81 1.67819
R44551 C8_P_btm.n518 C8_P_btm.t163 1.67819
R44552 C8_P_btm.n653 C8_P_btm.t253 1.67819
R44553 C8_P_btm.n450 C8_P_btm.t222 1.67819
R44554 C8_P_btm.n447 C8_P_btm.t161 1.67819
R44555 C8_P_btm.n444 C8_P_btm.t48 1.67819
R44556 C8_P_btm.n441 C8_P_btm.t189 1.67819
R44557 C8_P_btm.n438 C8_P_btm.t252 1.67819
R44558 C8_P_btm.n435 C8_P_btm.t194 1.67819
R44559 C8_P_btm.n432 C8_P_btm.t273 1.67819
R44560 C8_P_btm.n429 C8_P_btm.t66 1.67819
R44561 C8_P_btm.n426 C8_P_btm.t147 1.67819
R44562 C8_P_btm.n423 C8_P_btm.t94 1.67819
R44563 C8_P_btm.n420 C8_P_btm.t160 1.67819
R44564 C8_P_btm.n417 C8_P_btm.t107 1.67819
R44565 C8_P_btm.n414 C8_P_btm.t130 1.67819
R44566 C8_P_btm.n411 C8_P_btm.t272 1.67819
R44567 C8_P_btm.n408 C8_P_btm.t62 1.67819
R44568 C8_P_btm.n405 C8_P_btm.t255 1.67819
R44569 C8_P_btm.n402 C8_P_btm.t89 1.67819
R44570 C8_P_btm.n399 C8_P_btm.t118 1.67819
R44571 C8_P_btm.n396 C8_P_btm.t269 1.67819
R44572 C8_P_btm.n393 C8_P_btm.t105 1.67819
R44573 C8_P_btm.n390 C8_P_btm.t240 1.67819
R44574 C8_P_btm.n387 C8_P_btm.t59 1.67819
R44575 C8_P_btm.n384 C8_P_btm.t55 1.67819
R44576 C8_P_btm.n381 C8_P_btm.t210 1.67819
R44577 C8_P_btm.n378 C8_P_btm.t54 1.67819
R44578 C8_P_btm.n375 C8_P_btm.t223 1.67819
R44579 C8_P_btm.n372 C8_P_btm.t52 1.67819
R44580 C8_P_btm.n369 C8_P_btm.t237 1.67819
R44581 C8_P_btm.n363 C8_P_btm.t212 1.67819
R44582 C8_P_btm.n194 C8_P_btm.t109 1.67819
R44583 C8_P_btm.n197 C8_P_btm.t199 1.67819
R44584 C8_P_btm.n200 C8_P_btm.t47 1.67819
R44585 C8_P_btm.n203 C8_P_btm.t182 1.67819
R44586 C8_P_btm.n206 C8_P_btm.t243 1.67819
R44587 C8_P_btm.n209 C8_P_btm.t36 1.67819
R44588 C8_P_btm.n212 C8_P_btm.t216 1.67819
R44589 C8_P_btm.n215 C8_P_btm.t192 1.67819
R44590 C8_P_btm.n218 C8_P_btm.t78 1.67819
R44591 C8_P_btm.n221 C8_P_btm.t20 1.67819
R44592 C8_P_btm.n224 C8_P_btm.t65 1.67819
R44593 C8_P_btm.n227 C8_P_btm.t247 1.67819
R44594 C8_P_btm.n230 C8_P_btm.t43 1.67819
R44595 C8_P_btm.n233 C8_P_btm.t116 1.67819
R44596 C8_P_btm.n236 C8_P_btm.t30 1.67819
R44597 C8_P_btm.n239 C8_P_btm.t83 1.67819
R44598 C8_P_btm.n242 C8_P_btm.t137 1.67819
R44599 C8_P_btm.n245 C8_P_btm.t70 1.67819
R44600 C8_P_btm.n248 C8_P_btm.t260 1.67819
R44601 C8_P_btm.n251 C8_P_btm.t56 1.67819
R44602 C8_P_btm.n254 C8_P_btm.t129 1.67819
R44603 C8_P_btm.n257 C8_P_btm.t167 1.67819
R44604 C8_P_btm.n260 C8_P_btm.t97 1.67819
R44605 C8_P_btm.n263 C8_P_btm.t164 1.67819
R44606 C8_P_btm.n266 C8_P_btm.t226 1.67819
R44607 C8_P_btm.n269 C8_P_btm.t139 1.67819
R44608 C8_P_btm.n271 C8_P_btm.t197 1.67819
R44609 C8_P_btm.n277 C8_P_btm.t26 1.67819
R44610 C8_P_btm.n280 C8_P_btm.t232 1.67819
R44611 C8_P_btm.n283 C8_P_btm.t176 1.67819
R44612 C8_P_btm.n286 C8_P_btm.t111 1.67819
R44613 C8_P_btm.n289 C8_P_btm.t184 1.67819
R44614 C8_P_btm.n292 C8_P_btm.t23 1.67819
R44615 C8_P_btm.n295 C8_P_btm.t204 1.67819
R44616 C8_P_btm.n298 C8_P_btm.t266 1.67819
R44617 C8_P_btm.n301 C8_P_btm.t217 1.67819
R44618 C8_P_btm.n304 C8_P_btm.t156 1.67819
R44619 C8_P_btm.n307 C8_P_btm.t230 1.67819
R44620 C8_P_btm.n310 C8_P_btm.t171 1.67819
R44621 C8_P_btm.n313 C8_P_btm.t190 1.67819
R44622 C8_P_btm.n316 C8_P_btm.t201 1.67819
R44623 C8_P_btm.n319 C8_P_btm.t262 1.67819
R44624 C8_P_btm.n322 C8_P_btm.t72 1.67819
R44625 C8_P_btm.n325 C8_P_btm.t151 1.67819
R44626 C8_P_btm.n328 C8_P_btm.t85 1.67819
R44627 C8_P_btm.n331 C8_P_btm.t165 1.67819
R44628 C8_P_btm.n334 C8_P_btm.t119 1.67819
R44629 C8_P_btm.n337 C8_P_btm.t49 1.67819
R44630 C8_P_btm.n340 C8_P_btm.t121 1.67819
R44631 C8_P_btm.n343 C8_P_btm.t68 1.67819
R44632 C8_P_btm.n346 C8_P_btm.t25 1.67819
R44633 C8_P_btm.n349 C8_P_btm.t80 1.67819
R44634 C8_P_btm.n352 C8_P_btm.t27 1.67819
R44635 C8_P_btm.n355 C8_P_btm.t113 1.67819
R44636 C8_P_btm.n358 C8_P_btm.t40 1.67819
R44637 C8_P_btm.n84 C8_P_btm.n83 1.05569
R44638 C8_P_btm.n651 C8_P_btm.n101 1.05569
R44639 C8_P_btm.n152 C8_P_btm.n151 1.05569
R44640 C8_P_btm.n150 C8_P_btm.n149 1.05569
R44641 C8_P_btm.n361 C8_P_btm.n360 1.05569
R44642 C8_P_btm.n275 C8_P_btm.n107 1.05569
R44643 C8_P_btm.n14 C8_P_btm.n12 1.0005
R44644 C8_P_btm.n15 C8_P_btm.n11 1.0005
R44645 C8_P_btm.n877 C8_P_btm.n10 1.0005
R44646 C8_P_btm.n877 C8_P_btm.n876 1.0005
R44647 C8_P_btm.n18 C8_P_btm.n15 1.0005
R44648 C8_P_btm.n866 C8_P_btm.n14 1.0005
R44649 C8_P_btm.n866 C8_P_btm.n865 1.0005
R44650 C8_P_btm.n839 C8_P_btm.n18 1.0005
R44651 C8_P_btm.n876 C8_P_btm.n16 1.0005
R44652 C8_P_btm.n23 C8_P_btm.n16 1.0005
R44653 C8_P_btm.n839 C8_P_btm.n22 1.0005
R44654 C8_P_btm.n865 C8_P_btm.n19 1.0005
R44655 C8_P_btm.n824 C8_P_btm.n19 1.0005
R44656 C8_P_btm.n26 C8_P_btm.n22 1.0005
R44657 C8_P_btm.n25 C8_P_btm.n23 1.0005
R44658 C8_P_btm.n39 C8_P_btm.n25 1.0005
R44659 C8_P_btm.n33 C8_P_btm.n26 1.0005
R44660 C8_P_btm.n824 C8_P_btm.n823 1.0005
R44661 C8_P_btm.n823 C8_P_btm.n27 1.0005
R44662 C8_P_btm.n33 C8_P_btm.n30 1.0005
R44663 C8_P_btm.n40 C8_P_btm.n39 1.0005
R44664 C8_P_btm.n42 C8_P_btm.n40 1.0005
R44665 C8_P_btm.n43 C8_P_btm.n30 1.0005
R44666 C8_P_btm.n793 C8_P_btm.n27 1.0005
R44667 C8_P_btm.n793 C8_P_btm.n792 1.0005
R44668 C8_P_btm.n50 C8_P_btm.n43 1.0005
R44669 C8_P_btm.n56 C8_P_btm.n42 1.0005
R44670 C8_P_btm.n57 C8_P_btm.n56 1.0005
R44671 C8_P_btm.n50 C8_P_btm.n47 1.0005
R44672 C8_P_btm.n792 C8_P_btm.n44 1.0005
R44673 C8_P_btm.n762 C8_P_btm.n44 1.0005
R44674 C8_P_btm.n60 C8_P_btm.n47 1.0005
R44675 C8_P_btm.n59 C8_P_btm.n57 1.0005
R44676 C8_P_btm.n69 C8_P_btm.n59 1.0005
R44677 C8_P_btm.n70 C8_P_btm.n60 1.0005
R44678 C8_P_btm.n762 C8_P_btm.n761 1.0005
R44679 C8_P_btm.n761 C8_P_btm.n61 1.0005
R44680 C8_P_btm.n70 C8_P_btm.n64 1.0005
R44681 C8_P_btm.n69 C8_P_btm.n65 1.0005
R44682 C8_P_btm.n66 C8_P_btm.n58 1.0005
R44683 C8_P_btm.n68 C8_P_btm.n67 1.0005
R44684 C8_P_btm.n455 C8_P_btm.n106 1.0005
R44685 C8_P_btm.n456 C8_P_btm.n105 1.0005
R44686 C8_P_btm.n457 C8_P_btm.n104 1.0005
R44687 C8_P_btm.n459 C8_P_btm.n457 1.0005
R44688 C8_P_btm.n460 C8_P_btm.n456 1.0005
R44689 C8_P_btm.n636 C8_P_btm.n455 1.0005
R44690 C8_P_btm.n636 C8_P_btm.n635 1.0005
R44691 C8_P_btm.n463 C8_P_btm.n460 1.0005
R44692 C8_P_btm.n625 C8_P_btm.n459 1.0005
R44693 C8_P_btm.n625 C8_P_btm.n624 1.0005
R44694 C8_P_btm.n598 C8_P_btm.n463 1.0005
R44695 C8_P_btm.n635 C8_P_btm.n461 1.0005
R44696 C8_P_btm.n468 C8_P_btm.n461 1.0005
R44697 C8_P_btm.n598 C8_P_btm.n467 1.0005
R44698 C8_P_btm.n624 C8_P_btm.n464 1.0005
R44699 C8_P_btm.n583 C8_P_btm.n464 1.0005
R44700 C8_P_btm.n471 C8_P_btm.n467 1.0005
R44701 C8_P_btm.n470 C8_P_btm.n468 1.0005
R44702 C8_P_btm.n484 C8_P_btm.n470 1.0005
R44703 C8_P_btm.n478 C8_P_btm.n471 1.0005
R44704 C8_P_btm.n583 C8_P_btm.n582 1.0005
R44705 C8_P_btm.n582 C8_P_btm.n472 1.0005
R44706 C8_P_btm.n478 C8_P_btm.n475 1.0005
R44707 C8_P_btm.n485 C8_P_btm.n484 1.0005
R44708 C8_P_btm.n487 C8_P_btm.n485 1.0005
R44709 C8_P_btm.n488 C8_P_btm.n475 1.0005
R44710 C8_P_btm.n552 C8_P_btm.n472 1.0005
R44711 C8_P_btm.n552 C8_P_btm.n551 1.0005
R44712 C8_P_btm.n495 C8_P_btm.n488 1.0005
R44713 C8_P_btm.n501 C8_P_btm.n487 1.0005
R44714 C8_P_btm.n502 C8_P_btm.n501 1.0005
R44715 C8_P_btm.n495 C8_P_btm.n492 1.0005
R44716 C8_P_btm.n551 C8_P_btm.n489 1.0005
R44717 C8_P_btm.n521 C8_P_btm.n489 1.0005
R44718 C8_P_btm.n505 C8_P_btm.n492 1.0005
R44719 C8_P_btm.n504 C8_P_btm.n502 1.0005
R44720 C8_P_btm.n507 C8_P_btm.n504 1.0005
R44721 C8_P_btm.n506 C8_P_btm.n505 1.0005
R44722 C8_P_btm.n521 C8_P_btm.n520 1.0005
R44723 C8_P_btm.n516 C8_P_btm.n491 1.0005
R44724 C8_P_btm.n534 C8_P_btm.n533 1.0005
R44725 C8_P_btm.n533 C8_P_btm.n503 1.0005
R44726 C8_P_btm.n547 C8_P_btm.n546 1.0005
R44727 C8_P_btm.n546 C8_P_btm.n491 1.0005
R44728 C8_P_btm.n564 C8_P_btm.n486 1.0005
R44729 C8_P_btm.n534 C8_P_btm.n486 1.0005
R44730 C8_P_btm.n577 C8_P_btm.n474 1.0005
R44731 C8_P_btm.n547 C8_P_btm.n474 1.0005
R44732 C8_P_btm.n565 C8_P_btm.n469 1.0005
R44733 C8_P_btm.n565 C8_P_btm.n564 1.0005
R44734 C8_P_btm.n578 C8_P_btm.n466 1.0005
R44735 C8_P_btm.n578 C8_P_btm.n577 1.0005
R44736 C8_P_btm.n607 C8_P_btm.n595 1.0005
R44737 C8_P_btm.n595 C8_P_btm.n469 1.0005
R44738 C8_P_btm.n620 C8_P_btm.n619 1.0005
R44739 C8_P_btm.n619 C8_P_btm.n466 1.0005
R44740 C8_P_btm.n606 C8_P_btm.n597 1.0005
R44741 C8_P_btm.n607 C8_P_btm.n606 1.0005
R44742 C8_P_btm.n648 C8_P_btm.n458 1.0005
R44743 C8_P_btm.n620 C8_P_btm.n458 1.0005
R44744 C8_P_btm.n668 C8_P_btm.n454 1.0005
R44745 C8_P_btm.n597 C8_P_btm.n454 1.0005
R44746 C8_P_btm.n649 C8_P_btm.n103 1.0005
R44747 C8_P_btm.n649 C8_P_btm.n648 1.0005
R44748 C8_P_btm.n650 C8_P_btm.n102 1.0005
R44749 C8_P_btm.n108 C8_P_btm.n106 1.0005
R44750 C8_P_btm.n109 C8_P_btm.n105 1.0005
R44751 C8_P_btm.n110 C8_P_btm.n104 1.0005
R44752 C8_P_btm.n111 C8_P_btm.n103 1.0005
R44753 C8_P_btm.n112 C8_P_btm.n102 1.0005
R44754 C8_P_btm.n113 C8_P_btm.n101 1.0005
R44755 C8_P_btm.n114 C8_P_btm.n100 1.0005
R44756 C8_P_btm.n115 C8_P_btm.n99 1.0005
R44757 C8_P_btm.n116 C8_P_btm.n98 1.0005
R44758 C8_P_btm.n117 C8_P_btm.n97 1.0005
R44759 C8_P_btm.n118 C8_P_btm.n96 1.0005
R44760 C8_P_btm.n119 C8_P_btm.n95 1.0005
R44761 C8_P_btm.n120 C8_P_btm.n94 1.0005
R44762 C8_P_btm.n121 C8_P_btm.n93 1.0005
R44763 C8_P_btm.n122 C8_P_btm.n92 1.0005
R44764 C8_P_btm.n123 C8_P_btm.n91 1.0005
R44765 C8_P_btm.n124 C8_P_btm.n90 1.0005
R44766 C8_P_btm.n125 C8_P_btm.n89 1.0005
R44767 C8_P_btm.n126 C8_P_btm.n88 1.0005
R44768 C8_P_btm.n127 C8_P_btm.n87 1.0005
R44769 C8_P_btm.n128 C8_P_btm.n86 1.0005
R44770 C8_P_btm.n129 C8_P_btm.n85 1.0005
R44771 C8_P_btm.n130 C8_P_btm.n84 1.0005
R44772 C8_P_btm.n131 C8_P_btm.n67 1.0005
R44773 C8_P_btm.n132 C8_P_btm.n66 1.0005
R44774 C8_P_btm.n133 C8_P_btm.n65 1.0005
R44775 C8_P_btm.n134 C8_P_btm.n64 1.0005
R44776 C8_P_btm.n366 C8_P_btm.n61 1.0005
R44777 C8_P_btm.n366 C8_P_btm.n365 1.0005
R44778 C8_P_btm.n192 C8_P_btm.n134 1.0005
R44779 C8_P_btm.n191 C8_P_btm.n133 1.0005
R44780 C8_P_btm.n190 C8_P_btm.n132 1.0005
R44781 C8_P_btm.n189 C8_P_btm.n131 1.0005
R44782 C8_P_btm.n188 C8_P_btm.n130 1.0005
R44783 C8_P_btm.n187 C8_P_btm.n129 1.0005
R44784 C8_P_btm.n186 C8_P_btm.n128 1.0005
R44785 C8_P_btm.n185 C8_P_btm.n127 1.0005
R44786 C8_P_btm.n184 C8_P_btm.n126 1.0005
R44787 C8_P_btm.n183 C8_P_btm.n125 1.0005
R44788 C8_P_btm.n182 C8_P_btm.n124 1.0005
R44789 C8_P_btm.n181 C8_P_btm.n123 1.0005
R44790 C8_P_btm.n180 C8_P_btm.n122 1.0005
R44791 C8_P_btm.n179 C8_P_btm.n121 1.0005
R44792 C8_P_btm.n178 C8_P_btm.n120 1.0005
R44793 C8_P_btm.n177 C8_P_btm.n119 1.0005
R44794 C8_P_btm.n176 C8_P_btm.n118 1.0005
R44795 C8_P_btm.n175 C8_P_btm.n117 1.0005
R44796 C8_P_btm.n174 C8_P_btm.n116 1.0005
R44797 C8_P_btm.n173 C8_P_btm.n115 1.0005
R44798 C8_P_btm.n172 C8_P_btm.n114 1.0005
R44799 C8_P_btm.n171 C8_P_btm.n113 1.0005
R44800 C8_P_btm.n170 C8_P_btm.n112 1.0005
R44801 C8_P_btm.n169 C8_P_btm.n111 1.0005
R44802 C8_P_btm.n168 C8_P_btm.n110 1.0005
R44803 C8_P_btm.n167 C8_P_btm.n109 1.0005
R44804 C8_P_btm.n273 C8_P_btm.n108 1.0005
R44805 C8_P_btm.n274 C8_P_btm.n273 1.0005
R44806 C8_P_btm.n167 C8_P_btm.n164 1.0005
R44807 C8_P_btm.n168 C8_P_btm.n163 1.0005
R44808 C8_P_btm.n169 C8_P_btm.n162 1.0005
R44809 C8_P_btm.n170 C8_P_btm.n161 1.0005
R44810 C8_P_btm.n171 C8_P_btm.n160 1.0005
R44811 C8_P_btm.n172 C8_P_btm.n159 1.0005
R44812 C8_P_btm.n173 C8_P_btm.n158 1.0005
R44813 C8_P_btm.n174 C8_P_btm.n157 1.0005
R44814 C8_P_btm.n175 C8_P_btm.n156 1.0005
R44815 C8_P_btm.n176 C8_P_btm.n155 1.0005
R44816 C8_P_btm.n177 C8_P_btm.n154 1.0005
R44817 C8_P_btm.n178 C8_P_btm.n153 1.0005
R44818 C8_P_btm.n179 C8_P_btm.n152 1.0005
R44819 C8_P_btm.n180 C8_P_btm.n149 1.0005
R44820 C8_P_btm.n181 C8_P_btm.n148 1.0005
R44821 C8_P_btm.n182 C8_P_btm.n147 1.0005
R44822 C8_P_btm.n183 C8_P_btm.n146 1.0005
R44823 C8_P_btm.n184 C8_P_btm.n145 1.0005
R44824 C8_P_btm.n185 C8_P_btm.n144 1.0005
R44825 C8_P_btm.n186 C8_P_btm.n143 1.0005
R44826 C8_P_btm.n187 C8_P_btm.n142 1.0005
R44827 C8_P_btm.n188 C8_P_btm.n141 1.0005
R44828 C8_P_btm.n189 C8_P_btm.n140 1.0005
R44829 C8_P_btm.n190 C8_P_btm.n139 1.0005
R44830 C8_P_btm.n191 C8_P_btm.n138 1.0005
R44831 C8_P_btm.n192 C8_P_btm.n137 1.0005
R44832 C8_P_btm.n365 C8_P_btm.n135 1.0005
R44833 C8_P_btm.n453 C8_P_btm.n107 1.0005
R44834 C8_P_btm.n361 C8_P_btm.n63 1.0005
R44835 C8_P_btm.n756 C8_P_btm.n63 1.0005
R44836 C8_P_btm.n669 C8_P_btm.n453 1.0005
R44837 C8_P_btm.n669 C8_P_btm.n668 1.0005
R44838 C8_P_btm.n757 C8_P_btm.n756 1.0005
R44839 C8_P_btm.n757 C8_P_btm.n46 1.0005
R44840 C8_P_btm.n774 C8_P_btm.n58 1.0005
R44841 C8_P_btm.n775 C8_P_btm.n774 1.0005
R44842 C8_P_btm.n787 C8_P_btm.n46 1.0005
R44843 C8_P_btm.n788 C8_P_btm.n787 1.0005
R44844 C8_P_btm.n775 C8_P_btm.n41 1.0005
R44845 C8_P_btm.n805 C8_P_btm.n41 1.0005
R44846 C8_P_btm.n788 C8_P_btm.n29 1.0005
R44847 C8_P_btm.n818 C8_P_btm.n29 1.0005
R44848 C8_P_btm.n806 C8_P_btm.n805 1.0005
R44849 C8_P_btm.n806 C8_P_btm.n24 1.0005
R44850 C8_P_btm.n819 C8_P_btm.n818 1.0005
R44851 C8_P_btm.n819 C8_P_btm.n21 1.0005
R44852 C8_P_btm.n836 C8_P_btm.n24 1.0005
R44853 C8_P_btm.n848 C8_P_btm.n836 1.0005
R44854 C8_P_btm.n860 C8_P_btm.n21 1.0005
R44855 C8_P_btm.n861 C8_P_btm.n860 1.0005
R44856 C8_P_btm.n848 C8_P_btm.n847 1.0005
R44857 C8_P_btm.n847 C8_P_btm.n838 1.0005
R44858 C8_P_btm.n861 C8_P_btm.n13 1.0005
R44859 C8_P_btm.n889 C8_P_btm.n13 1.0005
R44860 C8_P_btm.n838 C8_P_btm.n9 1.0005
R44861 C8_P_btm.n902 C8_P_btm.n9 1.0005
R44862 C8_P_btm.n890 C8_P_btm.n889 1.0005
R44863 C8_P_btm.n903 C8_P_btm.n902 1.0005
R44864 C8_P_btm.n151 C8_P_btm.n150 0.733338
R44865 C8_P_btm.n83 C8_P_btm.n82 0.679419
R44866 C8_P_btm.n519 C8_P_btm.n517 0.679419
R44867 C8_P_btm.n509 C8_P_btm.n508 0.679419
R44868 C8_P_btm.n532 C8_P_btm.n531 0.679419
R44869 C8_P_btm.n523 C8_P_btm.n522 0.679419
R44870 C8_P_btm.n545 C8_P_btm.n544 0.679419
R44871 C8_P_btm.n536 C8_P_btm.n535 0.679419
R44872 C8_P_btm.n494 C8_P_btm.n493 0.679419
R44873 C8_P_btm.n550 C8_P_btm.n548 0.679419
R44874 C8_P_btm.n554 C8_P_btm.n553 0.679419
R44875 C8_P_btm.n563 C8_P_btm.n562 0.679419
R44876 C8_P_btm.n567 C8_P_btm.n566 0.679419
R44877 C8_P_btm.n576 C8_P_btm.n575 0.679419
R44878 C8_P_btm.n581 C8_P_btm.n579 0.679419
R44879 C8_P_btm.n477 C8_P_btm.n476 0.679419
R44880 C8_P_btm.n594 C8_P_btm.n593 0.679419
R44881 C8_P_btm.n585 C8_P_btm.n584 0.679419
R44882 C8_P_btm.n618 C8_P_btm.n617 0.679419
R44883 C8_P_btm.n609 C8_P_btm.n608 0.679419
R44884 C8_P_btm.n605 C8_P_btm.n604 0.679419
R44885 C8_P_btm.n623 C8_P_btm.n621 0.679419
R44886 C8_P_btm.n627 C8_P_btm.n626 0.679419
R44887 C8_P_btm.n596 C8_P_btm.n462 0.679419
R44888 C8_P_btm.n638 C8_P_btm.n637 0.679419
R44889 C8_P_btm.n647 C8_P_btm.n646 0.679419
R44890 C8_P_btm.n652 C8_P_btm.n651 0.679419
R44891 C8_P_btm.n667 C8_P_btm.n666 0.679419
R44892 C8_P_btm.n360 C8_P_btm.n359 0.679419
R44893 C8_P_btm.n276 C8_P_btm.n275 0.679419
R44894 C8_P_btm.n166 C8_P_btm.n165 0.679419
R44895 C8_P_btm.n364 C8_P_btm.n362 0.679419
R44896 C8_P_btm.n368 C8_P_btm.n367 0.679419
R44897 C8_P_btm.n452 C8_P_btm.n451 0.679419
R44898 C8_P_btm.n671 C8_P_btm.n670 0.679419
R44899 C8_P_btm.n755 C8_P_btm.n754 0.679419
R44900 C8_P_btm.n760 C8_P_btm.n758 0.679419
R44901 C8_P_btm.n773 C8_P_btm.n772 0.679419
R44902 C8_P_btm.n764 C8_P_btm.n763 0.679419
R44903 C8_P_btm.n786 C8_P_btm.n785 0.679419
R44904 C8_P_btm.n777 C8_P_btm.n776 0.679419
R44905 C8_P_btm.n49 C8_P_btm.n48 0.679419
R44906 C8_P_btm.n791 C8_P_btm.n789 0.679419
R44907 C8_P_btm.n795 C8_P_btm.n794 0.679419
R44908 C8_P_btm.n804 C8_P_btm.n803 0.679419
R44909 C8_P_btm.n808 C8_P_btm.n807 0.679419
R44910 C8_P_btm.n817 C8_P_btm.n816 0.679419
R44911 C8_P_btm.n822 C8_P_btm.n820 0.679419
R44912 C8_P_btm.n32 C8_P_btm.n31 0.679419
R44913 C8_P_btm.n835 C8_P_btm.n834 0.679419
R44914 C8_P_btm.n826 C8_P_btm.n825 0.679419
R44915 C8_P_btm.n859 C8_P_btm.n858 0.679419
R44916 C8_P_btm.n850 C8_P_btm.n849 0.679419
R44917 C8_P_btm.n846 C8_P_btm.n845 0.679419
R44918 C8_P_btm.n864 C8_P_btm.n862 0.679419
R44919 C8_P_btm.n868 C8_P_btm.n867 0.679419
R44920 C8_P_btm.n837 C8_P_btm.n17 0.679419
R44921 C8_P_btm.n879 C8_P_btm.n878 0.679419
R44922 C8_P_btm.n888 C8_P_btm.n887 0.679419
R44923 C8_P_btm.n892 C8_P_btm.n891 0.679419
R44924 C8_P_btm.n901 C8_P_btm.n900 0.679419
R44925 C8_P_btm.n80 C8_P_btm.n79 0.6255
R44926 C8_P_btm.n515 C8_P_btm.n514 0.6255
R44927 C8_P_btm.n512 C8_P_btm.n511 0.6255
R44928 C8_P_btm.n529 C8_P_btm.n528 0.6255
R44929 C8_P_btm.n526 C8_P_btm.n525 0.6255
R44930 C8_P_btm.n542 C8_P_btm.n541 0.6255
R44931 C8_P_btm.n539 C8_P_btm.n538 0.6255
R44932 C8_P_btm.n500 C8_P_btm.n498 0.6255
R44933 C8_P_btm.n496 C8_P_btm.n490 0.6255
R44934 C8_P_btm.n557 C8_P_btm.n556 0.6255
R44935 C8_P_btm.n560 C8_P_btm.n559 0.6255
R44936 C8_P_btm.n570 C8_P_btm.n569 0.6255
R44937 C8_P_btm.n573 C8_P_btm.n572 0.6255
R44938 C8_P_btm.n479 C8_P_btm.n473 0.6255
R44939 C8_P_btm.n483 C8_P_btm.n481 0.6255
R44940 C8_P_btm.n591 C8_P_btm.n590 0.6255
R44941 C8_P_btm.n588 C8_P_btm.n587 0.6255
R44942 C8_P_btm.n615 C8_P_btm.n614 0.6255
R44943 C8_P_btm.n612 C8_P_btm.n611 0.6255
R44944 C8_P_btm.n602 C8_P_btm.n601 0.6255
R44945 C8_P_btm.n599 C8_P_btm.n465 0.6255
R44946 C8_P_btm.n630 C8_P_btm.n629 0.6255
R44947 C8_P_btm.n634 C8_P_btm.n632 0.6255
R44948 C8_P_btm.n641 C8_P_btm.n640 0.6255
R44949 C8_P_btm.n644 C8_P_btm.n643 0.6255
R44950 C8_P_btm.n655 C8_P_btm.n654 0.6255
R44951 C8_P_btm.n658 C8_P_btm.n657 0.6255
R44952 C8_P_btm.n661 C8_P_btm.n660 0.6255
R44953 C8_P_btm.n664 C8_P_btm.n663 0.6255
R44954 C8_P_btm.n357 C8_P_btm.n356 0.6255
R44955 C8_P_btm.n354 C8_P_btm.n353 0.6255
R44956 C8_P_btm.n351 C8_P_btm.n350 0.6255
R44957 C8_P_btm.n348 C8_P_btm.n347 0.6255
R44958 C8_P_btm.n345 C8_P_btm.n344 0.6255
R44959 C8_P_btm.n342 C8_P_btm.n341 0.6255
R44960 C8_P_btm.n339 C8_P_btm.n338 0.6255
R44961 C8_P_btm.n336 C8_P_btm.n335 0.6255
R44962 C8_P_btm.n333 C8_P_btm.n332 0.6255
R44963 C8_P_btm.n330 C8_P_btm.n329 0.6255
R44964 C8_P_btm.n327 C8_P_btm.n326 0.6255
R44965 C8_P_btm.n324 C8_P_btm.n323 0.6255
R44966 C8_P_btm.n321 C8_P_btm.n320 0.6255
R44967 C8_P_btm.n318 C8_P_btm.n317 0.6255
R44968 C8_P_btm.n315 C8_P_btm.n314 0.6255
R44969 C8_P_btm.n312 C8_P_btm.n311 0.6255
R44970 C8_P_btm.n309 C8_P_btm.n308 0.6255
R44971 C8_P_btm.n306 C8_P_btm.n305 0.6255
R44972 C8_P_btm.n303 C8_P_btm.n302 0.6255
R44973 C8_P_btm.n300 C8_P_btm.n299 0.6255
R44974 C8_P_btm.n297 C8_P_btm.n296 0.6255
R44975 C8_P_btm.n294 C8_P_btm.n293 0.6255
R44976 C8_P_btm.n291 C8_P_btm.n290 0.6255
R44977 C8_P_btm.n288 C8_P_btm.n287 0.6255
R44978 C8_P_btm.n285 C8_P_btm.n284 0.6255
R44979 C8_P_btm.n282 C8_P_btm.n281 0.6255
R44980 C8_P_btm.n279 C8_P_btm.n278 0.6255
R44981 C8_P_btm.n272 C8_P_btm.n270 0.6255
R44982 C8_P_btm.n268 C8_P_btm.n267 0.6255
R44983 C8_P_btm.n265 C8_P_btm.n264 0.6255
R44984 C8_P_btm.n262 C8_P_btm.n261 0.6255
R44985 C8_P_btm.n259 C8_P_btm.n258 0.6255
R44986 C8_P_btm.n256 C8_P_btm.n255 0.6255
R44987 C8_P_btm.n253 C8_P_btm.n252 0.6255
R44988 C8_P_btm.n250 C8_P_btm.n249 0.6255
R44989 C8_P_btm.n247 C8_P_btm.n246 0.6255
R44990 C8_P_btm.n244 C8_P_btm.n243 0.6255
R44991 C8_P_btm.n241 C8_P_btm.n240 0.6255
R44992 C8_P_btm.n238 C8_P_btm.n237 0.6255
R44993 C8_P_btm.n235 C8_P_btm.n234 0.6255
R44994 C8_P_btm.n232 C8_P_btm.n231 0.6255
R44995 C8_P_btm.n229 C8_P_btm.n228 0.6255
R44996 C8_P_btm.n226 C8_P_btm.n225 0.6255
R44997 C8_P_btm.n223 C8_P_btm.n222 0.6255
R44998 C8_P_btm.n220 C8_P_btm.n219 0.6255
R44999 C8_P_btm.n217 C8_P_btm.n216 0.6255
R45000 C8_P_btm.n214 C8_P_btm.n213 0.6255
R45001 C8_P_btm.n211 C8_P_btm.n210 0.6255
R45002 C8_P_btm.n208 C8_P_btm.n207 0.6255
R45003 C8_P_btm.n205 C8_P_btm.n204 0.6255
R45004 C8_P_btm.n202 C8_P_btm.n201 0.6255
R45005 C8_P_btm.n199 C8_P_btm.n198 0.6255
R45006 C8_P_btm.n196 C8_P_btm.n195 0.6255
R45007 C8_P_btm.n193 C8_P_btm.n136 0.6255
R45008 C8_P_btm.n371 C8_P_btm.n370 0.6255
R45009 C8_P_btm.n374 C8_P_btm.n373 0.6255
R45010 C8_P_btm.n377 C8_P_btm.n376 0.6255
R45011 C8_P_btm.n380 C8_P_btm.n379 0.6255
R45012 C8_P_btm.n383 C8_P_btm.n382 0.6255
R45013 C8_P_btm.n386 C8_P_btm.n385 0.6255
R45014 C8_P_btm.n389 C8_P_btm.n388 0.6255
R45015 C8_P_btm.n392 C8_P_btm.n391 0.6255
R45016 C8_P_btm.n395 C8_P_btm.n394 0.6255
R45017 C8_P_btm.n398 C8_P_btm.n397 0.6255
R45018 C8_P_btm.n401 C8_P_btm.n400 0.6255
R45019 C8_P_btm.n404 C8_P_btm.n403 0.6255
R45020 C8_P_btm.n407 C8_P_btm.n406 0.6255
R45021 C8_P_btm.n410 C8_P_btm.n409 0.6255
R45022 C8_P_btm.n413 C8_P_btm.n412 0.6255
R45023 C8_P_btm.n416 C8_P_btm.n415 0.6255
R45024 C8_P_btm.n419 C8_P_btm.n418 0.6255
R45025 C8_P_btm.n422 C8_P_btm.n421 0.6255
R45026 C8_P_btm.n425 C8_P_btm.n424 0.6255
R45027 C8_P_btm.n428 C8_P_btm.n427 0.6255
R45028 C8_P_btm.n431 C8_P_btm.n430 0.6255
R45029 C8_P_btm.n434 C8_P_btm.n433 0.6255
R45030 C8_P_btm.n437 C8_P_btm.n436 0.6255
R45031 C8_P_btm.n440 C8_P_btm.n439 0.6255
R45032 C8_P_btm.n443 C8_P_btm.n442 0.6255
R45033 C8_P_btm.n446 C8_P_btm.n445 0.6255
R45034 C8_P_btm.n449 C8_P_btm.n448 0.6255
R45035 C8_P_btm.n674 C8_P_btm.n673 0.6255
R45036 C8_P_btm.n677 C8_P_btm.n676 0.6255
R45037 C8_P_btm.n680 C8_P_btm.n679 0.6255
R45038 C8_P_btm.n683 C8_P_btm.n682 0.6255
R45039 C8_P_btm.n686 C8_P_btm.n685 0.6255
R45040 C8_P_btm.n689 C8_P_btm.n688 0.6255
R45041 C8_P_btm.n692 C8_P_btm.n691 0.6255
R45042 C8_P_btm.n695 C8_P_btm.n694 0.6255
R45043 C8_P_btm.n698 C8_P_btm.n697 0.6255
R45044 C8_P_btm.n701 C8_P_btm.n700 0.6255
R45045 C8_P_btm.n704 C8_P_btm.n703 0.6255
R45046 C8_P_btm.n707 C8_P_btm.n706 0.6255
R45047 C8_P_btm.n710 C8_P_btm.n709 0.6255
R45048 C8_P_btm.n713 C8_P_btm.n712 0.6255
R45049 C8_P_btm.n716 C8_P_btm.n715 0.6255
R45050 C8_P_btm.n719 C8_P_btm.n718 0.6255
R45051 C8_P_btm.n722 C8_P_btm.n721 0.6255
R45052 C8_P_btm.n725 C8_P_btm.n724 0.6255
R45053 C8_P_btm.n728 C8_P_btm.n727 0.6255
R45054 C8_P_btm.n731 C8_P_btm.n730 0.6255
R45055 C8_P_btm.n734 C8_P_btm.n733 0.6255
R45056 C8_P_btm.n737 C8_P_btm.n736 0.6255
R45057 C8_P_btm.n740 C8_P_btm.n739 0.6255
R45058 C8_P_btm.n743 C8_P_btm.n742 0.6255
R45059 C8_P_btm.n746 C8_P_btm.n745 0.6255
R45060 C8_P_btm.n749 C8_P_btm.n748 0.6255
R45061 C8_P_btm.n752 C8_P_btm.n751 0.6255
R45062 C8_P_btm.n71 C8_P_btm.n62 0.6255
R45063 C8_P_btm.n74 C8_P_btm.n73 0.6255
R45064 C8_P_btm.n77 C8_P_btm.n76 0.6255
R45065 C8_P_btm.n770 C8_P_btm.n769 0.6255
R45066 C8_P_btm.n767 C8_P_btm.n766 0.6255
R45067 C8_P_btm.n783 C8_P_btm.n782 0.6255
R45068 C8_P_btm.n780 C8_P_btm.n779 0.6255
R45069 C8_P_btm.n55 C8_P_btm.n53 0.6255
R45070 C8_P_btm.n51 C8_P_btm.n45 0.6255
R45071 C8_P_btm.n798 C8_P_btm.n797 0.6255
R45072 C8_P_btm.n801 C8_P_btm.n800 0.6255
R45073 C8_P_btm.n811 C8_P_btm.n810 0.6255
R45074 C8_P_btm.n814 C8_P_btm.n813 0.6255
R45075 C8_P_btm.n34 C8_P_btm.n28 0.6255
R45076 C8_P_btm.n38 C8_P_btm.n36 0.6255
R45077 C8_P_btm.n832 C8_P_btm.n831 0.6255
R45078 C8_P_btm.n829 C8_P_btm.n828 0.6255
R45079 C8_P_btm.n856 C8_P_btm.n855 0.6255
R45080 C8_P_btm.n853 C8_P_btm.n852 0.6255
R45081 C8_P_btm.n843 C8_P_btm.n842 0.6255
R45082 C8_P_btm.n840 C8_P_btm.n20 0.6255
R45083 C8_P_btm.n871 C8_P_btm.n870 0.6255
R45084 C8_P_btm.n875 C8_P_btm.n873 0.6255
R45085 C8_P_btm.n882 C8_P_btm.n881 0.6255
R45086 C8_P_btm.n885 C8_P_btm.n884 0.6255
R45087 C8_P_btm.n895 C8_P_btm.n894 0.6255
R45088 C8_P_btm.n898 C8_P_btm.n897 0.6255
R45089 C8_P_btm.n82 C8_P_btm.n68 0.109875
R45090 C8_P_btm.n80 C8_P_btm.n68 0.109875
R45091 C8_P_btm.n520 C8_P_btm.n515 0.109875
R45092 C8_P_btm.n520 C8_P_btm.n519 0.109875
R45093 C8_P_btm.n512 C8_P_btm.n506 0.109875
R45094 C8_P_btm.n514 C8_P_btm.n506 0.109875
R45095 C8_P_btm.n509 C8_P_btm.n507 0.109875
R45096 C8_P_btm.n511 C8_P_btm.n507 0.109875
R45097 C8_P_btm.n531 C8_P_btm.n504 0.109875
R45098 C8_P_btm.n529 C8_P_btm.n504 0.109875
R45099 C8_P_btm.n528 C8_P_btm.n505 0.109875
R45100 C8_P_btm.n526 C8_P_btm.n505 0.109875
R45101 C8_P_btm.n525 C8_P_btm.n521 0.109875
R45102 C8_P_btm.n523 C8_P_btm.n521 0.109875
R45103 C8_P_btm.n542 C8_P_btm.n489 0.109875
R45104 C8_P_btm.n544 C8_P_btm.n489 0.109875
R45105 C8_P_btm.n539 C8_P_btm.n492 0.109875
R45106 C8_P_btm.n541 C8_P_btm.n492 0.109875
R45107 C8_P_btm.n536 C8_P_btm.n502 0.109875
R45108 C8_P_btm.n538 C8_P_btm.n502 0.109875
R45109 C8_P_btm.n501 C8_P_btm.n494 0.109875
R45110 C8_P_btm.n501 C8_P_btm.n500 0.109875
R45111 C8_P_btm.n498 C8_P_btm.n495 0.109875
R45112 C8_P_btm.n496 C8_P_btm.n495 0.109875
R45113 C8_P_btm.n551 C8_P_btm.n490 0.109875
R45114 C8_P_btm.n551 C8_P_btm.n550 0.109875
R45115 C8_P_btm.n556 C8_P_btm.n552 0.109875
R45116 C8_P_btm.n554 C8_P_btm.n552 0.109875
R45117 C8_P_btm.n559 C8_P_btm.n488 0.109875
R45118 C8_P_btm.n557 C8_P_btm.n488 0.109875
R45119 C8_P_btm.n562 C8_P_btm.n487 0.109875
R45120 C8_P_btm.n560 C8_P_btm.n487 0.109875
R45121 C8_P_btm.n567 C8_P_btm.n485 0.109875
R45122 C8_P_btm.n569 C8_P_btm.n485 0.109875
R45123 C8_P_btm.n570 C8_P_btm.n475 0.109875
R45124 C8_P_btm.n572 C8_P_btm.n475 0.109875
R45125 C8_P_btm.n573 C8_P_btm.n472 0.109875
R45126 C8_P_btm.n575 C8_P_btm.n472 0.109875
R45127 C8_P_btm.n582 C8_P_btm.n473 0.109875
R45128 C8_P_btm.n582 C8_P_btm.n581 0.109875
R45129 C8_P_btm.n481 C8_P_btm.n478 0.109875
R45130 C8_P_btm.n479 C8_P_btm.n478 0.109875
R45131 C8_P_btm.n484 C8_P_btm.n477 0.109875
R45132 C8_P_btm.n484 C8_P_btm.n483 0.109875
R45133 C8_P_btm.n593 C8_P_btm.n470 0.109875
R45134 C8_P_btm.n591 C8_P_btm.n470 0.109875
R45135 C8_P_btm.n590 C8_P_btm.n471 0.109875
R45136 C8_P_btm.n588 C8_P_btm.n471 0.109875
R45137 C8_P_btm.n587 C8_P_btm.n583 0.109875
R45138 C8_P_btm.n585 C8_P_btm.n583 0.109875
R45139 C8_P_btm.n615 C8_P_btm.n464 0.109875
R45140 C8_P_btm.n617 C8_P_btm.n464 0.109875
R45141 C8_P_btm.n612 C8_P_btm.n467 0.109875
R45142 C8_P_btm.n614 C8_P_btm.n467 0.109875
R45143 C8_P_btm.n609 C8_P_btm.n468 0.109875
R45144 C8_P_btm.n611 C8_P_btm.n468 0.109875
R45145 C8_P_btm.n604 C8_P_btm.n461 0.109875
R45146 C8_P_btm.n602 C8_P_btm.n461 0.109875
R45147 C8_P_btm.n601 C8_P_btm.n598 0.109875
R45148 C8_P_btm.n599 C8_P_btm.n598 0.109875
R45149 C8_P_btm.n624 C8_P_btm.n465 0.109875
R45150 C8_P_btm.n624 C8_P_btm.n623 0.109875
R45151 C8_P_btm.n629 C8_P_btm.n625 0.109875
R45152 C8_P_btm.n627 C8_P_btm.n625 0.109875
R45153 C8_P_btm.n632 C8_P_btm.n463 0.109875
R45154 C8_P_btm.n630 C8_P_btm.n463 0.109875
R45155 C8_P_btm.n635 C8_P_btm.n462 0.109875
R45156 C8_P_btm.n635 C8_P_btm.n634 0.109875
R45157 C8_P_btm.n638 C8_P_btm.n636 0.109875
R45158 C8_P_btm.n640 C8_P_btm.n636 0.109875
R45159 C8_P_btm.n641 C8_P_btm.n460 0.109875
R45160 C8_P_btm.n643 C8_P_btm.n460 0.109875
R45161 C8_P_btm.n644 C8_P_btm.n459 0.109875
R45162 C8_P_btm.n646 C8_P_btm.n459 0.109875
R45163 C8_P_btm.n654 C8_P_btm.n650 0.109875
R45164 C8_P_btm.n652 C8_P_btm.n650 0.109875
R45165 C8_P_btm.n657 C8_P_btm.n649 0.109875
R45166 C8_P_btm.n655 C8_P_btm.n649 0.109875
R45167 C8_P_btm.n660 C8_P_btm.n457 0.109875
R45168 C8_P_btm.n658 C8_P_btm.n457 0.109875
R45169 C8_P_btm.n663 C8_P_btm.n456 0.109875
R45170 C8_P_btm.n661 C8_P_btm.n456 0.109875
R45171 C8_P_btm.n666 C8_P_btm.n455 0.109875
R45172 C8_P_btm.n664 C8_P_btm.n455 0.109875
R45173 C8_P_btm.n357 C8_P_btm.n135 0.109875
R45174 C8_P_btm.n359 C8_P_btm.n135 0.109875
R45175 C8_P_btm.n354 C8_P_btm.n137 0.109875
R45176 C8_P_btm.n356 C8_P_btm.n137 0.109875
R45177 C8_P_btm.n351 C8_P_btm.n138 0.109875
R45178 C8_P_btm.n353 C8_P_btm.n138 0.109875
R45179 C8_P_btm.n348 C8_P_btm.n139 0.109875
R45180 C8_P_btm.n350 C8_P_btm.n139 0.109875
R45181 C8_P_btm.n345 C8_P_btm.n140 0.109875
R45182 C8_P_btm.n347 C8_P_btm.n140 0.109875
R45183 C8_P_btm.n342 C8_P_btm.n141 0.109875
R45184 C8_P_btm.n344 C8_P_btm.n141 0.109875
R45185 C8_P_btm.n339 C8_P_btm.n142 0.109875
R45186 C8_P_btm.n341 C8_P_btm.n142 0.109875
R45187 C8_P_btm.n336 C8_P_btm.n143 0.109875
R45188 C8_P_btm.n338 C8_P_btm.n143 0.109875
R45189 C8_P_btm.n333 C8_P_btm.n144 0.109875
R45190 C8_P_btm.n335 C8_P_btm.n144 0.109875
R45191 C8_P_btm.n330 C8_P_btm.n145 0.109875
R45192 C8_P_btm.n332 C8_P_btm.n145 0.109875
R45193 C8_P_btm.n327 C8_P_btm.n146 0.109875
R45194 C8_P_btm.n329 C8_P_btm.n146 0.109875
R45195 C8_P_btm.n324 C8_P_btm.n147 0.109875
R45196 C8_P_btm.n326 C8_P_btm.n147 0.109875
R45197 C8_P_btm.n321 C8_P_btm.n148 0.109875
R45198 C8_P_btm.n323 C8_P_btm.n148 0.109875
R45199 C8_P_btm.n318 C8_P_btm.n149 0.109875
R45200 C8_P_btm.n320 C8_P_btm.n149 0.109875
R45201 C8_P_btm.n315 C8_P_btm.n152 0.109875
R45202 C8_P_btm.n317 C8_P_btm.n152 0.109875
R45203 C8_P_btm.n312 C8_P_btm.n153 0.109875
R45204 C8_P_btm.n314 C8_P_btm.n153 0.109875
R45205 C8_P_btm.n309 C8_P_btm.n154 0.109875
R45206 C8_P_btm.n311 C8_P_btm.n154 0.109875
R45207 C8_P_btm.n306 C8_P_btm.n155 0.109875
R45208 C8_P_btm.n308 C8_P_btm.n155 0.109875
R45209 C8_P_btm.n303 C8_P_btm.n156 0.109875
R45210 C8_P_btm.n305 C8_P_btm.n156 0.109875
R45211 C8_P_btm.n300 C8_P_btm.n157 0.109875
R45212 C8_P_btm.n302 C8_P_btm.n157 0.109875
R45213 C8_P_btm.n297 C8_P_btm.n158 0.109875
R45214 C8_P_btm.n299 C8_P_btm.n158 0.109875
R45215 C8_P_btm.n294 C8_P_btm.n159 0.109875
R45216 C8_P_btm.n296 C8_P_btm.n159 0.109875
R45217 C8_P_btm.n291 C8_P_btm.n160 0.109875
R45218 C8_P_btm.n293 C8_P_btm.n160 0.109875
R45219 C8_P_btm.n288 C8_P_btm.n161 0.109875
R45220 C8_P_btm.n290 C8_P_btm.n161 0.109875
R45221 C8_P_btm.n285 C8_P_btm.n162 0.109875
R45222 C8_P_btm.n287 C8_P_btm.n162 0.109875
R45223 C8_P_btm.n282 C8_P_btm.n163 0.109875
R45224 C8_P_btm.n284 C8_P_btm.n163 0.109875
R45225 C8_P_btm.n279 C8_P_btm.n164 0.109875
R45226 C8_P_btm.n281 C8_P_btm.n164 0.109875
R45227 C8_P_btm.n276 C8_P_btm.n274 0.109875
R45228 C8_P_btm.n278 C8_P_btm.n274 0.109875
R45229 C8_P_btm.n273 C8_P_btm.n166 0.109875
R45230 C8_P_btm.n273 C8_P_btm.n272 0.109875
R45231 C8_P_btm.n270 C8_P_btm.n167 0.109875
R45232 C8_P_btm.n268 C8_P_btm.n167 0.109875
R45233 C8_P_btm.n267 C8_P_btm.n168 0.109875
R45234 C8_P_btm.n265 C8_P_btm.n168 0.109875
R45235 C8_P_btm.n264 C8_P_btm.n169 0.109875
R45236 C8_P_btm.n262 C8_P_btm.n169 0.109875
R45237 C8_P_btm.n261 C8_P_btm.n170 0.109875
R45238 C8_P_btm.n259 C8_P_btm.n170 0.109875
R45239 C8_P_btm.n258 C8_P_btm.n171 0.109875
R45240 C8_P_btm.n256 C8_P_btm.n171 0.109875
R45241 C8_P_btm.n255 C8_P_btm.n172 0.109875
R45242 C8_P_btm.n253 C8_P_btm.n172 0.109875
R45243 C8_P_btm.n252 C8_P_btm.n173 0.109875
R45244 C8_P_btm.n250 C8_P_btm.n173 0.109875
R45245 C8_P_btm.n249 C8_P_btm.n174 0.109875
R45246 C8_P_btm.n247 C8_P_btm.n174 0.109875
R45247 C8_P_btm.n246 C8_P_btm.n175 0.109875
R45248 C8_P_btm.n244 C8_P_btm.n175 0.109875
R45249 C8_P_btm.n243 C8_P_btm.n176 0.109875
R45250 C8_P_btm.n241 C8_P_btm.n176 0.109875
R45251 C8_P_btm.n240 C8_P_btm.n177 0.109875
R45252 C8_P_btm.n238 C8_P_btm.n177 0.109875
R45253 C8_P_btm.n237 C8_P_btm.n178 0.109875
R45254 C8_P_btm.n235 C8_P_btm.n178 0.109875
R45255 C8_P_btm.n234 C8_P_btm.n179 0.109875
R45256 C8_P_btm.n232 C8_P_btm.n179 0.109875
R45257 C8_P_btm.n231 C8_P_btm.n180 0.109875
R45258 C8_P_btm.n229 C8_P_btm.n180 0.109875
R45259 C8_P_btm.n228 C8_P_btm.n181 0.109875
R45260 C8_P_btm.n226 C8_P_btm.n181 0.109875
R45261 C8_P_btm.n225 C8_P_btm.n182 0.109875
R45262 C8_P_btm.n223 C8_P_btm.n182 0.109875
R45263 C8_P_btm.n222 C8_P_btm.n183 0.109875
R45264 C8_P_btm.n220 C8_P_btm.n183 0.109875
R45265 C8_P_btm.n219 C8_P_btm.n184 0.109875
R45266 C8_P_btm.n217 C8_P_btm.n184 0.109875
R45267 C8_P_btm.n216 C8_P_btm.n185 0.109875
R45268 C8_P_btm.n214 C8_P_btm.n185 0.109875
R45269 C8_P_btm.n213 C8_P_btm.n186 0.109875
R45270 C8_P_btm.n211 C8_P_btm.n186 0.109875
R45271 C8_P_btm.n210 C8_P_btm.n187 0.109875
R45272 C8_P_btm.n208 C8_P_btm.n187 0.109875
R45273 C8_P_btm.n207 C8_P_btm.n188 0.109875
R45274 C8_P_btm.n205 C8_P_btm.n188 0.109875
R45275 C8_P_btm.n204 C8_P_btm.n189 0.109875
R45276 C8_P_btm.n202 C8_P_btm.n189 0.109875
R45277 C8_P_btm.n201 C8_P_btm.n190 0.109875
R45278 C8_P_btm.n199 C8_P_btm.n190 0.109875
R45279 C8_P_btm.n198 C8_P_btm.n191 0.109875
R45280 C8_P_btm.n196 C8_P_btm.n191 0.109875
R45281 C8_P_btm.n195 C8_P_btm.n192 0.109875
R45282 C8_P_btm.n193 C8_P_btm.n192 0.109875
R45283 C8_P_btm.n365 C8_P_btm.n136 0.109875
R45284 C8_P_btm.n365 C8_P_btm.n364 0.109875
R45285 C8_P_btm.n370 C8_P_btm.n366 0.109875
R45286 C8_P_btm.n368 C8_P_btm.n366 0.109875
R45287 C8_P_btm.n373 C8_P_btm.n134 0.109875
R45288 C8_P_btm.n371 C8_P_btm.n134 0.109875
R45289 C8_P_btm.n376 C8_P_btm.n133 0.109875
R45290 C8_P_btm.n374 C8_P_btm.n133 0.109875
R45291 C8_P_btm.n379 C8_P_btm.n132 0.109875
R45292 C8_P_btm.n377 C8_P_btm.n132 0.109875
R45293 C8_P_btm.n382 C8_P_btm.n131 0.109875
R45294 C8_P_btm.n380 C8_P_btm.n131 0.109875
R45295 C8_P_btm.n385 C8_P_btm.n130 0.109875
R45296 C8_P_btm.n383 C8_P_btm.n130 0.109875
R45297 C8_P_btm.n388 C8_P_btm.n129 0.109875
R45298 C8_P_btm.n386 C8_P_btm.n129 0.109875
R45299 C8_P_btm.n391 C8_P_btm.n128 0.109875
R45300 C8_P_btm.n389 C8_P_btm.n128 0.109875
R45301 C8_P_btm.n394 C8_P_btm.n127 0.109875
R45302 C8_P_btm.n392 C8_P_btm.n127 0.109875
R45303 C8_P_btm.n397 C8_P_btm.n126 0.109875
R45304 C8_P_btm.n395 C8_P_btm.n126 0.109875
R45305 C8_P_btm.n400 C8_P_btm.n125 0.109875
R45306 C8_P_btm.n398 C8_P_btm.n125 0.109875
R45307 C8_P_btm.n403 C8_P_btm.n124 0.109875
R45308 C8_P_btm.n401 C8_P_btm.n124 0.109875
R45309 C8_P_btm.n406 C8_P_btm.n123 0.109875
R45310 C8_P_btm.n404 C8_P_btm.n123 0.109875
R45311 C8_P_btm.n409 C8_P_btm.n122 0.109875
R45312 C8_P_btm.n407 C8_P_btm.n122 0.109875
R45313 C8_P_btm.n412 C8_P_btm.n121 0.109875
R45314 C8_P_btm.n410 C8_P_btm.n121 0.109875
R45315 C8_P_btm.n415 C8_P_btm.n120 0.109875
R45316 C8_P_btm.n413 C8_P_btm.n120 0.109875
R45317 C8_P_btm.n418 C8_P_btm.n119 0.109875
R45318 C8_P_btm.n416 C8_P_btm.n119 0.109875
R45319 C8_P_btm.n421 C8_P_btm.n118 0.109875
R45320 C8_P_btm.n419 C8_P_btm.n118 0.109875
R45321 C8_P_btm.n424 C8_P_btm.n117 0.109875
R45322 C8_P_btm.n422 C8_P_btm.n117 0.109875
R45323 C8_P_btm.n427 C8_P_btm.n116 0.109875
R45324 C8_P_btm.n425 C8_P_btm.n116 0.109875
R45325 C8_P_btm.n430 C8_P_btm.n115 0.109875
R45326 C8_P_btm.n428 C8_P_btm.n115 0.109875
R45327 C8_P_btm.n433 C8_P_btm.n114 0.109875
R45328 C8_P_btm.n431 C8_P_btm.n114 0.109875
R45329 C8_P_btm.n436 C8_P_btm.n113 0.109875
R45330 C8_P_btm.n434 C8_P_btm.n113 0.109875
R45331 C8_P_btm.n439 C8_P_btm.n112 0.109875
R45332 C8_P_btm.n437 C8_P_btm.n112 0.109875
R45333 C8_P_btm.n442 C8_P_btm.n111 0.109875
R45334 C8_P_btm.n440 C8_P_btm.n111 0.109875
R45335 C8_P_btm.n445 C8_P_btm.n110 0.109875
R45336 C8_P_btm.n443 C8_P_btm.n110 0.109875
R45337 C8_P_btm.n448 C8_P_btm.n109 0.109875
R45338 C8_P_btm.n446 C8_P_btm.n109 0.109875
R45339 C8_P_btm.n451 C8_P_btm.n108 0.109875
R45340 C8_P_btm.n449 C8_P_btm.n108 0.109875
R45341 C8_P_btm.n671 C8_P_btm.n106 0.109875
R45342 C8_P_btm.n673 C8_P_btm.n106 0.109875
R45343 C8_P_btm.n674 C8_P_btm.n105 0.109875
R45344 C8_P_btm.n676 C8_P_btm.n105 0.109875
R45345 C8_P_btm.n677 C8_P_btm.n104 0.109875
R45346 C8_P_btm.n679 C8_P_btm.n104 0.109875
R45347 C8_P_btm.n680 C8_P_btm.n103 0.109875
R45348 C8_P_btm.n682 C8_P_btm.n103 0.109875
R45349 C8_P_btm.n683 C8_P_btm.n102 0.109875
R45350 C8_P_btm.n685 C8_P_btm.n102 0.109875
R45351 C8_P_btm.n686 C8_P_btm.n101 0.109875
R45352 C8_P_btm.n688 C8_P_btm.n101 0.109875
R45353 C8_P_btm.n689 C8_P_btm.n100 0.109875
R45354 C8_P_btm.n691 C8_P_btm.n100 0.109875
R45355 C8_P_btm.n692 C8_P_btm.n99 0.109875
R45356 C8_P_btm.n694 C8_P_btm.n99 0.109875
R45357 C8_P_btm.n695 C8_P_btm.n98 0.109875
R45358 C8_P_btm.n697 C8_P_btm.n98 0.109875
R45359 C8_P_btm.n698 C8_P_btm.n97 0.109875
R45360 C8_P_btm.n700 C8_P_btm.n97 0.109875
R45361 C8_P_btm.n701 C8_P_btm.n96 0.109875
R45362 C8_P_btm.n703 C8_P_btm.n96 0.109875
R45363 C8_P_btm.n704 C8_P_btm.n95 0.109875
R45364 C8_P_btm.n706 C8_P_btm.n95 0.109875
R45365 C8_P_btm.n707 C8_P_btm.n94 0.109875
R45366 C8_P_btm.n709 C8_P_btm.n94 0.109875
R45367 C8_P_btm.n710 C8_P_btm.n93 0.109875
R45368 C8_P_btm.n712 C8_P_btm.n93 0.109875
R45369 C8_P_btm.n713 C8_P_btm.n92 0.109875
R45370 C8_P_btm.n715 C8_P_btm.n92 0.109875
R45371 C8_P_btm.n716 C8_P_btm.n91 0.109875
R45372 C8_P_btm.n718 C8_P_btm.n91 0.109875
R45373 C8_P_btm.n719 C8_P_btm.n90 0.109875
R45374 C8_P_btm.n721 C8_P_btm.n90 0.109875
R45375 C8_P_btm.n722 C8_P_btm.n89 0.109875
R45376 C8_P_btm.n724 C8_P_btm.n89 0.109875
R45377 C8_P_btm.n725 C8_P_btm.n88 0.109875
R45378 C8_P_btm.n727 C8_P_btm.n88 0.109875
R45379 C8_P_btm.n728 C8_P_btm.n87 0.109875
R45380 C8_P_btm.n730 C8_P_btm.n87 0.109875
R45381 C8_P_btm.n731 C8_P_btm.n86 0.109875
R45382 C8_P_btm.n733 C8_P_btm.n86 0.109875
R45383 C8_P_btm.n734 C8_P_btm.n85 0.109875
R45384 C8_P_btm.n736 C8_P_btm.n85 0.109875
R45385 C8_P_btm.n737 C8_P_btm.n84 0.109875
R45386 C8_P_btm.n739 C8_P_btm.n84 0.109875
R45387 C8_P_btm.n740 C8_P_btm.n67 0.109875
R45388 C8_P_btm.n742 C8_P_btm.n67 0.109875
R45389 C8_P_btm.n743 C8_P_btm.n66 0.109875
R45390 C8_P_btm.n745 C8_P_btm.n66 0.109875
R45391 C8_P_btm.n746 C8_P_btm.n65 0.109875
R45392 C8_P_btm.n748 C8_P_btm.n65 0.109875
R45393 C8_P_btm.n749 C8_P_btm.n64 0.109875
R45394 C8_P_btm.n751 C8_P_btm.n64 0.109875
R45395 C8_P_btm.n752 C8_P_btm.n61 0.109875
R45396 C8_P_btm.n754 C8_P_btm.n61 0.109875
R45397 C8_P_btm.n761 C8_P_btm.n62 0.109875
R45398 C8_P_btm.n761 C8_P_btm.n760 0.109875
R45399 C8_P_btm.n73 C8_P_btm.n70 0.109875
R45400 C8_P_btm.n71 C8_P_btm.n70 0.109875
R45401 C8_P_btm.n76 C8_P_btm.n69 0.109875
R45402 C8_P_btm.n74 C8_P_btm.n69 0.109875
R45403 C8_P_btm.n79 C8_P_btm.n58 0.109875
R45404 C8_P_btm.n77 C8_P_btm.n58 0.109875
R45405 C8_P_btm.n772 C8_P_btm.n59 0.109875
R45406 C8_P_btm.n770 C8_P_btm.n59 0.109875
R45407 C8_P_btm.n769 C8_P_btm.n60 0.109875
R45408 C8_P_btm.n767 C8_P_btm.n60 0.109875
R45409 C8_P_btm.n766 C8_P_btm.n762 0.109875
R45410 C8_P_btm.n764 C8_P_btm.n762 0.109875
R45411 C8_P_btm.n783 C8_P_btm.n44 0.109875
R45412 C8_P_btm.n785 C8_P_btm.n44 0.109875
R45413 C8_P_btm.n780 C8_P_btm.n47 0.109875
R45414 C8_P_btm.n782 C8_P_btm.n47 0.109875
R45415 C8_P_btm.n777 C8_P_btm.n57 0.109875
R45416 C8_P_btm.n779 C8_P_btm.n57 0.109875
R45417 C8_P_btm.n56 C8_P_btm.n49 0.109875
R45418 C8_P_btm.n56 C8_P_btm.n55 0.109875
R45419 C8_P_btm.n53 C8_P_btm.n50 0.109875
R45420 C8_P_btm.n51 C8_P_btm.n50 0.109875
R45421 C8_P_btm.n792 C8_P_btm.n45 0.109875
R45422 C8_P_btm.n792 C8_P_btm.n791 0.109875
R45423 C8_P_btm.n797 C8_P_btm.n793 0.109875
R45424 C8_P_btm.n795 C8_P_btm.n793 0.109875
R45425 C8_P_btm.n800 C8_P_btm.n43 0.109875
R45426 C8_P_btm.n798 C8_P_btm.n43 0.109875
R45427 C8_P_btm.n803 C8_P_btm.n42 0.109875
R45428 C8_P_btm.n801 C8_P_btm.n42 0.109875
R45429 C8_P_btm.n808 C8_P_btm.n40 0.109875
R45430 C8_P_btm.n810 C8_P_btm.n40 0.109875
R45431 C8_P_btm.n811 C8_P_btm.n30 0.109875
R45432 C8_P_btm.n813 C8_P_btm.n30 0.109875
R45433 C8_P_btm.n814 C8_P_btm.n27 0.109875
R45434 C8_P_btm.n816 C8_P_btm.n27 0.109875
R45435 C8_P_btm.n823 C8_P_btm.n28 0.109875
R45436 C8_P_btm.n823 C8_P_btm.n822 0.109875
R45437 C8_P_btm.n36 C8_P_btm.n33 0.109875
R45438 C8_P_btm.n34 C8_P_btm.n33 0.109875
R45439 C8_P_btm.n39 C8_P_btm.n32 0.109875
R45440 C8_P_btm.n39 C8_P_btm.n38 0.109875
R45441 C8_P_btm.n834 C8_P_btm.n25 0.109875
R45442 C8_P_btm.n832 C8_P_btm.n25 0.109875
R45443 C8_P_btm.n831 C8_P_btm.n26 0.109875
R45444 C8_P_btm.n829 C8_P_btm.n26 0.109875
R45445 C8_P_btm.n828 C8_P_btm.n824 0.109875
R45446 C8_P_btm.n826 C8_P_btm.n824 0.109875
R45447 C8_P_btm.n856 C8_P_btm.n19 0.109875
R45448 C8_P_btm.n858 C8_P_btm.n19 0.109875
R45449 C8_P_btm.n853 C8_P_btm.n22 0.109875
R45450 C8_P_btm.n855 C8_P_btm.n22 0.109875
R45451 C8_P_btm.n850 C8_P_btm.n23 0.109875
R45452 C8_P_btm.n852 C8_P_btm.n23 0.109875
R45453 C8_P_btm.n845 C8_P_btm.n16 0.109875
R45454 C8_P_btm.n843 C8_P_btm.n16 0.109875
R45455 C8_P_btm.n842 C8_P_btm.n839 0.109875
R45456 C8_P_btm.n840 C8_P_btm.n839 0.109875
R45457 C8_P_btm.n865 C8_P_btm.n20 0.109875
R45458 C8_P_btm.n865 C8_P_btm.n864 0.109875
R45459 C8_P_btm.n870 C8_P_btm.n866 0.109875
R45460 C8_P_btm.n868 C8_P_btm.n866 0.109875
R45461 C8_P_btm.n873 C8_P_btm.n18 0.109875
R45462 C8_P_btm.n871 C8_P_btm.n18 0.109875
R45463 C8_P_btm.n876 C8_P_btm.n17 0.109875
R45464 C8_P_btm.n876 C8_P_btm.n875 0.109875
R45465 C8_P_btm.n879 C8_P_btm.n877 0.109875
R45466 C8_P_btm.n881 C8_P_btm.n877 0.109875
R45467 C8_P_btm.n882 C8_P_btm.n15 0.109875
R45468 C8_P_btm.n884 C8_P_btm.n15 0.109875
R45469 C8_P_btm.n885 C8_P_btm.n14 0.109875
R45470 C8_P_btm.n887 C8_P_btm.n14 0.109875
R45471 C8_P_btm.n894 C8_P_btm.n12 0.109875
R45472 C8_P_btm.n892 C8_P_btm.n12 0.109875
R45473 C8_P_btm.n897 C8_P_btm.n11 0.109875
R45474 C8_P_btm.n895 C8_P_btm.n11 0.109875
R45475 C8_P_btm.n900 C8_P_btm.n10 0.109875
R45476 C8_P_btm.n898 C8_P_btm.n10 0.109875
R45477 C8_P_btm.n517 C8_P_btm.n516 0.0556875
R45478 C8_P_btm.n508 C8_P_btm.n503 0.0556875
R45479 C8_P_btm.n533 C8_P_btm.n532 0.0556875
R45480 C8_P_btm.n522 C8_P_btm.n491 0.0556875
R45481 C8_P_btm.n546 C8_P_btm.n545 0.0556875
R45482 C8_P_btm.n535 C8_P_btm.n534 0.0556875
R45483 C8_P_btm.n493 C8_P_btm.n486 0.0556875
R45484 C8_P_btm.n548 C8_P_btm.n547 0.0556875
R45485 C8_P_btm.n553 C8_P_btm.n474 0.0556875
R45486 C8_P_btm.n564 C8_P_btm.n563 0.0556875
R45487 C8_P_btm.n566 C8_P_btm.n565 0.0556875
R45488 C8_P_btm.n577 C8_P_btm.n576 0.0556875
R45489 C8_P_btm.n579 C8_P_btm.n578 0.0556875
R45490 C8_P_btm.n476 C8_P_btm.n469 0.0556875
R45491 C8_P_btm.n595 C8_P_btm.n594 0.0556875
R45492 C8_P_btm.n584 C8_P_btm.n466 0.0556875
R45493 C8_P_btm.n619 C8_P_btm.n618 0.0556875
R45494 C8_P_btm.n608 C8_P_btm.n607 0.0556875
R45495 C8_P_btm.n606 C8_P_btm.n605 0.0556875
R45496 C8_P_btm.n621 C8_P_btm.n620 0.0556875
R45497 C8_P_btm.n626 C8_P_btm.n458 0.0556875
R45498 C8_P_btm.n597 C8_P_btm.n596 0.0556875
R45499 C8_P_btm.n637 C8_P_btm.n454 0.0556875
R45500 C8_P_btm.n648 C8_P_btm.n647 0.0556875
R45501 C8_P_btm.n668 C8_P_btm.n667 0.0556875
R45502 C8_P_btm.n165 C8_P_btm.n107 0.0556875
R45503 C8_P_btm.n362 C8_P_btm.n361 0.0556875
R45504 C8_P_btm.n367 C8_P_btm.n63 0.0556875
R45505 C8_P_btm.n453 C8_P_btm.n452 0.0556875
R45506 C8_P_btm.n670 C8_P_btm.n669 0.0556875
R45507 C8_P_btm.n756 C8_P_btm.n755 0.0556875
R45508 C8_P_btm.n758 C8_P_btm.n757 0.0556875
R45509 C8_P_btm.n774 C8_P_btm.n773 0.0556875
R45510 C8_P_btm.n763 C8_P_btm.n46 0.0556875
R45511 C8_P_btm.n787 C8_P_btm.n786 0.0556875
R45512 C8_P_btm.n776 C8_P_btm.n775 0.0556875
R45513 C8_P_btm.n48 C8_P_btm.n41 0.0556875
R45514 C8_P_btm.n789 C8_P_btm.n788 0.0556875
R45515 C8_P_btm.n794 C8_P_btm.n29 0.0556875
R45516 C8_P_btm.n805 C8_P_btm.n804 0.0556875
R45517 C8_P_btm.n807 C8_P_btm.n806 0.0556875
R45518 C8_P_btm.n818 C8_P_btm.n817 0.0556875
R45519 C8_P_btm.n820 C8_P_btm.n819 0.0556875
R45520 C8_P_btm.n31 C8_P_btm.n24 0.0556875
R45521 C8_P_btm.n836 C8_P_btm.n835 0.0556875
R45522 C8_P_btm.n825 C8_P_btm.n21 0.0556875
R45523 C8_P_btm.n860 C8_P_btm.n859 0.0556875
R45524 C8_P_btm.n849 C8_P_btm.n848 0.0556875
R45525 C8_P_btm.n847 C8_P_btm.n846 0.0556875
R45526 C8_P_btm.n862 C8_P_btm.n861 0.0556875
R45527 C8_P_btm.n867 C8_P_btm.n13 0.0556875
R45528 C8_P_btm.n838 C8_P_btm.n837 0.0556875
R45529 C8_P_btm.n878 C8_P_btm.n9 0.0556875
R45530 C8_P_btm.n889 C8_P_btm.n888 0.0556875
R45531 C8_P_btm.n891 C8_P_btm.n890 0.0556875
R45532 C8_P_btm.n902 C8_P_btm.n901 0.0556875
R45533 C9_N_btm C9_N_btm.n15 82.1151
R45534 C9_N_btm.n2 C9_N_btm.n0 33.0802
R45535 C9_N_btm.n6 C9_N_btm.n5 32.3614
R45536 C9_N_btm.n4 C9_N_btm.n3 32.3614
R45537 C9_N_btm.n2 C9_N_btm.n1 32.3614
R45538 C9_N_btm.n10 C9_N_btm.n6 24.0265
R45539 C9_N_btm.n11 C9_N_btm.t4 23.0826
R45540 C9_N_btm.n14 C9_N_btm.n12 15.4287
R45541 C9_N_btm.n9 C9_N_btm.n7 15.3784
R45542 C9_N_btm.n14 C9_N_btm.n13 14.9755
R45543 C9_N_btm.n9 C9_N_btm.n8 14.894
R45544 C9_N_btm.n15 C9_N_btm.n11 7.16717
R45545 C9_N_btm C9_N_btm.n1886 6.55675
R45546 C9_N_btm.n10 C9_N_btm.n9 5.71404
R45547 C9_N_btm.n15 C9_N_btm.n14 5.62029
R45548 C9_N_btm.n17 C9_N_btm.t530 5.03712
R45549 C9_N_btm.n18 C9_N_btm.t532 5.03712
R45550 C9_N_btm.n19 C9_N_btm.t533 5.03712
R45551 C9_N_btm.n20 C9_N_btm.t536 5.03712
R45552 C9_N_btm.n333 C9_N_btm.t531 5.03712
R45553 C9_N_btm.n332 C9_N_btm.t528 5.03712
R45554 C9_N_btm.n318 C9_N_btm.t535 5.03712
R45555 C9_N_btm.n317 C9_N_btm.t525 5.03712
R45556 C9_N_btm.n315 C9_N_btm.t527 5.03712
R45557 C9_N_btm.n348 C9_N_btm.t534 5.03712
R45558 C9_N_btm.n1870 C9_N_btm.t526 5.03712
R45559 C9_N_btm.n1882 C9_N_btm.n1881 4.60698
R45560 C9_N_btm.n1883 C9_N_btm.n1882 4.60698
R45561 C9_N_btm.n1879 C9_N_btm.n1878 4.60698
R45562 C9_N_btm.n1880 C9_N_btm.n1879 4.60698
R45563 C9_N_btm.n1876 C9_N_btm.n1875 4.60698
R45564 C9_N_btm.n1877 C9_N_btm.n1876 4.60698
R45565 C9_N_btm.n1873 C9_N_btm.n1872 4.60698
R45566 C9_N_btm.n1874 C9_N_btm.n1873 4.60698
R45567 C9_N_btm.n1867 C9_N_btm.n1866 4.60698
R45568 C9_N_btm.n1866 C9_N_btm.n1865 4.60698
R45569 C9_N_btm.n1864 C9_N_btm.n1863 4.60698
R45570 C9_N_btm.n1863 C9_N_btm.n1862 4.60698
R45571 C9_N_btm.n1861 C9_N_btm.n1860 4.60698
R45572 C9_N_btm.n1860 C9_N_btm.n1859 4.60698
R45573 C9_N_btm.n1858 C9_N_btm.n1857 4.60698
R45574 C9_N_btm.n1857 C9_N_btm.n1856 4.60698
R45575 C9_N_btm.n1852 C9_N_btm.n1851 4.60698
R45576 C9_N_btm.n1851 C9_N_btm.n26 4.60698
R45577 C9_N_btm.n1849 C9_N_btm.n1848 4.60698
R45578 C9_N_btm.n1850 C9_N_btm.n1849 4.60698
R45579 C9_N_btm.n1846 C9_N_btm.n1845 4.60698
R45580 C9_N_btm.n1847 C9_N_btm.n1846 4.60698
R45581 C9_N_btm.n1843 C9_N_btm.n1842 4.60698
R45582 C9_N_btm.n1844 C9_N_btm.n1843 4.60698
R45583 C9_N_btm.n1838 C9_N_btm.n1837 4.60698
R45584 C9_N_btm.n1837 C9_N_btm.n30 4.60698
R45585 C9_N_btm.n1809 C9_N_btm.n1808 4.60698
R45586 C9_N_btm.n1810 C9_N_btm.n1809 4.60698
R45587 C9_N_btm.n1812 C9_N_btm.n1811 4.60698
R45588 C9_N_btm.n1813 C9_N_btm.n1812 4.60698
R45589 C9_N_btm.n1815 C9_N_btm.n1814 4.60698
R45590 C9_N_btm.n1816 C9_N_btm.n1815 4.60698
R45591 C9_N_btm.n1823 C9_N_btm.n1822 4.60698
R45592 C9_N_btm.n1822 C9_N_btm.n1821 4.60698
R45593 C9_N_btm.n1826 C9_N_btm.n1825 4.60698
R45594 C9_N_btm.n1825 C9_N_btm.n1824 4.60698
R45595 C9_N_btm.n1829 C9_N_btm.n1828 4.60698
R45596 C9_N_btm.n1828 C9_N_btm.n1827 4.60698
R45597 C9_N_btm.n1832 C9_N_btm.n1831 4.60698
R45598 C9_N_btm.n1831 C9_N_btm.n1830 4.60698
R45599 C9_N_btm.n1791 C9_N_btm.n1790 4.60698
R45600 C9_N_btm.n1792 C9_N_btm.n1791 4.60698
R45601 C9_N_btm.n1794 C9_N_btm.n1793 4.60698
R45602 C9_N_btm.n1795 C9_N_btm.n1794 4.60698
R45603 C9_N_btm.n1797 C9_N_btm.n1796 4.60698
R45604 C9_N_btm.n1798 C9_N_btm.n1797 4.60698
R45605 C9_N_btm.n1800 C9_N_btm.n1799 4.60698
R45606 C9_N_btm.n1801 C9_N_btm.n1800 4.60698
R45607 C9_N_btm.n55 C9_N_btm.n54 4.60698
R45608 C9_N_btm.n54 C9_N_btm.n45 4.60698
R45609 C9_N_btm.n52 C9_N_btm.n51 4.60698
R45610 C9_N_btm.n53 C9_N_btm.n52 4.60698
R45611 C9_N_btm.n49 C9_N_btm.n48 4.60698
R45612 C9_N_btm.n50 C9_N_btm.n49 4.60698
R45613 C9_N_btm.n1786 C9_N_btm.n1785 4.60698
R45614 C9_N_btm.n1785 C9_N_btm.n40 4.60698
R45615 C9_N_btm.n1780 C9_N_btm.n1779 4.60698
R45616 C9_N_btm.n1779 C9_N_btm.n1778 4.60698
R45617 C9_N_btm.n1777 C9_N_btm.n1776 4.60698
R45618 C9_N_btm.n1776 C9_N_btm.n1775 4.60698
R45619 C9_N_btm.n1774 C9_N_btm.n1773 4.60698
R45620 C9_N_btm.n1773 C9_N_btm.n1772 4.60698
R45621 C9_N_btm.n1771 C9_N_btm.n1770 4.60698
R45622 C9_N_btm.n1770 C9_N_btm.n1769 4.60698
R45623 C9_N_btm.n1763 C9_N_btm.n1762 4.60698
R45624 C9_N_btm.n1764 C9_N_btm.n1763 4.60698
R45625 C9_N_btm.n1760 C9_N_btm.n1759 4.60698
R45626 C9_N_btm.n1761 C9_N_btm.n1760 4.60698
R45627 C9_N_btm.n1757 C9_N_btm.n1756 4.60698
R45628 C9_N_btm.n1758 C9_N_btm.n1757 4.60698
R45629 C9_N_btm.n1754 C9_N_btm.n1753 4.60698
R45630 C9_N_btm.n1755 C9_N_btm.n1754 4.60698
R45631 C9_N_btm.n1749 C9_N_btm.n1748 4.60698
R45632 C9_N_btm.n1748 C9_N_btm.n63 4.60698
R45633 C9_N_btm.n72 C9_N_btm.n71 4.60698
R45634 C9_N_btm.n73 C9_N_btm.n72 4.60698
R45635 C9_N_btm.n75 C9_N_btm.n74 4.60698
R45636 C9_N_btm.n76 C9_N_btm.n75 4.60698
R45637 C9_N_btm.n78 C9_N_btm.n77 4.60698
R45638 C9_N_btm.n77 C9_N_btm.n68 4.60698
R45639 C9_N_btm.n1734 C9_N_btm.n1733 4.60698
R45640 C9_N_btm.n1733 C9_N_btm.n1732 4.60698
R45641 C9_N_btm.n1737 C9_N_btm.n1736 4.60698
R45642 C9_N_btm.n1736 C9_N_btm.n1735 4.60698
R45643 C9_N_btm.n1740 C9_N_btm.n1739 4.60698
R45644 C9_N_btm.n1739 C9_N_btm.n1738 4.60698
R45645 C9_N_btm.n1743 C9_N_btm.n1742 4.60698
R45646 C9_N_btm.n1742 C9_N_btm.n1741 4.60698
R45647 C9_N_btm.n1717 C9_N_btm.n1716 4.60698
R45648 C9_N_btm.n1718 C9_N_btm.n1717 4.60698
R45649 C9_N_btm.n1720 C9_N_btm.n1719 4.60698
R45650 C9_N_btm.n1721 C9_N_btm.n1720 4.60698
R45651 C9_N_btm.n1723 C9_N_btm.n1722 4.60698
R45652 C9_N_btm.n1724 C9_N_btm.n1723 4.60698
R45653 C9_N_btm.n1726 C9_N_btm.n1725 4.60698
R45654 C9_N_btm.n1727 C9_N_btm.n1726 4.60698
R45655 C9_N_btm.n101 C9_N_btm.n100 4.60698
R45656 C9_N_btm.n100 C9_N_btm.n91 4.60698
R45657 C9_N_btm.n98 C9_N_btm.n97 4.60698
R45658 C9_N_btm.n99 C9_N_btm.n98 4.60698
R45659 C9_N_btm.n95 C9_N_btm.n94 4.60698
R45660 C9_N_btm.n96 C9_N_btm.n95 4.60698
R45661 C9_N_btm.n1712 C9_N_btm.n1711 4.60698
R45662 C9_N_btm.n1711 C9_N_btm.n86 4.60698
R45663 C9_N_btm.n1706 C9_N_btm.n1705 4.60698
R45664 C9_N_btm.n1705 C9_N_btm.n1704 4.60698
R45665 C9_N_btm.n1703 C9_N_btm.n1702 4.60698
R45666 C9_N_btm.n1702 C9_N_btm.n1701 4.60698
R45667 C9_N_btm.n1700 C9_N_btm.n1699 4.60698
R45668 C9_N_btm.n1699 C9_N_btm.n1698 4.60698
R45669 C9_N_btm.n1697 C9_N_btm.n1696 4.60698
R45670 C9_N_btm.n1696 C9_N_btm.n1695 4.60698
R45671 C9_N_btm.n1689 C9_N_btm.n1688 4.60698
R45672 C9_N_btm.n1690 C9_N_btm.n1689 4.60698
R45673 C9_N_btm.n1686 C9_N_btm.n1685 4.60698
R45674 C9_N_btm.n1687 C9_N_btm.n1686 4.60698
R45675 C9_N_btm.n1683 C9_N_btm.n1682 4.60698
R45676 C9_N_btm.n1684 C9_N_btm.n1683 4.60698
R45677 C9_N_btm.n1680 C9_N_btm.n1679 4.60698
R45678 C9_N_btm.n1681 C9_N_btm.n1680 4.60698
R45679 C9_N_btm.n1675 C9_N_btm.n1674 4.60698
R45680 C9_N_btm.n1674 C9_N_btm.n109 4.60698
R45681 C9_N_btm.n118 C9_N_btm.n117 4.60698
R45682 C9_N_btm.n119 C9_N_btm.n118 4.60698
R45683 C9_N_btm.n121 C9_N_btm.n120 4.60698
R45684 C9_N_btm.n122 C9_N_btm.n121 4.60698
R45685 C9_N_btm.n124 C9_N_btm.n123 4.60698
R45686 C9_N_btm.n123 C9_N_btm.n114 4.60698
R45687 C9_N_btm.n1660 C9_N_btm.n1659 4.60698
R45688 C9_N_btm.n1659 C9_N_btm.n1658 4.60698
R45689 C9_N_btm.n1663 C9_N_btm.n1662 4.60698
R45690 C9_N_btm.n1662 C9_N_btm.n1661 4.60698
R45691 C9_N_btm.n1666 C9_N_btm.n1665 4.60698
R45692 C9_N_btm.n1665 C9_N_btm.n1664 4.60698
R45693 C9_N_btm.n1669 C9_N_btm.n1668 4.60698
R45694 C9_N_btm.n1668 C9_N_btm.n1667 4.60698
R45695 C9_N_btm.n1642 C9_N_btm.n1641 4.60698
R45696 C9_N_btm.n1643 C9_N_btm.n1642 4.60698
R45697 C9_N_btm.n1645 C9_N_btm.n1644 4.60698
R45698 C9_N_btm.n1646 C9_N_btm.n1645 4.60698
R45699 C9_N_btm.n1648 C9_N_btm.n1647 4.60698
R45700 C9_N_btm.n1649 C9_N_btm.n1648 4.60698
R45701 C9_N_btm.n1651 C9_N_btm.n1650 4.60698
R45702 C9_N_btm.n1652 C9_N_btm.n1651 4.60698
R45703 C9_N_btm.n1654 C9_N_btm.n1653 4.60698
R45704 C9_N_btm.n1653 C9_N_btm.n128 4.60698
R45705 C9_N_btm.n674 C9_N_btm.n673 4.60698
R45706 C9_N_btm.n673 C9_N_btm.n672 4.60698
R45707 C9_N_btm.n671 C9_N_btm.n670 4.60698
R45708 C9_N_btm.n670 C9_N_btm.n669 4.60698
R45709 C9_N_btm.n668 C9_N_btm.n667 4.60698
R45710 C9_N_btm.n667 C9_N_btm.n666 4.60698
R45711 C9_N_btm.n665 C9_N_btm.n664 4.60698
R45712 C9_N_btm.n664 C9_N_btm.n663 4.60698
R45713 C9_N_btm.n662 C9_N_btm.n661 4.60698
R45714 C9_N_btm.n661 C9_N_btm.n660 4.60698
R45715 C9_N_btm.n659 C9_N_btm.n658 4.60698
R45716 C9_N_btm.n658 C9_N_btm.n657 4.60698
R45717 C9_N_btm.n656 C9_N_btm.n655 4.60698
R45718 C9_N_btm.n655 C9_N_btm.n654 4.60698
R45719 C9_N_btm.n653 C9_N_btm.n652 4.60698
R45720 C9_N_btm.n652 C9_N_btm.n651 4.60698
R45721 C9_N_btm.n650 C9_N_btm.n649 4.60698
R45722 C9_N_btm.n649 C9_N_btm.n648 4.60698
R45723 C9_N_btm.n647 C9_N_btm.n646 4.60698
R45724 C9_N_btm.n646 C9_N_btm.n645 4.60698
R45725 C9_N_btm.n644 C9_N_btm.n643 4.60698
R45726 C9_N_btm.n643 C9_N_btm.n642 4.60698
R45727 C9_N_btm.n641 C9_N_btm.n640 4.60698
R45728 C9_N_btm.n640 C9_N_btm.n639 4.60698
R45729 C9_N_btm.n638 C9_N_btm.n637 4.60698
R45730 C9_N_btm.n637 C9_N_btm.n636 4.60698
R45731 C9_N_btm.n732 C9_N_btm.n731 4.60698
R45732 C9_N_btm.n733 C9_N_btm.n732 4.60698
R45733 C9_N_btm.n729 C9_N_btm.n728 4.60698
R45734 C9_N_btm.n730 C9_N_btm.n729 4.60698
R45735 C9_N_btm.n726 C9_N_btm.n725 4.60698
R45736 C9_N_btm.n727 C9_N_btm.n726 4.60698
R45737 C9_N_btm.n723 C9_N_btm.n722 4.60698
R45738 C9_N_btm.n724 C9_N_btm.n723 4.60698
R45739 C9_N_btm.n720 C9_N_btm.n719 4.60698
R45740 C9_N_btm.n721 C9_N_btm.n720 4.60698
R45741 C9_N_btm.n717 C9_N_btm.n716 4.60698
R45742 C9_N_btm.n718 C9_N_btm.n717 4.60698
R45743 C9_N_btm.n714 C9_N_btm.n713 4.60698
R45744 C9_N_btm.n715 C9_N_btm.n714 4.60698
R45745 C9_N_btm.n711 C9_N_btm.n710 4.60698
R45746 C9_N_btm.n712 C9_N_btm.n711 4.60698
R45747 C9_N_btm.n708 C9_N_btm.n707 4.60698
R45748 C9_N_btm.n709 C9_N_btm.n708 4.60698
R45749 C9_N_btm.n705 C9_N_btm.n704 4.60698
R45750 C9_N_btm.n706 C9_N_btm.n705 4.60698
R45751 C9_N_btm.n702 C9_N_btm.n701 4.60698
R45752 C9_N_btm.n703 C9_N_btm.n702 4.60698
R45753 C9_N_btm.n699 C9_N_btm.n698 4.60698
R45754 C9_N_btm.n700 C9_N_btm.n699 4.60698
R45755 C9_N_btm.n696 C9_N_btm.n695 4.60698
R45756 C9_N_btm.n697 C9_N_btm.n696 4.60698
R45757 C9_N_btm.n693 C9_N_btm.n692 4.60698
R45758 C9_N_btm.n694 C9_N_btm.n693 4.60698
R45759 C9_N_btm.n690 C9_N_btm.n689 4.60698
R45760 C9_N_btm.n691 C9_N_btm.n690 4.60698
R45761 C9_N_btm.n687 C9_N_btm.n686 4.60698
R45762 C9_N_btm.n688 C9_N_btm.n687 4.60698
R45763 C9_N_btm.n684 C9_N_btm.n683 4.60698
R45764 C9_N_btm.n685 C9_N_btm.n684 4.60698
R45765 C9_N_btm.n681 C9_N_btm.n680 4.60698
R45766 C9_N_btm.n682 C9_N_btm.n681 4.60698
R45767 C9_N_btm.n1637 C9_N_btm.n1636 4.60698
R45768 C9_N_btm.n1636 C9_N_btm.n133 4.60698
R45769 C9_N_btm.n1631 C9_N_btm.n1630 4.60698
R45770 C9_N_btm.n1630 C9_N_btm.n1629 4.60698
R45771 C9_N_btm.n1628 C9_N_btm.n1627 4.60698
R45772 C9_N_btm.n1627 C9_N_btm.n1626 4.60698
R45773 C9_N_btm.n1625 C9_N_btm.n1624 4.60698
R45774 C9_N_btm.n1624 C9_N_btm.n1623 4.60698
R45775 C9_N_btm.n1622 C9_N_btm.n1621 4.60698
R45776 C9_N_btm.n1621 C9_N_btm.n1620 4.60698
R45777 C9_N_btm.n1619 C9_N_btm.n1618 4.60698
R45778 C9_N_btm.n1618 C9_N_btm.n1617 4.60698
R45779 C9_N_btm.n1616 C9_N_btm.n1615 4.60698
R45780 C9_N_btm.n1615 C9_N_btm.n1614 4.60698
R45781 C9_N_btm.n1613 C9_N_btm.n1612 4.60698
R45782 C9_N_btm.n1612 C9_N_btm.n1611 4.60698
R45783 C9_N_btm.n1610 C9_N_btm.n1609 4.60698
R45784 C9_N_btm.n1609 C9_N_btm.n1608 4.60698
R45785 C9_N_btm.n1607 C9_N_btm.n1606 4.60698
R45786 C9_N_btm.n1606 C9_N_btm.n1605 4.60698
R45787 C9_N_btm.n1604 C9_N_btm.n1603 4.60698
R45788 C9_N_btm.n1603 C9_N_btm.n1602 4.60698
R45789 C9_N_btm.n1601 C9_N_btm.n1600 4.60698
R45790 C9_N_btm.n1600 C9_N_btm.n1599 4.60698
R45791 C9_N_btm.n1598 C9_N_btm.n1597 4.60698
R45792 C9_N_btm.n1597 C9_N_btm.n1596 4.60698
R45793 C9_N_btm.n1595 C9_N_btm.n1594 4.60698
R45794 C9_N_btm.n1594 C9_N_btm.n1593 4.60698
R45795 C9_N_btm.n1592 C9_N_btm.n1591 4.60698
R45796 C9_N_btm.n1591 C9_N_btm.n1590 4.60698
R45797 C9_N_btm.n1589 C9_N_btm.n1588 4.60698
R45798 C9_N_btm.n1588 C9_N_btm.n1587 4.60698
R45799 C9_N_btm.n1586 C9_N_btm.n1585 4.60698
R45800 C9_N_btm.n1585 C9_N_btm.n1584 4.60698
R45801 C9_N_btm.n1583 C9_N_btm.n1582 4.60698
R45802 C9_N_btm.n1582 C9_N_btm.n1581 4.60698
R45803 C9_N_btm.n1580 C9_N_btm.n1579 4.60698
R45804 C9_N_btm.n1579 C9_N_btm.n1578 4.60698
R45805 C9_N_btm.n1577 C9_N_btm.n1576 4.60698
R45806 C9_N_btm.n1576 C9_N_btm.n1575 4.60698
R45807 C9_N_btm.n1574 C9_N_btm.n1573 4.60698
R45808 C9_N_btm.n1573 C9_N_btm.n1572 4.60698
R45809 C9_N_btm.n1571 C9_N_btm.n1570 4.60698
R45810 C9_N_btm.n1570 C9_N_btm.n1569 4.60698
R45811 C9_N_btm.n1568 C9_N_btm.n1567 4.60698
R45812 C9_N_btm.n1567 C9_N_btm.n1566 4.60698
R45813 C9_N_btm.n1565 C9_N_btm.n1564 4.60698
R45814 C9_N_btm.n1564 C9_N_btm.n1563 4.60698
R45815 C9_N_btm.n1562 C9_N_btm.n1561 4.60698
R45816 C9_N_btm.n1561 C9_N_btm.n1560 4.60698
R45817 C9_N_btm.n1559 C9_N_btm.n1558 4.60698
R45818 C9_N_btm.n1558 C9_N_btm.n1557 4.60698
R45819 C9_N_btm.n1556 C9_N_btm.n1555 4.60698
R45820 C9_N_btm.n1555 C9_N_btm.n1554 4.60698
R45821 C9_N_btm.n1553 C9_N_btm.n1552 4.60698
R45822 C9_N_btm.n1552 C9_N_btm.n1551 4.60698
R45823 C9_N_btm.n1550 C9_N_btm.n1549 4.60698
R45824 C9_N_btm.n1549 C9_N_btm.n1548 4.60698
R45825 C9_N_btm.n1547 C9_N_btm.n1546 4.60698
R45826 C9_N_btm.n1546 C9_N_btm.n1545 4.60698
R45827 C9_N_btm.n1544 C9_N_btm.n1543 4.60698
R45828 C9_N_btm.n1543 C9_N_btm.n1542 4.60698
R45829 C9_N_btm.n1541 C9_N_btm.n1540 4.60698
R45830 C9_N_btm.n1540 C9_N_btm.n1539 4.60698
R45831 C9_N_btm.n1538 C9_N_btm.n1537 4.60698
R45832 C9_N_btm.n1537 C9_N_btm.n1536 4.60698
R45833 C9_N_btm.n1535 C9_N_btm.n1534 4.60698
R45834 C9_N_btm.n1534 C9_N_btm.n1533 4.60698
R45835 C9_N_btm.n1532 C9_N_btm.n1531 4.60698
R45836 C9_N_btm.n1531 C9_N_btm.n1530 4.60698
R45837 C9_N_btm.n1529 C9_N_btm.n1528 4.60698
R45838 C9_N_btm.n1528 C9_N_btm.n1527 4.60698
R45839 C9_N_btm.n1526 C9_N_btm.n1525 4.60698
R45840 C9_N_btm.n1525 C9_N_btm.n1524 4.60698
R45841 C9_N_btm.n1523 C9_N_btm.n1522 4.60698
R45842 C9_N_btm.n1522 C9_N_btm.n1521 4.60698
R45843 C9_N_btm.n1520 C9_N_btm.n1519 4.60698
R45844 C9_N_btm.n1519 C9_N_btm.n1518 4.60698
R45845 C9_N_btm.n1517 C9_N_btm.n1516 4.60698
R45846 C9_N_btm.n1516 C9_N_btm.n1515 4.60698
R45847 C9_N_btm.n1514 C9_N_btm.n1513 4.60698
R45848 C9_N_btm.n1513 C9_N_btm.n1512 4.60698
R45849 C9_N_btm.n1506 C9_N_btm.n1505 4.60698
R45850 C9_N_btm.n1507 C9_N_btm.n1506 4.60698
R45851 C9_N_btm.n1503 C9_N_btm.n1502 4.60698
R45852 C9_N_btm.n1504 C9_N_btm.n1503 4.60698
R45853 C9_N_btm.n1500 C9_N_btm.n1499 4.60698
R45854 C9_N_btm.n1501 C9_N_btm.n1500 4.60698
R45855 C9_N_btm.n1497 C9_N_btm.n1496 4.60698
R45856 C9_N_btm.n1498 C9_N_btm.n1497 4.60698
R45857 C9_N_btm.n1494 C9_N_btm.n1493 4.60698
R45858 C9_N_btm.n1495 C9_N_btm.n1494 4.60698
R45859 C9_N_btm.n1491 C9_N_btm.n1490 4.60698
R45860 C9_N_btm.n1492 C9_N_btm.n1491 4.60698
R45861 C9_N_btm.n1488 C9_N_btm.n1487 4.60698
R45862 C9_N_btm.n1489 C9_N_btm.n1488 4.60698
R45863 C9_N_btm.n1485 C9_N_btm.n1484 4.60698
R45864 C9_N_btm.n1486 C9_N_btm.n1485 4.60698
R45865 C9_N_btm.n1482 C9_N_btm.n1481 4.60698
R45866 C9_N_btm.n1483 C9_N_btm.n1482 4.60698
R45867 C9_N_btm.n1479 C9_N_btm.n1478 4.60698
R45868 C9_N_btm.n1480 C9_N_btm.n1479 4.60698
R45869 C9_N_btm.n1476 C9_N_btm.n1475 4.60698
R45870 C9_N_btm.n1477 C9_N_btm.n1476 4.60698
R45871 C9_N_btm.n1473 C9_N_btm.n1472 4.60698
R45872 C9_N_btm.n1474 C9_N_btm.n1473 4.60698
R45873 C9_N_btm.n1470 C9_N_btm.n1469 4.60698
R45874 C9_N_btm.n1471 C9_N_btm.n1470 4.60698
R45875 C9_N_btm.n1467 C9_N_btm.n1466 4.60698
R45876 C9_N_btm.n1468 C9_N_btm.n1467 4.60698
R45877 C9_N_btm.n1464 C9_N_btm.n1463 4.60698
R45878 C9_N_btm.n1465 C9_N_btm.n1464 4.60698
R45879 C9_N_btm.n1461 C9_N_btm.n1460 4.60698
R45880 C9_N_btm.n1462 C9_N_btm.n1461 4.60698
R45881 C9_N_btm.n1458 C9_N_btm.n1457 4.60698
R45882 C9_N_btm.n1459 C9_N_btm.n1458 4.60698
R45883 C9_N_btm.n1455 C9_N_btm.n1454 4.60698
R45884 C9_N_btm.n1456 C9_N_btm.n1455 4.60698
R45885 C9_N_btm.n1452 C9_N_btm.n1451 4.60698
R45886 C9_N_btm.n1453 C9_N_btm.n1452 4.60698
R45887 C9_N_btm.n1449 C9_N_btm.n1448 4.60698
R45888 C9_N_btm.n1450 C9_N_btm.n1449 4.60698
R45889 C9_N_btm.n1446 C9_N_btm.n1445 4.60698
R45890 C9_N_btm.n1447 C9_N_btm.n1446 4.60698
R45891 C9_N_btm.n1443 C9_N_btm.n1442 4.60698
R45892 C9_N_btm.n1444 C9_N_btm.n1443 4.60698
R45893 C9_N_btm.n1440 C9_N_btm.n1439 4.60698
R45894 C9_N_btm.n1441 C9_N_btm.n1440 4.60698
R45895 C9_N_btm.n1437 C9_N_btm.n1436 4.60698
R45896 C9_N_btm.n1438 C9_N_btm.n1437 4.60698
R45897 C9_N_btm.n1434 C9_N_btm.n1433 4.60698
R45898 C9_N_btm.n1435 C9_N_btm.n1434 4.60698
R45899 C9_N_btm.n1431 C9_N_btm.n1430 4.60698
R45900 C9_N_btm.n1432 C9_N_btm.n1431 4.60698
R45901 C9_N_btm.n1428 C9_N_btm.n1427 4.60698
R45902 C9_N_btm.n1429 C9_N_btm.n1428 4.60698
R45903 C9_N_btm.n1425 C9_N_btm.n1424 4.60698
R45904 C9_N_btm.n1426 C9_N_btm.n1425 4.60698
R45905 C9_N_btm.n1422 C9_N_btm.n1421 4.60698
R45906 C9_N_btm.n1423 C9_N_btm.n1422 4.60698
R45907 C9_N_btm.n1419 C9_N_btm.n1418 4.60698
R45908 C9_N_btm.n1420 C9_N_btm.n1419 4.60698
R45909 C9_N_btm.n1416 C9_N_btm.n1415 4.60698
R45910 C9_N_btm.n1417 C9_N_btm.n1416 4.60698
R45911 C9_N_btm.n1413 C9_N_btm.n1412 4.60698
R45912 C9_N_btm.n1414 C9_N_btm.n1413 4.60698
R45913 C9_N_btm.n1410 C9_N_btm.n1409 4.60698
R45914 C9_N_btm.n1411 C9_N_btm.n1410 4.60698
R45915 C9_N_btm.n1407 C9_N_btm.n1406 4.60698
R45916 C9_N_btm.n1408 C9_N_btm.n1407 4.60698
R45917 C9_N_btm.n1404 C9_N_btm.n1403 4.60698
R45918 C9_N_btm.n1405 C9_N_btm.n1404 4.60698
R45919 C9_N_btm.n1401 C9_N_btm.n1400 4.60698
R45920 C9_N_btm.n1402 C9_N_btm.n1401 4.60698
R45921 C9_N_btm.n1398 C9_N_btm.n1397 4.60698
R45922 C9_N_btm.n1399 C9_N_btm.n1398 4.60698
R45923 C9_N_btm.n1395 C9_N_btm.n1394 4.60698
R45924 C9_N_btm.n1396 C9_N_btm.n1395 4.60698
R45925 C9_N_btm.n1392 C9_N_btm.n1391 4.60698
R45926 C9_N_btm.n1393 C9_N_btm.n1392 4.60698
R45927 C9_N_btm.n1389 C9_N_btm.n1388 4.60698
R45928 C9_N_btm.n1390 C9_N_btm.n1389 4.60698
R45929 C9_N_btm.n1384 C9_N_btm.n1383 4.60698
R45930 C9_N_btm.n1383 C9_N_btm.n840 4.60698
R45931 C9_N_btm.n921 C9_N_btm.n920 4.60698
R45932 C9_N_btm.n922 C9_N_btm.n921 4.60698
R45933 C9_N_btm.n924 C9_N_btm.n923 4.60698
R45934 C9_N_btm.n925 C9_N_btm.n924 4.60698
R45935 C9_N_btm.n927 C9_N_btm.n926 4.60698
R45936 C9_N_btm.n928 C9_N_btm.n927 4.60698
R45937 C9_N_btm.n930 C9_N_btm.n929 4.60698
R45938 C9_N_btm.n931 C9_N_btm.n930 4.60698
R45939 C9_N_btm.n933 C9_N_btm.n932 4.60698
R45940 C9_N_btm.n934 C9_N_btm.n933 4.60698
R45941 C9_N_btm.n936 C9_N_btm.n935 4.60698
R45942 C9_N_btm.n937 C9_N_btm.n936 4.60698
R45943 C9_N_btm.n939 C9_N_btm.n938 4.60698
R45944 C9_N_btm.n940 C9_N_btm.n939 4.60698
R45945 C9_N_btm.n942 C9_N_btm.n941 4.60698
R45946 C9_N_btm.n943 C9_N_btm.n942 4.60698
R45947 C9_N_btm.n945 C9_N_btm.n944 4.60698
R45948 C9_N_btm.n946 C9_N_btm.n945 4.60698
R45949 C9_N_btm.n948 C9_N_btm.n947 4.60698
R45950 C9_N_btm.n949 C9_N_btm.n948 4.60698
R45951 C9_N_btm.n951 C9_N_btm.n950 4.60698
R45952 C9_N_btm.n952 C9_N_btm.n951 4.60698
R45953 C9_N_btm.n954 C9_N_btm.n953 4.60698
R45954 C9_N_btm.n955 C9_N_btm.n954 4.60698
R45955 C9_N_btm.n957 C9_N_btm.n956 4.60698
R45956 C9_N_btm.n958 C9_N_btm.n957 4.60698
R45957 C9_N_btm.n960 C9_N_btm.n959 4.60698
R45958 C9_N_btm.n961 C9_N_btm.n960 4.60698
R45959 C9_N_btm.n963 C9_N_btm.n962 4.60698
R45960 C9_N_btm.n964 C9_N_btm.n963 4.60698
R45961 C9_N_btm.n966 C9_N_btm.n965 4.60698
R45962 C9_N_btm.n967 C9_N_btm.n966 4.60698
R45963 C9_N_btm.n969 C9_N_btm.n968 4.60698
R45964 C9_N_btm.n970 C9_N_btm.n969 4.60698
R45965 C9_N_btm.n972 C9_N_btm.n971 4.60698
R45966 C9_N_btm.n973 C9_N_btm.n972 4.60698
R45967 C9_N_btm.n975 C9_N_btm.n974 4.60698
R45968 C9_N_btm.n976 C9_N_btm.n975 4.60698
R45969 C9_N_btm.n978 C9_N_btm.n977 4.60698
R45970 C9_N_btm.n979 C9_N_btm.n978 4.60698
R45971 C9_N_btm.n981 C9_N_btm.n980 4.60698
R45972 C9_N_btm.n982 C9_N_btm.n981 4.60698
R45973 C9_N_btm.n984 C9_N_btm.n983 4.60698
R45974 C9_N_btm.n985 C9_N_btm.n984 4.60698
R45975 C9_N_btm.n987 C9_N_btm.n986 4.60698
R45976 C9_N_btm.n988 C9_N_btm.n987 4.60698
R45977 C9_N_btm.n990 C9_N_btm.n989 4.60698
R45978 C9_N_btm.n991 C9_N_btm.n990 4.60698
R45979 C9_N_btm.n993 C9_N_btm.n992 4.60698
R45980 C9_N_btm.n994 C9_N_btm.n993 4.60698
R45981 C9_N_btm.n996 C9_N_btm.n995 4.60698
R45982 C9_N_btm.n997 C9_N_btm.n996 4.60698
R45983 C9_N_btm.n999 C9_N_btm.n998 4.60698
R45984 C9_N_btm.n1000 C9_N_btm.n999 4.60698
R45985 C9_N_btm.n1002 C9_N_btm.n1001 4.60698
R45986 C9_N_btm.n1003 C9_N_btm.n1002 4.60698
R45987 C9_N_btm.n1005 C9_N_btm.n1004 4.60698
R45988 C9_N_btm.n1006 C9_N_btm.n1005 4.60698
R45989 C9_N_btm.n1008 C9_N_btm.n1007 4.60698
R45990 C9_N_btm.n1009 C9_N_btm.n1008 4.60698
R45991 C9_N_btm.n1011 C9_N_btm.n1010 4.60698
R45992 C9_N_btm.n1012 C9_N_btm.n1011 4.60698
R45993 C9_N_btm.n1014 C9_N_btm.n1013 4.60698
R45994 C9_N_btm.n1015 C9_N_btm.n1014 4.60698
R45995 C9_N_btm.n1017 C9_N_btm.n1016 4.60698
R45996 C9_N_btm.n1018 C9_N_btm.n1017 4.60698
R45997 C9_N_btm.n1020 C9_N_btm.n1019 4.60698
R45998 C9_N_btm.n1021 C9_N_btm.n1020 4.60698
R45999 C9_N_btm.n1023 C9_N_btm.n1022 4.60698
R46000 C9_N_btm.n1024 C9_N_btm.n1023 4.60698
R46001 C9_N_btm.n1026 C9_N_btm.n1025 4.60698
R46002 C9_N_btm.n1027 C9_N_btm.n1026 4.60698
R46003 C9_N_btm.n1029 C9_N_btm.n1028 4.60698
R46004 C9_N_btm.n1030 C9_N_btm.n1029 4.60698
R46005 C9_N_btm.n1032 C9_N_btm.n1031 4.60698
R46006 C9_N_btm.n1033 C9_N_btm.n1032 4.60698
R46007 C9_N_btm.n1035 C9_N_btm.n1034 4.60698
R46008 C9_N_btm.n1034 C9_N_btm.n881 4.60698
R46009 C9_N_btm.n1261 C9_N_btm.n1260 4.60698
R46010 C9_N_btm.n1260 C9_N_btm.n1259 4.60698
R46011 C9_N_btm.n1264 C9_N_btm.n1263 4.60698
R46012 C9_N_btm.n1263 C9_N_btm.n1262 4.60698
R46013 C9_N_btm.n1267 C9_N_btm.n1266 4.60698
R46014 C9_N_btm.n1266 C9_N_btm.n1265 4.60698
R46015 C9_N_btm.n1270 C9_N_btm.n1269 4.60698
R46016 C9_N_btm.n1269 C9_N_btm.n1268 4.60698
R46017 C9_N_btm.n1273 C9_N_btm.n1272 4.60698
R46018 C9_N_btm.n1272 C9_N_btm.n1271 4.60698
R46019 C9_N_btm.n1276 C9_N_btm.n1275 4.60698
R46020 C9_N_btm.n1275 C9_N_btm.n1274 4.60698
R46021 C9_N_btm.n1279 C9_N_btm.n1278 4.60698
R46022 C9_N_btm.n1278 C9_N_btm.n1277 4.60698
R46023 C9_N_btm.n1282 C9_N_btm.n1281 4.60698
R46024 C9_N_btm.n1281 C9_N_btm.n1280 4.60698
R46025 C9_N_btm.n1285 C9_N_btm.n1284 4.60698
R46026 C9_N_btm.n1284 C9_N_btm.n1283 4.60698
R46027 C9_N_btm.n1288 C9_N_btm.n1287 4.60698
R46028 C9_N_btm.n1287 C9_N_btm.n1286 4.60698
R46029 C9_N_btm.n1291 C9_N_btm.n1290 4.60698
R46030 C9_N_btm.n1290 C9_N_btm.n1289 4.60698
R46031 C9_N_btm.n1294 C9_N_btm.n1293 4.60698
R46032 C9_N_btm.n1293 C9_N_btm.n1292 4.60698
R46033 C9_N_btm.n1297 C9_N_btm.n1296 4.60698
R46034 C9_N_btm.n1296 C9_N_btm.n1295 4.60698
R46035 C9_N_btm.n1300 C9_N_btm.n1299 4.60698
R46036 C9_N_btm.n1299 C9_N_btm.n1298 4.60698
R46037 C9_N_btm.n1303 C9_N_btm.n1302 4.60698
R46038 C9_N_btm.n1302 C9_N_btm.n1301 4.60698
R46039 C9_N_btm.n1306 C9_N_btm.n1305 4.60698
R46040 C9_N_btm.n1305 C9_N_btm.n1304 4.60698
R46041 C9_N_btm.n1309 C9_N_btm.n1308 4.60698
R46042 C9_N_btm.n1308 C9_N_btm.n1307 4.60698
R46043 C9_N_btm.n1312 C9_N_btm.n1311 4.60698
R46044 C9_N_btm.n1311 C9_N_btm.n1310 4.60698
R46045 C9_N_btm.n1315 C9_N_btm.n1314 4.60698
R46046 C9_N_btm.n1314 C9_N_btm.n1313 4.60698
R46047 C9_N_btm.n1318 C9_N_btm.n1317 4.60698
R46048 C9_N_btm.n1317 C9_N_btm.n1316 4.60698
R46049 C9_N_btm.n1321 C9_N_btm.n1320 4.60698
R46050 C9_N_btm.n1320 C9_N_btm.n1319 4.60698
R46051 C9_N_btm.n1324 C9_N_btm.n1323 4.60698
R46052 C9_N_btm.n1323 C9_N_btm.n1322 4.60698
R46053 C9_N_btm.n1327 C9_N_btm.n1326 4.60698
R46054 C9_N_btm.n1326 C9_N_btm.n1325 4.60698
R46055 C9_N_btm.n1330 C9_N_btm.n1329 4.60698
R46056 C9_N_btm.n1329 C9_N_btm.n1328 4.60698
R46057 C9_N_btm.n1333 C9_N_btm.n1332 4.60698
R46058 C9_N_btm.n1332 C9_N_btm.n1331 4.60698
R46059 C9_N_btm.n1336 C9_N_btm.n1335 4.60698
R46060 C9_N_btm.n1335 C9_N_btm.n1334 4.60698
R46061 C9_N_btm.n1339 C9_N_btm.n1338 4.60698
R46062 C9_N_btm.n1338 C9_N_btm.n1337 4.60698
R46063 C9_N_btm.n1342 C9_N_btm.n1341 4.60698
R46064 C9_N_btm.n1341 C9_N_btm.n1340 4.60698
R46065 C9_N_btm.n1345 C9_N_btm.n1344 4.60698
R46066 C9_N_btm.n1344 C9_N_btm.n1343 4.60698
R46067 C9_N_btm.n1348 C9_N_btm.n1347 4.60698
R46068 C9_N_btm.n1347 C9_N_btm.n1346 4.60698
R46069 C9_N_btm.n1351 C9_N_btm.n1350 4.60698
R46070 C9_N_btm.n1350 C9_N_btm.n1349 4.60698
R46071 C9_N_btm.n1354 C9_N_btm.n1353 4.60698
R46072 C9_N_btm.n1353 C9_N_btm.n1352 4.60698
R46073 C9_N_btm.n1357 C9_N_btm.n1356 4.60698
R46074 C9_N_btm.n1356 C9_N_btm.n1355 4.60698
R46075 C9_N_btm.n1360 C9_N_btm.n1359 4.60698
R46076 C9_N_btm.n1359 C9_N_btm.n1358 4.60698
R46077 C9_N_btm.n1363 C9_N_btm.n1362 4.60698
R46078 C9_N_btm.n1362 C9_N_btm.n1361 4.60698
R46079 C9_N_btm.n1366 C9_N_btm.n1365 4.60698
R46080 C9_N_btm.n1365 C9_N_btm.n1364 4.60698
R46081 C9_N_btm.n1369 C9_N_btm.n1368 4.60698
R46082 C9_N_btm.n1368 C9_N_btm.n1367 4.60698
R46083 C9_N_btm.n1372 C9_N_btm.n1371 4.60698
R46084 C9_N_btm.n1371 C9_N_btm.n1370 4.60698
R46085 C9_N_btm.n1375 C9_N_btm.n1374 4.60698
R46086 C9_N_btm.n1374 C9_N_btm.n1373 4.60698
R46087 C9_N_btm.n1378 C9_N_btm.n1377 4.60698
R46088 C9_N_btm.n1377 C9_N_btm.n1376 4.60698
R46089 C9_N_btm.n1138 C9_N_btm.n1137 4.60698
R46090 C9_N_btm.n1137 C9_N_btm.n1136 4.60698
R46091 C9_N_btm.n1141 C9_N_btm.n1140 4.60698
R46092 C9_N_btm.n1140 C9_N_btm.n1139 4.60698
R46093 C9_N_btm.n1144 C9_N_btm.n1143 4.60698
R46094 C9_N_btm.n1143 C9_N_btm.n1142 4.60698
R46095 C9_N_btm.n1147 C9_N_btm.n1146 4.60698
R46096 C9_N_btm.n1146 C9_N_btm.n1145 4.60698
R46097 C9_N_btm.n1150 C9_N_btm.n1149 4.60698
R46098 C9_N_btm.n1149 C9_N_btm.n1148 4.60698
R46099 C9_N_btm.n1153 C9_N_btm.n1152 4.60698
R46100 C9_N_btm.n1152 C9_N_btm.n1151 4.60698
R46101 C9_N_btm.n1156 C9_N_btm.n1155 4.60698
R46102 C9_N_btm.n1155 C9_N_btm.n1154 4.60698
R46103 C9_N_btm.n1159 C9_N_btm.n1158 4.60698
R46104 C9_N_btm.n1158 C9_N_btm.n1157 4.60698
R46105 C9_N_btm.n1162 C9_N_btm.n1161 4.60698
R46106 C9_N_btm.n1161 C9_N_btm.n1160 4.60698
R46107 C9_N_btm.n1165 C9_N_btm.n1164 4.60698
R46108 C9_N_btm.n1164 C9_N_btm.n1163 4.60698
R46109 C9_N_btm.n1168 C9_N_btm.n1167 4.60698
R46110 C9_N_btm.n1167 C9_N_btm.n1166 4.60698
R46111 C9_N_btm.n1171 C9_N_btm.n1170 4.60698
R46112 C9_N_btm.n1170 C9_N_btm.n1169 4.60698
R46113 C9_N_btm.n1173 C9_N_btm.n1172 4.60698
R46114 C9_N_btm.n1174 C9_N_btm.n1173 4.60698
R46115 C9_N_btm.n1176 C9_N_btm.n1175 4.60698
R46116 C9_N_btm.n1177 C9_N_btm.n1176 4.60698
R46117 C9_N_btm.n1179 C9_N_btm.n1178 4.60698
R46118 C9_N_btm.n1180 C9_N_btm.n1179 4.60698
R46119 C9_N_btm.n1182 C9_N_btm.n1181 4.60698
R46120 C9_N_btm.n1183 C9_N_btm.n1182 4.60698
R46121 C9_N_btm.n1185 C9_N_btm.n1184 4.60698
R46122 C9_N_btm.n1186 C9_N_btm.n1185 4.60698
R46123 C9_N_btm.n1188 C9_N_btm.n1187 4.60698
R46124 C9_N_btm.n1189 C9_N_btm.n1188 4.60698
R46125 C9_N_btm.n1191 C9_N_btm.n1190 4.60698
R46126 C9_N_btm.n1192 C9_N_btm.n1191 4.60698
R46127 C9_N_btm.n1194 C9_N_btm.n1193 4.60698
R46128 C9_N_btm.n1195 C9_N_btm.n1194 4.60698
R46129 C9_N_btm.n1197 C9_N_btm.n1196 4.60698
R46130 C9_N_btm.n1198 C9_N_btm.n1197 4.60698
R46131 C9_N_btm.n1200 C9_N_btm.n1199 4.60698
R46132 C9_N_btm.n1201 C9_N_btm.n1200 4.60698
R46133 C9_N_btm.n1203 C9_N_btm.n1202 4.60698
R46134 C9_N_btm.n1204 C9_N_btm.n1203 4.60698
R46135 C9_N_btm.n1206 C9_N_btm.n1205 4.60698
R46136 C9_N_btm.n1207 C9_N_btm.n1206 4.60698
R46137 C9_N_btm.n1209 C9_N_btm.n1208 4.60698
R46138 C9_N_btm.n1210 C9_N_btm.n1209 4.60698
R46139 C9_N_btm.n1212 C9_N_btm.n1211 4.60698
R46140 C9_N_btm.n1213 C9_N_btm.n1212 4.60698
R46141 C9_N_btm.n1215 C9_N_btm.n1214 4.60698
R46142 C9_N_btm.n1216 C9_N_btm.n1215 4.60698
R46143 C9_N_btm.n1219 C9_N_btm.n1218 4.60698
R46144 C9_N_btm.n1218 C9_N_btm.n1217 4.60698
R46145 C9_N_btm.n1081 C9_N_btm.n1080 4.60698
R46146 C9_N_btm.n1082 C9_N_btm.n1081 4.60698
R46147 C9_N_btm.n1084 C9_N_btm.n1083 4.60698
R46148 C9_N_btm.n1085 C9_N_btm.n1084 4.60698
R46149 C9_N_btm.n1087 C9_N_btm.n1086 4.60698
R46150 C9_N_btm.n1088 C9_N_btm.n1087 4.60698
R46151 C9_N_btm.n1090 C9_N_btm.n1089 4.60698
R46152 C9_N_btm.n1091 C9_N_btm.n1090 4.60698
R46153 C9_N_btm.n1093 C9_N_btm.n1092 4.60698
R46154 C9_N_btm.n1094 C9_N_btm.n1093 4.60698
R46155 C9_N_btm.n1096 C9_N_btm.n1095 4.60698
R46156 C9_N_btm.n1097 C9_N_btm.n1096 4.60698
R46157 C9_N_btm.n1099 C9_N_btm.n1098 4.60698
R46158 C9_N_btm.n1100 C9_N_btm.n1099 4.60698
R46159 C9_N_btm.n1102 C9_N_btm.n1101 4.60698
R46160 C9_N_btm.n1103 C9_N_btm.n1102 4.60698
R46161 C9_N_btm.n1105 C9_N_btm.n1104 4.60698
R46162 C9_N_btm.n1106 C9_N_btm.n1105 4.60698
R46163 C9_N_btm.n1108 C9_N_btm.n1107 4.60698
R46164 C9_N_btm.n1109 C9_N_btm.n1108 4.60698
R46165 C9_N_btm.n1111 C9_N_btm.n1110 4.60698
R46166 C9_N_btm.n1112 C9_N_btm.n1111 4.60698
R46167 C9_N_btm.n1114 C9_N_btm.n1113 4.60698
R46168 C9_N_btm.n1115 C9_N_btm.n1114 4.60698
R46169 C9_N_btm.n1117 C9_N_btm.n1116 4.60698
R46170 C9_N_btm.n1118 C9_N_btm.n1117 4.60698
R46171 C9_N_btm.n1120 C9_N_btm.n1119 4.60698
R46172 C9_N_btm.n1121 C9_N_btm.n1120 4.60698
R46173 C9_N_btm.n1222 C9_N_btm.n1221 4.60698
R46174 C9_N_btm.n1221 C9_N_btm.n1220 4.60698
R46175 C9_N_btm.n1225 C9_N_btm.n1224 4.60698
R46176 C9_N_btm.n1224 C9_N_btm.n1223 4.60698
R46177 C9_N_btm.n1228 C9_N_btm.n1227 4.60698
R46178 C9_N_btm.n1227 C9_N_btm.n1226 4.60698
R46179 C9_N_btm.n1231 C9_N_btm.n1230 4.60698
R46180 C9_N_btm.n1230 C9_N_btm.n1229 4.60698
R46181 C9_N_btm.n1234 C9_N_btm.n1233 4.60698
R46182 C9_N_btm.n1233 C9_N_btm.n1232 4.60698
R46183 C9_N_btm.n1237 C9_N_btm.n1236 4.60698
R46184 C9_N_btm.n1236 C9_N_btm.n1235 4.60698
R46185 C9_N_btm.n1240 C9_N_btm.n1239 4.60698
R46186 C9_N_btm.n1239 C9_N_btm.n1238 4.60698
R46187 C9_N_btm.n1243 C9_N_btm.n1242 4.60698
R46188 C9_N_btm.n1242 C9_N_btm.n1241 4.60698
R46189 C9_N_btm.n1246 C9_N_btm.n1245 4.60698
R46190 C9_N_btm.n1245 C9_N_btm.n1244 4.60698
R46191 C9_N_btm.n1249 C9_N_btm.n1248 4.60698
R46192 C9_N_btm.n1248 C9_N_btm.n1247 4.60698
R46193 C9_N_btm.n1252 C9_N_btm.n1251 4.60698
R46194 C9_N_btm.n1251 C9_N_btm.n1250 4.60698
R46195 C9_N_btm.n1255 C9_N_btm.n1254 4.60698
R46196 C9_N_btm.n1254 C9_N_btm.n1253 4.60698
R46197 C9_N_btm.n795 C9_N_btm.n794 4.60698
R46198 C9_N_btm.n796 C9_N_btm.n795 4.60698
R46199 C9_N_btm.n792 C9_N_btm.n791 4.60698
R46200 C9_N_btm.n793 C9_N_btm.n792 4.60698
R46201 C9_N_btm.n789 C9_N_btm.n788 4.60698
R46202 C9_N_btm.n790 C9_N_btm.n789 4.60698
R46203 C9_N_btm.n786 C9_N_btm.n785 4.60698
R46204 C9_N_btm.n787 C9_N_btm.n786 4.60698
R46205 C9_N_btm.n783 C9_N_btm.n782 4.60698
R46206 C9_N_btm.n784 C9_N_btm.n783 4.60698
R46207 C9_N_btm.n780 C9_N_btm.n779 4.60698
R46208 C9_N_btm.n781 C9_N_btm.n780 4.60698
R46209 C9_N_btm.n777 C9_N_btm.n776 4.60698
R46210 C9_N_btm.n778 C9_N_btm.n777 4.60698
R46211 C9_N_btm.n774 C9_N_btm.n773 4.60698
R46212 C9_N_btm.n775 C9_N_btm.n774 4.60698
R46213 C9_N_btm.n771 C9_N_btm.n770 4.60698
R46214 C9_N_btm.n772 C9_N_btm.n771 4.60698
R46215 C9_N_btm.n768 C9_N_btm.n767 4.60698
R46216 C9_N_btm.n769 C9_N_btm.n768 4.60698
R46217 C9_N_btm.n765 C9_N_btm.n764 4.60698
R46218 C9_N_btm.n766 C9_N_btm.n765 4.60698
R46219 C9_N_btm.n762 C9_N_btm.n761 4.60698
R46220 C9_N_btm.n763 C9_N_btm.n762 4.60698
R46221 C9_N_btm.n759 C9_N_btm.n758 4.60698
R46222 C9_N_btm.n760 C9_N_btm.n759 4.60698
R46223 C9_N_btm.n756 C9_N_btm.n755 4.60698
R46224 C9_N_btm.n757 C9_N_btm.n756 4.60698
R46225 C9_N_btm.n753 C9_N_btm.n752 4.60698
R46226 C9_N_btm.n754 C9_N_btm.n753 4.60698
R46227 C9_N_btm.n750 C9_N_btm.n749 4.60698
R46228 C9_N_btm.n751 C9_N_btm.n750 4.60698
R46229 C9_N_btm.n747 C9_N_btm.n746 4.60698
R46230 C9_N_btm.n748 C9_N_btm.n747 4.60698
R46231 C9_N_btm.n744 C9_N_btm.n743 4.60698
R46232 C9_N_btm.n745 C9_N_btm.n744 4.60698
R46233 C9_N_btm.n741 C9_N_btm.n740 4.60698
R46234 C9_N_btm.n742 C9_N_btm.n741 4.60698
R46235 C9_N_btm.n605 C9_N_btm.n604 4.60698
R46236 C9_N_btm.n604 C9_N_btm.n603 4.60698
R46237 C9_N_btm.n602 C9_N_btm.n601 4.60698
R46238 C9_N_btm.n601 C9_N_btm.n600 4.60698
R46239 C9_N_btm.n599 C9_N_btm.n598 4.60698
R46240 C9_N_btm.n598 C9_N_btm.n597 4.60698
R46241 C9_N_btm.n596 C9_N_btm.n595 4.60698
R46242 C9_N_btm.n595 C9_N_btm.n594 4.60698
R46243 C9_N_btm.n593 C9_N_btm.n592 4.60698
R46244 C9_N_btm.n592 C9_N_btm.n591 4.60698
R46245 C9_N_btm.n590 C9_N_btm.n589 4.60698
R46246 C9_N_btm.n589 C9_N_btm.n588 4.60698
R46247 C9_N_btm.n587 C9_N_btm.n586 4.60698
R46248 C9_N_btm.n586 C9_N_btm.n585 4.60698
R46249 C9_N_btm.n584 C9_N_btm.n583 4.60698
R46250 C9_N_btm.n583 C9_N_btm.n582 4.60698
R46251 C9_N_btm.n581 C9_N_btm.n580 4.60698
R46252 C9_N_btm.n580 C9_N_btm.n579 4.60698
R46253 C9_N_btm.n578 C9_N_btm.n577 4.60698
R46254 C9_N_btm.n577 C9_N_btm.n576 4.60698
R46255 C9_N_btm.n575 C9_N_btm.n574 4.60698
R46256 C9_N_btm.n574 C9_N_btm.n573 4.60698
R46257 C9_N_btm.n572 C9_N_btm.n571 4.60698
R46258 C9_N_btm.n571 C9_N_btm.n570 4.60698
R46259 C9_N_btm.n569 C9_N_btm.n568 4.60698
R46260 C9_N_btm.n568 C9_N_btm.n567 4.60698
R46261 C9_N_btm.n566 C9_N_btm.n565 4.60698
R46262 C9_N_btm.n565 C9_N_btm.n564 4.60698
R46263 C9_N_btm.n563 C9_N_btm.n562 4.60698
R46264 C9_N_btm.n562 C9_N_btm.n561 4.60698
R46265 C9_N_btm.n560 C9_N_btm.n559 4.60698
R46266 C9_N_btm.n559 C9_N_btm.n558 4.60698
R46267 C9_N_btm.n557 C9_N_btm.n556 4.60698
R46268 C9_N_btm.n556 C9_N_btm.n555 4.60698
R46269 C9_N_btm.n554 C9_N_btm.n553 4.60698
R46270 C9_N_btm.n553 C9_N_btm.n552 4.60698
R46271 C9_N_btm.n548 C9_N_btm.n547 4.60698
R46272 C9_N_btm.n547 C9_N_btm.n211 4.60698
R46273 C9_N_btm.n545 C9_N_btm.n544 4.60698
R46274 C9_N_btm.n546 C9_N_btm.n545 4.60698
R46275 C9_N_btm.n542 C9_N_btm.n541 4.60698
R46276 C9_N_btm.n543 C9_N_btm.n542 4.60698
R46277 C9_N_btm.n539 C9_N_btm.n538 4.60698
R46278 C9_N_btm.n540 C9_N_btm.n539 4.60698
R46279 C9_N_btm.n533 C9_N_btm.n532 4.60698
R46280 C9_N_btm.n532 C9_N_btm.n531 4.60698
R46281 C9_N_btm.n530 C9_N_btm.n529 4.60698
R46282 C9_N_btm.n529 C9_N_btm.n528 4.60698
R46283 C9_N_btm.n527 C9_N_btm.n526 4.60698
R46284 C9_N_btm.n526 C9_N_btm.n525 4.60698
R46285 C9_N_btm.n524 C9_N_btm.n523 4.60698
R46286 C9_N_btm.n523 C9_N_btm.n522 4.60698
R46287 C9_N_btm.n514 C9_N_btm.n513 4.60698
R46288 C9_N_btm.n515 C9_N_btm.n514 4.60698
R46289 C9_N_btm.n511 C9_N_btm.n510 4.60698
R46290 C9_N_btm.n512 C9_N_btm.n511 4.60698
R46291 C9_N_btm.n508 C9_N_btm.n507 4.60698
R46292 C9_N_btm.n509 C9_N_btm.n508 4.60698
R46293 C9_N_btm.n505 C9_N_btm.n504 4.60698
R46294 C9_N_btm.n506 C9_N_btm.n505 4.60698
R46295 C9_N_btm.n500 C9_N_btm.n499 4.60698
R46296 C9_N_btm.n499 C9_N_btm.n224 4.60698
R46297 C9_N_btm.n233 C9_N_btm.n232 4.60698
R46298 C9_N_btm.n234 C9_N_btm.n233 4.60698
R46299 C9_N_btm.n236 C9_N_btm.n235 4.60698
R46300 C9_N_btm.n237 C9_N_btm.n236 4.60698
R46301 C9_N_btm.n239 C9_N_btm.n238 4.60698
R46302 C9_N_btm.n238 C9_N_btm.n229 4.60698
R46303 C9_N_btm.n485 C9_N_btm.n484 4.60698
R46304 C9_N_btm.n484 C9_N_btm.n483 4.60698
R46305 C9_N_btm.n488 C9_N_btm.n487 4.60698
R46306 C9_N_btm.n487 C9_N_btm.n486 4.60698
R46307 C9_N_btm.n491 C9_N_btm.n490 4.60698
R46308 C9_N_btm.n490 C9_N_btm.n489 4.60698
R46309 C9_N_btm.n494 C9_N_btm.n493 4.60698
R46310 C9_N_btm.n493 C9_N_btm.n492 4.60698
R46311 C9_N_btm.n468 C9_N_btm.n467 4.60698
R46312 C9_N_btm.n469 C9_N_btm.n468 4.60698
R46313 C9_N_btm.n471 C9_N_btm.n470 4.60698
R46314 C9_N_btm.n472 C9_N_btm.n471 4.60698
R46315 C9_N_btm.n474 C9_N_btm.n473 4.60698
R46316 C9_N_btm.n475 C9_N_btm.n474 4.60698
R46317 C9_N_btm.n477 C9_N_btm.n476 4.60698
R46318 C9_N_btm.n478 C9_N_btm.n477 4.60698
R46319 C9_N_btm.n262 C9_N_btm.n261 4.60698
R46320 C9_N_btm.n261 C9_N_btm.n252 4.60698
R46321 C9_N_btm.n259 C9_N_btm.n258 4.60698
R46322 C9_N_btm.n260 C9_N_btm.n259 4.60698
R46323 C9_N_btm.n256 C9_N_btm.n255 4.60698
R46324 C9_N_btm.n257 C9_N_btm.n256 4.60698
R46325 C9_N_btm.n463 C9_N_btm.n462 4.60698
R46326 C9_N_btm.n462 C9_N_btm.n247 4.60698
R46327 C9_N_btm.n457 C9_N_btm.n456 4.60698
R46328 C9_N_btm.n456 C9_N_btm.n455 4.60698
R46329 C9_N_btm.n454 C9_N_btm.n453 4.60698
R46330 C9_N_btm.n453 C9_N_btm.n452 4.60698
R46331 C9_N_btm.n451 C9_N_btm.n450 4.60698
R46332 C9_N_btm.n450 C9_N_btm.n449 4.60698
R46333 C9_N_btm.n448 C9_N_btm.n447 4.60698
R46334 C9_N_btm.n447 C9_N_btm.n446 4.60698
R46335 C9_N_btm.n440 C9_N_btm.n439 4.60698
R46336 C9_N_btm.n441 C9_N_btm.n440 4.60698
R46337 C9_N_btm.n437 C9_N_btm.n436 4.60698
R46338 C9_N_btm.n438 C9_N_btm.n437 4.60698
R46339 C9_N_btm.n434 C9_N_btm.n433 4.60698
R46340 C9_N_btm.n435 C9_N_btm.n434 4.60698
R46341 C9_N_btm.n431 C9_N_btm.n430 4.60698
R46342 C9_N_btm.n432 C9_N_btm.n431 4.60698
R46343 C9_N_btm.n426 C9_N_btm.n425 4.60698
R46344 C9_N_btm.n425 C9_N_btm.n270 4.60698
R46345 C9_N_btm.n279 C9_N_btm.n278 4.60698
R46346 C9_N_btm.n280 C9_N_btm.n279 4.60698
R46347 C9_N_btm.n282 C9_N_btm.n281 4.60698
R46348 C9_N_btm.n283 C9_N_btm.n282 4.60698
R46349 C9_N_btm.n285 C9_N_btm.n284 4.60698
R46350 C9_N_btm.n284 C9_N_btm.n275 4.60698
R46351 C9_N_btm.n411 C9_N_btm.n410 4.60698
R46352 C9_N_btm.n410 C9_N_btm.n409 4.60698
R46353 C9_N_btm.n414 C9_N_btm.n413 4.60698
R46354 C9_N_btm.n413 C9_N_btm.n412 4.60698
R46355 C9_N_btm.n417 C9_N_btm.n416 4.60698
R46356 C9_N_btm.n416 C9_N_btm.n415 4.60698
R46357 C9_N_btm.n420 C9_N_btm.n419 4.60698
R46358 C9_N_btm.n419 C9_N_btm.n418 4.60698
R46359 C9_N_btm.n394 C9_N_btm.n393 4.60698
R46360 C9_N_btm.n395 C9_N_btm.n394 4.60698
R46361 C9_N_btm.n397 C9_N_btm.n396 4.60698
R46362 C9_N_btm.n398 C9_N_btm.n397 4.60698
R46363 C9_N_btm.n400 C9_N_btm.n399 4.60698
R46364 C9_N_btm.n401 C9_N_btm.n400 4.60698
R46365 C9_N_btm.n403 C9_N_btm.n402 4.60698
R46366 C9_N_btm.n404 C9_N_btm.n403 4.60698
R46367 C9_N_btm.n308 C9_N_btm.n307 4.60698
R46368 C9_N_btm.n307 C9_N_btm.n298 4.60698
R46369 C9_N_btm.n305 C9_N_btm.n304 4.60698
R46370 C9_N_btm.n306 C9_N_btm.n305 4.60698
R46371 C9_N_btm.n302 C9_N_btm.n301 4.60698
R46372 C9_N_btm.n303 C9_N_btm.n302 4.60698
R46373 C9_N_btm.n389 C9_N_btm.n388 4.60698
R46374 C9_N_btm.n388 C9_N_btm.n293 4.60698
R46375 C9_N_btm.n383 C9_N_btm.n382 4.60698
R46376 C9_N_btm.n382 C9_N_btm.n381 4.60698
R46377 C9_N_btm.n380 C9_N_btm.n379 4.60698
R46378 C9_N_btm.n379 C9_N_btm.n378 4.60698
R46379 C9_N_btm.n377 C9_N_btm.n376 4.60698
R46380 C9_N_btm.n376 C9_N_btm.n375 4.60698
R46381 C9_N_btm.n374 C9_N_btm.n373 4.60698
R46382 C9_N_btm.n373 C9_N_btm.n372 4.60698
R46383 C9_N_btm.n366 C9_N_btm.n365 4.60698
R46384 C9_N_btm.n367 C9_N_btm.n366 4.60698
R46385 C9_N_btm.n363 C9_N_btm.n362 4.60698
R46386 C9_N_btm.n364 C9_N_btm.n363 4.60698
R46387 C9_N_btm.n360 C9_N_btm.n359 4.60698
R46388 C9_N_btm.n361 C9_N_btm.n360 4.60698
R46389 C9_N_btm.n357 C9_N_btm.n356 4.60698
R46390 C9_N_btm.n358 C9_N_btm.n357 4.60698
R46391 C9_N_btm.n352 C9_N_btm.n351 4.60698
R46392 C9_N_btm.n351 C9_N_btm.n316 4.60698
R46393 C9_N_btm.n324 C9_N_btm.n323 4.60698
R46394 C9_N_btm.n325 C9_N_btm.n324 4.60698
R46395 C9_N_btm.n327 C9_N_btm.n326 4.60698
R46396 C9_N_btm.n328 C9_N_btm.n327 4.60698
R46397 C9_N_btm.n330 C9_N_btm.n329 4.60698
R46398 C9_N_btm.n329 C9_N_btm.n320 4.60698
R46399 C9_N_btm.n337 C9_N_btm.n336 4.60698
R46400 C9_N_btm.n336 C9_N_btm.n335 4.60698
R46401 C9_N_btm.n340 C9_N_btm.n339 4.60698
R46402 C9_N_btm.n339 C9_N_btm.n338 4.60698
R46403 C9_N_btm.n343 C9_N_btm.n342 4.60698
R46404 C9_N_btm.n342 C9_N_btm.n341 4.60698
R46405 C9_N_btm.n346 C9_N_btm.n345 4.60698
R46406 C9_N_btm.n345 C9_N_btm.n344 4.60698
R46407 C9_N_btm.n738 C9_N_btm.n737 4.60698
R46408 C9_N_btm.n739 C9_N_btm.n738 4.60698
R46409 C9_N_btm.n735 C9_N_btm.n734 4.60698
R46410 C9_N_btm.n736 C9_N_btm.n735 4.60698
R46411 C9_N_btm.n1886 C9_N_btm.t529 4.03712
R46412 C9_N_btm.n1884 C9_N_btm.t447 3.98193
R46413 C9_N_btm.n1855 C9_N_btm.t271 3.98193
R46414 C9_N_btm.n1804 C9_N_btm.t322 3.98193
R46415 C9_N_btm.n1817 C9_N_btm.t138 3.98193
R46416 C9_N_btm.n1820 C9_N_btm.t191 3.98193
R46417 C9_N_btm.n1802 C9_N_btm.t237 3.98193
R46418 C9_N_btm.n44 C9_N_btm.t51 3.98193
R46419 C9_N_btm.n1768 C9_N_btm.t98 3.98193
R46420 C9_N_btm.n1765 C9_N_btm.t451 3.98193
R46421 C9_N_btm.n67 C9_N_btm.t488 3.98193
R46422 C9_N_btm.n1731 C9_N_btm.t17 3.98193
R46423 C9_N_btm.n1728 C9_N_btm.t370 3.98193
R46424 C9_N_btm.n90 C9_N_btm.t419 3.98193
R46425 C9_N_btm.n1694 C9_N_btm.t245 3.98193
R46426 C9_N_btm.n1691 C9_N_btm.t283 3.98193
R46427 C9_N_btm.n113 C9_N_btm.t335 3.98193
R46428 C9_N_btm.n1657 C9_N_btm.t159 3.98193
R46429 C9_N_btm.n635 C9_N_btm.t223 3.98193
R46430 C9_N_btm.n1511 C9_N_btm.t23 3.98193
R46431 C9_N_btm.n1508 C9_N_btm.t67 3.98193
R46432 C9_N_btm.n880 C9_N_btm.t100 3.98193
R46433 C9_N_btm.n1258 C9_N_btm.t155 3.98193
R46434 C9_N_btm.n841 C9_N_btm.t133 3.98193
R46435 C9_N_btm.n1079 C9_N_btm.t350 3.98193
R46436 C9_N_btm.n1122 C9_N_btm.t193 3.98193
R46437 C9_N_btm.n1256 C9_N_btm.t489 3.98193
R46438 C9_N_btm.n1379 C9_N_btm.t408 3.98193
R46439 C9_N_btm.n1382 C9_N_btm.t224 3.98193
R46440 C9_N_btm.n1387 C9_N_btm.t194 3.98193
R46441 C9_N_btm.n797 C9_N_btm.t492 3.98193
R46442 C9_N_btm.n551 C9_N_btm.t158 3.98193
R46443 C9_N_btm.n518 C9_N_btm.t101 3.98193
R46444 C9_N_btm.n521 C9_N_btm.t282 3.98193
R46445 C9_N_btm.n516 C9_N_btm.t244 3.98193
R46446 C9_N_btm.n228 C9_N_btm.t192 3.98193
R46447 C9_N_btm.n482 C9_N_btm.t369 3.98193
R46448 C9_N_btm.n479 C9_N_btm.t323 3.98193
R46449 C9_N_btm.n251 C9_N_btm.t487 3.98193
R46450 C9_N_btm.n445 C9_N_btm.t450 3.98193
R46451 C9_N_btm.n442 C9_N_btm.t402 3.98193
R46452 C9_N_btm.n274 C9_N_btm.t48 3.98193
R46453 C9_N_btm.n408 C9_N_btm.t361 3.98193
R46454 C9_N_btm.n405 C9_N_btm.t511 3.98193
R46455 C9_N_btm.n297 C9_N_btm.t137 3.98193
R46456 C9_N_btm.n371 C9_N_btm.t85 3.98193
R46457 C9_N_btm.n368 C9_N_btm.t270 3.98193
R46458 C9_N_btm.n319 C9_N_btm.t227 3.98193
R46459 C9_N_btm.n334 C9_N_btm.t397 3.98193
R46460 C9_N_btm.n347 C9_N_btm.t346 3.98193
R46461 C9_N_btm.n350 C9_N_btm.t171 3.98193
R46462 C9_N_btm.n355 C9_N_btm.t215 3.98193
R46463 C9_N_btm.n384 C9_N_btm.t28 3.98193
R46464 C9_N_btm.n387 C9_N_btm.t76 3.98193
R46465 C9_N_btm.n392 C9_N_btm.t127 3.98193
R46466 C9_N_btm.n421 C9_N_btm.t470 3.98193
R46467 C9_N_btm.n424 C9_N_btm.t22 3.98193
R46468 C9_N_btm.n429 C9_N_btm.t349 3.98193
R46469 C9_N_btm.n458 C9_N_btm.t389 3.98193
R46470 C9_N_btm.n461 C9_N_btm.t436 3.98193
R46471 C9_N_btm.n466 C9_N_btm.t260 3.98193
R46472 C9_N_btm.n495 C9_N_btm.t311 3.98193
R46473 C9_N_btm.n498 C9_N_btm.t128 3.98193
R46474 C9_N_btm.n503 C9_N_btm.t183 3.98193
R46475 C9_N_btm.n534 C9_N_btm.t229 3.98193
R46476 C9_N_btm.n537 C9_N_btm.t43 3.98193
R46477 C9_N_btm.n606 C9_N_btm.t309 3.98193
R46478 C9_N_btm.n1632 C9_N_btm.t57 3.98193
R46479 C9_N_btm.n1635 C9_N_btm.t337 3.98193
R46480 C9_N_btm.n1640 C9_N_btm.t80 3.98193
R46481 C9_N_btm.n1670 C9_N_btm.t422 3.98193
R46482 C9_N_btm.n1673 C9_N_btm.t177 3.98193
R46483 C9_N_btm.n1678 C9_N_btm.t491 3.98193
R46484 C9_N_btm.n1707 C9_N_btm.t315 3.98193
R46485 C9_N_btm.n1710 C9_N_btm.t116 3.98193
R46486 C9_N_btm.n1715 C9_N_btm.t391 3.98193
R46487 C9_N_btm.n1744 C9_N_btm.t141 3.98193
R46488 C9_N_btm.n1747 C9_N_btm.t476 3.98193
R46489 C9_N_btm.n1752 C9_N_btm.t286 3.98193
R46490 C9_N_btm.n1781 C9_N_btm.t33 3.98193
R46491 C9_N_btm.n1784 C9_N_btm.t372 3.98193
R46492 C9_N_btm.n1789 C9_N_btm.t252 3.98193
R46493 C9_N_btm.n1833 C9_N_btm.t454 3.98193
R46494 C9_N_btm.n1836 C9_N_btm.t264 3.98193
R46495 C9_N_btm.n1841 C9_N_btm.t263 3.98193
R46496 C9_N_btm.n1868 C9_N_btm.t352 3.98193
R46497 C9_N_btm.n1871 C9_N_btm.t91 3.98193
R46498 C9_N_btm.n11 C9_N_btm.n10 3.91717
R46499 C9_N_btm.n5 C9_N_btm.t6 3.57113
R46500 C9_N_btm.n5 C9_N_btm.t8 3.57113
R46501 C9_N_btm.n3 C9_N_btm.t12 3.57113
R46502 C9_N_btm.n3 C9_N_btm.t5 3.57113
R46503 C9_N_btm.n1 C9_N_btm.t10 3.57113
R46504 C9_N_btm.n1 C9_N_btm.t9 3.57113
R46505 C9_N_btm.n0 C9_N_btm.t11 3.57113
R46506 C9_N_btm.n0 C9_N_btm.t7 3.57113
R46507 C9_N_btm.n7 C9_N_btm.t1 2.4755
R46508 C9_N_btm.n7 C9_N_btm.t2 2.4755
R46509 C9_N_btm.n13 C9_N_btm.t539 2.4755
R46510 C9_N_btm.n13 C9_N_btm.t538 2.4755
R46511 C9_N_btm.n12 C9_N_btm.t537 2.4755
R46512 C9_N_btm.n12 C9_N_btm.t540 2.4755
R46513 C9_N_btm.n8 C9_N_btm.t0 2.4755
R46514 C9_N_btm.n8 C9_N_btm.t3 2.4755
R46515 C9_N_btm.n1882 C9_N_btm.t313 1.67819
R46516 C9_N_btm.n1879 C9_N_btm.t196 1.67819
R46517 C9_N_btm.n1876 C9_N_btm.t357 1.67819
R46518 C9_N_btm.n1873 C9_N_btm.t242 1.67819
R46519 C9_N_btm.n1866 C9_N_btm.t479 1.67819
R46520 C9_N_btm.n1863 C9_N_btm.t72 1.67819
R46521 C9_N_btm.n1860 C9_N_btm.t41 1.67819
R46522 C9_N_btm.n1857 C9_N_btm.t129 1.67819
R46523 C9_N_btm.n1851 C9_N_btm.t185 1.67819
R46524 C9_N_btm.n1849 C9_N_btm.t290 1.67819
R46525 C9_N_btm.n1846 C9_N_btm.t268 1.67819
R46526 C9_N_btm.n1843 C9_N_btm.t157 1.67819
R46527 C9_N_btm.n1837 C9_N_btm.t401 1.67819
R46528 C9_N_btm.n1809 C9_N_btm.t15 1.67819
R46529 C9_N_btm.n1812 C9_N_btm.t413 1.67819
R46530 C9_N_btm.n1815 C9_N_btm.t25 1.67819
R46531 C9_N_btm.n1822 C9_N_btm.t44 1.67819
R46532 C9_N_btm.n1825 C9_N_btm.t458 1.67819
R46533 C9_N_btm.n1828 C9_N_btm.t509 1.67819
R46534 C9_N_btm.n1831 C9_N_btm.t66 1.67819
R46535 C9_N_btm.n1791 C9_N_btm.t261 1.67819
R46536 C9_N_btm.n1794 C9_N_btm.t376 1.67819
R46537 C9_N_btm.n1797 C9_N_btm.t27 1.67819
R46538 C9_N_btm.n1800 C9_N_btm.t89 1.67819
R46539 C9_N_btm.n54 C9_N_btm.t440 1.67819
R46540 C9_N_btm.n52 C9_N_btm.t331 1.67819
R46541 C9_N_btm.n49 C9_N_btm.t94 1.67819
R46542 C9_N_btm.n1785 C9_N_btm.t190 1.67819
R46543 C9_N_btm.n1779 C9_N_btm.t182 1.67819
R46544 C9_N_btm.n1776 C9_N_btm.t293 1.67819
R46545 C9_N_btm.n1773 C9_N_btm.t377 1.67819
R46546 C9_N_btm.n1770 C9_N_btm.t481 1.67819
R46547 C9_N_btm.n1763 C9_N_btm.t316 1.67819
R46548 C9_N_btm.n1760 C9_N_btm.t198 1.67819
R46549 C9_N_btm.n1757 C9_N_btm.t146 1.67819
R46550 C9_N_btm.n1754 C9_N_btm.t430 1.67819
R46551 C9_N_btm.n1748 C9_N_btm.t86 1.67819
R46552 C9_N_btm.n72 C9_N_btm.t211 1.67819
R46553 C9_N_btm.n75 C9_N_btm.t508 1.67819
R46554 C9_N_btm.n77 C9_N_btm.t364 1.67819
R46555 C9_N_btm.n1733 C9_N_btm.t403 1.67819
R46556 C9_N_btm.n1736 C9_N_btm.t296 1.67819
R46557 C9_N_btm.n1739 C9_N_btm.t394 1.67819
R46558 C9_N_btm.n1742 C9_N_btm.t281 1.67819
R46559 C9_N_btm.n1717 C9_N_btm.t379 1.67819
R46560 C9_N_btm.n1720 C9_N_btm.t501 1.67819
R46561 C9_N_btm.n1723 C9_N_btm.t110 1.67819
R46562 C9_N_btm.n1726 C9_N_btm.t230 1.67819
R46563 C9_N_btm.n100 C9_N_btm.t274 1.67819
R46564 C9_N_btm.n98 C9_N_btm.t170 1.67819
R46565 C9_N_btm.n95 C9_N_btm.t319 1.67819
R46566 C9_N_btm.n1711 C9_N_btm.t203 1.67819
R46567 C9_N_btm.n1705 C9_N_btm.t449 1.67819
R46568 C9_N_btm.n1702 C9_N_btm.t38 1.67819
R46569 C9_N_btm.n1699 C9_N_btm.t189 1.67819
R46570 C9_N_btm.n1696 C9_N_btm.t92 1.67819
R46571 C9_N_btm.n1689 C9_N_btm.t142 1.67819
R46572 C9_N_btm.n1686 C9_N_btm.t248 1.67819
R46573 C9_N_btm.n1683 C9_N_btm.t231 1.67819
R46574 C9_N_btm.n1680 C9_N_btm.t114 1.67819
R46575 C9_N_btm.n1674 C9_N_btm.t312 1.67819
R46576 C9_N_btm.n118 C9_N_btm.t426 1.67819
R46577 C9_N_btm.n121 C9_N_btm.t74 1.67819
R46578 C9_N_btm.n123 C9_N_btm.t517 1.67819
R46579 C9_N_btm.n1659 C9_N_btm.t167 1.67819
R46580 C9_N_btm.n1662 C9_N_btm.t429 1.67819
R46581 C9_N_btm.n1665 C9_N_btm.t145 1.67819
R46582 C9_N_btm.n1668 C9_N_btm.t29 1.67819
R46583 C9_N_btm.n1642 C9_N_btm.t228 1.67819
R46584 C9_N_btm.n1645 C9_N_btm.t341 1.67819
R46585 C9_N_btm.n1648 C9_N_btm.t469 1.67819
R46586 C9_N_btm.n1651 C9_N_btm.t119 1.67819
R46587 C9_N_btm.n1653 C9_N_btm.t204 1.67819
R46588 C9_N_btm.n673 C9_N_btm.t31 1.67819
R46589 C9_N_btm.n670 C9_N_btm.t148 1.67819
R46590 C9_N_btm.n667 C9_N_btm.t291 1.67819
R46591 C9_N_btm.n664 C9_N_btm.t356 1.67819
R46592 C9_N_btm.n661 C9_N_btm.t241 1.67819
R46593 C9_N_btm.n658 C9_N_btm.t90 1.67819
R46594 C9_N_btm.n655 C9_N_btm.t214 1.67819
R46595 C9_N_btm.n652 C9_N_btm.t325 1.67819
R46596 C9_N_btm.n649 C9_N_btm.t161 1.67819
R46597 C9_N_btm.n646 C9_N_btm.t304 1.67819
R46598 C9_N_btm.n643 C9_N_btm.t411 1.67819
R46599 C9_N_btm.n640 C9_N_btm.t499 1.67819
R46600 C9_N_btm.n637 C9_N_btm.t383 1.67819
R46601 C9_N_btm.n732 C9_N_btm.t37 1.67819
R46602 C9_N_btm.n729 C9_N_btm.t207 1.67819
R46603 C9_N_btm.n726 C9_N_btm.t61 1.67819
R46604 C9_N_btm.n723 C9_N_btm.t233 1.67819
R46605 C9_N_btm.n720 C9_N_btm.t236 1.67819
R46606 C9_N_btm.n717 C9_N_btm.t496 1.67819
R46607 C9_N_btm.n714 C9_N_btm.t143 1.67819
R46608 C9_N_btm.n711 C9_N_btm.t503 1.67819
R46609 C9_N_btm.n708 C9_N_btm.t441 1.67819
R46610 C9_N_btm.n705 C9_N_btm.t54 1.67819
R46611 C9_N_btm.n702 C9_N_btm.t466 1.67819
R46612 C9_N_btm.n699 C9_N_btm.t105 1.67819
R46613 C9_N_btm.n696 C9_N_btm.t486 1.67819
R46614 C9_N_btm.n693 C9_N_btm.t382 1.67819
R46615 C9_N_btm.n690 C9_N_btm.t24 1.67819
R46616 C9_N_btm.n687 C9_N_btm.t410 1.67819
R46617 C9_N_btm.n684 C9_N_btm.t303 1.67819
R46618 C9_N_btm.n681 C9_N_btm.t247 1.67819
R46619 C9_N_btm.n1636 C9_N_btm.t471 1.67819
R46620 C9_N_btm.n1630 C9_N_btm.t139 1.67819
R46621 C9_N_btm.n1627 C9_N_btm.t255 1.67819
R46622 C9_N_btm.n1624 C9_N_btm.t348 1.67819
R46623 C9_N_btm.n1621 C9_N_btm.t456 1.67819
R46624 C9_N_btm.n1618 C9_N_btm.t68 1.67819
R46625 C9_N_btm.n1615 C9_N_btm.t433 1.67819
R46626 C9_N_btm.n1612 C9_N_btm.t504 1.67819
R46627 C9_N_btm.n1609 C9_N_btm.t162 1.67819
R46628 C9_N_btm.n1606 C9_N_btm.t505 1.67819
R46629 C9_N_btm.n1603 C9_N_btm.t99 1.67819
R46630 C9_N_btm.n1600 C9_N_btm.t482 1.67819
R46631 C9_N_btm.n1597 C9_N_btm.t75 1.67819
R46632 C9_N_btm.n1594 C9_N_btm.t195 1.67819
R46633 C9_N_btm.n1591 C9_N_btm.t49 1.67819
R46634 C9_N_btm.n1588 C9_N_btm.t174 1.67819
R46635 C9_N_btm.n1585 C9_N_btm.t277 1.67819
R46636 C9_N_btm.n1582 C9_N_btm.t107 1.67819
R46637 C9_N_btm.n1579 C9_N_btm.t522 1.67819
R46638 C9_N_btm.n1576 C9_N_btm.t82 1.67819
R46639 C9_N_btm.n1573 C9_N_btm.t201 1.67819
R46640 C9_N_btm.n1570 C9_N_btm.t345 1.67819
R46641 C9_N_btm.n1567 C9_N_btm.t180 1.67819
R46642 C9_N_btm.n1564 C9_N_btm.t285 1.67819
R46643 C9_N_btm.n1561 C9_N_btm.t396 1.67819
R46644 C9_N_btm.n1558 C9_N_btm.t259 1.67819
R46645 C9_N_btm.n1555 C9_N_btm.t374 1.67819
R46646 C9_N_btm.n1552 C9_N_btm.t210 1.67819
R46647 C9_N_btm.n1549 C9_N_btm.t351 1.67819
R46648 C9_N_btm.n1546 C9_N_btm.t459 1.67819
R46649 C9_N_btm.n1543 C9_N_btm.t320 1.67819
R46650 C9_N_btm.n1540 C9_N_btm.t453 1.67819
R46651 C9_N_btm.n1537 C9_N_btm.t39 1.67819
R46652 C9_N_btm.n1534 C9_N_btm.t399 1.67819
R46653 C9_N_btm.n1531 C9_N_btm.t58 1.67819
R46654 C9_N_btm.n1528 C9_N_btm.t130 1.67819
R46655 C9_N_btm.n1525 C9_N_btm.t480 1.67819
R46656 C9_N_btm.n1522 C9_N_btm.t73 1.67819
R46657 C9_N_btm.n1519 C9_N_btm.t461 1.67819
R46658 C9_N_btm.n1516 C9_N_btm.t45 1.67819
R46659 C9_N_btm.n1513 C9_N_btm.t173 1.67819
R46660 C9_N_btm.n1506 C9_N_btm.t217 1.67819
R46661 C9_N_btm.n1503 C9_N_btm.t93 1.67819
R46662 C9_N_btm.n1500 C9_N_btm.t19 1.67819
R46663 C9_N_btm.n1497 C9_N_btm.t123 1.67819
R46664 C9_N_btm.n1494 C9_N_btm.t354 1.67819
R46665 C9_N_btm.n1491 C9_N_btm.t184 1.67819
R46666 C9_N_btm.n1488 C9_N_btm.t35 1.67819
R46667 C9_N_btm.n1485 C9_N_btm.t448 1.67819
R46668 C9_N_btm.n1482 C9_N_btm.t83 1.67819
R46669 C9_N_btm.n1479 C9_N_btm.t490 1.67819
R46670 C9_N_btm.n1476 C9_N_btm.t366 1.67819
R46671 C9_N_btm.n1473 C9_N_btm.t187 1.67819
R46672 C9_N_btm.n1470 C9_N_btm.t390 1.67819
R46673 C9_N_btm.n1467 C9_N_btm.t523 1.67819
R46674 C9_N_btm.n1464 C9_N_btm.t423 1.67819
R46675 C9_N_btm.n1461 C9_N_btm.t310 1.67819
R46676 C9_N_btm.n1458 C9_N_btm.t445 1.67819
R46677 C9_N_btm.n1455 C9_N_btm.t336 1.67819
R46678 C9_N_btm.n1452 C9_N_btm.t226 1.67819
R46679 C9_N_btm.n1449 C9_N_btm.t384 1.67819
R46680 C9_N_btm.n1446 C9_N_btm.t510 1.67819
R46681 C9_N_btm.n1443 C9_N_btm.t132 1.67819
R46682 C9_N_btm.n1440 C9_N_btm.t306 1.67819
R46683 C9_N_btm.n1437 C9_N_btm.t165 1.67819
R46684 C9_N_btm.n1434 C9_N_btm.t328 1.67819
R46685 C9_N_btm.n1431 C9_N_btm.t219 1.67819
R46686 C9_N_btm.n1428 C9_N_btm.t70 1.67819
R46687 C9_N_btm.n1425 C9_N_btm.t251 1.67819
R46688 C9_N_btm.n1422 C9_N_btm.t125 1.67819
R46689 C9_N_btm.n1419 C9_N_btm.t298 1.67819
R46690 C9_N_btm.n1416 C9_N_btm.t153 1.67819
R46691 C9_N_btm.n1413 C9_N_btm.t36 1.67819
R46692 C9_N_btm.n1410 C9_N_btm.t206 1.67819
R46693 C9_N_btm.n1407 C9_N_btm.t60 1.67819
R46694 C9_N_btm.n1404 C9_N_btm.t473 1.67819
R46695 C9_N_btm.n1401 C9_N_btm.t118 1.67819
R46696 C9_N_btm.n1398 C9_N_btm.t495 1.67819
R46697 C9_N_btm.n1395 C9_N_btm.t387 1.67819
R46698 C9_N_btm.n1392 C9_N_btm.t444 1.67819
R46699 C9_N_btm.n1389 C9_N_btm.t334 1.67819
R46700 C9_N_btm.n1383 C9_N_btm.t363 1.67819
R46701 C9_N_btm.n921 C9_N_btm.t467 1.67819
R46702 C9_N_btm.n924 C9_N_btm.t427 1.67819
R46703 C9_N_btm.n927 C9_N_btm.t267 1.67819
R46704 C9_N_btm.n930 C9_N_btm.t156 1.67819
R46705 C9_N_btm.n933 C9_N_btm.t26 1.67819
R46706 C9_N_btm.n936 C9_N_btm.t96 1.67819
R46707 C9_N_btm.n939 C9_N_btm.t288 1.67819
R46708 C9_N_btm.n942 C9_N_btm.t71 1.67819
R46709 C9_N_btm.n945 C9_N_btm.t513 1.67819
R46710 C9_N_btm.n948 C9_N_btm.t42 1.67819
R46711 C9_N_btm.n951 C9_N_btm.t168 1.67819
R46712 C9_N_btm.n954 C9_N_btm.t273 1.67819
R46713 C9_N_btm.n957 C9_N_btm.t102 1.67819
R46714 C9_N_btm.n960 C9_N_btm.t512 1.67819
R46715 C9_N_btm.n963 C9_N_btm.t365 1.67819
R46716 C9_N_btm.n966 C9_N_btm.t521 1.67819
R46717 C9_N_btm.n969 C9_N_btm.t338 1.67819
R46718 C9_N_btm.n972 C9_N_btm.t176 1.67819
R46719 C9_N_btm.n975 C9_N_btm.t280 1.67819
R46720 C9_N_btm.n978 C9_N_btm.t424 1.67819
R46721 C9_N_btm.n981 C9_N_btm.t256 1.67819
R46722 C9_N_btm.n984 C9_N_btm.t371 1.67819
R46723 C9_N_btm.n987 C9_N_btm.t477 1.67819
R46724 C9_N_btm.n990 C9_N_btm.t347 1.67819
R46725 C9_N_btm.n993 C9_N_btm.t455 1.67819
R46726 C9_N_btm.n996 C9_N_btm.t292 1.67819
R46727 C9_N_btm.n999 C9_N_btm.t432 1.67819
R46728 C9_N_btm.n1002 C9_N_btm.t262 1.67819
R46729 C9_N_btm.n1005 C9_N_btm.t393 1.67819
R46730 C9_N_btm.n1008 C9_N_btm.t344 1.67819
R46731 C9_N_btm.n1011 C9_N_btm.t124 1.67819
R46732 C9_N_btm.n1014 C9_N_btm.t478 1.67819
R46733 C9_N_btm.n1017 C9_N_btm.t69 1.67819
R46734 C9_N_btm.n1020 C9_N_btm.t218 1.67819
R46735 C9_N_btm.n1023 C9_N_btm.t40 1.67819
R46736 C9_N_btm.n1026 C9_N_btm.t164 1.67819
R46737 C9_N_btm.n1029 C9_N_btm.t13 1.67819
R46738 C9_N_btm.n1032 C9_N_btm.t131 1.67819
R46739 C9_N_btm.n1034 C9_N_btm.t249 1.67819
R46740 C9_N_btm.n1260 C9_N_btm.t299 1.67819
R46741 C9_N_btm.n1263 C9_N_btm.t186 1.67819
R46742 C9_N_btm.n1266 C9_N_btm.t63 1.67819
R46743 C9_N_btm.n1269 C9_N_btm.t209 1.67819
R46744 C9_N_btm.n1272 C9_N_btm.t84 1.67819
R46745 C9_N_btm.n1275 C9_N_btm.t258 1.67819
R46746 C9_N_btm.n1278 C9_N_btm.t239 1.67819
R46747 C9_N_btm.n1281 C9_N_btm.t405 1.67819
R46748 C9_N_btm.n1284 C9_N_btm.t179 1.67819
R46749 C9_N_btm.n1287 C9_N_btm.t55 1.67819
R46750 C9_N_btm.n1290 C9_N_btm.t442 1.67819
R46751 C9_N_btm.n1293 C9_N_btm.t59 1.67819
R46752 C9_N_btm.n1296 C9_N_btm.t472 1.67819
R46753 C9_N_btm.n1299 C9_N_btm.t339 1.67819
R46754 C9_N_btm.n1302 C9_N_btm.t494 1.67819
R46755 C9_N_btm.n1305 C9_N_btm.t386 1.67819
R46756 C9_N_btm.n1308 C9_N_btm.t483 1.67819
R46757 C9_N_btm.n1311 C9_N_btm.t420 1.67819
R46758 C9_N_btm.n1314 C9_N_btm.t308 1.67819
R46759 C9_N_btm.n1317 C9_N_btm.t465 1.67819
R46760 C9_N_btm.n1320 C9_N_btm.t332 1.67819
R46761 C9_N_btm.n1323 C9_N_btm.t222 1.67819
R46762 C9_N_btm.n1326 C9_N_btm.t381 1.67819
R46763 C9_N_btm.n1329 C9_N_btm.t355 1.67819
R46764 C9_N_btm.n1332 C9_N_btm.t409 1.67819
R46765 C9_N_btm.n1335 C9_N_btm.t301 1.67819
R46766 C9_N_btm.n1338 C9_N_btm.t160 1.67819
R46767 C9_N_btm.n1341 C9_N_btm.t324 1.67819
R46768 C9_N_btm.n1344 C9_N_btm.t212 1.67819
R46769 C9_N_btm.n1347 C9_N_btm.t87 1.67819
R46770 C9_N_btm.n1350 C9_N_btm.t238 1.67819
R46771 C9_N_btm.n1353 C9_N_btm.t246 1.67819
R46772 C9_N_btm.n1356 C9_N_btm.t287 1.67819
R46773 C9_N_btm.n1359 C9_N_btm.t147 1.67819
R46774 C9_N_btm.n1362 C9_N_btm.t30 1.67819
R46775 C9_N_btm.n1365 C9_N_btm.t202 1.67819
R46776 C9_N_btm.n1368 C9_N_btm.t112 1.67819
R46777 C9_N_btm.n1371 C9_N_btm.t468 1.67819
R46778 C9_N_btm.n1374 C9_N_btm.t136 1.67819
R46779 C9_N_btm.n1377 C9_N_btm.t21 1.67819
R46780 C9_N_btm.n1137 C9_N_btm.t272 1.67819
R46781 C9_N_btm.n1140 C9_N_btm.t385 1.67819
R46782 C9_N_btm.n1143 C9_N_btm.t300 1.67819
R46783 C9_N_btm.n1146 C9_N_btm.t407 1.67819
R46784 C9_N_btm.n1149 C9_N_btm.t20 1.67819
R46785 C9_N_btm.n1152 C9_N_btm.t380 1.67819
R46786 C9_N_btm.n1155 C9_N_btm.t485 1.67819
R46787 C9_N_btm.n1158 C9_N_btm.t103 1.67819
R46788 C9_N_btm.n1161 C9_N_btm.t463 1.67819
R46789 C9_N_btm.n1164 C9_N_btm.t52 1.67819
R46790 C9_N_btm.n1167 C9_N_btm.t438 1.67819
R46791 C9_N_btm.n1170 C9_N_btm.t113 1.67819
R46792 C9_N_btm.n1173 C9_N_btm.t140 1.67819
R46793 C9_N_btm.n1176 C9_N_btm.t493 1.67819
R46794 C9_N_btm.n1179 C9_N_btm.t115 1.67819
R46795 C9_N_btm.n1182 C9_N_btm.t232 1.67819
R46796 C9_N_btm.n1185 C9_N_btm.t502 1.67819
R46797 C9_N_btm.n1188 C9_N_btm.t205 1.67819
R46798 C9_N_btm.n1191 C9_N_btm.t34 1.67819
R46799 C9_N_btm.n1194 C9_N_btm.t152 1.67819
R46800 C9_N_btm.n1197 C9_N_btm.t294 1.67819
R46801 C9_N_btm.n1200 C9_N_btm.t122 1.67819
R46802 C9_N_btm.n1203 C9_N_btm.t250 1.67819
R46803 C9_N_btm.n1206 C9_N_btm.t358 1.67819
R46804 C9_N_btm.n1209 C9_N_btm.t216 1.67819
R46805 C9_N_btm.n1212 C9_N_btm.t327 1.67819
R46806 C9_N_btm.n1215 C9_N_btm.t163 1.67819
R46807 C9_N_btm.n1218 C9_N_btm.t305 1.67819
R46808 C9_N_btm.n1081 C9_N_btm.t208 1.67819
R46809 C9_N_btm.n1084 C9_N_btm.t373 1.67819
R46810 C9_N_btm.n1087 C9_N_btm.t257 1.67819
R46811 C9_N_btm.n1090 C9_N_btm.t395 1.67819
R46812 C9_N_btm.n1093 C9_N_btm.t284 1.67819
R46813 C9_N_btm.n1096 C9_N_btm.t178 1.67819
R46814 C9_N_btm.n1099 C9_N_btm.t342 1.67819
R46815 C9_N_btm.n1102 C9_N_btm.t200 1.67819
R46816 C9_N_btm.n1105 C9_N_btm.t81 1.67819
R46817 C9_N_btm.n1108 C9_N_btm.t520 1.67819
R46818 C9_N_btm.n1111 C9_N_btm.t106 1.67819
R46819 C9_N_btm.n1114 C9_N_btm.t276 1.67819
R46820 C9_N_btm.n1117 C9_N_btm.t172 1.67819
R46821 C9_N_btm.n1120 C9_N_btm.t46 1.67819
R46822 C9_N_btm.n1221 C9_N_btm.t415 1.67819
R46823 C9_N_btm.n1224 C9_N_btm.t266 1.67819
R46824 C9_N_btm.n1227 C9_N_btm.t404 1.67819
R46825 C9_N_btm.n1230 C9_N_btm.t515 1.67819
R46826 C9_N_btm.n1233 C9_N_btm.t360 1.67819
R46827 C9_N_btm.n1236 C9_N_btm.t462 1.67819
R46828 C9_N_btm.n1239 C9_N_btm.t77 1.67819
R46829 C9_N_btm.n1242 C9_N_btm.t437 1.67819
R46830 C9_N_btm.n1245 C9_N_btm.t56 1.67819
R46831 C9_N_btm.n1248 C9_N_btm.t417 1.67819
R46832 C9_N_btm.n1251 C9_N_btm.t121 1.67819
R46833 C9_N_btm.n1254 C9_N_btm.t111 1.67819
R46834 C9_N_btm.n795 C9_N_btm.t117 1.67819
R46835 C9_N_btm.n792 C9_N_btm.t254 1.67819
R46836 C9_N_btm.n789 C9_N_btm.t418 1.67819
R46837 C9_N_btm.n786 C9_N_btm.t120 1.67819
R46838 C9_N_btm.n783 C9_N_btm.t439 1.67819
R46839 C9_N_btm.n780 C9_N_btm.t78 1.67819
R46840 C9_N_btm.n777 C9_N_btm.t464 1.67819
R46841 C9_N_btm.n774 C9_N_btm.t362 1.67819
R46842 C9_N_btm.n771 C9_N_btm.t18 1.67819
R46843 C9_N_btm.n768 C9_N_btm.t406 1.67819
R46844 C9_N_btm.n765 C9_N_btm.t269 1.67819
R46845 C9_N_btm.n762 C9_N_btm.t416 1.67819
R46846 C9_N_btm.n759 C9_N_btm.t307 1.67819
R46847 C9_N_btm.n756 C9_N_btm.t166 1.67819
R46848 C9_N_btm.n753 C9_N_btm.t329 1.67819
R46849 C9_N_btm.n750 C9_N_btm.t220 1.67819
R46850 C9_N_btm.n747 C9_N_btm.t359 1.67819
R46851 C9_N_btm.n744 C9_N_btm.t253 1.67819
R46852 C9_N_btm.n741 C9_N_btm.t126 1.67819
R46853 C9_N_btm.n604 C9_N_btm.t421 1.67819
R46854 C9_N_btm.n601 C9_N_btm.t435 1.67819
R46855 C9_N_btm.n598 C9_N_btm.t388 1.67819
R46856 C9_N_btm.n595 C9_N_btm.t497 1.67819
R46857 C9_N_btm.n592 C9_N_btm.t340 1.67819
R46858 C9_N_btm.n589 C9_N_btm.t474 1.67819
R46859 C9_N_btm.n586 C9_N_btm.t62 1.67819
R46860 C9_N_btm.n583 C9_N_btm.t443 1.67819
R46861 C9_N_btm.n580 C9_N_btm.t109 1.67819
R46862 C9_N_btm.n577 C9_N_btm.t181 1.67819
R46863 C9_N_btm.n574 C9_N_btm.t398 1.67819
R46864 C9_N_btm.n571 C9_N_btm.t289 1.67819
R46865 C9_N_btm.n568 C9_N_btm.t524 1.67819
R46866 C9_N_btm.n565 C9_N_btm.t88 1.67819
R46867 C9_N_btm.n562 C9_N_btm.t213 1.67819
R46868 C9_N_btm.n559 C9_N_btm.t516 1.67819
R46869 C9_N_btm.n556 C9_N_btm.t507 1.67819
R46870 C9_N_btm.n553 C9_N_btm.t302 1.67819
R46871 C9_N_btm.n547 C9_N_btm.t514 1.67819
R46872 C9_N_btm.n545 C9_N_btm.t134 1.67819
R46873 C9_N_btm.n542 C9_N_btm.t16 1.67819
R46874 C9_N_btm.n539 C9_N_btm.t169 1.67819
R46875 C9_N_btm.n532 C9_N_btm.t343 1.67819
R46876 C9_N_btm.n529 C9_N_btm.t199 1.67819
R46877 C9_N_btm.n526 C9_N_btm.t317 1.67819
R46878 C9_N_btm.n523 C9_N_btm.t428 1.67819
R46879 C9_N_btm.n514 C9_N_btm.t378 1.67819
R46880 C9_N_btm.n511 C9_N_btm.t265 1.67819
R46881 C9_N_btm.n508 C9_N_btm.t151 1.67819
R46882 C9_N_btm.n505 C9_N_btm.t295 1.67819
R46883 C9_N_btm.n499 C9_N_btm.t500 1.67819
R46884 C9_N_btm.n233 C9_N_btm.t97 1.67819
R46885 C9_N_btm.n236 C9_N_btm.t225 1.67819
R46886 C9_N_btm.n238 C9_N_btm.t333 1.67819
R46887 C9_N_btm.n484 C9_N_btm.t506 1.67819
R46888 C9_N_btm.n487 C9_N_btm.t392 1.67819
R46889 C9_N_btm.n490 C9_N_btm.t279 1.67819
R46890 C9_N_btm.n493 C9_N_btm.t425 1.67819
R46891 C9_N_btm.n468 C9_N_btm.t375 1.67819
R46892 C9_N_btm.n471 C9_N_btm.t235 1.67819
R46893 C9_N_btm.n474 C9_N_btm.t353 1.67819
R46894 C9_N_btm.n477 C9_N_btm.t460 1.67819
R46895 C9_N_btm.n261 C9_N_btm.t108 1.67819
R46896 C9_N_btm.n259 C9_N_btm.t50 1.67819
R46897 C9_N_btm.n256 C9_N_btm.t414 1.67819
R46898 C9_N_btm.n462 C9_N_btm.t53 1.67819
R46899 C9_N_btm.n456 C9_N_btm.t498 1.67819
R46900 C9_N_btm.n453 C9_N_btm.t368 1.67819
R46901 C9_N_btm.n450 C9_N_btm.t475 1.67819
R46902 C9_N_btm.n447 C9_N_btm.t65 1.67819
R46903 C9_N_btm.n440 C9_N_btm.t14 1.67819
R46904 C9_N_btm.n437 C9_N_btm.t434 1.67819
R46905 C9_N_btm.n434 C9_N_btm.t321 1.67819
R46906 C9_N_btm.n431 C9_N_btm.t457 1.67819
R46907 C9_N_btm.n425 C9_N_btm.t104 1.67819
R46908 C9_N_btm.n279 C9_N_btm.t484 1.67819
R46909 C9_N_btm.n282 C9_N_btm.t79 1.67819
R46910 C9_N_btm.n284 C9_N_btm.t197 1.67819
R46911 C9_N_btm.n410 C9_N_btm.t149 1.67819
R46912 C9_N_btm.n413 C9_N_btm.t32 1.67819
R46913 C9_N_btm.n416 C9_N_btm.t446 1.67819
R46914 C9_N_btm.n419 C9_N_btm.t240 1.67819
R46915 C9_N_btm.n394 C9_N_btm.t314 1.67819
R46916 C9_N_btm.n397 C9_N_btm.t95 1.67819
R46917 C9_N_btm.n400 C9_N_btm.t221 1.67819
R46918 C9_N_btm.n403 C9_N_btm.t330 1.67819
R46919 C9_N_btm.n307 C9_N_btm.t278 1.67819
R46920 C9_N_btm.n305 C9_N_btm.t175 1.67819
R46921 C9_N_btm.n302 C9_N_btm.t47 1.67819
R46922 C9_N_btm.n388 C9_N_btm.t519 1.67819
R46923 C9_N_btm.n382 C9_N_btm.t144 1.67819
R46924 C9_N_btm.n379 C9_N_btm.t400 1.67819
R46925 C9_N_btm.n376 C9_N_btm.t243 1.67819
R46926 C9_N_btm.n373 C9_N_btm.t234 1.67819
R46927 C9_N_btm.n366 C9_N_btm.t412 1.67819
R46928 C9_N_btm.n363 C9_N_btm.t150 1.67819
R46929 C9_N_btm.n360 C9_N_btm.t188 1.67819
R46930 C9_N_btm.n357 C9_N_btm.t326 1.67819
R46931 C9_N_btm.n351 C9_N_btm.t275 1.67819
R46932 C9_N_btm.n324 C9_N_btm.t135 1.67819
R46933 C9_N_btm.n327 C9_N_btm.t518 1.67819
R46934 C9_N_btm.n329 C9_N_btm.t367 1.67819
R46935 C9_N_btm.n336 C9_N_btm.t64 1.67819
R46936 C9_N_btm.n339 C9_N_btm.t431 1.67819
R46937 C9_N_btm.n342 C9_N_btm.t318 1.67819
R46938 C9_N_btm.n345 C9_N_btm.t452 1.67819
R46939 C9_N_btm.n738 C9_N_btm.t297 1.67819
R46940 C9_N_btm.n735 C9_N_btm.t154 1.67819
R46941 C9_N_btm.n1123 C9_N_btm.n1122 1.05569
R46942 C9_N_btm.n1079 C9_N_btm.n1050 1.05569
R46943 C9_N_btm.n1257 C9_N_btm.n1256 1.05569
R46944 C9_N_btm.n1380 C9_N_btm.n841 1.05569
R46945 C9_N_btm.n607 C9_N_btm.n606 1.05569
R46946 C9_N_btm.n635 C9_N_btm.n610 1.05569
R46947 C9_N_btm.n22 C9_N_btm.n20 1.0005
R46948 C9_N_btm.n23 C9_N_btm.n19 1.0005
R46949 C9_N_btm.n24 C9_N_btm.n18 1.0005
R46950 C9_N_btm.n1854 C9_N_btm.n17 1.0005
R46951 C9_N_btm.n1854 C9_N_btm.n1853 1.0005
R46952 C9_N_btm.n27 C9_N_btm.n24 1.0005
R46953 C9_N_btm.n28 C9_N_btm.n23 1.0005
R46954 C9_N_btm.n1840 C9_N_btm.n22 1.0005
R46955 C9_N_btm.n1840 C9_N_btm.n1839 1.0005
R46956 C9_N_btm.n1807 C9_N_btm.n28 1.0005
R46957 C9_N_btm.n1806 C9_N_btm.n27 1.0005
R46958 C9_N_btm.n1853 C9_N_btm.n25 1.0005
R46959 C9_N_btm.n34 C9_N_btm.n25 1.0005
R46960 C9_N_btm.n1806 C9_N_btm.n33 1.0005
R46961 C9_N_btm.n1807 C9_N_btm.n32 1.0005
R46962 C9_N_btm.n1839 C9_N_btm.n29 1.0005
R46963 C9_N_btm.n1788 C9_N_btm.n29 1.0005
R46964 C9_N_btm.n38 C9_N_btm.n32 1.0005
R46965 C9_N_btm.n37 C9_N_btm.n33 1.0005
R46966 C9_N_btm.n36 C9_N_btm.n34 1.0005
R46967 C9_N_btm.n56 C9_N_btm.n36 1.0005
R46968 C9_N_btm.n46 C9_N_btm.n37 1.0005
R46969 C9_N_btm.n47 C9_N_btm.n38 1.0005
R46970 C9_N_btm.n1788 C9_N_btm.n1787 1.0005
R46971 C9_N_btm.n1787 C9_N_btm.n39 1.0005
R46972 C9_N_btm.n47 C9_N_btm.n42 1.0005
R46973 C9_N_btm.n46 C9_N_btm.n43 1.0005
R46974 C9_N_btm.n57 C9_N_btm.n56 1.0005
R46975 C9_N_btm.n59 C9_N_btm.n57 1.0005
R46976 C9_N_btm.n60 C9_N_btm.n43 1.0005
R46977 C9_N_btm.n61 C9_N_btm.n42 1.0005
R46978 C9_N_btm.n1751 C9_N_btm.n39 1.0005
R46979 C9_N_btm.n1751 C9_N_btm.n1750 1.0005
R46980 C9_N_btm.n70 C9_N_btm.n61 1.0005
R46981 C9_N_btm.n69 C9_N_btm.n60 1.0005
R46982 C9_N_btm.n79 C9_N_btm.n59 1.0005
R46983 C9_N_btm.n80 C9_N_btm.n79 1.0005
R46984 C9_N_btm.n69 C9_N_btm.n66 1.0005
R46985 C9_N_btm.n70 C9_N_btm.n65 1.0005
R46986 C9_N_btm.n1750 C9_N_btm.n62 1.0005
R46987 C9_N_btm.n1714 C9_N_btm.n62 1.0005
R46988 C9_N_btm.n84 C9_N_btm.n65 1.0005
R46989 C9_N_btm.n83 C9_N_btm.n66 1.0005
R46990 C9_N_btm.n82 C9_N_btm.n80 1.0005
R46991 C9_N_btm.n102 C9_N_btm.n82 1.0005
R46992 C9_N_btm.n92 C9_N_btm.n83 1.0005
R46993 C9_N_btm.n93 C9_N_btm.n84 1.0005
R46994 C9_N_btm.n1714 C9_N_btm.n1713 1.0005
R46995 C9_N_btm.n1713 C9_N_btm.n85 1.0005
R46996 C9_N_btm.n93 C9_N_btm.n88 1.0005
R46997 C9_N_btm.n92 C9_N_btm.n89 1.0005
R46998 C9_N_btm.n103 C9_N_btm.n102 1.0005
R46999 C9_N_btm.n105 C9_N_btm.n103 1.0005
R47000 C9_N_btm.n106 C9_N_btm.n89 1.0005
R47001 C9_N_btm.n107 C9_N_btm.n88 1.0005
R47002 C9_N_btm.n1677 C9_N_btm.n85 1.0005
R47003 C9_N_btm.n1677 C9_N_btm.n1676 1.0005
R47004 C9_N_btm.n116 C9_N_btm.n107 1.0005
R47005 C9_N_btm.n115 C9_N_btm.n106 1.0005
R47006 C9_N_btm.n125 C9_N_btm.n105 1.0005
R47007 C9_N_btm.n126 C9_N_btm.n125 1.0005
R47008 C9_N_btm.n115 C9_N_btm.n112 1.0005
R47009 C9_N_btm.n116 C9_N_btm.n111 1.0005
R47010 C9_N_btm.n1676 C9_N_btm.n108 1.0005
R47011 C9_N_btm.n1639 C9_N_btm.n108 1.0005
R47012 C9_N_btm.n131 C9_N_btm.n111 1.0005
R47013 C9_N_btm.n130 C9_N_btm.n112 1.0005
R47014 C9_N_btm.n129 C9_N_btm.n126 1.0005
R47015 C9_N_btm.n1656 C9_N_btm.n1655 1.0005
R47016 C9_N_btm.n634 C9_N_btm.n611 1.0005
R47017 C9_N_btm.n633 C9_N_btm.n612 1.0005
R47018 C9_N_btm.n632 C9_N_btm.n613 1.0005
R47019 C9_N_btm.n631 C9_N_btm.n614 1.0005
R47020 C9_N_btm.n630 C9_N_btm.n615 1.0005
R47021 C9_N_btm.n629 C9_N_btm.n616 1.0005
R47022 C9_N_btm.n628 C9_N_btm.n617 1.0005
R47023 C9_N_btm.n627 C9_N_btm.n618 1.0005
R47024 C9_N_btm.n626 C9_N_btm.n619 1.0005
R47025 C9_N_btm.n625 C9_N_btm.n620 1.0005
R47026 C9_N_btm.n624 C9_N_btm.n621 1.0005
R47027 C9_N_btm.n623 C9_N_btm.n622 1.0005
R47028 C9_N_btm.n676 C9_N_btm.n675 1.0005
R47029 C9_N_btm.n1655 C9_N_btm.n127 1.0005
R47030 C9_N_btm.n677 C9_N_btm.n129 1.0005
R47031 C9_N_btm.n678 C9_N_btm.n130 1.0005
R47032 C9_N_btm.n679 C9_N_btm.n131 1.0005
R47033 C9_N_btm.n1639 C9_N_btm.n1638 1.0005
R47034 C9_N_btm.n1638 C9_N_btm.n132 1.0005
R47035 C9_N_btm.n679 C9_N_btm.n135 1.0005
R47036 C9_N_btm.n678 C9_N_btm.n136 1.0005
R47037 C9_N_btm.n677 C9_N_btm.n137 1.0005
R47038 C9_N_btm.n138 C9_N_btm.n127 1.0005
R47039 C9_N_btm.n676 C9_N_btm.n139 1.0005
R47040 C9_N_btm.n622 C9_N_btm.n140 1.0005
R47041 C9_N_btm.n621 C9_N_btm.n141 1.0005
R47042 C9_N_btm.n620 C9_N_btm.n142 1.0005
R47043 C9_N_btm.n619 C9_N_btm.n143 1.0005
R47044 C9_N_btm.n618 C9_N_btm.n144 1.0005
R47045 C9_N_btm.n617 C9_N_btm.n145 1.0005
R47046 C9_N_btm.n616 C9_N_btm.n146 1.0005
R47047 C9_N_btm.n615 C9_N_btm.n147 1.0005
R47048 C9_N_btm.n614 C9_N_btm.n148 1.0005
R47049 C9_N_btm.n613 C9_N_btm.n149 1.0005
R47050 C9_N_btm.n612 C9_N_btm.n150 1.0005
R47051 C9_N_btm.n611 C9_N_btm.n151 1.0005
R47052 C9_N_btm.n610 C9_N_btm.n152 1.0005
R47053 C9_N_btm.n800 C9_N_btm.n173 1.0005
R47054 C9_N_btm.n801 C9_N_btm.n172 1.0005
R47055 C9_N_btm.n802 C9_N_btm.n171 1.0005
R47056 C9_N_btm.n803 C9_N_btm.n170 1.0005
R47057 C9_N_btm.n804 C9_N_btm.n169 1.0005
R47058 C9_N_btm.n805 C9_N_btm.n168 1.0005
R47059 C9_N_btm.n806 C9_N_btm.n167 1.0005
R47060 C9_N_btm.n807 C9_N_btm.n166 1.0005
R47061 C9_N_btm.n808 C9_N_btm.n165 1.0005
R47062 C9_N_btm.n809 C9_N_btm.n164 1.0005
R47063 C9_N_btm.n810 C9_N_btm.n163 1.0005
R47064 C9_N_btm.n811 C9_N_btm.n162 1.0005
R47065 C9_N_btm.n812 C9_N_btm.n161 1.0005
R47066 C9_N_btm.n813 C9_N_btm.n160 1.0005
R47067 C9_N_btm.n814 C9_N_btm.n159 1.0005
R47068 C9_N_btm.n815 C9_N_btm.n158 1.0005
R47069 C9_N_btm.n816 C9_N_btm.n157 1.0005
R47070 C9_N_btm.n817 C9_N_btm.n156 1.0005
R47071 C9_N_btm.n818 C9_N_btm.n155 1.0005
R47072 C9_N_btm.n819 C9_N_btm.n154 1.0005
R47073 C9_N_btm.n820 C9_N_btm.n153 1.0005
R47074 C9_N_btm.n821 C9_N_btm.n152 1.0005
R47075 C9_N_btm.n822 C9_N_btm.n151 1.0005
R47076 C9_N_btm.n823 C9_N_btm.n150 1.0005
R47077 C9_N_btm.n824 C9_N_btm.n149 1.0005
R47078 C9_N_btm.n825 C9_N_btm.n148 1.0005
R47079 C9_N_btm.n826 C9_N_btm.n147 1.0005
R47080 C9_N_btm.n827 C9_N_btm.n146 1.0005
R47081 C9_N_btm.n828 C9_N_btm.n145 1.0005
R47082 C9_N_btm.n829 C9_N_btm.n144 1.0005
R47083 C9_N_btm.n830 C9_N_btm.n143 1.0005
R47084 C9_N_btm.n831 C9_N_btm.n142 1.0005
R47085 C9_N_btm.n832 C9_N_btm.n141 1.0005
R47086 C9_N_btm.n833 C9_N_btm.n140 1.0005
R47087 C9_N_btm.n834 C9_N_btm.n139 1.0005
R47088 C9_N_btm.n835 C9_N_btm.n138 1.0005
R47089 C9_N_btm.n836 C9_N_btm.n137 1.0005
R47090 C9_N_btm.n837 C9_N_btm.n136 1.0005
R47091 C9_N_btm.n838 C9_N_btm.n135 1.0005
R47092 C9_N_btm.n1386 C9_N_btm.n132 1.0005
R47093 C9_N_btm.n1386 C9_N_btm.n1385 1.0005
R47094 C9_N_btm.n919 C9_N_btm.n838 1.0005
R47095 C9_N_btm.n918 C9_N_btm.n837 1.0005
R47096 C9_N_btm.n917 C9_N_btm.n836 1.0005
R47097 C9_N_btm.n916 C9_N_btm.n835 1.0005
R47098 C9_N_btm.n915 C9_N_btm.n834 1.0005
R47099 C9_N_btm.n914 C9_N_btm.n833 1.0005
R47100 C9_N_btm.n913 C9_N_btm.n832 1.0005
R47101 C9_N_btm.n912 C9_N_btm.n831 1.0005
R47102 C9_N_btm.n911 C9_N_btm.n830 1.0005
R47103 C9_N_btm.n910 C9_N_btm.n829 1.0005
R47104 C9_N_btm.n909 C9_N_btm.n828 1.0005
R47105 C9_N_btm.n908 C9_N_btm.n827 1.0005
R47106 C9_N_btm.n907 C9_N_btm.n826 1.0005
R47107 C9_N_btm.n906 C9_N_btm.n825 1.0005
R47108 C9_N_btm.n905 C9_N_btm.n824 1.0005
R47109 C9_N_btm.n904 C9_N_btm.n823 1.0005
R47110 C9_N_btm.n903 C9_N_btm.n822 1.0005
R47111 C9_N_btm.n902 C9_N_btm.n821 1.0005
R47112 C9_N_btm.n901 C9_N_btm.n820 1.0005
R47113 C9_N_btm.n900 C9_N_btm.n819 1.0005
R47114 C9_N_btm.n899 C9_N_btm.n818 1.0005
R47115 C9_N_btm.n898 C9_N_btm.n817 1.0005
R47116 C9_N_btm.n897 C9_N_btm.n816 1.0005
R47117 C9_N_btm.n896 C9_N_btm.n815 1.0005
R47118 C9_N_btm.n895 C9_N_btm.n814 1.0005
R47119 C9_N_btm.n894 C9_N_btm.n813 1.0005
R47120 C9_N_btm.n893 C9_N_btm.n812 1.0005
R47121 C9_N_btm.n892 C9_N_btm.n811 1.0005
R47122 C9_N_btm.n891 C9_N_btm.n810 1.0005
R47123 C9_N_btm.n890 C9_N_btm.n809 1.0005
R47124 C9_N_btm.n889 C9_N_btm.n808 1.0005
R47125 C9_N_btm.n888 C9_N_btm.n807 1.0005
R47126 C9_N_btm.n887 C9_N_btm.n806 1.0005
R47127 C9_N_btm.n886 C9_N_btm.n805 1.0005
R47128 C9_N_btm.n885 C9_N_btm.n804 1.0005
R47129 C9_N_btm.n884 C9_N_btm.n803 1.0005
R47130 C9_N_btm.n883 C9_N_btm.n802 1.0005
R47131 C9_N_btm.n882 C9_N_btm.n801 1.0005
R47132 C9_N_btm.n1036 C9_N_btm.n800 1.0005
R47133 C9_N_btm.n1037 C9_N_btm.n1036 1.0005
R47134 C9_N_btm.n882 C9_N_btm.n879 1.0005
R47135 C9_N_btm.n883 C9_N_btm.n878 1.0005
R47136 C9_N_btm.n884 C9_N_btm.n877 1.0005
R47137 C9_N_btm.n885 C9_N_btm.n876 1.0005
R47138 C9_N_btm.n886 C9_N_btm.n875 1.0005
R47139 C9_N_btm.n887 C9_N_btm.n874 1.0005
R47140 C9_N_btm.n888 C9_N_btm.n873 1.0005
R47141 C9_N_btm.n889 C9_N_btm.n872 1.0005
R47142 C9_N_btm.n890 C9_N_btm.n871 1.0005
R47143 C9_N_btm.n891 C9_N_btm.n870 1.0005
R47144 C9_N_btm.n892 C9_N_btm.n869 1.0005
R47145 C9_N_btm.n893 C9_N_btm.n868 1.0005
R47146 C9_N_btm.n894 C9_N_btm.n867 1.0005
R47147 C9_N_btm.n895 C9_N_btm.n866 1.0005
R47148 C9_N_btm.n896 C9_N_btm.n865 1.0005
R47149 C9_N_btm.n897 C9_N_btm.n864 1.0005
R47150 C9_N_btm.n898 C9_N_btm.n863 1.0005
R47151 C9_N_btm.n899 C9_N_btm.n862 1.0005
R47152 C9_N_btm.n900 C9_N_btm.n861 1.0005
R47153 C9_N_btm.n901 C9_N_btm.n860 1.0005
R47154 C9_N_btm.n902 C9_N_btm.n859 1.0005
R47155 C9_N_btm.n903 C9_N_btm.n858 1.0005
R47156 C9_N_btm.n904 C9_N_btm.n857 1.0005
R47157 C9_N_btm.n905 C9_N_btm.n856 1.0005
R47158 C9_N_btm.n906 C9_N_btm.n855 1.0005
R47159 C9_N_btm.n907 C9_N_btm.n854 1.0005
R47160 C9_N_btm.n908 C9_N_btm.n853 1.0005
R47161 C9_N_btm.n909 C9_N_btm.n852 1.0005
R47162 C9_N_btm.n910 C9_N_btm.n851 1.0005
R47163 C9_N_btm.n911 C9_N_btm.n850 1.0005
R47164 C9_N_btm.n912 C9_N_btm.n849 1.0005
R47165 C9_N_btm.n913 C9_N_btm.n848 1.0005
R47166 C9_N_btm.n914 C9_N_btm.n847 1.0005
R47167 C9_N_btm.n915 C9_N_btm.n846 1.0005
R47168 C9_N_btm.n916 C9_N_btm.n845 1.0005
R47169 C9_N_btm.n917 C9_N_btm.n844 1.0005
R47170 C9_N_btm.n918 C9_N_btm.n843 1.0005
R47171 C9_N_btm.n919 C9_N_btm.n842 1.0005
R47172 C9_N_btm.n1385 C9_N_btm.n839 1.0005
R47173 C9_N_btm.n1135 C9_N_btm.n839 1.0005
R47174 C9_N_btm.n1134 C9_N_btm.n842 1.0005
R47175 C9_N_btm.n1133 C9_N_btm.n843 1.0005
R47176 C9_N_btm.n1132 C9_N_btm.n844 1.0005
R47177 C9_N_btm.n1131 C9_N_btm.n845 1.0005
R47178 C9_N_btm.n1130 C9_N_btm.n846 1.0005
R47179 C9_N_btm.n1129 C9_N_btm.n847 1.0005
R47180 C9_N_btm.n1128 C9_N_btm.n848 1.0005
R47181 C9_N_btm.n1127 C9_N_btm.n849 1.0005
R47182 C9_N_btm.n1126 C9_N_btm.n850 1.0005
R47183 C9_N_btm.n1125 C9_N_btm.n851 1.0005
R47184 C9_N_btm.n1124 C9_N_btm.n852 1.0005
R47185 C9_N_btm.n1123 C9_N_btm.n853 1.0005
R47186 C9_N_btm.n1064 C9_N_btm.n854 1.0005
R47187 C9_N_btm.n1063 C9_N_btm.n855 1.0005
R47188 C9_N_btm.n1062 C9_N_btm.n856 1.0005
R47189 C9_N_btm.n1061 C9_N_btm.n857 1.0005
R47190 C9_N_btm.n1060 C9_N_btm.n858 1.0005
R47191 C9_N_btm.n1059 C9_N_btm.n859 1.0005
R47192 C9_N_btm.n1058 C9_N_btm.n860 1.0005
R47193 C9_N_btm.n1057 C9_N_btm.n861 1.0005
R47194 C9_N_btm.n1056 C9_N_btm.n862 1.0005
R47195 C9_N_btm.n1055 C9_N_btm.n863 1.0005
R47196 C9_N_btm.n1054 C9_N_btm.n864 1.0005
R47197 C9_N_btm.n1053 C9_N_btm.n865 1.0005
R47198 C9_N_btm.n1052 C9_N_btm.n866 1.0005
R47199 C9_N_btm.n1051 C9_N_btm.n867 1.0005
R47200 C9_N_btm.n1078 C9_N_btm.n1051 1.0005
R47201 C9_N_btm.n1077 C9_N_btm.n1052 1.0005
R47202 C9_N_btm.n1076 C9_N_btm.n1053 1.0005
R47203 C9_N_btm.n1075 C9_N_btm.n1054 1.0005
R47204 C9_N_btm.n1074 C9_N_btm.n1055 1.0005
R47205 C9_N_btm.n1073 C9_N_btm.n1056 1.0005
R47206 C9_N_btm.n1072 C9_N_btm.n1057 1.0005
R47207 C9_N_btm.n1071 C9_N_btm.n1058 1.0005
R47208 C9_N_btm.n1070 C9_N_btm.n1059 1.0005
R47209 C9_N_btm.n1069 C9_N_btm.n1060 1.0005
R47210 C9_N_btm.n1068 C9_N_btm.n1061 1.0005
R47211 C9_N_btm.n1067 C9_N_btm.n1062 1.0005
R47212 C9_N_btm.n1066 C9_N_btm.n1063 1.0005
R47213 C9_N_btm.n1065 C9_N_btm.n1064 1.0005
R47214 C9_N_btm.n1050 C9_N_btm.n868 1.0005
R47215 C9_N_btm.n1049 C9_N_btm.n869 1.0005
R47216 C9_N_btm.n1048 C9_N_btm.n870 1.0005
R47217 C9_N_btm.n1047 C9_N_btm.n871 1.0005
R47218 C9_N_btm.n1046 C9_N_btm.n872 1.0005
R47219 C9_N_btm.n1045 C9_N_btm.n873 1.0005
R47220 C9_N_btm.n1044 C9_N_btm.n874 1.0005
R47221 C9_N_btm.n1043 C9_N_btm.n875 1.0005
R47222 C9_N_btm.n1042 C9_N_btm.n876 1.0005
R47223 C9_N_btm.n1041 C9_N_btm.n877 1.0005
R47224 C9_N_btm.n1040 C9_N_btm.n878 1.0005
R47225 C9_N_btm.n1039 C9_N_btm.n879 1.0005
R47226 C9_N_btm.n1038 C9_N_btm.n1037 1.0005
R47227 C9_N_btm.n1381 C9_N_btm.n1380 1.0005
R47228 C9_N_btm.n1509 C9_N_btm.n799 1.0005
R47229 C9_N_btm.n1257 C9_N_btm.n799 1.0005
R47230 C9_N_btm.n1633 C9_N_btm.n134 1.0005
R47231 C9_N_btm.n1381 C9_N_btm.n134 1.0005
R47232 C9_N_btm.n175 C9_N_btm.n173 1.0005
R47233 C9_N_btm.n176 C9_N_btm.n172 1.0005
R47234 C9_N_btm.n177 C9_N_btm.n171 1.0005
R47235 C9_N_btm.n178 C9_N_btm.n170 1.0005
R47236 C9_N_btm.n179 C9_N_btm.n169 1.0005
R47237 C9_N_btm.n180 C9_N_btm.n168 1.0005
R47238 C9_N_btm.n181 C9_N_btm.n167 1.0005
R47239 C9_N_btm.n182 C9_N_btm.n166 1.0005
R47240 C9_N_btm.n183 C9_N_btm.n165 1.0005
R47241 C9_N_btm.n184 C9_N_btm.n164 1.0005
R47242 C9_N_btm.n185 C9_N_btm.n163 1.0005
R47243 C9_N_btm.n186 C9_N_btm.n162 1.0005
R47244 C9_N_btm.n187 C9_N_btm.n161 1.0005
R47245 C9_N_btm.n188 C9_N_btm.n160 1.0005
R47246 C9_N_btm.n189 C9_N_btm.n159 1.0005
R47247 C9_N_btm.n190 C9_N_btm.n158 1.0005
R47248 C9_N_btm.n191 C9_N_btm.n157 1.0005
R47249 C9_N_btm.n192 C9_N_btm.n156 1.0005
R47250 C9_N_btm.n193 C9_N_btm.n192 1.0005
R47251 C9_N_btm.n194 C9_N_btm.n191 1.0005
R47252 C9_N_btm.n195 C9_N_btm.n190 1.0005
R47253 C9_N_btm.n196 C9_N_btm.n189 1.0005
R47254 C9_N_btm.n197 C9_N_btm.n188 1.0005
R47255 C9_N_btm.n198 C9_N_btm.n187 1.0005
R47256 C9_N_btm.n199 C9_N_btm.n186 1.0005
R47257 C9_N_btm.n200 C9_N_btm.n185 1.0005
R47258 C9_N_btm.n201 C9_N_btm.n184 1.0005
R47259 C9_N_btm.n202 C9_N_btm.n183 1.0005
R47260 C9_N_btm.n203 C9_N_btm.n182 1.0005
R47261 C9_N_btm.n204 C9_N_btm.n181 1.0005
R47262 C9_N_btm.n205 C9_N_btm.n180 1.0005
R47263 C9_N_btm.n206 C9_N_btm.n179 1.0005
R47264 C9_N_btm.n207 C9_N_btm.n178 1.0005
R47265 C9_N_btm.n208 C9_N_btm.n177 1.0005
R47266 C9_N_btm.n209 C9_N_btm.n176 1.0005
R47267 C9_N_btm.n550 C9_N_btm.n175 1.0005
R47268 C9_N_btm.n550 C9_N_btm.n549 1.0005
R47269 C9_N_btm.n212 C9_N_btm.n209 1.0005
R47270 C9_N_btm.n213 C9_N_btm.n208 1.0005
R47271 C9_N_btm.n214 C9_N_btm.n207 1.0005
R47272 C9_N_btm.n216 C9_N_btm.n214 1.0005
R47273 C9_N_btm.n217 C9_N_btm.n213 1.0005
R47274 C9_N_btm.n218 C9_N_btm.n212 1.0005
R47275 C9_N_btm.n549 C9_N_btm.n210 1.0005
R47276 C9_N_btm.n220 C9_N_btm.n210 1.0005
R47277 C9_N_btm.n221 C9_N_btm.n218 1.0005
R47278 C9_N_btm.n222 C9_N_btm.n217 1.0005
R47279 C9_N_btm.n502 C9_N_btm.n216 1.0005
R47280 C9_N_btm.n502 C9_N_btm.n501 1.0005
R47281 C9_N_btm.n231 C9_N_btm.n222 1.0005
R47282 C9_N_btm.n230 C9_N_btm.n221 1.0005
R47283 C9_N_btm.n240 C9_N_btm.n220 1.0005
R47284 C9_N_btm.n241 C9_N_btm.n240 1.0005
R47285 C9_N_btm.n230 C9_N_btm.n227 1.0005
R47286 C9_N_btm.n231 C9_N_btm.n226 1.0005
R47287 C9_N_btm.n501 C9_N_btm.n223 1.0005
R47288 C9_N_btm.n465 C9_N_btm.n223 1.0005
R47289 C9_N_btm.n245 C9_N_btm.n226 1.0005
R47290 C9_N_btm.n244 C9_N_btm.n227 1.0005
R47291 C9_N_btm.n243 C9_N_btm.n241 1.0005
R47292 C9_N_btm.n263 C9_N_btm.n243 1.0005
R47293 C9_N_btm.n253 C9_N_btm.n244 1.0005
R47294 C9_N_btm.n254 C9_N_btm.n245 1.0005
R47295 C9_N_btm.n465 C9_N_btm.n464 1.0005
R47296 C9_N_btm.n464 C9_N_btm.n246 1.0005
R47297 C9_N_btm.n254 C9_N_btm.n249 1.0005
R47298 C9_N_btm.n253 C9_N_btm.n250 1.0005
R47299 C9_N_btm.n264 C9_N_btm.n263 1.0005
R47300 C9_N_btm.n266 C9_N_btm.n264 1.0005
R47301 C9_N_btm.n267 C9_N_btm.n250 1.0005
R47302 C9_N_btm.n268 C9_N_btm.n249 1.0005
R47303 C9_N_btm.n428 C9_N_btm.n246 1.0005
R47304 C9_N_btm.n428 C9_N_btm.n427 1.0005
R47305 C9_N_btm.n277 C9_N_btm.n268 1.0005
R47306 C9_N_btm.n276 C9_N_btm.n267 1.0005
R47307 C9_N_btm.n286 C9_N_btm.n266 1.0005
R47308 C9_N_btm.n287 C9_N_btm.n286 1.0005
R47309 C9_N_btm.n276 C9_N_btm.n273 1.0005
R47310 C9_N_btm.n277 C9_N_btm.n272 1.0005
R47311 C9_N_btm.n427 C9_N_btm.n269 1.0005
R47312 C9_N_btm.n391 C9_N_btm.n269 1.0005
R47313 C9_N_btm.n291 C9_N_btm.n272 1.0005
R47314 C9_N_btm.n290 C9_N_btm.n273 1.0005
R47315 C9_N_btm.n289 C9_N_btm.n287 1.0005
R47316 C9_N_btm.n309 C9_N_btm.n289 1.0005
R47317 C9_N_btm.n299 C9_N_btm.n290 1.0005
R47318 C9_N_btm.n300 C9_N_btm.n291 1.0005
R47319 C9_N_btm.n391 C9_N_btm.n390 1.0005
R47320 C9_N_btm.n390 C9_N_btm.n292 1.0005
R47321 C9_N_btm.n300 C9_N_btm.n295 1.0005
R47322 C9_N_btm.n299 C9_N_btm.n296 1.0005
R47323 C9_N_btm.n310 C9_N_btm.n309 1.0005
R47324 C9_N_btm.n312 C9_N_btm.n310 1.0005
R47325 C9_N_btm.n313 C9_N_btm.n296 1.0005
R47326 C9_N_btm.n314 C9_N_btm.n295 1.0005
R47327 C9_N_btm.n354 C9_N_btm.n292 1.0005
R47328 C9_N_btm.n354 C9_N_btm.n353 1.0005
R47329 C9_N_btm.n322 C9_N_btm.n314 1.0005
R47330 C9_N_btm.n321 C9_N_btm.n313 1.0005
R47331 C9_N_btm.n331 C9_N_btm.n312 1.0005
R47332 C9_N_btm.n332 C9_N_btm.n331 1.0005
R47333 C9_N_btm.n321 C9_N_btm.n318 1.0005
R47334 C9_N_btm.n322 C9_N_btm.n317 1.0005
R47335 C9_N_btm.n353 C9_N_btm.n315 1.0005
R47336 C9_N_btm.n349 C9_N_btm.n348 1.0005
R47337 C9_N_btm.n333 C9_N_btm.n311 1.0005
R47338 C9_N_btm.n369 C9_N_btm.n311 1.0005
R47339 C9_N_btm.n349 C9_N_btm.n294 1.0005
R47340 C9_N_btm.n385 C9_N_btm.n294 1.0005
R47341 C9_N_btm.n370 C9_N_btm.n369 1.0005
R47342 C9_N_btm.n370 C9_N_btm.n288 1.0005
R47343 C9_N_btm.n386 C9_N_btm.n385 1.0005
R47344 C9_N_btm.n386 C9_N_btm.n271 1.0005
R47345 C9_N_btm.n406 C9_N_btm.n288 1.0005
R47346 C9_N_btm.n407 C9_N_btm.n406 1.0005
R47347 C9_N_btm.n422 C9_N_btm.n271 1.0005
R47348 C9_N_btm.n423 C9_N_btm.n422 1.0005
R47349 C9_N_btm.n407 C9_N_btm.n265 1.0005
R47350 C9_N_btm.n443 C9_N_btm.n265 1.0005
R47351 C9_N_btm.n423 C9_N_btm.n248 1.0005
R47352 C9_N_btm.n459 C9_N_btm.n248 1.0005
R47353 C9_N_btm.n444 C9_N_btm.n443 1.0005
R47354 C9_N_btm.n444 C9_N_btm.n242 1.0005
R47355 C9_N_btm.n460 C9_N_btm.n459 1.0005
R47356 C9_N_btm.n460 C9_N_btm.n225 1.0005
R47357 C9_N_btm.n480 C9_N_btm.n242 1.0005
R47358 C9_N_btm.n481 C9_N_btm.n480 1.0005
R47359 C9_N_btm.n496 C9_N_btm.n225 1.0005
R47360 C9_N_btm.n497 C9_N_btm.n496 1.0005
R47361 C9_N_btm.n481 C9_N_btm.n219 1.0005
R47362 C9_N_btm.n517 C9_N_btm.n219 1.0005
R47363 C9_N_btm.n497 C9_N_btm.n215 1.0005
R47364 C9_N_btm.n535 C9_N_btm.n215 1.0005
R47365 C9_N_btm.n520 C9_N_btm.n517 1.0005
R47366 C9_N_btm.n520 C9_N_btm.n519 1.0005
R47367 C9_N_btm.n536 C9_N_btm.n535 1.0005
R47368 C9_N_btm.n536 C9_N_btm.n206 1.0005
R47369 C9_N_btm.n519 C9_N_btm.n174 1.0005
R47370 C9_N_btm.n798 C9_N_btm.n174 1.0005
R47371 C9_N_btm.n607 C9_N_btm.n155 1.0005
R47372 C9_N_btm.n608 C9_N_btm.n154 1.0005
R47373 C9_N_btm.n609 C9_N_btm.n153 1.0005
R47374 C9_N_btm.n1510 C9_N_btm.n798 1.0005
R47375 C9_N_btm.n1510 C9_N_btm.n1509 1.0005
R47376 C9_N_btm.n1634 C9_N_btm.n110 1.0005
R47377 C9_N_btm.n1634 C9_N_btm.n1633 1.0005
R47378 C9_N_btm.n1672 C9_N_btm.n1671 1.0005
R47379 C9_N_btm.n1671 C9_N_btm.n110 1.0005
R47380 C9_N_btm.n1692 C9_N_btm.n104 1.0005
R47381 C9_N_btm.n1656 C9_N_btm.n104 1.0005
R47382 C9_N_btm.n1708 C9_N_btm.n87 1.0005
R47383 C9_N_btm.n1672 C9_N_btm.n87 1.0005
R47384 C9_N_btm.n1693 C9_N_btm.n81 1.0005
R47385 C9_N_btm.n1693 C9_N_btm.n1692 1.0005
R47386 C9_N_btm.n1709 C9_N_btm.n64 1.0005
R47387 C9_N_btm.n1709 C9_N_btm.n1708 1.0005
R47388 C9_N_btm.n1730 C9_N_btm.n1729 1.0005
R47389 C9_N_btm.n1729 C9_N_btm.n81 1.0005
R47390 C9_N_btm.n1746 C9_N_btm.n1745 1.0005
R47391 C9_N_btm.n1745 C9_N_btm.n64 1.0005
R47392 C9_N_btm.n1766 C9_N_btm.n58 1.0005
R47393 C9_N_btm.n1730 C9_N_btm.n58 1.0005
R47394 C9_N_btm.n1782 C9_N_btm.n41 1.0005
R47395 C9_N_btm.n1746 C9_N_btm.n41 1.0005
R47396 C9_N_btm.n1767 C9_N_btm.n35 1.0005
R47397 C9_N_btm.n1767 C9_N_btm.n1766 1.0005
R47398 C9_N_btm.n1783 C9_N_btm.n31 1.0005
R47399 C9_N_btm.n1783 C9_N_btm.n1782 1.0005
R47400 C9_N_btm.n1819 C9_N_btm.n1803 1.0005
R47401 C9_N_btm.n1803 C9_N_btm.n35 1.0005
R47402 C9_N_btm.n1835 C9_N_btm.n1834 1.0005
R47403 C9_N_btm.n1834 C9_N_btm.n31 1.0005
R47404 C9_N_btm.n1818 C9_N_btm.n1805 1.0005
R47405 C9_N_btm.n1819 C9_N_btm.n1818 1.0005
R47406 C9_N_btm.n1869 C9_N_btm.n21 1.0005
R47407 C9_N_btm.n1835 C9_N_btm.n21 1.0005
R47408 C9_N_btm.n1885 C9_N_btm.n16 1.0005
R47409 C9_N_btm.n1805 C9_N_btm.n16 1.0005
R47410 C9_N_btm.n1870 C9_N_btm.n1869 1.0005
R47411 C9_N_btm.n1886 C9_N_btm.n1885 1.0005
R47412 C9_N_btm.n4 C9_N_btm.n2 0.688
R47413 C9_N_btm.n1122 C9_N_btm.n1121 0.679419
R47414 C9_N_btm.n1080 C9_N_btm.n1079 0.679419
R47415 C9_N_btm.n1256 C9_N_btm.n1255 0.679419
R47416 C9_N_btm.n1136 C9_N_btm.n841 0.679419
R47417 C9_N_btm.n1379 C9_N_btm.n1378 0.679419
R47418 C9_N_btm.n1259 C9_N_btm.n1258 0.679419
R47419 C9_N_btm.n881 C9_N_btm.n880 0.679419
R47420 C9_N_btm.n1384 C9_N_btm.n1382 0.679419
R47421 C9_N_btm.n1388 C9_N_btm.n1387 0.679419
R47422 C9_N_btm.n1508 C9_N_btm.n1507 0.679419
R47423 C9_N_btm.n347 C9_N_btm.n346 0.679419
R47424 C9_N_btm.n335 C9_N_btm.n334 0.679419
R47425 C9_N_btm.n320 C9_N_btm.n319 0.679419
R47426 C9_N_btm.n352 C9_N_btm.n350 0.679419
R47427 C9_N_btm.n356 C9_N_btm.n355 0.679419
R47428 C9_N_btm.n368 C9_N_btm.n367 0.679419
R47429 C9_N_btm.n372 C9_N_btm.n371 0.679419
R47430 C9_N_btm.n384 C9_N_btm.n383 0.679419
R47431 C9_N_btm.n389 C9_N_btm.n387 0.679419
R47432 C9_N_btm.n298 C9_N_btm.n297 0.679419
R47433 C9_N_btm.n405 C9_N_btm.n404 0.679419
R47434 C9_N_btm.n393 C9_N_btm.n392 0.679419
R47435 C9_N_btm.n421 C9_N_btm.n420 0.679419
R47436 C9_N_btm.n409 C9_N_btm.n408 0.679419
R47437 C9_N_btm.n275 C9_N_btm.n274 0.679419
R47438 C9_N_btm.n426 C9_N_btm.n424 0.679419
R47439 C9_N_btm.n430 C9_N_btm.n429 0.679419
R47440 C9_N_btm.n442 C9_N_btm.n441 0.679419
R47441 C9_N_btm.n446 C9_N_btm.n445 0.679419
R47442 C9_N_btm.n458 C9_N_btm.n457 0.679419
R47443 C9_N_btm.n463 C9_N_btm.n461 0.679419
R47444 C9_N_btm.n252 C9_N_btm.n251 0.679419
R47445 C9_N_btm.n479 C9_N_btm.n478 0.679419
R47446 C9_N_btm.n467 C9_N_btm.n466 0.679419
R47447 C9_N_btm.n495 C9_N_btm.n494 0.679419
R47448 C9_N_btm.n483 C9_N_btm.n482 0.679419
R47449 C9_N_btm.n229 C9_N_btm.n228 0.679419
R47450 C9_N_btm.n500 C9_N_btm.n498 0.679419
R47451 C9_N_btm.n504 C9_N_btm.n503 0.679419
R47452 C9_N_btm.n516 C9_N_btm.n515 0.679419
R47453 C9_N_btm.n522 C9_N_btm.n521 0.679419
R47454 C9_N_btm.n534 C9_N_btm.n533 0.679419
R47455 C9_N_btm.n538 C9_N_btm.n537 0.679419
R47456 C9_N_btm.n518 C9_N_btm.n211 0.679419
R47457 C9_N_btm.n552 C9_N_btm.n551 0.679419
R47458 C9_N_btm.n606 C9_N_btm.n605 0.679419
R47459 C9_N_btm.n797 C9_N_btm.n796 0.679419
R47460 C9_N_btm.n1512 C9_N_btm.n1511 0.679419
R47461 C9_N_btm.n1632 C9_N_btm.n1631 0.679419
R47462 C9_N_btm.n1637 C9_N_btm.n1635 0.679419
R47463 C9_N_btm.n636 C9_N_btm.n635 0.679419
R47464 C9_N_btm.n1641 C9_N_btm.n1640 0.679419
R47465 C9_N_btm.n1670 C9_N_btm.n1669 0.679419
R47466 C9_N_btm.n1658 C9_N_btm.n1657 0.679419
R47467 C9_N_btm.n114 C9_N_btm.n113 0.679419
R47468 C9_N_btm.n1675 C9_N_btm.n1673 0.679419
R47469 C9_N_btm.n1679 C9_N_btm.n1678 0.679419
R47470 C9_N_btm.n1691 C9_N_btm.n1690 0.679419
R47471 C9_N_btm.n1695 C9_N_btm.n1694 0.679419
R47472 C9_N_btm.n1707 C9_N_btm.n1706 0.679419
R47473 C9_N_btm.n1712 C9_N_btm.n1710 0.679419
R47474 C9_N_btm.n91 C9_N_btm.n90 0.679419
R47475 C9_N_btm.n1728 C9_N_btm.n1727 0.679419
R47476 C9_N_btm.n1716 C9_N_btm.n1715 0.679419
R47477 C9_N_btm.n1744 C9_N_btm.n1743 0.679419
R47478 C9_N_btm.n1732 C9_N_btm.n1731 0.679419
R47479 C9_N_btm.n68 C9_N_btm.n67 0.679419
R47480 C9_N_btm.n1749 C9_N_btm.n1747 0.679419
R47481 C9_N_btm.n1753 C9_N_btm.n1752 0.679419
R47482 C9_N_btm.n1765 C9_N_btm.n1764 0.679419
R47483 C9_N_btm.n1769 C9_N_btm.n1768 0.679419
R47484 C9_N_btm.n1781 C9_N_btm.n1780 0.679419
R47485 C9_N_btm.n1786 C9_N_btm.n1784 0.679419
R47486 C9_N_btm.n45 C9_N_btm.n44 0.679419
R47487 C9_N_btm.n1802 C9_N_btm.n1801 0.679419
R47488 C9_N_btm.n1790 C9_N_btm.n1789 0.679419
R47489 C9_N_btm.n1833 C9_N_btm.n1832 0.679419
R47490 C9_N_btm.n1821 C9_N_btm.n1820 0.679419
R47491 C9_N_btm.n1817 C9_N_btm.n1816 0.679419
R47492 C9_N_btm.n1838 C9_N_btm.n1836 0.679419
R47493 C9_N_btm.n1842 C9_N_btm.n1841 0.679419
R47494 C9_N_btm.n1804 C9_N_btm.n26 0.679419
R47495 C9_N_btm.n1856 C9_N_btm.n1855 0.679419
R47496 C9_N_btm.n1868 C9_N_btm.n1867 0.679419
R47497 C9_N_btm.n1872 C9_N_btm.n1871 0.679419
R47498 C9_N_btm.n1884 C9_N_btm.n1883 0.679419
R47499 C9_N_btm.n6 C9_N_btm.n4 0.672375
R47500 C9_N_btm.n1119 C9_N_btm.n1118 0.6255
R47501 C9_N_btm.n1116 C9_N_btm.n1115 0.6255
R47502 C9_N_btm.n1113 C9_N_btm.n1112 0.6255
R47503 C9_N_btm.n1110 C9_N_btm.n1109 0.6255
R47504 C9_N_btm.n1107 C9_N_btm.n1106 0.6255
R47505 C9_N_btm.n1104 C9_N_btm.n1103 0.6255
R47506 C9_N_btm.n1101 C9_N_btm.n1100 0.6255
R47507 C9_N_btm.n1098 C9_N_btm.n1097 0.6255
R47508 C9_N_btm.n1095 C9_N_btm.n1094 0.6255
R47509 C9_N_btm.n1092 C9_N_btm.n1091 0.6255
R47510 C9_N_btm.n1089 C9_N_btm.n1088 0.6255
R47511 C9_N_btm.n1086 C9_N_btm.n1085 0.6255
R47512 C9_N_btm.n1083 C9_N_btm.n1082 0.6255
R47513 C9_N_btm.n1253 C9_N_btm.n1252 0.6255
R47514 C9_N_btm.n1250 C9_N_btm.n1249 0.6255
R47515 C9_N_btm.n1247 C9_N_btm.n1246 0.6255
R47516 C9_N_btm.n1244 C9_N_btm.n1243 0.6255
R47517 C9_N_btm.n1241 C9_N_btm.n1240 0.6255
R47518 C9_N_btm.n1238 C9_N_btm.n1237 0.6255
R47519 C9_N_btm.n1235 C9_N_btm.n1234 0.6255
R47520 C9_N_btm.n1232 C9_N_btm.n1231 0.6255
R47521 C9_N_btm.n1229 C9_N_btm.n1228 0.6255
R47522 C9_N_btm.n1226 C9_N_btm.n1225 0.6255
R47523 C9_N_btm.n1223 C9_N_btm.n1222 0.6255
R47524 C9_N_btm.n1220 C9_N_btm.n1219 0.6255
R47525 C9_N_btm.n1217 C9_N_btm.n1216 0.6255
R47526 C9_N_btm.n1214 C9_N_btm.n1213 0.6255
R47527 C9_N_btm.n1211 C9_N_btm.n1210 0.6255
R47528 C9_N_btm.n1208 C9_N_btm.n1207 0.6255
R47529 C9_N_btm.n1205 C9_N_btm.n1204 0.6255
R47530 C9_N_btm.n1202 C9_N_btm.n1201 0.6255
R47531 C9_N_btm.n1199 C9_N_btm.n1198 0.6255
R47532 C9_N_btm.n1196 C9_N_btm.n1195 0.6255
R47533 C9_N_btm.n1193 C9_N_btm.n1192 0.6255
R47534 C9_N_btm.n1190 C9_N_btm.n1189 0.6255
R47535 C9_N_btm.n1187 C9_N_btm.n1186 0.6255
R47536 C9_N_btm.n1184 C9_N_btm.n1183 0.6255
R47537 C9_N_btm.n1181 C9_N_btm.n1180 0.6255
R47538 C9_N_btm.n1178 C9_N_btm.n1177 0.6255
R47539 C9_N_btm.n1175 C9_N_btm.n1174 0.6255
R47540 C9_N_btm.n1172 C9_N_btm.n1171 0.6255
R47541 C9_N_btm.n1169 C9_N_btm.n1168 0.6255
R47542 C9_N_btm.n1166 C9_N_btm.n1165 0.6255
R47543 C9_N_btm.n1163 C9_N_btm.n1162 0.6255
R47544 C9_N_btm.n1160 C9_N_btm.n1159 0.6255
R47545 C9_N_btm.n1157 C9_N_btm.n1156 0.6255
R47546 C9_N_btm.n1154 C9_N_btm.n1153 0.6255
R47547 C9_N_btm.n1151 C9_N_btm.n1150 0.6255
R47548 C9_N_btm.n1148 C9_N_btm.n1147 0.6255
R47549 C9_N_btm.n1145 C9_N_btm.n1144 0.6255
R47550 C9_N_btm.n1142 C9_N_btm.n1141 0.6255
R47551 C9_N_btm.n1139 C9_N_btm.n1138 0.6255
R47552 C9_N_btm.n1376 C9_N_btm.n1375 0.6255
R47553 C9_N_btm.n1373 C9_N_btm.n1372 0.6255
R47554 C9_N_btm.n1370 C9_N_btm.n1369 0.6255
R47555 C9_N_btm.n1367 C9_N_btm.n1366 0.6255
R47556 C9_N_btm.n1364 C9_N_btm.n1363 0.6255
R47557 C9_N_btm.n1361 C9_N_btm.n1360 0.6255
R47558 C9_N_btm.n1358 C9_N_btm.n1357 0.6255
R47559 C9_N_btm.n1355 C9_N_btm.n1354 0.6255
R47560 C9_N_btm.n1352 C9_N_btm.n1351 0.6255
R47561 C9_N_btm.n1349 C9_N_btm.n1348 0.6255
R47562 C9_N_btm.n1346 C9_N_btm.n1345 0.6255
R47563 C9_N_btm.n1343 C9_N_btm.n1342 0.6255
R47564 C9_N_btm.n1340 C9_N_btm.n1339 0.6255
R47565 C9_N_btm.n1337 C9_N_btm.n1336 0.6255
R47566 C9_N_btm.n1334 C9_N_btm.n1333 0.6255
R47567 C9_N_btm.n1331 C9_N_btm.n1330 0.6255
R47568 C9_N_btm.n1328 C9_N_btm.n1327 0.6255
R47569 C9_N_btm.n1325 C9_N_btm.n1324 0.6255
R47570 C9_N_btm.n1322 C9_N_btm.n1321 0.6255
R47571 C9_N_btm.n1319 C9_N_btm.n1318 0.6255
R47572 C9_N_btm.n1316 C9_N_btm.n1315 0.6255
R47573 C9_N_btm.n1313 C9_N_btm.n1312 0.6255
R47574 C9_N_btm.n1310 C9_N_btm.n1309 0.6255
R47575 C9_N_btm.n1307 C9_N_btm.n1306 0.6255
R47576 C9_N_btm.n1304 C9_N_btm.n1303 0.6255
R47577 C9_N_btm.n1301 C9_N_btm.n1300 0.6255
R47578 C9_N_btm.n1298 C9_N_btm.n1297 0.6255
R47579 C9_N_btm.n1295 C9_N_btm.n1294 0.6255
R47580 C9_N_btm.n1292 C9_N_btm.n1291 0.6255
R47581 C9_N_btm.n1289 C9_N_btm.n1288 0.6255
R47582 C9_N_btm.n1286 C9_N_btm.n1285 0.6255
R47583 C9_N_btm.n1283 C9_N_btm.n1282 0.6255
R47584 C9_N_btm.n1280 C9_N_btm.n1279 0.6255
R47585 C9_N_btm.n1277 C9_N_btm.n1276 0.6255
R47586 C9_N_btm.n1274 C9_N_btm.n1273 0.6255
R47587 C9_N_btm.n1271 C9_N_btm.n1270 0.6255
R47588 C9_N_btm.n1268 C9_N_btm.n1267 0.6255
R47589 C9_N_btm.n1265 C9_N_btm.n1264 0.6255
R47590 C9_N_btm.n1262 C9_N_btm.n1261 0.6255
R47591 C9_N_btm.n1035 C9_N_btm.n1033 0.6255
R47592 C9_N_btm.n1031 C9_N_btm.n1030 0.6255
R47593 C9_N_btm.n1028 C9_N_btm.n1027 0.6255
R47594 C9_N_btm.n1025 C9_N_btm.n1024 0.6255
R47595 C9_N_btm.n1022 C9_N_btm.n1021 0.6255
R47596 C9_N_btm.n1019 C9_N_btm.n1018 0.6255
R47597 C9_N_btm.n1016 C9_N_btm.n1015 0.6255
R47598 C9_N_btm.n1013 C9_N_btm.n1012 0.6255
R47599 C9_N_btm.n1010 C9_N_btm.n1009 0.6255
R47600 C9_N_btm.n1007 C9_N_btm.n1006 0.6255
R47601 C9_N_btm.n1004 C9_N_btm.n1003 0.6255
R47602 C9_N_btm.n1001 C9_N_btm.n1000 0.6255
R47603 C9_N_btm.n998 C9_N_btm.n997 0.6255
R47604 C9_N_btm.n995 C9_N_btm.n994 0.6255
R47605 C9_N_btm.n992 C9_N_btm.n991 0.6255
R47606 C9_N_btm.n989 C9_N_btm.n988 0.6255
R47607 C9_N_btm.n986 C9_N_btm.n985 0.6255
R47608 C9_N_btm.n983 C9_N_btm.n982 0.6255
R47609 C9_N_btm.n980 C9_N_btm.n979 0.6255
R47610 C9_N_btm.n977 C9_N_btm.n976 0.6255
R47611 C9_N_btm.n974 C9_N_btm.n973 0.6255
R47612 C9_N_btm.n971 C9_N_btm.n970 0.6255
R47613 C9_N_btm.n968 C9_N_btm.n967 0.6255
R47614 C9_N_btm.n965 C9_N_btm.n964 0.6255
R47615 C9_N_btm.n962 C9_N_btm.n961 0.6255
R47616 C9_N_btm.n959 C9_N_btm.n958 0.6255
R47617 C9_N_btm.n956 C9_N_btm.n955 0.6255
R47618 C9_N_btm.n953 C9_N_btm.n952 0.6255
R47619 C9_N_btm.n950 C9_N_btm.n949 0.6255
R47620 C9_N_btm.n947 C9_N_btm.n946 0.6255
R47621 C9_N_btm.n944 C9_N_btm.n943 0.6255
R47622 C9_N_btm.n941 C9_N_btm.n940 0.6255
R47623 C9_N_btm.n938 C9_N_btm.n937 0.6255
R47624 C9_N_btm.n935 C9_N_btm.n934 0.6255
R47625 C9_N_btm.n932 C9_N_btm.n931 0.6255
R47626 C9_N_btm.n929 C9_N_btm.n928 0.6255
R47627 C9_N_btm.n926 C9_N_btm.n925 0.6255
R47628 C9_N_btm.n923 C9_N_btm.n922 0.6255
R47629 C9_N_btm.n920 C9_N_btm.n840 0.6255
R47630 C9_N_btm.n1391 C9_N_btm.n1390 0.6255
R47631 C9_N_btm.n1394 C9_N_btm.n1393 0.6255
R47632 C9_N_btm.n1397 C9_N_btm.n1396 0.6255
R47633 C9_N_btm.n1400 C9_N_btm.n1399 0.6255
R47634 C9_N_btm.n1403 C9_N_btm.n1402 0.6255
R47635 C9_N_btm.n1406 C9_N_btm.n1405 0.6255
R47636 C9_N_btm.n1409 C9_N_btm.n1408 0.6255
R47637 C9_N_btm.n1412 C9_N_btm.n1411 0.6255
R47638 C9_N_btm.n1415 C9_N_btm.n1414 0.6255
R47639 C9_N_btm.n1418 C9_N_btm.n1417 0.6255
R47640 C9_N_btm.n1421 C9_N_btm.n1420 0.6255
R47641 C9_N_btm.n1424 C9_N_btm.n1423 0.6255
R47642 C9_N_btm.n1427 C9_N_btm.n1426 0.6255
R47643 C9_N_btm.n1430 C9_N_btm.n1429 0.6255
R47644 C9_N_btm.n1433 C9_N_btm.n1432 0.6255
R47645 C9_N_btm.n1436 C9_N_btm.n1435 0.6255
R47646 C9_N_btm.n1439 C9_N_btm.n1438 0.6255
R47647 C9_N_btm.n1442 C9_N_btm.n1441 0.6255
R47648 C9_N_btm.n1445 C9_N_btm.n1444 0.6255
R47649 C9_N_btm.n1448 C9_N_btm.n1447 0.6255
R47650 C9_N_btm.n1451 C9_N_btm.n1450 0.6255
R47651 C9_N_btm.n1454 C9_N_btm.n1453 0.6255
R47652 C9_N_btm.n1457 C9_N_btm.n1456 0.6255
R47653 C9_N_btm.n1460 C9_N_btm.n1459 0.6255
R47654 C9_N_btm.n1463 C9_N_btm.n1462 0.6255
R47655 C9_N_btm.n1466 C9_N_btm.n1465 0.6255
R47656 C9_N_btm.n1469 C9_N_btm.n1468 0.6255
R47657 C9_N_btm.n1472 C9_N_btm.n1471 0.6255
R47658 C9_N_btm.n1475 C9_N_btm.n1474 0.6255
R47659 C9_N_btm.n1478 C9_N_btm.n1477 0.6255
R47660 C9_N_btm.n1481 C9_N_btm.n1480 0.6255
R47661 C9_N_btm.n1484 C9_N_btm.n1483 0.6255
R47662 C9_N_btm.n1487 C9_N_btm.n1486 0.6255
R47663 C9_N_btm.n1490 C9_N_btm.n1489 0.6255
R47664 C9_N_btm.n1493 C9_N_btm.n1492 0.6255
R47665 C9_N_btm.n1496 C9_N_btm.n1495 0.6255
R47666 C9_N_btm.n1499 C9_N_btm.n1498 0.6255
R47667 C9_N_btm.n1502 C9_N_btm.n1501 0.6255
R47668 C9_N_btm.n1505 C9_N_btm.n1504 0.6255
R47669 C9_N_btm.n344 C9_N_btm.n343 0.6255
R47670 C9_N_btm.n341 C9_N_btm.n340 0.6255
R47671 C9_N_btm.n338 C9_N_btm.n337 0.6255
R47672 C9_N_btm.n330 C9_N_btm.n328 0.6255
R47673 C9_N_btm.n326 C9_N_btm.n325 0.6255
R47674 C9_N_btm.n323 C9_N_btm.n316 0.6255
R47675 C9_N_btm.n359 C9_N_btm.n358 0.6255
R47676 C9_N_btm.n362 C9_N_btm.n361 0.6255
R47677 C9_N_btm.n365 C9_N_btm.n364 0.6255
R47678 C9_N_btm.n375 C9_N_btm.n374 0.6255
R47679 C9_N_btm.n378 C9_N_btm.n377 0.6255
R47680 C9_N_btm.n381 C9_N_btm.n380 0.6255
R47681 C9_N_btm.n301 C9_N_btm.n293 0.6255
R47682 C9_N_btm.n304 C9_N_btm.n303 0.6255
R47683 C9_N_btm.n308 C9_N_btm.n306 0.6255
R47684 C9_N_btm.n402 C9_N_btm.n401 0.6255
R47685 C9_N_btm.n399 C9_N_btm.n398 0.6255
R47686 C9_N_btm.n396 C9_N_btm.n395 0.6255
R47687 C9_N_btm.n418 C9_N_btm.n417 0.6255
R47688 C9_N_btm.n415 C9_N_btm.n414 0.6255
R47689 C9_N_btm.n412 C9_N_btm.n411 0.6255
R47690 C9_N_btm.n285 C9_N_btm.n283 0.6255
R47691 C9_N_btm.n281 C9_N_btm.n280 0.6255
R47692 C9_N_btm.n278 C9_N_btm.n270 0.6255
R47693 C9_N_btm.n433 C9_N_btm.n432 0.6255
R47694 C9_N_btm.n436 C9_N_btm.n435 0.6255
R47695 C9_N_btm.n439 C9_N_btm.n438 0.6255
R47696 C9_N_btm.n449 C9_N_btm.n448 0.6255
R47697 C9_N_btm.n452 C9_N_btm.n451 0.6255
R47698 C9_N_btm.n455 C9_N_btm.n454 0.6255
R47699 C9_N_btm.n255 C9_N_btm.n247 0.6255
R47700 C9_N_btm.n258 C9_N_btm.n257 0.6255
R47701 C9_N_btm.n262 C9_N_btm.n260 0.6255
R47702 C9_N_btm.n476 C9_N_btm.n475 0.6255
R47703 C9_N_btm.n473 C9_N_btm.n472 0.6255
R47704 C9_N_btm.n470 C9_N_btm.n469 0.6255
R47705 C9_N_btm.n492 C9_N_btm.n491 0.6255
R47706 C9_N_btm.n489 C9_N_btm.n488 0.6255
R47707 C9_N_btm.n486 C9_N_btm.n485 0.6255
R47708 C9_N_btm.n239 C9_N_btm.n237 0.6255
R47709 C9_N_btm.n235 C9_N_btm.n234 0.6255
R47710 C9_N_btm.n232 C9_N_btm.n224 0.6255
R47711 C9_N_btm.n507 C9_N_btm.n506 0.6255
R47712 C9_N_btm.n510 C9_N_btm.n509 0.6255
R47713 C9_N_btm.n513 C9_N_btm.n512 0.6255
R47714 C9_N_btm.n525 C9_N_btm.n524 0.6255
R47715 C9_N_btm.n528 C9_N_btm.n527 0.6255
R47716 C9_N_btm.n531 C9_N_btm.n530 0.6255
R47717 C9_N_btm.n541 C9_N_btm.n540 0.6255
R47718 C9_N_btm.n544 C9_N_btm.n543 0.6255
R47719 C9_N_btm.n548 C9_N_btm.n546 0.6255
R47720 C9_N_btm.n555 C9_N_btm.n554 0.6255
R47721 C9_N_btm.n558 C9_N_btm.n557 0.6255
R47722 C9_N_btm.n561 C9_N_btm.n560 0.6255
R47723 C9_N_btm.n564 C9_N_btm.n563 0.6255
R47724 C9_N_btm.n567 C9_N_btm.n566 0.6255
R47725 C9_N_btm.n570 C9_N_btm.n569 0.6255
R47726 C9_N_btm.n573 C9_N_btm.n572 0.6255
R47727 C9_N_btm.n576 C9_N_btm.n575 0.6255
R47728 C9_N_btm.n579 C9_N_btm.n578 0.6255
R47729 C9_N_btm.n582 C9_N_btm.n581 0.6255
R47730 C9_N_btm.n585 C9_N_btm.n584 0.6255
R47731 C9_N_btm.n588 C9_N_btm.n587 0.6255
R47732 C9_N_btm.n591 C9_N_btm.n590 0.6255
R47733 C9_N_btm.n594 C9_N_btm.n593 0.6255
R47734 C9_N_btm.n597 C9_N_btm.n596 0.6255
R47735 C9_N_btm.n600 C9_N_btm.n599 0.6255
R47736 C9_N_btm.n603 C9_N_btm.n602 0.6255
R47737 C9_N_btm.n734 C9_N_btm.n733 0.6255
R47738 C9_N_btm.n737 C9_N_btm.n736 0.6255
R47739 C9_N_btm.n740 C9_N_btm.n739 0.6255
R47740 C9_N_btm.n743 C9_N_btm.n742 0.6255
R47741 C9_N_btm.n746 C9_N_btm.n745 0.6255
R47742 C9_N_btm.n749 C9_N_btm.n748 0.6255
R47743 C9_N_btm.n752 C9_N_btm.n751 0.6255
R47744 C9_N_btm.n755 C9_N_btm.n754 0.6255
R47745 C9_N_btm.n758 C9_N_btm.n757 0.6255
R47746 C9_N_btm.n761 C9_N_btm.n760 0.6255
R47747 C9_N_btm.n764 C9_N_btm.n763 0.6255
R47748 C9_N_btm.n767 C9_N_btm.n766 0.6255
R47749 C9_N_btm.n770 C9_N_btm.n769 0.6255
R47750 C9_N_btm.n773 C9_N_btm.n772 0.6255
R47751 C9_N_btm.n776 C9_N_btm.n775 0.6255
R47752 C9_N_btm.n779 C9_N_btm.n778 0.6255
R47753 C9_N_btm.n782 C9_N_btm.n781 0.6255
R47754 C9_N_btm.n785 C9_N_btm.n784 0.6255
R47755 C9_N_btm.n788 C9_N_btm.n787 0.6255
R47756 C9_N_btm.n791 C9_N_btm.n790 0.6255
R47757 C9_N_btm.n794 C9_N_btm.n793 0.6255
R47758 C9_N_btm.n1515 C9_N_btm.n1514 0.6255
R47759 C9_N_btm.n1518 C9_N_btm.n1517 0.6255
R47760 C9_N_btm.n1521 C9_N_btm.n1520 0.6255
R47761 C9_N_btm.n1524 C9_N_btm.n1523 0.6255
R47762 C9_N_btm.n1527 C9_N_btm.n1526 0.6255
R47763 C9_N_btm.n1530 C9_N_btm.n1529 0.6255
R47764 C9_N_btm.n1533 C9_N_btm.n1532 0.6255
R47765 C9_N_btm.n1536 C9_N_btm.n1535 0.6255
R47766 C9_N_btm.n1539 C9_N_btm.n1538 0.6255
R47767 C9_N_btm.n1542 C9_N_btm.n1541 0.6255
R47768 C9_N_btm.n1545 C9_N_btm.n1544 0.6255
R47769 C9_N_btm.n1548 C9_N_btm.n1547 0.6255
R47770 C9_N_btm.n1551 C9_N_btm.n1550 0.6255
R47771 C9_N_btm.n1554 C9_N_btm.n1553 0.6255
R47772 C9_N_btm.n1557 C9_N_btm.n1556 0.6255
R47773 C9_N_btm.n1560 C9_N_btm.n1559 0.6255
R47774 C9_N_btm.n1563 C9_N_btm.n1562 0.6255
R47775 C9_N_btm.n1566 C9_N_btm.n1565 0.6255
R47776 C9_N_btm.n1569 C9_N_btm.n1568 0.6255
R47777 C9_N_btm.n1572 C9_N_btm.n1571 0.6255
R47778 C9_N_btm.n1575 C9_N_btm.n1574 0.6255
R47779 C9_N_btm.n1578 C9_N_btm.n1577 0.6255
R47780 C9_N_btm.n1581 C9_N_btm.n1580 0.6255
R47781 C9_N_btm.n1584 C9_N_btm.n1583 0.6255
R47782 C9_N_btm.n1587 C9_N_btm.n1586 0.6255
R47783 C9_N_btm.n1590 C9_N_btm.n1589 0.6255
R47784 C9_N_btm.n1593 C9_N_btm.n1592 0.6255
R47785 C9_N_btm.n1596 C9_N_btm.n1595 0.6255
R47786 C9_N_btm.n1599 C9_N_btm.n1598 0.6255
R47787 C9_N_btm.n1602 C9_N_btm.n1601 0.6255
R47788 C9_N_btm.n1605 C9_N_btm.n1604 0.6255
R47789 C9_N_btm.n1608 C9_N_btm.n1607 0.6255
R47790 C9_N_btm.n1611 C9_N_btm.n1610 0.6255
R47791 C9_N_btm.n1614 C9_N_btm.n1613 0.6255
R47792 C9_N_btm.n1617 C9_N_btm.n1616 0.6255
R47793 C9_N_btm.n1620 C9_N_btm.n1619 0.6255
R47794 C9_N_btm.n1623 C9_N_btm.n1622 0.6255
R47795 C9_N_btm.n1626 C9_N_btm.n1625 0.6255
R47796 C9_N_btm.n1629 C9_N_btm.n1628 0.6255
R47797 C9_N_btm.n680 C9_N_btm.n133 0.6255
R47798 C9_N_btm.n683 C9_N_btm.n682 0.6255
R47799 C9_N_btm.n686 C9_N_btm.n685 0.6255
R47800 C9_N_btm.n689 C9_N_btm.n688 0.6255
R47801 C9_N_btm.n692 C9_N_btm.n691 0.6255
R47802 C9_N_btm.n695 C9_N_btm.n694 0.6255
R47803 C9_N_btm.n698 C9_N_btm.n697 0.6255
R47804 C9_N_btm.n701 C9_N_btm.n700 0.6255
R47805 C9_N_btm.n704 C9_N_btm.n703 0.6255
R47806 C9_N_btm.n707 C9_N_btm.n706 0.6255
R47807 C9_N_btm.n710 C9_N_btm.n709 0.6255
R47808 C9_N_btm.n713 C9_N_btm.n712 0.6255
R47809 C9_N_btm.n716 C9_N_btm.n715 0.6255
R47810 C9_N_btm.n719 C9_N_btm.n718 0.6255
R47811 C9_N_btm.n722 C9_N_btm.n721 0.6255
R47812 C9_N_btm.n725 C9_N_btm.n724 0.6255
R47813 C9_N_btm.n728 C9_N_btm.n727 0.6255
R47814 C9_N_btm.n731 C9_N_btm.n730 0.6255
R47815 C9_N_btm.n639 C9_N_btm.n638 0.6255
R47816 C9_N_btm.n642 C9_N_btm.n641 0.6255
R47817 C9_N_btm.n645 C9_N_btm.n644 0.6255
R47818 C9_N_btm.n648 C9_N_btm.n647 0.6255
R47819 C9_N_btm.n651 C9_N_btm.n650 0.6255
R47820 C9_N_btm.n654 C9_N_btm.n653 0.6255
R47821 C9_N_btm.n657 C9_N_btm.n656 0.6255
R47822 C9_N_btm.n660 C9_N_btm.n659 0.6255
R47823 C9_N_btm.n663 C9_N_btm.n662 0.6255
R47824 C9_N_btm.n666 C9_N_btm.n665 0.6255
R47825 C9_N_btm.n669 C9_N_btm.n668 0.6255
R47826 C9_N_btm.n672 C9_N_btm.n671 0.6255
R47827 C9_N_btm.n674 C9_N_btm.n128 0.6255
R47828 C9_N_btm.n1654 C9_N_btm.n1652 0.6255
R47829 C9_N_btm.n1650 C9_N_btm.n1649 0.6255
R47830 C9_N_btm.n1647 C9_N_btm.n1646 0.6255
R47831 C9_N_btm.n1644 C9_N_btm.n1643 0.6255
R47832 C9_N_btm.n1667 C9_N_btm.n1666 0.6255
R47833 C9_N_btm.n1664 C9_N_btm.n1663 0.6255
R47834 C9_N_btm.n1661 C9_N_btm.n1660 0.6255
R47835 C9_N_btm.n124 C9_N_btm.n122 0.6255
R47836 C9_N_btm.n120 C9_N_btm.n119 0.6255
R47837 C9_N_btm.n117 C9_N_btm.n109 0.6255
R47838 C9_N_btm.n1682 C9_N_btm.n1681 0.6255
R47839 C9_N_btm.n1685 C9_N_btm.n1684 0.6255
R47840 C9_N_btm.n1688 C9_N_btm.n1687 0.6255
R47841 C9_N_btm.n1698 C9_N_btm.n1697 0.6255
R47842 C9_N_btm.n1701 C9_N_btm.n1700 0.6255
R47843 C9_N_btm.n1704 C9_N_btm.n1703 0.6255
R47844 C9_N_btm.n94 C9_N_btm.n86 0.6255
R47845 C9_N_btm.n97 C9_N_btm.n96 0.6255
R47846 C9_N_btm.n101 C9_N_btm.n99 0.6255
R47847 C9_N_btm.n1725 C9_N_btm.n1724 0.6255
R47848 C9_N_btm.n1722 C9_N_btm.n1721 0.6255
R47849 C9_N_btm.n1719 C9_N_btm.n1718 0.6255
R47850 C9_N_btm.n1741 C9_N_btm.n1740 0.6255
R47851 C9_N_btm.n1738 C9_N_btm.n1737 0.6255
R47852 C9_N_btm.n1735 C9_N_btm.n1734 0.6255
R47853 C9_N_btm.n78 C9_N_btm.n76 0.6255
R47854 C9_N_btm.n74 C9_N_btm.n73 0.6255
R47855 C9_N_btm.n71 C9_N_btm.n63 0.6255
R47856 C9_N_btm.n1756 C9_N_btm.n1755 0.6255
R47857 C9_N_btm.n1759 C9_N_btm.n1758 0.6255
R47858 C9_N_btm.n1762 C9_N_btm.n1761 0.6255
R47859 C9_N_btm.n1772 C9_N_btm.n1771 0.6255
R47860 C9_N_btm.n1775 C9_N_btm.n1774 0.6255
R47861 C9_N_btm.n1778 C9_N_btm.n1777 0.6255
R47862 C9_N_btm.n48 C9_N_btm.n40 0.6255
R47863 C9_N_btm.n51 C9_N_btm.n50 0.6255
R47864 C9_N_btm.n55 C9_N_btm.n53 0.6255
R47865 C9_N_btm.n1799 C9_N_btm.n1798 0.6255
R47866 C9_N_btm.n1796 C9_N_btm.n1795 0.6255
R47867 C9_N_btm.n1793 C9_N_btm.n1792 0.6255
R47868 C9_N_btm.n1830 C9_N_btm.n1829 0.6255
R47869 C9_N_btm.n1827 C9_N_btm.n1826 0.6255
R47870 C9_N_btm.n1824 C9_N_btm.n1823 0.6255
R47871 C9_N_btm.n1814 C9_N_btm.n1813 0.6255
R47872 C9_N_btm.n1811 C9_N_btm.n1810 0.6255
R47873 C9_N_btm.n1808 C9_N_btm.n30 0.6255
R47874 C9_N_btm.n1845 C9_N_btm.n1844 0.6255
R47875 C9_N_btm.n1848 C9_N_btm.n1847 0.6255
R47876 C9_N_btm.n1852 C9_N_btm.n1850 0.6255
R47877 C9_N_btm.n1859 C9_N_btm.n1858 0.6255
R47878 C9_N_btm.n1862 C9_N_btm.n1861 0.6255
R47879 C9_N_btm.n1865 C9_N_btm.n1864 0.6255
R47880 C9_N_btm.n1875 C9_N_btm.n1874 0.6255
R47881 C9_N_btm.n1878 C9_N_btm.n1877 0.6255
R47882 C9_N_btm.n1881 C9_N_btm.n1880 0.6255
R47883 C9_N_btm.n1119 C9_N_btm.n1065 0.109875
R47884 C9_N_btm.n1121 C9_N_btm.n1065 0.109875
R47885 C9_N_btm.n1116 C9_N_btm.n1066 0.109875
R47886 C9_N_btm.n1118 C9_N_btm.n1066 0.109875
R47887 C9_N_btm.n1113 C9_N_btm.n1067 0.109875
R47888 C9_N_btm.n1115 C9_N_btm.n1067 0.109875
R47889 C9_N_btm.n1110 C9_N_btm.n1068 0.109875
R47890 C9_N_btm.n1112 C9_N_btm.n1068 0.109875
R47891 C9_N_btm.n1107 C9_N_btm.n1069 0.109875
R47892 C9_N_btm.n1109 C9_N_btm.n1069 0.109875
R47893 C9_N_btm.n1104 C9_N_btm.n1070 0.109875
R47894 C9_N_btm.n1106 C9_N_btm.n1070 0.109875
R47895 C9_N_btm.n1101 C9_N_btm.n1071 0.109875
R47896 C9_N_btm.n1103 C9_N_btm.n1071 0.109875
R47897 C9_N_btm.n1098 C9_N_btm.n1072 0.109875
R47898 C9_N_btm.n1100 C9_N_btm.n1072 0.109875
R47899 C9_N_btm.n1095 C9_N_btm.n1073 0.109875
R47900 C9_N_btm.n1097 C9_N_btm.n1073 0.109875
R47901 C9_N_btm.n1092 C9_N_btm.n1074 0.109875
R47902 C9_N_btm.n1094 C9_N_btm.n1074 0.109875
R47903 C9_N_btm.n1089 C9_N_btm.n1075 0.109875
R47904 C9_N_btm.n1091 C9_N_btm.n1075 0.109875
R47905 C9_N_btm.n1086 C9_N_btm.n1076 0.109875
R47906 C9_N_btm.n1088 C9_N_btm.n1076 0.109875
R47907 C9_N_btm.n1083 C9_N_btm.n1077 0.109875
R47908 C9_N_btm.n1085 C9_N_btm.n1077 0.109875
R47909 C9_N_btm.n1080 C9_N_btm.n1078 0.109875
R47910 C9_N_btm.n1082 C9_N_btm.n1078 0.109875
R47911 C9_N_btm.n1255 C9_N_btm.n1038 0.109875
R47912 C9_N_btm.n1253 C9_N_btm.n1038 0.109875
R47913 C9_N_btm.n1252 C9_N_btm.n1039 0.109875
R47914 C9_N_btm.n1250 C9_N_btm.n1039 0.109875
R47915 C9_N_btm.n1249 C9_N_btm.n1040 0.109875
R47916 C9_N_btm.n1247 C9_N_btm.n1040 0.109875
R47917 C9_N_btm.n1246 C9_N_btm.n1041 0.109875
R47918 C9_N_btm.n1244 C9_N_btm.n1041 0.109875
R47919 C9_N_btm.n1243 C9_N_btm.n1042 0.109875
R47920 C9_N_btm.n1241 C9_N_btm.n1042 0.109875
R47921 C9_N_btm.n1240 C9_N_btm.n1043 0.109875
R47922 C9_N_btm.n1238 C9_N_btm.n1043 0.109875
R47923 C9_N_btm.n1237 C9_N_btm.n1044 0.109875
R47924 C9_N_btm.n1235 C9_N_btm.n1044 0.109875
R47925 C9_N_btm.n1234 C9_N_btm.n1045 0.109875
R47926 C9_N_btm.n1232 C9_N_btm.n1045 0.109875
R47927 C9_N_btm.n1231 C9_N_btm.n1046 0.109875
R47928 C9_N_btm.n1229 C9_N_btm.n1046 0.109875
R47929 C9_N_btm.n1228 C9_N_btm.n1047 0.109875
R47930 C9_N_btm.n1226 C9_N_btm.n1047 0.109875
R47931 C9_N_btm.n1225 C9_N_btm.n1048 0.109875
R47932 C9_N_btm.n1223 C9_N_btm.n1048 0.109875
R47933 C9_N_btm.n1222 C9_N_btm.n1049 0.109875
R47934 C9_N_btm.n1220 C9_N_btm.n1049 0.109875
R47935 C9_N_btm.n1219 C9_N_btm.n1050 0.109875
R47936 C9_N_btm.n1217 C9_N_btm.n1050 0.109875
R47937 C9_N_btm.n1216 C9_N_btm.n1051 0.109875
R47938 C9_N_btm.n1214 C9_N_btm.n1051 0.109875
R47939 C9_N_btm.n1213 C9_N_btm.n1052 0.109875
R47940 C9_N_btm.n1211 C9_N_btm.n1052 0.109875
R47941 C9_N_btm.n1210 C9_N_btm.n1053 0.109875
R47942 C9_N_btm.n1208 C9_N_btm.n1053 0.109875
R47943 C9_N_btm.n1207 C9_N_btm.n1054 0.109875
R47944 C9_N_btm.n1205 C9_N_btm.n1054 0.109875
R47945 C9_N_btm.n1204 C9_N_btm.n1055 0.109875
R47946 C9_N_btm.n1202 C9_N_btm.n1055 0.109875
R47947 C9_N_btm.n1201 C9_N_btm.n1056 0.109875
R47948 C9_N_btm.n1199 C9_N_btm.n1056 0.109875
R47949 C9_N_btm.n1198 C9_N_btm.n1057 0.109875
R47950 C9_N_btm.n1196 C9_N_btm.n1057 0.109875
R47951 C9_N_btm.n1195 C9_N_btm.n1058 0.109875
R47952 C9_N_btm.n1193 C9_N_btm.n1058 0.109875
R47953 C9_N_btm.n1192 C9_N_btm.n1059 0.109875
R47954 C9_N_btm.n1190 C9_N_btm.n1059 0.109875
R47955 C9_N_btm.n1189 C9_N_btm.n1060 0.109875
R47956 C9_N_btm.n1187 C9_N_btm.n1060 0.109875
R47957 C9_N_btm.n1186 C9_N_btm.n1061 0.109875
R47958 C9_N_btm.n1184 C9_N_btm.n1061 0.109875
R47959 C9_N_btm.n1183 C9_N_btm.n1062 0.109875
R47960 C9_N_btm.n1181 C9_N_btm.n1062 0.109875
R47961 C9_N_btm.n1180 C9_N_btm.n1063 0.109875
R47962 C9_N_btm.n1178 C9_N_btm.n1063 0.109875
R47963 C9_N_btm.n1177 C9_N_btm.n1064 0.109875
R47964 C9_N_btm.n1175 C9_N_btm.n1064 0.109875
R47965 C9_N_btm.n1174 C9_N_btm.n1123 0.109875
R47966 C9_N_btm.n1172 C9_N_btm.n1123 0.109875
R47967 C9_N_btm.n1171 C9_N_btm.n1124 0.109875
R47968 C9_N_btm.n1169 C9_N_btm.n1124 0.109875
R47969 C9_N_btm.n1168 C9_N_btm.n1125 0.109875
R47970 C9_N_btm.n1166 C9_N_btm.n1125 0.109875
R47971 C9_N_btm.n1165 C9_N_btm.n1126 0.109875
R47972 C9_N_btm.n1163 C9_N_btm.n1126 0.109875
R47973 C9_N_btm.n1162 C9_N_btm.n1127 0.109875
R47974 C9_N_btm.n1160 C9_N_btm.n1127 0.109875
R47975 C9_N_btm.n1159 C9_N_btm.n1128 0.109875
R47976 C9_N_btm.n1157 C9_N_btm.n1128 0.109875
R47977 C9_N_btm.n1156 C9_N_btm.n1129 0.109875
R47978 C9_N_btm.n1154 C9_N_btm.n1129 0.109875
R47979 C9_N_btm.n1153 C9_N_btm.n1130 0.109875
R47980 C9_N_btm.n1151 C9_N_btm.n1130 0.109875
R47981 C9_N_btm.n1150 C9_N_btm.n1131 0.109875
R47982 C9_N_btm.n1148 C9_N_btm.n1131 0.109875
R47983 C9_N_btm.n1147 C9_N_btm.n1132 0.109875
R47984 C9_N_btm.n1145 C9_N_btm.n1132 0.109875
R47985 C9_N_btm.n1144 C9_N_btm.n1133 0.109875
R47986 C9_N_btm.n1142 C9_N_btm.n1133 0.109875
R47987 C9_N_btm.n1141 C9_N_btm.n1134 0.109875
R47988 C9_N_btm.n1139 C9_N_btm.n1134 0.109875
R47989 C9_N_btm.n1138 C9_N_btm.n1135 0.109875
R47990 C9_N_btm.n1136 C9_N_btm.n1135 0.109875
R47991 C9_N_btm.n1376 C9_N_btm.n839 0.109875
R47992 C9_N_btm.n1378 C9_N_btm.n839 0.109875
R47993 C9_N_btm.n1373 C9_N_btm.n842 0.109875
R47994 C9_N_btm.n1375 C9_N_btm.n842 0.109875
R47995 C9_N_btm.n1370 C9_N_btm.n843 0.109875
R47996 C9_N_btm.n1372 C9_N_btm.n843 0.109875
R47997 C9_N_btm.n1367 C9_N_btm.n844 0.109875
R47998 C9_N_btm.n1369 C9_N_btm.n844 0.109875
R47999 C9_N_btm.n1364 C9_N_btm.n845 0.109875
R48000 C9_N_btm.n1366 C9_N_btm.n845 0.109875
R48001 C9_N_btm.n1361 C9_N_btm.n846 0.109875
R48002 C9_N_btm.n1363 C9_N_btm.n846 0.109875
R48003 C9_N_btm.n1358 C9_N_btm.n847 0.109875
R48004 C9_N_btm.n1360 C9_N_btm.n847 0.109875
R48005 C9_N_btm.n1355 C9_N_btm.n848 0.109875
R48006 C9_N_btm.n1357 C9_N_btm.n848 0.109875
R48007 C9_N_btm.n1352 C9_N_btm.n849 0.109875
R48008 C9_N_btm.n1354 C9_N_btm.n849 0.109875
R48009 C9_N_btm.n1349 C9_N_btm.n850 0.109875
R48010 C9_N_btm.n1351 C9_N_btm.n850 0.109875
R48011 C9_N_btm.n1346 C9_N_btm.n851 0.109875
R48012 C9_N_btm.n1348 C9_N_btm.n851 0.109875
R48013 C9_N_btm.n1343 C9_N_btm.n852 0.109875
R48014 C9_N_btm.n1345 C9_N_btm.n852 0.109875
R48015 C9_N_btm.n1340 C9_N_btm.n853 0.109875
R48016 C9_N_btm.n1342 C9_N_btm.n853 0.109875
R48017 C9_N_btm.n1337 C9_N_btm.n854 0.109875
R48018 C9_N_btm.n1339 C9_N_btm.n854 0.109875
R48019 C9_N_btm.n1334 C9_N_btm.n855 0.109875
R48020 C9_N_btm.n1336 C9_N_btm.n855 0.109875
R48021 C9_N_btm.n1331 C9_N_btm.n856 0.109875
R48022 C9_N_btm.n1333 C9_N_btm.n856 0.109875
R48023 C9_N_btm.n1328 C9_N_btm.n857 0.109875
R48024 C9_N_btm.n1330 C9_N_btm.n857 0.109875
R48025 C9_N_btm.n1325 C9_N_btm.n858 0.109875
R48026 C9_N_btm.n1327 C9_N_btm.n858 0.109875
R48027 C9_N_btm.n1322 C9_N_btm.n859 0.109875
R48028 C9_N_btm.n1324 C9_N_btm.n859 0.109875
R48029 C9_N_btm.n1319 C9_N_btm.n860 0.109875
R48030 C9_N_btm.n1321 C9_N_btm.n860 0.109875
R48031 C9_N_btm.n1316 C9_N_btm.n861 0.109875
R48032 C9_N_btm.n1318 C9_N_btm.n861 0.109875
R48033 C9_N_btm.n1313 C9_N_btm.n862 0.109875
R48034 C9_N_btm.n1315 C9_N_btm.n862 0.109875
R48035 C9_N_btm.n1310 C9_N_btm.n863 0.109875
R48036 C9_N_btm.n1312 C9_N_btm.n863 0.109875
R48037 C9_N_btm.n1307 C9_N_btm.n864 0.109875
R48038 C9_N_btm.n1309 C9_N_btm.n864 0.109875
R48039 C9_N_btm.n1304 C9_N_btm.n865 0.109875
R48040 C9_N_btm.n1306 C9_N_btm.n865 0.109875
R48041 C9_N_btm.n1301 C9_N_btm.n866 0.109875
R48042 C9_N_btm.n1303 C9_N_btm.n866 0.109875
R48043 C9_N_btm.n1298 C9_N_btm.n867 0.109875
R48044 C9_N_btm.n1300 C9_N_btm.n867 0.109875
R48045 C9_N_btm.n1295 C9_N_btm.n868 0.109875
R48046 C9_N_btm.n1297 C9_N_btm.n868 0.109875
R48047 C9_N_btm.n1292 C9_N_btm.n869 0.109875
R48048 C9_N_btm.n1294 C9_N_btm.n869 0.109875
R48049 C9_N_btm.n1289 C9_N_btm.n870 0.109875
R48050 C9_N_btm.n1291 C9_N_btm.n870 0.109875
R48051 C9_N_btm.n1286 C9_N_btm.n871 0.109875
R48052 C9_N_btm.n1288 C9_N_btm.n871 0.109875
R48053 C9_N_btm.n1283 C9_N_btm.n872 0.109875
R48054 C9_N_btm.n1285 C9_N_btm.n872 0.109875
R48055 C9_N_btm.n1280 C9_N_btm.n873 0.109875
R48056 C9_N_btm.n1282 C9_N_btm.n873 0.109875
R48057 C9_N_btm.n1277 C9_N_btm.n874 0.109875
R48058 C9_N_btm.n1279 C9_N_btm.n874 0.109875
R48059 C9_N_btm.n1274 C9_N_btm.n875 0.109875
R48060 C9_N_btm.n1276 C9_N_btm.n875 0.109875
R48061 C9_N_btm.n1271 C9_N_btm.n876 0.109875
R48062 C9_N_btm.n1273 C9_N_btm.n876 0.109875
R48063 C9_N_btm.n1268 C9_N_btm.n877 0.109875
R48064 C9_N_btm.n1270 C9_N_btm.n877 0.109875
R48065 C9_N_btm.n1265 C9_N_btm.n878 0.109875
R48066 C9_N_btm.n1267 C9_N_btm.n878 0.109875
R48067 C9_N_btm.n1262 C9_N_btm.n879 0.109875
R48068 C9_N_btm.n1264 C9_N_btm.n879 0.109875
R48069 C9_N_btm.n1259 C9_N_btm.n1037 0.109875
R48070 C9_N_btm.n1261 C9_N_btm.n1037 0.109875
R48071 C9_N_btm.n1036 C9_N_btm.n881 0.109875
R48072 C9_N_btm.n1036 C9_N_btm.n1035 0.109875
R48073 C9_N_btm.n1033 C9_N_btm.n882 0.109875
R48074 C9_N_btm.n1031 C9_N_btm.n882 0.109875
R48075 C9_N_btm.n1030 C9_N_btm.n883 0.109875
R48076 C9_N_btm.n1028 C9_N_btm.n883 0.109875
R48077 C9_N_btm.n1027 C9_N_btm.n884 0.109875
R48078 C9_N_btm.n1025 C9_N_btm.n884 0.109875
R48079 C9_N_btm.n1024 C9_N_btm.n885 0.109875
R48080 C9_N_btm.n1022 C9_N_btm.n885 0.109875
R48081 C9_N_btm.n1021 C9_N_btm.n886 0.109875
R48082 C9_N_btm.n1019 C9_N_btm.n886 0.109875
R48083 C9_N_btm.n1018 C9_N_btm.n887 0.109875
R48084 C9_N_btm.n1016 C9_N_btm.n887 0.109875
R48085 C9_N_btm.n1015 C9_N_btm.n888 0.109875
R48086 C9_N_btm.n1013 C9_N_btm.n888 0.109875
R48087 C9_N_btm.n1012 C9_N_btm.n889 0.109875
R48088 C9_N_btm.n1010 C9_N_btm.n889 0.109875
R48089 C9_N_btm.n1009 C9_N_btm.n890 0.109875
R48090 C9_N_btm.n1007 C9_N_btm.n890 0.109875
R48091 C9_N_btm.n1006 C9_N_btm.n891 0.109875
R48092 C9_N_btm.n1004 C9_N_btm.n891 0.109875
R48093 C9_N_btm.n1003 C9_N_btm.n892 0.109875
R48094 C9_N_btm.n1001 C9_N_btm.n892 0.109875
R48095 C9_N_btm.n1000 C9_N_btm.n893 0.109875
R48096 C9_N_btm.n998 C9_N_btm.n893 0.109875
R48097 C9_N_btm.n997 C9_N_btm.n894 0.109875
R48098 C9_N_btm.n995 C9_N_btm.n894 0.109875
R48099 C9_N_btm.n994 C9_N_btm.n895 0.109875
R48100 C9_N_btm.n992 C9_N_btm.n895 0.109875
R48101 C9_N_btm.n991 C9_N_btm.n896 0.109875
R48102 C9_N_btm.n989 C9_N_btm.n896 0.109875
R48103 C9_N_btm.n988 C9_N_btm.n897 0.109875
R48104 C9_N_btm.n986 C9_N_btm.n897 0.109875
R48105 C9_N_btm.n985 C9_N_btm.n898 0.109875
R48106 C9_N_btm.n983 C9_N_btm.n898 0.109875
R48107 C9_N_btm.n982 C9_N_btm.n899 0.109875
R48108 C9_N_btm.n980 C9_N_btm.n899 0.109875
R48109 C9_N_btm.n979 C9_N_btm.n900 0.109875
R48110 C9_N_btm.n977 C9_N_btm.n900 0.109875
R48111 C9_N_btm.n976 C9_N_btm.n901 0.109875
R48112 C9_N_btm.n974 C9_N_btm.n901 0.109875
R48113 C9_N_btm.n973 C9_N_btm.n902 0.109875
R48114 C9_N_btm.n971 C9_N_btm.n902 0.109875
R48115 C9_N_btm.n970 C9_N_btm.n903 0.109875
R48116 C9_N_btm.n968 C9_N_btm.n903 0.109875
R48117 C9_N_btm.n967 C9_N_btm.n904 0.109875
R48118 C9_N_btm.n965 C9_N_btm.n904 0.109875
R48119 C9_N_btm.n964 C9_N_btm.n905 0.109875
R48120 C9_N_btm.n962 C9_N_btm.n905 0.109875
R48121 C9_N_btm.n961 C9_N_btm.n906 0.109875
R48122 C9_N_btm.n959 C9_N_btm.n906 0.109875
R48123 C9_N_btm.n958 C9_N_btm.n907 0.109875
R48124 C9_N_btm.n956 C9_N_btm.n907 0.109875
R48125 C9_N_btm.n955 C9_N_btm.n908 0.109875
R48126 C9_N_btm.n953 C9_N_btm.n908 0.109875
R48127 C9_N_btm.n952 C9_N_btm.n909 0.109875
R48128 C9_N_btm.n950 C9_N_btm.n909 0.109875
R48129 C9_N_btm.n949 C9_N_btm.n910 0.109875
R48130 C9_N_btm.n947 C9_N_btm.n910 0.109875
R48131 C9_N_btm.n946 C9_N_btm.n911 0.109875
R48132 C9_N_btm.n944 C9_N_btm.n911 0.109875
R48133 C9_N_btm.n943 C9_N_btm.n912 0.109875
R48134 C9_N_btm.n941 C9_N_btm.n912 0.109875
R48135 C9_N_btm.n940 C9_N_btm.n913 0.109875
R48136 C9_N_btm.n938 C9_N_btm.n913 0.109875
R48137 C9_N_btm.n937 C9_N_btm.n914 0.109875
R48138 C9_N_btm.n935 C9_N_btm.n914 0.109875
R48139 C9_N_btm.n934 C9_N_btm.n915 0.109875
R48140 C9_N_btm.n932 C9_N_btm.n915 0.109875
R48141 C9_N_btm.n931 C9_N_btm.n916 0.109875
R48142 C9_N_btm.n929 C9_N_btm.n916 0.109875
R48143 C9_N_btm.n928 C9_N_btm.n917 0.109875
R48144 C9_N_btm.n926 C9_N_btm.n917 0.109875
R48145 C9_N_btm.n925 C9_N_btm.n918 0.109875
R48146 C9_N_btm.n923 C9_N_btm.n918 0.109875
R48147 C9_N_btm.n922 C9_N_btm.n919 0.109875
R48148 C9_N_btm.n920 C9_N_btm.n919 0.109875
R48149 C9_N_btm.n1385 C9_N_btm.n840 0.109875
R48150 C9_N_btm.n1385 C9_N_btm.n1384 0.109875
R48151 C9_N_btm.n1390 C9_N_btm.n1386 0.109875
R48152 C9_N_btm.n1388 C9_N_btm.n1386 0.109875
R48153 C9_N_btm.n1393 C9_N_btm.n838 0.109875
R48154 C9_N_btm.n1391 C9_N_btm.n838 0.109875
R48155 C9_N_btm.n1396 C9_N_btm.n837 0.109875
R48156 C9_N_btm.n1394 C9_N_btm.n837 0.109875
R48157 C9_N_btm.n1399 C9_N_btm.n836 0.109875
R48158 C9_N_btm.n1397 C9_N_btm.n836 0.109875
R48159 C9_N_btm.n1402 C9_N_btm.n835 0.109875
R48160 C9_N_btm.n1400 C9_N_btm.n835 0.109875
R48161 C9_N_btm.n1405 C9_N_btm.n834 0.109875
R48162 C9_N_btm.n1403 C9_N_btm.n834 0.109875
R48163 C9_N_btm.n1408 C9_N_btm.n833 0.109875
R48164 C9_N_btm.n1406 C9_N_btm.n833 0.109875
R48165 C9_N_btm.n1411 C9_N_btm.n832 0.109875
R48166 C9_N_btm.n1409 C9_N_btm.n832 0.109875
R48167 C9_N_btm.n1414 C9_N_btm.n831 0.109875
R48168 C9_N_btm.n1412 C9_N_btm.n831 0.109875
R48169 C9_N_btm.n1417 C9_N_btm.n830 0.109875
R48170 C9_N_btm.n1415 C9_N_btm.n830 0.109875
R48171 C9_N_btm.n1420 C9_N_btm.n829 0.109875
R48172 C9_N_btm.n1418 C9_N_btm.n829 0.109875
R48173 C9_N_btm.n1423 C9_N_btm.n828 0.109875
R48174 C9_N_btm.n1421 C9_N_btm.n828 0.109875
R48175 C9_N_btm.n1426 C9_N_btm.n827 0.109875
R48176 C9_N_btm.n1424 C9_N_btm.n827 0.109875
R48177 C9_N_btm.n1429 C9_N_btm.n826 0.109875
R48178 C9_N_btm.n1427 C9_N_btm.n826 0.109875
R48179 C9_N_btm.n1432 C9_N_btm.n825 0.109875
R48180 C9_N_btm.n1430 C9_N_btm.n825 0.109875
R48181 C9_N_btm.n1435 C9_N_btm.n824 0.109875
R48182 C9_N_btm.n1433 C9_N_btm.n824 0.109875
R48183 C9_N_btm.n1438 C9_N_btm.n823 0.109875
R48184 C9_N_btm.n1436 C9_N_btm.n823 0.109875
R48185 C9_N_btm.n1441 C9_N_btm.n822 0.109875
R48186 C9_N_btm.n1439 C9_N_btm.n822 0.109875
R48187 C9_N_btm.n1444 C9_N_btm.n821 0.109875
R48188 C9_N_btm.n1442 C9_N_btm.n821 0.109875
R48189 C9_N_btm.n1447 C9_N_btm.n820 0.109875
R48190 C9_N_btm.n1445 C9_N_btm.n820 0.109875
R48191 C9_N_btm.n1450 C9_N_btm.n819 0.109875
R48192 C9_N_btm.n1448 C9_N_btm.n819 0.109875
R48193 C9_N_btm.n1453 C9_N_btm.n818 0.109875
R48194 C9_N_btm.n1451 C9_N_btm.n818 0.109875
R48195 C9_N_btm.n1456 C9_N_btm.n817 0.109875
R48196 C9_N_btm.n1454 C9_N_btm.n817 0.109875
R48197 C9_N_btm.n1459 C9_N_btm.n816 0.109875
R48198 C9_N_btm.n1457 C9_N_btm.n816 0.109875
R48199 C9_N_btm.n1462 C9_N_btm.n815 0.109875
R48200 C9_N_btm.n1460 C9_N_btm.n815 0.109875
R48201 C9_N_btm.n1465 C9_N_btm.n814 0.109875
R48202 C9_N_btm.n1463 C9_N_btm.n814 0.109875
R48203 C9_N_btm.n1468 C9_N_btm.n813 0.109875
R48204 C9_N_btm.n1466 C9_N_btm.n813 0.109875
R48205 C9_N_btm.n1471 C9_N_btm.n812 0.109875
R48206 C9_N_btm.n1469 C9_N_btm.n812 0.109875
R48207 C9_N_btm.n1474 C9_N_btm.n811 0.109875
R48208 C9_N_btm.n1472 C9_N_btm.n811 0.109875
R48209 C9_N_btm.n1477 C9_N_btm.n810 0.109875
R48210 C9_N_btm.n1475 C9_N_btm.n810 0.109875
R48211 C9_N_btm.n1480 C9_N_btm.n809 0.109875
R48212 C9_N_btm.n1478 C9_N_btm.n809 0.109875
R48213 C9_N_btm.n1483 C9_N_btm.n808 0.109875
R48214 C9_N_btm.n1481 C9_N_btm.n808 0.109875
R48215 C9_N_btm.n1486 C9_N_btm.n807 0.109875
R48216 C9_N_btm.n1484 C9_N_btm.n807 0.109875
R48217 C9_N_btm.n1489 C9_N_btm.n806 0.109875
R48218 C9_N_btm.n1487 C9_N_btm.n806 0.109875
R48219 C9_N_btm.n1492 C9_N_btm.n805 0.109875
R48220 C9_N_btm.n1490 C9_N_btm.n805 0.109875
R48221 C9_N_btm.n1495 C9_N_btm.n804 0.109875
R48222 C9_N_btm.n1493 C9_N_btm.n804 0.109875
R48223 C9_N_btm.n1498 C9_N_btm.n803 0.109875
R48224 C9_N_btm.n1496 C9_N_btm.n803 0.109875
R48225 C9_N_btm.n1501 C9_N_btm.n802 0.109875
R48226 C9_N_btm.n1499 C9_N_btm.n802 0.109875
R48227 C9_N_btm.n1504 C9_N_btm.n801 0.109875
R48228 C9_N_btm.n1502 C9_N_btm.n801 0.109875
R48229 C9_N_btm.n1507 C9_N_btm.n800 0.109875
R48230 C9_N_btm.n1505 C9_N_btm.n800 0.109875
R48231 C9_N_btm.n344 C9_N_btm.n315 0.109875
R48232 C9_N_btm.n346 C9_N_btm.n315 0.109875
R48233 C9_N_btm.n341 C9_N_btm.n317 0.109875
R48234 C9_N_btm.n343 C9_N_btm.n317 0.109875
R48235 C9_N_btm.n338 C9_N_btm.n318 0.109875
R48236 C9_N_btm.n340 C9_N_btm.n318 0.109875
R48237 C9_N_btm.n335 C9_N_btm.n332 0.109875
R48238 C9_N_btm.n337 C9_N_btm.n332 0.109875
R48239 C9_N_btm.n331 C9_N_btm.n320 0.109875
R48240 C9_N_btm.n331 C9_N_btm.n330 0.109875
R48241 C9_N_btm.n328 C9_N_btm.n321 0.109875
R48242 C9_N_btm.n326 C9_N_btm.n321 0.109875
R48243 C9_N_btm.n325 C9_N_btm.n322 0.109875
R48244 C9_N_btm.n323 C9_N_btm.n322 0.109875
R48245 C9_N_btm.n353 C9_N_btm.n316 0.109875
R48246 C9_N_btm.n353 C9_N_btm.n352 0.109875
R48247 C9_N_btm.n358 C9_N_btm.n354 0.109875
R48248 C9_N_btm.n356 C9_N_btm.n354 0.109875
R48249 C9_N_btm.n361 C9_N_btm.n314 0.109875
R48250 C9_N_btm.n359 C9_N_btm.n314 0.109875
R48251 C9_N_btm.n364 C9_N_btm.n313 0.109875
R48252 C9_N_btm.n362 C9_N_btm.n313 0.109875
R48253 C9_N_btm.n367 C9_N_btm.n312 0.109875
R48254 C9_N_btm.n365 C9_N_btm.n312 0.109875
R48255 C9_N_btm.n372 C9_N_btm.n310 0.109875
R48256 C9_N_btm.n374 C9_N_btm.n310 0.109875
R48257 C9_N_btm.n375 C9_N_btm.n296 0.109875
R48258 C9_N_btm.n377 C9_N_btm.n296 0.109875
R48259 C9_N_btm.n378 C9_N_btm.n295 0.109875
R48260 C9_N_btm.n380 C9_N_btm.n295 0.109875
R48261 C9_N_btm.n381 C9_N_btm.n292 0.109875
R48262 C9_N_btm.n383 C9_N_btm.n292 0.109875
R48263 C9_N_btm.n390 C9_N_btm.n293 0.109875
R48264 C9_N_btm.n390 C9_N_btm.n389 0.109875
R48265 C9_N_btm.n303 C9_N_btm.n300 0.109875
R48266 C9_N_btm.n301 C9_N_btm.n300 0.109875
R48267 C9_N_btm.n306 C9_N_btm.n299 0.109875
R48268 C9_N_btm.n304 C9_N_btm.n299 0.109875
R48269 C9_N_btm.n309 C9_N_btm.n298 0.109875
R48270 C9_N_btm.n309 C9_N_btm.n308 0.109875
R48271 C9_N_btm.n404 C9_N_btm.n289 0.109875
R48272 C9_N_btm.n402 C9_N_btm.n289 0.109875
R48273 C9_N_btm.n401 C9_N_btm.n290 0.109875
R48274 C9_N_btm.n399 C9_N_btm.n290 0.109875
R48275 C9_N_btm.n398 C9_N_btm.n291 0.109875
R48276 C9_N_btm.n396 C9_N_btm.n291 0.109875
R48277 C9_N_btm.n395 C9_N_btm.n391 0.109875
R48278 C9_N_btm.n393 C9_N_btm.n391 0.109875
R48279 C9_N_btm.n418 C9_N_btm.n269 0.109875
R48280 C9_N_btm.n420 C9_N_btm.n269 0.109875
R48281 C9_N_btm.n415 C9_N_btm.n272 0.109875
R48282 C9_N_btm.n417 C9_N_btm.n272 0.109875
R48283 C9_N_btm.n412 C9_N_btm.n273 0.109875
R48284 C9_N_btm.n414 C9_N_btm.n273 0.109875
R48285 C9_N_btm.n409 C9_N_btm.n287 0.109875
R48286 C9_N_btm.n411 C9_N_btm.n287 0.109875
R48287 C9_N_btm.n286 C9_N_btm.n275 0.109875
R48288 C9_N_btm.n286 C9_N_btm.n285 0.109875
R48289 C9_N_btm.n283 C9_N_btm.n276 0.109875
R48290 C9_N_btm.n281 C9_N_btm.n276 0.109875
R48291 C9_N_btm.n280 C9_N_btm.n277 0.109875
R48292 C9_N_btm.n278 C9_N_btm.n277 0.109875
R48293 C9_N_btm.n427 C9_N_btm.n270 0.109875
R48294 C9_N_btm.n427 C9_N_btm.n426 0.109875
R48295 C9_N_btm.n432 C9_N_btm.n428 0.109875
R48296 C9_N_btm.n430 C9_N_btm.n428 0.109875
R48297 C9_N_btm.n435 C9_N_btm.n268 0.109875
R48298 C9_N_btm.n433 C9_N_btm.n268 0.109875
R48299 C9_N_btm.n438 C9_N_btm.n267 0.109875
R48300 C9_N_btm.n436 C9_N_btm.n267 0.109875
R48301 C9_N_btm.n441 C9_N_btm.n266 0.109875
R48302 C9_N_btm.n439 C9_N_btm.n266 0.109875
R48303 C9_N_btm.n446 C9_N_btm.n264 0.109875
R48304 C9_N_btm.n448 C9_N_btm.n264 0.109875
R48305 C9_N_btm.n449 C9_N_btm.n250 0.109875
R48306 C9_N_btm.n451 C9_N_btm.n250 0.109875
R48307 C9_N_btm.n452 C9_N_btm.n249 0.109875
R48308 C9_N_btm.n454 C9_N_btm.n249 0.109875
R48309 C9_N_btm.n455 C9_N_btm.n246 0.109875
R48310 C9_N_btm.n457 C9_N_btm.n246 0.109875
R48311 C9_N_btm.n464 C9_N_btm.n247 0.109875
R48312 C9_N_btm.n464 C9_N_btm.n463 0.109875
R48313 C9_N_btm.n257 C9_N_btm.n254 0.109875
R48314 C9_N_btm.n255 C9_N_btm.n254 0.109875
R48315 C9_N_btm.n260 C9_N_btm.n253 0.109875
R48316 C9_N_btm.n258 C9_N_btm.n253 0.109875
R48317 C9_N_btm.n263 C9_N_btm.n252 0.109875
R48318 C9_N_btm.n263 C9_N_btm.n262 0.109875
R48319 C9_N_btm.n478 C9_N_btm.n243 0.109875
R48320 C9_N_btm.n476 C9_N_btm.n243 0.109875
R48321 C9_N_btm.n475 C9_N_btm.n244 0.109875
R48322 C9_N_btm.n473 C9_N_btm.n244 0.109875
R48323 C9_N_btm.n472 C9_N_btm.n245 0.109875
R48324 C9_N_btm.n470 C9_N_btm.n245 0.109875
R48325 C9_N_btm.n469 C9_N_btm.n465 0.109875
R48326 C9_N_btm.n467 C9_N_btm.n465 0.109875
R48327 C9_N_btm.n492 C9_N_btm.n223 0.109875
R48328 C9_N_btm.n494 C9_N_btm.n223 0.109875
R48329 C9_N_btm.n489 C9_N_btm.n226 0.109875
R48330 C9_N_btm.n491 C9_N_btm.n226 0.109875
R48331 C9_N_btm.n486 C9_N_btm.n227 0.109875
R48332 C9_N_btm.n488 C9_N_btm.n227 0.109875
R48333 C9_N_btm.n483 C9_N_btm.n241 0.109875
R48334 C9_N_btm.n485 C9_N_btm.n241 0.109875
R48335 C9_N_btm.n240 C9_N_btm.n229 0.109875
R48336 C9_N_btm.n240 C9_N_btm.n239 0.109875
R48337 C9_N_btm.n237 C9_N_btm.n230 0.109875
R48338 C9_N_btm.n235 C9_N_btm.n230 0.109875
R48339 C9_N_btm.n234 C9_N_btm.n231 0.109875
R48340 C9_N_btm.n232 C9_N_btm.n231 0.109875
R48341 C9_N_btm.n501 C9_N_btm.n224 0.109875
R48342 C9_N_btm.n501 C9_N_btm.n500 0.109875
R48343 C9_N_btm.n506 C9_N_btm.n502 0.109875
R48344 C9_N_btm.n504 C9_N_btm.n502 0.109875
R48345 C9_N_btm.n509 C9_N_btm.n222 0.109875
R48346 C9_N_btm.n507 C9_N_btm.n222 0.109875
R48347 C9_N_btm.n512 C9_N_btm.n221 0.109875
R48348 C9_N_btm.n510 C9_N_btm.n221 0.109875
R48349 C9_N_btm.n515 C9_N_btm.n220 0.109875
R48350 C9_N_btm.n513 C9_N_btm.n220 0.109875
R48351 C9_N_btm.n522 C9_N_btm.n210 0.109875
R48352 C9_N_btm.n524 C9_N_btm.n210 0.109875
R48353 C9_N_btm.n525 C9_N_btm.n218 0.109875
R48354 C9_N_btm.n527 C9_N_btm.n218 0.109875
R48355 C9_N_btm.n528 C9_N_btm.n217 0.109875
R48356 C9_N_btm.n530 C9_N_btm.n217 0.109875
R48357 C9_N_btm.n531 C9_N_btm.n216 0.109875
R48358 C9_N_btm.n533 C9_N_btm.n216 0.109875
R48359 C9_N_btm.n540 C9_N_btm.n214 0.109875
R48360 C9_N_btm.n538 C9_N_btm.n214 0.109875
R48361 C9_N_btm.n543 C9_N_btm.n213 0.109875
R48362 C9_N_btm.n541 C9_N_btm.n213 0.109875
R48363 C9_N_btm.n546 C9_N_btm.n212 0.109875
R48364 C9_N_btm.n544 C9_N_btm.n212 0.109875
R48365 C9_N_btm.n549 C9_N_btm.n211 0.109875
R48366 C9_N_btm.n549 C9_N_btm.n548 0.109875
R48367 C9_N_btm.n552 C9_N_btm.n550 0.109875
R48368 C9_N_btm.n554 C9_N_btm.n550 0.109875
R48369 C9_N_btm.n555 C9_N_btm.n209 0.109875
R48370 C9_N_btm.n557 C9_N_btm.n209 0.109875
R48371 C9_N_btm.n558 C9_N_btm.n208 0.109875
R48372 C9_N_btm.n560 C9_N_btm.n208 0.109875
R48373 C9_N_btm.n561 C9_N_btm.n207 0.109875
R48374 C9_N_btm.n563 C9_N_btm.n207 0.109875
R48375 C9_N_btm.n564 C9_N_btm.n206 0.109875
R48376 C9_N_btm.n566 C9_N_btm.n206 0.109875
R48377 C9_N_btm.n567 C9_N_btm.n205 0.109875
R48378 C9_N_btm.n569 C9_N_btm.n205 0.109875
R48379 C9_N_btm.n570 C9_N_btm.n204 0.109875
R48380 C9_N_btm.n572 C9_N_btm.n204 0.109875
R48381 C9_N_btm.n573 C9_N_btm.n203 0.109875
R48382 C9_N_btm.n575 C9_N_btm.n203 0.109875
R48383 C9_N_btm.n576 C9_N_btm.n202 0.109875
R48384 C9_N_btm.n578 C9_N_btm.n202 0.109875
R48385 C9_N_btm.n579 C9_N_btm.n201 0.109875
R48386 C9_N_btm.n581 C9_N_btm.n201 0.109875
R48387 C9_N_btm.n582 C9_N_btm.n200 0.109875
R48388 C9_N_btm.n584 C9_N_btm.n200 0.109875
R48389 C9_N_btm.n585 C9_N_btm.n199 0.109875
R48390 C9_N_btm.n587 C9_N_btm.n199 0.109875
R48391 C9_N_btm.n588 C9_N_btm.n198 0.109875
R48392 C9_N_btm.n590 C9_N_btm.n198 0.109875
R48393 C9_N_btm.n591 C9_N_btm.n197 0.109875
R48394 C9_N_btm.n593 C9_N_btm.n197 0.109875
R48395 C9_N_btm.n594 C9_N_btm.n196 0.109875
R48396 C9_N_btm.n596 C9_N_btm.n196 0.109875
R48397 C9_N_btm.n597 C9_N_btm.n195 0.109875
R48398 C9_N_btm.n599 C9_N_btm.n195 0.109875
R48399 C9_N_btm.n600 C9_N_btm.n194 0.109875
R48400 C9_N_btm.n602 C9_N_btm.n194 0.109875
R48401 C9_N_btm.n603 C9_N_btm.n193 0.109875
R48402 C9_N_btm.n605 C9_N_btm.n193 0.109875
R48403 C9_N_btm.n736 C9_N_btm.n609 0.109875
R48404 C9_N_btm.n734 C9_N_btm.n609 0.109875
R48405 C9_N_btm.n739 C9_N_btm.n608 0.109875
R48406 C9_N_btm.n737 C9_N_btm.n608 0.109875
R48407 C9_N_btm.n742 C9_N_btm.n607 0.109875
R48408 C9_N_btm.n740 C9_N_btm.n607 0.109875
R48409 C9_N_btm.n745 C9_N_btm.n192 0.109875
R48410 C9_N_btm.n743 C9_N_btm.n192 0.109875
R48411 C9_N_btm.n748 C9_N_btm.n191 0.109875
R48412 C9_N_btm.n746 C9_N_btm.n191 0.109875
R48413 C9_N_btm.n751 C9_N_btm.n190 0.109875
R48414 C9_N_btm.n749 C9_N_btm.n190 0.109875
R48415 C9_N_btm.n754 C9_N_btm.n189 0.109875
R48416 C9_N_btm.n752 C9_N_btm.n189 0.109875
R48417 C9_N_btm.n757 C9_N_btm.n188 0.109875
R48418 C9_N_btm.n755 C9_N_btm.n188 0.109875
R48419 C9_N_btm.n760 C9_N_btm.n187 0.109875
R48420 C9_N_btm.n758 C9_N_btm.n187 0.109875
R48421 C9_N_btm.n763 C9_N_btm.n186 0.109875
R48422 C9_N_btm.n761 C9_N_btm.n186 0.109875
R48423 C9_N_btm.n766 C9_N_btm.n185 0.109875
R48424 C9_N_btm.n764 C9_N_btm.n185 0.109875
R48425 C9_N_btm.n769 C9_N_btm.n184 0.109875
R48426 C9_N_btm.n767 C9_N_btm.n184 0.109875
R48427 C9_N_btm.n772 C9_N_btm.n183 0.109875
R48428 C9_N_btm.n770 C9_N_btm.n183 0.109875
R48429 C9_N_btm.n775 C9_N_btm.n182 0.109875
R48430 C9_N_btm.n773 C9_N_btm.n182 0.109875
R48431 C9_N_btm.n778 C9_N_btm.n181 0.109875
R48432 C9_N_btm.n776 C9_N_btm.n181 0.109875
R48433 C9_N_btm.n781 C9_N_btm.n180 0.109875
R48434 C9_N_btm.n779 C9_N_btm.n180 0.109875
R48435 C9_N_btm.n784 C9_N_btm.n179 0.109875
R48436 C9_N_btm.n782 C9_N_btm.n179 0.109875
R48437 C9_N_btm.n787 C9_N_btm.n178 0.109875
R48438 C9_N_btm.n785 C9_N_btm.n178 0.109875
R48439 C9_N_btm.n790 C9_N_btm.n177 0.109875
R48440 C9_N_btm.n788 C9_N_btm.n177 0.109875
R48441 C9_N_btm.n793 C9_N_btm.n176 0.109875
R48442 C9_N_btm.n791 C9_N_btm.n176 0.109875
R48443 C9_N_btm.n796 C9_N_btm.n175 0.109875
R48444 C9_N_btm.n794 C9_N_btm.n175 0.109875
R48445 C9_N_btm.n1512 C9_N_btm.n173 0.109875
R48446 C9_N_btm.n1514 C9_N_btm.n173 0.109875
R48447 C9_N_btm.n1515 C9_N_btm.n172 0.109875
R48448 C9_N_btm.n1517 C9_N_btm.n172 0.109875
R48449 C9_N_btm.n1518 C9_N_btm.n171 0.109875
R48450 C9_N_btm.n1520 C9_N_btm.n171 0.109875
R48451 C9_N_btm.n1521 C9_N_btm.n170 0.109875
R48452 C9_N_btm.n1523 C9_N_btm.n170 0.109875
R48453 C9_N_btm.n1524 C9_N_btm.n169 0.109875
R48454 C9_N_btm.n1526 C9_N_btm.n169 0.109875
R48455 C9_N_btm.n1527 C9_N_btm.n168 0.109875
R48456 C9_N_btm.n1529 C9_N_btm.n168 0.109875
R48457 C9_N_btm.n1530 C9_N_btm.n167 0.109875
R48458 C9_N_btm.n1532 C9_N_btm.n167 0.109875
R48459 C9_N_btm.n1533 C9_N_btm.n166 0.109875
R48460 C9_N_btm.n1535 C9_N_btm.n166 0.109875
R48461 C9_N_btm.n1536 C9_N_btm.n165 0.109875
R48462 C9_N_btm.n1538 C9_N_btm.n165 0.109875
R48463 C9_N_btm.n1539 C9_N_btm.n164 0.109875
R48464 C9_N_btm.n1541 C9_N_btm.n164 0.109875
R48465 C9_N_btm.n1542 C9_N_btm.n163 0.109875
R48466 C9_N_btm.n1544 C9_N_btm.n163 0.109875
R48467 C9_N_btm.n1545 C9_N_btm.n162 0.109875
R48468 C9_N_btm.n1547 C9_N_btm.n162 0.109875
R48469 C9_N_btm.n1548 C9_N_btm.n161 0.109875
R48470 C9_N_btm.n1550 C9_N_btm.n161 0.109875
R48471 C9_N_btm.n1551 C9_N_btm.n160 0.109875
R48472 C9_N_btm.n1553 C9_N_btm.n160 0.109875
R48473 C9_N_btm.n1554 C9_N_btm.n159 0.109875
R48474 C9_N_btm.n1556 C9_N_btm.n159 0.109875
R48475 C9_N_btm.n1557 C9_N_btm.n158 0.109875
R48476 C9_N_btm.n1559 C9_N_btm.n158 0.109875
R48477 C9_N_btm.n1560 C9_N_btm.n157 0.109875
R48478 C9_N_btm.n1562 C9_N_btm.n157 0.109875
R48479 C9_N_btm.n1563 C9_N_btm.n156 0.109875
R48480 C9_N_btm.n1565 C9_N_btm.n156 0.109875
R48481 C9_N_btm.n1566 C9_N_btm.n155 0.109875
R48482 C9_N_btm.n1568 C9_N_btm.n155 0.109875
R48483 C9_N_btm.n1569 C9_N_btm.n154 0.109875
R48484 C9_N_btm.n1571 C9_N_btm.n154 0.109875
R48485 C9_N_btm.n1572 C9_N_btm.n153 0.109875
R48486 C9_N_btm.n1574 C9_N_btm.n153 0.109875
R48487 C9_N_btm.n1575 C9_N_btm.n152 0.109875
R48488 C9_N_btm.n1577 C9_N_btm.n152 0.109875
R48489 C9_N_btm.n1578 C9_N_btm.n151 0.109875
R48490 C9_N_btm.n1580 C9_N_btm.n151 0.109875
R48491 C9_N_btm.n1581 C9_N_btm.n150 0.109875
R48492 C9_N_btm.n1583 C9_N_btm.n150 0.109875
R48493 C9_N_btm.n1584 C9_N_btm.n149 0.109875
R48494 C9_N_btm.n1586 C9_N_btm.n149 0.109875
R48495 C9_N_btm.n1587 C9_N_btm.n148 0.109875
R48496 C9_N_btm.n1589 C9_N_btm.n148 0.109875
R48497 C9_N_btm.n1590 C9_N_btm.n147 0.109875
R48498 C9_N_btm.n1592 C9_N_btm.n147 0.109875
R48499 C9_N_btm.n1593 C9_N_btm.n146 0.109875
R48500 C9_N_btm.n1595 C9_N_btm.n146 0.109875
R48501 C9_N_btm.n1596 C9_N_btm.n145 0.109875
R48502 C9_N_btm.n1598 C9_N_btm.n145 0.109875
R48503 C9_N_btm.n1599 C9_N_btm.n144 0.109875
R48504 C9_N_btm.n1601 C9_N_btm.n144 0.109875
R48505 C9_N_btm.n1602 C9_N_btm.n143 0.109875
R48506 C9_N_btm.n1604 C9_N_btm.n143 0.109875
R48507 C9_N_btm.n1605 C9_N_btm.n142 0.109875
R48508 C9_N_btm.n1607 C9_N_btm.n142 0.109875
R48509 C9_N_btm.n1608 C9_N_btm.n141 0.109875
R48510 C9_N_btm.n1610 C9_N_btm.n141 0.109875
R48511 C9_N_btm.n1611 C9_N_btm.n140 0.109875
R48512 C9_N_btm.n1613 C9_N_btm.n140 0.109875
R48513 C9_N_btm.n1614 C9_N_btm.n139 0.109875
R48514 C9_N_btm.n1616 C9_N_btm.n139 0.109875
R48515 C9_N_btm.n1617 C9_N_btm.n138 0.109875
R48516 C9_N_btm.n1619 C9_N_btm.n138 0.109875
R48517 C9_N_btm.n1620 C9_N_btm.n137 0.109875
R48518 C9_N_btm.n1622 C9_N_btm.n137 0.109875
R48519 C9_N_btm.n1623 C9_N_btm.n136 0.109875
R48520 C9_N_btm.n1625 C9_N_btm.n136 0.109875
R48521 C9_N_btm.n1626 C9_N_btm.n135 0.109875
R48522 C9_N_btm.n1628 C9_N_btm.n135 0.109875
R48523 C9_N_btm.n1629 C9_N_btm.n132 0.109875
R48524 C9_N_btm.n1631 C9_N_btm.n132 0.109875
R48525 C9_N_btm.n1638 C9_N_btm.n133 0.109875
R48526 C9_N_btm.n1638 C9_N_btm.n1637 0.109875
R48527 C9_N_btm.n682 C9_N_btm.n679 0.109875
R48528 C9_N_btm.n680 C9_N_btm.n679 0.109875
R48529 C9_N_btm.n685 C9_N_btm.n678 0.109875
R48530 C9_N_btm.n683 C9_N_btm.n678 0.109875
R48531 C9_N_btm.n688 C9_N_btm.n677 0.109875
R48532 C9_N_btm.n686 C9_N_btm.n677 0.109875
R48533 C9_N_btm.n691 C9_N_btm.n127 0.109875
R48534 C9_N_btm.n689 C9_N_btm.n127 0.109875
R48535 C9_N_btm.n694 C9_N_btm.n676 0.109875
R48536 C9_N_btm.n692 C9_N_btm.n676 0.109875
R48537 C9_N_btm.n697 C9_N_btm.n622 0.109875
R48538 C9_N_btm.n695 C9_N_btm.n622 0.109875
R48539 C9_N_btm.n700 C9_N_btm.n621 0.109875
R48540 C9_N_btm.n698 C9_N_btm.n621 0.109875
R48541 C9_N_btm.n703 C9_N_btm.n620 0.109875
R48542 C9_N_btm.n701 C9_N_btm.n620 0.109875
R48543 C9_N_btm.n706 C9_N_btm.n619 0.109875
R48544 C9_N_btm.n704 C9_N_btm.n619 0.109875
R48545 C9_N_btm.n709 C9_N_btm.n618 0.109875
R48546 C9_N_btm.n707 C9_N_btm.n618 0.109875
R48547 C9_N_btm.n712 C9_N_btm.n617 0.109875
R48548 C9_N_btm.n710 C9_N_btm.n617 0.109875
R48549 C9_N_btm.n715 C9_N_btm.n616 0.109875
R48550 C9_N_btm.n713 C9_N_btm.n616 0.109875
R48551 C9_N_btm.n718 C9_N_btm.n615 0.109875
R48552 C9_N_btm.n716 C9_N_btm.n615 0.109875
R48553 C9_N_btm.n721 C9_N_btm.n614 0.109875
R48554 C9_N_btm.n719 C9_N_btm.n614 0.109875
R48555 C9_N_btm.n724 C9_N_btm.n613 0.109875
R48556 C9_N_btm.n722 C9_N_btm.n613 0.109875
R48557 C9_N_btm.n727 C9_N_btm.n612 0.109875
R48558 C9_N_btm.n725 C9_N_btm.n612 0.109875
R48559 C9_N_btm.n730 C9_N_btm.n611 0.109875
R48560 C9_N_btm.n728 C9_N_btm.n611 0.109875
R48561 C9_N_btm.n733 C9_N_btm.n610 0.109875
R48562 C9_N_btm.n731 C9_N_btm.n610 0.109875
R48563 C9_N_btm.n636 C9_N_btm.n634 0.109875
R48564 C9_N_btm.n638 C9_N_btm.n634 0.109875
R48565 C9_N_btm.n639 C9_N_btm.n633 0.109875
R48566 C9_N_btm.n641 C9_N_btm.n633 0.109875
R48567 C9_N_btm.n642 C9_N_btm.n632 0.109875
R48568 C9_N_btm.n644 C9_N_btm.n632 0.109875
R48569 C9_N_btm.n645 C9_N_btm.n631 0.109875
R48570 C9_N_btm.n647 C9_N_btm.n631 0.109875
R48571 C9_N_btm.n648 C9_N_btm.n630 0.109875
R48572 C9_N_btm.n650 C9_N_btm.n630 0.109875
R48573 C9_N_btm.n651 C9_N_btm.n629 0.109875
R48574 C9_N_btm.n653 C9_N_btm.n629 0.109875
R48575 C9_N_btm.n654 C9_N_btm.n628 0.109875
R48576 C9_N_btm.n656 C9_N_btm.n628 0.109875
R48577 C9_N_btm.n657 C9_N_btm.n627 0.109875
R48578 C9_N_btm.n659 C9_N_btm.n627 0.109875
R48579 C9_N_btm.n660 C9_N_btm.n626 0.109875
R48580 C9_N_btm.n662 C9_N_btm.n626 0.109875
R48581 C9_N_btm.n663 C9_N_btm.n625 0.109875
R48582 C9_N_btm.n665 C9_N_btm.n625 0.109875
R48583 C9_N_btm.n666 C9_N_btm.n624 0.109875
R48584 C9_N_btm.n668 C9_N_btm.n624 0.109875
R48585 C9_N_btm.n669 C9_N_btm.n623 0.109875
R48586 C9_N_btm.n671 C9_N_btm.n623 0.109875
R48587 C9_N_btm.n675 C9_N_btm.n672 0.109875
R48588 C9_N_btm.n675 C9_N_btm.n674 0.109875
R48589 C9_N_btm.n1655 C9_N_btm.n128 0.109875
R48590 C9_N_btm.n1655 C9_N_btm.n1654 0.109875
R48591 C9_N_btm.n1652 C9_N_btm.n129 0.109875
R48592 C9_N_btm.n1650 C9_N_btm.n129 0.109875
R48593 C9_N_btm.n1649 C9_N_btm.n130 0.109875
R48594 C9_N_btm.n1647 C9_N_btm.n130 0.109875
R48595 C9_N_btm.n1646 C9_N_btm.n131 0.109875
R48596 C9_N_btm.n1644 C9_N_btm.n131 0.109875
R48597 C9_N_btm.n1643 C9_N_btm.n1639 0.109875
R48598 C9_N_btm.n1641 C9_N_btm.n1639 0.109875
R48599 C9_N_btm.n1667 C9_N_btm.n108 0.109875
R48600 C9_N_btm.n1669 C9_N_btm.n108 0.109875
R48601 C9_N_btm.n1664 C9_N_btm.n111 0.109875
R48602 C9_N_btm.n1666 C9_N_btm.n111 0.109875
R48603 C9_N_btm.n1661 C9_N_btm.n112 0.109875
R48604 C9_N_btm.n1663 C9_N_btm.n112 0.109875
R48605 C9_N_btm.n1658 C9_N_btm.n126 0.109875
R48606 C9_N_btm.n1660 C9_N_btm.n126 0.109875
R48607 C9_N_btm.n125 C9_N_btm.n114 0.109875
R48608 C9_N_btm.n125 C9_N_btm.n124 0.109875
R48609 C9_N_btm.n122 C9_N_btm.n115 0.109875
R48610 C9_N_btm.n120 C9_N_btm.n115 0.109875
R48611 C9_N_btm.n119 C9_N_btm.n116 0.109875
R48612 C9_N_btm.n117 C9_N_btm.n116 0.109875
R48613 C9_N_btm.n1676 C9_N_btm.n109 0.109875
R48614 C9_N_btm.n1676 C9_N_btm.n1675 0.109875
R48615 C9_N_btm.n1681 C9_N_btm.n1677 0.109875
R48616 C9_N_btm.n1679 C9_N_btm.n1677 0.109875
R48617 C9_N_btm.n1684 C9_N_btm.n107 0.109875
R48618 C9_N_btm.n1682 C9_N_btm.n107 0.109875
R48619 C9_N_btm.n1687 C9_N_btm.n106 0.109875
R48620 C9_N_btm.n1685 C9_N_btm.n106 0.109875
R48621 C9_N_btm.n1690 C9_N_btm.n105 0.109875
R48622 C9_N_btm.n1688 C9_N_btm.n105 0.109875
R48623 C9_N_btm.n1695 C9_N_btm.n103 0.109875
R48624 C9_N_btm.n1697 C9_N_btm.n103 0.109875
R48625 C9_N_btm.n1698 C9_N_btm.n89 0.109875
R48626 C9_N_btm.n1700 C9_N_btm.n89 0.109875
R48627 C9_N_btm.n1701 C9_N_btm.n88 0.109875
R48628 C9_N_btm.n1703 C9_N_btm.n88 0.109875
R48629 C9_N_btm.n1704 C9_N_btm.n85 0.109875
R48630 C9_N_btm.n1706 C9_N_btm.n85 0.109875
R48631 C9_N_btm.n1713 C9_N_btm.n86 0.109875
R48632 C9_N_btm.n1713 C9_N_btm.n1712 0.109875
R48633 C9_N_btm.n96 C9_N_btm.n93 0.109875
R48634 C9_N_btm.n94 C9_N_btm.n93 0.109875
R48635 C9_N_btm.n99 C9_N_btm.n92 0.109875
R48636 C9_N_btm.n97 C9_N_btm.n92 0.109875
R48637 C9_N_btm.n102 C9_N_btm.n91 0.109875
R48638 C9_N_btm.n102 C9_N_btm.n101 0.109875
R48639 C9_N_btm.n1727 C9_N_btm.n82 0.109875
R48640 C9_N_btm.n1725 C9_N_btm.n82 0.109875
R48641 C9_N_btm.n1724 C9_N_btm.n83 0.109875
R48642 C9_N_btm.n1722 C9_N_btm.n83 0.109875
R48643 C9_N_btm.n1721 C9_N_btm.n84 0.109875
R48644 C9_N_btm.n1719 C9_N_btm.n84 0.109875
R48645 C9_N_btm.n1718 C9_N_btm.n1714 0.109875
R48646 C9_N_btm.n1716 C9_N_btm.n1714 0.109875
R48647 C9_N_btm.n1741 C9_N_btm.n62 0.109875
R48648 C9_N_btm.n1743 C9_N_btm.n62 0.109875
R48649 C9_N_btm.n1738 C9_N_btm.n65 0.109875
R48650 C9_N_btm.n1740 C9_N_btm.n65 0.109875
R48651 C9_N_btm.n1735 C9_N_btm.n66 0.109875
R48652 C9_N_btm.n1737 C9_N_btm.n66 0.109875
R48653 C9_N_btm.n1732 C9_N_btm.n80 0.109875
R48654 C9_N_btm.n1734 C9_N_btm.n80 0.109875
R48655 C9_N_btm.n79 C9_N_btm.n68 0.109875
R48656 C9_N_btm.n79 C9_N_btm.n78 0.109875
R48657 C9_N_btm.n76 C9_N_btm.n69 0.109875
R48658 C9_N_btm.n74 C9_N_btm.n69 0.109875
R48659 C9_N_btm.n73 C9_N_btm.n70 0.109875
R48660 C9_N_btm.n71 C9_N_btm.n70 0.109875
R48661 C9_N_btm.n1750 C9_N_btm.n63 0.109875
R48662 C9_N_btm.n1750 C9_N_btm.n1749 0.109875
R48663 C9_N_btm.n1755 C9_N_btm.n1751 0.109875
R48664 C9_N_btm.n1753 C9_N_btm.n1751 0.109875
R48665 C9_N_btm.n1758 C9_N_btm.n61 0.109875
R48666 C9_N_btm.n1756 C9_N_btm.n61 0.109875
R48667 C9_N_btm.n1761 C9_N_btm.n60 0.109875
R48668 C9_N_btm.n1759 C9_N_btm.n60 0.109875
R48669 C9_N_btm.n1764 C9_N_btm.n59 0.109875
R48670 C9_N_btm.n1762 C9_N_btm.n59 0.109875
R48671 C9_N_btm.n1769 C9_N_btm.n57 0.109875
R48672 C9_N_btm.n1771 C9_N_btm.n57 0.109875
R48673 C9_N_btm.n1772 C9_N_btm.n43 0.109875
R48674 C9_N_btm.n1774 C9_N_btm.n43 0.109875
R48675 C9_N_btm.n1775 C9_N_btm.n42 0.109875
R48676 C9_N_btm.n1777 C9_N_btm.n42 0.109875
R48677 C9_N_btm.n1778 C9_N_btm.n39 0.109875
R48678 C9_N_btm.n1780 C9_N_btm.n39 0.109875
R48679 C9_N_btm.n1787 C9_N_btm.n40 0.109875
R48680 C9_N_btm.n1787 C9_N_btm.n1786 0.109875
R48681 C9_N_btm.n50 C9_N_btm.n47 0.109875
R48682 C9_N_btm.n48 C9_N_btm.n47 0.109875
R48683 C9_N_btm.n53 C9_N_btm.n46 0.109875
R48684 C9_N_btm.n51 C9_N_btm.n46 0.109875
R48685 C9_N_btm.n56 C9_N_btm.n45 0.109875
R48686 C9_N_btm.n56 C9_N_btm.n55 0.109875
R48687 C9_N_btm.n1801 C9_N_btm.n36 0.109875
R48688 C9_N_btm.n1799 C9_N_btm.n36 0.109875
R48689 C9_N_btm.n1798 C9_N_btm.n37 0.109875
R48690 C9_N_btm.n1796 C9_N_btm.n37 0.109875
R48691 C9_N_btm.n1795 C9_N_btm.n38 0.109875
R48692 C9_N_btm.n1793 C9_N_btm.n38 0.109875
R48693 C9_N_btm.n1792 C9_N_btm.n1788 0.109875
R48694 C9_N_btm.n1790 C9_N_btm.n1788 0.109875
R48695 C9_N_btm.n1830 C9_N_btm.n29 0.109875
R48696 C9_N_btm.n1832 C9_N_btm.n29 0.109875
R48697 C9_N_btm.n1827 C9_N_btm.n32 0.109875
R48698 C9_N_btm.n1829 C9_N_btm.n32 0.109875
R48699 C9_N_btm.n1824 C9_N_btm.n33 0.109875
R48700 C9_N_btm.n1826 C9_N_btm.n33 0.109875
R48701 C9_N_btm.n1821 C9_N_btm.n34 0.109875
R48702 C9_N_btm.n1823 C9_N_btm.n34 0.109875
R48703 C9_N_btm.n1816 C9_N_btm.n25 0.109875
R48704 C9_N_btm.n1814 C9_N_btm.n25 0.109875
R48705 C9_N_btm.n1813 C9_N_btm.n1806 0.109875
R48706 C9_N_btm.n1811 C9_N_btm.n1806 0.109875
R48707 C9_N_btm.n1810 C9_N_btm.n1807 0.109875
R48708 C9_N_btm.n1808 C9_N_btm.n1807 0.109875
R48709 C9_N_btm.n1839 C9_N_btm.n30 0.109875
R48710 C9_N_btm.n1839 C9_N_btm.n1838 0.109875
R48711 C9_N_btm.n1844 C9_N_btm.n1840 0.109875
R48712 C9_N_btm.n1842 C9_N_btm.n1840 0.109875
R48713 C9_N_btm.n1847 C9_N_btm.n28 0.109875
R48714 C9_N_btm.n1845 C9_N_btm.n28 0.109875
R48715 C9_N_btm.n1850 C9_N_btm.n27 0.109875
R48716 C9_N_btm.n1848 C9_N_btm.n27 0.109875
R48717 C9_N_btm.n1853 C9_N_btm.n26 0.109875
R48718 C9_N_btm.n1853 C9_N_btm.n1852 0.109875
R48719 C9_N_btm.n1856 C9_N_btm.n1854 0.109875
R48720 C9_N_btm.n1858 C9_N_btm.n1854 0.109875
R48721 C9_N_btm.n1859 C9_N_btm.n24 0.109875
R48722 C9_N_btm.n1861 C9_N_btm.n24 0.109875
R48723 C9_N_btm.n1862 C9_N_btm.n23 0.109875
R48724 C9_N_btm.n1864 C9_N_btm.n23 0.109875
R48725 C9_N_btm.n1865 C9_N_btm.n22 0.109875
R48726 C9_N_btm.n1867 C9_N_btm.n22 0.109875
R48727 C9_N_btm.n1874 C9_N_btm.n20 0.109875
R48728 C9_N_btm.n1872 C9_N_btm.n20 0.109875
R48729 C9_N_btm.n1877 C9_N_btm.n19 0.109875
R48730 C9_N_btm.n1875 C9_N_btm.n19 0.109875
R48731 C9_N_btm.n1880 C9_N_btm.n18 0.109875
R48732 C9_N_btm.n1878 C9_N_btm.n18 0.109875
R48733 C9_N_btm.n1883 C9_N_btm.n17 0.109875
R48734 C9_N_btm.n1881 C9_N_btm.n17 0.109875
R48735 C9_N_btm.n1380 C9_N_btm.n1379 0.0556875
R48736 C9_N_btm.n1258 C9_N_btm.n1257 0.0556875
R48737 C9_N_btm.n880 C9_N_btm.n799 0.0556875
R48738 C9_N_btm.n1382 C9_N_btm.n1381 0.0556875
R48739 C9_N_btm.n1387 C9_N_btm.n134 0.0556875
R48740 C9_N_btm.n1509 C9_N_btm.n1508 0.0556875
R48741 C9_N_btm.n348 C9_N_btm.n347 0.0556875
R48742 C9_N_btm.n334 C9_N_btm.n333 0.0556875
R48743 C9_N_btm.n319 C9_N_btm.n311 0.0556875
R48744 C9_N_btm.n350 C9_N_btm.n349 0.0556875
R48745 C9_N_btm.n355 C9_N_btm.n294 0.0556875
R48746 C9_N_btm.n369 C9_N_btm.n368 0.0556875
R48747 C9_N_btm.n371 C9_N_btm.n370 0.0556875
R48748 C9_N_btm.n385 C9_N_btm.n384 0.0556875
R48749 C9_N_btm.n387 C9_N_btm.n386 0.0556875
R48750 C9_N_btm.n297 C9_N_btm.n288 0.0556875
R48751 C9_N_btm.n406 C9_N_btm.n405 0.0556875
R48752 C9_N_btm.n392 C9_N_btm.n271 0.0556875
R48753 C9_N_btm.n422 C9_N_btm.n421 0.0556875
R48754 C9_N_btm.n408 C9_N_btm.n407 0.0556875
R48755 C9_N_btm.n274 C9_N_btm.n265 0.0556875
R48756 C9_N_btm.n424 C9_N_btm.n423 0.0556875
R48757 C9_N_btm.n429 C9_N_btm.n248 0.0556875
R48758 C9_N_btm.n443 C9_N_btm.n442 0.0556875
R48759 C9_N_btm.n445 C9_N_btm.n444 0.0556875
R48760 C9_N_btm.n459 C9_N_btm.n458 0.0556875
R48761 C9_N_btm.n461 C9_N_btm.n460 0.0556875
R48762 C9_N_btm.n251 C9_N_btm.n242 0.0556875
R48763 C9_N_btm.n480 C9_N_btm.n479 0.0556875
R48764 C9_N_btm.n466 C9_N_btm.n225 0.0556875
R48765 C9_N_btm.n496 C9_N_btm.n495 0.0556875
R48766 C9_N_btm.n482 C9_N_btm.n481 0.0556875
R48767 C9_N_btm.n228 C9_N_btm.n219 0.0556875
R48768 C9_N_btm.n498 C9_N_btm.n497 0.0556875
R48769 C9_N_btm.n503 C9_N_btm.n215 0.0556875
R48770 C9_N_btm.n517 C9_N_btm.n516 0.0556875
R48771 C9_N_btm.n521 C9_N_btm.n520 0.0556875
R48772 C9_N_btm.n535 C9_N_btm.n534 0.0556875
R48773 C9_N_btm.n537 C9_N_btm.n536 0.0556875
R48774 C9_N_btm.n519 C9_N_btm.n518 0.0556875
R48775 C9_N_btm.n551 C9_N_btm.n174 0.0556875
R48776 C9_N_btm.n798 C9_N_btm.n797 0.0556875
R48777 C9_N_btm.n1511 C9_N_btm.n1510 0.0556875
R48778 C9_N_btm.n1633 C9_N_btm.n1632 0.0556875
R48779 C9_N_btm.n1635 C9_N_btm.n1634 0.0556875
R48780 C9_N_btm.n1640 C9_N_btm.n110 0.0556875
R48781 C9_N_btm.n1671 C9_N_btm.n1670 0.0556875
R48782 C9_N_btm.n1657 C9_N_btm.n1656 0.0556875
R48783 C9_N_btm.n113 C9_N_btm.n104 0.0556875
R48784 C9_N_btm.n1673 C9_N_btm.n1672 0.0556875
R48785 C9_N_btm.n1678 C9_N_btm.n87 0.0556875
R48786 C9_N_btm.n1692 C9_N_btm.n1691 0.0556875
R48787 C9_N_btm.n1694 C9_N_btm.n1693 0.0556875
R48788 C9_N_btm.n1708 C9_N_btm.n1707 0.0556875
R48789 C9_N_btm.n1710 C9_N_btm.n1709 0.0556875
R48790 C9_N_btm.n90 C9_N_btm.n81 0.0556875
R48791 C9_N_btm.n1729 C9_N_btm.n1728 0.0556875
R48792 C9_N_btm.n1715 C9_N_btm.n64 0.0556875
R48793 C9_N_btm.n1745 C9_N_btm.n1744 0.0556875
R48794 C9_N_btm.n1731 C9_N_btm.n1730 0.0556875
R48795 C9_N_btm.n67 C9_N_btm.n58 0.0556875
R48796 C9_N_btm.n1747 C9_N_btm.n1746 0.0556875
R48797 C9_N_btm.n1752 C9_N_btm.n41 0.0556875
R48798 C9_N_btm.n1766 C9_N_btm.n1765 0.0556875
R48799 C9_N_btm.n1768 C9_N_btm.n1767 0.0556875
R48800 C9_N_btm.n1782 C9_N_btm.n1781 0.0556875
R48801 C9_N_btm.n1784 C9_N_btm.n1783 0.0556875
R48802 C9_N_btm.n44 C9_N_btm.n35 0.0556875
R48803 C9_N_btm.n1803 C9_N_btm.n1802 0.0556875
R48804 C9_N_btm.n1789 C9_N_btm.n31 0.0556875
R48805 C9_N_btm.n1834 C9_N_btm.n1833 0.0556875
R48806 C9_N_btm.n1820 C9_N_btm.n1819 0.0556875
R48807 C9_N_btm.n1818 C9_N_btm.n1817 0.0556875
R48808 C9_N_btm.n1836 C9_N_btm.n1835 0.0556875
R48809 C9_N_btm.n1841 C9_N_btm.n21 0.0556875
R48810 C9_N_btm.n1805 C9_N_btm.n1804 0.0556875
R48811 C9_N_btm.n1855 C9_N_btm.n16 0.0556875
R48812 C9_N_btm.n1869 C9_N_btm.n1868 0.0556875
R48813 C9_N_btm.n1871 C9_N_btm.n1870 0.0556875
R48814 C9_N_btm.n1885 C9_N_btm.n1884 0.0556875
R48815 C9_P_btm C9_P_btm.n15 82.1463
R48816 C9_P_btm.n2 C9_P_btm.n0 33.0802
R48817 C9_P_btm.n6 C9_P_btm.n5 32.3614
R48818 C9_P_btm.n4 C9_P_btm.n3 32.3614
R48819 C9_P_btm.n2 C9_P_btm.n1 32.3614
R48820 C9_P_btm.n10 C9_P_btm.n6 24.0265
R48821 C9_P_btm.n11 C9_P_btm.t4 23.0826
R48822 C9_P_btm.n14 C9_P_btm.n12 15.4287
R48823 C9_P_btm.n9 C9_P_btm.n7 15.3784
R48824 C9_P_btm.n14 C9_P_btm.n13 14.9755
R48825 C9_P_btm.n9 C9_P_btm.n8 14.894
R48826 C9_P_btm.n15 C9_P_btm.n11 7.16717
R48827 C9_P_btm C9_P_btm.n1886 6.5255
R48828 C9_P_btm.n10 C9_P_btm.n9 5.71404
R48829 C9_P_btm.n15 C9_P_btm.n14 5.62029
R48830 C9_P_btm.n17 C9_P_btm.t18 5.03712
R48831 C9_P_btm.n18 C9_P_btm.t16 5.03712
R48832 C9_P_btm.n19 C9_P_btm.t17 5.03712
R48833 C9_P_btm.n20 C9_P_btm.t21 5.03712
R48834 C9_P_btm.n1870 C9_P_btm.t22 5.03712
R48835 C9_P_btm.n1046 C9_P_btm.t13 5.03712
R48836 C9_P_btm.n1045 C9_P_btm.t24 5.03712
R48837 C9_P_btm.n1031 C9_P_btm.t15 5.03712
R48838 C9_P_btm.n1030 C9_P_btm.t20 5.03712
R48839 C9_P_btm.n1028 C9_P_btm.t19 5.03712
R48840 C9_P_btm.n1061 C9_P_btm.t14 5.03712
R48841 C9_P_btm.n1883 C9_P_btm.n1882 4.60698
R48842 C9_P_btm.n1882 C9_P_btm.n1881 4.60698
R48843 C9_P_btm.n1880 C9_P_btm.n1879 4.60698
R48844 C9_P_btm.n1879 C9_P_btm.n1878 4.60698
R48845 C9_P_btm.n1877 C9_P_btm.n1876 4.60698
R48846 C9_P_btm.n1876 C9_P_btm.n1875 4.60698
R48847 C9_P_btm.n1874 C9_P_btm.n1873 4.60698
R48848 C9_P_btm.n1873 C9_P_btm.n1872 4.60698
R48849 C9_P_btm.n1867 C9_P_btm.n1866 4.60698
R48850 C9_P_btm.n1866 C9_P_btm.n1865 4.60698
R48851 C9_P_btm.n1864 C9_P_btm.n1863 4.60698
R48852 C9_P_btm.n1863 C9_P_btm.n1862 4.60698
R48853 C9_P_btm.n1861 C9_P_btm.n1860 4.60698
R48854 C9_P_btm.n1860 C9_P_btm.n1859 4.60698
R48855 C9_P_btm.n1858 C9_P_btm.n1857 4.60698
R48856 C9_P_btm.n1857 C9_P_btm.n1856 4.60698
R48857 C9_P_btm.n1852 C9_P_btm.n1851 4.60698
R48858 C9_P_btm.n1851 C9_P_btm.n26 4.60698
R48859 C9_P_btm.n1849 C9_P_btm.n1848 4.60698
R48860 C9_P_btm.n1850 C9_P_btm.n1849 4.60698
R48861 C9_P_btm.n1846 C9_P_btm.n1845 4.60698
R48862 C9_P_btm.n1847 C9_P_btm.n1846 4.60698
R48863 C9_P_btm.n1843 C9_P_btm.n1842 4.60698
R48864 C9_P_btm.n1844 C9_P_btm.n1843 4.60698
R48865 C9_P_btm.n1838 C9_P_btm.n1837 4.60698
R48866 C9_P_btm.n1837 C9_P_btm.n30 4.60698
R48867 C9_P_btm.n1809 C9_P_btm.n1808 4.60698
R48868 C9_P_btm.n1810 C9_P_btm.n1809 4.60698
R48869 C9_P_btm.n1812 C9_P_btm.n1811 4.60698
R48870 C9_P_btm.n1813 C9_P_btm.n1812 4.60698
R48871 C9_P_btm.n1815 C9_P_btm.n1814 4.60698
R48872 C9_P_btm.n1816 C9_P_btm.n1815 4.60698
R48873 C9_P_btm.n1823 C9_P_btm.n1822 4.60698
R48874 C9_P_btm.n1822 C9_P_btm.n1821 4.60698
R48875 C9_P_btm.n1826 C9_P_btm.n1825 4.60698
R48876 C9_P_btm.n1825 C9_P_btm.n1824 4.60698
R48877 C9_P_btm.n1829 C9_P_btm.n1828 4.60698
R48878 C9_P_btm.n1828 C9_P_btm.n1827 4.60698
R48879 C9_P_btm.n1832 C9_P_btm.n1831 4.60698
R48880 C9_P_btm.n1831 C9_P_btm.n1830 4.60698
R48881 C9_P_btm.n1791 C9_P_btm.n1790 4.60698
R48882 C9_P_btm.n1792 C9_P_btm.n1791 4.60698
R48883 C9_P_btm.n1794 C9_P_btm.n1793 4.60698
R48884 C9_P_btm.n1795 C9_P_btm.n1794 4.60698
R48885 C9_P_btm.n1797 C9_P_btm.n1796 4.60698
R48886 C9_P_btm.n1798 C9_P_btm.n1797 4.60698
R48887 C9_P_btm.n1800 C9_P_btm.n1799 4.60698
R48888 C9_P_btm.n1801 C9_P_btm.n1800 4.60698
R48889 C9_P_btm.n55 C9_P_btm.n54 4.60698
R48890 C9_P_btm.n54 C9_P_btm.n45 4.60698
R48891 C9_P_btm.n52 C9_P_btm.n51 4.60698
R48892 C9_P_btm.n53 C9_P_btm.n52 4.60698
R48893 C9_P_btm.n49 C9_P_btm.n48 4.60698
R48894 C9_P_btm.n50 C9_P_btm.n49 4.60698
R48895 C9_P_btm.n1786 C9_P_btm.n1785 4.60698
R48896 C9_P_btm.n1785 C9_P_btm.n40 4.60698
R48897 C9_P_btm.n1780 C9_P_btm.n1779 4.60698
R48898 C9_P_btm.n1779 C9_P_btm.n1778 4.60698
R48899 C9_P_btm.n1777 C9_P_btm.n1776 4.60698
R48900 C9_P_btm.n1776 C9_P_btm.n1775 4.60698
R48901 C9_P_btm.n1774 C9_P_btm.n1773 4.60698
R48902 C9_P_btm.n1773 C9_P_btm.n1772 4.60698
R48903 C9_P_btm.n1771 C9_P_btm.n1770 4.60698
R48904 C9_P_btm.n1770 C9_P_btm.n1769 4.60698
R48905 C9_P_btm.n1763 C9_P_btm.n1762 4.60698
R48906 C9_P_btm.n1764 C9_P_btm.n1763 4.60698
R48907 C9_P_btm.n1760 C9_P_btm.n1759 4.60698
R48908 C9_P_btm.n1761 C9_P_btm.n1760 4.60698
R48909 C9_P_btm.n1757 C9_P_btm.n1756 4.60698
R48910 C9_P_btm.n1758 C9_P_btm.n1757 4.60698
R48911 C9_P_btm.n1754 C9_P_btm.n1753 4.60698
R48912 C9_P_btm.n1755 C9_P_btm.n1754 4.60698
R48913 C9_P_btm.n1749 C9_P_btm.n1748 4.60698
R48914 C9_P_btm.n1748 C9_P_btm.n63 4.60698
R48915 C9_P_btm.n72 C9_P_btm.n71 4.60698
R48916 C9_P_btm.n73 C9_P_btm.n72 4.60698
R48917 C9_P_btm.n75 C9_P_btm.n74 4.60698
R48918 C9_P_btm.n76 C9_P_btm.n75 4.60698
R48919 C9_P_btm.n78 C9_P_btm.n77 4.60698
R48920 C9_P_btm.n77 C9_P_btm.n68 4.60698
R48921 C9_P_btm.n1734 C9_P_btm.n1733 4.60698
R48922 C9_P_btm.n1733 C9_P_btm.n1732 4.60698
R48923 C9_P_btm.n1737 C9_P_btm.n1736 4.60698
R48924 C9_P_btm.n1736 C9_P_btm.n1735 4.60698
R48925 C9_P_btm.n1740 C9_P_btm.n1739 4.60698
R48926 C9_P_btm.n1739 C9_P_btm.n1738 4.60698
R48927 C9_P_btm.n1743 C9_P_btm.n1742 4.60698
R48928 C9_P_btm.n1742 C9_P_btm.n1741 4.60698
R48929 C9_P_btm.n1717 C9_P_btm.n1716 4.60698
R48930 C9_P_btm.n1718 C9_P_btm.n1717 4.60698
R48931 C9_P_btm.n1720 C9_P_btm.n1719 4.60698
R48932 C9_P_btm.n1721 C9_P_btm.n1720 4.60698
R48933 C9_P_btm.n1723 C9_P_btm.n1722 4.60698
R48934 C9_P_btm.n1724 C9_P_btm.n1723 4.60698
R48935 C9_P_btm.n1726 C9_P_btm.n1725 4.60698
R48936 C9_P_btm.n1727 C9_P_btm.n1726 4.60698
R48937 C9_P_btm.n101 C9_P_btm.n100 4.60698
R48938 C9_P_btm.n100 C9_P_btm.n91 4.60698
R48939 C9_P_btm.n98 C9_P_btm.n97 4.60698
R48940 C9_P_btm.n99 C9_P_btm.n98 4.60698
R48941 C9_P_btm.n95 C9_P_btm.n94 4.60698
R48942 C9_P_btm.n96 C9_P_btm.n95 4.60698
R48943 C9_P_btm.n1712 C9_P_btm.n1711 4.60698
R48944 C9_P_btm.n1711 C9_P_btm.n86 4.60698
R48945 C9_P_btm.n1706 C9_P_btm.n1705 4.60698
R48946 C9_P_btm.n1705 C9_P_btm.n1704 4.60698
R48947 C9_P_btm.n1703 C9_P_btm.n1702 4.60698
R48948 C9_P_btm.n1702 C9_P_btm.n1701 4.60698
R48949 C9_P_btm.n1700 C9_P_btm.n1699 4.60698
R48950 C9_P_btm.n1699 C9_P_btm.n1698 4.60698
R48951 C9_P_btm.n1697 C9_P_btm.n1696 4.60698
R48952 C9_P_btm.n1696 C9_P_btm.n1695 4.60698
R48953 C9_P_btm.n1689 C9_P_btm.n1688 4.60698
R48954 C9_P_btm.n1690 C9_P_btm.n1689 4.60698
R48955 C9_P_btm.n1686 C9_P_btm.n1685 4.60698
R48956 C9_P_btm.n1687 C9_P_btm.n1686 4.60698
R48957 C9_P_btm.n1683 C9_P_btm.n1682 4.60698
R48958 C9_P_btm.n1684 C9_P_btm.n1683 4.60698
R48959 C9_P_btm.n1680 C9_P_btm.n1679 4.60698
R48960 C9_P_btm.n1681 C9_P_btm.n1680 4.60698
R48961 C9_P_btm.n1675 C9_P_btm.n1674 4.60698
R48962 C9_P_btm.n1674 C9_P_btm.n109 4.60698
R48963 C9_P_btm.n118 C9_P_btm.n117 4.60698
R48964 C9_P_btm.n119 C9_P_btm.n118 4.60698
R48965 C9_P_btm.n121 C9_P_btm.n120 4.60698
R48966 C9_P_btm.n122 C9_P_btm.n121 4.60698
R48967 C9_P_btm.n124 C9_P_btm.n123 4.60698
R48968 C9_P_btm.n123 C9_P_btm.n114 4.60698
R48969 C9_P_btm.n1660 C9_P_btm.n1659 4.60698
R48970 C9_P_btm.n1659 C9_P_btm.n1658 4.60698
R48971 C9_P_btm.n1663 C9_P_btm.n1662 4.60698
R48972 C9_P_btm.n1662 C9_P_btm.n1661 4.60698
R48973 C9_P_btm.n1666 C9_P_btm.n1665 4.60698
R48974 C9_P_btm.n1665 C9_P_btm.n1664 4.60698
R48975 C9_P_btm.n1669 C9_P_btm.n1668 4.60698
R48976 C9_P_btm.n1668 C9_P_btm.n1667 4.60698
R48977 C9_P_btm.n1642 C9_P_btm.n1641 4.60698
R48978 C9_P_btm.n1643 C9_P_btm.n1642 4.60698
R48979 C9_P_btm.n1645 C9_P_btm.n1644 4.60698
R48980 C9_P_btm.n1646 C9_P_btm.n1645 4.60698
R48981 C9_P_btm.n1648 C9_P_btm.n1647 4.60698
R48982 C9_P_btm.n1649 C9_P_btm.n1648 4.60698
R48983 C9_P_btm.n1651 C9_P_btm.n1650 4.60698
R48984 C9_P_btm.n1652 C9_P_btm.n1651 4.60698
R48985 C9_P_btm.n1653 C9_P_btm.n128 4.60698
R48986 C9_P_btm.n1654 C9_P_btm.n1653 4.60698
R48987 C9_P_btm.n1384 C9_P_btm.n1383 4.60698
R48988 C9_P_btm.n1385 C9_P_btm.n1384 4.60698
R48989 C9_P_btm.n1381 C9_P_btm.n1380 4.60698
R48990 C9_P_btm.n1382 C9_P_btm.n1381 4.60698
R48991 C9_P_btm.n1378 C9_P_btm.n1377 4.60698
R48992 C9_P_btm.n1379 C9_P_btm.n1378 4.60698
R48993 C9_P_btm.n1375 C9_P_btm.n1374 4.60698
R48994 C9_P_btm.n1376 C9_P_btm.n1375 4.60698
R48995 C9_P_btm.n1372 C9_P_btm.n1371 4.60698
R48996 C9_P_btm.n1373 C9_P_btm.n1372 4.60698
R48997 C9_P_btm.n1369 C9_P_btm.n1368 4.60698
R48998 C9_P_btm.n1370 C9_P_btm.n1369 4.60698
R48999 C9_P_btm.n1366 C9_P_btm.n1365 4.60698
R49000 C9_P_btm.n1367 C9_P_btm.n1366 4.60698
R49001 C9_P_btm.n1363 C9_P_btm.n1362 4.60698
R49002 C9_P_btm.n1364 C9_P_btm.n1363 4.60698
R49003 C9_P_btm.n1360 C9_P_btm.n1359 4.60698
R49004 C9_P_btm.n1361 C9_P_btm.n1360 4.60698
R49005 C9_P_btm.n1357 C9_P_btm.n1356 4.60698
R49006 C9_P_btm.n1358 C9_P_btm.n1357 4.60698
R49007 C9_P_btm.n1354 C9_P_btm.n1353 4.60698
R49008 C9_P_btm.n1355 C9_P_btm.n1354 4.60698
R49009 C9_P_btm.n1351 C9_P_btm.n1350 4.60698
R49010 C9_P_btm.n1352 C9_P_btm.n1351 4.60698
R49011 C9_P_btm.n1348 C9_P_btm.n1347 4.60698
R49012 C9_P_btm.n1349 C9_P_btm.n1348 4.60698
R49013 C9_P_btm.n1444 C9_P_btm.n1443 4.60698
R49014 C9_P_btm.n1443 C9_P_btm.n1442 4.60698
R49015 C9_P_btm.n1440 C9_P_btm.n1439 4.60698
R49016 C9_P_btm.n1441 C9_P_btm.n1440 4.60698
R49017 C9_P_btm.n1437 C9_P_btm.n1436 4.60698
R49018 C9_P_btm.n1438 C9_P_btm.n1437 4.60698
R49019 C9_P_btm.n1434 C9_P_btm.n1433 4.60698
R49020 C9_P_btm.n1435 C9_P_btm.n1434 4.60698
R49021 C9_P_btm.n1431 C9_P_btm.n1430 4.60698
R49022 C9_P_btm.n1432 C9_P_btm.n1431 4.60698
R49023 C9_P_btm.n1428 C9_P_btm.n1427 4.60698
R49024 C9_P_btm.n1429 C9_P_btm.n1428 4.60698
R49025 C9_P_btm.n1425 C9_P_btm.n1424 4.60698
R49026 C9_P_btm.n1426 C9_P_btm.n1425 4.60698
R49027 C9_P_btm.n1422 C9_P_btm.n1421 4.60698
R49028 C9_P_btm.n1423 C9_P_btm.n1422 4.60698
R49029 C9_P_btm.n1419 C9_P_btm.n1418 4.60698
R49030 C9_P_btm.n1420 C9_P_btm.n1419 4.60698
R49031 C9_P_btm.n1416 C9_P_btm.n1415 4.60698
R49032 C9_P_btm.n1417 C9_P_btm.n1416 4.60698
R49033 C9_P_btm.n1413 C9_P_btm.n1412 4.60698
R49034 C9_P_btm.n1414 C9_P_btm.n1413 4.60698
R49035 C9_P_btm.n1410 C9_P_btm.n1409 4.60698
R49036 C9_P_btm.n1411 C9_P_btm.n1410 4.60698
R49037 C9_P_btm.n1407 C9_P_btm.n1406 4.60698
R49038 C9_P_btm.n1408 C9_P_btm.n1407 4.60698
R49039 C9_P_btm.n1404 C9_P_btm.n1403 4.60698
R49040 C9_P_btm.n1405 C9_P_btm.n1404 4.60698
R49041 C9_P_btm.n1401 C9_P_btm.n1400 4.60698
R49042 C9_P_btm.n1402 C9_P_btm.n1401 4.60698
R49043 C9_P_btm.n1398 C9_P_btm.n1397 4.60698
R49044 C9_P_btm.n1399 C9_P_btm.n1398 4.60698
R49045 C9_P_btm.n1395 C9_P_btm.n1394 4.60698
R49046 C9_P_btm.n1396 C9_P_btm.n1395 4.60698
R49047 C9_P_btm.n1392 C9_P_btm.n1391 4.60698
R49048 C9_P_btm.n1393 C9_P_btm.n1392 4.60698
R49049 C9_P_btm.n1637 C9_P_btm.n1636 4.60698
R49050 C9_P_btm.n1636 C9_P_btm.n133 4.60698
R49051 C9_P_btm.n1631 C9_P_btm.n1630 4.60698
R49052 C9_P_btm.n1630 C9_P_btm.n1629 4.60698
R49053 C9_P_btm.n1628 C9_P_btm.n1627 4.60698
R49054 C9_P_btm.n1627 C9_P_btm.n1626 4.60698
R49055 C9_P_btm.n1625 C9_P_btm.n1624 4.60698
R49056 C9_P_btm.n1624 C9_P_btm.n1623 4.60698
R49057 C9_P_btm.n1622 C9_P_btm.n1621 4.60698
R49058 C9_P_btm.n1621 C9_P_btm.n1620 4.60698
R49059 C9_P_btm.n1619 C9_P_btm.n1618 4.60698
R49060 C9_P_btm.n1618 C9_P_btm.n1617 4.60698
R49061 C9_P_btm.n1616 C9_P_btm.n1615 4.60698
R49062 C9_P_btm.n1615 C9_P_btm.n1614 4.60698
R49063 C9_P_btm.n1613 C9_P_btm.n1612 4.60698
R49064 C9_P_btm.n1612 C9_P_btm.n1611 4.60698
R49065 C9_P_btm.n1610 C9_P_btm.n1609 4.60698
R49066 C9_P_btm.n1609 C9_P_btm.n1608 4.60698
R49067 C9_P_btm.n1607 C9_P_btm.n1606 4.60698
R49068 C9_P_btm.n1606 C9_P_btm.n1605 4.60698
R49069 C9_P_btm.n1604 C9_P_btm.n1603 4.60698
R49070 C9_P_btm.n1603 C9_P_btm.n1602 4.60698
R49071 C9_P_btm.n1601 C9_P_btm.n1600 4.60698
R49072 C9_P_btm.n1600 C9_P_btm.n1599 4.60698
R49073 C9_P_btm.n1598 C9_P_btm.n1597 4.60698
R49074 C9_P_btm.n1597 C9_P_btm.n1596 4.60698
R49075 C9_P_btm.n1595 C9_P_btm.n1594 4.60698
R49076 C9_P_btm.n1594 C9_P_btm.n1593 4.60698
R49077 C9_P_btm.n1592 C9_P_btm.n1591 4.60698
R49078 C9_P_btm.n1591 C9_P_btm.n1590 4.60698
R49079 C9_P_btm.n1589 C9_P_btm.n1588 4.60698
R49080 C9_P_btm.n1588 C9_P_btm.n1587 4.60698
R49081 C9_P_btm.n1586 C9_P_btm.n1585 4.60698
R49082 C9_P_btm.n1585 C9_P_btm.n1584 4.60698
R49083 C9_P_btm.n1583 C9_P_btm.n1582 4.60698
R49084 C9_P_btm.n1582 C9_P_btm.n1581 4.60698
R49085 C9_P_btm.n1580 C9_P_btm.n1579 4.60698
R49086 C9_P_btm.n1579 C9_P_btm.n1578 4.60698
R49087 C9_P_btm.n1577 C9_P_btm.n1576 4.60698
R49088 C9_P_btm.n1576 C9_P_btm.n1575 4.60698
R49089 C9_P_btm.n1574 C9_P_btm.n1573 4.60698
R49090 C9_P_btm.n1573 C9_P_btm.n1572 4.60698
R49091 C9_P_btm.n1571 C9_P_btm.n1570 4.60698
R49092 C9_P_btm.n1570 C9_P_btm.n1569 4.60698
R49093 C9_P_btm.n1568 C9_P_btm.n1567 4.60698
R49094 C9_P_btm.n1567 C9_P_btm.n1566 4.60698
R49095 C9_P_btm.n1565 C9_P_btm.n1564 4.60698
R49096 C9_P_btm.n1564 C9_P_btm.n1563 4.60698
R49097 C9_P_btm.n1562 C9_P_btm.n1561 4.60698
R49098 C9_P_btm.n1561 C9_P_btm.n1560 4.60698
R49099 C9_P_btm.n1559 C9_P_btm.n1558 4.60698
R49100 C9_P_btm.n1558 C9_P_btm.n1557 4.60698
R49101 C9_P_btm.n1556 C9_P_btm.n1555 4.60698
R49102 C9_P_btm.n1555 C9_P_btm.n1554 4.60698
R49103 C9_P_btm.n1553 C9_P_btm.n1552 4.60698
R49104 C9_P_btm.n1552 C9_P_btm.n1551 4.60698
R49105 C9_P_btm.n1550 C9_P_btm.n1549 4.60698
R49106 C9_P_btm.n1549 C9_P_btm.n1548 4.60698
R49107 C9_P_btm.n1547 C9_P_btm.n1546 4.60698
R49108 C9_P_btm.n1546 C9_P_btm.n1545 4.60698
R49109 C9_P_btm.n1544 C9_P_btm.n1543 4.60698
R49110 C9_P_btm.n1543 C9_P_btm.n1542 4.60698
R49111 C9_P_btm.n1541 C9_P_btm.n1540 4.60698
R49112 C9_P_btm.n1540 C9_P_btm.n1539 4.60698
R49113 C9_P_btm.n1538 C9_P_btm.n1537 4.60698
R49114 C9_P_btm.n1537 C9_P_btm.n1536 4.60698
R49115 C9_P_btm.n1535 C9_P_btm.n1534 4.60698
R49116 C9_P_btm.n1534 C9_P_btm.n1533 4.60698
R49117 C9_P_btm.n1532 C9_P_btm.n1531 4.60698
R49118 C9_P_btm.n1531 C9_P_btm.n1530 4.60698
R49119 C9_P_btm.n1529 C9_P_btm.n1528 4.60698
R49120 C9_P_btm.n1528 C9_P_btm.n1527 4.60698
R49121 C9_P_btm.n1526 C9_P_btm.n1525 4.60698
R49122 C9_P_btm.n1525 C9_P_btm.n1524 4.60698
R49123 C9_P_btm.n1523 C9_P_btm.n1522 4.60698
R49124 C9_P_btm.n1522 C9_P_btm.n1521 4.60698
R49125 C9_P_btm.n1520 C9_P_btm.n1519 4.60698
R49126 C9_P_btm.n1519 C9_P_btm.n1518 4.60698
R49127 C9_P_btm.n1517 C9_P_btm.n1516 4.60698
R49128 C9_P_btm.n1516 C9_P_btm.n1515 4.60698
R49129 C9_P_btm.n1514 C9_P_btm.n1513 4.60698
R49130 C9_P_btm.n1513 C9_P_btm.n1512 4.60698
R49131 C9_P_btm.n1506 C9_P_btm.n1505 4.60698
R49132 C9_P_btm.n1507 C9_P_btm.n1506 4.60698
R49133 C9_P_btm.n1503 C9_P_btm.n1502 4.60698
R49134 C9_P_btm.n1504 C9_P_btm.n1503 4.60698
R49135 C9_P_btm.n1500 C9_P_btm.n1499 4.60698
R49136 C9_P_btm.n1501 C9_P_btm.n1500 4.60698
R49137 C9_P_btm.n1497 C9_P_btm.n1496 4.60698
R49138 C9_P_btm.n1498 C9_P_btm.n1497 4.60698
R49139 C9_P_btm.n1494 C9_P_btm.n1493 4.60698
R49140 C9_P_btm.n1495 C9_P_btm.n1494 4.60698
R49141 C9_P_btm.n1491 C9_P_btm.n1490 4.60698
R49142 C9_P_btm.n1492 C9_P_btm.n1491 4.60698
R49143 C9_P_btm.n1488 C9_P_btm.n1487 4.60698
R49144 C9_P_btm.n1489 C9_P_btm.n1488 4.60698
R49145 C9_P_btm.n1485 C9_P_btm.n1484 4.60698
R49146 C9_P_btm.n1486 C9_P_btm.n1485 4.60698
R49147 C9_P_btm.n1482 C9_P_btm.n1481 4.60698
R49148 C9_P_btm.n1483 C9_P_btm.n1482 4.60698
R49149 C9_P_btm.n1479 C9_P_btm.n1478 4.60698
R49150 C9_P_btm.n1480 C9_P_btm.n1479 4.60698
R49151 C9_P_btm.n1476 C9_P_btm.n1475 4.60698
R49152 C9_P_btm.n1477 C9_P_btm.n1476 4.60698
R49153 C9_P_btm.n1473 C9_P_btm.n1472 4.60698
R49154 C9_P_btm.n1474 C9_P_btm.n1473 4.60698
R49155 C9_P_btm.n1470 C9_P_btm.n1469 4.60698
R49156 C9_P_btm.n1471 C9_P_btm.n1470 4.60698
R49157 C9_P_btm.n1467 C9_P_btm.n1466 4.60698
R49158 C9_P_btm.n1468 C9_P_btm.n1467 4.60698
R49159 C9_P_btm.n1464 C9_P_btm.n1463 4.60698
R49160 C9_P_btm.n1465 C9_P_btm.n1464 4.60698
R49161 C9_P_btm.n1461 C9_P_btm.n1460 4.60698
R49162 C9_P_btm.n1462 C9_P_btm.n1461 4.60698
R49163 C9_P_btm.n1458 C9_P_btm.n1457 4.60698
R49164 C9_P_btm.n1459 C9_P_btm.n1458 4.60698
R49165 C9_P_btm.n1455 C9_P_btm.n1454 4.60698
R49166 C9_P_btm.n1456 C9_P_btm.n1455 4.60698
R49167 C9_P_btm.n1452 C9_P_btm.n1451 4.60698
R49168 C9_P_btm.n1453 C9_P_btm.n1452 4.60698
R49169 C9_P_btm.n1315 C9_P_btm.n1314 4.60698
R49170 C9_P_btm.n1316 C9_P_btm.n1315 4.60698
R49171 C9_P_btm.n1312 C9_P_btm.n1311 4.60698
R49172 C9_P_btm.n1313 C9_P_btm.n1312 4.60698
R49173 C9_P_btm.n1309 C9_P_btm.n1308 4.60698
R49174 C9_P_btm.n1310 C9_P_btm.n1309 4.60698
R49175 C9_P_btm.n1306 C9_P_btm.n1305 4.60698
R49176 C9_P_btm.n1307 C9_P_btm.n1306 4.60698
R49177 C9_P_btm.n1303 C9_P_btm.n1302 4.60698
R49178 C9_P_btm.n1304 C9_P_btm.n1303 4.60698
R49179 C9_P_btm.n1300 C9_P_btm.n1299 4.60698
R49180 C9_P_btm.n1301 C9_P_btm.n1300 4.60698
R49181 C9_P_btm.n1297 C9_P_btm.n1296 4.60698
R49182 C9_P_btm.n1298 C9_P_btm.n1297 4.60698
R49183 C9_P_btm.n1294 C9_P_btm.n1293 4.60698
R49184 C9_P_btm.n1295 C9_P_btm.n1294 4.60698
R49185 C9_P_btm.n1291 C9_P_btm.n1290 4.60698
R49186 C9_P_btm.n1292 C9_P_btm.n1291 4.60698
R49187 C9_P_btm.n1288 C9_P_btm.n1287 4.60698
R49188 C9_P_btm.n1289 C9_P_btm.n1288 4.60698
R49189 C9_P_btm.n1285 C9_P_btm.n1284 4.60698
R49190 C9_P_btm.n1286 C9_P_btm.n1285 4.60698
R49191 C9_P_btm.n1282 C9_P_btm.n1281 4.60698
R49192 C9_P_btm.n1283 C9_P_btm.n1282 4.60698
R49193 C9_P_btm.n1279 C9_P_btm.n1278 4.60698
R49194 C9_P_btm.n1280 C9_P_btm.n1279 4.60698
R49195 C9_P_btm.n1277 C9_P_btm.n1276 4.60698
R49196 C9_P_btm.n1276 C9_P_btm.n1275 4.60698
R49197 C9_P_btm.n1274 C9_P_btm.n1273 4.60698
R49198 C9_P_btm.n1273 C9_P_btm.n1272 4.60698
R49199 C9_P_btm.n1271 C9_P_btm.n1270 4.60698
R49200 C9_P_btm.n1270 C9_P_btm.n1269 4.60698
R49201 C9_P_btm.n1268 C9_P_btm.n1267 4.60698
R49202 C9_P_btm.n1267 C9_P_btm.n1266 4.60698
R49203 C9_P_btm.n1265 C9_P_btm.n1264 4.60698
R49204 C9_P_btm.n1264 C9_P_btm.n1263 4.60698
R49205 C9_P_btm.n1259 C9_P_btm.n1258 4.60698
R49206 C9_P_btm.n1258 C9_P_btm.n922 4.60698
R49207 C9_P_btm.n1256 C9_P_btm.n1255 4.60698
R49208 C9_P_btm.n1257 C9_P_btm.n1256 4.60698
R49209 C9_P_btm.n1253 C9_P_btm.n1252 4.60698
R49210 C9_P_btm.n1254 C9_P_btm.n1253 4.60698
R49211 C9_P_btm.n1250 C9_P_btm.n1249 4.60698
R49212 C9_P_btm.n1251 C9_P_btm.n1250 4.60698
R49213 C9_P_btm.n1244 C9_P_btm.n1243 4.60698
R49214 C9_P_btm.n1243 C9_P_btm.n1242 4.60698
R49215 C9_P_btm.n1241 C9_P_btm.n1240 4.60698
R49216 C9_P_btm.n1240 C9_P_btm.n1239 4.60698
R49217 C9_P_btm.n1238 C9_P_btm.n1237 4.60698
R49218 C9_P_btm.n1237 C9_P_btm.n1236 4.60698
R49219 C9_P_btm.n1235 C9_P_btm.n1234 4.60698
R49220 C9_P_btm.n1234 C9_P_btm.n1233 4.60698
R49221 C9_P_btm.n1227 C9_P_btm.n1226 4.60698
R49222 C9_P_btm.n1228 C9_P_btm.n1227 4.60698
R49223 C9_P_btm.n1224 C9_P_btm.n1223 4.60698
R49224 C9_P_btm.n1225 C9_P_btm.n1224 4.60698
R49225 C9_P_btm.n1221 C9_P_btm.n1220 4.60698
R49226 C9_P_btm.n1222 C9_P_btm.n1221 4.60698
R49227 C9_P_btm.n1218 C9_P_btm.n1217 4.60698
R49228 C9_P_btm.n1219 C9_P_btm.n1218 4.60698
R49229 C9_P_btm.n1213 C9_P_btm.n1212 4.60698
R49230 C9_P_btm.n1212 C9_P_btm.n937 4.60698
R49231 C9_P_btm.n946 C9_P_btm.n945 4.60698
R49232 C9_P_btm.n947 C9_P_btm.n946 4.60698
R49233 C9_P_btm.n949 C9_P_btm.n948 4.60698
R49234 C9_P_btm.n950 C9_P_btm.n949 4.60698
R49235 C9_P_btm.n952 C9_P_btm.n951 4.60698
R49236 C9_P_btm.n951 C9_P_btm.n942 4.60698
R49237 C9_P_btm.n1198 C9_P_btm.n1197 4.60698
R49238 C9_P_btm.n1197 C9_P_btm.n1196 4.60698
R49239 C9_P_btm.n1201 C9_P_btm.n1200 4.60698
R49240 C9_P_btm.n1200 C9_P_btm.n1199 4.60698
R49241 C9_P_btm.n1204 C9_P_btm.n1203 4.60698
R49242 C9_P_btm.n1203 C9_P_btm.n1202 4.60698
R49243 C9_P_btm.n1207 C9_P_btm.n1206 4.60698
R49244 C9_P_btm.n1206 C9_P_btm.n1205 4.60698
R49245 C9_P_btm.n1181 C9_P_btm.n1180 4.60698
R49246 C9_P_btm.n1182 C9_P_btm.n1181 4.60698
R49247 C9_P_btm.n1184 C9_P_btm.n1183 4.60698
R49248 C9_P_btm.n1185 C9_P_btm.n1184 4.60698
R49249 C9_P_btm.n1187 C9_P_btm.n1186 4.60698
R49250 C9_P_btm.n1188 C9_P_btm.n1187 4.60698
R49251 C9_P_btm.n1190 C9_P_btm.n1189 4.60698
R49252 C9_P_btm.n1191 C9_P_btm.n1190 4.60698
R49253 C9_P_btm.n975 C9_P_btm.n974 4.60698
R49254 C9_P_btm.n974 C9_P_btm.n965 4.60698
R49255 C9_P_btm.n972 C9_P_btm.n971 4.60698
R49256 C9_P_btm.n973 C9_P_btm.n972 4.60698
R49257 C9_P_btm.n969 C9_P_btm.n968 4.60698
R49258 C9_P_btm.n970 C9_P_btm.n969 4.60698
R49259 C9_P_btm.n1176 C9_P_btm.n1175 4.60698
R49260 C9_P_btm.n1175 C9_P_btm.n960 4.60698
R49261 C9_P_btm.n1170 C9_P_btm.n1169 4.60698
R49262 C9_P_btm.n1169 C9_P_btm.n1168 4.60698
R49263 C9_P_btm.n1167 C9_P_btm.n1166 4.60698
R49264 C9_P_btm.n1166 C9_P_btm.n1165 4.60698
R49265 C9_P_btm.n1164 C9_P_btm.n1163 4.60698
R49266 C9_P_btm.n1163 C9_P_btm.n1162 4.60698
R49267 C9_P_btm.n1161 C9_P_btm.n1160 4.60698
R49268 C9_P_btm.n1160 C9_P_btm.n1159 4.60698
R49269 C9_P_btm.n1153 C9_P_btm.n1152 4.60698
R49270 C9_P_btm.n1154 C9_P_btm.n1153 4.60698
R49271 C9_P_btm.n1150 C9_P_btm.n1149 4.60698
R49272 C9_P_btm.n1151 C9_P_btm.n1150 4.60698
R49273 C9_P_btm.n1147 C9_P_btm.n1146 4.60698
R49274 C9_P_btm.n1148 C9_P_btm.n1147 4.60698
R49275 C9_P_btm.n1144 C9_P_btm.n1143 4.60698
R49276 C9_P_btm.n1145 C9_P_btm.n1144 4.60698
R49277 C9_P_btm.n1139 C9_P_btm.n1138 4.60698
R49278 C9_P_btm.n1138 C9_P_btm.n983 4.60698
R49279 C9_P_btm.n992 C9_P_btm.n991 4.60698
R49280 C9_P_btm.n993 C9_P_btm.n992 4.60698
R49281 C9_P_btm.n995 C9_P_btm.n994 4.60698
R49282 C9_P_btm.n996 C9_P_btm.n995 4.60698
R49283 C9_P_btm.n998 C9_P_btm.n997 4.60698
R49284 C9_P_btm.n997 C9_P_btm.n988 4.60698
R49285 C9_P_btm.n1124 C9_P_btm.n1123 4.60698
R49286 C9_P_btm.n1123 C9_P_btm.n1122 4.60698
R49287 C9_P_btm.n1127 C9_P_btm.n1126 4.60698
R49288 C9_P_btm.n1126 C9_P_btm.n1125 4.60698
R49289 C9_P_btm.n1130 C9_P_btm.n1129 4.60698
R49290 C9_P_btm.n1129 C9_P_btm.n1128 4.60698
R49291 C9_P_btm.n1133 C9_P_btm.n1132 4.60698
R49292 C9_P_btm.n1132 C9_P_btm.n1131 4.60698
R49293 C9_P_btm.n1107 C9_P_btm.n1106 4.60698
R49294 C9_P_btm.n1108 C9_P_btm.n1107 4.60698
R49295 C9_P_btm.n1110 C9_P_btm.n1109 4.60698
R49296 C9_P_btm.n1111 C9_P_btm.n1110 4.60698
R49297 C9_P_btm.n1113 C9_P_btm.n1112 4.60698
R49298 C9_P_btm.n1114 C9_P_btm.n1113 4.60698
R49299 C9_P_btm.n1116 C9_P_btm.n1115 4.60698
R49300 C9_P_btm.n1117 C9_P_btm.n1116 4.60698
R49301 C9_P_btm.n1021 C9_P_btm.n1020 4.60698
R49302 C9_P_btm.n1020 C9_P_btm.n1011 4.60698
R49303 C9_P_btm.n1018 C9_P_btm.n1017 4.60698
R49304 C9_P_btm.n1019 C9_P_btm.n1018 4.60698
R49305 C9_P_btm.n1015 C9_P_btm.n1014 4.60698
R49306 C9_P_btm.n1016 C9_P_btm.n1015 4.60698
R49307 C9_P_btm.n1102 C9_P_btm.n1101 4.60698
R49308 C9_P_btm.n1101 C9_P_btm.n1006 4.60698
R49309 C9_P_btm.n1096 C9_P_btm.n1095 4.60698
R49310 C9_P_btm.n1095 C9_P_btm.n1094 4.60698
R49311 C9_P_btm.n1093 C9_P_btm.n1092 4.60698
R49312 C9_P_btm.n1092 C9_P_btm.n1091 4.60698
R49313 C9_P_btm.n1090 C9_P_btm.n1089 4.60698
R49314 C9_P_btm.n1089 C9_P_btm.n1088 4.60698
R49315 C9_P_btm.n1087 C9_P_btm.n1086 4.60698
R49316 C9_P_btm.n1086 C9_P_btm.n1085 4.60698
R49317 C9_P_btm.n1079 C9_P_btm.n1078 4.60698
R49318 C9_P_btm.n1080 C9_P_btm.n1079 4.60698
R49319 C9_P_btm.n1076 C9_P_btm.n1075 4.60698
R49320 C9_P_btm.n1077 C9_P_btm.n1076 4.60698
R49321 C9_P_btm.n1073 C9_P_btm.n1072 4.60698
R49322 C9_P_btm.n1074 C9_P_btm.n1073 4.60698
R49323 C9_P_btm.n1070 C9_P_btm.n1069 4.60698
R49324 C9_P_btm.n1071 C9_P_btm.n1070 4.60698
R49325 C9_P_btm.n1065 C9_P_btm.n1064 4.60698
R49326 C9_P_btm.n1064 C9_P_btm.n1029 4.60698
R49327 C9_P_btm.n1037 C9_P_btm.n1036 4.60698
R49328 C9_P_btm.n1038 C9_P_btm.n1037 4.60698
R49329 C9_P_btm.n1040 C9_P_btm.n1039 4.60698
R49330 C9_P_btm.n1041 C9_P_btm.n1040 4.60698
R49331 C9_P_btm.n1043 C9_P_btm.n1042 4.60698
R49332 C9_P_btm.n1042 C9_P_btm.n1033 4.60698
R49333 C9_P_btm.n1049 C9_P_btm.n1048 4.60698
R49334 C9_P_btm.n1050 C9_P_btm.n1049 4.60698
R49335 C9_P_btm.n1052 C9_P_btm.n1051 4.60698
R49336 C9_P_btm.n1053 C9_P_btm.n1052 4.60698
R49337 C9_P_btm.n1055 C9_P_btm.n1054 4.60698
R49338 C9_P_btm.n1056 C9_P_btm.n1055 4.60698
R49339 C9_P_btm.n1058 C9_P_btm.n1057 4.60698
R49340 C9_P_btm.n1059 C9_P_btm.n1058 4.60698
R49341 C9_P_btm.n1450 C9_P_btm.n1449 4.60698
R49342 C9_P_btm.n1449 C9_P_btm.n1448 4.60698
R49343 C9_P_btm.n1447 C9_P_btm.n1446 4.60698
R49344 C9_P_btm.n1446 C9_P_btm.n1445 4.60698
R49345 C9_P_btm.n881 C9_P_btm.n880 4.60698
R49346 C9_P_btm.n882 C9_P_btm.n881 4.60698
R49347 C9_P_btm.n878 C9_P_btm.n877 4.60698
R49348 C9_P_btm.n879 C9_P_btm.n878 4.60698
R49349 C9_P_btm.n875 C9_P_btm.n874 4.60698
R49350 C9_P_btm.n876 C9_P_btm.n875 4.60698
R49351 C9_P_btm.n872 C9_P_btm.n871 4.60698
R49352 C9_P_btm.n873 C9_P_btm.n872 4.60698
R49353 C9_P_btm.n869 C9_P_btm.n868 4.60698
R49354 C9_P_btm.n870 C9_P_btm.n869 4.60698
R49355 C9_P_btm.n866 C9_P_btm.n865 4.60698
R49356 C9_P_btm.n867 C9_P_btm.n866 4.60698
R49357 C9_P_btm.n863 C9_P_btm.n862 4.60698
R49358 C9_P_btm.n864 C9_P_btm.n863 4.60698
R49359 C9_P_btm.n860 C9_P_btm.n859 4.60698
R49360 C9_P_btm.n861 C9_P_btm.n860 4.60698
R49361 C9_P_btm.n857 C9_P_btm.n856 4.60698
R49362 C9_P_btm.n858 C9_P_btm.n857 4.60698
R49363 C9_P_btm.n854 C9_P_btm.n853 4.60698
R49364 C9_P_btm.n855 C9_P_btm.n854 4.60698
R49365 C9_P_btm.n851 C9_P_btm.n850 4.60698
R49366 C9_P_btm.n852 C9_P_btm.n851 4.60698
R49367 C9_P_btm.n848 C9_P_btm.n847 4.60698
R49368 C9_P_btm.n849 C9_P_btm.n848 4.60698
R49369 C9_P_btm.n845 C9_P_btm.n844 4.60698
R49370 C9_P_btm.n846 C9_P_btm.n845 4.60698
R49371 C9_P_btm.n842 C9_P_btm.n841 4.60698
R49372 C9_P_btm.n843 C9_P_btm.n842 4.60698
R49373 C9_P_btm.n839 C9_P_btm.n838 4.60698
R49374 C9_P_btm.n840 C9_P_btm.n839 4.60698
R49375 C9_P_btm.n836 C9_P_btm.n835 4.60698
R49376 C9_P_btm.n837 C9_P_btm.n836 4.60698
R49377 C9_P_btm.n833 C9_P_btm.n832 4.60698
R49378 C9_P_btm.n834 C9_P_btm.n833 4.60698
R49379 C9_P_btm.n830 C9_P_btm.n829 4.60698
R49380 C9_P_btm.n831 C9_P_btm.n830 4.60698
R49381 C9_P_btm.n827 C9_P_btm.n826 4.60698
R49382 C9_P_btm.n828 C9_P_btm.n827 4.60698
R49383 C9_P_btm.n824 C9_P_btm.n823 4.60698
R49384 C9_P_btm.n825 C9_P_btm.n824 4.60698
R49385 C9_P_btm.n821 C9_P_btm.n820 4.60698
R49386 C9_P_btm.n822 C9_P_btm.n821 4.60698
R49387 C9_P_btm.n818 C9_P_btm.n817 4.60698
R49388 C9_P_btm.n819 C9_P_btm.n818 4.60698
R49389 C9_P_btm.n815 C9_P_btm.n814 4.60698
R49390 C9_P_btm.n816 C9_P_btm.n815 4.60698
R49391 C9_P_btm.n812 C9_P_btm.n811 4.60698
R49392 C9_P_btm.n813 C9_P_btm.n812 4.60698
R49393 C9_P_btm.n809 C9_P_btm.n808 4.60698
R49394 C9_P_btm.n810 C9_P_btm.n809 4.60698
R49395 C9_P_btm.n806 C9_P_btm.n805 4.60698
R49396 C9_P_btm.n807 C9_P_btm.n806 4.60698
R49397 C9_P_btm.n803 C9_P_btm.n802 4.60698
R49398 C9_P_btm.n804 C9_P_btm.n803 4.60698
R49399 C9_P_btm.n800 C9_P_btm.n799 4.60698
R49400 C9_P_btm.n801 C9_P_btm.n800 4.60698
R49401 C9_P_btm.n797 C9_P_btm.n796 4.60698
R49402 C9_P_btm.n798 C9_P_btm.n797 4.60698
R49403 C9_P_btm.n794 C9_P_btm.n793 4.60698
R49404 C9_P_btm.n795 C9_P_btm.n794 4.60698
R49405 C9_P_btm.n791 C9_P_btm.n790 4.60698
R49406 C9_P_btm.n792 C9_P_btm.n791 4.60698
R49407 C9_P_btm.n788 C9_P_btm.n787 4.60698
R49408 C9_P_btm.n789 C9_P_btm.n788 4.60698
R49409 C9_P_btm.n785 C9_P_btm.n784 4.60698
R49410 C9_P_btm.n786 C9_P_btm.n785 4.60698
R49411 C9_P_btm.n782 C9_P_btm.n781 4.60698
R49412 C9_P_btm.n783 C9_P_btm.n782 4.60698
R49413 C9_P_btm.n779 C9_P_btm.n778 4.60698
R49414 C9_P_btm.n780 C9_P_btm.n779 4.60698
R49415 C9_P_btm.n776 C9_P_btm.n775 4.60698
R49416 C9_P_btm.n777 C9_P_btm.n776 4.60698
R49417 C9_P_btm.n773 C9_P_btm.n772 4.60698
R49418 C9_P_btm.n774 C9_P_btm.n773 4.60698
R49419 C9_P_btm.n770 C9_P_btm.n769 4.60698
R49420 C9_P_btm.n771 C9_P_btm.n770 4.60698
R49421 C9_P_btm.n767 C9_P_btm.n766 4.60698
R49422 C9_P_btm.n768 C9_P_btm.n767 4.60698
R49423 C9_P_btm.n764 C9_P_btm.n763 4.60698
R49424 C9_P_btm.n765 C9_P_btm.n764 4.60698
R49425 C9_P_btm.n759 C9_P_btm.n758 4.60698
R49426 C9_P_btm.n758 C9_P_btm.n215 4.60698
R49427 C9_P_btm.n296 C9_P_btm.n295 4.60698
R49428 C9_P_btm.n297 C9_P_btm.n296 4.60698
R49429 C9_P_btm.n299 C9_P_btm.n298 4.60698
R49430 C9_P_btm.n300 C9_P_btm.n299 4.60698
R49431 C9_P_btm.n302 C9_P_btm.n301 4.60698
R49432 C9_P_btm.n303 C9_P_btm.n302 4.60698
R49433 C9_P_btm.n305 C9_P_btm.n304 4.60698
R49434 C9_P_btm.n306 C9_P_btm.n305 4.60698
R49435 C9_P_btm.n308 C9_P_btm.n307 4.60698
R49436 C9_P_btm.n309 C9_P_btm.n308 4.60698
R49437 C9_P_btm.n311 C9_P_btm.n310 4.60698
R49438 C9_P_btm.n312 C9_P_btm.n311 4.60698
R49439 C9_P_btm.n314 C9_P_btm.n313 4.60698
R49440 C9_P_btm.n315 C9_P_btm.n314 4.60698
R49441 C9_P_btm.n317 C9_P_btm.n316 4.60698
R49442 C9_P_btm.n318 C9_P_btm.n317 4.60698
R49443 C9_P_btm.n320 C9_P_btm.n319 4.60698
R49444 C9_P_btm.n321 C9_P_btm.n320 4.60698
R49445 C9_P_btm.n323 C9_P_btm.n322 4.60698
R49446 C9_P_btm.n324 C9_P_btm.n323 4.60698
R49447 C9_P_btm.n326 C9_P_btm.n325 4.60698
R49448 C9_P_btm.n327 C9_P_btm.n326 4.60698
R49449 C9_P_btm.n329 C9_P_btm.n328 4.60698
R49450 C9_P_btm.n330 C9_P_btm.n329 4.60698
R49451 C9_P_btm.n332 C9_P_btm.n331 4.60698
R49452 C9_P_btm.n333 C9_P_btm.n332 4.60698
R49453 C9_P_btm.n335 C9_P_btm.n334 4.60698
R49454 C9_P_btm.n336 C9_P_btm.n335 4.60698
R49455 C9_P_btm.n338 C9_P_btm.n337 4.60698
R49456 C9_P_btm.n339 C9_P_btm.n338 4.60698
R49457 C9_P_btm.n341 C9_P_btm.n340 4.60698
R49458 C9_P_btm.n342 C9_P_btm.n341 4.60698
R49459 C9_P_btm.n344 C9_P_btm.n343 4.60698
R49460 C9_P_btm.n345 C9_P_btm.n344 4.60698
R49461 C9_P_btm.n347 C9_P_btm.n346 4.60698
R49462 C9_P_btm.n348 C9_P_btm.n347 4.60698
R49463 C9_P_btm.n350 C9_P_btm.n349 4.60698
R49464 C9_P_btm.n351 C9_P_btm.n350 4.60698
R49465 C9_P_btm.n353 C9_P_btm.n352 4.60698
R49466 C9_P_btm.n354 C9_P_btm.n353 4.60698
R49467 C9_P_btm.n356 C9_P_btm.n355 4.60698
R49468 C9_P_btm.n357 C9_P_btm.n356 4.60698
R49469 C9_P_btm.n359 C9_P_btm.n358 4.60698
R49470 C9_P_btm.n360 C9_P_btm.n359 4.60698
R49471 C9_P_btm.n362 C9_P_btm.n361 4.60698
R49472 C9_P_btm.n363 C9_P_btm.n362 4.60698
R49473 C9_P_btm.n365 C9_P_btm.n364 4.60698
R49474 C9_P_btm.n366 C9_P_btm.n365 4.60698
R49475 C9_P_btm.n368 C9_P_btm.n367 4.60698
R49476 C9_P_btm.n369 C9_P_btm.n368 4.60698
R49477 C9_P_btm.n371 C9_P_btm.n370 4.60698
R49478 C9_P_btm.n372 C9_P_btm.n371 4.60698
R49479 C9_P_btm.n374 C9_P_btm.n373 4.60698
R49480 C9_P_btm.n375 C9_P_btm.n374 4.60698
R49481 C9_P_btm.n377 C9_P_btm.n376 4.60698
R49482 C9_P_btm.n378 C9_P_btm.n377 4.60698
R49483 C9_P_btm.n380 C9_P_btm.n379 4.60698
R49484 C9_P_btm.n381 C9_P_btm.n380 4.60698
R49485 C9_P_btm.n383 C9_P_btm.n382 4.60698
R49486 C9_P_btm.n384 C9_P_btm.n383 4.60698
R49487 C9_P_btm.n386 C9_P_btm.n385 4.60698
R49488 C9_P_btm.n387 C9_P_btm.n386 4.60698
R49489 C9_P_btm.n389 C9_P_btm.n388 4.60698
R49490 C9_P_btm.n390 C9_P_btm.n389 4.60698
R49491 C9_P_btm.n392 C9_P_btm.n391 4.60698
R49492 C9_P_btm.n393 C9_P_btm.n392 4.60698
R49493 C9_P_btm.n395 C9_P_btm.n394 4.60698
R49494 C9_P_btm.n396 C9_P_btm.n395 4.60698
R49495 C9_P_btm.n398 C9_P_btm.n397 4.60698
R49496 C9_P_btm.n399 C9_P_btm.n398 4.60698
R49497 C9_P_btm.n401 C9_P_btm.n400 4.60698
R49498 C9_P_btm.n402 C9_P_btm.n401 4.60698
R49499 C9_P_btm.n404 C9_P_btm.n403 4.60698
R49500 C9_P_btm.n405 C9_P_btm.n404 4.60698
R49501 C9_P_btm.n407 C9_P_btm.n406 4.60698
R49502 C9_P_btm.n408 C9_P_btm.n407 4.60698
R49503 C9_P_btm.n410 C9_P_btm.n409 4.60698
R49504 C9_P_btm.n409 C9_P_btm.n256 4.60698
R49505 C9_P_btm.n636 C9_P_btm.n635 4.60698
R49506 C9_P_btm.n635 C9_P_btm.n634 4.60698
R49507 C9_P_btm.n639 C9_P_btm.n638 4.60698
R49508 C9_P_btm.n638 C9_P_btm.n637 4.60698
R49509 C9_P_btm.n642 C9_P_btm.n641 4.60698
R49510 C9_P_btm.n641 C9_P_btm.n640 4.60698
R49511 C9_P_btm.n645 C9_P_btm.n644 4.60698
R49512 C9_P_btm.n644 C9_P_btm.n643 4.60698
R49513 C9_P_btm.n648 C9_P_btm.n647 4.60698
R49514 C9_P_btm.n647 C9_P_btm.n646 4.60698
R49515 C9_P_btm.n651 C9_P_btm.n650 4.60698
R49516 C9_P_btm.n650 C9_P_btm.n649 4.60698
R49517 C9_P_btm.n654 C9_P_btm.n653 4.60698
R49518 C9_P_btm.n653 C9_P_btm.n652 4.60698
R49519 C9_P_btm.n657 C9_P_btm.n656 4.60698
R49520 C9_P_btm.n656 C9_P_btm.n655 4.60698
R49521 C9_P_btm.n660 C9_P_btm.n659 4.60698
R49522 C9_P_btm.n659 C9_P_btm.n658 4.60698
R49523 C9_P_btm.n663 C9_P_btm.n662 4.60698
R49524 C9_P_btm.n662 C9_P_btm.n661 4.60698
R49525 C9_P_btm.n666 C9_P_btm.n665 4.60698
R49526 C9_P_btm.n665 C9_P_btm.n664 4.60698
R49527 C9_P_btm.n669 C9_P_btm.n668 4.60698
R49528 C9_P_btm.n668 C9_P_btm.n667 4.60698
R49529 C9_P_btm.n672 C9_P_btm.n671 4.60698
R49530 C9_P_btm.n671 C9_P_btm.n670 4.60698
R49531 C9_P_btm.n675 C9_P_btm.n674 4.60698
R49532 C9_P_btm.n674 C9_P_btm.n673 4.60698
R49533 C9_P_btm.n678 C9_P_btm.n677 4.60698
R49534 C9_P_btm.n677 C9_P_btm.n676 4.60698
R49535 C9_P_btm.n681 C9_P_btm.n680 4.60698
R49536 C9_P_btm.n680 C9_P_btm.n679 4.60698
R49537 C9_P_btm.n684 C9_P_btm.n683 4.60698
R49538 C9_P_btm.n683 C9_P_btm.n682 4.60698
R49539 C9_P_btm.n687 C9_P_btm.n686 4.60698
R49540 C9_P_btm.n686 C9_P_btm.n685 4.60698
R49541 C9_P_btm.n690 C9_P_btm.n689 4.60698
R49542 C9_P_btm.n689 C9_P_btm.n688 4.60698
R49543 C9_P_btm.n693 C9_P_btm.n692 4.60698
R49544 C9_P_btm.n692 C9_P_btm.n691 4.60698
R49545 C9_P_btm.n696 C9_P_btm.n695 4.60698
R49546 C9_P_btm.n695 C9_P_btm.n694 4.60698
R49547 C9_P_btm.n699 C9_P_btm.n698 4.60698
R49548 C9_P_btm.n698 C9_P_btm.n697 4.60698
R49549 C9_P_btm.n702 C9_P_btm.n701 4.60698
R49550 C9_P_btm.n701 C9_P_btm.n700 4.60698
R49551 C9_P_btm.n705 C9_P_btm.n704 4.60698
R49552 C9_P_btm.n704 C9_P_btm.n703 4.60698
R49553 C9_P_btm.n708 C9_P_btm.n707 4.60698
R49554 C9_P_btm.n707 C9_P_btm.n706 4.60698
R49555 C9_P_btm.n711 C9_P_btm.n710 4.60698
R49556 C9_P_btm.n710 C9_P_btm.n709 4.60698
R49557 C9_P_btm.n714 C9_P_btm.n713 4.60698
R49558 C9_P_btm.n713 C9_P_btm.n712 4.60698
R49559 C9_P_btm.n717 C9_P_btm.n716 4.60698
R49560 C9_P_btm.n716 C9_P_btm.n715 4.60698
R49561 C9_P_btm.n720 C9_P_btm.n719 4.60698
R49562 C9_P_btm.n719 C9_P_btm.n718 4.60698
R49563 C9_P_btm.n723 C9_P_btm.n722 4.60698
R49564 C9_P_btm.n722 C9_P_btm.n721 4.60698
R49565 C9_P_btm.n726 C9_P_btm.n725 4.60698
R49566 C9_P_btm.n725 C9_P_btm.n724 4.60698
R49567 C9_P_btm.n729 C9_P_btm.n728 4.60698
R49568 C9_P_btm.n728 C9_P_btm.n727 4.60698
R49569 C9_P_btm.n732 C9_P_btm.n731 4.60698
R49570 C9_P_btm.n731 C9_P_btm.n730 4.60698
R49571 C9_P_btm.n735 C9_P_btm.n734 4.60698
R49572 C9_P_btm.n734 C9_P_btm.n733 4.60698
R49573 C9_P_btm.n738 C9_P_btm.n737 4.60698
R49574 C9_P_btm.n737 C9_P_btm.n736 4.60698
R49575 C9_P_btm.n741 C9_P_btm.n740 4.60698
R49576 C9_P_btm.n740 C9_P_btm.n739 4.60698
R49577 C9_P_btm.n744 C9_P_btm.n743 4.60698
R49578 C9_P_btm.n743 C9_P_btm.n742 4.60698
R49579 C9_P_btm.n747 C9_P_btm.n746 4.60698
R49580 C9_P_btm.n746 C9_P_btm.n745 4.60698
R49581 C9_P_btm.n750 C9_P_btm.n749 4.60698
R49582 C9_P_btm.n749 C9_P_btm.n748 4.60698
R49583 C9_P_btm.n753 C9_P_btm.n752 4.60698
R49584 C9_P_btm.n752 C9_P_btm.n751 4.60698
R49585 C9_P_btm.n512 C9_P_btm.n511 4.60698
R49586 C9_P_btm.n513 C9_P_btm.n512 4.60698
R49587 C9_P_btm.n515 C9_P_btm.n514 4.60698
R49588 C9_P_btm.n516 C9_P_btm.n515 4.60698
R49589 C9_P_btm.n518 C9_P_btm.n517 4.60698
R49590 C9_P_btm.n519 C9_P_btm.n518 4.60698
R49591 C9_P_btm.n521 C9_P_btm.n520 4.60698
R49592 C9_P_btm.n522 C9_P_btm.n521 4.60698
R49593 C9_P_btm.n524 C9_P_btm.n523 4.60698
R49594 C9_P_btm.n525 C9_P_btm.n524 4.60698
R49595 C9_P_btm.n527 C9_P_btm.n526 4.60698
R49596 C9_P_btm.n528 C9_P_btm.n527 4.60698
R49597 C9_P_btm.n530 C9_P_btm.n529 4.60698
R49598 C9_P_btm.n531 C9_P_btm.n530 4.60698
R49599 C9_P_btm.n533 C9_P_btm.n532 4.60698
R49600 C9_P_btm.n534 C9_P_btm.n533 4.60698
R49601 C9_P_btm.n536 C9_P_btm.n535 4.60698
R49602 C9_P_btm.n537 C9_P_btm.n536 4.60698
R49603 C9_P_btm.n539 C9_P_btm.n538 4.60698
R49604 C9_P_btm.n540 C9_P_btm.n539 4.60698
R49605 C9_P_btm.n542 C9_P_btm.n541 4.60698
R49606 C9_P_btm.n543 C9_P_btm.n542 4.60698
R49607 C9_P_btm.n545 C9_P_btm.n544 4.60698
R49608 C9_P_btm.n546 C9_P_btm.n545 4.60698
R49609 C9_P_btm.n548 C9_P_btm.n547 4.60698
R49610 C9_P_btm.n549 C9_P_btm.n548 4.60698
R49611 C9_P_btm.n551 C9_P_btm.n550 4.60698
R49612 C9_P_btm.n552 C9_P_btm.n551 4.60698
R49613 C9_P_btm.n554 C9_P_btm.n553 4.60698
R49614 C9_P_btm.n555 C9_P_btm.n554 4.60698
R49615 C9_P_btm.n557 C9_P_btm.n556 4.60698
R49616 C9_P_btm.n558 C9_P_btm.n557 4.60698
R49617 C9_P_btm.n560 C9_P_btm.n559 4.60698
R49618 C9_P_btm.n561 C9_P_btm.n560 4.60698
R49619 C9_P_btm.n563 C9_P_btm.n562 4.60698
R49620 C9_P_btm.n564 C9_P_btm.n563 4.60698
R49621 C9_P_btm.n566 C9_P_btm.n565 4.60698
R49622 C9_P_btm.n567 C9_P_btm.n566 4.60698
R49623 C9_P_btm.n569 C9_P_btm.n568 4.60698
R49624 C9_P_btm.n570 C9_P_btm.n569 4.60698
R49625 C9_P_btm.n572 C9_P_btm.n571 4.60698
R49626 C9_P_btm.n573 C9_P_btm.n572 4.60698
R49627 C9_P_btm.n575 C9_P_btm.n574 4.60698
R49628 C9_P_btm.n576 C9_P_btm.n575 4.60698
R49629 C9_P_btm.n578 C9_P_btm.n577 4.60698
R49630 C9_P_btm.n579 C9_P_btm.n578 4.60698
R49631 C9_P_btm.n581 C9_P_btm.n580 4.60698
R49632 C9_P_btm.n582 C9_P_btm.n581 4.60698
R49633 C9_P_btm.n584 C9_P_btm.n583 4.60698
R49634 C9_P_btm.n585 C9_P_btm.n584 4.60698
R49635 C9_P_btm.n587 C9_P_btm.n586 4.60698
R49636 C9_P_btm.n588 C9_P_btm.n587 4.60698
R49637 C9_P_btm.n590 C9_P_btm.n589 4.60698
R49638 C9_P_btm.n591 C9_P_btm.n590 4.60698
R49639 C9_P_btm.n593 C9_P_btm.n592 4.60698
R49640 C9_P_btm.n594 C9_P_btm.n593 4.60698
R49641 C9_P_btm.n457 C9_P_btm.n456 4.60698
R49642 C9_P_btm.n456 C9_P_btm.n455 4.60698
R49643 C9_P_btm.n460 C9_P_btm.n459 4.60698
R49644 C9_P_btm.n459 C9_P_btm.n458 4.60698
R49645 C9_P_btm.n463 C9_P_btm.n462 4.60698
R49646 C9_P_btm.n462 C9_P_btm.n461 4.60698
R49647 C9_P_btm.n466 C9_P_btm.n465 4.60698
R49648 C9_P_btm.n465 C9_P_btm.n464 4.60698
R49649 C9_P_btm.n469 C9_P_btm.n468 4.60698
R49650 C9_P_btm.n468 C9_P_btm.n467 4.60698
R49651 C9_P_btm.n472 C9_P_btm.n471 4.60698
R49652 C9_P_btm.n471 C9_P_btm.n470 4.60698
R49653 C9_P_btm.n475 C9_P_btm.n474 4.60698
R49654 C9_P_btm.n474 C9_P_btm.n473 4.60698
R49655 C9_P_btm.n478 C9_P_btm.n477 4.60698
R49656 C9_P_btm.n477 C9_P_btm.n476 4.60698
R49657 C9_P_btm.n481 C9_P_btm.n480 4.60698
R49658 C9_P_btm.n480 C9_P_btm.n479 4.60698
R49659 C9_P_btm.n484 C9_P_btm.n483 4.60698
R49660 C9_P_btm.n483 C9_P_btm.n482 4.60698
R49661 C9_P_btm.n487 C9_P_btm.n486 4.60698
R49662 C9_P_btm.n486 C9_P_btm.n485 4.60698
R49663 C9_P_btm.n490 C9_P_btm.n489 4.60698
R49664 C9_P_btm.n489 C9_P_btm.n488 4.60698
R49665 C9_P_btm.n493 C9_P_btm.n492 4.60698
R49666 C9_P_btm.n492 C9_P_btm.n491 4.60698
R49667 C9_P_btm.n496 C9_P_btm.n495 4.60698
R49668 C9_P_btm.n495 C9_P_btm.n494 4.60698
R49669 C9_P_btm.n596 C9_P_btm.n595 4.60698
R49670 C9_P_btm.n597 C9_P_btm.n596 4.60698
R49671 C9_P_btm.n599 C9_P_btm.n598 4.60698
R49672 C9_P_btm.n600 C9_P_btm.n599 4.60698
R49673 C9_P_btm.n602 C9_P_btm.n601 4.60698
R49674 C9_P_btm.n603 C9_P_btm.n602 4.60698
R49675 C9_P_btm.n605 C9_P_btm.n604 4.60698
R49676 C9_P_btm.n606 C9_P_btm.n605 4.60698
R49677 C9_P_btm.n608 C9_P_btm.n607 4.60698
R49678 C9_P_btm.n609 C9_P_btm.n608 4.60698
R49679 C9_P_btm.n611 C9_P_btm.n610 4.60698
R49680 C9_P_btm.n612 C9_P_btm.n611 4.60698
R49681 C9_P_btm.n614 C9_P_btm.n613 4.60698
R49682 C9_P_btm.n615 C9_P_btm.n614 4.60698
R49683 C9_P_btm.n617 C9_P_btm.n616 4.60698
R49684 C9_P_btm.n618 C9_P_btm.n617 4.60698
R49685 C9_P_btm.n620 C9_P_btm.n619 4.60698
R49686 C9_P_btm.n621 C9_P_btm.n620 4.60698
R49687 C9_P_btm.n623 C9_P_btm.n622 4.60698
R49688 C9_P_btm.n624 C9_P_btm.n623 4.60698
R49689 C9_P_btm.n626 C9_P_btm.n625 4.60698
R49690 C9_P_btm.n627 C9_P_btm.n626 4.60698
R49691 C9_P_btm.n629 C9_P_btm.n628 4.60698
R49692 C9_P_btm.n630 C9_P_btm.n629 4.60698
R49693 C9_P_btm.n1886 C9_P_btm.t23 4.03712
R49694 C9_P_btm.n1884 C9_P_btm.t354 3.98193
R49695 C9_P_btm.n1871 C9_P_btm.t272 3.98193
R49696 C9_P_btm.n1855 C9_P_btm.t101 3.98193
R49697 C9_P_btm.n1804 C9_P_btm.t487 3.98193
R49698 C9_P_btm.n1817 C9_P_btm.t157 3.98193
R49699 C9_P_btm.n1820 C9_P_btm.t119 3.98193
R49700 C9_P_btm.n1802 C9_P_btm.t514 3.98193
R49701 C9_P_btm.n44 C9_P_btm.t231 3.98193
R49702 C9_P_btm.n1768 C9_P_btm.t190 3.98193
R49703 C9_P_btm.n1765 C9_P_btm.t345 3.98193
R49704 C9_P_btm.n67 C9_P_btm.t304 3.98193
R49705 C9_P_btm.n1731 C9_P_btm.t530 3.98193
R49706 C9_P_btm.n1728 C9_P_btm.t432 3.98193
R49707 C9_P_btm.n90 C9_P_btm.t384 3.98193
R49708 C9_P_btm.n1694 C9_P_btm.t259 3.98193
R49709 C9_P_btm.n1691 C9_P_btm.t102 3.98193
R49710 C9_P_btm.n113 C9_P_btm.t473 3.98193
R49711 C9_P_btm.n1657 C9_P_btm.t140 3.98193
R49712 C9_P_btm.n1346 C9_P_btm.t220 3.98193
R49713 C9_P_btm.n1511 C9_P_btm.t115 3.98193
R49714 C9_P_btm.n1508 C9_P_btm.t104 3.98193
R49715 C9_P_btm.n1317 C9_P_btm.t191 3.98193
R49716 C9_P_btm.n1262 C9_P_btm.t47 3.98193
R49717 C9_P_btm.n930 C9_P_btm.t86 3.98193
R49718 C9_P_btm.n1232 C9_P_btm.t420 3.98193
R49719 C9_P_btm.n1229 C9_P_btm.t472 3.98193
R49720 C9_P_btm.n941 C9_P_btm.t53 3.98193
R49721 C9_P_btm.n1195 C9_P_btm.t335 3.98193
R49722 C9_P_btm.n1192 C9_P_btm.t383 3.98193
R49723 C9_P_btm.n964 C9_P_btm.t210 3.98193
R49724 C9_P_btm.n1158 C9_P_btm.t528 3.98193
R49725 C9_P_btm.n1155 C9_P_btm.t303 3.98193
R49726 C9_P_btm.n987 C9_P_btm.t144 3.98193
R49727 C9_P_btm.n1121 C9_P_btm.t519 3.98193
R49728 C9_P_btm.n1118 C9_P_btm.t288 3.98193
R49729 C9_P_btm.n1010 C9_P_btm.t399 3.98193
R49730 C9_P_btm.n1084 C9_P_btm.t114 3.98193
R49731 C9_P_btm.n1081 C9_P_btm.t436 3.98193
R49732 C9_P_btm.n1032 C9_P_btm.t486 3.98193
R49733 C9_P_btm.n1047 C9_P_btm.t306 3.98193
R49734 C9_P_btm.n1060 C9_P_btm.t251 3.98193
R49735 C9_P_btm.n1063 C9_P_btm.t421 3.98193
R49736 C9_P_btm.n1068 C9_P_btm.t372 3.98193
R49737 C9_P_btm.n1097 C9_P_btm.t51 3.98193
R49738 C9_P_btm.n1100 C9_P_btm.t508 3.98193
R49739 C9_P_btm.n1105 C9_P_btm.t455 3.98193
R49740 C9_P_btm.n1134 C9_P_btm.t129 3.98193
R49741 C9_P_btm.n1137 C9_P_btm.t82 3.98193
R49742 C9_P_btm.n1142 C9_P_btm.t502 3.98193
R49743 C9_P_btm.n1171 C9_P_btm.t200 3.98193
R49744 C9_P_btm.n1174 C9_P_btm.t168 3.98193
R49745 C9_P_btm.n1179 C9_P_btm.t322 3.98193
R49746 C9_P_btm.n1208 C9_P_btm.t279 3.98193
R49747 C9_P_btm.n1211 C9_P_btm.t451 3.98193
R49748 C9_P_btm.n1216 C9_P_btm.t409 3.98193
R49749 C9_P_btm.n1245 C9_P_btm.t363 3.98193
R49750 C9_P_btm.n1248 C9_P_btm.t301 3.98193
R49751 C9_P_btm.n883 C9_P_btm.t31 3.98193
R49752 C9_P_btm.n255 C9_P_btm.t443 3.98193
R49753 C9_P_btm.n633 C9_P_btm.t494 3.98193
R49754 C9_P_btm.n454 C9_P_btm.t185 3.98193
R49755 C9_P_btm.n497 C9_P_btm.t26 3.98193
R49756 C9_P_btm.n631 C9_P_btm.t321 3.98193
R49757 C9_P_btm.n216 C9_P_btm.t527 3.98193
R49758 C9_P_btm.n754 C9_P_btm.t313 3.98193
R49759 C9_P_btm.n757 C9_P_btm.t138 3.98193
R49760 C9_P_btm.n762 C9_P_btm.t151 3.98193
R49761 C9_P_btm.n1632 C9_P_btm.t320 3.98193
R49762 C9_P_btm.n1635 C9_P_btm.t194 3.98193
R49763 C9_P_btm.n1640 C9_P_btm.t280 3.98193
R49764 C9_P_btm.n1670 C9_P_btm.t474 3.98193
R49765 C9_P_btm.n1673 C9_P_btm.t201 3.98193
R49766 C9_P_btm.n1678 C9_P_btm.t385 3.98193
R49767 C9_P_btm.n1707 C9_P_btm.t71 3.98193
R49768 C9_P_btm.n1710 C9_P_btm.t302 3.98193
R49769 C9_P_btm.n1715 C9_P_btm.t497 3.98193
R49770 C9_P_btm.n1744 C9_P_btm.t225 3.98193
R49771 C9_P_btm.n1747 C9_P_btm.t410 3.98193
R49772 C9_P_btm.n1752 C9_P_btm.t90 3.98193
R49773 C9_P_btm.n1781 C9_P_btm.t323 3.98193
R49774 C9_P_btm.n1784 C9_P_btm.t117 3.98193
R49775 C9_P_btm.n1789 C9_P_btm.t512 3.98193
R49776 C9_P_btm.n1833 C9_P_btm.t433 3.98193
R49777 C9_P_btm.n1836 C9_P_btm.t351 3.98193
R49778 C9_P_btm.n1841 C9_P_btm.t344 3.98193
R49779 C9_P_btm.n1868 C9_P_btm.t27 3.98193
R49780 C9_P_btm.n11 C9_P_btm.n10 3.91717
R49781 C9_P_btm.n5 C9_P_btm.t5 3.57113
R49782 C9_P_btm.n5 C9_P_btm.t8 3.57113
R49783 C9_P_btm.n3 C9_P_btm.t9 3.57113
R49784 C9_P_btm.n3 C9_P_btm.t10 3.57113
R49785 C9_P_btm.n1 C9_P_btm.t11 3.57113
R49786 C9_P_btm.n1 C9_P_btm.t12 3.57113
R49787 C9_P_btm.n0 C9_P_btm.t7 3.57113
R49788 C9_P_btm.n0 C9_P_btm.t6 3.57113
R49789 C9_P_btm.n7 C9_P_btm.t2 2.4755
R49790 C9_P_btm.n7 C9_P_btm.t3 2.4755
R49791 C9_P_btm.n13 C9_P_btm.t540 2.4755
R49792 C9_P_btm.n13 C9_P_btm.t539 2.4755
R49793 C9_P_btm.n12 C9_P_btm.t538 2.4755
R49794 C9_P_btm.n12 C9_P_btm.t537 2.4755
R49795 C9_P_btm.n8 C9_P_btm.t1 2.4755
R49796 C9_P_btm.n8 C9_P_btm.t0 2.4755
R49797 C9_P_btm.n1882 C9_P_btm.t215 1.67819
R49798 C9_P_btm.n1879 C9_P_btm.t398 1.67819
R49799 C9_P_btm.n1876 C9_P_btm.t260 1.67819
R49800 C9_P_btm.n1873 C9_P_btm.t404 1.67819
R49801 C9_P_btm.n1866 C9_P_btm.t173 1.67819
R49802 C9_P_btm.n1863 C9_P_btm.t274 1.67819
R49803 C9_P_btm.n1860 C9_P_btm.t278 1.67819
R49804 C9_P_btm.n1857 C9_P_btm.t388 1.67819
R49805 C9_P_btm.n1851 C9_P_btm.t336 1.67819
R49806 C9_P_btm.n1849 C9_P_btm.t256 1.67819
R49807 C9_P_btm.n1846 C9_P_btm.t95 1.67819
R49808 C9_P_btm.n1843 C9_P_btm.t490 1.67819
R49809 C9_P_btm.n1837 C9_P_btm.t499 1.67819
R49810 C9_P_btm.n1809 C9_P_btm.t352 1.67819
R49811 C9_P_btm.n1812 C9_P_btm.t408 1.67819
R49812 C9_P_btm.n1815 C9_P_btm.t516 1.67819
R49813 C9_P_btm.n1822 C9_P_btm.t479 1.67819
R49814 C9_P_btm.n1825 C9_P_btm.t362 1.67819
R49815 C9_P_btm.n1828 C9_P_btm.t177 1.67819
R49816 C9_P_btm.n1831 C9_P_btm.t62 1.67819
R49817 C9_P_btm.n1791 C9_P_btm.t379 1.67819
R49818 C9_P_btm.n1794 C9_P_btm.t511 1.67819
R49819 C9_P_btm.n1797 C9_P_btm.t315 1.67819
R49820 C9_P_btm.n1800 C9_P_btm.t424 1.67819
R49821 C9_P_btm.n54 C9_P_btm.t96 1.67819
R49822 C9_P_btm.n52 C9_P_btm.t492 1.67819
R49823 C9_P_btm.n49 C9_P_btm.t252 1.67819
R49824 C9_P_btm.n1785 C9_P_btm.t153 1.67819
R49825 C9_P_btm.n1779 C9_P_btm.t468 1.67819
R49826 C9_P_btm.n1776 C9_P_btm.t73 1.67819
R49827 C9_P_btm.n1773 C9_P_btm.t442 1.67819
R49828 C9_P_btm.n1770 C9_P_btm.t108 1.67819
R49829 C9_P_btm.n1763 C9_P_btm.t211 1.67819
R49830 C9_P_btm.n1760 C9_P_btm.t254 1.67819
R49831 C9_P_btm.n1757 C9_P_btm.t329 1.67819
R49832 C9_P_btm.n1754 C9_P_btm.t218 1.67819
R49833 C9_P_btm.n1748 C9_P_btm.t44 1.67819
R49834 C9_P_btm.n72 C9_P_btm.t163 1.67819
R49835 C9_P_btm.n75 C9_P_btm.t63 1.67819
R49836 C9_P_btm.n77 C9_P_btm.t179 1.67819
R49837 C9_P_btm.n1733 C9_P_btm.t132 1.67819
R49838 C9_P_btm.n1736 C9_P_btm.t42 1.67819
R49839 C9_P_btm.n1739 C9_P_btm.t475 1.67819
R49840 C9_P_btm.n1742 C9_P_btm.t358 1.67819
R49841 C9_P_btm.n1717 C9_P_btm.t124 1.67819
R49842 C9_P_btm.n1720 C9_P_btm.t233 1.67819
R49843 C9_P_btm.n1723 C9_P_btm.t196 1.67819
R49844 C9_P_btm.n1726 C9_P_btm.t293 1.67819
R49845 C9_P_btm.n100 C9_P_btm.t520 1.67819
R49846 C9_P_btm.n98 C9_P_btm.t154 1.67819
R49847 C9_P_btm.n95 C9_P_btm.t105 1.67819
R49848 C9_P_btm.n1711 C9_P_btm.t440 1.67819
R49849 C9_P_btm.n1705 C9_P_btm.t199 1.67819
R49850 C9_P_btm.n1702 C9_P_btm.t307 1.67819
R49851 C9_P_btm.n1699 C9_P_btm.t310 1.67819
R49852 C9_P_btm.n1696 C9_P_btm.t422 1.67819
R49853 C9_P_btm.n1689 C9_P_btm.t373 1.67819
R49854 C9_P_btm.n1686 C9_P_btm.t264 1.67819
R49855 C9_P_btm.n1683 C9_P_btm.t130 1.67819
R49856 C9_P_btm.n1680 C9_P_btm.t34 1.67819
R49857 C9_P_btm.n1674 C9_P_btm.t332 1.67819
R49858 C9_P_btm.n118 C9_P_btm.t447 1.67819
R49859 C9_P_btm.n121 C9_P_btm.t217 1.67819
R49860 C9_P_btm.n123 C9_P_btm.t327 1.67819
R49861 C9_P_btm.n1659 C9_P_btm.t509 1.67819
R49862 C9_P_btm.n1662 C9_P_btm.t390 1.67819
R49863 C9_P_btm.n1665 C9_P_btm.t205 1.67819
R49864 C9_P_btm.n1668 C9_P_btm.t111 1.67819
R49865 C9_P_btm.n1642 C9_P_btm.t417 1.67819
R49866 C9_P_btm.n1645 C9_P_btm.t109 1.67819
R49867 C9_P_btm.n1648 C9_P_btm.t341 1.67819
R49868 C9_P_btm.n1651 C9_P_btm.t458 1.67819
R49869 C9_P_btm.n1653 C9_P_btm.t88 1.67819
R49870 C9_P_btm.n1384 C9_P_btm.t431 1.67819
R49871 C9_P_btm.n1381 C9_P_btm.t35 1.67819
R49872 C9_P_btm.n1378 C9_P_btm.t176 1.67819
R49873 C9_P_btm.n1375 C9_P_btm.t70 1.67819
R49874 C9_P_btm.n1372 C9_P_btm.t125 1.67819
R49875 C9_P_btm.n1369 C9_P_btm.t495 1.67819
R49876 C9_P_btm.n1366 C9_P_btm.t99 1.67819
R49877 C9_P_btm.n1363 C9_P_btm.t202 1.67819
R49878 C9_P_btm.n1360 C9_P_btm.t56 1.67819
R49879 C9_P_btm.n1357 C9_P_btm.t184 1.67819
R49880 C9_P_btm.n1354 C9_P_btm.t283 1.67819
R49881 C9_P_btm.n1351 C9_P_btm.t134 1.67819
R49882 C9_P_btm.n1348 C9_P_btm.t532 1.67819
R49883 C9_P_btm.n1443 C9_P_btm.t167 1.67819
R49884 C9_P_btm.n1440 C9_P_btm.t311 1.67819
R49885 C9_P_btm.n1437 C9_P_btm.t187 1.67819
R49886 C9_P_btm.n1434 C9_P_btm.t333 1.67819
R49887 C9_P_btm.n1431 C9_P_btm.t240 1.67819
R49888 C9_P_btm.n1428 C9_P_btm.t110 1.67819
R49889 C9_P_btm.n1425 C9_P_btm.t522 1.67819
R49890 C9_P_btm.n1422 C9_P_btm.t161 1.67819
R49891 C9_P_btm.n1419 C9_P_btm.t43 1.67819
R49892 C9_P_btm.n1416 C9_P_btm.t180 1.67819
R49893 C9_P_btm.n1413 C9_P_btm.t66 1.67819
R49894 C9_P_btm.n1410 C9_P_btm.t222 1.67819
R49895 C9_P_btm.n1407 C9_P_btm.t92 1.67819
R49896 C9_P_btm.n1404 C9_P_btm.t489 1.67819
R49897 C9_P_btm.n1401 C9_P_btm.t149 1.67819
R49898 C9_P_btm.n1398 C9_P_btm.t38 1.67819
R49899 C9_P_btm.n1395 C9_P_btm.t400 1.67819
R49900 C9_P_btm.n1392 C9_P_btm.t247 1.67819
R49901 C9_P_btm.n1636 C9_P_btm.t146 1.67819
R49902 C9_P_btm.n1630 C9_P_btm.t462 1.67819
R49903 C9_P_btm.n1627 C9_P_btm.t68 1.67819
R49904 C9_P_btm.n1624 C9_P_btm.t355 1.67819
R49905 C9_P_btm.n1621 C9_P_btm.t471 1.67819
R49906 C9_P_btm.n1618 C9_P_btm.t106 1.67819
R49907 C9_P_btm.n1615 C9_P_btm.t439 1.67819
R49908 C9_P_btm.n1612 C9_P_btm.t100 1.67819
R49909 C9_P_btm.n1609 C9_P_btm.t186 1.67819
R49910 C9_P_btm.n1606 C9_P_btm.t94 1.67819
R49911 C9_P_btm.n1603 C9_P_btm.t136 1.67819
R49912 C9_P_btm.n1600 C9_P_btm.t507 1.67819
R49913 C9_P_btm.n1597 C9_P_btm.t232 1.67819
R49914 C9_P_btm.n1594 C9_P_btm.t208 1.67819
R49915 C9_P_btm.n1591 C9_P_btm.t236 1.67819
R49916 C9_P_btm.n1588 C9_P_btm.t193 1.67819
R49917 C9_P_btm.n1585 C9_P_btm.t289 1.67819
R49918 C9_P_btm.n1582 C9_P_btm.t143 1.67819
R49919 C9_P_btm.n1579 C9_P_btm.t266 1.67819
R49920 C9_P_btm.n1576 C9_P_btm.t268 1.67819
R49921 C9_P_btm.n1573 C9_P_btm.t213 1.67819
R49922 C9_P_btm.n1570 C9_P_btm.t347 1.67819
R49923 C9_P_btm.n1567 C9_P_btm.t533 1.67819
R49924 C9_P_btm.n1564 C9_P_btm.t295 1.67819
R49925 C9_P_btm.n1561 C9_P_btm.t411 1.67819
R49926 C9_P_btm.n1558 C9_P_btm.t277 1.67819
R49927 C9_P_btm.n1555 C9_P_btm.t381 1.67819
R49928 C9_P_btm.n1552 C9_P_btm.t226 1.67819
R49929 C9_P_btm.n1549 C9_P_btm.t359 1.67819
R49930 C9_P_btm.n1546 C9_P_btm.t476 1.67819
R49931 C9_P_btm.n1543 C9_P_btm.t326 1.67819
R49932 C9_P_btm.n1540 C9_P_btm.t470 1.67819
R49933 C9_P_btm.n1537 C9_P_btm.t76 1.67819
R49934 C9_P_btm.n1534 C9_P_btm.t416 1.67819
R49935 C9_P_btm.n1531 C9_P_btm.t52 1.67819
R49936 C9_P_btm.n1528 C9_P_btm.t165 1.67819
R49937 C9_P_btm.n1525 C9_P_btm.t506 1.67819
R49938 C9_P_btm.n1522 C9_P_btm.t227 1.67819
R49939 C9_P_btm.n1519 C9_P_btm.t480 1.67819
R49940 C9_P_btm.n1516 C9_P_btm.t81 1.67819
R49941 C9_P_btm.n1513 C9_P_btm.t524 1.67819
R49942 C9_P_btm.n1506 C9_P_btm.t238 1.67819
R49943 C9_P_btm.n1503 C9_P_btm.t128 1.67819
R49944 C9_P_btm.n1500 C9_P_btm.t25 1.67819
R49945 C9_P_btm.n1497 C9_P_btm.t160 1.67819
R49946 C9_P_btm.n1494 C9_P_btm.t41 1.67819
R49947 C9_P_btm.n1491 C9_P_btm.t198 1.67819
R49948 C9_P_btm.n1488 C9_P_btm.t65 1.67819
R49949 C9_P_btm.n1485 C9_P_btm.t461 1.67819
R49950 C9_P_btm.n1482 C9_P_btm.t121 1.67819
R49951 C9_P_btm.n1479 C9_P_btm.t517 1.67819
R49952 C9_P_btm.n1476 C9_P_btm.t370 1.67819
R49953 C9_P_btm.n1473 C9_P_btm.t324 1.67819
R49954 C9_P_btm.n1470 C9_P_btm.t405 1.67819
R49955 C9_P_btm.n1467 C9_P_btm.t273 1.67819
R49956 C9_P_btm.n1464 C9_P_btm.t429 1.67819
R49957 C9_P_btm.n1461 C9_P_btm.t318 1.67819
R49958 C9_P_btm.n1458 C9_P_btm.t456 1.67819
R49959 C9_P_btm.n1455 C9_P_btm.t339 1.67819
R49960 C9_P_btm.n1452 C9_P_btm.t267 1.67819
R49961 C9_P_btm.n1315 C9_P_btm.t286 1.67819
R49962 C9_P_btm.n1312 C9_P_btm.t401 1.67819
R49963 C9_P_btm.n1309 C9_P_btm.t265 1.67819
R49964 C9_P_btm.n1306 C9_P_btm.t374 1.67819
R49965 C9_P_btm.n1303 C9_P_btm.t212 1.67819
R49966 C9_P_btm.n1300 C9_P_btm.t346 1.67819
R49967 C9_P_btm.n1297 C9_P_btm.t464 1.67819
R49968 C9_P_btm.n1294 C9_P_btm.t317 1.67819
R49969 C9_P_btm.n1291 C9_P_btm.t453 1.67819
R49970 C9_P_btm.n1288 C9_P_btm.t60 1.67819
R49971 C9_P_btm.n1285 C9_P_btm.t403 1.67819
R49972 C9_P_btm.n1282 C9_P_btm.t245 1.67819
R49973 C9_P_btm.n1279 C9_P_btm.t155 1.67819
R49974 C9_P_btm.n1276 C9_P_btm.t493 1.67819
R49975 C9_P_btm.n1273 C9_P_btm.t98 1.67819
R49976 C9_P_btm.n1270 C9_P_btm.t465 1.67819
R49977 C9_P_btm.n1267 C9_P_btm.t72 1.67819
R49978 C9_P_btm.n1264 C9_P_btm.t182 1.67819
R49979 C9_P_btm.n1258 C9_P_btm.t216 1.67819
R49980 C9_P_btm.n1256 C9_P_btm.t500 1.67819
R49981 C9_P_btm.n1253 C9_P_btm.t521 1.67819
R49982 C9_P_btm.n1250 C9_P_btm.t145 1.67819
R49983 C9_P_btm.n1243 C9_P_btm.t481 1.67819
R49984 C9_P_btm.n1240 C9_P_btm.t331 1.67819
R49985 C9_P_btm.n1237 C9_P_btm.t446 1.67819
R49986 C9_P_btm.n1234 C9_P_btm.t228 1.67819
R49987 C9_P_btm.n1227 C9_P_btm.t107 1.67819
R49988 C9_P_btm.n1224 C9_P_btm.t510 1.67819
R49989 C9_P_btm.n1221 C9_P_btm.t378 1.67819
R49990 C9_P_btm.n1218 C9_P_btm.t30 1.67819
R49991 C9_P_btm.n1212 C9_P_btm.t59 1.67819
R49992 C9_P_btm.n946 C9_P_btm.t426 1.67819
R49993 C9_P_btm.n949 C9_P_btm.t28 1.67819
R49994 C9_P_btm.n951 C9_P_btm.t152 1.67819
R49995 C9_P_btm.n1197 C9_P_btm.t482 1.67819
R49996 C9_P_btm.n1200 C9_P_btm.t365 1.67819
R49997 C9_P_btm.n1203 C9_P_btm.t526 1.67819
R49998 C9_P_btm.n1206 C9_P_btm.t389 1.67819
R49999 C9_P_btm.n1181 C9_P_btm.t437 1.67819
R50000 C9_P_btm.n1184 C9_P_btm.t297 1.67819
R50001 C9_P_btm.n1187 C9_P_btm.t413 1.67819
R50002 C9_P_btm.n1190 C9_P_btm.t37 1.67819
R50003 C9_P_btm.n974 C9_P_btm.t342 1.67819
R50004 C9_P_btm.n972 C9_P_btm.t298 1.67819
R50005 C9_P_btm.n969 C9_P_btm.t139 1.67819
R50006 C9_P_btm.n1175 C9_P_btm.t263 1.67819
R50007 C9_P_btm.n1169 C9_P_btm.t309 1.67819
R50008 C9_P_btm.n1166 C9_P_btm.t183 1.67819
R50009 C9_P_btm.n1163 C9_P_btm.t282 1.67819
R50010 C9_P_btm.n1160 C9_P_btm.t392 1.67819
R50011 C9_P_btm.n1153 C9_P_btm.t441 1.67819
R50012 C9_P_btm.n1150 C9_P_btm.t328 1.67819
R50013 C9_P_btm.n1147 C9_P_btm.t219 1.67819
R50014 C9_P_btm.n1144 C9_P_btm.t356 1.67819
R50015 C9_P_btm.n1138 C9_P_btm.t195 1.67819
R50016 C9_P_btm.n992 C9_P_btm.t243 1.67819
R50017 C9_P_btm.n995 C9_P_btm.t172 1.67819
R50018 C9_P_btm.n997 C9_P_btm.t270 1.67819
R50019 C9_P_btm.n1123 C9_P_btm.t314 1.67819
R50020 C9_P_btm.n1126 C9_P_btm.t206 1.67819
R50021 C9_P_btm.n1129 C9_P_btm.t113 1.67819
R50022 C9_P_btm.n1132 C9_P_btm.t246 1.67819
R50023 C9_P_btm.n1107 C9_P_btm.t61 1.67819
R50024 C9_P_btm.n1110 C9_P_btm.t428 1.67819
R50025 C9_P_btm.n1113 C9_P_btm.t32 1.67819
R50026 C9_P_btm.n1116 C9_P_btm.t156 1.67819
R50027 C9_P_btm.n1020 C9_P_btm.t197 1.67819
R50028 C9_P_btm.n1018 C9_P_btm.t83 1.67819
R50029 C9_P_btm.n1015 C9_P_btm.t483 1.67819
R50030 C9_P_btm.n1101 C9_P_btm.t239 1.67819
R50031 C9_P_btm.n1095 C9_P_btm.t164 1.67819
R50032 C9_P_btm.n1092 C9_P_btm.t45 1.67819
R50033 C9_P_btm.n1089 C9_P_btm.t133 1.67819
R50034 C9_P_btm.n1086 C9_P_btm.t253 1.67819
R50035 C9_P_btm.n1079 C9_P_btm.t69 1.67819
R50036 C9_P_btm.n1076 C9_P_btm.t463 1.67819
R50037 C9_P_btm.n1073 C9_P_btm.t343 1.67819
R50038 C9_P_btm.n1070 C9_P_btm.t491 1.67819
R50039 C9_P_btm.n1064 C9_P_btm.t244 1.67819
R50040 C9_P_btm.n1037 C9_P_btm.t393 1.67819
R50041 C9_P_btm.n1040 C9_P_btm.t39 1.67819
R50042 C9_P_btm.n1042 C9_P_btm.t299 1.67819
R50043 C9_P_btm.n1049 C9_P_btm.t444 1.67819
R50044 C9_P_btm.n1052 C9_P_btm.t330 1.67819
R50045 C9_P_btm.n1055 C9_P_btm.t230 1.67819
R50046 C9_P_btm.n1058 C9_P_btm.t361 1.67819
R50047 C9_P_btm.n1449 C9_P_btm.t394 1.67819
R50048 C9_P_btm.n1446 C9_P_btm.t534 1.67819
R50049 C9_P_btm.n881 C9_P_btm.t147 1.67819
R50050 C9_P_btm.n878 C9_P_btm.t29 1.67819
R50051 C9_P_btm.n875 C9_P_btm.t425 1.67819
R50052 C9_P_btm.n872 C9_P_btm.t57 1.67819
R50053 C9_P_btm.n869 C9_P_btm.t449 1.67819
R50054 C9_P_btm.n866 C9_P_btm.t242 1.67819
R50055 C9_P_btm.n863 C9_P_btm.t484 1.67819
R50056 C9_P_btm.n860 C9_P_btm.t366 1.67819
R50057 C9_P_btm.n857 C9_P_btm.t116 1.67819
R50058 C9_P_btm.n854 C9_P_btm.t418 1.67819
R50059 C9_P_btm.n851 C9_P_btm.t281 1.67819
R50060 C9_P_btm.n848 C9_P_btm.t423 1.67819
R50061 C9_P_btm.n845 C9_P_btm.t312 1.67819
R50062 C9_P_btm.n842 C9_P_btm.t188 1.67819
R50063 C9_P_btm.n839 C9_P_btm.t334 1.67819
R50064 C9_P_btm.n836 C9_P_btm.t241 1.67819
R50065 C9_P_btm.n833 C9_P_btm.t364 1.67819
R50066 C9_P_btm.n830 C9_P_btm.t255 1.67819
R50067 C9_P_btm.n827 C9_P_btm.t162 1.67819
R50068 C9_P_btm.n824 C9_P_btm.t305 1.67819
R50069 C9_P_btm.n821 C9_P_btm.t181 1.67819
R50070 C9_P_btm.n818 C9_P_btm.t67 1.67819
R50071 C9_P_btm.n815 C9_P_btm.t223 1.67819
R50072 C9_P_btm.n812 C9_P_btm.t91 1.67819
R50073 C9_P_btm.n809 C9_P_btm.t250 1.67819
R50074 C9_P_btm.n806 C9_P_btm.t150 1.67819
R50075 C9_P_btm.n803 C9_P_btm.t46 1.67819
R50076 C9_P_btm.n800 C9_P_btm.t175 1.67819
R50077 C9_P_btm.n797 C9_P_btm.t58 1.67819
R50078 C9_P_btm.n794 C9_P_btm.t450 1.67819
R50079 C9_P_btm.n791 C9_P_btm.t85 1.67819
R50080 C9_P_btm.n788 C9_P_btm.t485 1.67819
R50081 C9_P_btm.n785 C9_P_btm.t142 1.67819
R50082 C9_P_btm.n782 C9_P_btm.t518 1.67819
R50083 C9_P_btm.n779 C9_P_btm.t391 1.67819
R50084 C9_P_btm.n776 C9_P_btm.t221 1.67819
R50085 C9_P_btm.n773 C9_P_btm.t419 1.67819
R50086 C9_P_btm.n770 C9_P_btm.t308 1.67819
R50087 C9_P_btm.n767 C9_P_btm.t380 1.67819
R50088 C9_P_btm.n764 C9_P_btm.t276 1.67819
R50089 C9_P_btm.n758 C9_P_btm.t536 1.67819
R50090 C9_P_btm.n296 C9_P_btm.t371 1.67819
R50091 C9_P_btm.n299 C9_P_btm.t452 1.67819
R50092 C9_P_btm.n302 C9_P_btm.t353 1.67819
R50093 C9_P_btm.n305 C9_P_btm.t496 1.67819
R50094 C9_P_btm.n308 C9_P_btm.t158 1.67819
R50095 C9_P_btm.n311 C9_P_btm.t438 1.67819
R50096 C9_P_btm.n314 C9_P_btm.t74 1.67819
R50097 C9_P_btm.n317 C9_P_btm.t414 1.67819
R50098 C9_P_btm.n320 C9_P_btm.t49 1.67819
R50099 C9_P_btm.n323 C9_P_btm.t386 1.67819
R50100 C9_P_btm.n326 C9_P_btm.t504 1.67819
R50101 C9_P_btm.n329 C9_P_btm.t224 1.67819
R50102 C9_P_btm.n332 C9_P_btm.t445 1.67819
R50103 C9_P_btm.n335 C9_P_btm.t79 1.67819
R50104 C9_P_btm.n338 C9_P_btm.t192 1.67819
R50105 C9_P_btm.n341 C9_P_btm.t229 1.67819
R50106 C9_P_btm.n344 C9_P_btm.t169 1.67819
R50107 C9_P_btm.n347 C9_P_btm.t55 1.67819
R50108 C9_P_btm.n350 C9_P_btm.t258 1.67819
R50109 C9_P_btm.n353 C9_P_btm.t350 1.67819
R50110 C9_P_btm.n356 C9_P_btm.t84 1.67819
R50111 C9_P_btm.n359 C9_P_btm.t531 1.67819
R50112 C9_P_btm.n362 C9_P_btm.t294 1.67819
R50113 C9_P_btm.n365 C9_P_btm.t174 1.67819
R50114 C9_P_btm.n368 C9_P_btm.t275 1.67819
R50115 C9_P_btm.n371 C9_P_btm.t122 1.67819
R50116 C9_P_btm.n374 C9_P_btm.t249 1.67819
R50117 C9_P_btm.n377 C9_P_btm.t357 1.67819
R50118 C9_P_btm.n380 C9_P_btm.t214 1.67819
R50119 C9_P_btm.n383 C9_P_btm.t348 1.67819
R50120 C9_P_btm.n386 C9_P_btm.t466 1.67819
R50121 C9_P_btm.n389 C9_P_btm.t296 1.67819
R50122 C9_P_btm.n392 C9_P_btm.t412 1.67819
R50123 C9_P_btm.n395 C9_P_btm.t48 1.67819
R50124 C9_P_btm.n398 C9_P_btm.t382 1.67819
R50125 C9_P_btm.n401 C9_P_btm.t503 1.67819
R50126 C9_P_btm.n404 C9_P_btm.t360 1.67819
R50127 C9_P_btm.n407 C9_P_btm.t477 1.67819
R50128 C9_P_btm.n409 C9_P_btm.t78 1.67819
R50129 C9_P_btm.n635 C9_P_btm.t123 1.67819
R50130 C9_P_btm.n638 C9_P_btm.t529 1.67819
R50131 C9_P_btm.n641 C9_P_btm.t406 1.67819
R50132 C9_P_btm.n644 C9_P_btm.t33 1.67819
R50133 C9_P_btm.n647 C9_P_btm.t430 1.67819
R50134 C9_P_btm.n650 C9_P_btm.t87 1.67819
R50135 C9_P_btm.n653 C9_P_btm.t457 1.67819
R50136 C9_P_btm.n656 C9_P_btm.t340 1.67819
R50137 C9_P_btm.n659 C9_P_btm.t54 1.67819
R50138 C9_P_btm.n662 C9_P_btm.t395 1.67819
R50139 C9_P_btm.n665 C9_P_btm.t535 1.67819
R50140 C9_P_btm.n668 C9_P_btm.t402 1.67819
R50141 C9_P_btm.n671 C9_P_btm.t287 1.67819
R50142 C9_P_btm.n674 C9_P_btm.t171 1.67819
R50143 C9_P_btm.n677 C9_P_btm.t316 1.67819
R50144 C9_P_btm.n680 C9_P_btm.t207 1.67819
R50145 C9_P_btm.n683 C9_P_btm.t337 1.67819
R50146 C9_P_btm.n686 C9_P_btm.t257 1.67819
R50147 C9_P_btm.n689 C9_P_btm.t135 1.67819
R50148 C9_P_btm.n692 C9_P_btm.t284 1.67819
R50149 C9_P_btm.n695 C9_P_btm.t166 1.67819
R50150 C9_P_btm.n698 C9_P_btm.t93 1.67819
R50151 C9_P_btm.n701 C9_P_btm.t203 1.67819
R50152 C9_P_btm.n704 C9_P_btm.t77 1.67819
R50153 C9_P_btm.n707 C9_P_btm.t234 1.67819
R50154 C9_P_btm.n710 C9_P_btm.t126 1.67819
R50155 C9_P_btm.n713 C9_P_btm.t501 1.67819
R50156 C9_P_btm.n716 C9_P_btm.t159 1.67819
R50157 C9_P_btm.n719 C9_P_btm.t36 1.67819
R50158 C9_P_btm.n722 C9_P_btm.t434 1.67819
R50159 C9_P_btm.n725 C9_P_btm.t64 1.67819
R50160 C9_P_btm.n728 C9_P_btm.t459 1.67819
R50161 C9_P_btm.n731 C9_P_btm.t513 1.67819
R50162 C9_P_btm.n734 C9_P_btm.t488 1.67819
R50163 C9_P_btm.n737 C9_P_btm.t368 1.67819
R50164 C9_P_btm.n740 C9_P_btm.t515 1.67819
R50165 C9_P_btm.n743 C9_P_btm.t396 1.67819
R50166 C9_P_btm.n746 C9_P_btm.t285 1.67819
R50167 C9_P_btm.n749 C9_P_btm.t300 1.67819
R50168 C9_P_btm.n752 C9_P_btm.t448 1.67819
R50169 C9_P_btm.n512 C9_P_btm.t148 1.67819
R50170 C9_P_btm.n515 C9_P_btm.t248 1.67819
R50171 C9_P_btm.n518 C9_P_btm.t137 1.67819
R50172 C9_P_btm.n521 C9_P_btm.t292 1.67819
R50173 C9_P_btm.n524 C9_P_btm.t367 1.67819
R50174 C9_P_btm.n527 C9_P_btm.t209 1.67819
R50175 C9_P_btm.n530 C9_P_btm.t319 1.67819
R50176 C9_P_btm.n533 C9_P_btm.t454 1.67819
R50177 C9_P_btm.n536 C9_P_btm.t291 1.67819
R50178 C9_P_btm.n539 C9_P_btm.t407 1.67819
R50179 C9_P_btm.n542 C9_P_btm.t271 1.67819
R50180 C9_P_btm.n545 C9_P_btm.t376 1.67819
R50181 C9_P_btm.n548 C9_P_btm.t498 1.67819
R50182 C9_P_btm.n551 C9_P_btm.t325 1.67819
R50183 C9_P_btm.n554 C9_P_btm.t469 1.67819
R50184 C9_P_btm.n557 C9_P_btm.t75 1.67819
R50185 C9_P_btm.n560 C9_P_btm.t415 1.67819
R50186 C9_P_btm.n563 C9_P_btm.t50 1.67819
R50187 C9_P_btm.n566 C9_P_btm.t387 1.67819
R50188 C9_P_btm.n569 C9_P_btm.t505 1.67819
R50189 C9_P_btm.n572 C9_P_btm.t131 1.67819
R50190 C9_P_btm.n575 C9_P_btm.t478 1.67819
R50191 C9_P_btm.n578 C9_P_btm.t80 1.67819
R50192 C9_P_btm.n581 C9_P_btm.t523 1.67819
R50193 C9_P_btm.n584 C9_P_btm.t112 1.67819
R50194 C9_P_btm.n587 C9_P_btm.t170 1.67819
R50195 C9_P_btm.n590 C9_P_btm.t189 1.67819
R50196 C9_P_btm.n593 C9_P_btm.t141 1.67819
R50197 C9_P_btm.n456 C9_P_btm.t97 1.67819
R50198 C9_P_btm.n459 C9_P_btm.t204 1.67819
R50199 C9_P_btm.n462 C9_P_btm.t103 1.67819
R50200 C9_P_btm.n465 C9_P_btm.t237 1.67819
R50201 C9_P_btm.n468 C9_P_btm.t127 1.67819
R50202 C9_P_btm.n471 C9_P_btm.t262 1.67819
R50203 C9_P_btm.n474 C9_P_btm.t178 1.67819
R50204 C9_P_btm.n477 C9_P_btm.t40 1.67819
R50205 C9_P_btm.n480 C9_P_btm.t435 1.67819
R50206 C9_P_btm.n483 C9_P_btm.t89 1.67819
R50207 C9_P_btm.n486 C9_P_btm.t460 1.67819
R50208 C9_P_btm.n489 C9_P_btm.t120 1.67819
R50209 C9_P_btm.n492 C9_P_btm.t118 1.67819
R50210 C9_P_btm.n495 C9_P_btm.t369 1.67819
R50211 C9_P_btm.n596 C9_P_btm.t377 1.67819
R50212 C9_P_btm.n599 C9_P_btm.t235 1.67819
R50213 C9_P_btm.n602 C9_P_btm.t261 1.67819
R50214 C9_P_btm.n605 C9_P_btm.t338 1.67819
R50215 C9_P_btm.n608 C9_P_btm.t525 1.67819
R50216 C9_P_btm.n611 C9_P_btm.t290 1.67819
R50217 C9_P_btm.n614 C9_P_btm.t427 1.67819
R50218 C9_P_btm.n617 C9_P_btm.t269 1.67819
R50219 C9_P_btm.n620 C9_P_btm.t375 1.67819
R50220 C9_P_btm.n623 C9_P_btm.t397 1.67819
R50221 C9_P_btm.n626 C9_P_btm.t349 1.67819
R50222 C9_P_btm.n629 C9_P_btm.t467 1.67819
R50223 C9_P_btm.n1318 C9_P_btm.n1317 1.05569
R50224 C9_P_btm.n498 C9_P_btm.n497 1.05569
R50225 C9_P_btm.n454 C9_P_btm.n425 1.05569
R50226 C9_P_btm.n632 C9_P_btm.n631 1.05569
R50227 C9_P_btm.n755 C9_P_btm.n216 1.05569
R50228 C9_P_btm.n1346 C9_P_btm.n1321 1.05569
R50229 C9_P_btm.n22 C9_P_btm.n20 1.0005
R50230 C9_P_btm.n23 C9_P_btm.n19 1.0005
R50231 C9_P_btm.n24 C9_P_btm.n18 1.0005
R50232 C9_P_btm.n1854 C9_P_btm.n17 1.0005
R50233 C9_P_btm.n1854 C9_P_btm.n1853 1.0005
R50234 C9_P_btm.n27 C9_P_btm.n24 1.0005
R50235 C9_P_btm.n28 C9_P_btm.n23 1.0005
R50236 C9_P_btm.n1840 C9_P_btm.n22 1.0005
R50237 C9_P_btm.n1840 C9_P_btm.n1839 1.0005
R50238 C9_P_btm.n1807 C9_P_btm.n28 1.0005
R50239 C9_P_btm.n1806 C9_P_btm.n27 1.0005
R50240 C9_P_btm.n1853 C9_P_btm.n25 1.0005
R50241 C9_P_btm.n34 C9_P_btm.n25 1.0005
R50242 C9_P_btm.n1806 C9_P_btm.n33 1.0005
R50243 C9_P_btm.n1807 C9_P_btm.n32 1.0005
R50244 C9_P_btm.n1839 C9_P_btm.n29 1.0005
R50245 C9_P_btm.n1788 C9_P_btm.n29 1.0005
R50246 C9_P_btm.n38 C9_P_btm.n32 1.0005
R50247 C9_P_btm.n37 C9_P_btm.n33 1.0005
R50248 C9_P_btm.n36 C9_P_btm.n34 1.0005
R50249 C9_P_btm.n56 C9_P_btm.n36 1.0005
R50250 C9_P_btm.n46 C9_P_btm.n37 1.0005
R50251 C9_P_btm.n47 C9_P_btm.n38 1.0005
R50252 C9_P_btm.n1788 C9_P_btm.n1787 1.0005
R50253 C9_P_btm.n1787 C9_P_btm.n39 1.0005
R50254 C9_P_btm.n47 C9_P_btm.n42 1.0005
R50255 C9_P_btm.n46 C9_P_btm.n43 1.0005
R50256 C9_P_btm.n57 C9_P_btm.n56 1.0005
R50257 C9_P_btm.n59 C9_P_btm.n57 1.0005
R50258 C9_P_btm.n60 C9_P_btm.n43 1.0005
R50259 C9_P_btm.n61 C9_P_btm.n42 1.0005
R50260 C9_P_btm.n1751 C9_P_btm.n39 1.0005
R50261 C9_P_btm.n1751 C9_P_btm.n1750 1.0005
R50262 C9_P_btm.n70 C9_P_btm.n61 1.0005
R50263 C9_P_btm.n69 C9_P_btm.n60 1.0005
R50264 C9_P_btm.n79 C9_P_btm.n59 1.0005
R50265 C9_P_btm.n80 C9_P_btm.n79 1.0005
R50266 C9_P_btm.n69 C9_P_btm.n66 1.0005
R50267 C9_P_btm.n70 C9_P_btm.n65 1.0005
R50268 C9_P_btm.n1750 C9_P_btm.n62 1.0005
R50269 C9_P_btm.n1714 C9_P_btm.n62 1.0005
R50270 C9_P_btm.n84 C9_P_btm.n65 1.0005
R50271 C9_P_btm.n83 C9_P_btm.n66 1.0005
R50272 C9_P_btm.n82 C9_P_btm.n80 1.0005
R50273 C9_P_btm.n102 C9_P_btm.n82 1.0005
R50274 C9_P_btm.n92 C9_P_btm.n83 1.0005
R50275 C9_P_btm.n93 C9_P_btm.n84 1.0005
R50276 C9_P_btm.n1714 C9_P_btm.n1713 1.0005
R50277 C9_P_btm.n1713 C9_P_btm.n85 1.0005
R50278 C9_P_btm.n93 C9_P_btm.n88 1.0005
R50279 C9_P_btm.n92 C9_P_btm.n89 1.0005
R50280 C9_P_btm.n103 C9_P_btm.n102 1.0005
R50281 C9_P_btm.n105 C9_P_btm.n103 1.0005
R50282 C9_P_btm.n106 C9_P_btm.n89 1.0005
R50283 C9_P_btm.n107 C9_P_btm.n88 1.0005
R50284 C9_P_btm.n1677 C9_P_btm.n85 1.0005
R50285 C9_P_btm.n1677 C9_P_btm.n1676 1.0005
R50286 C9_P_btm.n116 C9_P_btm.n107 1.0005
R50287 C9_P_btm.n115 C9_P_btm.n106 1.0005
R50288 C9_P_btm.n125 C9_P_btm.n105 1.0005
R50289 C9_P_btm.n126 C9_P_btm.n125 1.0005
R50290 C9_P_btm.n115 C9_P_btm.n112 1.0005
R50291 C9_P_btm.n116 C9_P_btm.n111 1.0005
R50292 C9_P_btm.n1676 C9_P_btm.n108 1.0005
R50293 C9_P_btm.n1639 C9_P_btm.n108 1.0005
R50294 C9_P_btm.n131 C9_P_btm.n111 1.0005
R50295 C9_P_btm.n130 C9_P_btm.n112 1.0005
R50296 C9_P_btm.n129 C9_P_btm.n126 1.0005
R50297 C9_P_btm.n1656 C9_P_btm.n1655 1.0005
R50298 C9_P_btm.n1345 C9_P_btm.n1322 1.0005
R50299 C9_P_btm.n1344 C9_P_btm.n1323 1.0005
R50300 C9_P_btm.n1343 C9_P_btm.n1324 1.0005
R50301 C9_P_btm.n1342 C9_P_btm.n1325 1.0005
R50302 C9_P_btm.n1341 C9_P_btm.n1326 1.0005
R50303 C9_P_btm.n1340 C9_P_btm.n1327 1.0005
R50304 C9_P_btm.n1339 C9_P_btm.n1328 1.0005
R50305 C9_P_btm.n1338 C9_P_btm.n1329 1.0005
R50306 C9_P_btm.n1337 C9_P_btm.n1330 1.0005
R50307 C9_P_btm.n1336 C9_P_btm.n1331 1.0005
R50308 C9_P_btm.n1335 C9_P_btm.n1332 1.0005
R50309 C9_P_btm.n1334 C9_P_btm.n1333 1.0005
R50310 C9_P_btm.n1387 C9_P_btm.n1386 1.0005
R50311 C9_P_btm.n1655 C9_P_btm.n127 1.0005
R50312 C9_P_btm.n1388 C9_P_btm.n129 1.0005
R50313 C9_P_btm.n1389 C9_P_btm.n130 1.0005
R50314 C9_P_btm.n1390 C9_P_btm.n131 1.0005
R50315 C9_P_btm.n1639 C9_P_btm.n1638 1.0005
R50316 C9_P_btm.n1638 C9_P_btm.n132 1.0005
R50317 C9_P_btm.n1390 C9_P_btm.n135 1.0005
R50318 C9_P_btm.n1389 C9_P_btm.n136 1.0005
R50319 C9_P_btm.n1388 C9_P_btm.n137 1.0005
R50320 C9_P_btm.n138 C9_P_btm.n127 1.0005
R50321 C9_P_btm.n1387 C9_P_btm.n139 1.0005
R50322 C9_P_btm.n1333 C9_P_btm.n140 1.0005
R50323 C9_P_btm.n1332 C9_P_btm.n141 1.0005
R50324 C9_P_btm.n1331 C9_P_btm.n142 1.0005
R50325 C9_P_btm.n1330 C9_P_btm.n143 1.0005
R50326 C9_P_btm.n1329 C9_P_btm.n144 1.0005
R50327 C9_P_btm.n1328 C9_P_btm.n145 1.0005
R50328 C9_P_btm.n1327 C9_P_btm.n146 1.0005
R50329 C9_P_btm.n1326 C9_P_btm.n147 1.0005
R50330 C9_P_btm.n1325 C9_P_btm.n148 1.0005
R50331 C9_P_btm.n1324 C9_P_btm.n149 1.0005
R50332 C9_P_btm.n1323 C9_P_btm.n150 1.0005
R50333 C9_P_btm.n1322 C9_P_btm.n151 1.0005
R50334 C9_P_btm.n1321 C9_P_btm.n152 1.0005
R50335 C9_P_btm.n886 C9_P_btm.n173 1.0005
R50336 C9_P_btm.n887 C9_P_btm.n172 1.0005
R50337 C9_P_btm.n888 C9_P_btm.n171 1.0005
R50338 C9_P_btm.n889 C9_P_btm.n170 1.0005
R50339 C9_P_btm.n890 C9_P_btm.n169 1.0005
R50340 C9_P_btm.n891 C9_P_btm.n168 1.0005
R50341 C9_P_btm.n892 C9_P_btm.n167 1.0005
R50342 C9_P_btm.n893 C9_P_btm.n166 1.0005
R50343 C9_P_btm.n894 C9_P_btm.n165 1.0005
R50344 C9_P_btm.n895 C9_P_btm.n164 1.0005
R50345 C9_P_btm.n896 C9_P_btm.n163 1.0005
R50346 C9_P_btm.n897 C9_P_btm.n162 1.0005
R50347 C9_P_btm.n898 C9_P_btm.n161 1.0005
R50348 C9_P_btm.n899 C9_P_btm.n160 1.0005
R50349 C9_P_btm.n900 C9_P_btm.n159 1.0005
R50350 C9_P_btm.n901 C9_P_btm.n158 1.0005
R50351 C9_P_btm.n902 C9_P_btm.n157 1.0005
R50352 C9_P_btm.n903 C9_P_btm.n156 1.0005
R50353 C9_P_btm.n904 C9_P_btm.n903 1.0005
R50354 C9_P_btm.n905 C9_P_btm.n902 1.0005
R50355 C9_P_btm.n906 C9_P_btm.n901 1.0005
R50356 C9_P_btm.n907 C9_P_btm.n900 1.0005
R50357 C9_P_btm.n908 C9_P_btm.n899 1.0005
R50358 C9_P_btm.n909 C9_P_btm.n898 1.0005
R50359 C9_P_btm.n910 C9_P_btm.n897 1.0005
R50360 C9_P_btm.n911 C9_P_btm.n896 1.0005
R50361 C9_P_btm.n912 C9_P_btm.n895 1.0005
R50362 C9_P_btm.n913 C9_P_btm.n894 1.0005
R50363 C9_P_btm.n914 C9_P_btm.n893 1.0005
R50364 C9_P_btm.n915 C9_P_btm.n892 1.0005
R50365 C9_P_btm.n916 C9_P_btm.n891 1.0005
R50366 C9_P_btm.n917 C9_P_btm.n890 1.0005
R50367 C9_P_btm.n918 C9_P_btm.n889 1.0005
R50368 C9_P_btm.n919 C9_P_btm.n888 1.0005
R50369 C9_P_btm.n920 C9_P_btm.n887 1.0005
R50370 C9_P_btm.n1261 C9_P_btm.n886 1.0005
R50371 C9_P_btm.n1261 C9_P_btm.n1260 1.0005
R50372 C9_P_btm.n923 C9_P_btm.n920 1.0005
R50373 C9_P_btm.n924 C9_P_btm.n919 1.0005
R50374 C9_P_btm.n925 C9_P_btm.n918 1.0005
R50375 C9_P_btm.n927 C9_P_btm.n925 1.0005
R50376 C9_P_btm.n928 C9_P_btm.n924 1.0005
R50377 C9_P_btm.n929 C9_P_btm.n923 1.0005
R50378 C9_P_btm.n1260 C9_P_btm.n921 1.0005
R50379 C9_P_btm.n933 C9_P_btm.n921 1.0005
R50380 C9_P_btm.n934 C9_P_btm.n929 1.0005
R50381 C9_P_btm.n935 C9_P_btm.n928 1.0005
R50382 C9_P_btm.n1215 C9_P_btm.n927 1.0005
R50383 C9_P_btm.n1215 C9_P_btm.n1214 1.0005
R50384 C9_P_btm.n944 C9_P_btm.n935 1.0005
R50385 C9_P_btm.n943 C9_P_btm.n934 1.0005
R50386 C9_P_btm.n953 C9_P_btm.n933 1.0005
R50387 C9_P_btm.n954 C9_P_btm.n953 1.0005
R50388 C9_P_btm.n943 C9_P_btm.n940 1.0005
R50389 C9_P_btm.n944 C9_P_btm.n939 1.0005
R50390 C9_P_btm.n1214 C9_P_btm.n936 1.0005
R50391 C9_P_btm.n1178 C9_P_btm.n936 1.0005
R50392 C9_P_btm.n958 C9_P_btm.n939 1.0005
R50393 C9_P_btm.n957 C9_P_btm.n940 1.0005
R50394 C9_P_btm.n956 C9_P_btm.n954 1.0005
R50395 C9_P_btm.n976 C9_P_btm.n956 1.0005
R50396 C9_P_btm.n966 C9_P_btm.n957 1.0005
R50397 C9_P_btm.n967 C9_P_btm.n958 1.0005
R50398 C9_P_btm.n1178 C9_P_btm.n1177 1.0005
R50399 C9_P_btm.n1177 C9_P_btm.n959 1.0005
R50400 C9_P_btm.n967 C9_P_btm.n962 1.0005
R50401 C9_P_btm.n966 C9_P_btm.n963 1.0005
R50402 C9_P_btm.n977 C9_P_btm.n976 1.0005
R50403 C9_P_btm.n979 C9_P_btm.n977 1.0005
R50404 C9_P_btm.n980 C9_P_btm.n963 1.0005
R50405 C9_P_btm.n981 C9_P_btm.n962 1.0005
R50406 C9_P_btm.n1141 C9_P_btm.n959 1.0005
R50407 C9_P_btm.n1141 C9_P_btm.n1140 1.0005
R50408 C9_P_btm.n990 C9_P_btm.n981 1.0005
R50409 C9_P_btm.n989 C9_P_btm.n980 1.0005
R50410 C9_P_btm.n999 C9_P_btm.n979 1.0005
R50411 C9_P_btm.n1000 C9_P_btm.n999 1.0005
R50412 C9_P_btm.n989 C9_P_btm.n986 1.0005
R50413 C9_P_btm.n990 C9_P_btm.n985 1.0005
R50414 C9_P_btm.n1140 C9_P_btm.n982 1.0005
R50415 C9_P_btm.n1104 C9_P_btm.n982 1.0005
R50416 C9_P_btm.n1004 C9_P_btm.n985 1.0005
R50417 C9_P_btm.n1003 C9_P_btm.n986 1.0005
R50418 C9_P_btm.n1002 C9_P_btm.n1000 1.0005
R50419 C9_P_btm.n1022 C9_P_btm.n1002 1.0005
R50420 C9_P_btm.n1012 C9_P_btm.n1003 1.0005
R50421 C9_P_btm.n1013 C9_P_btm.n1004 1.0005
R50422 C9_P_btm.n1104 C9_P_btm.n1103 1.0005
R50423 C9_P_btm.n1103 C9_P_btm.n1005 1.0005
R50424 C9_P_btm.n1013 C9_P_btm.n1008 1.0005
R50425 C9_P_btm.n1012 C9_P_btm.n1009 1.0005
R50426 C9_P_btm.n1023 C9_P_btm.n1022 1.0005
R50427 C9_P_btm.n1025 C9_P_btm.n1023 1.0005
R50428 C9_P_btm.n1026 C9_P_btm.n1009 1.0005
R50429 C9_P_btm.n1027 C9_P_btm.n1008 1.0005
R50430 C9_P_btm.n1067 C9_P_btm.n1005 1.0005
R50431 C9_P_btm.n1067 C9_P_btm.n1066 1.0005
R50432 C9_P_btm.n1035 C9_P_btm.n1027 1.0005
R50433 C9_P_btm.n1034 C9_P_btm.n1026 1.0005
R50434 C9_P_btm.n1044 C9_P_btm.n1025 1.0005
R50435 C9_P_btm.n1045 C9_P_btm.n1044 1.0005
R50436 C9_P_btm.n1034 C9_P_btm.n1031 1.0005
R50437 C9_P_btm.n1035 C9_P_btm.n1030 1.0005
R50438 C9_P_btm.n1066 C9_P_btm.n1028 1.0005
R50439 C9_P_btm.n1062 C9_P_btm.n1061 1.0005
R50440 C9_P_btm.n1082 C9_P_btm.n1024 1.0005
R50441 C9_P_btm.n1046 C9_P_btm.n1024 1.0005
R50442 C9_P_btm.n1098 C9_P_btm.n1007 1.0005
R50443 C9_P_btm.n1062 C9_P_btm.n1007 1.0005
R50444 C9_P_btm.n1083 C9_P_btm.n1001 1.0005
R50445 C9_P_btm.n1083 C9_P_btm.n1082 1.0005
R50446 C9_P_btm.n1099 C9_P_btm.n984 1.0005
R50447 C9_P_btm.n1099 C9_P_btm.n1098 1.0005
R50448 C9_P_btm.n1120 C9_P_btm.n1119 1.0005
R50449 C9_P_btm.n1119 C9_P_btm.n1001 1.0005
R50450 C9_P_btm.n1136 C9_P_btm.n1135 1.0005
R50451 C9_P_btm.n1135 C9_P_btm.n984 1.0005
R50452 C9_P_btm.n1156 C9_P_btm.n978 1.0005
R50453 C9_P_btm.n1120 C9_P_btm.n978 1.0005
R50454 C9_P_btm.n1172 C9_P_btm.n961 1.0005
R50455 C9_P_btm.n1136 C9_P_btm.n961 1.0005
R50456 C9_P_btm.n1157 C9_P_btm.n955 1.0005
R50457 C9_P_btm.n1157 C9_P_btm.n1156 1.0005
R50458 C9_P_btm.n1173 C9_P_btm.n938 1.0005
R50459 C9_P_btm.n1173 C9_P_btm.n1172 1.0005
R50460 C9_P_btm.n1194 C9_P_btm.n1193 1.0005
R50461 C9_P_btm.n1193 C9_P_btm.n955 1.0005
R50462 C9_P_btm.n1210 C9_P_btm.n1209 1.0005
R50463 C9_P_btm.n1209 C9_P_btm.n938 1.0005
R50464 C9_P_btm.n1230 C9_P_btm.n932 1.0005
R50465 C9_P_btm.n1194 C9_P_btm.n932 1.0005
R50466 C9_P_btm.n1246 C9_P_btm.n926 1.0005
R50467 C9_P_btm.n1210 C9_P_btm.n926 1.0005
R50468 C9_P_btm.n1231 C9_P_btm.n931 1.0005
R50469 C9_P_btm.n1231 C9_P_btm.n1230 1.0005
R50470 C9_P_btm.n1247 C9_P_btm.n917 1.0005
R50471 C9_P_btm.n1247 C9_P_btm.n1246 1.0005
R50472 C9_P_btm.n1509 C9_P_btm.n885 1.0005
R50473 C9_P_btm.n931 C9_P_btm.n885 1.0005
R50474 C9_P_btm.n1318 C9_P_btm.n155 1.0005
R50475 C9_P_btm.n1319 C9_P_btm.n154 1.0005
R50476 C9_P_btm.n1320 C9_P_btm.n153 1.0005
R50477 C9_P_btm.n175 C9_P_btm.n173 1.0005
R50478 C9_P_btm.n176 C9_P_btm.n172 1.0005
R50479 C9_P_btm.n177 C9_P_btm.n171 1.0005
R50480 C9_P_btm.n178 C9_P_btm.n170 1.0005
R50481 C9_P_btm.n179 C9_P_btm.n169 1.0005
R50482 C9_P_btm.n180 C9_P_btm.n168 1.0005
R50483 C9_P_btm.n181 C9_P_btm.n167 1.0005
R50484 C9_P_btm.n182 C9_P_btm.n166 1.0005
R50485 C9_P_btm.n183 C9_P_btm.n165 1.0005
R50486 C9_P_btm.n184 C9_P_btm.n164 1.0005
R50487 C9_P_btm.n185 C9_P_btm.n163 1.0005
R50488 C9_P_btm.n186 C9_P_btm.n162 1.0005
R50489 C9_P_btm.n187 C9_P_btm.n161 1.0005
R50490 C9_P_btm.n188 C9_P_btm.n160 1.0005
R50491 C9_P_btm.n189 C9_P_btm.n159 1.0005
R50492 C9_P_btm.n190 C9_P_btm.n158 1.0005
R50493 C9_P_btm.n191 C9_P_btm.n157 1.0005
R50494 C9_P_btm.n192 C9_P_btm.n156 1.0005
R50495 C9_P_btm.n193 C9_P_btm.n155 1.0005
R50496 C9_P_btm.n194 C9_P_btm.n154 1.0005
R50497 C9_P_btm.n195 C9_P_btm.n153 1.0005
R50498 C9_P_btm.n196 C9_P_btm.n152 1.0005
R50499 C9_P_btm.n197 C9_P_btm.n151 1.0005
R50500 C9_P_btm.n198 C9_P_btm.n150 1.0005
R50501 C9_P_btm.n199 C9_P_btm.n149 1.0005
R50502 C9_P_btm.n200 C9_P_btm.n148 1.0005
R50503 C9_P_btm.n201 C9_P_btm.n147 1.0005
R50504 C9_P_btm.n202 C9_P_btm.n146 1.0005
R50505 C9_P_btm.n203 C9_P_btm.n145 1.0005
R50506 C9_P_btm.n204 C9_P_btm.n144 1.0005
R50507 C9_P_btm.n205 C9_P_btm.n143 1.0005
R50508 C9_P_btm.n206 C9_P_btm.n142 1.0005
R50509 C9_P_btm.n207 C9_P_btm.n141 1.0005
R50510 C9_P_btm.n208 C9_P_btm.n140 1.0005
R50511 C9_P_btm.n209 C9_P_btm.n139 1.0005
R50512 C9_P_btm.n210 C9_P_btm.n138 1.0005
R50513 C9_P_btm.n211 C9_P_btm.n137 1.0005
R50514 C9_P_btm.n212 C9_P_btm.n136 1.0005
R50515 C9_P_btm.n213 C9_P_btm.n135 1.0005
R50516 C9_P_btm.n761 C9_P_btm.n132 1.0005
R50517 C9_P_btm.n761 C9_P_btm.n760 1.0005
R50518 C9_P_btm.n294 C9_P_btm.n213 1.0005
R50519 C9_P_btm.n293 C9_P_btm.n212 1.0005
R50520 C9_P_btm.n292 C9_P_btm.n211 1.0005
R50521 C9_P_btm.n291 C9_P_btm.n210 1.0005
R50522 C9_P_btm.n290 C9_P_btm.n209 1.0005
R50523 C9_P_btm.n289 C9_P_btm.n208 1.0005
R50524 C9_P_btm.n288 C9_P_btm.n207 1.0005
R50525 C9_P_btm.n287 C9_P_btm.n206 1.0005
R50526 C9_P_btm.n286 C9_P_btm.n205 1.0005
R50527 C9_P_btm.n285 C9_P_btm.n204 1.0005
R50528 C9_P_btm.n284 C9_P_btm.n203 1.0005
R50529 C9_P_btm.n283 C9_P_btm.n202 1.0005
R50530 C9_P_btm.n282 C9_P_btm.n201 1.0005
R50531 C9_P_btm.n281 C9_P_btm.n200 1.0005
R50532 C9_P_btm.n280 C9_P_btm.n199 1.0005
R50533 C9_P_btm.n279 C9_P_btm.n198 1.0005
R50534 C9_P_btm.n278 C9_P_btm.n197 1.0005
R50535 C9_P_btm.n277 C9_P_btm.n196 1.0005
R50536 C9_P_btm.n276 C9_P_btm.n195 1.0005
R50537 C9_P_btm.n275 C9_P_btm.n194 1.0005
R50538 C9_P_btm.n274 C9_P_btm.n193 1.0005
R50539 C9_P_btm.n273 C9_P_btm.n192 1.0005
R50540 C9_P_btm.n272 C9_P_btm.n191 1.0005
R50541 C9_P_btm.n271 C9_P_btm.n190 1.0005
R50542 C9_P_btm.n270 C9_P_btm.n189 1.0005
R50543 C9_P_btm.n269 C9_P_btm.n188 1.0005
R50544 C9_P_btm.n268 C9_P_btm.n187 1.0005
R50545 C9_P_btm.n267 C9_P_btm.n186 1.0005
R50546 C9_P_btm.n266 C9_P_btm.n185 1.0005
R50547 C9_P_btm.n265 C9_P_btm.n184 1.0005
R50548 C9_P_btm.n264 C9_P_btm.n183 1.0005
R50549 C9_P_btm.n263 C9_P_btm.n182 1.0005
R50550 C9_P_btm.n262 C9_P_btm.n181 1.0005
R50551 C9_P_btm.n261 C9_P_btm.n180 1.0005
R50552 C9_P_btm.n260 C9_P_btm.n179 1.0005
R50553 C9_P_btm.n259 C9_P_btm.n178 1.0005
R50554 C9_P_btm.n258 C9_P_btm.n177 1.0005
R50555 C9_P_btm.n257 C9_P_btm.n176 1.0005
R50556 C9_P_btm.n411 C9_P_btm.n175 1.0005
R50557 C9_P_btm.n412 C9_P_btm.n411 1.0005
R50558 C9_P_btm.n257 C9_P_btm.n254 1.0005
R50559 C9_P_btm.n258 C9_P_btm.n253 1.0005
R50560 C9_P_btm.n259 C9_P_btm.n252 1.0005
R50561 C9_P_btm.n260 C9_P_btm.n251 1.0005
R50562 C9_P_btm.n261 C9_P_btm.n250 1.0005
R50563 C9_P_btm.n262 C9_P_btm.n249 1.0005
R50564 C9_P_btm.n263 C9_P_btm.n248 1.0005
R50565 C9_P_btm.n264 C9_P_btm.n247 1.0005
R50566 C9_P_btm.n265 C9_P_btm.n246 1.0005
R50567 C9_P_btm.n266 C9_P_btm.n245 1.0005
R50568 C9_P_btm.n267 C9_P_btm.n244 1.0005
R50569 C9_P_btm.n268 C9_P_btm.n243 1.0005
R50570 C9_P_btm.n269 C9_P_btm.n242 1.0005
R50571 C9_P_btm.n270 C9_P_btm.n241 1.0005
R50572 C9_P_btm.n271 C9_P_btm.n240 1.0005
R50573 C9_P_btm.n272 C9_P_btm.n239 1.0005
R50574 C9_P_btm.n273 C9_P_btm.n238 1.0005
R50575 C9_P_btm.n274 C9_P_btm.n237 1.0005
R50576 C9_P_btm.n275 C9_P_btm.n236 1.0005
R50577 C9_P_btm.n276 C9_P_btm.n235 1.0005
R50578 C9_P_btm.n277 C9_P_btm.n234 1.0005
R50579 C9_P_btm.n278 C9_P_btm.n233 1.0005
R50580 C9_P_btm.n279 C9_P_btm.n232 1.0005
R50581 C9_P_btm.n280 C9_P_btm.n231 1.0005
R50582 C9_P_btm.n281 C9_P_btm.n230 1.0005
R50583 C9_P_btm.n282 C9_P_btm.n229 1.0005
R50584 C9_P_btm.n283 C9_P_btm.n228 1.0005
R50585 C9_P_btm.n284 C9_P_btm.n227 1.0005
R50586 C9_P_btm.n285 C9_P_btm.n226 1.0005
R50587 C9_P_btm.n286 C9_P_btm.n225 1.0005
R50588 C9_P_btm.n287 C9_P_btm.n224 1.0005
R50589 C9_P_btm.n288 C9_P_btm.n223 1.0005
R50590 C9_P_btm.n289 C9_P_btm.n222 1.0005
R50591 C9_P_btm.n290 C9_P_btm.n221 1.0005
R50592 C9_P_btm.n291 C9_P_btm.n220 1.0005
R50593 C9_P_btm.n292 C9_P_btm.n219 1.0005
R50594 C9_P_btm.n293 C9_P_btm.n218 1.0005
R50595 C9_P_btm.n294 C9_P_btm.n217 1.0005
R50596 C9_P_btm.n760 C9_P_btm.n214 1.0005
R50597 C9_P_btm.n510 C9_P_btm.n214 1.0005
R50598 C9_P_btm.n509 C9_P_btm.n217 1.0005
R50599 C9_P_btm.n508 C9_P_btm.n218 1.0005
R50600 C9_P_btm.n507 C9_P_btm.n219 1.0005
R50601 C9_P_btm.n506 C9_P_btm.n220 1.0005
R50602 C9_P_btm.n505 C9_P_btm.n221 1.0005
R50603 C9_P_btm.n504 C9_P_btm.n222 1.0005
R50604 C9_P_btm.n503 C9_P_btm.n223 1.0005
R50605 C9_P_btm.n502 C9_P_btm.n224 1.0005
R50606 C9_P_btm.n501 C9_P_btm.n225 1.0005
R50607 C9_P_btm.n500 C9_P_btm.n226 1.0005
R50608 C9_P_btm.n499 C9_P_btm.n227 1.0005
R50609 C9_P_btm.n498 C9_P_btm.n228 1.0005
R50610 C9_P_btm.n439 C9_P_btm.n229 1.0005
R50611 C9_P_btm.n438 C9_P_btm.n230 1.0005
R50612 C9_P_btm.n437 C9_P_btm.n231 1.0005
R50613 C9_P_btm.n436 C9_P_btm.n232 1.0005
R50614 C9_P_btm.n435 C9_P_btm.n233 1.0005
R50615 C9_P_btm.n434 C9_P_btm.n234 1.0005
R50616 C9_P_btm.n433 C9_P_btm.n235 1.0005
R50617 C9_P_btm.n432 C9_P_btm.n236 1.0005
R50618 C9_P_btm.n431 C9_P_btm.n237 1.0005
R50619 C9_P_btm.n430 C9_P_btm.n238 1.0005
R50620 C9_P_btm.n429 C9_P_btm.n239 1.0005
R50621 C9_P_btm.n428 C9_P_btm.n240 1.0005
R50622 C9_P_btm.n427 C9_P_btm.n241 1.0005
R50623 C9_P_btm.n426 C9_P_btm.n242 1.0005
R50624 C9_P_btm.n453 C9_P_btm.n426 1.0005
R50625 C9_P_btm.n452 C9_P_btm.n427 1.0005
R50626 C9_P_btm.n451 C9_P_btm.n428 1.0005
R50627 C9_P_btm.n450 C9_P_btm.n429 1.0005
R50628 C9_P_btm.n449 C9_P_btm.n430 1.0005
R50629 C9_P_btm.n448 C9_P_btm.n431 1.0005
R50630 C9_P_btm.n447 C9_P_btm.n432 1.0005
R50631 C9_P_btm.n446 C9_P_btm.n433 1.0005
R50632 C9_P_btm.n445 C9_P_btm.n434 1.0005
R50633 C9_P_btm.n444 C9_P_btm.n435 1.0005
R50634 C9_P_btm.n443 C9_P_btm.n436 1.0005
R50635 C9_P_btm.n442 C9_P_btm.n437 1.0005
R50636 C9_P_btm.n441 C9_P_btm.n438 1.0005
R50637 C9_P_btm.n440 C9_P_btm.n439 1.0005
R50638 C9_P_btm.n425 C9_P_btm.n243 1.0005
R50639 C9_P_btm.n424 C9_P_btm.n244 1.0005
R50640 C9_P_btm.n423 C9_P_btm.n245 1.0005
R50641 C9_P_btm.n422 C9_P_btm.n246 1.0005
R50642 C9_P_btm.n421 C9_P_btm.n247 1.0005
R50643 C9_P_btm.n420 C9_P_btm.n248 1.0005
R50644 C9_P_btm.n419 C9_P_btm.n249 1.0005
R50645 C9_P_btm.n418 C9_P_btm.n250 1.0005
R50646 C9_P_btm.n417 C9_P_btm.n251 1.0005
R50647 C9_P_btm.n416 C9_P_btm.n252 1.0005
R50648 C9_P_btm.n415 C9_P_btm.n253 1.0005
R50649 C9_P_btm.n414 C9_P_btm.n254 1.0005
R50650 C9_P_btm.n413 C9_P_btm.n412 1.0005
R50651 C9_P_btm.n756 C9_P_btm.n755 1.0005
R50652 C9_P_btm.n632 C9_P_btm.n174 1.0005
R50653 C9_P_btm.n884 C9_P_btm.n174 1.0005
R50654 C9_P_btm.n756 C9_P_btm.n134 1.0005
R50655 C9_P_btm.n1633 C9_P_btm.n134 1.0005
R50656 C9_P_btm.n1510 C9_P_btm.n884 1.0005
R50657 C9_P_btm.n1510 C9_P_btm.n1509 1.0005
R50658 C9_P_btm.n1634 C9_P_btm.n1633 1.0005
R50659 C9_P_btm.n1634 C9_P_btm.n110 1.0005
R50660 C9_P_btm.n1671 C9_P_btm.n110 1.0005
R50661 C9_P_btm.n1672 C9_P_btm.n1671 1.0005
R50662 C9_P_btm.n1656 C9_P_btm.n104 1.0005
R50663 C9_P_btm.n1692 C9_P_btm.n104 1.0005
R50664 C9_P_btm.n1672 C9_P_btm.n87 1.0005
R50665 C9_P_btm.n1708 C9_P_btm.n87 1.0005
R50666 C9_P_btm.n1693 C9_P_btm.n1692 1.0005
R50667 C9_P_btm.n1693 C9_P_btm.n81 1.0005
R50668 C9_P_btm.n1709 C9_P_btm.n1708 1.0005
R50669 C9_P_btm.n1709 C9_P_btm.n64 1.0005
R50670 C9_P_btm.n1729 C9_P_btm.n81 1.0005
R50671 C9_P_btm.n1730 C9_P_btm.n1729 1.0005
R50672 C9_P_btm.n1745 C9_P_btm.n64 1.0005
R50673 C9_P_btm.n1746 C9_P_btm.n1745 1.0005
R50674 C9_P_btm.n1730 C9_P_btm.n58 1.0005
R50675 C9_P_btm.n1766 C9_P_btm.n58 1.0005
R50676 C9_P_btm.n1746 C9_P_btm.n41 1.0005
R50677 C9_P_btm.n1782 C9_P_btm.n41 1.0005
R50678 C9_P_btm.n1767 C9_P_btm.n1766 1.0005
R50679 C9_P_btm.n1767 C9_P_btm.n35 1.0005
R50680 C9_P_btm.n1783 C9_P_btm.n1782 1.0005
R50681 C9_P_btm.n1783 C9_P_btm.n31 1.0005
R50682 C9_P_btm.n1803 C9_P_btm.n35 1.0005
R50683 C9_P_btm.n1819 C9_P_btm.n1803 1.0005
R50684 C9_P_btm.n1834 C9_P_btm.n31 1.0005
R50685 C9_P_btm.n1835 C9_P_btm.n1834 1.0005
R50686 C9_P_btm.n1819 C9_P_btm.n1818 1.0005
R50687 C9_P_btm.n1818 C9_P_btm.n1805 1.0005
R50688 C9_P_btm.n1835 C9_P_btm.n21 1.0005
R50689 C9_P_btm.n1869 C9_P_btm.n21 1.0005
R50690 C9_P_btm.n1805 C9_P_btm.n16 1.0005
R50691 C9_P_btm.n1885 C9_P_btm.n16 1.0005
R50692 C9_P_btm.n1870 C9_P_btm.n1869 1.0005
R50693 C9_P_btm.n1886 C9_P_btm.n1885 1.0005
R50694 C9_P_btm.n4 C9_P_btm.n2 0.688
R50695 C9_P_btm.n1060 C9_P_btm.n1059 0.679419
R50696 C9_P_btm.n1048 C9_P_btm.n1047 0.679419
R50697 C9_P_btm.n1033 C9_P_btm.n1032 0.679419
R50698 C9_P_btm.n1065 C9_P_btm.n1063 0.679419
R50699 C9_P_btm.n1069 C9_P_btm.n1068 0.679419
R50700 C9_P_btm.n1081 C9_P_btm.n1080 0.679419
R50701 C9_P_btm.n1085 C9_P_btm.n1084 0.679419
R50702 C9_P_btm.n1097 C9_P_btm.n1096 0.679419
R50703 C9_P_btm.n1102 C9_P_btm.n1100 0.679419
R50704 C9_P_btm.n1011 C9_P_btm.n1010 0.679419
R50705 C9_P_btm.n1118 C9_P_btm.n1117 0.679419
R50706 C9_P_btm.n1106 C9_P_btm.n1105 0.679419
R50707 C9_P_btm.n1134 C9_P_btm.n1133 0.679419
R50708 C9_P_btm.n1122 C9_P_btm.n1121 0.679419
R50709 C9_P_btm.n988 C9_P_btm.n987 0.679419
R50710 C9_P_btm.n1139 C9_P_btm.n1137 0.679419
R50711 C9_P_btm.n1143 C9_P_btm.n1142 0.679419
R50712 C9_P_btm.n1155 C9_P_btm.n1154 0.679419
R50713 C9_P_btm.n1159 C9_P_btm.n1158 0.679419
R50714 C9_P_btm.n1171 C9_P_btm.n1170 0.679419
R50715 C9_P_btm.n1176 C9_P_btm.n1174 0.679419
R50716 C9_P_btm.n965 C9_P_btm.n964 0.679419
R50717 C9_P_btm.n1192 C9_P_btm.n1191 0.679419
R50718 C9_P_btm.n1180 C9_P_btm.n1179 0.679419
R50719 C9_P_btm.n1208 C9_P_btm.n1207 0.679419
R50720 C9_P_btm.n1196 C9_P_btm.n1195 0.679419
R50721 C9_P_btm.n942 C9_P_btm.n941 0.679419
R50722 C9_P_btm.n1213 C9_P_btm.n1211 0.679419
R50723 C9_P_btm.n1217 C9_P_btm.n1216 0.679419
R50724 C9_P_btm.n1229 C9_P_btm.n1228 0.679419
R50725 C9_P_btm.n1233 C9_P_btm.n1232 0.679419
R50726 C9_P_btm.n1245 C9_P_btm.n1244 0.679419
R50727 C9_P_btm.n1249 C9_P_btm.n1248 0.679419
R50728 C9_P_btm.n930 C9_P_btm.n922 0.679419
R50729 C9_P_btm.n1263 C9_P_btm.n1262 0.679419
R50730 C9_P_btm.n1317 C9_P_btm.n1316 0.679419
R50731 C9_P_btm.n1508 C9_P_btm.n1507 0.679419
R50732 C9_P_btm.n497 C9_P_btm.n496 0.679419
R50733 C9_P_btm.n455 C9_P_btm.n454 0.679419
R50734 C9_P_btm.n631 C9_P_btm.n630 0.679419
R50735 C9_P_btm.n511 C9_P_btm.n216 0.679419
R50736 C9_P_btm.n754 C9_P_btm.n753 0.679419
R50737 C9_P_btm.n634 C9_P_btm.n633 0.679419
R50738 C9_P_btm.n256 C9_P_btm.n255 0.679419
R50739 C9_P_btm.n759 C9_P_btm.n757 0.679419
R50740 C9_P_btm.n763 C9_P_btm.n762 0.679419
R50741 C9_P_btm.n883 C9_P_btm.n882 0.679419
R50742 C9_P_btm.n1512 C9_P_btm.n1511 0.679419
R50743 C9_P_btm.n1632 C9_P_btm.n1631 0.679419
R50744 C9_P_btm.n1637 C9_P_btm.n1635 0.679419
R50745 C9_P_btm.n1347 C9_P_btm.n1346 0.679419
R50746 C9_P_btm.n1641 C9_P_btm.n1640 0.679419
R50747 C9_P_btm.n1670 C9_P_btm.n1669 0.679419
R50748 C9_P_btm.n1658 C9_P_btm.n1657 0.679419
R50749 C9_P_btm.n114 C9_P_btm.n113 0.679419
R50750 C9_P_btm.n1675 C9_P_btm.n1673 0.679419
R50751 C9_P_btm.n1679 C9_P_btm.n1678 0.679419
R50752 C9_P_btm.n1691 C9_P_btm.n1690 0.679419
R50753 C9_P_btm.n1695 C9_P_btm.n1694 0.679419
R50754 C9_P_btm.n1707 C9_P_btm.n1706 0.679419
R50755 C9_P_btm.n1712 C9_P_btm.n1710 0.679419
R50756 C9_P_btm.n91 C9_P_btm.n90 0.679419
R50757 C9_P_btm.n1728 C9_P_btm.n1727 0.679419
R50758 C9_P_btm.n1716 C9_P_btm.n1715 0.679419
R50759 C9_P_btm.n1744 C9_P_btm.n1743 0.679419
R50760 C9_P_btm.n1732 C9_P_btm.n1731 0.679419
R50761 C9_P_btm.n68 C9_P_btm.n67 0.679419
R50762 C9_P_btm.n1749 C9_P_btm.n1747 0.679419
R50763 C9_P_btm.n1753 C9_P_btm.n1752 0.679419
R50764 C9_P_btm.n1765 C9_P_btm.n1764 0.679419
R50765 C9_P_btm.n1769 C9_P_btm.n1768 0.679419
R50766 C9_P_btm.n1781 C9_P_btm.n1780 0.679419
R50767 C9_P_btm.n1786 C9_P_btm.n1784 0.679419
R50768 C9_P_btm.n45 C9_P_btm.n44 0.679419
R50769 C9_P_btm.n1802 C9_P_btm.n1801 0.679419
R50770 C9_P_btm.n1790 C9_P_btm.n1789 0.679419
R50771 C9_P_btm.n1833 C9_P_btm.n1832 0.679419
R50772 C9_P_btm.n1821 C9_P_btm.n1820 0.679419
R50773 C9_P_btm.n1817 C9_P_btm.n1816 0.679419
R50774 C9_P_btm.n1838 C9_P_btm.n1836 0.679419
R50775 C9_P_btm.n1842 C9_P_btm.n1841 0.679419
R50776 C9_P_btm.n1804 C9_P_btm.n26 0.679419
R50777 C9_P_btm.n1856 C9_P_btm.n1855 0.679419
R50778 C9_P_btm.n1868 C9_P_btm.n1867 0.679419
R50779 C9_P_btm.n1872 C9_P_btm.n1871 0.679419
R50780 C9_P_btm.n1884 C9_P_btm.n1883 0.679419
R50781 C9_P_btm.n6 C9_P_btm.n4 0.672375
R50782 C9_P_btm.n1057 C9_P_btm.n1056 0.6255
R50783 C9_P_btm.n1054 C9_P_btm.n1053 0.6255
R50784 C9_P_btm.n1051 C9_P_btm.n1050 0.6255
R50785 C9_P_btm.n1043 C9_P_btm.n1041 0.6255
R50786 C9_P_btm.n1039 C9_P_btm.n1038 0.6255
R50787 C9_P_btm.n1036 C9_P_btm.n1029 0.6255
R50788 C9_P_btm.n1072 C9_P_btm.n1071 0.6255
R50789 C9_P_btm.n1075 C9_P_btm.n1074 0.6255
R50790 C9_P_btm.n1078 C9_P_btm.n1077 0.6255
R50791 C9_P_btm.n1088 C9_P_btm.n1087 0.6255
R50792 C9_P_btm.n1091 C9_P_btm.n1090 0.6255
R50793 C9_P_btm.n1094 C9_P_btm.n1093 0.6255
R50794 C9_P_btm.n1014 C9_P_btm.n1006 0.6255
R50795 C9_P_btm.n1017 C9_P_btm.n1016 0.6255
R50796 C9_P_btm.n1021 C9_P_btm.n1019 0.6255
R50797 C9_P_btm.n1115 C9_P_btm.n1114 0.6255
R50798 C9_P_btm.n1112 C9_P_btm.n1111 0.6255
R50799 C9_P_btm.n1109 C9_P_btm.n1108 0.6255
R50800 C9_P_btm.n1131 C9_P_btm.n1130 0.6255
R50801 C9_P_btm.n1128 C9_P_btm.n1127 0.6255
R50802 C9_P_btm.n1125 C9_P_btm.n1124 0.6255
R50803 C9_P_btm.n998 C9_P_btm.n996 0.6255
R50804 C9_P_btm.n994 C9_P_btm.n993 0.6255
R50805 C9_P_btm.n991 C9_P_btm.n983 0.6255
R50806 C9_P_btm.n1146 C9_P_btm.n1145 0.6255
R50807 C9_P_btm.n1149 C9_P_btm.n1148 0.6255
R50808 C9_P_btm.n1152 C9_P_btm.n1151 0.6255
R50809 C9_P_btm.n1162 C9_P_btm.n1161 0.6255
R50810 C9_P_btm.n1165 C9_P_btm.n1164 0.6255
R50811 C9_P_btm.n1168 C9_P_btm.n1167 0.6255
R50812 C9_P_btm.n968 C9_P_btm.n960 0.6255
R50813 C9_P_btm.n971 C9_P_btm.n970 0.6255
R50814 C9_P_btm.n975 C9_P_btm.n973 0.6255
R50815 C9_P_btm.n1189 C9_P_btm.n1188 0.6255
R50816 C9_P_btm.n1186 C9_P_btm.n1185 0.6255
R50817 C9_P_btm.n1183 C9_P_btm.n1182 0.6255
R50818 C9_P_btm.n1205 C9_P_btm.n1204 0.6255
R50819 C9_P_btm.n1202 C9_P_btm.n1201 0.6255
R50820 C9_P_btm.n1199 C9_P_btm.n1198 0.6255
R50821 C9_P_btm.n952 C9_P_btm.n950 0.6255
R50822 C9_P_btm.n948 C9_P_btm.n947 0.6255
R50823 C9_P_btm.n945 C9_P_btm.n937 0.6255
R50824 C9_P_btm.n1220 C9_P_btm.n1219 0.6255
R50825 C9_P_btm.n1223 C9_P_btm.n1222 0.6255
R50826 C9_P_btm.n1226 C9_P_btm.n1225 0.6255
R50827 C9_P_btm.n1236 C9_P_btm.n1235 0.6255
R50828 C9_P_btm.n1239 C9_P_btm.n1238 0.6255
R50829 C9_P_btm.n1242 C9_P_btm.n1241 0.6255
R50830 C9_P_btm.n1252 C9_P_btm.n1251 0.6255
R50831 C9_P_btm.n1255 C9_P_btm.n1254 0.6255
R50832 C9_P_btm.n1259 C9_P_btm.n1257 0.6255
R50833 C9_P_btm.n1266 C9_P_btm.n1265 0.6255
R50834 C9_P_btm.n1269 C9_P_btm.n1268 0.6255
R50835 C9_P_btm.n1272 C9_P_btm.n1271 0.6255
R50836 C9_P_btm.n1275 C9_P_btm.n1274 0.6255
R50837 C9_P_btm.n1278 C9_P_btm.n1277 0.6255
R50838 C9_P_btm.n1281 C9_P_btm.n1280 0.6255
R50839 C9_P_btm.n1284 C9_P_btm.n1283 0.6255
R50840 C9_P_btm.n1287 C9_P_btm.n1286 0.6255
R50841 C9_P_btm.n1290 C9_P_btm.n1289 0.6255
R50842 C9_P_btm.n1293 C9_P_btm.n1292 0.6255
R50843 C9_P_btm.n1296 C9_P_btm.n1295 0.6255
R50844 C9_P_btm.n1299 C9_P_btm.n1298 0.6255
R50845 C9_P_btm.n1302 C9_P_btm.n1301 0.6255
R50846 C9_P_btm.n1305 C9_P_btm.n1304 0.6255
R50847 C9_P_btm.n1308 C9_P_btm.n1307 0.6255
R50848 C9_P_btm.n1311 C9_P_btm.n1310 0.6255
R50849 C9_P_btm.n1314 C9_P_btm.n1313 0.6255
R50850 C9_P_btm.n1445 C9_P_btm.n1444 0.6255
R50851 C9_P_btm.n1448 C9_P_btm.n1447 0.6255
R50852 C9_P_btm.n1451 C9_P_btm.n1450 0.6255
R50853 C9_P_btm.n1454 C9_P_btm.n1453 0.6255
R50854 C9_P_btm.n1457 C9_P_btm.n1456 0.6255
R50855 C9_P_btm.n1460 C9_P_btm.n1459 0.6255
R50856 C9_P_btm.n1463 C9_P_btm.n1462 0.6255
R50857 C9_P_btm.n1466 C9_P_btm.n1465 0.6255
R50858 C9_P_btm.n1469 C9_P_btm.n1468 0.6255
R50859 C9_P_btm.n1472 C9_P_btm.n1471 0.6255
R50860 C9_P_btm.n1475 C9_P_btm.n1474 0.6255
R50861 C9_P_btm.n1478 C9_P_btm.n1477 0.6255
R50862 C9_P_btm.n1481 C9_P_btm.n1480 0.6255
R50863 C9_P_btm.n1484 C9_P_btm.n1483 0.6255
R50864 C9_P_btm.n1487 C9_P_btm.n1486 0.6255
R50865 C9_P_btm.n1490 C9_P_btm.n1489 0.6255
R50866 C9_P_btm.n1493 C9_P_btm.n1492 0.6255
R50867 C9_P_btm.n1496 C9_P_btm.n1495 0.6255
R50868 C9_P_btm.n1499 C9_P_btm.n1498 0.6255
R50869 C9_P_btm.n1502 C9_P_btm.n1501 0.6255
R50870 C9_P_btm.n1505 C9_P_btm.n1504 0.6255
R50871 C9_P_btm.n494 C9_P_btm.n493 0.6255
R50872 C9_P_btm.n491 C9_P_btm.n490 0.6255
R50873 C9_P_btm.n488 C9_P_btm.n487 0.6255
R50874 C9_P_btm.n485 C9_P_btm.n484 0.6255
R50875 C9_P_btm.n482 C9_P_btm.n481 0.6255
R50876 C9_P_btm.n479 C9_P_btm.n478 0.6255
R50877 C9_P_btm.n476 C9_P_btm.n475 0.6255
R50878 C9_P_btm.n473 C9_P_btm.n472 0.6255
R50879 C9_P_btm.n470 C9_P_btm.n469 0.6255
R50880 C9_P_btm.n467 C9_P_btm.n466 0.6255
R50881 C9_P_btm.n464 C9_P_btm.n463 0.6255
R50882 C9_P_btm.n461 C9_P_btm.n460 0.6255
R50883 C9_P_btm.n458 C9_P_btm.n457 0.6255
R50884 C9_P_btm.n628 C9_P_btm.n627 0.6255
R50885 C9_P_btm.n625 C9_P_btm.n624 0.6255
R50886 C9_P_btm.n622 C9_P_btm.n621 0.6255
R50887 C9_P_btm.n619 C9_P_btm.n618 0.6255
R50888 C9_P_btm.n616 C9_P_btm.n615 0.6255
R50889 C9_P_btm.n613 C9_P_btm.n612 0.6255
R50890 C9_P_btm.n610 C9_P_btm.n609 0.6255
R50891 C9_P_btm.n607 C9_P_btm.n606 0.6255
R50892 C9_P_btm.n604 C9_P_btm.n603 0.6255
R50893 C9_P_btm.n601 C9_P_btm.n600 0.6255
R50894 C9_P_btm.n598 C9_P_btm.n597 0.6255
R50895 C9_P_btm.n595 C9_P_btm.n594 0.6255
R50896 C9_P_btm.n592 C9_P_btm.n591 0.6255
R50897 C9_P_btm.n589 C9_P_btm.n588 0.6255
R50898 C9_P_btm.n586 C9_P_btm.n585 0.6255
R50899 C9_P_btm.n583 C9_P_btm.n582 0.6255
R50900 C9_P_btm.n580 C9_P_btm.n579 0.6255
R50901 C9_P_btm.n577 C9_P_btm.n576 0.6255
R50902 C9_P_btm.n574 C9_P_btm.n573 0.6255
R50903 C9_P_btm.n571 C9_P_btm.n570 0.6255
R50904 C9_P_btm.n568 C9_P_btm.n567 0.6255
R50905 C9_P_btm.n565 C9_P_btm.n564 0.6255
R50906 C9_P_btm.n562 C9_P_btm.n561 0.6255
R50907 C9_P_btm.n559 C9_P_btm.n558 0.6255
R50908 C9_P_btm.n556 C9_P_btm.n555 0.6255
R50909 C9_P_btm.n553 C9_P_btm.n552 0.6255
R50910 C9_P_btm.n550 C9_P_btm.n549 0.6255
R50911 C9_P_btm.n547 C9_P_btm.n546 0.6255
R50912 C9_P_btm.n544 C9_P_btm.n543 0.6255
R50913 C9_P_btm.n541 C9_P_btm.n540 0.6255
R50914 C9_P_btm.n538 C9_P_btm.n537 0.6255
R50915 C9_P_btm.n535 C9_P_btm.n534 0.6255
R50916 C9_P_btm.n532 C9_P_btm.n531 0.6255
R50917 C9_P_btm.n529 C9_P_btm.n528 0.6255
R50918 C9_P_btm.n526 C9_P_btm.n525 0.6255
R50919 C9_P_btm.n523 C9_P_btm.n522 0.6255
R50920 C9_P_btm.n520 C9_P_btm.n519 0.6255
R50921 C9_P_btm.n517 C9_P_btm.n516 0.6255
R50922 C9_P_btm.n514 C9_P_btm.n513 0.6255
R50923 C9_P_btm.n751 C9_P_btm.n750 0.6255
R50924 C9_P_btm.n748 C9_P_btm.n747 0.6255
R50925 C9_P_btm.n745 C9_P_btm.n744 0.6255
R50926 C9_P_btm.n742 C9_P_btm.n741 0.6255
R50927 C9_P_btm.n739 C9_P_btm.n738 0.6255
R50928 C9_P_btm.n736 C9_P_btm.n735 0.6255
R50929 C9_P_btm.n733 C9_P_btm.n732 0.6255
R50930 C9_P_btm.n730 C9_P_btm.n729 0.6255
R50931 C9_P_btm.n727 C9_P_btm.n726 0.6255
R50932 C9_P_btm.n724 C9_P_btm.n723 0.6255
R50933 C9_P_btm.n721 C9_P_btm.n720 0.6255
R50934 C9_P_btm.n718 C9_P_btm.n717 0.6255
R50935 C9_P_btm.n715 C9_P_btm.n714 0.6255
R50936 C9_P_btm.n712 C9_P_btm.n711 0.6255
R50937 C9_P_btm.n709 C9_P_btm.n708 0.6255
R50938 C9_P_btm.n706 C9_P_btm.n705 0.6255
R50939 C9_P_btm.n703 C9_P_btm.n702 0.6255
R50940 C9_P_btm.n700 C9_P_btm.n699 0.6255
R50941 C9_P_btm.n697 C9_P_btm.n696 0.6255
R50942 C9_P_btm.n694 C9_P_btm.n693 0.6255
R50943 C9_P_btm.n691 C9_P_btm.n690 0.6255
R50944 C9_P_btm.n688 C9_P_btm.n687 0.6255
R50945 C9_P_btm.n685 C9_P_btm.n684 0.6255
R50946 C9_P_btm.n682 C9_P_btm.n681 0.6255
R50947 C9_P_btm.n679 C9_P_btm.n678 0.6255
R50948 C9_P_btm.n676 C9_P_btm.n675 0.6255
R50949 C9_P_btm.n673 C9_P_btm.n672 0.6255
R50950 C9_P_btm.n670 C9_P_btm.n669 0.6255
R50951 C9_P_btm.n667 C9_P_btm.n666 0.6255
R50952 C9_P_btm.n664 C9_P_btm.n663 0.6255
R50953 C9_P_btm.n661 C9_P_btm.n660 0.6255
R50954 C9_P_btm.n658 C9_P_btm.n657 0.6255
R50955 C9_P_btm.n655 C9_P_btm.n654 0.6255
R50956 C9_P_btm.n652 C9_P_btm.n651 0.6255
R50957 C9_P_btm.n649 C9_P_btm.n648 0.6255
R50958 C9_P_btm.n646 C9_P_btm.n645 0.6255
R50959 C9_P_btm.n643 C9_P_btm.n642 0.6255
R50960 C9_P_btm.n640 C9_P_btm.n639 0.6255
R50961 C9_P_btm.n637 C9_P_btm.n636 0.6255
R50962 C9_P_btm.n410 C9_P_btm.n408 0.6255
R50963 C9_P_btm.n406 C9_P_btm.n405 0.6255
R50964 C9_P_btm.n403 C9_P_btm.n402 0.6255
R50965 C9_P_btm.n400 C9_P_btm.n399 0.6255
R50966 C9_P_btm.n397 C9_P_btm.n396 0.6255
R50967 C9_P_btm.n394 C9_P_btm.n393 0.6255
R50968 C9_P_btm.n391 C9_P_btm.n390 0.6255
R50969 C9_P_btm.n388 C9_P_btm.n387 0.6255
R50970 C9_P_btm.n385 C9_P_btm.n384 0.6255
R50971 C9_P_btm.n382 C9_P_btm.n381 0.6255
R50972 C9_P_btm.n379 C9_P_btm.n378 0.6255
R50973 C9_P_btm.n376 C9_P_btm.n375 0.6255
R50974 C9_P_btm.n373 C9_P_btm.n372 0.6255
R50975 C9_P_btm.n370 C9_P_btm.n369 0.6255
R50976 C9_P_btm.n367 C9_P_btm.n366 0.6255
R50977 C9_P_btm.n364 C9_P_btm.n363 0.6255
R50978 C9_P_btm.n361 C9_P_btm.n360 0.6255
R50979 C9_P_btm.n358 C9_P_btm.n357 0.6255
R50980 C9_P_btm.n355 C9_P_btm.n354 0.6255
R50981 C9_P_btm.n352 C9_P_btm.n351 0.6255
R50982 C9_P_btm.n349 C9_P_btm.n348 0.6255
R50983 C9_P_btm.n346 C9_P_btm.n345 0.6255
R50984 C9_P_btm.n343 C9_P_btm.n342 0.6255
R50985 C9_P_btm.n340 C9_P_btm.n339 0.6255
R50986 C9_P_btm.n337 C9_P_btm.n336 0.6255
R50987 C9_P_btm.n334 C9_P_btm.n333 0.6255
R50988 C9_P_btm.n331 C9_P_btm.n330 0.6255
R50989 C9_P_btm.n328 C9_P_btm.n327 0.6255
R50990 C9_P_btm.n325 C9_P_btm.n324 0.6255
R50991 C9_P_btm.n322 C9_P_btm.n321 0.6255
R50992 C9_P_btm.n319 C9_P_btm.n318 0.6255
R50993 C9_P_btm.n316 C9_P_btm.n315 0.6255
R50994 C9_P_btm.n313 C9_P_btm.n312 0.6255
R50995 C9_P_btm.n310 C9_P_btm.n309 0.6255
R50996 C9_P_btm.n307 C9_P_btm.n306 0.6255
R50997 C9_P_btm.n304 C9_P_btm.n303 0.6255
R50998 C9_P_btm.n301 C9_P_btm.n300 0.6255
R50999 C9_P_btm.n298 C9_P_btm.n297 0.6255
R51000 C9_P_btm.n295 C9_P_btm.n215 0.6255
R51001 C9_P_btm.n766 C9_P_btm.n765 0.6255
R51002 C9_P_btm.n769 C9_P_btm.n768 0.6255
R51003 C9_P_btm.n772 C9_P_btm.n771 0.6255
R51004 C9_P_btm.n775 C9_P_btm.n774 0.6255
R51005 C9_P_btm.n778 C9_P_btm.n777 0.6255
R51006 C9_P_btm.n781 C9_P_btm.n780 0.6255
R51007 C9_P_btm.n784 C9_P_btm.n783 0.6255
R51008 C9_P_btm.n787 C9_P_btm.n786 0.6255
R51009 C9_P_btm.n790 C9_P_btm.n789 0.6255
R51010 C9_P_btm.n793 C9_P_btm.n792 0.6255
R51011 C9_P_btm.n796 C9_P_btm.n795 0.6255
R51012 C9_P_btm.n799 C9_P_btm.n798 0.6255
R51013 C9_P_btm.n802 C9_P_btm.n801 0.6255
R51014 C9_P_btm.n805 C9_P_btm.n804 0.6255
R51015 C9_P_btm.n808 C9_P_btm.n807 0.6255
R51016 C9_P_btm.n811 C9_P_btm.n810 0.6255
R51017 C9_P_btm.n814 C9_P_btm.n813 0.6255
R51018 C9_P_btm.n817 C9_P_btm.n816 0.6255
R51019 C9_P_btm.n820 C9_P_btm.n819 0.6255
R51020 C9_P_btm.n823 C9_P_btm.n822 0.6255
R51021 C9_P_btm.n826 C9_P_btm.n825 0.6255
R51022 C9_P_btm.n829 C9_P_btm.n828 0.6255
R51023 C9_P_btm.n832 C9_P_btm.n831 0.6255
R51024 C9_P_btm.n835 C9_P_btm.n834 0.6255
R51025 C9_P_btm.n838 C9_P_btm.n837 0.6255
R51026 C9_P_btm.n841 C9_P_btm.n840 0.6255
R51027 C9_P_btm.n844 C9_P_btm.n843 0.6255
R51028 C9_P_btm.n847 C9_P_btm.n846 0.6255
R51029 C9_P_btm.n850 C9_P_btm.n849 0.6255
R51030 C9_P_btm.n853 C9_P_btm.n852 0.6255
R51031 C9_P_btm.n856 C9_P_btm.n855 0.6255
R51032 C9_P_btm.n859 C9_P_btm.n858 0.6255
R51033 C9_P_btm.n862 C9_P_btm.n861 0.6255
R51034 C9_P_btm.n865 C9_P_btm.n864 0.6255
R51035 C9_P_btm.n868 C9_P_btm.n867 0.6255
R51036 C9_P_btm.n871 C9_P_btm.n870 0.6255
R51037 C9_P_btm.n874 C9_P_btm.n873 0.6255
R51038 C9_P_btm.n877 C9_P_btm.n876 0.6255
R51039 C9_P_btm.n880 C9_P_btm.n879 0.6255
R51040 C9_P_btm.n1515 C9_P_btm.n1514 0.6255
R51041 C9_P_btm.n1518 C9_P_btm.n1517 0.6255
R51042 C9_P_btm.n1521 C9_P_btm.n1520 0.6255
R51043 C9_P_btm.n1524 C9_P_btm.n1523 0.6255
R51044 C9_P_btm.n1527 C9_P_btm.n1526 0.6255
R51045 C9_P_btm.n1530 C9_P_btm.n1529 0.6255
R51046 C9_P_btm.n1533 C9_P_btm.n1532 0.6255
R51047 C9_P_btm.n1536 C9_P_btm.n1535 0.6255
R51048 C9_P_btm.n1539 C9_P_btm.n1538 0.6255
R51049 C9_P_btm.n1542 C9_P_btm.n1541 0.6255
R51050 C9_P_btm.n1545 C9_P_btm.n1544 0.6255
R51051 C9_P_btm.n1548 C9_P_btm.n1547 0.6255
R51052 C9_P_btm.n1551 C9_P_btm.n1550 0.6255
R51053 C9_P_btm.n1554 C9_P_btm.n1553 0.6255
R51054 C9_P_btm.n1557 C9_P_btm.n1556 0.6255
R51055 C9_P_btm.n1560 C9_P_btm.n1559 0.6255
R51056 C9_P_btm.n1563 C9_P_btm.n1562 0.6255
R51057 C9_P_btm.n1566 C9_P_btm.n1565 0.6255
R51058 C9_P_btm.n1569 C9_P_btm.n1568 0.6255
R51059 C9_P_btm.n1572 C9_P_btm.n1571 0.6255
R51060 C9_P_btm.n1575 C9_P_btm.n1574 0.6255
R51061 C9_P_btm.n1578 C9_P_btm.n1577 0.6255
R51062 C9_P_btm.n1581 C9_P_btm.n1580 0.6255
R51063 C9_P_btm.n1584 C9_P_btm.n1583 0.6255
R51064 C9_P_btm.n1587 C9_P_btm.n1586 0.6255
R51065 C9_P_btm.n1590 C9_P_btm.n1589 0.6255
R51066 C9_P_btm.n1593 C9_P_btm.n1592 0.6255
R51067 C9_P_btm.n1596 C9_P_btm.n1595 0.6255
R51068 C9_P_btm.n1599 C9_P_btm.n1598 0.6255
R51069 C9_P_btm.n1602 C9_P_btm.n1601 0.6255
R51070 C9_P_btm.n1605 C9_P_btm.n1604 0.6255
R51071 C9_P_btm.n1608 C9_P_btm.n1607 0.6255
R51072 C9_P_btm.n1611 C9_P_btm.n1610 0.6255
R51073 C9_P_btm.n1614 C9_P_btm.n1613 0.6255
R51074 C9_P_btm.n1617 C9_P_btm.n1616 0.6255
R51075 C9_P_btm.n1620 C9_P_btm.n1619 0.6255
R51076 C9_P_btm.n1623 C9_P_btm.n1622 0.6255
R51077 C9_P_btm.n1626 C9_P_btm.n1625 0.6255
R51078 C9_P_btm.n1629 C9_P_btm.n1628 0.6255
R51079 C9_P_btm.n1391 C9_P_btm.n133 0.6255
R51080 C9_P_btm.n1394 C9_P_btm.n1393 0.6255
R51081 C9_P_btm.n1397 C9_P_btm.n1396 0.6255
R51082 C9_P_btm.n1400 C9_P_btm.n1399 0.6255
R51083 C9_P_btm.n1403 C9_P_btm.n1402 0.6255
R51084 C9_P_btm.n1406 C9_P_btm.n1405 0.6255
R51085 C9_P_btm.n1409 C9_P_btm.n1408 0.6255
R51086 C9_P_btm.n1412 C9_P_btm.n1411 0.6255
R51087 C9_P_btm.n1415 C9_P_btm.n1414 0.6255
R51088 C9_P_btm.n1418 C9_P_btm.n1417 0.6255
R51089 C9_P_btm.n1421 C9_P_btm.n1420 0.6255
R51090 C9_P_btm.n1424 C9_P_btm.n1423 0.6255
R51091 C9_P_btm.n1427 C9_P_btm.n1426 0.6255
R51092 C9_P_btm.n1430 C9_P_btm.n1429 0.6255
R51093 C9_P_btm.n1433 C9_P_btm.n1432 0.6255
R51094 C9_P_btm.n1436 C9_P_btm.n1435 0.6255
R51095 C9_P_btm.n1439 C9_P_btm.n1438 0.6255
R51096 C9_P_btm.n1442 C9_P_btm.n1441 0.6255
R51097 C9_P_btm.n1350 C9_P_btm.n1349 0.6255
R51098 C9_P_btm.n1353 C9_P_btm.n1352 0.6255
R51099 C9_P_btm.n1356 C9_P_btm.n1355 0.6255
R51100 C9_P_btm.n1359 C9_P_btm.n1358 0.6255
R51101 C9_P_btm.n1362 C9_P_btm.n1361 0.6255
R51102 C9_P_btm.n1365 C9_P_btm.n1364 0.6255
R51103 C9_P_btm.n1368 C9_P_btm.n1367 0.6255
R51104 C9_P_btm.n1371 C9_P_btm.n1370 0.6255
R51105 C9_P_btm.n1374 C9_P_btm.n1373 0.6255
R51106 C9_P_btm.n1377 C9_P_btm.n1376 0.6255
R51107 C9_P_btm.n1380 C9_P_btm.n1379 0.6255
R51108 C9_P_btm.n1383 C9_P_btm.n1382 0.6255
R51109 C9_P_btm.n1385 C9_P_btm.n128 0.6255
R51110 C9_P_btm.n1654 C9_P_btm.n1652 0.6255
R51111 C9_P_btm.n1650 C9_P_btm.n1649 0.6255
R51112 C9_P_btm.n1647 C9_P_btm.n1646 0.6255
R51113 C9_P_btm.n1644 C9_P_btm.n1643 0.6255
R51114 C9_P_btm.n1667 C9_P_btm.n1666 0.6255
R51115 C9_P_btm.n1664 C9_P_btm.n1663 0.6255
R51116 C9_P_btm.n1661 C9_P_btm.n1660 0.6255
R51117 C9_P_btm.n124 C9_P_btm.n122 0.6255
R51118 C9_P_btm.n120 C9_P_btm.n119 0.6255
R51119 C9_P_btm.n117 C9_P_btm.n109 0.6255
R51120 C9_P_btm.n1682 C9_P_btm.n1681 0.6255
R51121 C9_P_btm.n1685 C9_P_btm.n1684 0.6255
R51122 C9_P_btm.n1688 C9_P_btm.n1687 0.6255
R51123 C9_P_btm.n1698 C9_P_btm.n1697 0.6255
R51124 C9_P_btm.n1701 C9_P_btm.n1700 0.6255
R51125 C9_P_btm.n1704 C9_P_btm.n1703 0.6255
R51126 C9_P_btm.n94 C9_P_btm.n86 0.6255
R51127 C9_P_btm.n97 C9_P_btm.n96 0.6255
R51128 C9_P_btm.n101 C9_P_btm.n99 0.6255
R51129 C9_P_btm.n1725 C9_P_btm.n1724 0.6255
R51130 C9_P_btm.n1722 C9_P_btm.n1721 0.6255
R51131 C9_P_btm.n1719 C9_P_btm.n1718 0.6255
R51132 C9_P_btm.n1741 C9_P_btm.n1740 0.6255
R51133 C9_P_btm.n1738 C9_P_btm.n1737 0.6255
R51134 C9_P_btm.n1735 C9_P_btm.n1734 0.6255
R51135 C9_P_btm.n78 C9_P_btm.n76 0.6255
R51136 C9_P_btm.n74 C9_P_btm.n73 0.6255
R51137 C9_P_btm.n71 C9_P_btm.n63 0.6255
R51138 C9_P_btm.n1756 C9_P_btm.n1755 0.6255
R51139 C9_P_btm.n1759 C9_P_btm.n1758 0.6255
R51140 C9_P_btm.n1762 C9_P_btm.n1761 0.6255
R51141 C9_P_btm.n1772 C9_P_btm.n1771 0.6255
R51142 C9_P_btm.n1775 C9_P_btm.n1774 0.6255
R51143 C9_P_btm.n1778 C9_P_btm.n1777 0.6255
R51144 C9_P_btm.n48 C9_P_btm.n40 0.6255
R51145 C9_P_btm.n51 C9_P_btm.n50 0.6255
R51146 C9_P_btm.n55 C9_P_btm.n53 0.6255
R51147 C9_P_btm.n1799 C9_P_btm.n1798 0.6255
R51148 C9_P_btm.n1796 C9_P_btm.n1795 0.6255
R51149 C9_P_btm.n1793 C9_P_btm.n1792 0.6255
R51150 C9_P_btm.n1830 C9_P_btm.n1829 0.6255
R51151 C9_P_btm.n1827 C9_P_btm.n1826 0.6255
R51152 C9_P_btm.n1824 C9_P_btm.n1823 0.6255
R51153 C9_P_btm.n1814 C9_P_btm.n1813 0.6255
R51154 C9_P_btm.n1811 C9_P_btm.n1810 0.6255
R51155 C9_P_btm.n1808 C9_P_btm.n30 0.6255
R51156 C9_P_btm.n1845 C9_P_btm.n1844 0.6255
R51157 C9_P_btm.n1848 C9_P_btm.n1847 0.6255
R51158 C9_P_btm.n1852 C9_P_btm.n1850 0.6255
R51159 C9_P_btm.n1859 C9_P_btm.n1858 0.6255
R51160 C9_P_btm.n1862 C9_P_btm.n1861 0.6255
R51161 C9_P_btm.n1865 C9_P_btm.n1864 0.6255
R51162 C9_P_btm.n1875 C9_P_btm.n1874 0.6255
R51163 C9_P_btm.n1878 C9_P_btm.n1877 0.6255
R51164 C9_P_btm.n1881 C9_P_btm.n1880 0.6255
R51165 C9_P_btm.n1057 C9_P_btm.n1028 0.109875
R51166 C9_P_btm.n1059 C9_P_btm.n1028 0.109875
R51167 C9_P_btm.n1054 C9_P_btm.n1030 0.109875
R51168 C9_P_btm.n1056 C9_P_btm.n1030 0.109875
R51169 C9_P_btm.n1051 C9_P_btm.n1031 0.109875
R51170 C9_P_btm.n1053 C9_P_btm.n1031 0.109875
R51171 C9_P_btm.n1048 C9_P_btm.n1045 0.109875
R51172 C9_P_btm.n1050 C9_P_btm.n1045 0.109875
R51173 C9_P_btm.n1044 C9_P_btm.n1033 0.109875
R51174 C9_P_btm.n1044 C9_P_btm.n1043 0.109875
R51175 C9_P_btm.n1041 C9_P_btm.n1034 0.109875
R51176 C9_P_btm.n1039 C9_P_btm.n1034 0.109875
R51177 C9_P_btm.n1038 C9_P_btm.n1035 0.109875
R51178 C9_P_btm.n1036 C9_P_btm.n1035 0.109875
R51179 C9_P_btm.n1066 C9_P_btm.n1029 0.109875
R51180 C9_P_btm.n1066 C9_P_btm.n1065 0.109875
R51181 C9_P_btm.n1071 C9_P_btm.n1067 0.109875
R51182 C9_P_btm.n1069 C9_P_btm.n1067 0.109875
R51183 C9_P_btm.n1074 C9_P_btm.n1027 0.109875
R51184 C9_P_btm.n1072 C9_P_btm.n1027 0.109875
R51185 C9_P_btm.n1077 C9_P_btm.n1026 0.109875
R51186 C9_P_btm.n1075 C9_P_btm.n1026 0.109875
R51187 C9_P_btm.n1080 C9_P_btm.n1025 0.109875
R51188 C9_P_btm.n1078 C9_P_btm.n1025 0.109875
R51189 C9_P_btm.n1085 C9_P_btm.n1023 0.109875
R51190 C9_P_btm.n1087 C9_P_btm.n1023 0.109875
R51191 C9_P_btm.n1088 C9_P_btm.n1009 0.109875
R51192 C9_P_btm.n1090 C9_P_btm.n1009 0.109875
R51193 C9_P_btm.n1091 C9_P_btm.n1008 0.109875
R51194 C9_P_btm.n1093 C9_P_btm.n1008 0.109875
R51195 C9_P_btm.n1094 C9_P_btm.n1005 0.109875
R51196 C9_P_btm.n1096 C9_P_btm.n1005 0.109875
R51197 C9_P_btm.n1103 C9_P_btm.n1006 0.109875
R51198 C9_P_btm.n1103 C9_P_btm.n1102 0.109875
R51199 C9_P_btm.n1016 C9_P_btm.n1013 0.109875
R51200 C9_P_btm.n1014 C9_P_btm.n1013 0.109875
R51201 C9_P_btm.n1019 C9_P_btm.n1012 0.109875
R51202 C9_P_btm.n1017 C9_P_btm.n1012 0.109875
R51203 C9_P_btm.n1022 C9_P_btm.n1011 0.109875
R51204 C9_P_btm.n1022 C9_P_btm.n1021 0.109875
R51205 C9_P_btm.n1117 C9_P_btm.n1002 0.109875
R51206 C9_P_btm.n1115 C9_P_btm.n1002 0.109875
R51207 C9_P_btm.n1114 C9_P_btm.n1003 0.109875
R51208 C9_P_btm.n1112 C9_P_btm.n1003 0.109875
R51209 C9_P_btm.n1111 C9_P_btm.n1004 0.109875
R51210 C9_P_btm.n1109 C9_P_btm.n1004 0.109875
R51211 C9_P_btm.n1108 C9_P_btm.n1104 0.109875
R51212 C9_P_btm.n1106 C9_P_btm.n1104 0.109875
R51213 C9_P_btm.n1131 C9_P_btm.n982 0.109875
R51214 C9_P_btm.n1133 C9_P_btm.n982 0.109875
R51215 C9_P_btm.n1128 C9_P_btm.n985 0.109875
R51216 C9_P_btm.n1130 C9_P_btm.n985 0.109875
R51217 C9_P_btm.n1125 C9_P_btm.n986 0.109875
R51218 C9_P_btm.n1127 C9_P_btm.n986 0.109875
R51219 C9_P_btm.n1122 C9_P_btm.n1000 0.109875
R51220 C9_P_btm.n1124 C9_P_btm.n1000 0.109875
R51221 C9_P_btm.n999 C9_P_btm.n988 0.109875
R51222 C9_P_btm.n999 C9_P_btm.n998 0.109875
R51223 C9_P_btm.n996 C9_P_btm.n989 0.109875
R51224 C9_P_btm.n994 C9_P_btm.n989 0.109875
R51225 C9_P_btm.n993 C9_P_btm.n990 0.109875
R51226 C9_P_btm.n991 C9_P_btm.n990 0.109875
R51227 C9_P_btm.n1140 C9_P_btm.n983 0.109875
R51228 C9_P_btm.n1140 C9_P_btm.n1139 0.109875
R51229 C9_P_btm.n1145 C9_P_btm.n1141 0.109875
R51230 C9_P_btm.n1143 C9_P_btm.n1141 0.109875
R51231 C9_P_btm.n1148 C9_P_btm.n981 0.109875
R51232 C9_P_btm.n1146 C9_P_btm.n981 0.109875
R51233 C9_P_btm.n1151 C9_P_btm.n980 0.109875
R51234 C9_P_btm.n1149 C9_P_btm.n980 0.109875
R51235 C9_P_btm.n1154 C9_P_btm.n979 0.109875
R51236 C9_P_btm.n1152 C9_P_btm.n979 0.109875
R51237 C9_P_btm.n1159 C9_P_btm.n977 0.109875
R51238 C9_P_btm.n1161 C9_P_btm.n977 0.109875
R51239 C9_P_btm.n1162 C9_P_btm.n963 0.109875
R51240 C9_P_btm.n1164 C9_P_btm.n963 0.109875
R51241 C9_P_btm.n1165 C9_P_btm.n962 0.109875
R51242 C9_P_btm.n1167 C9_P_btm.n962 0.109875
R51243 C9_P_btm.n1168 C9_P_btm.n959 0.109875
R51244 C9_P_btm.n1170 C9_P_btm.n959 0.109875
R51245 C9_P_btm.n1177 C9_P_btm.n960 0.109875
R51246 C9_P_btm.n1177 C9_P_btm.n1176 0.109875
R51247 C9_P_btm.n970 C9_P_btm.n967 0.109875
R51248 C9_P_btm.n968 C9_P_btm.n967 0.109875
R51249 C9_P_btm.n973 C9_P_btm.n966 0.109875
R51250 C9_P_btm.n971 C9_P_btm.n966 0.109875
R51251 C9_P_btm.n976 C9_P_btm.n965 0.109875
R51252 C9_P_btm.n976 C9_P_btm.n975 0.109875
R51253 C9_P_btm.n1191 C9_P_btm.n956 0.109875
R51254 C9_P_btm.n1189 C9_P_btm.n956 0.109875
R51255 C9_P_btm.n1188 C9_P_btm.n957 0.109875
R51256 C9_P_btm.n1186 C9_P_btm.n957 0.109875
R51257 C9_P_btm.n1185 C9_P_btm.n958 0.109875
R51258 C9_P_btm.n1183 C9_P_btm.n958 0.109875
R51259 C9_P_btm.n1182 C9_P_btm.n1178 0.109875
R51260 C9_P_btm.n1180 C9_P_btm.n1178 0.109875
R51261 C9_P_btm.n1205 C9_P_btm.n936 0.109875
R51262 C9_P_btm.n1207 C9_P_btm.n936 0.109875
R51263 C9_P_btm.n1202 C9_P_btm.n939 0.109875
R51264 C9_P_btm.n1204 C9_P_btm.n939 0.109875
R51265 C9_P_btm.n1199 C9_P_btm.n940 0.109875
R51266 C9_P_btm.n1201 C9_P_btm.n940 0.109875
R51267 C9_P_btm.n1196 C9_P_btm.n954 0.109875
R51268 C9_P_btm.n1198 C9_P_btm.n954 0.109875
R51269 C9_P_btm.n953 C9_P_btm.n942 0.109875
R51270 C9_P_btm.n953 C9_P_btm.n952 0.109875
R51271 C9_P_btm.n950 C9_P_btm.n943 0.109875
R51272 C9_P_btm.n948 C9_P_btm.n943 0.109875
R51273 C9_P_btm.n947 C9_P_btm.n944 0.109875
R51274 C9_P_btm.n945 C9_P_btm.n944 0.109875
R51275 C9_P_btm.n1214 C9_P_btm.n937 0.109875
R51276 C9_P_btm.n1214 C9_P_btm.n1213 0.109875
R51277 C9_P_btm.n1219 C9_P_btm.n1215 0.109875
R51278 C9_P_btm.n1217 C9_P_btm.n1215 0.109875
R51279 C9_P_btm.n1222 C9_P_btm.n935 0.109875
R51280 C9_P_btm.n1220 C9_P_btm.n935 0.109875
R51281 C9_P_btm.n1225 C9_P_btm.n934 0.109875
R51282 C9_P_btm.n1223 C9_P_btm.n934 0.109875
R51283 C9_P_btm.n1228 C9_P_btm.n933 0.109875
R51284 C9_P_btm.n1226 C9_P_btm.n933 0.109875
R51285 C9_P_btm.n1233 C9_P_btm.n921 0.109875
R51286 C9_P_btm.n1235 C9_P_btm.n921 0.109875
R51287 C9_P_btm.n1236 C9_P_btm.n929 0.109875
R51288 C9_P_btm.n1238 C9_P_btm.n929 0.109875
R51289 C9_P_btm.n1239 C9_P_btm.n928 0.109875
R51290 C9_P_btm.n1241 C9_P_btm.n928 0.109875
R51291 C9_P_btm.n1242 C9_P_btm.n927 0.109875
R51292 C9_P_btm.n1244 C9_P_btm.n927 0.109875
R51293 C9_P_btm.n1251 C9_P_btm.n925 0.109875
R51294 C9_P_btm.n1249 C9_P_btm.n925 0.109875
R51295 C9_P_btm.n1254 C9_P_btm.n924 0.109875
R51296 C9_P_btm.n1252 C9_P_btm.n924 0.109875
R51297 C9_P_btm.n1257 C9_P_btm.n923 0.109875
R51298 C9_P_btm.n1255 C9_P_btm.n923 0.109875
R51299 C9_P_btm.n1260 C9_P_btm.n922 0.109875
R51300 C9_P_btm.n1260 C9_P_btm.n1259 0.109875
R51301 C9_P_btm.n1263 C9_P_btm.n1261 0.109875
R51302 C9_P_btm.n1265 C9_P_btm.n1261 0.109875
R51303 C9_P_btm.n1266 C9_P_btm.n920 0.109875
R51304 C9_P_btm.n1268 C9_P_btm.n920 0.109875
R51305 C9_P_btm.n1269 C9_P_btm.n919 0.109875
R51306 C9_P_btm.n1271 C9_P_btm.n919 0.109875
R51307 C9_P_btm.n1272 C9_P_btm.n918 0.109875
R51308 C9_P_btm.n1274 C9_P_btm.n918 0.109875
R51309 C9_P_btm.n1275 C9_P_btm.n917 0.109875
R51310 C9_P_btm.n1277 C9_P_btm.n917 0.109875
R51311 C9_P_btm.n1278 C9_P_btm.n916 0.109875
R51312 C9_P_btm.n1280 C9_P_btm.n916 0.109875
R51313 C9_P_btm.n1281 C9_P_btm.n915 0.109875
R51314 C9_P_btm.n1283 C9_P_btm.n915 0.109875
R51315 C9_P_btm.n1284 C9_P_btm.n914 0.109875
R51316 C9_P_btm.n1286 C9_P_btm.n914 0.109875
R51317 C9_P_btm.n1287 C9_P_btm.n913 0.109875
R51318 C9_P_btm.n1289 C9_P_btm.n913 0.109875
R51319 C9_P_btm.n1290 C9_P_btm.n912 0.109875
R51320 C9_P_btm.n1292 C9_P_btm.n912 0.109875
R51321 C9_P_btm.n1293 C9_P_btm.n911 0.109875
R51322 C9_P_btm.n1295 C9_P_btm.n911 0.109875
R51323 C9_P_btm.n1296 C9_P_btm.n910 0.109875
R51324 C9_P_btm.n1298 C9_P_btm.n910 0.109875
R51325 C9_P_btm.n1299 C9_P_btm.n909 0.109875
R51326 C9_P_btm.n1301 C9_P_btm.n909 0.109875
R51327 C9_P_btm.n1302 C9_P_btm.n908 0.109875
R51328 C9_P_btm.n1304 C9_P_btm.n908 0.109875
R51329 C9_P_btm.n1305 C9_P_btm.n907 0.109875
R51330 C9_P_btm.n1307 C9_P_btm.n907 0.109875
R51331 C9_P_btm.n1308 C9_P_btm.n906 0.109875
R51332 C9_P_btm.n1310 C9_P_btm.n906 0.109875
R51333 C9_P_btm.n1311 C9_P_btm.n905 0.109875
R51334 C9_P_btm.n1313 C9_P_btm.n905 0.109875
R51335 C9_P_btm.n1314 C9_P_btm.n904 0.109875
R51336 C9_P_btm.n1316 C9_P_btm.n904 0.109875
R51337 C9_P_btm.n1447 C9_P_btm.n1320 0.109875
R51338 C9_P_btm.n1445 C9_P_btm.n1320 0.109875
R51339 C9_P_btm.n1450 C9_P_btm.n1319 0.109875
R51340 C9_P_btm.n1448 C9_P_btm.n1319 0.109875
R51341 C9_P_btm.n1453 C9_P_btm.n1318 0.109875
R51342 C9_P_btm.n1451 C9_P_btm.n1318 0.109875
R51343 C9_P_btm.n1456 C9_P_btm.n903 0.109875
R51344 C9_P_btm.n1454 C9_P_btm.n903 0.109875
R51345 C9_P_btm.n1459 C9_P_btm.n902 0.109875
R51346 C9_P_btm.n1457 C9_P_btm.n902 0.109875
R51347 C9_P_btm.n1462 C9_P_btm.n901 0.109875
R51348 C9_P_btm.n1460 C9_P_btm.n901 0.109875
R51349 C9_P_btm.n1465 C9_P_btm.n900 0.109875
R51350 C9_P_btm.n1463 C9_P_btm.n900 0.109875
R51351 C9_P_btm.n1468 C9_P_btm.n899 0.109875
R51352 C9_P_btm.n1466 C9_P_btm.n899 0.109875
R51353 C9_P_btm.n1471 C9_P_btm.n898 0.109875
R51354 C9_P_btm.n1469 C9_P_btm.n898 0.109875
R51355 C9_P_btm.n1474 C9_P_btm.n897 0.109875
R51356 C9_P_btm.n1472 C9_P_btm.n897 0.109875
R51357 C9_P_btm.n1477 C9_P_btm.n896 0.109875
R51358 C9_P_btm.n1475 C9_P_btm.n896 0.109875
R51359 C9_P_btm.n1480 C9_P_btm.n895 0.109875
R51360 C9_P_btm.n1478 C9_P_btm.n895 0.109875
R51361 C9_P_btm.n1483 C9_P_btm.n894 0.109875
R51362 C9_P_btm.n1481 C9_P_btm.n894 0.109875
R51363 C9_P_btm.n1486 C9_P_btm.n893 0.109875
R51364 C9_P_btm.n1484 C9_P_btm.n893 0.109875
R51365 C9_P_btm.n1489 C9_P_btm.n892 0.109875
R51366 C9_P_btm.n1487 C9_P_btm.n892 0.109875
R51367 C9_P_btm.n1492 C9_P_btm.n891 0.109875
R51368 C9_P_btm.n1490 C9_P_btm.n891 0.109875
R51369 C9_P_btm.n1495 C9_P_btm.n890 0.109875
R51370 C9_P_btm.n1493 C9_P_btm.n890 0.109875
R51371 C9_P_btm.n1498 C9_P_btm.n889 0.109875
R51372 C9_P_btm.n1496 C9_P_btm.n889 0.109875
R51373 C9_P_btm.n1501 C9_P_btm.n888 0.109875
R51374 C9_P_btm.n1499 C9_P_btm.n888 0.109875
R51375 C9_P_btm.n1504 C9_P_btm.n887 0.109875
R51376 C9_P_btm.n1502 C9_P_btm.n887 0.109875
R51377 C9_P_btm.n1507 C9_P_btm.n886 0.109875
R51378 C9_P_btm.n1505 C9_P_btm.n886 0.109875
R51379 C9_P_btm.n494 C9_P_btm.n440 0.109875
R51380 C9_P_btm.n496 C9_P_btm.n440 0.109875
R51381 C9_P_btm.n491 C9_P_btm.n441 0.109875
R51382 C9_P_btm.n493 C9_P_btm.n441 0.109875
R51383 C9_P_btm.n488 C9_P_btm.n442 0.109875
R51384 C9_P_btm.n490 C9_P_btm.n442 0.109875
R51385 C9_P_btm.n485 C9_P_btm.n443 0.109875
R51386 C9_P_btm.n487 C9_P_btm.n443 0.109875
R51387 C9_P_btm.n482 C9_P_btm.n444 0.109875
R51388 C9_P_btm.n484 C9_P_btm.n444 0.109875
R51389 C9_P_btm.n479 C9_P_btm.n445 0.109875
R51390 C9_P_btm.n481 C9_P_btm.n445 0.109875
R51391 C9_P_btm.n476 C9_P_btm.n446 0.109875
R51392 C9_P_btm.n478 C9_P_btm.n446 0.109875
R51393 C9_P_btm.n473 C9_P_btm.n447 0.109875
R51394 C9_P_btm.n475 C9_P_btm.n447 0.109875
R51395 C9_P_btm.n470 C9_P_btm.n448 0.109875
R51396 C9_P_btm.n472 C9_P_btm.n448 0.109875
R51397 C9_P_btm.n467 C9_P_btm.n449 0.109875
R51398 C9_P_btm.n469 C9_P_btm.n449 0.109875
R51399 C9_P_btm.n464 C9_P_btm.n450 0.109875
R51400 C9_P_btm.n466 C9_P_btm.n450 0.109875
R51401 C9_P_btm.n461 C9_P_btm.n451 0.109875
R51402 C9_P_btm.n463 C9_P_btm.n451 0.109875
R51403 C9_P_btm.n458 C9_P_btm.n452 0.109875
R51404 C9_P_btm.n460 C9_P_btm.n452 0.109875
R51405 C9_P_btm.n455 C9_P_btm.n453 0.109875
R51406 C9_P_btm.n457 C9_P_btm.n453 0.109875
R51407 C9_P_btm.n630 C9_P_btm.n413 0.109875
R51408 C9_P_btm.n628 C9_P_btm.n413 0.109875
R51409 C9_P_btm.n627 C9_P_btm.n414 0.109875
R51410 C9_P_btm.n625 C9_P_btm.n414 0.109875
R51411 C9_P_btm.n624 C9_P_btm.n415 0.109875
R51412 C9_P_btm.n622 C9_P_btm.n415 0.109875
R51413 C9_P_btm.n621 C9_P_btm.n416 0.109875
R51414 C9_P_btm.n619 C9_P_btm.n416 0.109875
R51415 C9_P_btm.n618 C9_P_btm.n417 0.109875
R51416 C9_P_btm.n616 C9_P_btm.n417 0.109875
R51417 C9_P_btm.n615 C9_P_btm.n418 0.109875
R51418 C9_P_btm.n613 C9_P_btm.n418 0.109875
R51419 C9_P_btm.n612 C9_P_btm.n419 0.109875
R51420 C9_P_btm.n610 C9_P_btm.n419 0.109875
R51421 C9_P_btm.n609 C9_P_btm.n420 0.109875
R51422 C9_P_btm.n607 C9_P_btm.n420 0.109875
R51423 C9_P_btm.n606 C9_P_btm.n421 0.109875
R51424 C9_P_btm.n604 C9_P_btm.n421 0.109875
R51425 C9_P_btm.n603 C9_P_btm.n422 0.109875
R51426 C9_P_btm.n601 C9_P_btm.n422 0.109875
R51427 C9_P_btm.n600 C9_P_btm.n423 0.109875
R51428 C9_P_btm.n598 C9_P_btm.n423 0.109875
R51429 C9_P_btm.n597 C9_P_btm.n424 0.109875
R51430 C9_P_btm.n595 C9_P_btm.n424 0.109875
R51431 C9_P_btm.n594 C9_P_btm.n425 0.109875
R51432 C9_P_btm.n592 C9_P_btm.n425 0.109875
R51433 C9_P_btm.n591 C9_P_btm.n426 0.109875
R51434 C9_P_btm.n589 C9_P_btm.n426 0.109875
R51435 C9_P_btm.n588 C9_P_btm.n427 0.109875
R51436 C9_P_btm.n586 C9_P_btm.n427 0.109875
R51437 C9_P_btm.n585 C9_P_btm.n428 0.109875
R51438 C9_P_btm.n583 C9_P_btm.n428 0.109875
R51439 C9_P_btm.n582 C9_P_btm.n429 0.109875
R51440 C9_P_btm.n580 C9_P_btm.n429 0.109875
R51441 C9_P_btm.n579 C9_P_btm.n430 0.109875
R51442 C9_P_btm.n577 C9_P_btm.n430 0.109875
R51443 C9_P_btm.n576 C9_P_btm.n431 0.109875
R51444 C9_P_btm.n574 C9_P_btm.n431 0.109875
R51445 C9_P_btm.n573 C9_P_btm.n432 0.109875
R51446 C9_P_btm.n571 C9_P_btm.n432 0.109875
R51447 C9_P_btm.n570 C9_P_btm.n433 0.109875
R51448 C9_P_btm.n568 C9_P_btm.n433 0.109875
R51449 C9_P_btm.n567 C9_P_btm.n434 0.109875
R51450 C9_P_btm.n565 C9_P_btm.n434 0.109875
R51451 C9_P_btm.n564 C9_P_btm.n435 0.109875
R51452 C9_P_btm.n562 C9_P_btm.n435 0.109875
R51453 C9_P_btm.n561 C9_P_btm.n436 0.109875
R51454 C9_P_btm.n559 C9_P_btm.n436 0.109875
R51455 C9_P_btm.n558 C9_P_btm.n437 0.109875
R51456 C9_P_btm.n556 C9_P_btm.n437 0.109875
R51457 C9_P_btm.n555 C9_P_btm.n438 0.109875
R51458 C9_P_btm.n553 C9_P_btm.n438 0.109875
R51459 C9_P_btm.n552 C9_P_btm.n439 0.109875
R51460 C9_P_btm.n550 C9_P_btm.n439 0.109875
R51461 C9_P_btm.n549 C9_P_btm.n498 0.109875
R51462 C9_P_btm.n547 C9_P_btm.n498 0.109875
R51463 C9_P_btm.n546 C9_P_btm.n499 0.109875
R51464 C9_P_btm.n544 C9_P_btm.n499 0.109875
R51465 C9_P_btm.n543 C9_P_btm.n500 0.109875
R51466 C9_P_btm.n541 C9_P_btm.n500 0.109875
R51467 C9_P_btm.n540 C9_P_btm.n501 0.109875
R51468 C9_P_btm.n538 C9_P_btm.n501 0.109875
R51469 C9_P_btm.n537 C9_P_btm.n502 0.109875
R51470 C9_P_btm.n535 C9_P_btm.n502 0.109875
R51471 C9_P_btm.n534 C9_P_btm.n503 0.109875
R51472 C9_P_btm.n532 C9_P_btm.n503 0.109875
R51473 C9_P_btm.n531 C9_P_btm.n504 0.109875
R51474 C9_P_btm.n529 C9_P_btm.n504 0.109875
R51475 C9_P_btm.n528 C9_P_btm.n505 0.109875
R51476 C9_P_btm.n526 C9_P_btm.n505 0.109875
R51477 C9_P_btm.n525 C9_P_btm.n506 0.109875
R51478 C9_P_btm.n523 C9_P_btm.n506 0.109875
R51479 C9_P_btm.n522 C9_P_btm.n507 0.109875
R51480 C9_P_btm.n520 C9_P_btm.n507 0.109875
R51481 C9_P_btm.n519 C9_P_btm.n508 0.109875
R51482 C9_P_btm.n517 C9_P_btm.n508 0.109875
R51483 C9_P_btm.n516 C9_P_btm.n509 0.109875
R51484 C9_P_btm.n514 C9_P_btm.n509 0.109875
R51485 C9_P_btm.n513 C9_P_btm.n510 0.109875
R51486 C9_P_btm.n511 C9_P_btm.n510 0.109875
R51487 C9_P_btm.n751 C9_P_btm.n214 0.109875
R51488 C9_P_btm.n753 C9_P_btm.n214 0.109875
R51489 C9_P_btm.n748 C9_P_btm.n217 0.109875
R51490 C9_P_btm.n750 C9_P_btm.n217 0.109875
R51491 C9_P_btm.n745 C9_P_btm.n218 0.109875
R51492 C9_P_btm.n747 C9_P_btm.n218 0.109875
R51493 C9_P_btm.n742 C9_P_btm.n219 0.109875
R51494 C9_P_btm.n744 C9_P_btm.n219 0.109875
R51495 C9_P_btm.n739 C9_P_btm.n220 0.109875
R51496 C9_P_btm.n741 C9_P_btm.n220 0.109875
R51497 C9_P_btm.n736 C9_P_btm.n221 0.109875
R51498 C9_P_btm.n738 C9_P_btm.n221 0.109875
R51499 C9_P_btm.n733 C9_P_btm.n222 0.109875
R51500 C9_P_btm.n735 C9_P_btm.n222 0.109875
R51501 C9_P_btm.n730 C9_P_btm.n223 0.109875
R51502 C9_P_btm.n732 C9_P_btm.n223 0.109875
R51503 C9_P_btm.n727 C9_P_btm.n224 0.109875
R51504 C9_P_btm.n729 C9_P_btm.n224 0.109875
R51505 C9_P_btm.n724 C9_P_btm.n225 0.109875
R51506 C9_P_btm.n726 C9_P_btm.n225 0.109875
R51507 C9_P_btm.n721 C9_P_btm.n226 0.109875
R51508 C9_P_btm.n723 C9_P_btm.n226 0.109875
R51509 C9_P_btm.n718 C9_P_btm.n227 0.109875
R51510 C9_P_btm.n720 C9_P_btm.n227 0.109875
R51511 C9_P_btm.n715 C9_P_btm.n228 0.109875
R51512 C9_P_btm.n717 C9_P_btm.n228 0.109875
R51513 C9_P_btm.n712 C9_P_btm.n229 0.109875
R51514 C9_P_btm.n714 C9_P_btm.n229 0.109875
R51515 C9_P_btm.n709 C9_P_btm.n230 0.109875
R51516 C9_P_btm.n711 C9_P_btm.n230 0.109875
R51517 C9_P_btm.n706 C9_P_btm.n231 0.109875
R51518 C9_P_btm.n708 C9_P_btm.n231 0.109875
R51519 C9_P_btm.n703 C9_P_btm.n232 0.109875
R51520 C9_P_btm.n705 C9_P_btm.n232 0.109875
R51521 C9_P_btm.n700 C9_P_btm.n233 0.109875
R51522 C9_P_btm.n702 C9_P_btm.n233 0.109875
R51523 C9_P_btm.n697 C9_P_btm.n234 0.109875
R51524 C9_P_btm.n699 C9_P_btm.n234 0.109875
R51525 C9_P_btm.n694 C9_P_btm.n235 0.109875
R51526 C9_P_btm.n696 C9_P_btm.n235 0.109875
R51527 C9_P_btm.n691 C9_P_btm.n236 0.109875
R51528 C9_P_btm.n693 C9_P_btm.n236 0.109875
R51529 C9_P_btm.n688 C9_P_btm.n237 0.109875
R51530 C9_P_btm.n690 C9_P_btm.n237 0.109875
R51531 C9_P_btm.n685 C9_P_btm.n238 0.109875
R51532 C9_P_btm.n687 C9_P_btm.n238 0.109875
R51533 C9_P_btm.n682 C9_P_btm.n239 0.109875
R51534 C9_P_btm.n684 C9_P_btm.n239 0.109875
R51535 C9_P_btm.n679 C9_P_btm.n240 0.109875
R51536 C9_P_btm.n681 C9_P_btm.n240 0.109875
R51537 C9_P_btm.n676 C9_P_btm.n241 0.109875
R51538 C9_P_btm.n678 C9_P_btm.n241 0.109875
R51539 C9_P_btm.n673 C9_P_btm.n242 0.109875
R51540 C9_P_btm.n675 C9_P_btm.n242 0.109875
R51541 C9_P_btm.n670 C9_P_btm.n243 0.109875
R51542 C9_P_btm.n672 C9_P_btm.n243 0.109875
R51543 C9_P_btm.n667 C9_P_btm.n244 0.109875
R51544 C9_P_btm.n669 C9_P_btm.n244 0.109875
R51545 C9_P_btm.n664 C9_P_btm.n245 0.109875
R51546 C9_P_btm.n666 C9_P_btm.n245 0.109875
R51547 C9_P_btm.n661 C9_P_btm.n246 0.109875
R51548 C9_P_btm.n663 C9_P_btm.n246 0.109875
R51549 C9_P_btm.n658 C9_P_btm.n247 0.109875
R51550 C9_P_btm.n660 C9_P_btm.n247 0.109875
R51551 C9_P_btm.n655 C9_P_btm.n248 0.109875
R51552 C9_P_btm.n657 C9_P_btm.n248 0.109875
R51553 C9_P_btm.n652 C9_P_btm.n249 0.109875
R51554 C9_P_btm.n654 C9_P_btm.n249 0.109875
R51555 C9_P_btm.n649 C9_P_btm.n250 0.109875
R51556 C9_P_btm.n651 C9_P_btm.n250 0.109875
R51557 C9_P_btm.n646 C9_P_btm.n251 0.109875
R51558 C9_P_btm.n648 C9_P_btm.n251 0.109875
R51559 C9_P_btm.n643 C9_P_btm.n252 0.109875
R51560 C9_P_btm.n645 C9_P_btm.n252 0.109875
R51561 C9_P_btm.n640 C9_P_btm.n253 0.109875
R51562 C9_P_btm.n642 C9_P_btm.n253 0.109875
R51563 C9_P_btm.n637 C9_P_btm.n254 0.109875
R51564 C9_P_btm.n639 C9_P_btm.n254 0.109875
R51565 C9_P_btm.n634 C9_P_btm.n412 0.109875
R51566 C9_P_btm.n636 C9_P_btm.n412 0.109875
R51567 C9_P_btm.n411 C9_P_btm.n256 0.109875
R51568 C9_P_btm.n411 C9_P_btm.n410 0.109875
R51569 C9_P_btm.n408 C9_P_btm.n257 0.109875
R51570 C9_P_btm.n406 C9_P_btm.n257 0.109875
R51571 C9_P_btm.n405 C9_P_btm.n258 0.109875
R51572 C9_P_btm.n403 C9_P_btm.n258 0.109875
R51573 C9_P_btm.n402 C9_P_btm.n259 0.109875
R51574 C9_P_btm.n400 C9_P_btm.n259 0.109875
R51575 C9_P_btm.n399 C9_P_btm.n260 0.109875
R51576 C9_P_btm.n397 C9_P_btm.n260 0.109875
R51577 C9_P_btm.n396 C9_P_btm.n261 0.109875
R51578 C9_P_btm.n394 C9_P_btm.n261 0.109875
R51579 C9_P_btm.n393 C9_P_btm.n262 0.109875
R51580 C9_P_btm.n391 C9_P_btm.n262 0.109875
R51581 C9_P_btm.n390 C9_P_btm.n263 0.109875
R51582 C9_P_btm.n388 C9_P_btm.n263 0.109875
R51583 C9_P_btm.n387 C9_P_btm.n264 0.109875
R51584 C9_P_btm.n385 C9_P_btm.n264 0.109875
R51585 C9_P_btm.n384 C9_P_btm.n265 0.109875
R51586 C9_P_btm.n382 C9_P_btm.n265 0.109875
R51587 C9_P_btm.n381 C9_P_btm.n266 0.109875
R51588 C9_P_btm.n379 C9_P_btm.n266 0.109875
R51589 C9_P_btm.n378 C9_P_btm.n267 0.109875
R51590 C9_P_btm.n376 C9_P_btm.n267 0.109875
R51591 C9_P_btm.n375 C9_P_btm.n268 0.109875
R51592 C9_P_btm.n373 C9_P_btm.n268 0.109875
R51593 C9_P_btm.n372 C9_P_btm.n269 0.109875
R51594 C9_P_btm.n370 C9_P_btm.n269 0.109875
R51595 C9_P_btm.n369 C9_P_btm.n270 0.109875
R51596 C9_P_btm.n367 C9_P_btm.n270 0.109875
R51597 C9_P_btm.n366 C9_P_btm.n271 0.109875
R51598 C9_P_btm.n364 C9_P_btm.n271 0.109875
R51599 C9_P_btm.n363 C9_P_btm.n272 0.109875
R51600 C9_P_btm.n361 C9_P_btm.n272 0.109875
R51601 C9_P_btm.n360 C9_P_btm.n273 0.109875
R51602 C9_P_btm.n358 C9_P_btm.n273 0.109875
R51603 C9_P_btm.n357 C9_P_btm.n274 0.109875
R51604 C9_P_btm.n355 C9_P_btm.n274 0.109875
R51605 C9_P_btm.n354 C9_P_btm.n275 0.109875
R51606 C9_P_btm.n352 C9_P_btm.n275 0.109875
R51607 C9_P_btm.n351 C9_P_btm.n276 0.109875
R51608 C9_P_btm.n349 C9_P_btm.n276 0.109875
R51609 C9_P_btm.n348 C9_P_btm.n277 0.109875
R51610 C9_P_btm.n346 C9_P_btm.n277 0.109875
R51611 C9_P_btm.n345 C9_P_btm.n278 0.109875
R51612 C9_P_btm.n343 C9_P_btm.n278 0.109875
R51613 C9_P_btm.n342 C9_P_btm.n279 0.109875
R51614 C9_P_btm.n340 C9_P_btm.n279 0.109875
R51615 C9_P_btm.n339 C9_P_btm.n280 0.109875
R51616 C9_P_btm.n337 C9_P_btm.n280 0.109875
R51617 C9_P_btm.n336 C9_P_btm.n281 0.109875
R51618 C9_P_btm.n334 C9_P_btm.n281 0.109875
R51619 C9_P_btm.n333 C9_P_btm.n282 0.109875
R51620 C9_P_btm.n331 C9_P_btm.n282 0.109875
R51621 C9_P_btm.n330 C9_P_btm.n283 0.109875
R51622 C9_P_btm.n328 C9_P_btm.n283 0.109875
R51623 C9_P_btm.n327 C9_P_btm.n284 0.109875
R51624 C9_P_btm.n325 C9_P_btm.n284 0.109875
R51625 C9_P_btm.n324 C9_P_btm.n285 0.109875
R51626 C9_P_btm.n322 C9_P_btm.n285 0.109875
R51627 C9_P_btm.n321 C9_P_btm.n286 0.109875
R51628 C9_P_btm.n319 C9_P_btm.n286 0.109875
R51629 C9_P_btm.n318 C9_P_btm.n287 0.109875
R51630 C9_P_btm.n316 C9_P_btm.n287 0.109875
R51631 C9_P_btm.n315 C9_P_btm.n288 0.109875
R51632 C9_P_btm.n313 C9_P_btm.n288 0.109875
R51633 C9_P_btm.n312 C9_P_btm.n289 0.109875
R51634 C9_P_btm.n310 C9_P_btm.n289 0.109875
R51635 C9_P_btm.n309 C9_P_btm.n290 0.109875
R51636 C9_P_btm.n307 C9_P_btm.n290 0.109875
R51637 C9_P_btm.n306 C9_P_btm.n291 0.109875
R51638 C9_P_btm.n304 C9_P_btm.n291 0.109875
R51639 C9_P_btm.n303 C9_P_btm.n292 0.109875
R51640 C9_P_btm.n301 C9_P_btm.n292 0.109875
R51641 C9_P_btm.n300 C9_P_btm.n293 0.109875
R51642 C9_P_btm.n298 C9_P_btm.n293 0.109875
R51643 C9_P_btm.n297 C9_P_btm.n294 0.109875
R51644 C9_P_btm.n295 C9_P_btm.n294 0.109875
R51645 C9_P_btm.n760 C9_P_btm.n215 0.109875
R51646 C9_P_btm.n760 C9_P_btm.n759 0.109875
R51647 C9_P_btm.n765 C9_P_btm.n761 0.109875
R51648 C9_P_btm.n763 C9_P_btm.n761 0.109875
R51649 C9_P_btm.n768 C9_P_btm.n213 0.109875
R51650 C9_P_btm.n766 C9_P_btm.n213 0.109875
R51651 C9_P_btm.n771 C9_P_btm.n212 0.109875
R51652 C9_P_btm.n769 C9_P_btm.n212 0.109875
R51653 C9_P_btm.n774 C9_P_btm.n211 0.109875
R51654 C9_P_btm.n772 C9_P_btm.n211 0.109875
R51655 C9_P_btm.n777 C9_P_btm.n210 0.109875
R51656 C9_P_btm.n775 C9_P_btm.n210 0.109875
R51657 C9_P_btm.n780 C9_P_btm.n209 0.109875
R51658 C9_P_btm.n778 C9_P_btm.n209 0.109875
R51659 C9_P_btm.n783 C9_P_btm.n208 0.109875
R51660 C9_P_btm.n781 C9_P_btm.n208 0.109875
R51661 C9_P_btm.n786 C9_P_btm.n207 0.109875
R51662 C9_P_btm.n784 C9_P_btm.n207 0.109875
R51663 C9_P_btm.n789 C9_P_btm.n206 0.109875
R51664 C9_P_btm.n787 C9_P_btm.n206 0.109875
R51665 C9_P_btm.n792 C9_P_btm.n205 0.109875
R51666 C9_P_btm.n790 C9_P_btm.n205 0.109875
R51667 C9_P_btm.n795 C9_P_btm.n204 0.109875
R51668 C9_P_btm.n793 C9_P_btm.n204 0.109875
R51669 C9_P_btm.n798 C9_P_btm.n203 0.109875
R51670 C9_P_btm.n796 C9_P_btm.n203 0.109875
R51671 C9_P_btm.n801 C9_P_btm.n202 0.109875
R51672 C9_P_btm.n799 C9_P_btm.n202 0.109875
R51673 C9_P_btm.n804 C9_P_btm.n201 0.109875
R51674 C9_P_btm.n802 C9_P_btm.n201 0.109875
R51675 C9_P_btm.n807 C9_P_btm.n200 0.109875
R51676 C9_P_btm.n805 C9_P_btm.n200 0.109875
R51677 C9_P_btm.n810 C9_P_btm.n199 0.109875
R51678 C9_P_btm.n808 C9_P_btm.n199 0.109875
R51679 C9_P_btm.n813 C9_P_btm.n198 0.109875
R51680 C9_P_btm.n811 C9_P_btm.n198 0.109875
R51681 C9_P_btm.n816 C9_P_btm.n197 0.109875
R51682 C9_P_btm.n814 C9_P_btm.n197 0.109875
R51683 C9_P_btm.n819 C9_P_btm.n196 0.109875
R51684 C9_P_btm.n817 C9_P_btm.n196 0.109875
R51685 C9_P_btm.n822 C9_P_btm.n195 0.109875
R51686 C9_P_btm.n820 C9_P_btm.n195 0.109875
R51687 C9_P_btm.n825 C9_P_btm.n194 0.109875
R51688 C9_P_btm.n823 C9_P_btm.n194 0.109875
R51689 C9_P_btm.n828 C9_P_btm.n193 0.109875
R51690 C9_P_btm.n826 C9_P_btm.n193 0.109875
R51691 C9_P_btm.n831 C9_P_btm.n192 0.109875
R51692 C9_P_btm.n829 C9_P_btm.n192 0.109875
R51693 C9_P_btm.n834 C9_P_btm.n191 0.109875
R51694 C9_P_btm.n832 C9_P_btm.n191 0.109875
R51695 C9_P_btm.n837 C9_P_btm.n190 0.109875
R51696 C9_P_btm.n835 C9_P_btm.n190 0.109875
R51697 C9_P_btm.n840 C9_P_btm.n189 0.109875
R51698 C9_P_btm.n838 C9_P_btm.n189 0.109875
R51699 C9_P_btm.n843 C9_P_btm.n188 0.109875
R51700 C9_P_btm.n841 C9_P_btm.n188 0.109875
R51701 C9_P_btm.n846 C9_P_btm.n187 0.109875
R51702 C9_P_btm.n844 C9_P_btm.n187 0.109875
R51703 C9_P_btm.n849 C9_P_btm.n186 0.109875
R51704 C9_P_btm.n847 C9_P_btm.n186 0.109875
R51705 C9_P_btm.n852 C9_P_btm.n185 0.109875
R51706 C9_P_btm.n850 C9_P_btm.n185 0.109875
R51707 C9_P_btm.n855 C9_P_btm.n184 0.109875
R51708 C9_P_btm.n853 C9_P_btm.n184 0.109875
R51709 C9_P_btm.n858 C9_P_btm.n183 0.109875
R51710 C9_P_btm.n856 C9_P_btm.n183 0.109875
R51711 C9_P_btm.n861 C9_P_btm.n182 0.109875
R51712 C9_P_btm.n859 C9_P_btm.n182 0.109875
R51713 C9_P_btm.n864 C9_P_btm.n181 0.109875
R51714 C9_P_btm.n862 C9_P_btm.n181 0.109875
R51715 C9_P_btm.n867 C9_P_btm.n180 0.109875
R51716 C9_P_btm.n865 C9_P_btm.n180 0.109875
R51717 C9_P_btm.n870 C9_P_btm.n179 0.109875
R51718 C9_P_btm.n868 C9_P_btm.n179 0.109875
R51719 C9_P_btm.n873 C9_P_btm.n178 0.109875
R51720 C9_P_btm.n871 C9_P_btm.n178 0.109875
R51721 C9_P_btm.n876 C9_P_btm.n177 0.109875
R51722 C9_P_btm.n874 C9_P_btm.n177 0.109875
R51723 C9_P_btm.n879 C9_P_btm.n176 0.109875
R51724 C9_P_btm.n877 C9_P_btm.n176 0.109875
R51725 C9_P_btm.n882 C9_P_btm.n175 0.109875
R51726 C9_P_btm.n880 C9_P_btm.n175 0.109875
R51727 C9_P_btm.n1512 C9_P_btm.n173 0.109875
R51728 C9_P_btm.n1514 C9_P_btm.n173 0.109875
R51729 C9_P_btm.n1515 C9_P_btm.n172 0.109875
R51730 C9_P_btm.n1517 C9_P_btm.n172 0.109875
R51731 C9_P_btm.n1518 C9_P_btm.n171 0.109875
R51732 C9_P_btm.n1520 C9_P_btm.n171 0.109875
R51733 C9_P_btm.n1521 C9_P_btm.n170 0.109875
R51734 C9_P_btm.n1523 C9_P_btm.n170 0.109875
R51735 C9_P_btm.n1524 C9_P_btm.n169 0.109875
R51736 C9_P_btm.n1526 C9_P_btm.n169 0.109875
R51737 C9_P_btm.n1527 C9_P_btm.n168 0.109875
R51738 C9_P_btm.n1529 C9_P_btm.n168 0.109875
R51739 C9_P_btm.n1530 C9_P_btm.n167 0.109875
R51740 C9_P_btm.n1532 C9_P_btm.n167 0.109875
R51741 C9_P_btm.n1533 C9_P_btm.n166 0.109875
R51742 C9_P_btm.n1535 C9_P_btm.n166 0.109875
R51743 C9_P_btm.n1536 C9_P_btm.n165 0.109875
R51744 C9_P_btm.n1538 C9_P_btm.n165 0.109875
R51745 C9_P_btm.n1539 C9_P_btm.n164 0.109875
R51746 C9_P_btm.n1541 C9_P_btm.n164 0.109875
R51747 C9_P_btm.n1542 C9_P_btm.n163 0.109875
R51748 C9_P_btm.n1544 C9_P_btm.n163 0.109875
R51749 C9_P_btm.n1545 C9_P_btm.n162 0.109875
R51750 C9_P_btm.n1547 C9_P_btm.n162 0.109875
R51751 C9_P_btm.n1548 C9_P_btm.n161 0.109875
R51752 C9_P_btm.n1550 C9_P_btm.n161 0.109875
R51753 C9_P_btm.n1551 C9_P_btm.n160 0.109875
R51754 C9_P_btm.n1553 C9_P_btm.n160 0.109875
R51755 C9_P_btm.n1554 C9_P_btm.n159 0.109875
R51756 C9_P_btm.n1556 C9_P_btm.n159 0.109875
R51757 C9_P_btm.n1557 C9_P_btm.n158 0.109875
R51758 C9_P_btm.n1559 C9_P_btm.n158 0.109875
R51759 C9_P_btm.n1560 C9_P_btm.n157 0.109875
R51760 C9_P_btm.n1562 C9_P_btm.n157 0.109875
R51761 C9_P_btm.n1563 C9_P_btm.n156 0.109875
R51762 C9_P_btm.n1565 C9_P_btm.n156 0.109875
R51763 C9_P_btm.n1566 C9_P_btm.n155 0.109875
R51764 C9_P_btm.n1568 C9_P_btm.n155 0.109875
R51765 C9_P_btm.n1569 C9_P_btm.n154 0.109875
R51766 C9_P_btm.n1571 C9_P_btm.n154 0.109875
R51767 C9_P_btm.n1572 C9_P_btm.n153 0.109875
R51768 C9_P_btm.n1574 C9_P_btm.n153 0.109875
R51769 C9_P_btm.n1575 C9_P_btm.n152 0.109875
R51770 C9_P_btm.n1577 C9_P_btm.n152 0.109875
R51771 C9_P_btm.n1578 C9_P_btm.n151 0.109875
R51772 C9_P_btm.n1580 C9_P_btm.n151 0.109875
R51773 C9_P_btm.n1581 C9_P_btm.n150 0.109875
R51774 C9_P_btm.n1583 C9_P_btm.n150 0.109875
R51775 C9_P_btm.n1584 C9_P_btm.n149 0.109875
R51776 C9_P_btm.n1586 C9_P_btm.n149 0.109875
R51777 C9_P_btm.n1587 C9_P_btm.n148 0.109875
R51778 C9_P_btm.n1589 C9_P_btm.n148 0.109875
R51779 C9_P_btm.n1590 C9_P_btm.n147 0.109875
R51780 C9_P_btm.n1592 C9_P_btm.n147 0.109875
R51781 C9_P_btm.n1593 C9_P_btm.n146 0.109875
R51782 C9_P_btm.n1595 C9_P_btm.n146 0.109875
R51783 C9_P_btm.n1596 C9_P_btm.n145 0.109875
R51784 C9_P_btm.n1598 C9_P_btm.n145 0.109875
R51785 C9_P_btm.n1599 C9_P_btm.n144 0.109875
R51786 C9_P_btm.n1601 C9_P_btm.n144 0.109875
R51787 C9_P_btm.n1602 C9_P_btm.n143 0.109875
R51788 C9_P_btm.n1604 C9_P_btm.n143 0.109875
R51789 C9_P_btm.n1605 C9_P_btm.n142 0.109875
R51790 C9_P_btm.n1607 C9_P_btm.n142 0.109875
R51791 C9_P_btm.n1608 C9_P_btm.n141 0.109875
R51792 C9_P_btm.n1610 C9_P_btm.n141 0.109875
R51793 C9_P_btm.n1611 C9_P_btm.n140 0.109875
R51794 C9_P_btm.n1613 C9_P_btm.n140 0.109875
R51795 C9_P_btm.n1614 C9_P_btm.n139 0.109875
R51796 C9_P_btm.n1616 C9_P_btm.n139 0.109875
R51797 C9_P_btm.n1617 C9_P_btm.n138 0.109875
R51798 C9_P_btm.n1619 C9_P_btm.n138 0.109875
R51799 C9_P_btm.n1620 C9_P_btm.n137 0.109875
R51800 C9_P_btm.n1622 C9_P_btm.n137 0.109875
R51801 C9_P_btm.n1623 C9_P_btm.n136 0.109875
R51802 C9_P_btm.n1625 C9_P_btm.n136 0.109875
R51803 C9_P_btm.n1626 C9_P_btm.n135 0.109875
R51804 C9_P_btm.n1628 C9_P_btm.n135 0.109875
R51805 C9_P_btm.n1629 C9_P_btm.n132 0.109875
R51806 C9_P_btm.n1631 C9_P_btm.n132 0.109875
R51807 C9_P_btm.n1638 C9_P_btm.n133 0.109875
R51808 C9_P_btm.n1638 C9_P_btm.n1637 0.109875
R51809 C9_P_btm.n1393 C9_P_btm.n1390 0.109875
R51810 C9_P_btm.n1391 C9_P_btm.n1390 0.109875
R51811 C9_P_btm.n1396 C9_P_btm.n1389 0.109875
R51812 C9_P_btm.n1394 C9_P_btm.n1389 0.109875
R51813 C9_P_btm.n1399 C9_P_btm.n1388 0.109875
R51814 C9_P_btm.n1397 C9_P_btm.n1388 0.109875
R51815 C9_P_btm.n1402 C9_P_btm.n127 0.109875
R51816 C9_P_btm.n1400 C9_P_btm.n127 0.109875
R51817 C9_P_btm.n1405 C9_P_btm.n1387 0.109875
R51818 C9_P_btm.n1403 C9_P_btm.n1387 0.109875
R51819 C9_P_btm.n1408 C9_P_btm.n1333 0.109875
R51820 C9_P_btm.n1406 C9_P_btm.n1333 0.109875
R51821 C9_P_btm.n1411 C9_P_btm.n1332 0.109875
R51822 C9_P_btm.n1409 C9_P_btm.n1332 0.109875
R51823 C9_P_btm.n1414 C9_P_btm.n1331 0.109875
R51824 C9_P_btm.n1412 C9_P_btm.n1331 0.109875
R51825 C9_P_btm.n1417 C9_P_btm.n1330 0.109875
R51826 C9_P_btm.n1415 C9_P_btm.n1330 0.109875
R51827 C9_P_btm.n1420 C9_P_btm.n1329 0.109875
R51828 C9_P_btm.n1418 C9_P_btm.n1329 0.109875
R51829 C9_P_btm.n1423 C9_P_btm.n1328 0.109875
R51830 C9_P_btm.n1421 C9_P_btm.n1328 0.109875
R51831 C9_P_btm.n1426 C9_P_btm.n1327 0.109875
R51832 C9_P_btm.n1424 C9_P_btm.n1327 0.109875
R51833 C9_P_btm.n1429 C9_P_btm.n1326 0.109875
R51834 C9_P_btm.n1427 C9_P_btm.n1326 0.109875
R51835 C9_P_btm.n1432 C9_P_btm.n1325 0.109875
R51836 C9_P_btm.n1430 C9_P_btm.n1325 0.109875
R51837 C9_P_btm.n1435 C9_P_btm.n1324 0.109875
R51838 C9_P_btm.n1433 C9_P_btm.n1324 0.109875
R51839 C9_P_btm.n1438 C9_P_btm.n1323 0.109875
R51840 C9_P_btm.n1436 C9_P_btm.n1323 0.109875
R51841 C9_P_btm.n1441 C9_P_btm.n1322 0.109875
R51842 C9_P_btm.n1439 C9_P_btm.n1322 0.109875
R51843 C9_P_btm.n1444 C9_P_btm.n1321 0.109875
R51844 C9_P_btm.n1442 C9_P_btm.n1321 0.109875
R51845 C9_P_btm.n1347 C9_P_btm.n1345 0.109875
R51846 C9_P_btm.n1349 C9_P_btm.n1345 0.109875
R51847 C9_P_btm.n1350 C9_P_btm.n1344 0.109875
R51848 C9_P_btm.n1352 C9_P_btm.n1344 0.109875
R51849 C9_P_btm.n1353 C9_P_btm.n1343 0.109875
R51850 C9_P_btm.n1355 C9_P_btm.n1343 0.109875
R51851 C9_P_btm.n1356 C9_P_btm.n1342 0.109875
R51852 C9_P_btm.n1358 C9_P_btm.n1342 0.109875
R51853 C9_P_btm.n1359 C9_P_btm.n1341 0.109875
R51854 C9_P_btm.n1361 C9_P_btm.n1341 0.109875
R51855 C9_P_btm.n1362 C9_P_btm.n1340 0.109875
R51856 C9_P_btm.n1364 C9_P_btm.n1340 0.109875
R51857 C9_P_btm.n1365 C9_P_btm.n1339 0.109875
R51858 C9_P_btm.n1367 C9_P_btm.n1339 0.109875
R51859 C9_P_btm.n1368 C9_P_btm.n1338 0.109875
R51860 C9_P_btm.n1370 C9_P_btm.n1338 0.109875
R51861 C9_P_btm.n1371 C9_P_btm.n1337 0.109875
R51862 C9_P_btm.n1373 C9_P_btm.n1337 0.109875
R51863 C9_P_btm.n1374 C9_P_btm.n1336 0.109875
R51864 C9_P_btm.n1376 C9_P_btm.n1336 0.109875
R51865 C9_P_btm.n1377 C9_P_btm.n1335 0.109875
R51866 C9_P_btm.n1379 C9_P_btm.n1335 0.109875
R51867 C9_P_btm.n1380 C9_P_btm.n1334 0.109875
R51868 C9_P_btm.n1382 C9_P_btm.n1334 0.109875
R51869 C9_P_btm.n1386 C9_P_btm.n1383 0.109875
R51870 C9_P_btm.n1386 C9_P_btm.n1385 0.109875
R51871 C9_P_btm.n1655 C9_P_btm.n128 0.109875
R51872 C9_P_btm.n1655 C9_P_btm.n1654 0.109875
R51873 C9_P_btm.n1652 C9_P_btm.n129 0.109875
R51874 C9_P_btm.n1650 C9_P_btm.n129 0.109875
R51875 C9_P_btm.n1649 C9_P_btm.n130 0.109875
R51876 C9_P_btm.n1647 C9_P_btm.n130 0.109875
R51877 C9_P_btm.n1646 C9_P_btm.n131 0.109875
R51878 C9_P_btm.n1644 C9_P_btm.n131 0.109875
R51879 C9_P_btm.n1643 C9_P_btm.n1639 0.109875
R51880 C9_P_btm.n1641 C9_P_btm.n1639 0.109875
R51881 C9_P_btm.n1667 C9_P_btm.n108 0.109875
R51882 C9_P_btm.n1669 C9_P_btm.n108 0.109875
R51883 C9_P_btm.n1664 C9_P_btm.n111 0.109875
R51884 C9_P_btm.n1666 C9_P_btm.n111 0.109875
R51885 C9_P_btm.n1661 C9_P_btm.n112 0.109875
R51886 C9_P_btm.n1663 C9_P_btm.n112 0.109875
R51887 C9_P_btm.n1658 C9_P_btm.n126 0.109875
R51888 C9_P_btm.n1660 C9_P_btm.n126 0.109875
R51889 C9_P_btm.n125 C9_P_btm.n114 0.109875
R51890 C9_P_btm.n125 C9_P_btm.n124 0.109875
R51891 C9_P_btm.n122 C9_P_btm.n115 0.109875
R51892 C9_P_btm.n120 C9_P_btm.n115 0.109875
R51893 C9_P_btm.n119 C9_P_btm.n116 0.109875
R51894 C9_P_btm.n117 C9_P_btm.n116 0.109875
R51895 C9_P_btm.n1676 C9_P_btm.n109 0.109875
R51896 C9_P_btm.n1676 C9_P_btm.n1675 0.109875
R51897 C9_P_btm.n1681 C9_P_btm.n1677 0.109875
R51898 C9_P_btm.n1679 C9_P_btm.n1677 0.109875
R51899 C9_P_btm.n1684 C9_P_btm.n107 0.109875
R51900 C9_P_btm.n1682 C9_P_btm.n107 0.109875
R51901 C9_P_btm.n1687 C9_P_btm.n106 0.109875
R51902 C9_P_btm.n1685 C9_P_btm.n106 0.109875
R51903 C9_P_btm.n1690 C9_P_btm.n105 0.109875
R51904 C9_P_btm.n1688 C9_P_btm.n105 0.109875
R51905 C9_P_btm.n1695 C9_P_btm.n103 0.109875
R51906 C9_P_btm.n1697 C9_P_btm.n103 0.109875
R51907 C9_P_btm.n1698 C9_P_btm.n89 0.109875
R51908 C9_P_btm.n1700 C9_P_btm.n89 0.109875
R51909 C9_P_btm.n1701 C9_P_btm.n88 0.109875
R51910 C9_P_btm.n1703 C9_P_btm.n88 0.109875
R51911 C9_P_btm.n1704 C9_P_btm.n85 0.109875
R51912 C9_P_btm.n1706 C9_P_btm.n85 0.109875
R51913 C9_P_btm.n1713 C9_P_btm.n86 0.109875
R51914 C9_P_btm.n1713 C9_P_btm.n1712 0.109875
R51915 C9_P_btm.n96 C9_P_btm.n93 0.109875
R51916 C9_P_btm.n94 C9_P_btm.n93 0.109875
R51917 C9_P_btm.n99 C9_P_btm.n92 0.109875
R51918 C9_P_btm.n97 C9_P_btm.n92 0.109875
R51919 C9_P_btm.n102 C9_P_btm.n91 0.109875
R51920 C9_P_btm.n102 C9_P_btm.n101 0.109875
R51921 C9_P_btm.n1727 C9_P_btm.n82 0.109875
R51922 C9_P_btm.n1725 C9_P_btm.n82 0.109875
R51923 C9_P_btm.n1724 C9_P_btm.n83 0.109875
R51924 C9_P_btm.n1722 C9_P_btm.n83 0.109875
R51925 C9_P_btm.n1721 C9_P_btm.n84 0.109875
R51926 C9_P_btm.n1719 C9_P_btm.n84 0.109875
R51927 C9_P_btm.n1718 C9_P_btm.n1714 0.109875
R51928 C9_P_btm.n1716 C9_P_btm.n1714 0.109875
R51929 C9_P_btm.n1741 C9_P_btm.n62 0.109875
R51930 C9_P_btm.n1743 C9_P_btm.n62 0.109875
R51931 C9_P_btm.n1738 C9_P_btm.n65 0.109875
R51932 C9_P_btm.n1740 C9_P_btm.n65 0.109875
R51933 C9_P_btm.n1735 C9_P_btm.n66 0.109875
R51934 C9_P_btm.n1737 C9_P_btm.n66 0.109875
R51935 C9_P_btm.n1732 C9_P_btm.n80 0.109875
R51936 C9_P_btm.n1734 C9_P_btm.n80 0.109875
R51937 C9_P_btm.n79 C9_P_btm.n68 0.109875
R51938 C9_P_btm.n79 C9_P_btm.n78 0.109875
R51939 C9_P_btm.n76 C9_P_btm.n69 0.109875
R51940 C9_P_btm.n74 C9_P_btm.n69 0.109875
R51941 C9_P_btm.n73 C9_P_btm.n70 0.109875
R51942 C9_P_btm.n71 C9_P_btm.n70 0.109875
R51943 C9_P_btm.n1750 C9_P_btm.n63 0.109875
R51944 C9_P_btm.n1750 C9_P_btm.n1749 0.109875
R51945 C9_P_btm.n1755 C9_P_btm.n1751 0.109875
R51946 C9_P_btm.n1753 C9_P_btm.n1751 0.109875
R51947 C9_P_btm.n1758 C9_P_btm.n61 0.109875
R51948 C9_P_btm.n1756 C9_P_btm.n61 0.109875
R51949 C9_P_btm.n1761 C9_P_btm.n60 0.109875
R51950 C9_P_btm.n1759 C9_P_btm.n60 0.109875
R51951 C9_P_btm.n1764 C9_P_btm.n59 0.109875
R51952 C9_P_btm.n1762 C9_P_btm.n59 0.109875
R51953 C9_P_btm.n1769 C9_P_btm.n57 0.109875
R51954 C9_P_btm.n1771 C9_P_btm.n57 0.109875
R51955 C9_P_btm.n1772 C9_P_btm.n43 0.109875
R51956 C9_P_btm.n1774 C9_P_btm.n43 0.109875
R51957 C9_P_btm.n1775 C9_P_btm.n42 0.109875
R51958 C9_P_btm.n1777 C9_P_btm.n42 0.109875
R51959 C9_P_btm.n1778 C9_P_btm.n39 0.109875
R51960 C9_P_btm.n1780 C9_P_btm.n39 0.109875
R51961 C9_P_btm.n1787 C9_P_btm.n40 0.109875
R51962 C9_P_btm.n1787 C9_P_btm.n1786 0.109875
R51963 C9_P_btm.n50 C9_P_btm.n47 0.109875
R51964 C9_P_btm.n48 C9_P_btm.n47 0.109875
R51965 C9_P_btm.n53 C9_P_btm.n46 0.109875
R51966 C9_P_btm.n51 C9_P_btm.n46 0.109875
R51967 C9_P_btm.n56 C9_P_btm.n45 0.109875
R51968 C9_P_btm.n56 C9_P_btm.n55 0.109875
R51969 C9_P_btm.n1801 C9_P_btm.n36 0.109875
R51970 C9_P_btm.n1799 C9_P_btm.n36 0.109875
R51971 C9_P_btm.n1798 C9_P_btm.n37 0.109875
R51972 C9_P_btm.n1796 C9_P_btm.n37 0.109875
R51973 C9_P_btm.n1795 C9_P_btm.n38 0.109875
R51974 C9_P_btm.n1793 C9_P_btm.n38 0.109875
R51975 C9_P_btm.n1792 C9_P_btm.n1788 0.109875
R51976 C9_P_btm.n1790 C9_P_btm.n1788 0.109875
R51977 C9_P_btm.n1830 C9_P_btm.n29 0.109875
R51978 C9_P_btm.n1832 C9_P_btm.n29 0.109875
R51979 C9_P_btm.n1827 C9_P_btm.n32 0.109875
R51980 C9_P_btm.n1829 C9_P_btm.n32 0.109875
R51981 C9_P_btm.n1824 C9_P_btm.n33 0.109875
R51982 C9_P_btm.n1826 C9_P_btm.n33 0.109875
R51983 C9_P_btm.n1821 C9_P_btm.n34 0.109875
R51984 C9_P_btm.n1823 C9_P_btm.n34 0.109875
R51985 C9_P_btm.n1816 C9_P_btm.n25 0.109875
R51986 C9_P_btm.n1814 C9_P_btm.n25 0.109875
R51987 C9_P_btm.n1813 C9_P_btm.n1806 0.109875
R51988 C9_P_btm.n1811 C9_P_btm.n1806 0.109875
R51989 C9_P_btm.n1810 C9_P_btm.n1807 0.109875
R51990 C9_P_btm.n1808 C9_P_btm.n1807 0.109875
R51991 C9_P_btm.n1839 C9_P_btm.n30 0.109875
R51992 C9_P_btm.n1839 C9_P_btm.n1838 0.109875
R51993 C9_P_btm.n1844 C9_P_btm.n1840 0.109875
R51994 C9_P_btm.n1842 C9_P_btm.n1840 0.109875
R51995 C9_P_btm.n1847 C9_P_btm.n28 0.109875
R51996 C9_P_btm.n1845 C9_P_btm.n28 0.109875
R51997 C9_P_btm.n1850 C9_P_btm.n27 0.109875
R51998 C9_P_btm.n1848 C9_P_btm.n27 0.109875
R51999 C9_P_btm.n1853 C9_P_btm.n26 0.109875
R52000 C9_P_btm.n1853 C9_P_btm.n1852 0.109875
R52001 C9_P_btm.n1856 C9_P_btm.n1854 0.109875
R52002 C9_P_btm.n1858 C9_P_btm.n1854 0.109875
R52003 C9_P_btm.n1859 C9_P_btm.n24 0.109875
R52004 C9_P_btm.n1861 C9_P_btm.n24 0.109875
R52005 C9_P_btm.n1862 C9_P_btm.n23 0.109875
R52006 C9_P_btm.n1864 C9_P_btm.n23 0.109875
R52007 C9_P_btm.n1865 C9_P_btm.n22 0.109875
R52008 C9_P_btm.n1867 C9_P_btm.n22 0.109875
R52009 C9_P_btm.n1874 C9_P_btm.n20 0.109875
R52010 C9_P_btm.n1872 C9_P_btm.n20 0.109875
R52011 C9_P_btm.n1877 C9_P_btm.n19 0.109875
R52012 C9_P_btm.n1875 C9_P_btm.n19 0.109875
R52013 C9_P_btm.n1880 C9_P_btm.n18 0.109875
R52014 C9_P_btm.n1878 C9_P_btm.n18 0.109875
R52015 C9_P_btm.n1883 C9_P_btm.n17 0.109875
R52016 C9_P_btm.n1881 C9_P_btm.n17 0.109875
R52017 C9_P_btm.n1061 C9_P_btm.n1060 0.0556875
R52018 C9_P_btm.n1047 C9_P_btm.n1046 0.0556875
R52019 C9_P_btm.n1032 C9_P_btm.n1024 0.0556875
R52020 C9_P_btm.n1063 C9_P_btm.n1062 0.0556875
R52021 C9_P_btm.n1068 C9_P_btm.n1007 0.0556875
R52022 C9_P_btm.n1082 C9_P_btm.n1081 0.0556875
R52023 C9_P_btm.n1084 C9_P_btm.n1083 0.0556875
R52024 C9_P_btm.n1098 C9_P_btm.n1097 0.0556875
R52025 C9_P_btm.n1100 C9_P_btm.n1099 0.0556875
R52026 C9_P_btm.n1010 C9_P_btm.n1001 0.0556875
R52027 C9_P_btm.n1119 C9_P_btm.n1118 0.0556875
R52028 C9_P_btm.n1105 C9_P_btm.n984 0.0556875
R52029 C9_P_btm.n1135 C9_P_btm.n1134 0.0556875
R52030 C9_P_btm.n1121 C9_P_btm.n1120 0.0556875
R52031 C9_P_btm.n987 C9_P_btm.n978 0.0556875
R52032 C9_P_btm.n1137 C9_P_btm.n1136 0.0556875
R52033 C9_P_btm.n1142 C9_P_btm.n961 0.0556875
R52034 C9_P_btm.n1156 C9_P_btm.n1155 0.0556875
R52035 C9_P_btm.n1158 C9_P_btm.n1157 0.0556875
R52036 C9_P_btm.n1172 C9_P_btm.n1171 0.0556875
R52037 C9_P_btm.n1174 C9_P_btm.n1173 0.0556875
R52038 C9_P_btm.n964 C9_P_btm.n955 0.0556875
R52039 C9_P_btm.n1193 C9_P_btm.n1192 0.0556875
R52040 C9_P_btm.n1179 C9_P_btm.n938 0.0556875
R52041 C9_P_btm.n1209 C9_P_btm.n1208 0.0556875
R52042 C9_P_btm.n1195 C9_P_btm.n1194 0.0556875
R52043 C9_P_btm.n941 C9_P_btm.n932 0.0556875
R52044 C9_P_btm.n1211 C9_P_btm.n1210 0.0556875
R52045 C9_P_btm.n1216 C9_P_btm.n926 0.0556875
R52046 C9_P_btm.n1230 C9_P_btm.n1229 0.0556875
R52047 C9_P_btm.n1232 C9_P_btm.n1231 0.0556875
R52048 C9_P_btm.n1246 C9_P_btm.n1245 0.0556875
R52049 C9_P_btm.n1248 C9_P_btm.n1247 0.0556875
R52050 C9_P_btm.n931 C9_P_btm.n930 0.0556875
R52051 C9_P_btm.n1262 C9_P_btm.n885 0.0556875
R52052 C9_P_btm.n1509 C9_P_btm.n1508 0.0556875
R52053 C9_P_btm.n755 C9_P_btm.n754 0.0556875
R52054 C9_P_btm.n633 C9_P_btm.n632 0.0556875
R52055 C9_P_btm.n255 C9_P_btm.n174 0.0556875
R52056 C9_P_btm.n757 C9_P_btm.n756 0.0556875
R52057 C9_P_btm.n762 C9_P_btm.n134 0.0556875
R52058 C9_P_btm.n884 C9_P_btm.n883 0.0556875
R52059 C9_P_btm.n1511 C9_P_btm.n1510 0.0556875
R52060 C9_P_btm.n1633 C9_P_btm.n1632 0.0556875
R52061 C9_P_btm.n1635 C9_P_btm.n1634 0.0556875
R52062 C9_P_btm.n1640 C9_P_btm.n110 0.0556875
R52063 C9_P_btm.n1671 C9_P_btm.n1670 0.0556875
R52064 C9_P_btm.n1657 C9_P_btm.n1656 0.0556875
R52065 C9_P_btm.n113 C9_P_btm.n104 0.0556875
R52066 C9_P_btm.n1673 C9_P_btm.n1672 0.0556875
R52067 C9_P_btm.n1678 C9_P_btm.n87 0.0556875
R52068 C9_P_btm.n1692 C9_P_btm.n1691 0.0556875
R52069 C9_P_btm.n1694 C9_P_btm.n1693 0.0556875
R52070 C9_P_btm.n1708 C9_P_btm.n1707 0.0556875
R52071 C9_P_btm.n1710 C9_P_btm.n1709 0.0556875
R52072 C9_P_btm.n90 C9_P_btm.n81 0.0556875
R52073 C9_P_btm.n1729 C9_P_btm.n1728 0.0556875
R52074 C9_P_btm.n1715 C9_P_btm.n64 0.0556875
R52075 C9_P_btm.n1745 C9_P_btm.n1744 0.0556875
R52076 C9_P_btm.n1731 C9_P_btm.n1730 0.0556875
R52077 C9_P_btm.n67 C9_P_btm.n58 0.0556875
R52078 C9_P_btm.n1747 C9_P_btm.n1746 0.0556875
R52079 C9_P_btm.n1752 C9_P_btm.n41 0.0556875
R52080 C9_P_btm.n1766 C9_P_btm.n1765 0.0556875
R52081 C9_P_btm.n1768 C9_P_btm.n1767 0.0556875
R52082 C9_P_btm.n1782 C9_P_btm.n1781 0.0556875
R52083 C9_P_btm.n1784 C9_P_btm.n1783 0.0556875
R52084 C9_P_btm.n44 C9_P_btm.n35 0.0556875
R52085 C9_P_btm.n1803 C9_P_btm.n1802 0.0556875
R52086 C9_P_btm.n1789 C9_P_btm.n31 0.0556875
R52087 C9_P_btm.n1834 C9_P_btm.n1833 0.0556875
R52088 C9_P_btm.n1820 C9_P_btm.n1819 0.0556875
R52089 C9_P_btm.n1818 C9_P_btm.n1817 0.0556875
R52090 C9_P_btm.n1836 C9_P_btm.n1835 0.0556875
R52091 C9_P_btm.n1841 C9_P_btm.n21 0.0556875
R52092 C9_P_btm.n1805 C9_P_btm.n1804 0.0556875
R52093 C9_P_btm.n1855 C9_P_btm.n16 0.0556875
R52094 C9_P_btm.n1869 C9_P_btm.n1868 0.0556875
R52095 C9_P_btm.n1871 C9_P_btm.n1870 0.0556875
R52096 C9_P_btm.n1885 C9_P_btm.n1884 0.0556875
R52097 a_n1123_35174.n16 a_n1123_35174.n0 21.0497
R52098 a_n1123_35174.n17 a_n1123_35174.n16 20.1816
R52099 a_n1123_35174.t5 a_n1123_35174.n2 10.7351
R52100 a_n1123_35174.n13 a_n1123_35174.t5 10.7351
R52101 a_n1123_35174.n7 a_n1123_35174.t6 10.7351
R52102 a_n1123_35174.t6 a_n1123_35174.n6 10.7351
R52103 a_n1123_35174.n13 a_n1123_35174.t7 10.7351
R52104 a_n1123_35174.t7 a_n1123_35174.n1 10.7351
R52105 a_n1123_35174.t4 a_n1123_35174.n7 10.7351
R52106 a_n1123_35174.n8 a_n1123_35174.t4 10.7351
R52107 a_n1123_35174.n16 a_n1123_35174.n15 8.273
R52108 a_n1123_35174.n14 a_n1123_35174.n2 6.92882
R52109 a_n1123_35174.n15 a_n1123_35174.n1 6.39231
R52110 a_n1123_35174.n11 a_n1123_35174.n2 5.96815
R52111 a_n1123_35174.n6 a_n1123_35174.n4 5.82388
R52112 a_n1123_35174.n6 a_n1123_35174.n5 5.73036
R52113 a_n1123_35174.n8 a_n1123_35174.n5 5.57405
R52114 a_n1123_35174.n0 a_n1123_35174.t2 4.9505
R52115 a_n1123_35174.n0 a_n1123_35174.t3 4.9505
R52116 a_n1123_35174.n17 a_n1123_35174.t1 4.9505
R52117 a_n1123_35174.t0 a_n1123_35174.n17 4.9505
R52118 a_n1123_35174.n14 a_n1123_35174.n13 3.29479
R52119 a_n1123_35174.n9 a_n1123_35174.n4 3.27414
R52120 a_n1123_35174.n11 a_n1123_35174.n10 3.26815
R52121 a_n1123_35174.n10 a_n1123_35174.n9 3.08441
R52122 a_n1123_35174.n7 a_n1123_35174.n5 2.93762
R52123 a_n1123_35174.n10 a_n1123_35174.n1 2.59444
R52124 a_n1123_35174.n9 a_n1123_35174.n8 2.38669
R52125 a_n1123_35174.n4 a_n1123_35174.n3 2.24404
R52126 a_n1123_35174.n12 a_n1123_35174.n11 2.23808
R52127 a_n1123_35174.n12 a_n1123_35174.n3 1.16457
R52128 a_n1123_35174.n13 a_n1123_35174.n12 0.785683
R52129 a_n1123_35174.n7 a_n1123_35174.n3 0.739928
R52130 a_n1123_35174.n15 a_n1123_35174.n14 0.34925
R52131 w_1375_34946.n37 w_1375_34946.n9 27635.6
R52132 w_1375_34946.n39 w_1375_34946.n35 14784.7
R52133 w_1375_34946.n36 w_1375_34946.n35 14784.7
R52134 w_1375_34946.n39 w_1375_34946.n34 14784.7
R52135 w_1375_34946.n34 w_1375_34946.n7 11195.3
R52136 w_1375_34946.n50 w_1375_34946.n48 3017.65
R52137 w_1375_34946.n59 w_1375_34946.n11 3017.65
R52138 w_1375_34946.n48 w_1375_34946.n11 3017.65
R52139 w_1375_34946.n60 w_1375_34946.n8 1757.65
R52140 w_1375_34946.n10 w_1375_34946.n7 1757.65
R52141 w_1375_34946.n36 w_1375_34946.n10 1711.76
R52142 w_1375_34946.n40 w_1375_34946.n33 1577.04
R52143 w_1375_34946.n41 w_1375_34946.n24 1373.85
R52144 w_1375_34946.n50 w_1375_34946.n8 1080
R52145 w_1375_34946.n32 w_1375_34946.n3 936.235
R52146 w_1375_34946.n63 w_1375_34946.t0 905.04
R52147 w_1375_34946.t0 w_1375_34946.n62 812.54
R52148 w_1375_34946.n39 w_1375_34946.t2 724.569
R52149 w_1375_34946.t5 w_1375_34946.n37 717.962
R52150 w_1375_34946.t2 w_1375_34946.n38 668.146
R52151 w_1375_34946.n38 w_1375_34946.t5 668.146
R52152 w_1375_34946.n65 w_1375_34946.n5 621.553
R52153 w_1375_34946.n24 w_1375_34946.n5 572.612
R52154 w_1375_34946.n63 w_1375_34946.n7 557.648
R52155 w_1375_34946.n63 w_1375_34946.n8 557.648
R52156 w_1375_34946.n61 w_1375_34946.n10 557.648
R52157 w_1375_34946.n61 w_1375_34946.n60 557.648
R52158 w_1375_34946.n33 w_1375_34946.n32 497.599
R52159 w_1375_34946.n58 w_1375_34946.n57 298.877
R52160 w_1375_34946.n53 w_1375_34946.n52 280.202
R52161 w_1375_34946.n56 w_1375_34946.n13 277.776
R52162 w_1375_34946.t1 w_1375_34946.n69 228.215
R52163 w_1375_34946.n41 w_1375_34946.n40 195.883
R52164 w_1375_34946.n12 w_1375_34946.n6 187.482
R52165 w_1375_34946.n66 w_1375_34946.n65 187.482
R52166 w_1375_34946.n66 w_1375_34946.n3 182.589
R52167 w_1375_34946.t10 w_1375_34946.n48 137.529
R52168 w_1375_34946.n51 w_1375_34946.n6 115.201
R52169 w_1375_34946.n62 w_1375_34946.n9 103.859
R52170 w_1375_34946.n61 w_1375_34946.n4 92.5005
R52171 w_1375_34946.n62 w_1375_34946.n61 92.5005
R52172 w_1375_34946.n64 w_1375_34946.n63 92.5005
R52173 w_1375_34946.t14 w_1375_34946.n9 75.2024
R52174 w_1375_34946.t16 w_1375_34946.t14 73.6677
R52175 w_1375_34946.t12 w_1375_34946.t10 73.6677
R52176 w_1375_34946.n17 w_1375_34946.t11 65.4041
R52177 w_1375_34946.n15 w_1375_34946.t15 62.5643
R52178 w_1375_34946.n20 w_1375_34946.t9 61.7296
R52179 w_1375_34946.n23 w_1375_34946.t3 61.7296
R52180 w_1375_34946.n28 w_1375_34946.t7 61.7296
R52181 w_1375_34946.t4 w_1375_34946.n25 61.7296
R52182 w_1375_34946.n60 w_1375_34946.n59 60.0005
R52183 w_1375_34946.n66 w_1375_34946.n4 59.4829
R52184 w_1375_34946.n12 w_1375_34946.n4 59.4829
R52185 w_1375_34946.n65 w_1375_34946.n64 59.4829
R52186 w_1375_34946.n64 w_1375_34946.n6 59.4829
R52187 w_1375_34946.n17 w_1375_34946.n16 56.8163
R52188 w_1375_34946.n22 w_1375_34946.n21 54.1123
R52189 w_1375_34946.n27 w_1375_34946.n26 54.1123
R52190 w_1375_34946.n49 w_1375_34946.t16 36.8341
R52191 w_1375_34946.n49 w_1375_34946.t12 36.8341
R52192 w_1375_34946.n57 w_1375_34946.n11 26.4291
R52193 w_1375_34946.n49 w_1375_34946.n11 26.4291
R52194 w_1375_34946.n51 w_1375_34946.n50 26.4291
R52195 w_1375_34946.n50 w_1375_34946.n49 26.4291
R52196 w_1375_34946.n53 w_1375_34946.n13 20.4805
R52197 w_1375_34946.n52 w_1375_34946.n51 16.9417
R52198 w_1375_34946.n68 w_1375_34946.n1 15.2505
R52199 w_1375_34946.n48 w_1375_34946.n13 13.2148
R52200 w_1375_34946.n59 w_1375_34946.n58 13.2148
R52201 w_1375_34946.n59 w_1375_34946.n9 13.2148
R52202 w_1375_34946.n57 w_1375_34946.n56 8.2968
R52203 w_1375_34946.n16 w_1375_34946.t17 8.12675
R52204 w_1375_34946.n16 w_1375_34946.t13 8.12675
R52205 w_1375_34946.t3 w_1375_34946.n22 7.61783
R52206 w_1375_34946.n22 w_1375_34946.t8 7.61783
R52207 w_1375_34946.n26 w_1375_34946.t4 7.61783
R52208 w_1375_34946.n26 w_1375_34946.t6 7.61783
R52209 w_1375_34946.n36 w_1375_34946.n3 6.60764
R52210 w_1375_34946.n37 w_1375_34946.n36 6.60764
R52211 w_1375_34946.n40 w_1375_34946.n39 6.60764
R52212 w_1375_34946.n31 w_1375_34946.n19 6.41545
R52213 w_1375_34946.n58 w_1375_34946.n12 6.4005
R52214 w_1375_34946.n44 w_1375_34946.n43 6.37679
R52215 w_1375_34946.n18 w_1375_34946.n17 2.72081
R52216 w_1375_34946.n31 w_1375_34946.n30 2.50632
R52217 w_1375_34946.n45 w_1375_34946.n44 2.12421
R52218 w_1375_34946.n34 w_1375_34946.n24 2.03347
R52219 w_1375_34946.n38 w_1375_34946.n34 2.03347
R52220 w_1375_34946.n35 w_1375_34946.n33 2.03347
R52221 w_1375_34946.n38 w_1375_34946.n35 2.03347
R52222 w_1375_34946.n56 w_1375_34946.n55 1.5505
R52223 w_1375_34946.n52 w_1375_34946.n47 1.5505
R52224 w_1375_34946.n55 w_1375_34946.n54 1.26141
R52225 w_1375_34946.n54 w_1375_34946.n53 1.03383
R52226 w_1375_34946.n42 w_1375_34946.n41 1.03383
R52227 w_1375_34946.n67 w_1375_34946.n66 1.03383
R52228 w_1375_34946.n15 w_1375_34946.n14 1.00774
R52229 w_1375_34946.n54 w_1375_34946.n47 0.938644
R52230 w_1375_34946.n27 w_1375_34946.n25 0.891526
R52231 w_1375_34946.n28 w_1375_34946.n27 0.891526
R52232 w_1375_34946.n23 w_1375_34946.n21 0.891526
R52233 w_1375_34946.n21 w_1375_34946.n20 0.891526
R52234 w_1375_34946.n43 w_1375_34946.n19 0.741479
R52235 w_1375_34946.n55 w_1375_34946.n14 0.542875
R52236 w_1375_34946.n46 w_1375_34946.n45 0.494823
R52237 w_1375_34946.n47 w_1375_34946.n46 0.441222
R52238 w_1375_34946.n46 w_1375_34946.n18 0.428803
R52239 w_1375_34946.n29 w_1375_34946.n1 0.286876
R52240 w_1375_34946.n30 w_1375_34946.n29 0.260999
R52241 w_1375_34946.n45 w_1375_34946.n0 0.253077
R52242 w_1375_34946.n32 w_1375_34946.n31 0.227329
R52243 w_1375_34946.n44 w_1375_34946.n5 0.227329
R52244 w_1375_34946.n29 w_1375_34946.n14 0.19304
R52245 w_1375_34946.n2 w_1375_34946.n1 0.178335
R52246 w_1375_34946.n69 w_1375_34946.n68 0.0711522
R52247 w_1375_34946.n2 w_1375_34946.n0 0.0700876
R52248 w_1375_34946.n18 w_1375_34946.n15 0.057539
R52249 w_1375_34946.n25 w_1375_34946.n19 0.0351737
R52250 w_1375_34946.n42 w_1375_34946.n23 0.0340082
R52251 w_1375_34946.n30 w_1375_34946.n28 0.0333481
R52252 w_1375_34946.n20 w_1375_34946.n2 0.0328427
R52253 w_1375_34946.n69 w_1375_34946.n0 0.0303913
R52254 w_1375_34946.n68 w_1375_34946.n67 0.0136119
R52255 w_1375_34946.n43 w_1375_34946.n42 0.0016655
R52256 w_1375_34946.n67 w_1375_34946.n2 0.00137413
R52257 a_22812_30659.n0 a_22812_30659.t9 756.547
R52258 a_22812_30659.n14 a_22812_30659.t5 756.226
R52259 a_22812_30659.n0 a_22812_30659.t17 756.226
R52260 a_22812_30659.n1 a_22812_30659.t10 756.226
R52261 a_22812_30659.n2 a_22812_30659.t16 756.226
R52262 a_22812_30659.n3 a_22812_30659.t6 756.226
R52263 a_22812_30659.n4 a_22812_30659.t8 756.226
R52264 a_22812_30659.n5 a_22812_30659.t4 756.226
R52265 a_22812_30659.n6 a_22812_30659.t12 756.226
R52266 a_22812_30659.n7 a_22812_30659.t18 756.226
R52267 a_22812_30659.n8 a_22812_30659.t14 756.226
R52268 a_22812_30659.n9 a_22812_30659.t19 756.226
R52269 a_22812_30659.n10 a_22812_30659.t15 756.226
R52270 a_22812_30659.n11 a_22812_30659.t11 756.226
R52271 a_22812_30659.n12 a_22812_30659.t7 756.226
R52272 a_22812_30659.n13 a_22812_30659.t13 756.226
R52273 a_22812_30659.n16 a_22812_30659.n15 380.32
R52274 a_22812_30659.n17 a_22812_30659.n16 185
R52275 a_22812_30659.n16 a_22812_30659.n14 102.317
R52276 a_22812_30659.n15 a_22812_30659.t3 26.5955
R52277 a_22812_30659.n15 a_22812_30659.t2 26.5955
R52278 a_22812_30659.t1 a_22812_30659.n17 24.9236
R52279 a_22812_30659.n17 a_22812_30659.t0 24.9236
R52280 a_22812_30659.n13 a_22812_30659.n12 0.3205
R52281 a_22812_30659.n12 a_22812_30659.n11 0.3205
R52282 a_22812_30659.n11 a_22812_30659.n10 0.3205
R52283 a_22812_30659.n10 a_22812_30659.n9 0.3205
R52284 a_22812_30659.n9 a_22812_30659.n8 0.3205
R52285 a_22812_30659.n8 a_22812_30659.n7 0.3205
R52286 a_22812_30659.n7 a_22812_30659.n6 0.3205
R52287 a_22812_30659.n6 a_22812_30659.n5 0.3205
R52288 a_22812_30659.n5 a_22812_30659.n4 0.3205
R52289 a_22812_30659.n4 a_22812_30659.n3 0.3205
R52290 a_22812_30659.n3 a_22812_30659.n2 0.3205
R52291 a_22812_30659.n2 a_22812_30659.n1 0.3205
R52292 a_22812_30659.n1 a_22812_30659.n0 0.3205
R52293 a_22812_30659.n14 a_22812_30659.n13 0.303833
R52294 VREF.n36 VREF.t4 67.0515
R52295 VREF.n0 VREF.t6 67.0515
R52296 VREF.n40 VREF.t52 66.3952
R52297 VREF.n39 VREF.t7 66.3952
R52298 VREF.n38 VREF.t10 66.3952
R52299 VREF.n37 VREF.t71 66.3952
R52300 VREF.n36 VREF.t51 66.3952
R52301 VREF.n4 VREF.t5 66.3952
R52302 VREF.n3 VREF.t72 66.3952
R52303 VREF.n2 VREF.t22 66.3952
R52304 VREF.n1 VREF.t70 66.3952
R52305 VREF.n0 VREF.t73 66.3952
R52306 VREF.n72 VREF.n71 38.8204
R52307 VREF.n71 VREF.t33 34.2201
R52308 VREF.n35 VREF.t65 34.2201
R52309 VREF.n70 VREF.n69 30.6495
R52310 VREF.n68 VREF.n67 30.6495
R52311 VREF.n66 VREF.n65 30.6495
R52312 VREF.n64 VREF.n63 30.6495
R52313 VREF.n62 VREF.n61 30.6495
R52314 VREF.n60 VREF.n59 30.6495
R52315 VREF.n58 VREF.n57 30.6495
R52316 VREF.n56 VREF.n55 30.6495
R52317 VREF.n54 VREF.n53 30.6495
R52318 VREF.n52 VREF.n51 30.6495
R52319 VREF.n50 VREF.n49 30.6495
R52320 VREF.n48 VREF.n47 30.6495
R52321 VREF.n46 VREF.n45 30.6495
R52322 VREF.n44 VREF.n43 30.6495
R52323 VREF.n42 VREF.n41 30.6495
R52324 VREF.n34 VREF.n33 30.6495
R52325 VREF.n32 VREF.n31 30.6495
R52326 VREF.n30 VREF.n29 30.6495
R52327 VREF.n28 VREF.n27 30.6495
R52328 VREF.n26 VREF.n25 30.6495
R52329 VREF.n24 VREF.n23 30.6495
R52330 VREF.n22 VREF.n21 30.6495
R52331 VREF.n20 VREF.n19 30.6495
R52332 VREF.n18 VREF.n17 30.6495
R52333 VREF.n16 VREF.n15 30.6495
R52334 VREF.n14 VREF.n13 30.6495
R52335 VREF.n12 VREF.n11 30.6495
R52336 VREF.n10 VREF.n9 30.6495
R52337 VREF.n8 VREF.n7 30.6495
R52338 VREF.n6 VREF.n5 30.6495
R52339 VREF.n72 VREF.n35 12.7128
R52340 VREF VREF.n72 5.39669
R52341 VREF.n69 VREF.t41 3.57113
R52342 VREF.n69 VREF.t46 3.57113
R52343 VREF.n67 VREF.t38 3.57113
R52344 VREF.n67 VREF.t35 3.57113
R52345 VREF.n65 VREF.t42 3.57113
R52346 VREF.n65 VREF.t39 3.57113
R52347 VREF.n63 VREF.t43 3.57113
R52348 VREF.n63 VREF.t44 3.57113
R52349 VREF.n61 VREF.t40 3.57113
R52350 VREF.n61 VREF.t36 3.57113
R52351 VREF.n59 VREF.t31 3.57113
R52352 VREF.n59 VREF.t34 3.57113
R52353 VREF.n57 VREF.t37 3.57113
R52354 VREF.n57 VREF.t45 3.57113
R52355 VREF.n55 VREF.t32 3.57113
R52356 VREF.n55 VREF.t24 3.57113
R52357 VREF.n53 VREF.t26 3.57113
R52358 VREF.n53 VREF.t30 3.57113
R52359 VREF.n51 VREF.t23 3.57113
R52360 VREF.n51 VREF.t28 3.57113
R52361 VREF.n49 VREF.t27 3.57113
R52362 VREF.n49 VREF.t29 3.57113
R52363 VREF.n47 VREF.t25 3.57113
R52364 VREF.n47 VREF.t48 3.57113
R52365 VREF.n45 VREF.t47 3.57113
R52366 VREF.n45 VREF.t49 3.57113
R52367 VREF.n43 VREF.t50 3.57113
R52368 VREF.n43 VREF.t9 3.57113
R52369 VREF.n41 VREF.t8 3.57113
R52370 VREF.n41 VREF.t19 3.57113
R52371 VREF.n33 VREF.t59 3.57113
R52372 VREF.n33 VREF.t57 3.57113
R52373 VREF.n31 VREF.t64 3.57113
R52374 VREF.n31 VREF.t58 3.57113
R52375 VREF.n29 VREF.t56 3.57113
R52376 VREF.n29 VREF.t62 3.57113
R52377 VREF.n27 VREF.t60 3.57113
R52378 VREF.n27 VREF.t53 3.57113
R52379 VREF.n25 VREF.t67 3.57113
R52380 VREF.n25 VREF.t55 3.57113
R52381 VREF.n23 VREF.t61 3.57113
R52382 VREF.n23 VREF.t63 3.57113
R52383 VREF.n21 VREF.t68 3.57113
R52384 VREF.n21 VREF.t54 3.57113
R52385 VREF.n19 VREF.t14 3.57113
R52386 VREF.n19 VREF.t66 3.57113
R52387 VREF.n17 VREF.t16 3.57113
R52388 VREF.n17 VREF.t11 3.57113
R52389 VREF.n15 VREF.t18 3.57113
R52390 VREF.n15 VREF.t15 3.57113
R52391 VREF.n13 VREF.t12 3.57113
R52392 VREF.n13 VREF.t17 3.57113
R52393 VREF.n11 VREF.t1 3.57113
R52394 VREF.n11 VREF.t13 3.57113
R52395 VREF.n9 VREF.t0 3.57113
R52396 VREF.n9 VREF.t3 3.57113
R52397 VREF.n7 VREF.t20 3.57113
R52398 VREF.n7 VREF.t2 3.57113
R52399 VREF.n5 VREF.t69 3.57113
R52400 VREF.n5 VREF.t21 3.57113
R52401 VREF.n44 VREF.n42 0.71925
R52402 VREF.n46 VREF.n44 0.71925
R52403 VREF.n50 VREF.n48 0.71925
R52404 VREF.n52 VREF.n50 0.71925
R52405 VREF.n56 VREF.n54 0.71925
R52406 VREF.n60 VREF.n58 0.71925
R52407 VREF.n62 VREF.n60 0.71925
R52408 VREF.n66 VREF.n64 0.71925
R52409 VREF.n70 VREF.n68 0.71925
R52410 VREF.n71 VREF.n70 0.71925
R52411 VREF.n8 VREF.n6 0.71925
R52412 VREF.n10 VREF.n8 0.71925
R52413 VREF.n14 VREF.n12 0.71925
R52414 VREF.n16 VREF.n14 0.71925
R52415 VREF.n20 VREF.n18 0.71925
R52416 VREF.n24 VREF.n22 0.71925
R52417 VREF.n26 VREF.n24 0.71925
R52418 VREF.n30 VREF.n28 0.71925
R52419 VREF.n34 VREF.n32 0.71925
R52420 VREF.n35 VREF.n34 0.71925
R52421 VREF.n38 VREF.n37 0.688
R52422 VREF.n48 VREF.n46 0.688
R52423 VREF.n54 VREF.n52 0.688
R52424 VREF.n58 VREF.n56 0.688
R52425 VREF.n64 VREF.n62 0.688
R52426 VREF.n68 VREF.n66 0.688
R52427 VREF.n2 VREF.n1 0.688
R52428 VREF.n12 VREF.n10 0.688
R52429 VREF.n18 VREF.n16 0.688
R52430 VREF.n22 VREF.n20 0.688
R52431 VREF.n28 VREF.n26 0.688
R52432 VREF.n32 VREF.n30 0.688
R52433 VREF.n37 VREF.n36 0.65675
R52434 VREF.n39 VREF.n38 0.65675
R52435 VREF.n40 VREF.n39 0.65675
R52436 VREF.n42 VREF.n40 0.65675
R52437 VREF.n1 VREF.n0 0.65675
R52438 VREF.n3 VREF.n2 0.65675
R52439 VREF.n4 VREF.n3 0.65675
R52440 VREF.n6 VREF.n4 0.65675
R52441 a_n53_44363.n20 a_n53_44363.n0 688.152
R52442 a_n53_44363.n12 a_n53_44363.t15 471.289
R52443 a_n53_44363.n10 a_n53_44363.t14 471.289
R52444 a_n53_44363.n8 a_n53_44363.t19 471.289
R52445 a_n53_44363.n6 a_n53_44363.t6 471.289
R52446 a_n53_44363.n5 a_n53_44363.t11 471.289
R52447 a_n53_44363.n3 a_n53_44363.t12 471.289
R52448 a_n53_44363.n2 a_n53_44363.t4 471.289
R52449 a_n53_44363.n1 a_n53_44363.t18 471.289
R52450 a_n53_44363.n16 a_n53_44363.t22 241.536
R52451 a_n53_44363.n14 a_n53_44363.t21 241.536
R52452 a_n53_44363.n4 a_n53_44363.n2 200.24
R52453 a_n53_44363.n7 a_n53_44363.n5 197.768
R52454 a_n53_44363.n9 a_n53_44363.n8 193.337
R52455 a_n53_44363.n21 a_n53_44363.n20 190.62
R52456 a_n53_44363.n19 a_n53_44363.n1 185.113
R52457 a_n53_44363.n11 a_n53_44363.n10 184.809
R52458 a_n53_44363.n13 a_n53_44363.n12 183.177
R52459 a_n53_44363.n7 a_n53_44363.n6 183.177
R52460 a_n53_44363.n4 a_n53_44363.n3 183.177
R52461 a_n53_44363.n17 a_n53_44363.n16 176.865
R52462 a_n53_44363.n15 a_n53_44363.n14 173.25
R52463 a_n53_44363.n16 a_n53_44363.t16 169.237
R52464 a_n53_44363.n14 a_n53_44363.t9 169.237
R52465 a_n53_44363.n12 a_n53_44363.t8 148.35
R52466 a_n53_44363.n10 a_n53_44363.t13 148.35
R52467 a_n53_44363.n8 a_n53_44363.t23 148.35
R52468 a_n53_44363.n6 a_n53_44363.t5 148.35
R52469 a_n53_44363.n5 a_n53_44363.t20 148.35
R52470 a_n53_44363.n3 a_n53_44363.t7 148.35
R52471 a_n53_44363.n2 a_n53_44363.t10 148.35
R52472 a_n53_44363.n1 a_n53_44363.t17 148.35
R52473 a_n53_44363.n21 a_n53_44363.t0 38.5719
R52474 a_n53_44363.t1 a_n53_44363.n21 38.5719
R52475 a_n53_44363.n0 a_n53_44363.t2 26.5955
R52476 a_n53_44363.n0 a_n53_44363.t3 26.5955
R52477 a_n53_44363.n15 a_n53_44363.n13 25.9869
R52478 a_n53_44363.n9 a_n53_44363.n7 13.2273
R52479 a_n53_44363.n17 a_n53_44363.n15 10.9167
R52480 a_n53_44363.n18 a_n53_44363.n17 10.5293
R52481 a_n53_44363.n18 a_n53_44363.n4 9.62704
R52482 a_n53_44363.n20 a_n53_44363.n19 9.59462
R52483 a_n53_44363.n13 a_n53_44363.n11 6.04462
R52484 a_n53_44363.n19 a_n53_44363.n18 5.58292
R52485 a_n53_44363.n11 a_n53_44363.n9 3.56506
R52486 a_13524_46832.n17 a_13524_46832.n0 620.551
R52487 a_13524_46832.t20 a_13524_46832.t18 618.109
R52488 a_13524_46832.t25 a_13524_46832.t17 547.874
R52489 a_13524_46832.t24 a_13524_46832.t6 397.286
R52490 a_13524_46832.n2 a_13524_46832.t13 377.248
R52491 a_13524_46832.n10 a_13524_46832.t20 361.37
R52492 a_13524_46832.n15 a_13524_46832.t24 353.377
R52493 a_13524_46832.n7 a_13524_46832.t4 322.747
R52494 a_13524_46832.n6 a_13524_46832.t5 305.267
R52495 a_13524_46832.n18 a_13524_46832.n17 258.063
R52496 a_13524_46832.n1 a_13524_46832.t14 229.369
R52497 a_13524_46832.n3 a_13524_46832.t22 223.327
R52498 a_13524_46832.n13 a_13524_46832.t16 212.081
R52499 a_13524_46832.n12 a_13524_46832.t12 212.081
R52500 a_13524_46832.n14 a_13524_46832.n13 205.014
R52501 a_13524_46832.n7 a_13524_46832.t10 194.213
R52502 a_13524_46832.n8 a_13524_46832.n5 192.095
R52503 a_13524_46832.n8 a_13524_46832.n7 188.018
R52504 a_13524_46832.n10 a_13524_46832.n9 180.667
R52505 a_13524_46832.n6 a_13524_46832.t21 179.823
R52506 a_13524_46832.n2 a_13524_46832.t9 174
R52507 a_13524_46832.n9 a_13524_46832.t23 173.34
R52508 a_13524_46832.n16 a_13524_46832.n1 169.988
R52509 a_13524_46832.n9 a_13524_46832.t15 162.81
R52510 a_13524_46832.n1 a_13524_46832.t7 157.07
R52511 a_13524_46832.n13 a_13524_46832.t19 139.78
R52512 a_13524_46832.n12 a_13524_46832.t11 139.78
R52513 a_13524_46832.n5 a_13524_46832.t8 130.27
R52514 a_13524_46832.n7 a_13524_46832.n6 126.803
R52515 a_13524_46832.n4 a_13524_46832.t25 123.43
R52516 a_13524_46832.n13 a_13524_46832.n12 61.346
R52517 a_13524_46832.n4 a_13524_46832.n3 41.3757
R52518 a_13524_46832.n18 a_13524_46832.t0 38.5719
R52519 a_13524_46832.t1 a_13524_46832.n18 38.5719
R52520 a_13524_46832.n0 a_13524_46832.t3 26.5955
R52521 a_13524_46832.n0 a_13524_46832.t2 26.5955
R52522 a_13524_46832.n5 a_13524_46832.n4 24.7519
R52523 a_13524_46832.n16 a_13524_46832.n15 20.0309
R52524 a_13524_46832.n17 a_13524_46832.n16 18.6592
R52525 a_13524_46832.n11 a_13524_46832.n10 7.55957
R52526 a_13524_46832.n11 a_13524_46832.n8 4.97577
R52527 a_13524_46832.n14 a_13524_46832.n11 3.15435
R52528 a_13524_46832.n15 a_13524_46832.n14 2.53724
R52529 a_13524_46832.n3 a_13524_46832.n2 1.78218
R52530 a_1053_45123.n9 a_1053_45123.t8 414.432
R52531 a_1053_45123.n11 a_1053_45123.t1 352.678
R52532 a_1053_45123.n9 a_1053_45123.t11 300.349
R52533 a_1053_45123.t0 a_1053_45123.n11 285.036
R52534 a_1053_45123.n1 a_1053_45123.t3 268.135
R52535 a_1053_45123.n7 a_1053_45123.t5 256.07
R52536 a_1053_45123.n2 a_1053_45123.t10 221.72
R52537 a_1053_45123.n4 a_1053_45123.t6 206.547
R52538 a_1053_45123.n0 a_1053_45123.t9 196.549
R52539 a_1053_45123.n6 a_1053_45123.n0 182.565
R52540 a_1053_45123.n8 a_1053_45123.n7 181.849
R52541 a_1053_45123.n5 a_1053_45123.n1 175.041
R52542 a_1053_45123.n5 a_1053_45123.n4 152
R52543 a_1053_45123.n7 a_1053_45123.t2 150.03
R52544 a_1053_45123.n3 a_1053_45123.t4 149.421
R52545 a_1053_45123.n0 a_1053_45123.t7 148.35
R52546 a_1053_45123.n10 a_1053_45123.n9 99.6442
R52547 a_1053_45123.n6 a_1053_45123.n5 42.2605
R52548 a_1053_45123.n2 a_1053_45123.n1 28.5635
R52549 a_1053_45123.n11 a_1053_45123.n10 26.2998
R52550 a_1053_45123.n3 a_1053_45123.n2 17.8524
R52551 a_1053_45123.n4 a_1053_45123.n3 17.8524
R52552 a_1053_45123.n10 a_1053_45123.n8 11.8527
R52553 a_1053_45123.n8 a_1053_45123.n6 1.71582
R52554 a_9096_45276.t3 a_9096_45276.t2 392.027
R52555 a_9096_45276.n2 a_9096_45276.t1 366.548
R52556 a_9096_45276.n1 a_9096_45276.t3 363.923
R52557 a_9096_45276.n0 a_9096_45276.t4 329.007
R52558 a_9096_45276.t0 a_9096_45276.n2 310.909
R52559 a_9096_45276.n0 a_9096_45276.t5 200.475
R52560 a_9096_45276.n1 a_9096_45276.n0 178.071
R52561 a_9096_45276.n2 a_9096_45276.n1 44.3015
R52562 SMPL_ON_P.n0 SMPL_ON_P.t9 260.322
R52563 SMPL_ON_P.n6 SMPL_ON_P.n4 244.069
R52564 SMPL_ON_P.n3 SMPL_ON_P.n2 236.589
R52565 SMPL_ON_P.n6 SMPL_ON_P.n5 204.893
R52566 SMPL_ON_P.n3 SMPL_ON_P.n1 200.321
R52567 SMPL_ON_P SMPL_ON_P.n0 184.986
R52568 SMPL_ON_P.n0 SMPL_ON_P.t8 175.169
R52569 SMPL_ON_P SMPL_ON_P.n7 71.5326
R52570 SMPL_ON_P.n7 SMPL_ON_P.n6 27.3803
R52571 SMPL_ON_P.n5 SMPL_ON_P.t7 26.5955
R52572 SMPL_ON_P.n5 SMPL_ON_P.t4 26.5955
R52573 SMPL_ON_P.n4 SMPL_ON_P.t5 26.5955
R52574 SMPL_ON_P.n4 SMPL_ON_P.t6 26.5955
R52575 SMPL_ON_P.n1 SMPL_ON_P.t2 24.9236
R52576 SMPL_ON_P.n1 SMPL_ON_P.t0 24.9236
R52577 SMPL_ON_P.n2 SMPL_ON_P.t3 24.9236
R52578 SMPL_ON_P.n2 SMPL_ON_P.t1 24.9236
R52579 SMPL_ON_P.n7 SMPL_ON_P.n3 24.8776
R52580 a_15730_45670.n7 a_15730_45670.t10 293.969
R52581 a_15730_45670.n12 a_15730_45670.t13 261.887
R52582 a_15730_45670.n3 a_15730_45670.n1 248.088
R52583 a_15730_45670.n19 a_15730_45670.t22 241.536
R52584 a_15730_45670.n14 a_15730_45670.t23 241.536
R52585 a_15730_45670.n15 a_15730_45670.t8 236.18
R52586 a_15730_45670.n5 a_15730_45670.t20 230.363
R52587 a_15730_45670.n9 a_15730_45670.t27 212.081
R52588 a_15730_45670.n10 a_15730_45670.t18 212.081
R52589 a_15730_45670.n3 a_15730_45670.n2 208.508
R52590 a_15730_45670.n20 a_15730_45670.n19 198.696
R52591 a_15730_45670.n16 a_15730_45670.n14 184.114
R52592 a_15730_45670.n17 a_15730_45670.n13 181.41
R52593 a_15730_45670.n16 a_15730_45670.n15 173.3
R52594 a_15730_45670.n19 a_15730_45670.t14 169.237
R52595 a_15730_45670.n14 a_15730_45670.t24 169.237
R52596 a_15730_45670.n6 a_15730_45670.n4 167.239
R52597 a_15730_45670.n15 a_15730_45670.t17 163.881
R52598 a_15730_45670.n8 a_15730_45670.n7 163.879
R52599 a_15730_45670.n6 a_15730_45670.n5 163.643
R52600 a_15730_45670.n18 a_15730_45670.n12 162.429
R52601 a_15730_45670.n5 a_15730_45670.t11 158.064
R52602 a_15730_45670.n12 a_15730_45670.t12 155.847
R52603 a_15730_45670.n13 a_15730_45670.t16 142.994
R52604 a_15730_45670.n9 a_15730_45670.t9 139.78
R52605 a_15730_45670.n10 a_15730_45670.t15 139.78
R52606 a_15730_45670.n7 a_15730_45670.t25 138.338
R52607 a_15730_45670.n24 a_15730_45670.n0 137.575
R52608 a_15730_45670.n4 a_15730_45670.t21 137.177
R52609 a_15730_45670.n13 a_15730_45670.t26 126.927
R52610 a_15730_45670.n4 a_15730_45670.t19 121.109
R52611 a_15730_45670.n25 a_15730_45670.n24 99.1749
R52612 a_15730_45670.n21 a_15730_45670.n11 94.1665
R52613 a_15730_45670.n11 a_15730_45670.n9 52.4879
R52614 a_15730_45670.n23 a_15730_45670.n3 38.4831
R52615 a_15730_45670.n1 a_15730_45670.t5 26.5955
R52616 a_15730_45670.n1 a_15730_45670.t6 26.5955
R52617 a_15730_45670.n2 a_15730_45670.t7 26.5955
R52618 a_15730_45670.n2 a_15730_45670.t4 26.5955
R52619 a_15730_45670.n0 a_15730_45670.t0 24.9236
R52620 a_15730_45670.n0 a_15730_45670.t1 24.9236
R52621 a_15730_45670.n25 a_15730_45670.t2 24.9236
R52622 a_15730_45670.t3 a_15730_45670.n25 24.9236
R52623 a_15730_45670.n23 a_15730_45670.n22 24.5725
R52624 a_15730_45670.n22 a_15730_45670.n21 17.2587
R52625 a_15730_45670.n21 a_15730_45670.n20 16.0611
R52626 a_15730_45670.n20 a_15730_45670.n18 15.5566
R52627 a_15730_45670.n24 a_15730_45670.n23 14.8665
R52628 a_15730_45670.n8 a_15730_45670.n6 12.8161
R52629 a_15730_45670.n11 a_15730_45670.n10 9.34851
R52630 a_15730_45670.n18 a_15730_45670.n17 6.78775
R52631 a_15730_45670.n17 a_15730_45670.n16 4.5029
R52632 a_15730_45670.n22 a_15730_45670.n8 1.52676
R52633 a_n1459_43236.n10 a_n1459_43236.n9 329.507
R52634 a_n1459_43236.n6 a_n1459_43236.n5 300.118
R52635 a_n1459_43236.n9 a_n1459_43236.n8 299.834
R52636 a_n1459_43236.n3 a_n1459_43236.n0 293.543
R52637 a_n1459_43236.n6 a_n1459_43236.n4 291.81
R52638 a_n1459_43236.n0 a_n1459_43236.t9 276.464
R52639 a_n1459_43236.n2 a_n1459_43236.t10 212.081
R52640 a_n1459_43236.n1 a_n1459_43236.t13 212.081
R52641 a_n1459_43236.n3 a_n1459_43236.n2 208.338
R52642 a_n1459_43236.n0 a_n1459_43236.t12 196.131
R52643 a_n1459_43236.n2 a_n1459_43236.t11 139.78
R52644 a_n1459_43236.n1 a_n1459_43236.t8 139.78
R52645 a_n1459_43236.n9 a_n1459_43236.n7 78.5231
R52646 a_n1459_43236.n2 a_n1459_43236.n1 61.346
R52647 a_n1459_43236.n8 a_n1459_43236.t3 26.5955
R52648 a_n1459_43236.n8 a_n1459_43236.t2 26.5955
R52649 a_n1459_43236.n5 a_n1459_43236.t6 26.5955
R52650 a_n1459_43236.n5 a_n1459_43236.t7 26.5955
R52651 a_n1459_43236.t0 a_n1459_43236.n10 26.5955
R52652 a_n1459_43236.n10 a_n1459_43236.t1 26.5955
R52653 a_n1459_43236.n4 a_n1459_43236.t5 24.9236
R52654 a_n1459_43236.n4 a_n1459_43236.t4 24.9236
R52655 a_n1459_43236.n7 a_n1459_43236.n3 18.2078
R52656 a_n1459_43236.n7 a_n1459_43236.n6 1.2805
R52657 VDAC_Ni VDAC_Ni.t9 388.632
R52658 VDAC_Ni.n3 VDAC_Ni.t10 231.123
R52659 VDAC_Ni.n2 VDAC_Ni.n0 104.255
R52660 VDAC_Ni.n2 VDAC_Ni.n1 103.96
R52661 VDAC_Ni.n3 VDAC_Ni.t0 50.8513
R52662 VDAC_Ni.n8 VDAC_Ni.n7 37.3168
R52663 VDAC_Ni.n6 VDAC_Ni.n5 37.3168
R52664 VDAC_Ni.n1 VDAC_Ni.t1 16.253
R52665 VDAC_Ni.n1 VDAC_Ni.t2 16.253
R52666 VDAC_Ni.n0 VDAC_Ni.t4 16.253
R52667 VDAC_Ni.n0 VDAC_Ni.t3 16.253
R52668 VDAC_Ni.n7 VDAC_Ni.t7 9.9005
R52669 VDAC_Ni.n7 VDAC_Ni.t8 9.9005
R52670 VDAC_Ni.n5 VDAC_Ni.t5 9.9005
R52671 VDAC_Ni.n5 VDAC_Ni.t6 9.9005
R52672 VDAC_Ni.n9 VDAC_Ni.n8 1.89332
R52673 VDAC_Ni.n4 VDAC_Ni.n2 1.5005
R52674 VDAC_Ni.n4 VDAC_Ni.n3 1.5005
R52675 VDAC_Ni.n6 VDAC_Ni.n4 0.328625
R52676 VDAC_Ni.n8 VDAC_Ni.n6 0.313
R52677 VDAC_Ni.n9 VDAC_Ni 0.016125
R52678 VDAC_Ni VDAC_Ni.n9 0.0112759
R52679 a_10259_42870.n6 a_10259_42870.t13 334.723
R52680 a_10259_42870.n12 a_10259_42870.t23 315.442
R52681 a_10259_42870.n16 a_10259_42870.t12 267.065
R52682 a_10259_42870.n4 a_10259_42870.t8 256.716
R52683 a_10259_42870.n2 a_10259_42870.n0 248.087
R52684 a_10259_42870.n7 a_10259_42870.t20 241.536
R52685 a_10259_42870.n8 a_10259_42870.t16 238.397
R52686 a_10259_42870.n3 a_10259_42870.t17 231.835
R52687 a_10259_42870.n12 a_10259_42870.t21 225.47
R52688 a_10259_42870.n13 a_10259_42870.t11 221.72
R52689 a_10259_42870.n14 a_10259_42870.t25 221.72
R52690 a_10259_42870.n2 a_10259_42870.n1 208.507
R52691 a_10259_42870.n6 a_10259_42870.t24 206.19
R52692 a_10259_42870.n17 a_10259_42870.n16 200.32
R52693 a_10259_42870.n5 a_10259_42870.n4 199.062
R52694 a_10259_42870.n8 a_10259_42870.t14 195.017
R52695 a_10259_42870.n20 a_10259_42870.n6 189.034
R52696 a_10259_42870.n11 a_10259_42870.n7 178.174
R52697 a_10259_42870.n18 a_10259_42870.n12 177.613
R52698 a_10259_42870.n10 a_10259_42870.n9 170.935
R52699 a_10259_42870.n7 a_10259_42870.t19 169.237
R52700 a_10259_42870.n17 a_10259_42870.n15 166.101
R52701 a_10259_42870.n5 a_10259_42870.n3 164.185
R52702 a_10259_42870.n10 a_10259_42870.n8 161.981
R52703 a_10259_42870.n4 a_10259_42870.t22 161.275
R52704 a_10259_42870.n3 a_10259_42870.t27 157.07
R52705 a_10259_42870.n13 a_10259_42870.t10 149.421
R52706 a_10259_42870.n14 a_10259_42870.t9 149.421
R52707 a_10259_42870.n16 a_10259_42870.t18 148.35
R52708 a_10259_42870.n25 a_10259_42870.n24 137.576
R52709 a_10259_42870.n9 a_10259_42870.t26 137.177
R52710 a_10259_42870.n9 a_10259_42870.t15 121.109
R52711 a_10259_42870.n24 a_10259_42870.n23 99.1759
R52712 a_10259_42870.n15 a_10259_42870.n13 37.4894
R52713 a_10259_42870.n15 a_10259_42870.n14 37.4894
R52714 a_10259_42870.n24 a_10259_42870.n22 36.0958
R52715 a_10259_42870.n0 a_10259_42870.t6 26.5955
R52716 a_10259_42870.n0 a_10259_42870.t5 26.5955
R52717 a_10259_42870.n1 a_10259_42870.t7 26.5955
R52718 a_10259_42870.n1 a_10259_42870.t4 26.5955
R52719 a_10259_42870.n23 a_10259_42870.t1 24.9236
R52720 a_10259_42870.n23 a_10259_42870.t0 24.9236
R52721 a_10259_42870.t3 a_10259_42870.n25 24.9236
R52722 a_10259_42870.n25 a_10259_42870.t2 24.9236
R52723 a_10259_42870.n22 a_10259_42870.n2 17.2539
R52724 a_10259_42870.n21 a_10259_42870.n5 16.1653
R52725 a_10259_42870.n21 a_10259_42870.n20 11.9043
R52726 a_10259_42870.n11 a_10259_42870.n10 10.3865
R52727 a_10259_42870.n22 a_10259_42870.n21 9.59462
R52728 a_10259_42870.n19 a_10259_42870.n18 8.61863
R52729 a_10259_42870.n18 a_10259_42870.n17 4.5005
R52730 a_10259_42870.n19 a_10259_42870.n11 2.74363
R52731 a_10259_42870.n20 a_10259_42870.n19 1.51149
R52732 C8_N_btm C8_N_btm.n8 66.3443
R52733 C8_N_btm.n8 C8_N_btm.n7 43.4801
R52734 C8_N_btm.n2 C8_N_btm.n0 33.0333
R52735 C8_N_btm.n2 C8_N_btm.n1 32.3614
R52736 C8_N_btm.n4 C8_N_btm.n2 21.6828
R52737 C8_N_btm.n4 C8_N_btm.n3 20.8888
R52738 C8_N_btm.n6 C8_N_btm.n5 20.8766
R52739 C8_N_btm.n6 C8_N_btm.n4 11.2088
R52740 C8_N_btm.n7 C8_N_btm.t3 9.9005
R52741 C8_N_btm.n7 C8_N_btm.t2 9.9005
R52742 C8_N_btm.n8 C8_N_btm.n6 8.45883
R52743 C8_N_btm C8_N_btm.n903 6.713
R52744 C8_N_btm.n10 C8_N_btm.t270 5.03712
R52745 C8_N_btm.n11 C8_N_btm.t263 5.03712
R52746 C8_N_btm.n12 C8_N_btm.t269 5.03712
R52747 C8_N_btm.n156 C8_N_btm.t264 5.03712
R52748 C8_N_btm.n160 C8_N_btm.t262 5.03712
R52749 C8_N_btm.n159 C8_N_btm.t265 5.03712
R52750 C8_N_btm.n173 C8_N_btm.t268 5.03712
R52751 C8_N_btm.n169 C8_N_btm.t267 5.03712
R52752 C8_N_btm.n890 C8_N_btm.t271 5.03712
R52753 C8_N_btm.n899 C8_N_btm.n898 4.60698
R52754 C8_N_btm.n900 C8_N_btm.n899 4.60698
R52755 C8_N_btm.n896 C8_N_btm.n895 4.60698
R52756 C8_N_btm.n897 C8_N_btm.n896 4.60698
R52757 C8_N_btm.n893 C8_N_btm.n892 4.60698
R52758 C8_N_btm.n894 C8_N_btm.n893 4.60698
R52759 C8_N_btm.n887 C8_N_btm.n886 4.60698
R52760 C8_N_btm.n886 C8_N_btm.n885 4.60698
R52761 C8_N_btm.n884 C8_N_btm.n883 4.60698
R52762 C8_N_btm.n883 C8_N_btm.n882 4.60698
R52763 C8_N_btm.n881 C8_N_btm.n880 4.60698
R52764 C8_N_btm.n880 C8_N_btm.n879 4.60698
R52765 C8_N_btm.n875 C8_N_btm.n874 4.60698
R52766 C8_N_btm.n874 C8_N_btm.n17 4.60698
R52767 C8_N_btm.n872 C8_N_btm.n871 4.60698
R52768 C8_N_btm.n873 C8_N_btm.n872 4.60698
R52769 C8_N_btm.n869 C8_N_btm.n868 4.60698
R52770 C8_N_btm.n870 C8_N_btm.n869 4.60698
R52771 C8_N_btm.n864 C8_N_btm.n863 4.60698
R52772 C8_N_btm.n863 C8_N_btm.n20 4.60698
R52773 C8_N_btm.n841 C8_N_btm.n840 4.60698
R52774 C8_N_btm.n842 C8_N_btm.n841 4.60698
R52775 C8_N_btm.n844 C8_N_btm.n843 4.60698
R52776 C8_N_btm.n845 C8_N_btm.n844 4.60698
R52777 C8_N_btm.n852 C8_N_btm.n851 4.60698
R52778 C8_N_btm.n851 C8_N_btm.n850 4.60698
R52779 C8_N_btm.n855 C8_N_btm.n854 4.60698
R52780 C8_N_btm.n854 C8_N_btm.n853 4.60698
R52781 C8_N_btm.n858 C8_N_btm.n857 4.60698
R52782 C8_N_btm.n857 C8_N_btm.n856 4.60698
R52783 C8_N_btm.n827 C8_N_btm.n826 4.60698
R52784 C8_N_btm.n828 C8_N_btm.n827 4.60698
R52785 C8_N_btm.n830 C8_N_btm.n829 4.60698
R52786 C8_N_btm.n831 C8_N_btm.n830 4.60698
R52787 C8_N_btm.n833 C8_N_btm.n832 4.60698
R52788 C8_N_btm.n834 C8_N_btm.n833 4.60698
R52789 C8_N_btm.n38 C8_N_btm.n37 4.60698
R52790 C8_N_btm.n37 C8_N_btm.n32 4.60698
R52791 C8_N_btm.n35 C8_N_btm.n34 4.60698
R52792 C8_N_btm.n36 C8_N_btm.n35 4.60698
R52793 C8_N_btm.n822 C8_N_btm.n821 4.60698
R52794 C8_N_btm.n821 C8_N_btm.n28 4.60698
R52795 C8_N_btm.n816 C8_N_btm.n815 4.60698
R52796 C8_N_btm.n815 C8_N_btm.n814 4.60698
R52797 C8_N_btm.n813 C8_N_btm.n812 4.60698
R52798 C8_N_btm.n812 C8_N_btm.n811 4.60698
R52799 C8_N_btm.n810 C8_N_btm.n809 4.60698
R52800 C8_N_btm.n809 C8_N_btm.n808 4.60698
R52801 C8_N_btm.n802 C8_N_btm.n801 4.60698
R52802 C8_N_btm.n803 C8_N_btm.n802 4.60698
R52803 C8_N_btm.n799 C8_N_btm.n798 4.60698
R52804 C8_N_btm.n800 C8_N_btm.n799 4.60698
R52805 C8_N_btm.n796 C8_N_btm.n795 4.60698
R52806 C8_N_btm.n797 C8_N_btm.n796 4.60698
R52807 C8_N_btm.n791 C8_N_btm.n790 4.60698
R52808 C8_N_btm.n790 C8_N_btm.n45 4.60698
R52809 C8_N_btm.n52 C8_N_btm.n51 4.60698
R52810 C8_N_btm.n53 C8_N_btm.n52 4.60698
R52811 C8_N_btm.n55 C8_N_btm.n54 4.60698
R52812 C8_N_btm.n54 C8_N_btm.n49 4.60698
R52813 C8_N_btm.n779 C8_N_btm.n778 4.60698
R52814 C8_N_btm.n778 C8_N_btm.n777 4.60698
R52815 C8_N_btm.n782 C8_N_btm.n781 4.60698
R52816 C8_N_btm.n781 C8_N_btm.n780 4.60698
R52817 C8_N_btm.n785 C8_N_btm.n784 4.60698
R52818 C8_N_btm.n784 C8_N_btm.n783 4.60698
R52819 C8_N_btm.n765 C8_N_btm.n764 4.60698
R52820 C8_N_btm.n766 C8_N_btm.n765 4.60698
R52821 C8_N_btm.n768 C8_N_btm.n767 4.60698
R52822 C8_N_btm.n769 C8_N_btm.n768 4.60698
R52823 C8_N_btm.n771 C8_N_btm.n770 4.60698
R52824 C8_N_btm.n772 C8_N_btm.n771 4.60698
R52825 C8_N_btm.n78 C8_N_btm.n77 4.60698
R52826 C8_N_btm.n79 C8_N_btm.n78 4.60698
R52827 C8_N_btm.n75 C8_N_btm.n74 4.60698
R52828 C8_N_btm.n76 C8_N_btm.n75 4.60698
R52829 C8_N_btm.n72 C8_N_btm.n71 4.60698
R52830 C8_N_btm.n73 C8_N_btm.n72 4.60698
R52831 C8_N_btm.n760 C8_N_btm.n759 4.60698
R52832 C8_N_btm.n759 C8_N_btm.n62 4.60698
R52833 C8_N_btm.n754 C8_N_btm.n753 4.60698
R52834 C8_N_btm.n753 C8_N_btm.n752 4.60698
R52835 C8_N_btm.n751 C8_N_btm.n750 4.60698
R52836 C8_N_btm.n750 C8_N_btm.n749 4.60698
R52837 C8_N_btm.n748 C8_N_btm.n747 4.60698
R52838 C8_N_btm.n747 C8_N_btm.n746 4.60698
R52839 C8_N_btm.n745 C8_N_btm.n744 4.60698
R52840 C8_N_btm.n744 C8_N_btm.n743 4.60698
R52841 C8_N_btm.n742 C8_N_btm.n741 4.60698
R52842 C8_N_btm.n741 C8_N_btm.n740 4.60698
R52843 C8_N_btm.n739 C8_N_btm.n738 4.60698
R52844 C8_N_btm.n738 C8_N_btm.n737 4.60698
R52845 C8_N_btm.n81 C8_N_btm.n80 4.60698
R52846 C8_N_btm.n82 C8_N_btm.n81 4.60698
R52847 C8_N_btm.n736 C8_N_btm.n735 4.60698
R52848 C8_N_btm.n735 C8_N_btm.n734 4.60698
R52849 C8_N_btm.n733 C8_N_btm.n732 4.60698
R52850 C8_N_btm.n732 C8_N_btm.n731 4.60698
R52851 C8_N_btm.n730 C8_N_btm.n729 4.60698
R52852 C8_N_btm.n729 C8_N_btm.n728 4.60698
R52853 C8_N_btm.n727 C8_N_btm.n726 4.60698
R52854 C8_N_btm.n726 C8_N_btm.n725 4.60698
R52855 C8_N_btm.n724 C8_N_btm.n723 4.60698
R52856 C8_N_btm.n723 C8_N_btm.n722 4.60698
R52857 C8_N_btm.n721 C8_N_btm.n720 4.60698
R52858 C8_N_btm.n720 C8_N_btm.n719 4.60698
R52859 C8_N_btm.n718 C8_N_btm.n717 4.60698
R52860 C8_N_btm.n717 C8_N_btm.n716 4.60698
R52861 C8_N_btm.n715 C8_N_btm.n714 4.60698
R52862 C8_N_btm.n714 C8_N_btm.n713 4.60698
R52863 C8_N_btm.n712 C8_N_btm.n711 4.60698
R52864 C8_N_btm.n711 C8_N_btm.n710 4.60698
R52865 C8_N_btm.n709 C8_N_btm.n708 4.60698
R52866 C8_N_btm.n708 C8_N_btm.n707 4.60698
R52867 C8_N_btm.n706 C8_N_btm.n705 4.60698
R52868 C8_N_btm.n705 C8_N_btm.n704 4.60698
R52869 C8_N_btm.n703 C8_N_btm.n702 4.60698
R52870 C8_N_btm.n702 C8_N_btm.n701 4.60698
R52871 C8_N_btm.n700 C8_N_btm.n699 4.60698
R52872 C8_N_btm.n699 C8_N_btm.n698 4.60698
R52873 C8_N_btm.n697 C8_N_btm.n696 4.60698
R52874 C8_N_btm.n696 C8_N_btm.n695 4.60698
R52875 C8_N_btm.n694 C8_N_btm.n693 4.60698
R52876 C8_N_btm.n693 C8_N_btm.n692 4.60698
R52877 C8_N_btm.n691 C8_N_btm.n690 4.60698
R52878 C8_N_btm.n690 C8_N_btm.n689 4.60698
R52879 C8_N_btm.n688 C8_N_btm.n687 4.60698
R52880 C8_N_btm.n687 C8_N_btm.n686 4.60698
R52881 C8_N_btm.n685 C8_N_btm.n684 4.60698
R52882 C8_N_btm.n684 C8_N_btm.n683 4.60698
R52883 C8_N_btm.n682 C8_N_btm.n681 4.60698
R52884 C8_N_btm.n681 C8_N_btm.n680 4.60698
R52885 C8_N_btm.n679 C8_N_btm.n678 4.60698
R52886 C8_N_btm.n678 C8_N_btm.n677 4.60698
R52887 C8_N_btm.n676 C8_N_btm.n675 4.60698
R52888 C8_N_btm.n675 C8_N_btm.n674 4.60698
R52889 C8_N_btm.n673 C8_N_btm.n672 4.60698
R52890 C8_N_btm.n672 C8_N_btm.n671 4.60698
R52891 C8_N_btm.n665 C8_N_btm.n664 4.60698
R52892 C8_N_btm.n666 C8_N_btm.n665 4.60698
R52893 C8_N_btm.n662 C8_N_btm.n661 4.60698
R52894 C8_N_btm.n663 C8_N_btm.n662 4.60698
R52895 C8_N_btm.n659 C8_N_btm.n658 4.60698
R52896 C8_N_btm.n660 C8_N_btm.n659 4.60698
R52897 C8_N_btm.n656 C8_N_btm.n655 4.60698
R52898 C8_N_btm.n657 C8_N_btm.n656 4.60698
R52899 C8_N_btm.n653 C8_N_btm.n652 4.60698
R52900 C8_N_btm.n654 C8_N_btm.n653 4.60698
R52901 C8_N_btm.n650 C8_N_btm.n649 4.60698
R52902 C8_N_btm.n651 C8_N_btm.n650 4.60698
R52903 C8_N_btm.n647 C8_N_btm.n646 4.60698
R52904 C8_N_btm.n648 C8_N_btm.n647 4.60698
R52905 C8_N_btm.n644 C8_N_btm.n643 4.60698
R52906 C8_N_btm.n645 C8_N_btm.n644 4.60698
R52907 C8_N_btm.n641 C8_N_btm.n640 4.60698
R52908 C8_N_btm.n642 C8_N_btm.n641 4.60698
R52909 C8_N_btm.n638 C8_N_btm.n637 4.60698
R52910 C8_N_btm.n639 C8_N_btm.n638 4.60698
R52911 C8_N_btm.n635 C8_N_btm.n634 4.60698
R52912 C8_N_btm.n636 C8_N_btm.n635 4.60698
R52913 C8_N_btm.n632 C8_N_btm.n631 4.60698
R52914 C8_N_btm.n633 C8_N_btm.n632 4.60698
R52915 C8_N_btm.n629 C8_N_btm.n628 4.60698
R52916 C8_N_btm.n630 C8_N_btm.n629 4.60698
R52917 C8_N_btm.n626 C8_N_btm.n625 4.60698
R52918 C8_N_btm.n627 C8_N_btm.n626 4.60698
R52919 C8_N_btm.n623 C8_N_btm.n622 4.60698
R52920 C8_N_btm.n624 C8_N_btm.n623 4.60698
R52921 C8_N_btm.n620 C8_N_btm.n619 4.60698
R52922 C8_N_btm.n621 C8_N_btm.n620 4.60698
R52923 C8_N_btm.n617 C8_N_btm.n616 4.60698
R52924 C8_N_btm.n618 C8_N_btm.n617 4.60698
R52925 C8_N_btm.n614 C8_N_btm.n613 4.60698
R52926 C8_N_btm.n615 C8_N_btm.n614 4.60698
R52927 C8_N_btm.n611 C8_N_btm.n610 4.60698
R52928 C8_N_btm.n612 C8_N_btm.n611 4.60698
R52929 C8_N_btm.n608 C8_N_btm.n607 4.60698
R52930 C8_N_btm.n609 C8_N_btm.n608 4.60698
R52931 C8_N_btm.n605 C8_N_btm.n604 4.60698
R52932 C8_N_btm.n606 C8_N_btm.n605 4.60698
R52933 C8_N_btm.n602 C8_N_btm.n601 4.60698
R52934 C8_N_btm.n603 C8_N_btm.n602 4.60698
R52935 C8_N_btm.n599 C8_N_btm.n598 4.60698
R52936 C8_N_btm.n600 C8_N_btm.n599 4.60698
R52937 C8_N_btm.n596 C8_N_btm.n595 4.60698
R52938 C8_N_btm.n597 C8_N_btm.n596 4.60698
R52939 C8_N_btm.n593 C8_N_btm.n592 4.60698
R52940 C8_N_btm.n594 C8_N_btm.n593 4.60698
R52941 C8_N_btm.n590 C8_N_btm.n589 4.60698
R52942 C8_N_btm.n591 C8_N_btm.n590 4.60698
R52943 C8_N_btm.n587 C8_N_btm.n586 4.60698
R52944 C8_N_btm.n588 C8_N_btm.n587 4.60698
R52945 C8_N_btm.n584 C8_N_btm.n583 4.60698
R52946 C8_N_btm.n585 C8_N_btm.n584 4.60698
R52947 C8_N_btm.n579 C8_N_btm.n578 4.60698
R52948 C8_N_btm.n578 C8_N_btm.n351 4.60698
R52949 C8_N_btm.n409 C8_N_btm.n408 4.60698
R52950 C8_N_btm.n410 C8_N_btm.n409 4.60698
R52951 C8_N_btm.n412 C8_N_btm.n411 4.60698
R52952 C8_N_btm.n413 C8_N_btm.n412 4.60698
R52953 C8_N_btm.n415 C8_N_btm.n414 4.60698
R52954 C8_N_btm.n416 C8_N_btm.n415 4.60698
R52955 C8_N_btm.n418 C8_N_btm.n417 4.60698
R52956 C8_N_btm.n419 C8_N_btm.n418 4.60698
R52957 C8_N_btm.n421 C8_N_btm.n420 4.60698
R52958 C8_N_btm.n422 C8_N_btm.n421 4.60698
R52959 C8_N_btm.n424 C8_N_btm.n423 4.60698
R52960 C8_N_btm.n425 C8_N_btm.n424 4.60698
R52961 C8_N_btm.n427 C8_N_btm.n426 4.60698
R52962 C8_N_btm.n428 C8_N_btm.n427 4.60698
R52963 C8_N_btm.n430 C8_N_btm.n429 4.60698
R52964 C8_N_btm.n431 C8_N_btm.n430 4.60698
R52965 C8_N_btm.n433 C8_N_btm.n432 4.60698
R52966 C8_N_btm.n434 C8_N_btm.n433 4.60698
R52967 C8_N_btm.n436 C8_N_btm.n435 4.60698
R52968 C8_N_btm.n437 C8_N_btm.n436 4.60698
R52969 C8_N_btm.n439 C8_N_btm.n438 4.60698
R52970 C8_N_btm.n440 C8_N_btm.n439 4.60698
R52971 C8_N_btm.n442 C8_N_btm.n441 4.60698
R52972 C8_N_btm.n443 C8_N_btm.n442 4.60698
R52973 C8_N_btm.n445 C8_N_btm.n444 4.60698
R52974 C8_N_btm.n446 C8_N_btm.n445 4.60698
R52975 C8_N_btm.n448 C8_N_btm.n447 4.60698
R52976 C8_N_btm.n449 C8_N_btm.n448 4.60698
R52977 C8_N_btm.n451 C8_N_btm.n450 4.60698
R52978 C8_N_btm.n452 C8_N_btm.n451 4.60698
R52979 C8_N_btm.n454 C8_N_btm.n453 4.60698
R52980 C8_N_btm.n455 C8_N_btm.n454 4.60698
R52981 C8_N_btm.n457 C8_N_btm.n456 4.60698
R52982 C8_N_btm.n458 C8_N_btm.n457 4.60698
R52983 C8_N_btm.n460 C8_N_btm.n459 4.60698
R52984 C8_N_btm.n461 C8_N_btm.n460 4.60698
R52985 C8_N_btm.n463 C8_N_btm.n462 4.60698
R52986 C8_N_btm.n464 C8_N_btm.n463 4.60698
R52987 C8_N_btm.n466 C8_N_btm.n465 4.60698
R52988 C8_N_btm.n467 C8_N_btm.n466 4.60698
R52989 C8_N_btm.n469 C8_N_btm.n468 4.60698
R52990 C8_N_btm.n470 C8_N_btm.n469 4.60698
R52991 C8_N_btm.n472 C8_N_btm.n471 4.60698
R52992 C8_N_btm.n473 C8_N_btm.n472 4.60698
R52993 C8_N_btm.n475 C8_N_btm.n474 4.60698
R52994 C8_N_btm.n476 C8_N_btm.n475 4.60698
R52995 C8_N_btm.n478 C8_N_btm.n477 4.60698
R52996 C8_N_btm.n479 C8_N_btm.n478 4.60698
R52997 C8_N_btm.n481 C8_N_btm.n480 4.60698
R52998 C8_N_btm.n482 C8_N_btm.n481 4.60698
R52999 C8_N_btm.n484 C8_N_btm.n483 4.60698
R53000 C8_N_btm.n485 C8_N_btm.n484 4.60698
R53001 C8_N_btm.n487 C8_N_btm.n486 4.60698
R53002 C8_N_btm.n486 C8_N_btm.n381 4.60698
R53003 C8_N_btm.n492 C8_N_btm.n491 4.60698
R53004 C8_N_btm.n493 C8_N_btm.n492 4.60698
R53005 C8_N_btm.n495 C8_N_btm.n494 4.60698
R53006 C8_N_btm.n496 C8_N_btm.n495 4.60698
R53007 C8_N_btm.n498 C8_N_btm.n497 4.60698
R53008 C8_N_btm.n499 C8_N_btm.n498 4.60698
R53009 C8_N_btm.n501 C8_N_btm.n500 4.60698
R53010 C8_N_btm.n502 C8_N_btm.n501 4.60698
R53011 C8_N_btm.n504 C8_N_btm.n503 4.60698
R53012 C8_N_btm.n505 C8_N_btm.n504 4.60698
R53013 C8_N_btm.n507 C8_N_btm.n506 4.60698
R53014 C8_N_btm.n508 C8_N_btm.n507 4.60698
R53015 C8_N_btm.n510 C8_N_btm.n509 4.60698
R53016 C8_N_btm.n511 C8_N_btm.n510 4.60698
R53017 C8_N_btm.n513 C8_N_btm.n512 4.60698
R53018 C8_N_btm.n514 C8_N_btm.n513 4.60698
R53019 C8_N_btm.n516 C8_N_btm.n515 4.60698
R53020 C8_N_btm.n517 C8_N_btm.n516 4.60698
R53021 C8_N_btm.n519 C8_N_btm.n518 4.60698
R53022 C8_N_btm.n520 C8_N_btm.n519 4.60698
R53023 C8_N_btm.n522 C8_N_btm.n521 4.60698
R53024 C8_N_btm.n523 C8_N_btm.n522 4.60698
R53025 C8_N_btm.n525 C8_N_btm.n524 4.60698
R53026 C8_N_btm.n526 C8_N_btm.n525 4.60698
R53027 C8_N_btm.n528 C8_N_btm.n527 4.60698
R53028 C8_N_btm.n529 C8_N_btm.n528 4.60698
R53029 C8_N_btm.n531 C8_N_btm.n530 4.60698
R53030 C8_N_btm.n532 C8_N_btm.n531 4.60698
R53031 C8_N_btm.n535 C8_N_btm.n534 4.60698
R53032 C8_N_btm.n534 C8_N_btm.n533 4.60698
R53033 C8_N_btm.n537 C8_N_btm.n536 4.60698
R53034 C8_N_btm.n538 C8_N_btm.n537 4.60698
R53035 C8_N_btm.n540 C8_N_btm.n539 4.60698
R53036 C8_N_btm.n541 C8_N_btm.n540 4.60698
R53037 C8_N_btm.n543 C8_N_btm.n542 4.60698
R53038 C8_N_btm.n544 C8_N_btm.n543 4.60698
R53039 C8_N_btm.n546 C8_N_btm.n545 4.60698
R53040 C8_N_btm.n547 C8_N_btm.n546 4.60698
R53041 C8_N_btm.n549 C8_N_btm.n548 4.60698
R53042 C8_N_btm.n550 C8_N_btm.n549 4.60698
R53043 C8_N_btm.n552 C8_N_btm.n551 4.60698
R53044 C8_N_btm.n553 C8_N_btm.n552 4.60698
R53045 C8_N_btm.n555 C8_N_btm.n554 4.60698
R53046 C8_N_btm.n556 C8_N_btm.n555 4.60698
R53047 C8_N_btm.n558 C8_N_btm.n557 4.60698
R53048 C8_N_btm.n559 C8_N_btm.n558 4.60698
R53049 C8_N_btm.n561 C8_N_btm.n560 4.60698
R53050 C8_N_btm.n562 C8_N_btm.n561 4.60698
R53051 C8_N_btm.n564 C8_N_btm.n563 4.60698
R53052 C8_N_btm.n565 C8_N_btm.n564 4.60698
R53053 C8_N_btm.n567 C8_N_btm.n566 4.60698
R53054 C8_N_btm.n568 C8_N_btm.n567 4.60698
R53055 C8_N_btm.n570 C8_N_btm.n569 4.60698
R53056 C8_N_btm.n571 C8_N_btm.n570 4.60698
R53057 C8_N_btm.n573 C8_N_btm.n572 4.60698
R53058 C8_N_btm.n574 C8_N_btm.n573 4.60698
R53059 C8_N_btm.n318 C8_N_btm.n317 4.60698
R53060 C8_N_btm.n319 C8_N_btm.n318 4.60698
R53061 C8_N_btm.n315 C8_N_btm.n314 4.60698
R53062 C8_N_btm.n316 C8_N_btm.n315 4.60698
R53063 C8_N_btm.n312 C8_N_btm.n311 4.60698
R53064 C8_N_btm.n313 C8_N_btm.n312 4.60698
R53065 C8_N_btm.n309 C8_N_btm.n308 4.60698
R53066 C8_N_btm.n310 C8_N_btm.n309 4.60698
R53067 C8_N_btm.n299 C8_N_btm.n298 4.60698
R53068 C8_N_btm.n298 C8_N_btm.n297 4.60698
R53069 C8_N_btm.n296 C8_N_btm.n295 4.60698
R53070 C8_N_btm.n295 C8_N_btm.n294 4.60698
R53071 C8_N_btm.n293 C8_N_btm.n292 4.60698
R53072 C8_N_btm.n292 C8_N_btm.n291 4.60698
R53073 C8_N_btm.n287 C8_N_btm.n286 4.60698
R53074 C8_N_btm.n286 C8_N_btm.n115 4.60698
R53075 C8_N_btm.n284 C8_N_btm.n283 4.60698
R53076 C8_N_btm.n285 C8_N_btm.n284 4.60698
R53077 C8_N_btm.n281 C8_N_btm.n280 4.60698
R53078 C8_N_btm.n282 C8_N_btm.n281 4.60698
R53079 C8_N_btm.n276 C8_N_btm.n275 4.60698
R53080 C8_N_btm.n275 C8_N_btm.n118 4.60698
R53081 C8_N_btm.n253 C8_N_btm.n252 4.60698
R53082 C8_N_btm.n254 C8_N_btm.n253 4.60698
R53083 C8_N_btm.n256 C8_N_btm.n255 4.60698
R53084 C8_N_btm.n257 C8_N_btm.n256 4.60698
R53085 C8_N_btm.n264 C8_N_btm.n263 4.60698
R53086 C8_N_btm.n263 C8_N_btm.n262 4.60698
R53087 C8_N_btm.n267 C8_N_btm.n266 4.60698
R53088 C8_N_btm.n266 C8_N_btm.n265 4.60698
R53089 C8_N_btm.n270 C8_N_btm.n269 4.60698
R53090 C8_N_btm.n269 C8_N_btm.n268 4.60698
R53091 C8_N_btm.n239 C8_N_btm.n238 4.60698
R53092 C8_N_btm.n240 C8_N_btm.n239 4.60698
R53093 C8_N_btm.n242 C8_N_btm.n241 4.60698
R53094 C8_N_btm.n243 C8_N_btm.n242 4.60698
R53095 C8_N_btm.n245 C8_N_btm.n244 4.60698
R53096 C8_N_btm.n246 C8_N_btm.n245 4.60698
R53097 C8_N_btm.n136 C8_N_btm.n135 4.60698
R53098 C8_N_btm.n135 C8_N_btm.n130 4.60698
R53099 C8_N_btm.n133 C8_N_btm.n132 4.60698
R53100 C8_N_btm.n134 C8_N_btm.n133 4.60698
R53101 C8_N_btm.n234 C8_N_btm.n233 4.60698
R53102 C8_N_btm.n233 C8_N_btm.n126 4.60698
R53103 C8_N_btm.n228 C8_N_btm.n227 4.60698
R53104 C8_N_btm.n227 C8_N_btm.n226 4.60698
R53105 C8_N_btm.n225 C8_N_btm.n224 4.60698
R53106 C8_N_btm.n224 C8_N_btm.n223 4.60698
R53107 C8_N_btm.n222 C8_N_btm.n221 4.60698
R53108 C8_N_btm.n221 C8_N_btm.n220 4.60698
R53109 C8_N_btm.n214 C8_N_btm.n213 4.60698
R53110 C8_N_btm.n215 C8_N_btm.n214 4.60698
R53111 C8_N_btm.n211 C8_N_btm.n210 4.60698
R53112 C8_N_btm.n212 C8_N_btm.n211 4.60698
R53113 C8_N_btm.n208 C8_N_btm.n207 4.60698
R53114 C8_N_btm.n209 C8_N_btm.n208 4.60698
R53115 C8_N_btm.n203 C8_N_btm.n202 4.60698
R53116 C8_N_btm.n202 C8_N_btm.n143 4.60698
R53117 C8_N_btm.n150 C8_N_btm.n149 4.60698
R53118 C8_N_btm.n151 C8_N_btm.n150 4.60698
R53119 C8_N_btm.n153 C8_N_btm.n152 4.60698
R53120 C8_N_btm.n152 C8_N_btm.n147 4.60698
R53121 C8_N_btm.n191 C8_N_btm.n190 4.60698
R53122 C8_N_btm.n190 C8_N_btm.n189 4.60698
R53123 C8_N_btm.n194 C8_N_btm.n193 4.60698
R53124 C8_N_btm.n193 C8_N_btm.n192 4.60698
R53125 C8_N_btm.n197 C8_N_btm.n196 4.60698
R53126 C8_N_btm.n196 C8_N_btm.n195 4.60698
R53127 C8_N_btm.n177 C8_N_btm.n176 4.60698
R53128 C8_N_btm.n178 C8_N_btm.n177 4.60698
R53129 C8_N_btm.n180 C8_N_btm.n179 4.60698
R53130 C8_N_btm.n181 C8_N_btm.n180 4.60698
R53131 C8_N_btm.n183 C8_N_btm.n182 4.60698
R53132 C8_N_btm.n184 C8_N_btm.n183 4.60698
R53133 C8_N_btm.n164 C8_N_btm.n163 4.60698
R53134 C8_N_btm.n163 C8_N_btm.n162 4.60698
R53135 C8_N_btm.n167 C8_N_btm.n166 4.60698
R53136 C8_N_btm.n166 C8_N_btm.n165 4.60698
R53137 C8_N_btm.n172 C8_N_btm.n171 4.60698
R53138 C8_N_btm.n171 C8_N_btm.n168 4.60698
R53139 C8_N_btm.n306 C8_N_btm.n305 4.60698
R53140 C8_N_btm.n307 C8_N_btm.n306 4.60698
R53141 C8_N_btm.n903 C8_N_btm.t266 4.03712
R53142 C8_N_btm.n901 C8_N_btm.t236 3.98193
R53143 C8_N_btm.n878 C8_N_btm.t137 3.98193
R53144 C8_N_btm.n837 C8_N_btm.t163 3.98193
R53145 C8_N_btm.n846 C8_N_btm.t76 3.98193
R53146 C8_N_btm.n849 C8_N_btm.t257 3.98193
R53147 C8_N_btm.n835 C8_N_btm.t248 3.98193
R53148 C8_N_btm.n31 C8_N_btm.t39 3.98193
R53149 C8_N_btm.n807 C8_N_btm.t61 3.98193
R53150 C8_N_btm.n804 C8_N_btm.t12 3.98193
R53151 C8_N_btm.n48 C8_N_btm.t144 3.98193
R53152 C8_N_btm.n776 C8_N_btm.t24 3.98193
R53153 C8_N_btm.n773 C8_N_btm.t192 3.98193
R53154 C8_N_btm.n83 C8_N_btm.t204 3.98193
R53155 C8_N_btm.n670 C8_N_btm.t261 3.98193
R53156 C8_N_btm.n667 C8_N_btm.t159 3.98193
R53157 C8_N_btm.n380 C8_N_btm.t187 3.98193
R53158 C8_N_btm.n490 C8_N_btm.t254 3.98193
R53159 C8_N_btm.n365 C8_N_btm.t149 3.98193
R53160 C8_N_btm.n366 C8_N_btm.t230 3.98193
R53161 C8_N_btm.n575 C8_N_btm.t9 3.98193
R53162 C8_N_btm.n577 C8_N_btm.t73 3.98193
R53163 C8_N_btm.n582 C8_N_btm.t53 3.98193
R53164 C8_N_btm.n320 C8_N_btm.t234 3.98193
R53165 C8_N_btm.n290 C8_N_btm.t209 3.98193
R53166 C8_N_btm.n249 C8_N_btm.t34 3.98193
R53167 C8_N_btm.n258 C8_N_btm.t14 3.98193
R53168 C8_N_btm.n261 C8_N_btm.t7 3.98193
R53169 C8_N_btm.n247 C8_N_btm.t72 3.98193
R53170 C8_N_btm.n129 C8_N_btm.t52 3.98193
R53171 C8_N_btm.n219 C8_N_btm.t132 3.98193
R53172 C8_N_btm.n216 C8_N_btm.t110 3.98193
R53173 C8_N_btm.n146 C8_N_btm.t89 3.98193
R53174 C8_N_btm.n188 C8_N_btm.t180 3.98193
R53175 C8_N_btm.n185 C8_N_btm.t148 3.98193
R53176 C8_N_btm.n161 C8_N_btm.t99 3.98193
R53177 C8_N_btm.n170 C8_N_btm.t138 3.98193
R53178 C8_N_btm.n175 C8_N_btm.t117 3.98193
R53179 C8_N_btm.n198 C8_N_btm.t77 3.98193
R53180 C8_N_btm.n201 C8_N_btm.t213 3.98193
R53181 C8_N_btm.n206 C8_N_btm.t19 3.98193
R53182 C8_N_btm.n229 C8_N_btm.t40 3.98193
R53183 C8_N_btm.n232 C8_N_btm.t214 3.98193
R53184 C8_N_btm.n237 C8_N_btm.t189 3.98193
R53185 C8_N_btm.n271 C8_N_btm.t140 3.98193
R53186 C8_N_btm.n274 C8_N_btm.t164 3.98193
R53187 C8_N_btm.n279 C8_N_btm.t193 3.98193
R53188 C8_N_btm.n300 C8_N_btm.t100 3.98193
R53189 C8_N_btm.n304 C8_N_btm.t256 3.98193
R53190 C8_N_btm.n755 C8_N_btm.t28 3.98193
R53191 C8_N_btm.n758 C8_N_btm.t111 3.98193
R53192 C8_N_btm.n763 C8_N_btm.t90 3.98193
R53193 C8_N_btm.n786 C8_N_btm.t181 3.98193
R53194 C8_N_btm.n789 C8_N_btm.t150 3.98193
R53195 C8_N_btm.n794 C8_N_btm.t260 3.98193
R53196 C8_N_btm.n817 C8_N_btm.t225 3.98193
R53197 C8_N_btm.n820 C8_N_btm.t197 3.98193
R53198 C8_N_btm.n825 C8_N_btm.t242 3.98193
R53199 C8_N_btm.n859 C8_N_btm.t10 3.98193
R53200 C8_N_btm.n862 C8_N_btm.t240 3.98193
R53201 C8_N_btm.n867 C8_N_btm.t65 3.98193
R53202 C8_N_btm.n888 C8_N_btm.t45 3.98193
R53203 C8_N_btm.n891 C8_N_btm.t124 3.98193
R53204 C8_N_btm.n1 C8_N_btm.t273 3.57113
R53205 C8_N_btm.n1 C8_N_btm.t272 3.57113
R53206 C8_N_btm.n0 C8_N_btm.t274 3.57113
R53207 C8_N_btm.n0 C8_N_btm.t275 3.57113
R53208 C8_N_btm.n3 C8_N_btm.t5 2.4755
R53209 C8_N_btm.n3 C8_N_btm.t4 2.4755
R53210 C8_N_btm.n5 C8_N_btm.t0 2.4755
R53211 C8_N_btm.n5 C8_N_btm.t1 2.4755
R53212 C8_N_btm.n899 C8_N_btm.t172 1.67819
R53213 C8_N_btm.n896 C8_N_btm.t143 1.67819
R53214 C8_N_btm.n893 C8_N_btm.t188 1.67819
R53215 C8_N_btm.n886 C8_N_btm.t255 1.67819
R53216 C8_N_btm.n883 C8_N_btm.t165 1.67819
R53217 C8_N_btm.n880 C8_N_btm.t84 1.67819
R53218 C8_N_btm.n874 C8_N_btm.t105 1.67819
R53219 C8_N_btm.n872 C8_N_btm.t194 1.67819
R53220 C8_N_btm.n869 C8_N_btm.t247 1.67819
R53221 C8_N_btm.n863 C8_N_btm.t36 1.67819
R53222 C8_N_btm.n841 C8_N_btm.t101 1.67819
R53223 C8_N_btm.n844 C8_N_btm.t54 1.67819
R53224 C8_N_btm.n851 C8_N_btm.t47 1.67819
R53225 C8_N_btm.n854 C8_N_btm.t251 1.67819
R53226 C8_N_btm.n857 C8_N_btm.t241 1.67819
R53227 C8_N_btm.n827 C8_N_btm.t79 1.67819
R53228 C8_N_btm.n830 C8_N_btm.t145 1.67819
R53229 C8_N_btm.n833 C8_N_btm.t67 1.67819
R53230 C8_N_btm.n37 C8_N_btm.t32 1.67819
R53231 C8_N_btm.n35 C8_N_btm.t63 1.67819
R53232 C8_N_btm.n821 C8_N_btm.t177 1.67819
R53233 C8_N_btm.n815 C8_N_btm.t22 1.67819
R53234 C8_N_btm.n812 C8_N_btm.t85 1.67819
R53235 C8_N_btm.n809 C8_N_btm.t58 1.67819
R53236 C8_N_btm.n802 C8_N_btm.t175 1.67819
R53237 C8_N_btm.n799 C8_N_btm.t103 1.67819
R53238 C8_N_btm.n796 C8_N_btm.t191 1.67819
R53239 C8_N_btm.n790 C8_N_btm.t215 1.67819
R53240 C8_N_btm.n52 C8_N_btm.t57 1.67819
R53241 C8_N_btm.n54 C8_N_btm.t199 1.67819
R53242 C8_N_btm.n778 C8_N_btm.t227 1.67819
R53243 C8_N_btm.n781 C8_N_btm.t48 1.67819
R53244 C8_N_btm.n784 C8_N_btm.t239 1.67819
R53245 C8_N_btm.n765 C8_N_btm.t141 1.67819
R53246 C8_N_btm.n768 C8_N_btm.t221 1.67819
R53247 C8_N_btm.n771 C8_N_btm.t128 1.67819
R53248 C8_N_btm.n78 C8_N_btm.t217 1.67819
R53249 C8_N_btm.n75 C8_N_btm.t153 1.67819
R53250 C8_N_btm.n72 C8_N_btm.t244 1.67819
R53251 C8_N_btm.n759 C8_N_btm.t167 1.67819
R53252 C8_N_btm.n753 C8_N_btm.t80 1.67819
R53253 C8_N_btm.n750 C8_N_btm.t146 1.67819
R53254 C8_N_btm.n747 C8_N_btm.t69 1.67819
R53255 C8_N_btm.n744 C8_N_btm.t249 1.67819
R53256 C8_N_btm.n741 C8_N_btm.t120 1.67819
R53257 C8_N_btm.n738 C8_N_btm.t109 1.67819
R53258 C8_N_btm.n81 C8_N_btm.t139 1.67819
R53259 C8_N_btm.n735 C8_N_btm.t166 1.67819
R53260 C8_N_btm.n732 C8_N_btm.t86 1.67819
R53261 C8_N_btm.n729 C8_N_btm.t151 1.67819
R53262 C8_N_btm.n726 C8_N_btm.t216 1.67819
R53263 C8_N_btm.n723 C8_N_btm.t123 1.67819
R53264 C8_N_btm.n720 C8_N_btm.t201 1.67819
R53265 C8_N_btm.n717 C8_N_btm.t115 1.67819
R53266 C8_N_btm.n714 C8_N_btm.t170 1.67819
R53267 C8_N_btm.n711 C8_N_btm.t6 1.67819
R53268 C8_N_btm.n708 C8_N_btm.t156 1.67819
R53269 C8_N_btm.n705 C8_N_btm.t220 1.67819
R53270 C8_N_btm.n702 C8_N_btm.t17 1.67819
R53271 C8_N_btm.n699 C8_N_btm.t208 1.67819
R53272 C8_N_btm.n696 C8_N_btm.t41 1.67819
R53273 C8_N_btm.n693 C8_N_btm.t179 1.67819
R53274 C8_N_btm.n690 C8_N_btm.t97 1.67819
R53275 C8_N_btm.n687 C8_N_btm.t44 1.67819
R53276 C8_N_btm.n684 C8_N_btm.t235 1.67819
R53277 C8_N_btm.n681 C8_N_btm.t42 1.67819
R53278 C8_N_btm.n678 C8_N_btm.t96 1.67819
R53279 C8_N_btm.n675 C8_N_btm.t18 1.67819
R53280 C8_N_btm.n672 C8_N_btm.t68 1.67819
R53281 C8_N_btm.n665 C8_N_btm.t91 1.67819
R53282 C8_N_btm.n662 C8_N_btm.t38 1.67819
R53283 C8_N_btm.n659 C8_N_btm.t161 1.67819
R53284 C8_N_btm.n656 C8_N_btm.t62 1.67819
R53285 C8_N_btm.n653 C8_N_btm.t186 1.67819
R53286 C8_N_btm.n650 C8_N_btm.t64 1.67819
R53287 C8_N_btm.n647 C8_N_btm.t15 1.67819
R53288 C8_N_btm.n644 C8_N_btm.t203 1.67819
R53289 C8_N_btm.n641 C8_N_btm.t121 1.67819
R53290 C8_N_btm.n638 C8_N_btm.t233 1.67819
R53291 C8_N_btm.n635 C8_N_btm.t37 1.67819
R53292 C8_N_btm.n632 C8_N_btm.t11 1.67819
R53293 C8_N_btm.n629 C8_N_btm.t183 1.67819
R53294 C8_N_btm.n626 C8_N_btm.t243 1.67819
R53295 C8_N_btm.n623 C8_N_btm.t196 1.67819
R53296 C8_N_btm.n620 C8_N_btm.t134 1.67819
R53297 C8_N_btm.n617 C8_N_btm.t228 1.67819
R53298 C8_N_btm.n614 C8_N_btm.t147 1.67819
R53299 C8_N_btm.n611 C8_N_btm.t8 1.67819
R53300 C8_N_btm.n608 C8_N_btm.t182 1.67819
R53301 C8_N_btm.n605 C8_N_btm.t106 1.67819
R53302 C8_N_btm.n602 C8_N_btm.t195 1.67819
R53303 C8_N_btm.n599 C8_N_btm.t131 1.67819
R53304 C8_N_btm.n596 C8_N_btm.t78 1.67819
R53305 C8_N_btm.n593 C8_N_btm.t142 1.67819
R53306 C8_N_btm.n590 C8_N_btm.t92 1.67819
R53307 C8_N_btm.n587 C8_N_btm.t176 1.67819
R53308 C8_N_btm.n584 C8_N_btm.t102 1.67819
R53309 C8_N_btm.n578 C8_N_btm.t122 1.67819
R53310 C8_N_btm.n409 C8_N_btm.t200 1.67819
R53311 C8_N_btm.n412 C8_N_btm.t114 1.67819
R53312 C8_N_btm.n415 C8_N_btm.t169 1.67819
R53313 C8_N_btm.n418 C8_N_btm.t258 1.67819
R53314 C8_N_btm.n421 C8_N_btm.t155 1.67819
R53315 C8_N_btm.n424 C8_N_btm.t219 1.67819
R53316 C8_N_btm.n427 C8_N_btm.t126 1.67819
R53317 C8_N_btm.n430 C8_N_btm.t207 1.67819
R53318 C8_N_btm.n433 C8_N_btm.t94 1.67819
R53319 C8_N_btm.n436 C8_N_btm.t178 1.67819
R53320 C8_N_btm.n439 C8_N_btm.t259 1.67819
R53321 C8_N_btm.n442 C8_N_btm.t160 1.67819
R53322 C8_N_btm.n445 C8_N_btm.t224 1.67819
R53323 C8_N_btm.n448 C8_N_btm.t31 1.67819
R53324 C8_N_btm.n451 C8_N_btm.t211 1.67819
R53325 C8_N_btm.n454 C8_N_btm.t23 1.67819
R53326 C8_N_btm.n457 C8_N_btm.t59 1.67819
R53327 C8_N_btm.n460 C8_N_btm.t218 1.67819
R53328 C8_N_btm.n463 C8_N_btm.t50 1.67819
R53329 C8_N_btm.n466 C8_N_btm.t229 1.67819
R53330 C8_N_btm.n469 C8_N_btm.t35 1.67819
R53331 C8_N_btm.n472 C8_N_btm.t88 1.67819
R53332 C8_N_btm.n475 C8_N_btm.t21 1.67819
R53333 C8_N_btm.n478 C8_N_btm.t83 1.67819
R53334 C8_N_btm.n481 C8_N_btm.t136 1.67819
R53335 C8_N_btm.n484 C8_N_btm.t60 1.67819
R53336 C8_N_btm.n486 C8_N_btm.t113 1.67819
R53337 C8_N_btm.n492 C8_N_btm.t29 1.67819
R53338 C8_N_btm.n495 C8_N_btm.t238 1.67819
R53339 C8_N_btm.n498 C8_N_btm.t56 1.67819
R53340 C8_N_btm.n501 C8_N_btm.t246 1.67819
R53341 C8_N_btm.n504 C8_N_btm.t93 1.67819
R53342 C8_N_btm.n507 C8_N_btm.t133 1.67819
R53343 C8_N_btm.n510 C8_N_btm.t210 1.67819
R53344 C8_N_btm.n513 C8_N_btm.t130 1.67819
R53345 C8_N_btm.n516 C8_N_btm.t222 1.67819
R53346 C8_N_btm.n519 C8_N_btm.t158 1.67819
R53347 C8_N_btm.n522 C8_N_btm.t237 1.67819
R53348 C8_N_btm.n525 C8_N_btm.t173 1.67819
R53349 C8_N_btm.n528 C8_N_btm.t118 1.67819
R53350 C8_N_btm.n531 C8_N_btm.t205 1.67819
R53351 C8_N_btm.n534 C8_N_btm.t125 1.67819
R53352 C8_N_btm.n537 C8_N_btm.t74 1.67819
R53353 C8_N_btm.n540 C8_N_btm.t154 1.67819
R53354 C8_N_btm.n543 C8_N_btm.t87 1.67819
R53355 C8_N_btm.n546 C8_N_btm.t168 1.67819
R53356 C8_N_btm.n549 C8_N_btm.t112 1.67819
R53357 C8_N_btm.n552 C8_N_btm.t49 1.67819
R53358 C8_N_btm.n555 C8_N_btm.t252 1.67819
R53359 C8_N_btm.n558 C8_N_btm.t71 1.67819
R53360 C8_N_btm.n561 C8_N_btm.t20 1.67819
R53361 C8_N_btm.n564 C8_N_btm.t81 1.67819
R53362 C8_N_btm.n567 C8_N_btm.t30 1.67819
R53363 C8_N_btm.n570 C8_N_btm.t107 1.67819
R53364 C8_N_btm.n573 C8_N_btm.t43 1.67819
R53365 C8_N_btm.n318 C8_N_btm.t152 1.67819
R53366 C8_N_btm.n315 C8_N_btm.t98 1.67819
R53367 C8_N_btm.n312 C8_N_btm.t185 1.67819
R53368 C8_N_btm.n309 C8_N_btm.t250 1.67819
R53369 C8_N_btm.n298 C8_N_btm.t157 1.67819
R53370 C8_N_btm.n295 C8_N_btm.t75 1.67819
R53371 C8_N_btm.n292 C8_N_btm.t127 1.67819
R53372 C8_N_btm.n286 C8_N_btm.t226 1.67819
R53373 C8_N_btm.n284 C8_N_btm.t162 1.67819
R53374 C8_N_btm.n281 C8_N_btm.t223 1.67819
R53375 C8_N_btm.n275 C8_N_btm.t232 1.67819
R53376 C8_N_btm.n253 C8_N_btm.t135 1.67819
R53377 C8_N_btm.n256 C8_N_btm.t198 1.67819
R53378 C8_N_btm.n263 C8_N_btm.t174 1.67819
R53379 C8_N_btm.n266 C8_N_btm.t119 1.67819
R53380 C8_N_btm.n269 C8_N_btm.t206 1.67819
R53381 C8_N_btm.n239 C8_N_btm.t33 1.67819
R53382 C8_N_btm.n242 C8_N_btm.t212 1.67819
R53383 C8_N_btm.n245 C8_N_btm.t26 1.67819
R53384 C8_N_btm.n135 C8_N_btm.t27 1.67819
R53385 C8_N_btm.n133 C8_N_btm.t184 1.67819
R53386 C8_N_btm.n233 C8_N_btm.t13 1.67819
R53387 C8_N_btm.n227 C8_N_btm.t95 1.67819
R53388 C8_N_btm.n224 C8_N_btm.t16 1.67819
R53389 C8_N_btm.n221 C8_N_btm.t66 1.67819
R53390 C8_N_btm.n214 C8_N_btm.t46 1.67819
R53391 C8_N_btm.n211 C8_N_btm.t245 1.67819
R53392 C8_N_btm.n208 C8_N_btm.t70 1.67819
R53393 C8_N_btm.n202 C8_N_btm.t51 1.67819
R53394 C8_N_btm.n150 C8_N_btm.t231 1.67819
R53395 C8_N_btm.n152 C8_N_btm.t25 1.67819
R53396 C8_N_btm.n190 C8_N_btm.t104 1.67819
R53397 C8_N_btm.n193 C8_N_btm.t55 1.67819
R53398 C8_N_btm.n196 C8_N_btm.t129 1.67819
R53399 C8_N_btm.n177 C8_N_btm.t108 1.67819
R53400 C8_N_btm.n180 C8_N_btm.t253 1.67819
R53401 C8_N_btm.n183 C8_N_btm.t82 1.67819
R53402 C8_N_btm.n163 C8_N_btm.t171 1.67819
R53403 C8_N_btm.n166 C8_N_btm.t116 1.67819
R53404 C8_N_btm.n171 C8_N_btm.t202 1.67819
R53405 C8_N_btm.n306 C8_N_btm.t190 1.67819
R53406 C8_N_btm.n84 C8_N_btm.n83 1.05569
R53407 C8_N_btm.n367 C8_N_btm.n366 1.05569
R53408 C8_N_btm.n365 C8_N_btm.n364 1.05569
R53409 C8_N_btm.n576 C8_N_btm.n575 1.05569
R53410 C8_N_btm.n490 C8_N_btm.n322 1.05569
R53411 C8_N_btm.n304 C8_N_btm.n101 1.05569
R53412 C8_N_btm.n14 C8_N_btm.n12 1.0005
R53413 C8_N_btm.n15 C8_N_btm.n11 1.0005
R53414 C8_N_btm.n877 C8_N_btm.n10 1.0005
R53415 C8_N_btm.n877 C8_N_btm.n876 1.0005
R53416 C8_N_btm.n18 C8_N_btm.n15 1.0005
R53417 C8_N_btm.n866 C8_N_btm.n14 1.0005
R53418 C8_N_btm.n866 C8_N_btm.n865 1.0005
R53419 C8_N_btm.n839 C8_N_btm.n18 1.0005
R53420 C8_N_btm.n876 C8_N_btm.n16 1.0005
R53421 C8_N_btm.n23 C8_N_btm.n16 1.0005
R53422 C8_N_btm.n839 C8_N_btm.n22 1.0005
R53423 C8_N_btm.n865 C8_N_btm.n19 1.0005
R53424 C8_N_btm.n824 C8_N_btm.n19 1.0005
R53425 C8_N_btm.n26 C8_N_btm.n22 1.0005
R53426 C8_N_btm.n25 C8_N_btm.n23 1.0005
R53427 C8_N_btm.n39 C8_N_btm.n25 1.0005
R53428 C8_N_btm.n33 C8_N_btm.n26 1.0005
R53429 C8_N_btm.n824 C8_N_btm.n823 1.0005
R53430 C8_N_btm.n823 C8_N_btm.n27 1.0005
R53431 C8_N_btm.n33 C8_N_btm.n30 1.0005
R53432 C8_N_btm.n40 C8_N_btm.n39 1.0005
R53433 C8_N_btm.n42 C8_N_btm.n40 1.0005
R53434 C8_N_btm.n43 C8_N_btm.n30 1.0005
R53435 C8_N_btm.n793 C8_N_btm.n27 1.0005
R53436 C8_N_btm.n793 C8_N_btm.n792 1.0005
R53437 C8_N_btm.n50 C8_N_btm.n43 1.0005
R53438 C8_N_btm.n56 C8_N_btm.n42 1.0005
R53439 C8_N_btm.n57 C8_N_btm.n56 1.0005
R53440 C8_N_btm.n50 C8_N_btm.n47 1.0005
R53441 C8_N_btm.n792 C8_N_btm.n44 1.0005
R53442 C8_N_btm.n762 C8_N_btm.n44 1.0005
R53443 C8_N_btm.n60 C8_N_btm.n47 1.0005
R53444 C8_N_btm.n59 C8_N_btm.n57 1.0005
R53445 C8_N_btm.n69 C8_N_btm.n59 1.0005
R53446 C8_N_btm.n70 C8_N_btm.n60 1.0005
R53447 C8_N_btm.n762 C8_N_btm.n761 1.0005
R53448 C8_N_btm.n761 C8_N_btm.n61 1.0005
R53449 C8_N_btm.n70 C8_N_btm.n64 1.0005
R53450 C8_N_btm.n69 C8_N_btm.n65 1.0005
R53451 C8_N_btm.n66 C8_N_btm.n58 1.0005
R53452 C8_N_btm.n68 C8_N_btm.n67 1.0005
R53453 C8_N_btm.n323 C8_N_btm.n106 1.0005
R53454 C8_N_btm.n324 C8_N_btm.n105 1.0005
R53455 C8_N_btm.n325 C8_N_btm.n104 1.0005
R53456 C8_N_btm.n326 C8_N_btm.n103 1.0005
R53457 C8_N_btm.n327 C8_N_btm.n102 1.0005
R53458 C8_N_btm.n328 C8_N_btm.n101 1.0005
R53459 C8_N_btm.n329 C8_N_btm.n100 1.0005
R53460 C8_N_btm.n330 C8_N_btm.n99 1.0005
R53461 C8_N_btm.n331 C8_N_btm.n98 1.0005
R53462 C8_N_btm.n332 C8_N_btm.n97 1.0005
R53463 C8_N_btm.n333 C8_N_btm.n96 1.0005
R53464 C8_N_btm.n334 C8_N_btm.n95 1.0005
R53465 C8_N_btm.n335 C8_N_btm.n94 1.0005
R53466 C8_N_btm.n336 C8_N_btm.n93 1.0005
R53467 C8_N_btm.n337 C8_N_btm.n92 1.0005
R53468 C8_N_btm.n338 C8_N_btm.n91 1.0005
R53469 C8_N_btm.n339 C8_N_btm.n90 1.0005
R53470 C8_N_btm.n340 C8_N_btm.n89 1.0005
R53471 C8_N_btm.n341 C8_N_btm.n88 1.0005
R53472 C8_N_btm.n342 C8_N_btm.n87 1.0005
R53473 C8_N_btm.n343 C8_N_btm.n86 1.0005
R53474 C8_N_btm.n344 C8_N_btm.n85 1.0005
R53475 C8_N_btm.n345 C8_N_btm.n84 1.0005
R53476 C8_N_btm.n346 C8_N_btm.n67 1.0005
R53477 C8_N_btm.n347 C8_N_btm.n66 1.0005
R53478 C8_N_btm.n348 C8_N_btm.n65 1.0005
R53479 C8_N_btm.n349 C8_N_btm.n64 1.0005
R53480 C8_N_btm.n581 C8_N_btm.n61 1.0005
R53481 C8_N_btm.n581 C8_N_btm.n580 1.0005
R53482 C8_N_btm.n407 C8_N_btm.n349 1.0005
R53483 C8_N_btm.n406 C8_N_btm.n348 1.0005
R53484 C8_N_btm.n405 C8_N_btm.n347 1.0005
R53485 C8_N_btm.n404 C8_N_btm.n346 1.0005
R53486 C8_N_btm.n403 C8_N_btm.n345 1.0005
R53487 C8_N_btm.n402 C8_N_btm.n344 1.0005
R53488 C8_N_btm.n401 C8_N_btm.n343 1.0005
R53489 C8_N_btm.n400 C8_N_btm.n342 1.0005
R53490 C8_N_btm.n399 C8_N_btm.n341 1.0005
R53491 C8_N_btm.n398 C8_N_btm.n340 1.0005
R53492 C8_N_btm.n397 C8_N_btm.n339 1.0005
R53493 C8_N_btm.n396 C8_N_btm.n338 1.0005
R53494 C8_N_btm.n395 C8_N_btm.n337 1.0005
R53495 C8_N_btm.n394 C8_N_btm.n336 1.0005
R53496 C8_N_btm.n393 C8_N_btm.n335 1.0005
R53497 C8_N_btm.n392 C8_N_btm.n334 1.0005
R53498 C8_N_btm.n391 C8_N_btm.n333 1.0005
R53499 C8_N_btm.n390 C8_N_btm.n332 1.0005
R53500 C8_N_btm.n389 C8_N_btm.n331 1.0005
R53501 C8_N_btm.n388 C8_N_btm.n330 1.0005
R53502 C8_N_btm.n387 C8_N_btm.n329 1.0005
R53503 C8_N_btm.n386 C8_N_btm.n328 1.0005
R53504 C8_N_btm.n385 C8_N_btm.n327 1.0005
R53505 C8_N_btm.n384 C8_N_btm.n326 1.0005
R53506 C8_N_btm.n383 C8_N_btm.n325 1.0005
R53507 C8_N_btm.n382 C8_N_btm.n324 1.0005
R53508 C8_N_btm.n488 C8_N_btm.n323 1.0005
R53509 C8_N_btm.n489 C8_N_btm.n488 1.0005
R53510 C8_N_btm.n382 C8_N_btm.n379 1.0005
R53511 C8_N_btm.n383 C8_N_btm.n378 1.0005
R53512 C8_N_btm.n384 C8_N_btm.n377 1.0005
R53513 C8_N_btm.n385 C8_N_btm.n376 1.0005
R53514 C8_N_btm.n386 C8_N_btm.n375 1.0005
R53515 C8_N_btm.n387 C8_N_btm.n374 1.0005
R53516 C8_N_btm.n388 C8_N_btm.n373 1.0005
R53517 C8_N_btm.n389 C8_N_btm.n372 1.0005
R53518 C8_N_btm.n390 C8_N_btm.n371 1.0005
R53519 C8_N_btm.n391 C8_N_btm.n370 1.0005
R53520 C8_N_btm.n392 C8_N_btm.n369 1.0005
R53521 C8_N_btm.n393 C8_N_btm.n368 1.0005
R53522 C8_N_btm.n394 C8_N_btm.n367 1.0005
R53523 C8_N_btm.n395 C8_N_btm.n364 1.0005
R53524 C8_N_btm.n396 C8_N_btm.n363 1.0005
R53525 C8_N_btm.n397 C8_N_btm.n362 1.0005
R53526 C8_N_btm.n398 C8_N_btm.n361 1.0005
R53527 C8_N_btm.n399 C8_N_btm.n360 1.0005
R53528 C8_N_btm.n400 C8_N_btm.n359 1.0005
R53529 C8_N_btm.n401 C8_N_btm.n358 1.0005
R53530 C8_N_btm.n402 C8_N_btm.n357 1.0005
R53531 C8_N_btm.n403 C8_N_btm.n356 1.0005
R53532 C8_N_btm.n404 C8_N_btm.n355 1.0005
R53533 C8_N_btm.n405 C8_N_btm.n354 1.0005
R53534 C8_N_btm.n406 C8_N_btm.n353 1.0005
R53535 C8_N_btm.n407 C8_N_btm.n352 1.0005
R53536 C8_N_btm.n580 C8_N_btm.n350 1.0005
R53537 C8_N_btm.n668 C8_N_btm.n322 1.0005
R53538 C8_N_btm.n756 C8_N_btm.n63 1.0005
R53539 C8_N_btm.n576 C8_N_btm.n63 1.0005
R53540 C8_N_btm.n108 C8_N_btm.n106 1.0005
R53541 C8_N_btm.n109 C8_N_btm.n105 1.0005
R53542 C8_N_btm.n110 C8_N_btm.n104 1.0005
R53543 C8_N_btm.n112 C8_N_btm.n110 1.0005
R53544 C8_N_btm.n113 C8_N_btm.n109 1.0005
R53545 C8_N_btm.n289 C8_N_btm.n108 1.0005
R53546 C8_N_btm.n289 C8_N_btm.n288 1.0005
R53547 C8_N_btm.n116 C8_N_btm.n113 1.0005
R53548 C8_N_btm.n278 C8_N_btm.n112 1.0005
R53549 C8_N_btm.n278 C8_N_btm.n277 1.0005
R53550 C8_N_btm.n251 C8_N_btm.n116 1.0005
R53551 C8_N_btm.n288 C8_N_btm.n114 1.0005
R53552 C8_N_btm.n121 C8_N_btm.n114 1.0005
R53553 C8_N_btm.n251 C8_N_btm.n120 1.0005
R53554 C8_N_btm.n277 C8_N_btm.n117 1.0005
R53555 C8_N_btm.n236 C8_N_btm.n117 1.0005
R53556 C8_N_btm.n124 C8_N_btm.n120 1.0005
R53557 C8_N_btm.n123 C8_N_btm.n121 1.0005
R53558 C8_N_btm.n137 C8_N_btm.n123 1.0005
R53559 C8_N_btm.n131 C8_N_btm.n124 1.0005
R53560 C8_N_btm.n236 C8_N_btm.n235 1.0005
R53561 C8_N_btm.n235 C8_N_btm.n125 1.0005
R53562 C8_N_btm.n131 C8_N_btm.n128 1.0005
R53563 C8_N_btm.n138 C8_N_btm.n137 1.0005
R53564 C8_N_btm.n140 C8_N_btm.n138 1.0005
R53565 C8_N_btm.n141 C8_N_btm.n128 1.0005
R53566 C8_N_btm.n205 C8_N_btm.n125 1.0005
R53567 C8_N_btm.n205 C8_N_btm.n204 1.0005
R53568 C8_N_btm.n148 C8_N_btm.n141 1.0005
R53569 C8_N_btm.n154 C8_N_btm.n140 1.0005
R53570 C8_N_btm.n155 C8_N_btm.n154 1.0005
R53571 C8_N_btm.n148 C8_N_btm.n145 1.0005
R53572 C8_N_btm.n204 C8_N_btm.n142 1.0005
R53573 C8_N_btm.n174 C8_N_btm.n142 1.0005
R53574 C8_N_btm.n158 C8_N_btm.n145 1.0005
R53575 C8_N_btm.n157 C8_N_btm.n155 1.0005
R53576 C8_N_btm.n160 C8_N_btm.n157 1.0005
R53577 C8_N_btm.n159 C8_N_btm.n158 1.0005
R53578 C8_N_btm.n174 C8_N_btm.n173 1.0005
R53579 C8_N_btm.n169 C8_N_btm.n144 1.0005
R53580 C8_N_btm.n186 C8_N_btm.n156 1.0005
R53581 C8_N_btm.n187 C8_N_btm.n186 1.0005
R53582 C8_N_btm.n199 C8_N_btm.n144 1.0005
R53583 C8_N_btm.n200 C8_N_btm.n199 1.0005
R53584 C8_N_btm.n187 C8_N_btm.n139 1.0005
R53585 C8_N_btm.n217 C8_N_btm.n139 1.0005
R53586 C8_N_btm.n200 C8_N_btm.n127 1.0005
R53587 C8_N_btm.n230 C8_N_btm.n127 1.0005
R53588 C8_N_btm.n218 C8_N_btm.n217 1.0005
R53589 C8_N_btm.n218 C8_N_btm.n122 1.0005
R53590 C8_N_btm.n231 C8_N_btm.n230 1.0005
R53591 C8_N_btm.n231 C8_N_btm.n119 1.0005
R53592 C8_N_btm.n248 C8_N_btm.n122 1.0005
R53593 C8_N_btm.n260 C8_N_btm.n248 1.0005
R53594 C8_N_btm.n272 C8_N_btm.n119 1.0005
R53595 C8_N_btm.n273 C8_N_btm.n272 1.0005
R53596 C8_N_btm.n260 C8_N_btm.n259 1.0005
R53597 C8_N_btm.n259 C8_N_btm.n250 1.0005
R53598 C8_N_btm.n273 C8_N_btm.n111 1.0005
R53599 C8_N_btm.n301 C8_N_btm.n111 1.0005
R53600 C8_N_btm.n250 C8_N_btm.n107 1.0005
R53601 C8_N_btm.n321 C8_N_btm.n107 1.0005
R53602 C8_N_btm.n302 C8_N_btm.n301 1.0005
R53603 C8_N_btm.n302 C8_N_btm.n103 1.0005
R53604 C8_N_btm.n303 C8_N_btm.n102 1.0005
R53605 C8_N_btm.n669 C8_N_btm.n321 1.0005
R53606 C8_N_btm.n669 C8_N_btm.n668 1.0005
R53607 C8_N_btm.n757 C8_N_btm.n46 1.0005
R53608 C8_N_btm.n757 C8_N_btm.n756 1.0005
R53609 C8_N_btm.n775 C8_N_btm.n774 1.0005
R53610 C8_N_btm.n774 C8_N_btm.n58 1.0005
R53611 C8_N_btm.n788 C8_N_btm.n787 1.0005
R53612 C8_N_btm.n787 C8_N_btm.n46 1.0005
R53613 C8_N_btm.n805 C8_N_btm.n41 1.0005
R53614 C8_N_btm.n775 C8_N_btm.n41 1.0005
R53615 C8_N_btm.n818 C8_N_btm.n29 1.0005
R53616 C8_N_btm.n788 C8_N_btm.n29 1.0005
R53617 C8_N_btm.n806 C8_N_btm.n24 1.0005
R53618 C8_N_btm.n806 C8_N_btm.n805 1.0005
R53619 C8_N_btm.n819 C8_N_btm.n21 1.0005
R53620 C8_N_btm.n819 C8_N_btm.n818 1.0005
R53621 C8_N_btm.n848 C8_N_btm.n836 1.0005
R53622 C8_N_btm.n836 C8_N_btm.n24 1.0005
R53623 C8_N_btm.n861 C8_N_btm.n860 1.0005
R53624 C8_N_btm.n860 C8_N_btm.n21 1.0005
R53625 C8_N_btm.n847 C8_N_btm.n838 1.0005
R53626 C8_N_btm.n848 C8_N_btm.n847 1.0005
R53627 C8_N_btm.n889 C8_N_btm.n13 1.0005
R53628 C8_N_btm.n861 C8_N_btm.n13 1.0005
R53629 C8_N_btm.n902 C8_N_btm.n9 1.0005
R53630 C8_N_btm.n838 C8_N_btm.n9 1.0005
R53631 C8_N_btm.n890 C8_N_btm.n889 1.0005
R53632 C8_N_btm.n903 C8_N_btm.n902 1.0005
R53633 C8_N_btm.n366 C8_N_btm.n365 0.733338
R53634 C8_N_btm.n83 C8_N_btm.n82 0.679419
R53635 C8_N_btm.n575 C8_N_btm.n574 0.679419
R53636 C8_N_btm.n491 C8_N_btm.n490 0.679419
R53637 C8_N_btm.n381 C8_N_btm.n380 0.679419
R53638 C8_N_btm.n579 C8_N_btm.n577 0.679419
R53639 C8_N_btm.n583 C8_N_btm.n582 0.679419
R53640 C8_N_btm.n667 C8_N_btm.n666 0.679419
R53641 C8_N_btm.n172 C8_N_btm.n170 0.679419
R53642 C8_N_btm.n162 C8_N_btm.n161 0.679419
R53643 C8_N_btm.n185 C8_N_btm.n184 0.679419
R53644 C8_N_btm.n176 C8_N_btm.n175 0.679419
R53645 C8_N_btm.n198 C8_N_btm.n197 0.679419
R53646 C8_N_btm.n189 C8_N_btm.n188 0.679419
R53647 C8_N_btm.n147 C8_N_btm.n146 0.679419
R53648 C8_N_btm.n203 C8_N_btm.n201 0.679419
R53649 C8_N_btm.n207 C8_N_btm.n206 0.679419
R53650 C8_N_btm.n216 C8_N_btm.n215 0.679419
R53651 C8_N_btm.n220 C8_N_btm.n219 0.679419
R53652 C8_N_btm.n229 C8_N_btm.n228 0.679419
R53653 C8_N_btm.n234 C8_N_btm.n232 0.679419
R53654 C8_N_btm.n130 C8_N_btm.n129 0.679419
R53655 C8_N_btm.n247 C8_N_btm.n246 0.679419
R53656 C8_N_btm.n238 C8_N_btm.n237 0.679419
R53657 C8_N_btm.n271 C8_N_btm.n270 0.679419
R53658 C8_N_btm.n262 C8_N_btm.n261 0.679419
R53659 C8_N_btm.n258 C8_N_btm.n257 0.679419
R53660 C8_N_btm.n276 C8_N_btm.n274 0.679419
R53661 C8_N_btm.n280 C8_N_btm.n279 0.679419
R53662 C8_N_btm.n249 C8_N_btm.n115 0.679419
R53663 C8_N_btm.n291 C8_N_btm.n290 0.679419
R53664 C8_N_btm.n300 C8_N_btm.n299 0.679419
R53665 C8_N_btm.n305 C8_N_btm.n304 0.679419
R53666 C8_N_btm.n320 C8_N_btm.n319 0.679419
R53667 C8_N_btm.n671 C8_N_btm.n670 0.679419
R53668 C8_N_btm.n755 C8_N_btm.n754 0.679419
R53669 C8_N_btm.n760 C8_N_btm.n758 0.679419
R53670 C8_N_btm.n773 C8_N_btm.n772 0.679419
R53671 C8_N_btm.n764 C8_N_btm.n763 0.679419
R53672 C8_N_btm.n786 C8_N_btm.n785 0.679419
R53673 C8_N_btm.n777 C8_N_btm.n776 0.679419
R53674 C8_N_btm.n49 C8_N_btm.n48 0.679419
R53675 C8_N_btm.n791 C8_N_btm.n789 0.679419
R53676 C8_N_btm.n795 C8_N_btm.n794 0.679419
R53677 C8_N_btm.n804 C8_N_btm.n803 0.679419
R53678 C8_N_btm.n808 C8_N_btm.n807 0.679419
R53679 C8_N_btm.n817 C8_N_btm.n816 0.679419
R53680 C8_N_btm.n822 C8_N_btm.n820 0.679419
R53681 C8_N_btm.n32 C8_N_btm.n31 0.679419
R53682 C8_N_btm.n835 C8_N_btm.n834 0.679419
R53683 C8_N_btm.n826 C8_N_btm.n825 0.679419
R53684 C8_N_btm.n859 C8_N_btm.n858 0.679419
R53685 C8_N_btm.n850 C8_N_btm.n849 0.679419
R53686 C8_N_btm.n846 C8_N_btm.n845 0.679419
R53687 C8_N_btm.n864 C8_N_btm.n862 0.679419
R53688 C8_N_btm.n868 C8_N_btm.n867 0.679419
R53689 C8_N_btm.n837 C8_N_btm.n17 0.679419
R53690 C8_N_btm.n879 C8_N_btm.n878 0.679419
R53691 C8_N_btm.n888 C8_N_btm.n887 0.679419
R53692 C8_N_btm.n892 C8_N_btm.n891 0.679419
R53693 C8_N_btm.n901 C8_N_btm.n900 0.679419
R53694 C8_N_btm.n80 C8_N_btm.n79 0.6255
R53695 C8_N_btm.n572 C8_N_btm.n571 0.6255
R53696 C8_N_btm.n569 C8_N_btm.n568 0.6255
R53697 C8_N_btm.n566 C8_N_btm.n565 0.6255
R53698 C8_N_btm.n563 C8_N_btm.n562 0.6255
R53699 C8_N_btm.n560 C8_N_btm.n559 0.6255
R53700 C8_N_btm.n557 C8_N_btm.n556 0.6255
R53701 C8_N_btm.n554 C8_N_btm.n553 0.6255
R53702 C8_N_btm.n551 C8_N_btm.n550 0.6255
R53703 C8_N_btm.n548 C8_N_btm.n547 0.6255
R53704 C8_N_btm.n545 C8_N_btm.n544 0.6255
R53705 C8_N_btm.n542 C8_N_btm.n541 0.6255
R53706 C8_N_btm.n539 C8_N_btm.n538 0.6255
R53707 C8_N_btm.n536 C8_N_btm.n535 0.6255
R53708 C8_N_btm.n533 C8_N_btm.n532 0.6255
R53709 C8_N_btm.n530 C8_N_btm.n529 0.6255
R53710 C8_N_btm.n527 C8_N_btm.n526 0.6255
R53711 C8_N_btm.n524 C8_N_btm.n523 0.6255
R53712 C8_N_btm.n521 C8_N_btm.n520 0.6255
R53713 C8_N_btm.n518 C8_N_btm.n517 0.6255
R53714 C8_N_btm.n515 C8_N_btm.n514 0.6255
R53715 C8_N_btm.n512 C8_N_btm.n511 0.6255
R53716 C8_N_btm.n509 C8_N_btm.n508 0.6255
R53717 C8_N_btm.n506 C8_N_btm.n505 0.6255
R53718 C8_N_btm.n503 C8_N_btm.n502 0.6255
R53719 C8_N_btm.n500 C8_N_btm.n499 0.6255
R53720 C8_N_btm.n497 C8_N_btm.n496 0.6255
R53721 C8_N_btm.n494 C8_N_btm.n493 0.6255
R53722 C8_N_btm.n487 C8_N_btm.n485 0.6255
R53723 C8_N_btm.n483 C8_N_btm.n482 0.6255
R53724 C8_N_btm.n480 C8_N_btm.n479 0.6255
R53725 C8_N_btm.n477 C8_N_btm.n476 0.6255
R53726 C8_N_btm.n474 C8_N_btm.n473 0.6255
R53727 C8_N_btm.n471 C8_N_btm.n470 0.6255
R53728 C8_N_btm.n468 C8_N_btm.n467 0.6255
R53729 C8_N_btm.n465 C8_N_btm.n464 0.6255
R53730 C8_N_btm.n462 C8_N_btm.n461 0.6255
R53731 C8_N_btm.n459 C8_N_btm.n458 0.6255
R53732 C8_N_btm.n456 C8_N_btm.n455 0.6255
R53733 C8_N_btm.n453 C8_N_btm.n452 0.6255
R53734 C8_N_btm.n450 C8_N_btm.n449 0.6255
R53735 C8_N_btm.n447 C8_N_btm.n446 0.6255
R53736 C8_N_btm.n444 C8_N_btm.n443 0.6255
R53737 C8_N_btm.n441 C8_N_btm.n440 0.6255
R53738 C8_N_btm.n438 C8_N_btm.n437 0.6255
R53739 C8_N_btm.n435 C8_N_btm.n434 0.6255
R53740 C8_N_btm.n432 C8_N_btm.n431 0.6255
R53741 C8_N_btm.n429 C8_N_btm.n428 0.6255
R53742 C8_N_btm.n426 C8_N_btm.n425 0.6255
R53743 C8_N_btm.n423 C8_N_btm.n422 0.6255
R53744 C8_N_btm.n420 C8_N_btm.n419 0.6255
R53745 C8_N_btm.n417 C8_N_btm.n416 0.6255
R53746 C8_N_btm.n414 C8_N_btm.n413 0.6255
R53747 C8_N_btm.n411 C8_N_btm.n410 0.6255
R53748 C8_N_btm.n408 C8_N_btm.n351 0.6255
R53749 C8_N_btm.n586 C8_N_btm.n585 0.6255
R53750 C8_N_btm.n589 C8_N_btm.n588 0.6255
R53751 C8_N_btm.n592 C8_N_btm.n591 0.6255
R53752 C8_N_btm.n595 C8_N_btm.n594 0.6255
R53753 C8_N_btm.n598 C8_N_btm.n597 0.6255
R53754 C8_N_btm.n601 C8_N_btm.n600 0.6255
R53755 C8_N_btm.n604 C8_N_btm.n603 0.6255
R53756 C8_N_btm.n607 C8_N_btm.n606 0.6255
R53757 C8_N_btm.n610 C8_N_btm.n609 0.6255
R53758 C8_N_btm.n613 C8_N_btm.n612 0.6255
R53759 C8_N_btm.n616 C8_N_btm.n615 0.6255
R53760 C8_N_btm.n619 C8_N_btm.n618 0.6255
R53761 C8_N_btm.n622 C8_N_btm.n621 0.6255
R53762 C8_N_btm.n625 C8_N_btm.n624 0.6255
R53763 C8_N_btm.n628 C8_N_btm.n627 0.6255
R53764 C8_N_btm.n631 C8_N_btm.n630 0.6255
R53765 C8_N_btm.n634 C8_N_btm.n633 0.6255
R53766 C8_N_btm.n637 C8_N_btm.n636 0.6255
R53767 C8_N_btm.n640 C8_N_btm.n639 0.6255
R53768 C8_N_btm.n643 C8_N_btm.n642 0.6255
R53769 C8_N_btm.n646 C8_N_btm.n645 0.6255
R53770 C8_N_btm.n649 C8_N_btm.n648 0.6255
R53771 C8_N_btm.n652 C8_N_btm.n651 0.6255
R53772 C8_N_btm.n655 C8_N_btm.n654 0.6255
R53773 C8_N_btm.n658 C8_N_btm.n657 0.6255
R53774 C8_N_btm.n661 C8_N_btm.n660 0.6255
R53775 C8_N_btm.n664 C8_N_btm.n663 0.6255
R53776 C8_N_btm.n168 C8_N_btm.n167 0.6255
R53777 C8_N_btm.n165 C8_N_btm.n164 0.6255
R53778 C8_N_btm.n182 C8_N_btm.n181 0.6255
R53779 C8_N_btm.n179 C8_N_btm.n178 0.6255
R53780 C8_N_btm.n195 C8_N_btm.n194 0.6255
R53781 C8_N_btm.n192 C8_N_btm.n191 0.6255
R53782 C8_N_btm.n153 C8_N_btm.n151 0.6255
R53783 C8_N_btm.n149 C8_N_btm.n143 0.6255
R53784 C8_N_btm.n210 C8_N_btm.n209 0.6255
R53785 C8_N_btm.n213 C8_N_btm.n212 0.6255
R53786 C8_N_btm.n223 C8_N_btm.n222 0.6255
R53787 C8_N_btm.n226 C8_N_btm.n225 0.6255
R53788 C8_N_btm.n132 C8_N_btm.n126 0.6255
R53789 C8_N_btm.n136 C8_N_btm.n134 0.6255
R53790 C8_N_btm.n244 C8_N_btm.n243 0.6255
R53791 C8_N_btm.n241 C8_N_btm.n240 0.6255
R53792 C8_N_btm.n268 C8_N_btm.n267 0.6255
R53793 C8_N_btm.n265 C8_N_btm.n264 0.6255
R53794 C8_N_btm.n255 C8_N_btm.n254 0.6255
R53795 C8_N_btm.n252 C8_N_btm.n118 0.6255
R53796 C8_N_btm.n283 C8_N_btm.n282 0.6255
R53797 C8_N_btm.n287 C8_N_btm.n285 0.6255
R53798 C8_N_btm.n294 C8_N_btm.n293 0.6255
R53799 C8_N_btm.n297 C8_N_btm.n296 0.6255
R53800 C8_N_btm.n308 C8_N_btm.n307 0.6255
R53801 C8_N_btm.n311 C8_N_btm.n310 0.6255
R53802 C8_N_btm.n314 C8_N_btm.n313 0.6255
R53803 C8_N_btm.n317 C8_N_btm.n316 0.6255
R53804 C8_N_btm.n674 C8_N_btm.n673 0.6255
R53805 C8_N_btm.n677 C8_N_btm.n676 0.6255
R53806 C8_N_btm.n680 C8_N_btm.n679 0.6255
R53807 C8_N_btm.n683 C8_N_btm.n682 0.6255
R53808 C8_N_btm.n686 C8_N_btm.n685 0.6255
R53809 C8_N_btm.n689 C8_N_btm.n688 0.6255
R53810 C8_N_btm.n692 C8_N_btm.n691 0.6255
R53811 C8_N_btm.n695 C8_N_btm.n694 0.6255
R53812 C8_N_btm.n698 C8_N_btm.n697 0.6255
R53813 C8_N_btm.n701 C8_N_btm.n700 0.6255
R53814 C8_N_btm.n704 C8_N_btm.n703 0.6255
R53815 C8_N_btm.n707 C8_N_btm.n706 0.6255
R53816 C8_N_btm.n710 C8_N_btm.n709 0.6255
R53817 C8_N_btm.n713 C8_N_btm.n712 0.6255
R53818 C8_N_btm.n716 C8_N_btm.n715 0.6255
R53819 C8_N_btm.n719 C8_N_btm.n718 0.6255
R53820 C8_N_btm.n722 C8_N_btm.n721 0.6255
R53821 C8_N_btm.n725 C8_N_btm.n724 0.6255
R53822 C8_N_btm.n728 C8_N_btm.n727 0.6255
R53823 C8_N_btm.n731 C8_N_btm.n730 0.6255
R53824 C8_N_btm.n734 C8_N_btm.n733 0.6255
R53825 C8_N_btm.n737 C8_N_btm.n736 0.6255
R53826 C8_N_btm.n740 C8_N_btm.n739 0.6255
R53827 C8_N_btm.n743 C8_N_btm.n742 0.6255
R53828 C8_N_btm.n746 C8_N_btm.n745 0.6255
R53829 C8_N_btm.n749 C8_N_btm.n748 0.6255
R53830 C8_N_btm.n752 C8_N_btm.n751 0.6255
R53831 C8_N_btm.n71 C8_N_btm.n62 0.6255
R53832 C8_N_btm.n74 C8_N_btm.n73 0.6255
R53833 C8_N_btm.n77 C8_N_btm.n76 0.6255
R53834 C8_N_btm.n770 C8_N_btm.n769 0.6255
R53835 C8_N_btm.n767 C8_N_btm.n766 0.6255
R53836 C8_N_btm.n783 C8_N_btm.n782 0.6255
R53837 C8_N_btm.n780 C8_N_btm.n779 0.6255
R53838 C8_N_btm.n55 C8_N_btm.n53 0.6255
R53839 C8_N_btm.n51 C8_N_btm.n45 0.6255
R53840 C8_N_btm.n798 C8_N_btm.n797 0.6255
R53841 C8_N_btm.n801 C8_N_btm.n800 0.6255
R53842 C8_N_btm.n811 C8_N_btm.n810 0.6255
R53843 C8_N_btm.n814 C8_N_btm.n813 0.6255
R53844 C8_N_btm.n34 C8_N_btm.n28 0.6255
R53845 C8_N_btm.n38 C8_N_btm.n36 0.6255
R53846 C8_N_btm.n832 C8_N_btm.n831 0.6255
R53847 C8_N_btm.n829 C8_N_btm.n828 0.6255
R53848 C8_N_btm.n856 C8_N_btm.n855 0.6255
R53849 C8_N_btm.n853 C8_N_btm.n852 0.6255
R53850 C8_N_btm.n843 C8_N_btm.n842 0.6255
R53851 C8_N_btm.n840 C8_N_btm.n20 0.6255
R53852 C8_N_btm.n871 C8_N_btm.n870 0.6255
R53853 C8_N_btm.n875 C8_N_btm.n873 0.6255
R53854 C8_N_btm.n882 C8_N_btm.n881 0.6255
R53855 C8_N_btm.n885 C8_N_btm.n884 0.6255
R53856 C8_N_btm.n895 C8_N_btm.n894 0.6255
R53857 C8_N_btm.n898 C8_N_btm.n897 0.6255
R53858 C8_N_btm.n82 C8_N_btm.n68 0.109875
R53859 C8_N_btm.n80 C8_N_btm.n68 0.109875
R53860 C8_N_btm.n572 C8_N_btm.n350 0.109875
R53861 C8_N_btm.n574 C8_N_btm.n350 0.109875
R53862 C8_N_btm.n569 C8_N_btm.n352 0.109875
R53863 C8_N_btm.n571 C8_N_btm.n352 0.109875
R53864 C8_N_btm.n566 C8_N_btm.n353 0.109875
R53865 C8_N_btm.n568 C8_N_btm.n353 0.109875
R53866 C8_N_btm.n563 C8_N_btm.n354 0.109875
R53867 C8_N_btm.n565 C8_N_btm.n354 0.109875
R53868 C8_N_btm.n560 C8_N_btm.n355 0.109875
R53869 C8_N_btm.n562 C8_N_btm.n355 0.109875
R53870 C8_N_btm.n557 C8_N_btm.n356 0.109875
R53871 C8_N_btm.n559 C8_N_btm.n356 0.109875
R53872 C8_N_btm.n554 C8_N_btm.n357 0.109875
R53873 C8_N_btm.n556 C8_N_btm.n357 0.109875
R53874 C8_N_btm.n551 C8_N_btm.n358 0.109875
R53875 C8_N_btm.n553 C8_N_btm.n358 0.109875
R53876 C8_N_btm.n548 C8_N_btm.n359 0.109875
R53877 C8_N_btm.n550 C8_N_btm.n359 0.109875
R53878 C8_N_btm.n545 C8_N_btm.n360 0.109875
R53879 C8_N_btm.n547 C8_N_btm.n360 0.109875
R53880 C8_N_btm.n542 C8_N_btm.n361 0.109875
R53881 C8_N_btm.n544 C8_N_btm.n361 0.109875
R53882 C8_N_btm.n539 C8_N_btm.n362 0.109875
R53883 C8_N_btm.n541 C8_N_btm.n362 0.109875
R53884 C8_N_btm.n536 C8_N_btm.n363 0.109875
R53885 C8_N_btm.n538 C8_N_btm.n363 0.109875
R53886 C8_N_btm.n533 C8_N_btm.n364 0.109875
R53887 C8_N_btm.n535 C8_N_btm.n364 0.109875
R53888 C8_N_btm.n530 C8_N_btm.n367 0.109875
R53889 C8_N_btm.n532 C8_N_btm.n367 0.109875
R53890 C8_N_btm.n527 C8_N_btm.n368 0.109875
R53891 C8_N_btm.n529 C8_N_btm.n368 0.109875
R53892 C8_N_btm.n524 C8_N_btm.n369 0.109875
R53893 C8_N_btm.n526 C8_N_btm.n369 0.109875
R53894 C8_N_btm.n521 C8_N_btm.n370 0.109875
R53895 C8_N_btm.n523 C8_N_btm.n370 0.109875
R53896 C8_N_btm.n518 C8_N_btm.n371 0.109875
R53897 C8_N_btm.n520 C8_N_btm.n371 0.109875
R53898 C8_N_btm.n515 C8_N_btm.n372 0.109875
R53899 C8_N_btm.n517 C8_N_btm.n372 0.109875
R53900 C8_N_btm.n512 C8_N_btm.n373 0.109875
R53901 C8_N_btm.n514 C8_N_btm.n373 0.109875
R53902 C8_N_btm.n509 C8_N_btm.n374 0.109875
R53903 C8_N_btm.n511 C8_N_btm.n374 0.109875
R53904 C8_N_btm.n506 C8_N_btm.n375 0.109875
R53905 C8_N_btm.n508 C8_N_btm.n375 0.109875
R53906 C8_N_btm.n503 C8_N_btm.n376 0.109875
R53907 C8_N_btm.n505 C8_N_btm.n376 0.109875
R53908 C8_N_btm.n500 C8_N_btm.n377 0.109875
R53909 C8_N_btm.n502 C8_N_btm.n377 0.109875
R53910 C8_N_btm.n497 C8_N_btm.n378 0.109875
R53911 C8_N_btm.n499 C8_N_btm.n378 0.109875
R53912 C8_N_btm.n494 C8_N_btm.n379 0.109875
R53913 C8_N_btm.n496 C8_N_btm.n379 0.109875
R53914 C8_N_btm.n491 C8_N_btm.n489 0.109875
R53915 C8_N_btm.n493 C8_N_btm.n489 0.109875
R53916 C8_N_btm.n488 C8_N_btm.n381 0.109875
R53917 C8_N_btm.n488 C8_N_btm.n487 0.109875
R53918 C8_N_btm.n485 C8_N_btm.n382 0.109875
R53919 C8_N_btm.n483 C8_N_btm.n382 0.109875
R53920 C8_N_btm.n482 C8_N_btm.n383 0.109875
R53921 C8_N_btm.n480 C8_N_btm.n383 0.109875
R53922 C8_N_btm.n479 C8_N_btm.n384 0.109875
R53923 C8_N_btm.n477 C8_N_btm.n384 0.109875
R53924 C8_N_btm.n476 C8_N_btm.n385 0.109875
R53925 C8_N_btm.n474 C8_N_btm.n385 0.109875
R53926 C8_N_btm.n473 C8_N_btm.n386 0.109875
R53927 C8_N_btm.n471 C8_N_btm.n386 0.109875
R53928 C8_N_btm.n470 C8_N_btm.n387 0.109875
R53929 C8_N_btm.n468 C8_N_btm.n387 0.109875
R53930 C8_N_btm.n467 C8_N_btm.n388 0.109875
R53931 C8_N_btm.n465 C8_N_btm.n388 0.109875
R53932 C8_N_btm.n464 C8_N_btm.n389 0.109875
R53933 C8_N_btm.n462 C8_N_btm.n389 0.109875
R53934 C8_N_btm.n461 C8_N_btm.n390 0.109875
R53935 C8_N_btm.n459 C8_N_btm.n390 0.109875
R53936 C8_N_btm.n458 C8_N_btm.n391 0.109875
R53937 C8_N_btm.n456 C8_N_btm.n391 0.109875
R53938 C8_N_btm.n455 C8_N_btm.n392 0.109875
R53939 C8_N_btm.n453 C8_N_btm.n392 0.109875
R53940 C8_N_btm.n452 C8_N_btm.n393 0.109875
R53941 C8_N_btm.n450 C8_N_btm.n393 0.109875
R53942 C8_N_btm.n449 C8_N_btm.n394 0.109875
R53943 C8_N_btm.n447 C8_N_btm.n394 0.109875
R53944 C8_N_btm.n446 C8_N_btm.n395 0.109875
R53945 C8_N_btm.n444 C8_N_btm.n395 0.109875
R53946 C8_N_btm.n443 C8_N_btm.n396 0.109875
R53947 C8_N_btm.n441 C8_N_btm.n396 0.109875
R53948 C8_N_btm.n440 C8_N_btm.n397 0.109875
R53949 C8_N_btm.n438 C8_N_btm.n397 0.109875
R53950 C8_N_btm.n437 C8_N_btm.n398 0.109875
R53951 C8_N_btm.n435 C8_N_btm.n398 0.109875
R53952 C8_N_btm.n434 C8_N_btm.n399 0.109875
R53953 C8_N_btm.n432 C8_N_btm.n399 0.109875
R53954 C8_N_btm.n431 C8_N_btm.n400 0.109875
R53955 C8_N_btm.n429 C8_N_btm.n400 0.109875
R53956 C8_N_btm.n428 C8_N_btm.n401 0.109875
R53957 C8_N_btm.n426 C8_N_btm.n401 0.109875
R53958 C8_N_btm.n425 C8_N_btm.n402 0.109875
R53959 C8_N_btm.n423 C8_N_btm.n402 0.109875
R53960 C8_N_btm.n422 C8_N_btm.n403 0.109875
R53961 C8_N_btm.n420 C8_N_btm.n403 0.109875
R53962 C8_N_btm.n419 C8_N_btm.n404 0.109875
R53963 C8_N_btm.n417 C8_N_btm.n404 0.109875
R53964 C8_N_btm.n416 C8_N_btm.n405 0.109875
R53965 C8_N_btm.n414 C8_N_btm.n405 0.109875
R53966 C8_N_btm.n413 C8_N_btm.n406 0.109875
R53967 C8_N_btm.n411 C8_N_btm.n406 0.109875
R53968 C8_N_btm.n410 C8_N_btm.n407 0.109875
R53969 C8_N_btm.n408 C8_N_btm.n407 0.109875
R53970 C8_N_btm.n580 C8_N_btm.n351 0.109875
R53971 C8_N_btm.n580 C8_N_btm.n579 0.109875
R53972 C8_N_btm.n585 C8_N_btm.n581 0.109875
R53973 C8_N_btm.n583 C8_N_btm.n581 0.109875
R53974 C8_N_btm.n588 C8_N_btm.n349 0.109875
R53975 C8_N_btm.n586 C8_N_btm.n349 0.109875
R53976 C8_N_btm.n591 C8_N_btm.n348 0.109875
R53977 C8_N_btm.n589 C8_N_btm.n348 0.109875
R53978 C8_N_btm.n594 C8_N_btm.n347 0.109875
R53979 C8_N_btm.n592 C8_N_btm.n347 0.109875
R53980 C8_N_btm.n597 C8_N_btm.n346 0.109875
R53981 C8_N_btm.n595 C8_N_btm.n346 0.109875
R53982 C8_N_btm.n600 C8_N_btm.n345 0.109875
R53983 C8_N_btm.n598 C8_N_btm.n345 0.109875
R53984 C8_N_btm.n603 C8_N_btm.n344 0.109875
R53985 C8_N_btm.n601 C8_N_btm.n344 0.109875
R53986 C8_N_btm.n606 C8_N_btm.n343 0.109875
R53987 C8_N_btm.n604 C8_N_btm.n343 0.109875
R53988 C8_N_btm.n609 C8_N_btm.n342 0.109875
R53989 C8_N_btm.n607 C8_N_btm.n342 0.109875
R53990 C8_N_btm.n612 C8_N_btm.n341 0.109875
R53991 C8_N_btm.n610 C8_N_btm.n341 0.109875
R53992 C8_N_btm.n615 C8_N_btm.n340 0.109875
R53993 C8_N_btm.n613 C8_N_btm.n340 0.109875
R53994 C8_N_btm.n618 C8_N_btm.n339 0.109875
R53995 C8_N_btm.n616 C8_N_btm.n339 0.109875
R53996 C8_N_btm.n621 C8_N_btm.n338 0.109875
R53997 C8_N_btm.n619 C8_N_btm.n338 0.109875
R53998 C8_N_btm.n624 C8_N_btm.n337 0.109875
R53999 C8_N_btm.n622 C8_N_btm.n337 0.109875
R54000 C8_N_btm.n627 C8_N_btm.n336 0.109875
R54001 C8_N_btm.n625 C8_N_btm.n336 0.109875
R54002 C8_N_btm.n630 C8_N_btm.n335 0.109875
R54003 C8_N_btm.n628 C8_N_btm.n335 0.109875
R54004 C8_N_btm.n633 C8_N_btm.n334 0.109875
R54005 C8_N_btm.n631 C8_N_btm.n334 0.109875
R54006 C8_N_btm.n636 C8_N_btm.n333 0.109875
R54007 C8_N_btm.n634 C8_N_btm.n333 0.109875
R54008 C8_N_btm.n639 C8_N_btm.n332 0.109875
R54009 C8_N_btm.n637 C8_N_btm.n332 0.109875
R54010 C8_N_btm.n642 C8_N_btm.n331 0.109875
R54011 C8_N_btm.n640 C8_N_btm.n331 0.109875
R54012 C8_N_btm.n645 C8_N_btm.n330 0.109875
R54013 C8_N_btm.n643 C8_N_btm.n330 0.109875
R54014 C8_N_btm.n648 C8_N_btm.n329 0.109875
R54015 C8_N_btm.n646 C8_N_btm.n329 0.109875
R54016 C8_N_btm.n651 C8_N_btm.n328 0.109875
R54017 C8_N_btm.n649 C8_N_btm.n328 0.109875
R54018 C8_N_btm.n654 C8_N_btm.n327 0.109875
R54019 C8_N_btm.n652 C8_N_btm.n327 0.109875
R54020 C8_N_btm.n657 C8_N_btm.n326 0.109875
R54021 C8_N_btm.n655 C8_N_btm.n326 0.109875
R54022 C8_N_btm.n660 C8_N_btm.n325 0.109875
R54023 C8_N_btm.n658 C8_N_btm.n325 0.109875
R54024 C8_N_btm.n663 C8_N_btm.n324 0.109875
R54025 C8_N_btm.n661 C8_N_btm.n324 0.109875
R54026 C8_N_btm.n666 C8_N_btm.n323 0.109875
R54027 C8_N_btm.n664 C8_N_btm.n323 0.109875
R54028 C8_N_btm.n173 C8_N_btm.n168 0.109875
R54029 C8_N_btm.n173 C8_N_btm.n172 0.109875
R54030 C8_N_btm.n165 C8_N_btm.n159 0.109875
R54031 C8_N_btm.n167 C8_N_btm.n159 0.109875
R54032 C8_N_btm.n162 C8_N_btm.n160 0.109875
R54033 C8_N_btm.n164 C8_N_btm.n160 0.109875
R54034 C8_N_btm.n184 C8_N_btm.n157 0.109875
R54035 C8_N_btm.n182 C8_N_btm.n157 0.109875
R54036 C8_N_btm.n181 C8_N_btm.n158 0.109875
R54037 C8_N_btm.n179 C8_N_btm.n158 0.109875
R54038 C8_N_btm.n178 C8_N_btm.n174 0.109875
R54039 C8_N_btm.n176 C8_N_btm.n174 0.109875
R54040 C8_N_btm.n195 C8_N_btm.n142 0.109875
R54041 C8_N_btm.n197 C8_N_btm.n142 0.109875
R54042 C8_N_btm.n192 C8_N_btm.n145 0.109875
R54043 C8_N_btm.n194 C8_N_btm.n145 0.109875
R54044 C8_N_btm.n189 C8_N_btm.n155 0.109875
R54045 C8_N_btm.n191 C8_N_btm.n155 0.109875
R54046 C8_N_btm.n154 C8_N_btm.n147 0.109875
R54047 C8_N_btm.n154 C8_N_btm.n153 0.109875
R54048 C8_N_btm.n151 C8_N_btm.n148 0.109875
R54049 C8_N_btm.n149 C8_N_btm.n148 0.109875
R54050 C8_N_btm.n204 C8_N_btm.n143 0.109875
R54051 C8_N_btm.n204 C8_N_btm.n203 0.109875
R54052 C8_N_btm.n209 C8_N_btm.n205 0.109875
R54053 C8_N_btm.n207 C8_N_btm.n205 0.109875
R54054 C8_N_btm.n212 C8_N_btm.n141 0.109875
R54055 C8_N_btm.n210 C8_N_btm.n141 0.109875
R54056 C8_N_btm.n215 C8_N_btm.n140 0.109875
R54057 C8_N_btm.n213 C8_N_btm.n140 0.109875
R54058 C8_N_btm.n220 C8_N_btm.n138 0.109875
R54059 C8_N_btm.n222 C8_N_btm.n138 0.109875
R54060 C8_N_btm.n223 C8_N_btm.n128 0.109875
R54061 C8_N_btm.n225 C8_N_btm.n128 0.109875
R54062 C8_N_btm.n226 C8_N_btm.n125 0.109875
R54063 C8_N_btm.n228 C8_N_btm.n125 0.109875
R54064 C8_N_btm.n235 C8_N_btm.n126 0.109875
R54065 C8_N_btm.n235 C8_N_btm.n234 0.109875
R54066 C8_N_btm.n134 C8_N_btm.n131 0.109875
R54067 C8_N_btm.n132 C8_N_btm.n131 0.109875
R54068 C8_N_btm.n137 C8_N_btm.n130 0.109875
R54069 C8_N_btm.n137 C8_N_btm.n136 0.109875
R54070 C8_N_btm.n246 C8_N_btm.n123 0.109875
R54071 C8_N_btm.n244 C8_N_btm.n123 0.109875
R54072 C8_N_btm.n243 C8_N_btm.n124 0.109875
R54073 C8_N_btm.n241 C8_N_btm.n124 0.109875
R54074 C8_N_btm.n240 C8_N_btm.n236 0.109875
R54075 C8_N_btm.n238 C8_N_btm.n236 0.109875
R54076 C8_N_btm.n268 C8_N_btm.n117 0.109875
R54077 C8_N_btm.n270 C8_N_btm.n117 0.109875
R54078 C8_N_btm.n265 C8_N_btm.n120 0.109875
R54079 C8_N_btm.n267 C8_N_btm.n120 0.109875
R54080 C8_N_btm.n262 C8_N_btm.n121 0.109875
R54081 C8_N_btm.n264 C8_N_btm.n121 0.109875
R54082 C8_N_btm.n257 C8_N_btm.n114 0.109875
R54083 C8_N_btm.n255 C8_N_btm.n114 0.109875
R54084 C8_N_btm.n254 C8_N_btm.n251 0.109875
R54085 C8_N_btm.n252 C8_N_btm.n251 0.109875
R54086 C8_N_btm.n277 C8_N_btm.n118 0.109875
R54087 C8_N_btm.n277 C8_N_btm.n276 0.109875
R54088 C8_N_btm.n282 C8_N_btm.n278 0.109875
R54089 C8_N_btm.n280 C8_N_btm.n278 0.109875
R54090 C8_N_btm.n285 C8_N_btm.n116 0.109875
R54091 C8_N_btm.n283 C8_N_btm.n116 0.109875
R54092 C8_N_btm.n288 C8_N_btm.n115 0.109875
R54093 C8_N_btm.n288 C8_N_btm.n287 0.109875
R54094 C8_N_btm.n291 C8_N_btm.n289 0.109875
R54095 C8_N_btm.n293 C8_N_btm.n289 0.109875
R54096 C8_N_btm.n294 C8_N_btm.n113 0.109875
R54097 C8_N_btm.n296 C8_N_btm.n113 0.109875
R54098 C8_N_btm.n297 C8_N_btm.n112 0.109875
R54099 C8_N_btm.n299 C8_N_btm.n112 0.109875
R54100 C8_N_btm.n307 C8_N_btm.n303 0.109875
R54101 C8_N_btm.n305 C8_N_btm.n303 0.109875
R54102 C8_N_btm.n310 C8_N_btm.n302 0.109875
R54103 C8_N_btm.n308 C8_N_btm.n302 0.109875
R54104 C8_N_btm.n313 C8_N_btm.n110 0.109875
R54105 C8_N_btm.n311 C8_N_btm.n110 0.109875
R54106 C8_N_btm.n316 C8_N_btm.n109 0.109875
R54107 C8_N_btm.n314 C8_N_btm.n109 0.109875
R54108 C8_N_btm.n319 C8_N_btm.n108 0.109875
R54109 C8_N_btm.n317 C8_N_btm.n108 0.109875
R54110 C8_N_btm.n671 C8_N_btm.n106 0.109875
R54111 C8_N_btm.n673 C8_N_btm.n106 0.109875
R54112 C8_N_btm.n674 C8_N_btm.n105 0.109875
R54113 C8_N_btm.n676 C8_N_btm.n105 0.109875
R54114 C8_N_btm.n677 C8_N_btm.n104 0.109875
R54115 C8_N_btm.n679 C8_N_btm.n104 0.109875
R54116 C8_N_btm.n680 C8_N_btm.n103 0.109875
R54117 C8_N_btm.n682 C8_N_btm.n103 0.109875
R54118 C8_N_btm.n683 C8_N_btm.n102 0.109875
R54119 C8_N_btm.n685 C8_N_btm.n102 0.109875
R54120 C8_N_btm.n686 C8_N_btm.n101 0.109875
R54121 C8_N_btm.n688 C8_N_btm.n101 0.109875
R54122 C8_N_btm.n689 C8_N_btm.n100 0.109875
R54123 C8_N_btm.n691 C8_N_btm.n100 0.109875
R54124 C8_N_btm.n692 C8_N_btm.n99 0.109875
R54125 C8_N_btm.n694 C8_N_btm.n99 0.109875
R54126 C8_N_btm.n695 C8_N_btm.n98 0.109875
R54127 C8_N_btm.n697 C8_N_btm.n98 0.109875
R54128 C8_N_btm.n698 C8_N_btm.n97 0.109875
R54129 C8_N_btm.n700 C8_N_btm.n97 0.109875
R54130 C8_N_btm.n701 C8_N_btm.n96 0.109875
R54131 C8_N_btm.n703 C8_N_btm.n96 0.109875
R54132 C8_N_btm.n704 C8_N_btm.n95 0.109875
R54133 C8_N_btm.n706 C8_N_btm.n95 0.109875
R54134 C8_N_btm.n707 C8_N_btm.n94 0.109875
R54135 C8_N_btm.n709 C8_N_btm.n94 0.109875
R54136 C8_N_btm.n710 C8_N_btm.n93 0.109875
R54137 C8_N_btm.n712 C8_N_btm.n93 0.109875
R54138 C8_N_btm.n713 C8_N_btm.n92 0.109875
R54139 C8_N_btm.n715 C8_N_btm.n92 0.109875
R54140 C8_N_btm.n716 C8_N_btm.n91 0.109875
R54141 C8_N_btm.n718 C8_N_btm.n91 0.109875
R54142 C8_N_btm.n719 C8_N_btm.n90 0.109875
R54143 C8_N_btm.n721 C8_N_btm.n90 0.109875
R54144 C8_N_btm.n722 C8_N_btm.n89 0.109875
R54145 C8_N_btm.n724 C8_N_btm.n89 0.109875
R54146 C8_N_btm.n725 C8_N_btm.n88 0.109875
R54147 C8_N_btm.n727 C8_N_btm.n88 0.109875
R54148 C8_N_btm.n728 C8_N_btm.n87 0.109875
R54149 C8_N_btm.n730 C8_N_btm.n87 0.109875
R54150 C8_N_btm.n731 C8_N_btm.n86 0.109875
R54151 C8_N_btm.n733 C8_N_btm.n86 0.109875
R54152 C8_N_btm.n734 C8_N_btm.n85 0.109875
R54153 C8_N_btm.n736 C8_N_btm.n85 0.109875
R54154 C8_N_btm.n737 C8_N_btm.n84 0.109875
R54155 C8_N_btm.n739 C8_N_btm.n84 0.109875
R54156 C8_N_btm.n740 C8_N_btm.n67 0.109875
R54157 C8_N_btm.n742 C8_N_btm.n67 0.109875
R54158 C8_N_btm.n743 C8_N_btm.n66 0.109875
R54159 C8_N_btm.n745 C8_N_btm.n66 0.109875
R54160 C8_N_btm.n746 C8_N_btm.n65 0.109875
R54161 C8_N_btm.n748 C8_N_btm.n65 0.109875
R54162 C8_N_btm.n749 C8_N_btm.n64 0.109875
R54163 C8_N_btm.n751 C8_N_btm.n64 0.109875
R54164 C8_N_btm.n752 C8_N_btm.n61 0.109875
R54165 C8_N_btm.n754 C8_N_btm.n61 0.109875
R54166 C8_N_btm.n761 C8_N_btm.n62 0.109875
R54167 C8_N_btm.n761 C8_N_btm.n760 0.109875
R54168 C8_N_btm.n73 C8_N_btm.n70 0.109875
R54169 C8_N_btm.n71 C8_N_btm.n70 0.109875
R54170 C8_N_btm.n76 C8_N_btm.n69 0.109875
R54171 C8_N_btm.n74 C8_N_btm.n69 0.109875
R54172 C8_N_btm.n79 C8_N_btm.n58 0.109875
R54173 C8_N_btm.n77 C8_N_btm.n58 0.109875
R54174 C8_N_btm.n772 C8_N_btm.n59 0.109875
R54175 C8_N_btm.n770 C8_N_btm.n59 0.109875
R54176 C8_N_btm.n769 C8_N_btm.n60 0.109875
R54177 C8_N_btm.n767 C8_N_btm.n60 0.109875
R54178 C8_N_btm.n766 C8_N_btm.n762 0.109875
R54179 C8_N_btm.n764 C8_N_btm.n762 0.109875
R54180 C8_N_btm.n783 C8_N_btm.n44 0.109875
R54181 C8_N_btm.n785 C8_N_btm.n44 0.109875
R54182 C8_N_btm.n780 C8_N_btm.n47 0.109875
R54183 C8_N_btm.n782 C8_N_btm.n47 0.109875
R54184 C8_N_btm.n777 C8_N_btm.n57 0.109875
R54185 C8_N_btm.n779 C8_N_btm.n57 0.109875
R54186 C8_N_btm.n56 C8_N_btm.n49 0.109875
R54187 C8_N_btm.n56 C8_N_btm.n55 0.109875
R54188 C8_N_btm.n53 C8_N_btm.n50 0.109875
R54189 C8_N_btm.n51 C8_N_btm.n50 0.109875
R54190 C8_N_btm.n792 C8_N_btm.n45 0.109875
R54191 C8_N_btm.n792 C8_N_btm.n791 0.109875
R54192 C8_N_btm.n797 C8_N_btm.n793 0.109875
R54193 C8_N_btm.n795 C8_N_btm.n793 0.109875
R54194 C8_N_btm.n800 C8_N_btm.n43 0.109875
R54195 C8_N_btm.n798 C8_N_btm.n43 0.109875
R54196 C8_N_btm.n803 C8_N_btm.n42 0.109875
R54197 C8_N_btm.n801 C8_N_btm.n42 0.109875
R54198 C8_N_btm.n808 C8_N_btm.n40 0.109875
R54199 C8_N_btm.n810 C8_N_btm.n40 0.109875
R54200 C8_N_btm.n811 C8_N_btm.n30 0.109875
R54201 C8_N_btm.n813 C8_N_btm.n30 0.109875
R54202 C8_N_btm.n814 C8_N_btm.n27 0.109875
R54203 C8_N_btm.n816 C8_N_btm.n27 0.109875
R54204 C8_N_btm.n823 C8_N_btm.n28 0.109875
R54205 C8_N_btm.n823 C8_N_btm.n822 0.109875
R54206 C8_N_btm.n36 C8_N_btm.n33 0.109875
R54207 C8_N_btm.n34 C8_N_btm.n33 0.109875
R54208 C8_N_btm.n39 C8_N_btm.n32 0.109875
R54209 C8_N_btm.n39 C8_N_btm.n38 0.109875
R54210 C8_N_btm.n834 C8_N_btm.n25 0.109875
R54211 C8_N_btm.n832 C8_N_btm.n25 0.109875
R54212 C8_N_btm.n831 C8_N_btm.n26 0.109875
R54213 C8_N_btm.n829 C8_N_btm.n26 0.109875
R54214 C8_N_btm.n828 C8_N_btm.n824 0.109875
R54215 C8_N_btm.n826 C8_N_btm.n824 0.109875
R54216 C8_N_btm.n856 C8_N_btm.n19 0.109875
R54217 C8_N_btm.n858 C8_N_btm.n19 0.109875
R54218 C8_N_btm.n853 C8_N_btm.n22 0.109875
R54219 C8_N_btm.n855 C8_N_btm.n22 0.109875
R54220 C8_N_btm.n850 C8_N_btm.n23 0.109875
R54221 C8_N_btm.n852 C8_N_btm.n23 0.109875
R54222 C8_N_btm.n845 C8_N_btm.n16 0.109875
R54223 C8_N_btm.n843 C8_N_btm.n16 0.109875
R54224 C8_N_btm.n842 C8_N_btm.n839 0.109875
R54225 C8_N_btm.n840 C8_N_btm.n839 0.109875
R54226 C8_N_btm.n865 C8_N_btm.n20 0.109875
R54227 C8_N_btm.n865 C8_N_btm.n864 0.109875
R54228 C8_N_btm.n870 C8_N_btm.n866 0.109875
R54229 C8_N_btm.n868 C8_N_btm.n866 0.109875
R54230 C8_N_btm.n873 C8_N_btm.n18 0.109875
R54231 C8_N_btm.n871 C8_N_btm.n18 0.109875
R54232 C8_N_btm.n876 C8_N_btm.n17 0.109875
R54233 C8_N_btm.n876 C8_N_btm.n875 0.109875
R54234 C8_N_btm.n879 C8_N_btm.n877 0.109875
R54235 C8_N_btm.n881 C8_N_btm.n877 0.109875
R54236 C8_N_btm.n882 C8_N_btm.n15 0.109875
R54237 C8_N_btm.n884 C8_N_btm.n15 0.109875
R54238 C8_N_btm.n885 C8_N_btm.n14 0.109875
R54239 C8_N_btm.n887 C8_N_btm.n14 0.109875
R54240 C8_N_btm.n894 C8_N_btm.n12 0.109875
R54241 C8_N_btm.n892 C8_N_btm.n12 0.109875
R54242 C8_N_btm.n897 C8_N_btm.n11 0.109875
R54243 C8_N_btm.n895 C8_N_btm.n11 0.109875
R54244 C8_N_btm.n900 C8_N_btm.n10 0.109875
R54245 C8_N_btm.n898 C8_N_btm.n10 0.109875
R54246 C8_N_btm.n380 C8_N_btm.n322 0.0556875
R54247 C8_N_btm.n577 C8_N_btm.n576 0.0556875
R54248 C8_N_btm.n582 C8_N_btm.n63 0.0556875
R54249 C8_N_btm.n668 C8_N_btm.n667 0.0556875
R54250 C8_N_btm.n170 C8_N_btm.n169 0.0556875
R54251 C8_N_btm.n161 C8_N_btm.n156 0.0556875
R54252 C8_N_btm.n186 C8_N_btm.n185 0.0556875
R54253 C8_N_btm.n175 C8_N_btm.n144 0.0556875
R54254 C8_N_btm.n199 C8_N_btm.n198 0.0556875
R54255 C8_N_btm.n188 C8_N_btm.n187 0.0556875
R54256 C8_N_btm.n146 C8_N_btm.n139 0.0556875
R54257 C8_N_btm.n201 C8_N_btm.n200 0.0556875
R54258 C8_N_btm.n206 C8_N_btm.n127 0.0556875
R54259 C8_N_btm.n217 C8_N_btm.n216 0.0556875
R54260 C8_N_btm.n219 C8_N_btm.n218 0.0556875
R54261 C8_N_btm.n230 C8_N_btm.n229 0.0556875
R54262 C8_N_btm.n232 C8_N_btm.n231 0.0556875
R54263 C8_N_btm.n129 C8_N_btm.n122 0.0556875
R54264 C8_N_btm.n248 C8_N_btm.n247 0.0556875
R54265 C8_N_btm.n237 C8_N_btm.n119 0.0556875
R54266 C8_N_btm.n272 C8_N_btm.n271 0.0556875
R54267 C8_N_btm.n261 C8_N_btm.n260 0.0556875
R54268 C8_N_btm.n259 C8_N_btm.n258 0.0556875
R54269 C8_N_btm.n274 C8_N_btm.n273 0.0556875
R54270 C8_N_btm.n279 C8_N_btm.n111 0.0556875
R54271 C8_N_btm.n250 C8_N_btm.n249 0.0556875
R54272 C8_N_btm.n290 C8_N_btm.n107 0.0556875
R54273 C8_N_btm.n301 C8_N_btm.n300 0.0556875
R54274 C8_N_btm.n321 C8_N_btm.n320 0.0556875
R54275 C8_N_btm.n670 C8_N_btm.n669 0.0556875
R54276 C8_N_btm.n756 C8_N_btm.n755 0.0556875
R54277 C8_N_btm.n758 C8_N_btm.n757 0.0556875
R54278 C8_N_btm.n774 C8_N_btm.n773 0.0556875
R54279 C8_N_btm.n763 C8_N_btm.n46 0.0556875
R54280 C8_N_btm.n787 C8_N_btm.n786 0.0556875
R54281 C8_N_btm.n776 C8_N_btm.n775 0.0556875
R54282 C8_N_btm.n48 C8_N_btm.n41 0.0556875
R54283 C8_N_btm.n789 C8_N_btm.n788 0.0556875
R54284 C8_N_btm.n794 C8_N_btm.n29 0.0556875
R54285 C8_N_btm.n805 C8_N_btm.n804 0.0556875
R54286 C8_N_btm.n807 C8_N_btm.n806 0.0556875
R54287 C8_N_btm.n818 C8_N_btm.n817 0.0556875
R54288 C8_N_btm.n820 C8_N_btm.n819 0.0556875
R54289 C8_N_btm.n31 C8_N_btm.n24 0.0556875
R54290 C8_N_btm.n836 C8_N_btm.n835 0.0556875
R54291 C8_N_btm.n825 C8_N_btm.n21 0.0556875
R54292 C8_N_btm.n860 C8_N_btm.n859 0.0556875
R54293 C8_N_btm.n849 C8_N_btm.n848 0.0556875
R54294 C8_N_btm.n847 C8_N_btm.n846 0.0556875
R54295 C8_N_btm.n862 C8_N_btm.n861 0.0556875
R54296 C8_N_btm.n867 C8_N_btm.n13 0.0556875
R54297 C8_N_btm.n838 C8_N_btm.n837 0.0556875
R54298 C8_N_btm.n878 C8_N_btm.n9 0.0556875
R54299 C8_N_btm.n889 C8_N_btm.n888 0.0556875
R54300 C8_N_btm.n891 C8_N_btm.n890 0.0556875
R54301 C8_N_btm.n902 C8_N_btm.n901 0.0556875
R54302 a_13273_44868.n8 a_13273_44868.t23 330.12
R54303 a_13273_44868.n6 a_13273_44868.t27 256.726
R54304 a_13273_44868.n2 a_13273_44868.n0 248.087
R54305 a_13273_44868.n19 a_13273_44868.t22 238.397
R54306 a_13273_44868.n3 a_13273_44868.t10 231.835
R54307 a_13273_44868.n15 a_13273_44868.t13 231.017
R54308 a_13273_44868.n13 a_13273_44868.t12 231.017
R54309 a_13273_44868.n20 a_13273_44868.t19 221.72
R54310 a_13273_44868.n21 a_13273_44868.t29 221.72
R54311 a_13273_44868.n4 a_13273_44868.t17 212.081
R54312 a_13273_44868.n5 a_13273_44868.t9 212.081
R54313 a_13273_44868.n2 a_13273_44868.n1 208.507
R54314 a_13273_44868.n17 a_13273_44868.n5 207.501
R54315 a_13273_44868.n8 a_13273_44868.t14 201.587
R54316 a_13273_44868.n19 a_13273_44868.t28 195.017
R54317 a_13273_44868.n23 a_13273_44868.n22 190.44
R54318 a_13273_44868.n23 a_13273_44868.n19 184.151
R54319 a_13273_44868.n7 a_13273_44868.t16 183.505
R54320 a_13273_44868.n9 a_13273_44868.n7 181.725
R54321 a_13273_44868.n12 a_13273_44868.n6 178.672
R54322 a_13273_44868.n14 a_13273_44868.n13 176.94
R54323 a_13273_44868.n18 a_13273_44868.n3 171.261
R54324 a_13273_44868.n9 a_13273_44868.n8 166.133
R54325 a_13273_44868.n16 a_13273_44868.n15 163.046
R54326 a_13273_44868.n11 a_13273_44868.n10 163.024
R54327 a_13273_44868.n6 a_13273_44868.t21 161.275
R54328 a_13273_44868.n15 a_13273_44868.t18 158.716
R54329 a_13273_44868.n13 a_13273_44868.t31 158.716
R54330 a_13273_44868.n3 a_13273_44868.t26 157.07
R54331 a_13273_44868.n20 a_13273_44868.t8 149.421
R54332 a_13273_44868.n21 a_13273_44868.t24 149.421
R54333 a_13273_44868.n4 a_13273_44868.t15 139.78
R54334 a_13273_44868.n5 a_13273_44868.t25 139.78
R54335 a_13273_44868.n28 a_13273_44868.n27 137.576
R54336 a_13273_44868.n10 a_13273_44868.t20 137.177
R54337 a_13273_44868.n10 a_13273_44868.t11 121.109
R54338 a_13273_44868.n7 a_13273_44868.t30 114.532
R54339 a_13273_44868.n27 a_13273_44868.n26 99.1759
R54340 a_13273_44868.n5 a_13273_44868.n4 62.8066
R54341 a_13273_44868.n22 a_13273_44868.n20 37.4894
R54342 a_13273_44868.n22 a_13273_44868.n21 37.4894
R54343 a_13273_44868.n25 a_13273_44868.n2 27.8685
R54344 a_13273_44868.n0 a_13273_44868.t5 26.5955
R54345 a_13273_44868.n0 a_13273_44868.t6 26.5955
R54346 a_13273_44868.n1 a_13273_44868.t4 26.5955
R54347 a_13273_44868.n1 a_13273_44868.t7 26.5955
R54348 a_13273_44868.n27 a_13273_44868.n25 25.4811
R54349 a_13273_44868.n26 a_13273_44868.t1 24.9236
R54350 a_13273_44868.n26 a_13273_44868.t0 24.9236
R54351 a_13273_44868.n28 a_13273_44868.t2 24.9236
R54352 a_13273_44868.t3 a_13273_44868.n28 24.9236
R54353 a_13273_44868.n16 a_13273_44868.n14 18.4164
R54354 a_13273_44868.n11 a_13273_44868.n9 15.6475
R54355 a_13273_44868.n17 a_13273_44868.n16 15.5666
R54356 a_13273_44868.n24 a_13273_44868.n18 12.3027
R54357 a_13273_44868.n24 a_13273_44868.n23 11.9579
R54358 a_13273_44868.n25 a_13273_44868.n24 10.416
R54359 a_13273_44868.n18 a_13273_44868.n17 4.5005
R54360 a_13273_44868.n12 a_13273_44868.n11 1.23264
R54361 a_13273_44868.n14 a_13273_44868.n12 0.1255
R54362 C7_N_btm C7_N_btm.n3 62.1151
R54363 C7_N_btm.n3 C7_N_btm.t2 53.6613
R54364 C7_N_btm.n1 C7_N_btm.n0 52.9499
R54365 C7_N_btm.n1 C7_N_btm.t137 23.6451
R54366 C7_N_btm.n2 C7_N_btm.t138 23.6328
R54367 C7_N_btm.n2 C7_N_btm.n1 11.2505
R54368 C7_N_btm.n3 C7_N_btm.n2 8.41717
R54369 C7_N_btm C7_N_btm.n344 7.05675
R54370 C7_N_btm.n5 C7_N_btm.t135 5.03712
R54371 C7_N_btm.n41 C7_N_btm.t132 5.03712
R54372 C7_N_btm.n34 C7_N_btm.t136 5.03712
R54373 C7_N_btm.n35 C7_N_btm.t131 5.03712
R54374 C7_N_btm.n337 C7_N_btm.t134 5.03712
R54375 C7_N_btm.n99 C7_N_btm.t22 4.76719
R54376 C7_N_btm.n15 C7_N_btm.t61 4.76719
R54377 C7_N_btm.n340 C7_N_btm.n339 4.60698
R54378 C7_N_btm.n341 C7_N_btm.n340 4.60698
R54379 C7_N_btm.n334 C7_N_btm.n333 4.60698
R54380 C7_N_btm.n333 C7_N_btm.n332 4.60698
R54381 C7_N_btm.n328 C7_N_btm.n327 4.60698
R54382 C7_N_btm.n327 C7_N_btm.n325 4.60698
R54383 C7_N_btm.n319 C7_N_btm.n318 4.60698
R54384 C7_N_btm.n320 C7_N_btm.n319 4.60698
R54385 C7_N_btm.n313 C7_N_btm.n312 4.60698
R54386 C7_N_btm.n312 C7_N_btm.n311 4.60698
R54387 C7_N_btm.n307 C7_N_btm.n306 4.60698
R54388 C7_N_btm.n306 C7_N_btm.n304 4.60698
R54389 C7_N_btm.n298 C7_N_btm.n297 4.60698
R54390 C7_N_btm.n299 C7_N_btm.n298 4.60698
R54391 C7_N_btm.n292 C7_N_btm.n291 4.60698
R54392 C7_N_btm.n291 C7_N_btm.n290 4.60698
R54393 C7_N_btm.n286 C7_N_btm.n285 4.60698
R54394 C7_N_btm.n285 C7_N_btm.n283 4.60698
R54395 C7_N_btm.n276 C7_N_btm.n275 4.60698
R54396 C7_N_btm.n277 C7_N_btm.n276 4.60698
R54397 C7_N_btm.n279 C7_N_btm.n278 4.60698
R54398 C7_N_btm.n278 C7_N_btm.n20 4.60698
R54399 C7_N_btm.n267 C7_N_btm.n266 4.60698
R54400 C7_N_btm.n266 C7_N_btm.n265 4.60698
R54401 C7_N_btm.n270 C7_N_btm.n269 4.60698
R54402 C7_N_btm.n269 C7_N_btm.n268 4.60698
R54403 C7_N_btm.n190 C7_N_btm.n189 4.60698
R54404 C7_N_btm.n189 C7_N_btm.n188 4.60698
R54405 C7_N_btm.n192 C7_N_btm.n191 4.60698
R54406 C7_N_btm.n193 C7_N_btm.n192 4.60698
R54407 C7_N_btm.n195 C7_N_btm.n194 4.60698
R54408 C7_N_btm.n196 C7_N_btm.n195 4.60698
R54409 C7_N_btm.n198 C7_N_btm.n197 4.60698
R54410 C7_N_btm.n199 C7_N_btm.n198 4.60698
R54411 C7_N_btm.n201 C7_N_btm.n200 4.60698
R54412 C7_N_btm.n202 C7_N_btm.n201 4.60698
R54413 C7_N_btm.n204 C7_N_btm.n203 4.60698
R54414 C7_N_btm.n205 C7_N_btm.n204 4.60698
R54415 C7_N_btm.n207 C7_N_btm.n206 4.60698
R54416 C7_N_btm.n208 C7_N_btm.n207 4.60698
R54417 C7_N_btm.n210 C7_N_btm.n209 4.60698
R54418 C7_N_btm.n211 C7_N_btm.n210 4.60698
R54419 C7_N_btm.n213 C7_N_btm.n212 4.60698
R54420 C7_N_btm.n214 C7_N_btm.n213 4.60698
R54421 C7_N_btm.n216 C7_N_btm.n215 4.60698
R54422 C7_N_btm.n217 C7_N_btm.n216 4.60698
R54423 C7_N_btm.n219 C7_N_btm.n218 4.60698
R54424 C7_N_btm.n220 C7_N_btm.n219 4.60698
R54425 C7_N_btm.n222 C7_N_btm.n221 4.60698
R54426 C7_N_btm.n223 C7_N_btm.n222 4.60698
R54427 C7_N_btm.n225 C7_N_btm.n224 4.60698
R54428 C7_N_btm.n226 C7_N_btm.n225 4.60698
R54429 C7_N_btm.n228 C7_N_btm.n227 4.60698
R54430 C7_N_btm.n229 C7_N_btm.n228 4.60698
R54431 C7_N_btm.n231 C7_N_btm.n230 4.60698
R54432 C7_N_btm.n232 C7_N_btm.n231 4.60698
R54433 C7_N_btm.n234 C7_N_btm.n233 4.60698
R54434 C7_N_btm.n235 C7_N_btm.n234 4.60698
R54435 C7_N_btm.n238 C7_N_btm.n237 4.60698
R54436 C7_N_btm.n237 C7_N_btm.n236 4.60698
R54437 C7_N_btm.n144 C7_N_btm.n143 4.60698
R54438 C7_N_btm.n145 C7_N_btm.n144 4.60698
R54439 C7_N_btm.n147 C7_N_btm.n146 4.60698
R54440 C7_N_btm.n148 C7_N_btm.n147 4.60698
R54441 C7_N_btm.n150 C7_N_btm.n149 4.60698
R54442 C7_N_btm.n151 C7_N_btm.n150 4.60698
R54443 C7_N_btm.n153 C7_N_btm.n152 4.60698
R54444 C7_N_btm.n154 C7_N_btm.n153 4.60698
R54445 C7_N_btm.n156 C7_N_btm.n155 4.60698
R54446 C7_N_btm.n157 C7_N_btm.n156 4.60698
R54447 C7_N_btm.n159 C7_N_btm.n158 4.60698
R54448 C7_N_btm.n160 C7_N_btm.n159 4.60698
R54449 C7_N_btm.n162 C7_N_btm.n161 4.60698
R54450 C7_N_btm.n163 C7_N_btm.n162 4.60698
R54451 C7_N_btm.n165 C7_N_btm.n164 4.60698
R54452 C7_N_btm.n166 C7_N_btm.n165 4.60698
R54453 C7_N_btm.n168 C7_N_btm.n167 4.60698
R54454 C7_N_btm.n169 C7_N_btm.n168 4.60698
R54455 C7_N_btm.n171 C7_N_btm.n170 4.60698
R54456 C7_N_btm.n172 C7_N_btm.n171 4.60698
R54457 C7_N_btm.n174 C7_N_btm.n173 4.60698
R54458 C7_N_btm.n175 C7_N_btm.n174 4.60698
R54459 C7_N_btm.n177 C7_N_btm.n176 4.60698
R54460 C7_N_btm.n178 C7_N_btm.n177 4.60698
R54461 C7_N_btm.n180 C7_N_btm.n179 4.60698
R54462 C7_N_btm.n181 C7_N_btm.n180 4.60698
R54463 C7_N_btm.n183 C7_N_btm.n182 4.60698
R54464 C7_N_btm.n184 C7_N_btm.n183 4.60698
R54465 C7_N_btm.n241 C7_N_btm.n240 4.60698
R54466 C7_N_btm.n240 C7_N_btm.n239 4.60698
R54467 C7_N_btm.n247 C7_N_btm.n246 4.60698
R54468 C7_N_btm.n246 C7_N_btm.n245 4.60698
R54469 C7_N_btm.n250 C7_N_btm.n249 4.60698
R54470 C7_N_btm.n249 C7_N_btm.n248 4.60698
R54471 C7_N_btm.n105 C7_N_btm.n104 4.60698
R54472 C7_N_btm.n106 C7_N_btm.n105 4.60698
R54473 C7_N_btm.n108 C7_N_btm.n107 4.60698
R54474 C7_N_btm.n109 C7_N_btm.n108 4.60698
R54475 C7_N_btm.n95 C7_N_btm.n94 4.60698
R54476 C7_N_btm.n94 C7_N_btm.n93 4.60698
R54477 C7_N_btm.n89 C7_N_btm.n88 4.60698
R54478 C7_N_btm.n88 C7_N_btm.n86 4.60698
R54479 C7_N_btm.n80 C7_N_btm.n79 4.60698
R54480 C7_N_btm.n81 C7_N_btm.n80 4.60698
R54481 C7_N_btm.n74 C7_N_btm.n73 4.60698
R54482 C7_N_btm.n73 C7_N_btm.n72 4.60698
R54483 C7_N_btm.n68 C7_N_btm.n67 4.60698
R54484 C7_N_btm.n67 C7_N_btm.n65 4.60698
R54485 C7_N_btm.n59 C7_N_btm.n58 4.60698
R54486 C7_N_btm.n60 C7_N_btm.n59 4.60698
R54487 C7_N_btm.n53 C7_N_btm.n52 4.60698
R54488 C7_N_btm.n52 C7_N_btm.n51 4.60698
R54489 C7_N_btm.n47 C7_N_btm.n46 4.60698
R54490 C7_N_btm.n46 C7_N_btm.n44 4.60698
R54491 C7_N_btm.n38 C7_N_btm.n37 4.60698
R54492 C7_N_btm.n39 C7_N_btm.n38 4.60698
R54493 C7_N_btm.n344 C7_N_btm.t133 4.03712
R54494 C7_N_btm.n342 C7_N_btm.t11 3.98193
R54495 C7_N_btm.n331 C7_N_btm.t96 3.98193
R54496 C7_N_btm.n324 C7_N_btm.t104 3.98193
R54497 C7_N_btm.n321 C7_N_btm.t66 3.98193
R54498 C7_N_btm.n310 C7_N_btm.t77 3.98193
R54499 C7_N_btm.n303 C7_N_btm.t89 3.98193
R54500 C7_N_btm.n300 C7_N_btm.t53 3.98193
R54501 C7_N_btm.n289 C7_N_btm.t60 3.98193
R54502 C7_N_btm.n282 C7_N_btm.t12 3.98193
R54503 C7_N_btm.n21 C7_N_btm.t67 3.98193
R54504 C7_N_btm.n142 C7_N_btm.t125 3.98193
R54505 C7_N_btm.n185 C7_N_btm.t119 3.98193
R54506 C7_N_btm.n242 C7_N_btm.t54 3.98193
R54507 C7_N_btm.n244 C7_N_btm.t68 3.98193
R54508 C7_N_btm.n110 C7_N_btm.t58 3.98193
R54509 C7_N_btm.n92 C7_N_btm.t50 3.98193
R54510 C7_N_btm.n85 C7_N_btm.t87 3.98193
R54511 C7_N_btm.n82 C7_N_btm.t74 3.98193
R54512 C7_N_btm.n71 C7_N_btm.t3 3.98193
R54513 C7_N_btm.n64 C7_N_btm.t103 3.98193
R54514 C7_N_btm.n61 C7_N_btm.t95 3.98193
R54515 C7_N_btm.n50 C7_N_btm.t114 3.98193
R54516 C7_N_btm.n43 C7_N_btm.t98 3.98193
R54517 C7_N_btm.n40 C7_N_btm.t49 3.98193
R54518 C7_N_btm.n36 C7_N_btm.t122 3.98193
R54519 C7_N_btm.n45 C7_N_btm.t4 3.98193
R54520 C7_N_btm.n54 C7_N_btm.t19 3.98193
R54521 C7_N_btm.n57 C7_N_btm.t101 3.98193
R54522 C7_N_btm.n66 C7_N_btm.t41 3.98193
R54523 C7_N_btm.n75 C7_N_btm.t127 3.98193
R54524 C7_N_btm.n78 C7_N_btm.t84 3.98193
R54525 C7_N_btm.n87 C7_N_btm.t93 3.98193
R54526 C7_N_btm.n96 C7_N_btm.t124 3.98193
R54527 C7_N_btm.n271 C7_N_btm.t105 3.98193
R54528 C7_N_btm.n274 C7_N_btm.t97 3.98193
R54529 C7_N_btm.n284 C7_N_btm.t86 3.98193
R54530 C7_N_btm.n293 C7_N_btm.t72 3.98193
R54531 C7_N_btm.n296 C7_N_btm.t42 3.98193
R54532 C7_N_btm.n305 C7_N_btm.t35 3.98193
R54533 C7_N_btm.n314 C7_N_btm.t25 3.98193
R54534 C7_N_btm.n317 C7_N_btm.t23 3.98193
R54535 C7_N_btm.n326 C7_N_btm.t126 3.98193
R54536 C7_N_btm.n335 C7_N_btm.t47 3.98193
R54537 C7_N_btm.n338 C7_N_btm.t85 3.98193
R54538 C7_N_btm.n103 C7_N_btm.t28 3.92851
R54539 C7_N_btm.n102 C7_N_btm.t69 3.92851
R54540 C7_N_btm.n101 C7_N_btm.t123 3.92851
R54541 C7_N_btm.n100 C7_N_btm.t75 3.92851
R54542 C7_N_btm.n99 C7_N_btm.t118 3.92851
R54543 C7_N_btm.n251 C7_N_btm.t121 3.92851
R54544 C7_N_btm.n252 C7_N_btm.t81 3.92851
R54545 C7_N_btm.n253 C7_N_btm.t57 3.92851
R54546 C7_N_btm.n254 C7_N_btm.t88 3.92851
R54547 C7_N_btm.n255 C7_N_btm.t63 3.92851
R54548 C7_N_btm.n256 C7_N_btm.t34 3.92851
R54549 C7_N_btm.n257 C7_N_btm.t71 3.92851
R54550 C7_N_btm.n258 C7_N_btm.t117 3.92851
R54551 C7_N_btm.n259 C7_N_btm.t55 3.92851
R54552 C7_N_btm.n260 C7_N_btm.t112 3.92851
R54553 C7_N_btm.n261 C7_N_btm.t16 3.92851
R54554 C7_N_btm.n262 C7_N_btm.t129 3.92851
R54555 C7_N_btm.n263 C7_N_btm.t31 3.92851
R54556 C7_N_btm.n264 C7_N_btm.t24 3.92851
R54557 C7_N_btm.n19 C7_N_btm.t107 3.92851
R54558 C7_N_btm.n18 C7_N_btm.t18 3.92851
R54559 C7_N_btm.n17 C7_N_btm.t52 3.92851
R54560 C7_N_btm.n16 C7_N_btm.t33 3.92851
R54561 C7_N_btm.n15 C7_N_btm.t43 3.92851
R54562 C7_N_btm.n0 C7_N_btm.t1 3.57113
R54563 C7_N_btm.n0 C7_N_btm.t0 3.57113
R54564 C7_N_btm.n340 C7_N_btm.t108 1.67819
R54565 C7_N_btm.n333 C7_N_btm.t70 1.67819
R54566 C7_N_btm.n327 C7_N_btm.t38 1.67819
R54567 C7_N_btm.n319 C7_N_btm.t40 1.67819
R54568 C7_N_btm.n312 C7_N_btm.t111 1.67819
R54569 C7_N_btm.n306 C7_N_btm.t64 1.67819
R54570 C7_N_btm.n298 C7_N_btm.t17 1.67819
R54571 C7_N_btm.n291 C7_N_btm.t29 1.67819
R54572 C7_N_btm.n285 C7_N_btm.t110 1.67819
R54573 C7_N_btm.n276 C7_N_btm.t115 1.67819
R54574 C7_N_btm.n278 C7_N_btm.t83 1.67819
R54575 C7_N_btm.n266 C7_N_btm.t37 1.67819
R54576 C7_N_btm.n269 C7_N_btm.t6 1.67819
R54577 C7_N_btm.n189 C7_N_btm.t92 1.67819
R54578 C7_N_btm.n192 C7_N_btm.t44 1.67819
R54579 C7_N_btm.n195 C7_N_btm.t80 1.67819
R54580 C7_N_btm.n198 C7_N_btm.t9 1.67819
R54581 C7_N_btm.n201 C7_N_btm.t13 1.67819
R54582 C7_N_btm.n204 C7_N_btm.t99 1.67819
R54583 C7_N_btm.n207 C7_N_btm.t5 1.67819
R54584 C7_N_btm.n210 C7_N_btm.t94 1.67819
R54585 C7_N_btm.n213 C7_N_btm.t46 1.67819
R54586 C7_N_btm.n216 C7_N_btm.t30 1.67819
R54587 C7_N_btm.n219 C7_N_btm.t116 1.67819
R54588 C7_N_btm.n222 C7_N_btm.t15 1.67819
R54589 C7_N_btm.n225 C7_N_btm.t51 1.67819
R54590 C7_N_btm.n228 C7_N_btm.t10 1.67819
R54591 C7_N_btm.n231 C7_N_btm.t39 1.67819
R54592 C7_N_btm.n234 C7_N_btm.t48 1.67819
R54593 C7_N_btm.n237 C7_N_btm.t32 1.67819
R54594 C7_N_btm.n144 C7_N_btm.t7 1.67819
R54595 C7_N_btm.n147 C7_N_btm.t82 1.67819
R54596 C7_N_btm.n150 C7_N_btm.t21 1.67819
R54597 C7_N_btm.n153 C7_N_btm.t128 1.67819
R54598 C7_N_btm.n156 C7_N_btm.t27 1.67819
R54599 C7_N_btm.n159 C7_N_btm.t76 1.67819
R54600 C7_N_btm.n162 C7_N_btm.t45 1.67819
R54601 C7_N_btm.n165 C7_N_btm.t65 1.67819
R54602 C7_N_btm.n168 C7_N_btm.t102 1.67819
R54603 C7_N_btm.n171 C7_N_btm.t20 1.67819
R54604 C7_N_btm.n174 C7_N_btm.t109 1.67819
R54605 C7_N_btm.n177 C7_N_btm.t113 1.67819
R54606 C7_N_btm.n180 C7_N_btm.t59 1.67819
R54607 C7_N_btm.n183 C7_N_btm.t91 1.67819
R54608 C7_N_btm.n240 C7_N_btm.t62 1.67819
R54609 C7_N_btm.n246 C7_N_btm.t100 1.67819
R54610 C7_N_btm.n249 C7_N_btm.t73 1.67819
R54611 C7_N_btm.n105 C7_N_btm.t130 1.67819
R54612 C7_N_btm.n108 C7_N_btm.t90 1.67819
R54613 C7_N_btm.n94 C7_N_btm.t79 1.67819
R54614 C7_N_btm.n88 C7_N_btm.t8 1.67819
R54615 C7_N_btm.n80 C7_N_btm.t106 1.67819
R54616 C7_N_btm.n73 C7_N_btm.t26 1.67819
R54617 C7_N_btm.n67 C7_N_btm.t14 1.67819
R54618 C7_N_btm.n59 C7_N_btm.t120 1.67819
R54619 C7_N_btm.n52 C7_N_btm.t56 1.67819
R54620 C7_N_btm.n46 C7_N_btm.t36 1.67819
R54621 C7_N_btm.n38 C7_N_btm.t78 1.67819
R54622 C7_N_btm.n186 C7_N_btm.n185 1.05569
R54623 C7_N_btm.n142 C7_N_btm.n113 1.05569
R54624 C7_N_btm.n243 C7_N_btm.n242 1.05569
R54625 C7_N_btm.n272 C7_N_btm.n21 1.05569
R54626 C7_N_btm.n330 C7_N_btm.n5 1.0005
R54627 C7_N_btm.n330 C7_N_btm.n329 1.0005
R54628 C7_N_btm.n329 C7_N_btm.n7 1.0005
R54629 C7_N_btm.n309 C7_N_btm.n7 1.0005
R54630 C7_N_btm.n309 C7_N_btm.n308 1.0005
R54631 C7_N_btm.n308 C7_N_btm.n10 1.0005
R54632 C7_N_btm.n288 C7_N_btm.n10 1.0005
R54633 C7_N_btm.n288 C7_N_btm.n287 1.0005
R54634 C7_N_btm.n287 C7_N_btm.n13 1.0005
R54635 C7_N_btm.n22 C7_N_btm.n13 1.0005
R54636 C7_N_btm.n187 C7_N_btm.n22 1.0005
R54637 C7_N_btm.n186 C7_N_btm.n14 1.0005
R54638 C7_N_btm.n141 C7_N_btm.n114 1.0005
R54639 C7_N_btm.n140 C7_N_btm.n115 1.0005
R54640 C7_N_btm.n139 C7_N_btm.n116 1.0005
R54641 C7_N_btm.n138 C7_N_btm.n117 1.0005
R54642 C7_N_btm.n137 C7_N_btm.n118 1.0005
R54643 C7_N_btm.n136 C7_N_btm.n119 1.0005
R54644 C7_N_btm.n135 C7_N_btm.n120 1.0005
R54645 C7_N_btm.n134 C7_N_btm.n121 1.0005
R54646 C7_N_btm.n133 C7_N_btm.n122 1.0005
R54647 C7_N_btm.n132 C7_N_btm.n123 1.0005
R54648 C7_N_btm.n131 C7_N_btm.n124 1.0005
R54649 C7_N_btm.n130 C7_N_btm.n125 1.0005
R54650 C7_N_btm.n129 C7_N_btm.n126 1.0005
R54651 C7_N_btm.n128 C7_N_btm.n127 1.0005
R54652 C7_N_btm.n112 C7_N_btm.n24 1.0005
R54653 C7_N_btm.n26 C7_N_btm.n24 1.0005
R54654 C7_N_btm.n91 C7_N_btm.n26 1.0005
R54655 C7_N_btm.n91 C7_N_btm.n90 1.0005
R54656 C7_N_btm.n90 C7_N_btm.n28 1.0005
R54657 C7_N_btm.n70 C7_N_btm.n28 1.0005
R54658 C7_N_btm.n70 C7_N_btm.n69 1.0005
R54659 C7_N_btm.n69 C7_N_btm.n31 1.0005
R54660 C7_N_btm.n49 C7_N_btm.n31 1.0005
R54661 C7_N_btm.n49 C7_N_btm.n48 1.0005
R54662 C7_N_btm.n48 C7_N_btm.n34 1.0005
R54663 C7_N_btm.n35 C7_N_btm.n33 1.0005
R54664 C7_N_btm.n42 C7_N_btm.n41 1.0005
R54665 C7_N_btm.n42 C7_N_btm.n32 1.0005
R54666 C7_N_btm.n55 C7_N_btm.n33 1.0005
R54667 C7_N_btm.n56 C7_N_btm.n55 1.0005
R54668 C7_N_btm.n62 C7_N_btm.n32 1.0005
R54669 C7_N_btm.n63 C7_N_btm.n62 1.0005
R54670 C7_N_btm.n56 C7_N_btm.n30 1.0005
R54671 C7_N_btm.n76 C7_N_btm.n30 1.0005
R54672 C7_N_btm.n63 C7_N_btm.n29 1.0005
R54673 C7_N_btm.n83 C7_N_btm.n29 1.0005
R54674 C7_N_btm.n77 C7_N_btm.n76 1.0005
R54675 C7_N_btm.n77 C7_N_btm.n27 1.0005
R54676 C7_N_btm.n84 C7_N_btm.n83 1.0005
R54677 C7_N_btm.n84 C7_N_btm.n25 1.0005
R54678 C7_N_btm.n97 C7_N_btm.n27 1.0005
R54679 C7_N_btm.n98 C7_N_btm.n97 1.0005
R54680 C7_N_btm.n111 C7_N_btm.n25 1.0005
R54681 C7_N_btm.n243 C7_N_btm.n111 1.0005
R54682 C7_N_btm.n98 C7_N_btm.n23 1.0005
R54683 C7_N_btm.n113 C7_N_btm.n23 1.0005
R54684 C7_N_btm.n273 C7_N_btm.n272 1.0005
R54685 C7_N_btm.n281 C7_N_btm.n280 1.0005
R54686 C7_N_btm.n280 C7_N_btm.n14 1.0005
R54687 C7_N_btm.n294 C7_N_btm.n12 1.0005
R54688 C7_N_btm.n273 C7_N_btm.n12 1.0005
R54689 C7_N_btm.n301 C7_N_btm.n11 1.0005
R54690 C7_N_btm.n281 C7_N_btm.n11 1.0005
R54691 C7_N_btm.n295 C7_N_btm.n9 1.0005
R54692 C7_N_btm.n295 C7_N_btm.n294 1.0005
R54693 C7_N_btm.n302 C7_N_btm.n8 1.0005
R54694 C7_N_btm.n302 C7_N_btm.n301 1.0005
R54695 C7_N_btm.n316 C7_N_btm.n315 1.0005
R54696 C7_N_btm.n315 C7_N_btm.n9 1.0005
R54697 C7_N_btm.n323 C7_N_btm.n322 1.0005
R54698 C7_N_btm.n322 C7_N_btm.n8 1.0005
R54699 C7_N_btm.n336 C7_N_btm.n6 1.0005
R54700 C7_N_btm.n316 C7_N_btm.n6 1.0005
R54701 C7_N_btm.n343 C7_N_btm.n4 1.0005
R54702 C7_N_btm.n323 C7_N_btm.n4 1.0005
R54703 C7_N_btm.n337 C7_N_btm.n336 1.0005
R54704 C7_N_btm.n344 C7_N_btm.n343 1.0005
R54705 C7_N_btm.n100 C7_N_btm.n99 0.840176
R54706 C7_N_btm.n101 C7_N_btm.n100 0.840176
R54707 C7_N_btm.n102 C7_N_btm.n101 0.840176
R54708 C7_N_btm.n103 C7_N_btm.n102 0.840176
R54709 C7_N_btm.n264 C7_N_btm.n263 0.840176
R54710 C7_N_btm.n263 C7_N_btm.n262 0.840176
R54711 C7_N_btm.n262 C7_N_btm.n261 0.840176
R54712 C7_N_btm.n261 C7_N_btm.n260 0.840176
R54713 C7_N_btm.n260 C7_N_btm.n259 0.840176
R54714 C7_N_btm.n259 C7_N_btm.n258 0.840176
R54715 C7_N_btm.n258 C7_N_btm.n257 0.840176
R54716 C7_N_btm.n257 C7_N_btm.n256 0.840176
R54717 C7_N_btm.n256 C7_N_btm.n255 0.840176
R54718 C7_N_btm.n255 C7_N_btm.n254 0.840176
R54719 C7_N_btm.n254 C7_N_btm.n253 0.840176
R54720 C7_N_btm.n253 C7_N_btm.n252 0.840176
R54721 C7_N_btm.n252 C7_N_btm.n251 0.840176
R54722 C7_N_btm.n16 C7_N_btm.n15 0.840176
R54723 C7_N_btm.n17 C7_N_btm.n16 0.840176
R54724 C7_N_btm.n18 C7_N_btm.n17 0.840176
R54725 C7_N_btm.n19 C7_N_btm.n18 0.840176
R54726 C7_N_btm.n104 C7_N_btm.n103 0.732838
R54727 C7_N_btm.n265 C7_N_btm.n264 0.732838
R54728 C7_N_btm.n251 C7_N_btm.n250 0.732838
R54729 C7_N_btm.n20 C7_N_btm.n19 0.732838
R54730 C7_N_btm.n185 C7_N_btm.n184 0.679419
R54731 C7_N_btm.n143 C7_N_btm.n142 0.679419
R54732 C7_N_btm.n37 C7_N_btm.n36 0.679419
R54733 C7_N_btm.n40 C7_N_btm.n39 0.679419
R54734 C7_N_btm.n44 C7_N_btm.n43 0.679419
R54735 C7_N_btm.n47 C7_N_btm.n45 0.679419
R54736 C7_N_btm.n54 C7_N_btm.n53 0.679419
R54737 C7_N_btm.n51 C7_N_btm.n50 0.679419
R54738 C7_N_btm.n61 C7_N_btm.n60 0.679419
R54739 C7_N_btm.n58 C7_N_btm.n57 0.679419
R54740 C7_N_btm.n68 C7_N_btm.n66 0.679419
R54741 C7_N_btm.n65 C7_N_btm.n64 0.679419
R54742 C7_N_btm.n72 C7_N_btm.n71 0.679419
R54743 C7_N_btm.n75 C7_N_btm.n74 0.679419
R54744 C7_N_btm.n79 C7_N_btm.n78 0.679419
R54745 C7_N_btm.n82 C7_N_btm.n81 0.679419
R54746 C7_N_btm.n86 C7_N_btm.n85 0.679419
R54747 C7_N_btm.n89 C7_N_btm.n87 0.679419
R54748 C7_N_btm.n96 C7_N_btm.n95 0.679419
R54749 C7_N_btm.n93 C7_N_btm.n92 0.679419
R54750 C7_N_btm.n110 C7_N_btm.n109 0.679419
R54751 C7_N_btm.n245 C7_N_btm.n244 0.679419
R54752 C7_N_btm.n242 C7_N_btm.n241 0.679419
R54753 C7_N_btm.n188 C7_N_btm.n21 0.679419
R54754 C7_N_btm.n271 C7_N_btm.n270 0.679419
R54755 C7_N_btm.n275 C7_N_btm.n274 0.679419
R54756 C7_N_btm.n286 C7_N_btm.n284 0.679419
R54757 C7_N_btm.n283 C7_N_btm.n282 0.679419
R54758 C7_N_btm.n290 C7_N_btm.n289 0.679419
R54759 C7_N_btm.n293 C7_N_btm.n292 0.679419
R54760 C7_N_btm.n297 C7_N_btm.n296 0.679419
R54761 C7_N_btm.n300 C7_N_btm.n299 0.679419
R54762 C7_N_btm.n304 C7_N_btm.n303 0.679419
R54763 C7_N_btm.n307 C7_N_btm.n305 0.679419
R54764 C7_N_btm.n314 C7_N_btm.n313 0.679419
R54765 C7_N_btm.n311 C7_N_btm.n310 0.679419
R54766 C7_N_btm.n321 C7_N_btm.n320 0.679419
R54767 C7_N_btm.n318 C7_N_btm.n317 0.679419
R54768 C7_N_btm.n328 C7_N_btm.n326 0.679419
R54769 C7_N_btm.n325 C7_N_btm.n324 0.679419
R54770 C7_N_btm.n332 C7_N_btm.n331 0.679419
R54771 C7_N_btm.n335 C7_N_btm.n334 0.679419
R54772 C7_N_btm.n339 C7_N_btm.n338 0.679419
R54773 C7_N_btm.n342 C7_N_btm.n341 0.679419
R54774 C7_N_btm.n182 C7_N_btm.n181 0.6255
R54775 C7_N_btm.n179 C7_N_btm.n178 0.6255
R54776 C7_N_btm.n176 C7_N_btm.n175 0.6255
R54777 C7_N_btm.n173 C7_N_btm.n172 0.6255
R54778 C7_N_btm.n170 C7_N_btm.n169 0.6255
R54779 C7_N_btm.n167 C7_N_btm.n166 0.6255
R54780 C7_N_btm.n164 C7_N_btm.n163 0.6255
R54781 C7_N_btm.n161 C7_N_btm.n160 0.6255
R54782 C7_N_btm.n158 C7_N_btm.n157 0.6255
R54783 C7_N_btm.n155 C7_N_btm.n154 0.6255
R54784 C7_N_btm.n152 C7_N_btm.n151 0.6255
R54785 C7_N_btm.n149 C7_N_btm.n148 0.6255
R54786 C7_N_btm.n146 C7_N_btm.n145 0.6255
R54787 C7_N_btm.n107 C7_N_btm.n106 0.6255
R54788 C7_N_btm.n248 C7_N_btm.n247 0.6255
R54789 C7_N_btm.n239 C7_N_btm.n238 0.6255
R54790 C7_N_btm.n236 C7_N_btm.n235 0.6255
R54791 C7_N_btm.n233 C7_N_btm.n232 0.6255
R54792 C7_N_btm.n230 C7_N_btm.n229 0.6255
R54793 C7_N_btm.n227 C7_N_btm.n226 0.6255
R54794 C7_N_btm.n224 C7_N_btm.n223 0.6255
R54795 C7_N_btm.n221 C7_N_btm.n220 0.6255
R54796 C7_N_btm.n218 C7_N_btm.n217 0.6255
R54797 C7_N_btm.n215 C7_N_btm.n214 0.6255
R54798 C7_N_btm.n212 C7_N_btm.n211 0.6255
R54799 C7_N_btm.n209 C7_N_btm.n208 0.6255
R54800 C7_N_btm.n206 C7_N_btm.n205 0.6255
R54801 C7_N_btm.n203 C7_N_btm.n202 0.6255
R54802 C7_N_btm.n200 C7_N_btm.n199 0.6255
R54803 C7_N_btm.n197 C7_N_btm.n196 0.6255
R54804 C7_N_btm.n194 C7_N_btm.n193 0.6255
R54805 C7_N_btm.n191 C7_N_btm.n190 0.6255
R54806 C7_N_btm.n268 C7_N_btm.n267 0.6255
R54807 C7_N_btm.n279 C7_N_btm.n277 0.6255
R54808 C7_N_btm.n182 C7_N_btm.n128 0.109875
R54809 C7_N_btm.n184 C7_N_btm.n128 0.109875
R54810 C7_N_btm.n179 C7_N_btm.n129 0.109875
R54811 C7_N_btm.n181 C7_N_btm.n129 0.109875
R54812 C7_N_btm.n176 C7_N_btm.n130 0.109875
R54813 C7_N_btm.n178 C7_N_btm.n130 0.109875
R54814 C7_N_btm.n173 C7_N_btm.n131 0.109875
R54815 C7_N_btm.n175 C7_N_btm.n131 0.109875
R54816 C7_N_btm.n170 C7_N_btm.n132 0.109875
R54817 C7_N_btm.n172 C7_N_btm.n132 0.109875
R54818 C7_N_btm.n167 C7_N_btm.n133 0.109875
R54819 C7_N_btm.n169 C7_N_btm.n133 0.109875
R54820 C7_N_btm.n164 C7_N_btm.n134 0.109875
R54821 C7_N_btm.n166 C7_N_btm.n134 0.109875
R54822 C7_N_btm.n161 C7_N_btm.n135 0.109875
R54823 C7_N_btm.n163 C7_N_btm.n135 0.109875
R54824 C7_N_btm.n158 C7_N_btm.n136 0.109875
R54825 C7_N_btm.n160 C7_N_btm.n136 0.109875
R54826 C7_N_btm.n155 C7_N_btm.n137 0.109875
R54827 C7_N_btm.n157 C7_N_btm.n137 0.109875
R54828 C7_N_btm.n152 C7_N_btm.n138 0.109875
R54829 C7_N_btm.n154 C7_N_btm.n138 0.109875
R54830 C7_N_btm.n149 C7_N_btm.n139 0.109875
R54831 C7_N_btm.n151 C7_N_btm.n139 0.109875
R54832 C7_N_btm.n146 C7_N_btm.n140 0.109875
R54833 C7_N_btm.n148 C7_N_btm.n140 0.109875
R54834 C7_N_btm.n143 C7_N_btm.n141 0.109875
R54835 C7_N_btm.n145 C7_N_btm.n141 0.109875
R54836 C7_N_btm.n39 C7_N_btm.n34 0.109875
R54837 C7_N_btm.n37 C7_N_btm.n34 0.109875
R54838 C7_N_btm.n48 C7_N_btm.n44 0.109875
R54839 C7_N_btm.n48 C7_N_btm.n47 0.109875
R54840 C7_N_btm.n51 C7_N_btm.n49 0.109875
R54841 C7_N_btm.n53 C7_N_btm.n49 0.109875
R54842 C7_N_btm.n60 C7_N_btm.n31 0.109875
R54843 C7_N_btm.n58 C7_N_btm.n31 0.109875
R54844 C7_N_btm.n69 C7_N_btm.n65 0.109875
R54845 C7_N_btm.n69 C7_N_btm.n68 0.109875
R54846 C7_N_btm.n72 C7_N_btm.n70 0.109875
R54847 C7_N_btm.n74 C7_N_btm.n70 0.109875
R54848 C7_N_btm.n81 C7_N_btm.n28 0.109875
R54849 C7_N_btm.n79 C7_N_btm.n28 0.109875
R54850 C7_N_btm.n90 C7_N_btm.n86 0.109875
R54851 C7_N_btm.n90 C7_N_btm.n89 0.109875
R54852 C7_N_btm.n93 C7_N_btm.n91 0.109875
R54853 C7_N_btm.n95 C7_N_btm.n91 0.109875
R54854 C7_N_btm.n109 C7_N_btm.n26 0.109875
R54855 C7_N_btm.n107 C7_N_btm.n26 0.109875
R54856 C7_N_btm.n106 C7_N_btm.n98 0.109875
R54857 C7_N_btm.n104 C7_N_btm.n98 0.109875
R54858 C7_N_btm.n248 C7_N_btm.n23 0.109875
R54859 C7_N_btm.n250 C7_N_btm.n23 0.109875
R54860 C7_N_btm.n245 C7_N_btm.n24 0.109875
R54861 C7_N_btm.n247 C7_N_btm.n24 0.109875
R54862 C7_N_btm.n241 C7_N_btm.n112 0.109875
R54863 C7_N_btm.n239 C7_N_btm.n112 0.109875
R54864 C7_N_btm.n238 C7_N_btm.n113 0.109875
R54865 C7_N_btm.n236 C7_N_btm.n113 0.109875
R54866 C7_N_btm.n235 C7_N_btm.n114 0.109875
R54867 C7_N_btm.n233 C7_N_btm.n114 0.109875
R54868 C7_N_btm.n232 C7_N_btm.n115 0.109875
R54869 C7_N_btm.n230 C7_N_btm.n115 0.109875
R54870 C7_N_btm.n229 C7_N_btm.n116 0.109875
R54871 C7_N_btm.n227 C7_N_btm.n116 0.109875
R54872 C7_N_btm.n226 C7_N_btm.n117 0.109875
R54873 C7_N_btm.n224 C7_N_btm.n117 0.109875
R54874 C7_N_btm.n223 C7_N_btm.n118 0.109875
R54875 C7_N_btm.n221 C7_N_btm.n118 0.109875
R54876 C7_N_btm.n220 C7_N_btm.n119 0.109875
R54877 C7_N_btm.n218 C7_N_btm.n119 0.109875
R54878 C7_N_btm.n217 C7_N_btm.n120 0.109875
R54879 C7_N_btm.n215 C7_N_btm.n120 0.109875
R54880 C7_N_btm.n214 C7_N_btm.n121 0.109875
R54881 C7_N_btm.n212 C7_N_btm.n121 0.109875
R54882 C7_N_btm.n211 C7_N_btm.n122 0.109875
R54883 C7_N_btm.n209 C7_N_btm.n122 0.109875
R54884 C7_N_btm.n208 C7_N_btm.n123 0.109875
R54885 C7_N_btm.n206 C7_N_btm.n123 0.109875
R54886 C7_N_btm.n205 C7_N_btm.n124 0.109875
R54887 C7_N_btm.n203 C7_N_btm.n124 0.109875
R54888 C7_N_btm.n202 C7_N_btm.n125 0.109875
R54889 C7_N_btm.n200 C7_N_btm.n125 0.109875
R54890 C7_N_btm.n199 C7_N_btm.n126 0.109875
R54891 C7_N_btm.n197 C7_N_btm.n126 0.109875
R54892 C7_N_btm.n196 C7_N_btm.n127 0.109875
R54893 C7_N_btm.n194 C7_N_btm.n127 0.109875
R54894 C7_N_btm.n193 C7_N_btm.n186 0.109875
R54895 C7_N_btm.n191 C7_N_btm.n186 0.109875
R54896 C7_N_btm.n190 C7_N_btm.n187 0.109875
R54897 C7_N_btm.n188 C7_N_btm.n187 0.109875
R54898 C7_N_btm.n268 C7_N_btm.n22 0.109875
R54899 C7_N_btm.n270 C7_N_btm.n22 0.109875
R54900 C7_N_btm.n265 C7_N_btm.n14 0.109875
R54901 C7_N_btm.n267 C7_N_btm.n14 0.109875
R54902 C7_N_btm.n280 C7_N_btm.n20 0.109875
R54903 C7_N_btm.n280 C7_N_btm.n279 0.109875
R54904 C7_N_btm.n277 C7_N_btm.n13 0.109875
R54905 C7_N_btm.n275 C7_N_btm.n13 0.109875
R54906 C7_N_btm.n287 C7_N_btm.n283 0.109875
R54907 C7_N_btm.n287 C7_N_btm.n286 0.109875
R54908 C7_N_btm.n290 C7_N_btm.n288 0.109875
R54909 C7_N_btm.n292 C7_N_btm.n288 0.109875
R54910 C7_N_btm.n299 C7_N_btm.n10 0.109875
R54911 C7_N_btm.n297 C7_N_btm.n10 0.109875
R54912 C7_N_btm.n308 C7_N_btm.n304 0.109875
R54913 C7_N_btm.n308 C7_N_btm.n307 0.109875
R54914 C7_N_btm.n311 C7_N_btm.n309 0.109875
R54915 C7_N_btm.n313 C7_N_btm.n309 0.109875
R54916 C7_N_btm.n320 C7_N_btm.n7 0.109875
R54917 C7_N_btm.n318 C7_N_btm.n7 0.109875
R54918 C7_N_btm.n329 C7_N_btm.n325 0.109875
R54919 C7_N_btm.n329 C7_N_btm.n328 0.109875
R54920 C7_N_btm.n332 C7_N_btm.n330 0.109875
R54921 C7_N_btm.n334 C7_N_btm.n330 0.109875
R54922 C7_N_btm.n341 C7_N_btm.n5 0.109875
R54923 C7_N_btm.n339 C7_N_btm.n5 0.109875
R54924 C7_N_btm.n36 C7_N_btm.n35 0.0556875
R54925 C7_N_btm.n41 C7_N_btm.n40 0.0556875
R54926 C7_N_btm.n43 C7_N_btm.n42 0.0556875
R54927 C7_N_btm.n45 C7_N_btm.n33 0.0556875
R54928 C7_N_btm.n55 C7_N_btm.n54 0.0556875
R54929 C7_N_btm.n50 C7_N_btm.n32 0.0556875
R54930 C7_N_btm.n62 C7_N_btm.n61 0.0556875
R54931 C7_N_btm.n57 C7_N_btm.n56 0.0556875
R54932 C7_N_btm.n66 C7_N_btm.n30 0.0556875
R54933 C7_N_btm.n64 C7_N_btm.n63 0.0556875
R54934 C7_N_btm.n71 C7_N_btm.n29 0.0556875
R54935 C7_N_btm.n76 C7_N_btm.n75 0.0556875
R54936 C7_N_btm.n78 C7_N_btm.n77 0.0556875
R54937 C7_N_btm.n83 C7_N_btm.n82 0.0556875
R54938 C7_N_btm.n85 C7_N_btm.n84 0.0556875
R54939 C7_N_btm.n87 C7_N_btm.n27 0.0556875
R54940 C7_N_btm.n97 C7_N_btm.n96 0.0556875
R54941 C7_N_btm.n92 C7_N_btm.n25 0.0556875
R54942 C7_N_btm.n111 C7_N_btm.n110 0.0556875
R54943 C7_N_btm.n244 C7_N_btm.n243 0.0556875
R54944 C7_N_btm.n272 C7_N_btm.n271 0.0556875
R54945 C7_N_btm.n274 C7_N_btm.n273 0.0556875
R54946 C7_N_btm.n284 C7_N_btm.n12 0.0556875
R54947 C7_N_btm.n282 C7_N_btm.n281 0.0556875
R54948 C7_N_btm.n289 C7_N_btm.n11 0.0556875
R54949 C7_N_btm.n294 C7_N_btm.n293 0.0556875
R54950 C7_N_btm.n296 C7_N_btm.n295 0.0556875
R54951 C7_N_btm.n301 C7_N_btm.n300 0.0556875
R54952 C7_N_btm.n303 C7_N_btm.n302 0.0556875
R54953 C7_N_btm.n305 C7_N_btm.n9 0.0556875
R54954 C7_N_btm.n315 C7_N_btm.n314 0.0556875
R54955 C7_N_btm.n310 C7_N_btm.n8 0.0556875
R54956 C7_N_btm.n322 C7_N_btm.n321 0.0556875
R54957 C7_N_btm.n317 C7_N_btm.n316 0.0556875
R54958 C7_N_btm.n326 C7_N_btm.n6 0.0556875
R54959 C7_N_btm.n324 C7_N_btm.n323 0.0556875
R54960 C7_N_btm.n331 C7_N_btm.n4 0.0556875
R54961 C7_N_btm.n336 C7_N_btm.n335 0.0556875
R54962 C7_N_btm.n338 C7_N_btm.n337 0.0556875
R54963 C7_N_btm.n343 C7_N_btm.n342 0.0556875
R54964 C7_P_btm C7_P_btm.n3 62.2088
R54965 C7_P_btm.n3 C7_P_btm.t0 53.6613
R54966 C7_P_btm.n1 C7_P_btm.n0 52.9499
R54967 C7_P_btm.n1 C7_P_btm.t137 23.6451
R54968 C7_P_btm.n2 C7_P_btm.t138 23.6328
R54969 C7_P_btm.n2 C7_P_btm.n1 11.2505
R54970 C7_P_btm.n3 C7_P_btm.n2 8.41717
R54971 C7_P_btm C7_P_btm.n344 6.963
R54972 C7_P_btm.n5 C7_P_btm.t7 5.03712
R54973 C7_P_btm.n337 C7_P_btm.t5 5.03712
R54974 C7_P_btm.n41 C7_P_btm.t4 5.03712
R54975 C7_P_btm.n34 C7_P_btm.t3 5.03712
R54976 C7_P_btm.n35 C7_P_btm.t8 5.03712
R54977 C7_P_btm.n99 C7_P_btm.t99 4.76719
R54978 C7_P_btm.n15 C7_P_btm.t75 4.76719
R54979 C7_P_btm.n341 C7_P_btm.n340 4.60698
R54980 C7_P_btm.n340 C7_P_btm.n339 4.60698
R54981 C7_P_btm.n334 C7_P_btm.n333 4.60698
R54982 C7_P_btm.n333 C7_P_btm.n332 4.60698
R54983 C7_P_btm.n328 C7_P_btm.n327 4.60698
R54984 C7_P_btm.n327 C7_P_btm.n325 4.60698
R54985 C7_P_btm.n319 C7_P_btm.n318 4.60698
R54986 C7_P_btm.n320 C7_P_btm.n319 4.60698
R54987 C7_P_btm.n313 C7_P_btm.n312 4.60698
R54988 C7_P_btm.n312 C7_P_btm.n311 4.60698
R54989 C7_P_btm.n307 C7_P_btm.n306 4.60698
R54990 C7_P_btm.n306 C7_P_btm.n304 4.60698
R54991 C7_P_btm.n298 C7_P_btm.n297 4.60698
R54992 C7_P_btm.n299 C7_P_btm.n298 4.60698
R54993 C7_P_btm.n292 C7_P_btm.n291 4.60698
R54994 C7_P_btm.n291 C7_P_btm.n290 4.60698
R54995 C7_P_btm.n286 C7_P_btm.n285 4.60698
R54996 C7_P_btm.n285 C7_P_btm.n283 4.60698
R54997 C7_P_btm.n276 C7_P_btm.n275 4.60698
R54998 C7_P_btm.n277 C7_P_btm.n276 4.60698
R54999 C7_P_btm.n279 C7_P_btm.n278 4.60698
R55000 C7_P_btm.n278 C7_P_btm.n20 4.60698
R55001 C7_P_btm.n266 C7_P_btm.n265 4.60698
R55002 C7_P_btm.n267 C7_P_btm.n266 4.60698
R55003 C7_P_btm.n270 C7_P_btm.n269 4.60698
R55004 C7_P_btm.n269 C7_P_btm.n268 4.60698
R55005 C7_P_btm.n189 C7_P_btm.n188 4.60698
R55006 C7_P_btm.n190 C7_P_btm.n189 4.60698
R55007 C7_P_btm.n192 C7_P_btm.n191 4.60698
R55008 C7_P_btm.n193 C7_P_btm.n192 4.60698
R55009 C7_P_btm.n195 C7_P_btm.n194 4.60698
R55010 C7_P_btm.n196 C7_P_btm.n195 4.60698
R55011 C7_P_btm.n198 C7_P_btm.n197 4.60698
R55012 C7_P_btm.n199 C7_P_btm.n198 4.60698
R55013 C7_P_btm.n201 C7_P_btm.n200 4.60698
R55014 C7_P_btm.n202 C7_P_btm.n201 4.60698
R55015 C7_P_btm.n204 C7_P_btm.n203 4.60698
R55016 C7_P_btm.n205 C7_P_btm.n204 4.60698
R55017 C7_P_btm.n207 C7_P_btm.n206 4.60698
R55018 C7_P_btm.n208 C7_P_btm.n207 4.60698
R55019 C7_P_btm.n210 C7_P_btm.n209 4.60698
R55020 C7_P_btm.n211 C7_P_btm.n210 4.60698
R55021 C7_P_btm.n213 C7_P_btm.n212 4.60698
R55022 C7_P_btm.n214 C7_P_btm.n213 4.60698
R55023 C7_P_btm.n216 C7_P_btm.n215 4.60698
R55024 C7_P_btm.n217 C7_P_btm.n216 4.60698
R55025 C7_P_btm.n219 C7_P_btm.n218 4.60698
R55026 C7_P_btm.n220 C7_P_btm.n219 4.60698
R55027 C7_P_btm.n222 C7_P_btm.n221 4.60698
R55028 C7_P_btm.n223 C7_P_btm.n222 4.60698
R55029 C7_P_btm.n225 C7_P_btm.n224 4.60698
R55030 C7_P_btm.n226 C7_P_btm.n225 4.60698
R55031 C7_P_btm.n228 C7_P_btm.n227 4.60698
R55032 C7_P_btm.n229 C7_P_btm.n228 4.60698
R55033 C7_P_btm.n231 C7_P_btm.n230 4.60698
R55034 C7_P_btm.n232 C7_P_btm.n231 4.60698
R55035 C7_P_btm.n234 C7_P_btm.n233 4.60698
R55036 C7_P_btm.n235 C7_P_btm.n234 4.60698
R55037 C7_P_btm.n237 C7_P_btm.n236 4.60698
R55038 C7_P_btm.n238 C7_P_btm.n237 4.60698
R55039 C7_P_btm.n145 C7_P_btm.n144 4.60698
R55040 C7_P_btm.n144 C7_P_btm.n143 4.60698
R55041 C7_P_btm.n148 C7_P_btm.n147 4.60698
R55042 C7_P_btm.n147 C7_P_btm.n146 4.60698
R55043 C7_P_btm.n151 C7_P_btm.n150 4.60698
R55044 C7_P_btm.n150 C7_P_btm.n149 4.60698
R55045 C7_P_btm.n154 C7_P_btm.n153 4.60698
R55046 C7_P_btm.n153 C7_P_btm.n152 4.60698
R55047 C7_P_btm.n157 C7_P_btm.n156 4.60698
R55048 C7_P_btm.n156 C7_P_btm.n155 4.60698
R55049 C7_P_btm.n160 C7_P_btm.n159 4.60698
R55050 C7_P_btm.n159 C7_P_btm.n158 4.60698
R55051 C7_P_btm.n163 C7_P_btm.n162 4.60698
R55052 C7_P_btm.n162 C7_P_btm.n161 4.60698
R55053 C7_P_btm.n166 C7_P_btm.n165 4.60698
R55054 C7_P_btm.n165 C7_P_btm.n164 4.60698
R55055 C7_P_btm.n169 C7_P_btm.n168 4.60698
R55056 C7_P_btm.n168 C7_P_btm.n167 4.60698
R55057 C7_P_btm.n172 C7_P_btm.n171 4.60698
R55058 C7_P_btm.n171 C7_P_btm.n170 4.60698
R55059 C7_P_btm.n175 C7_P_btm.n174 4.60698
R55060 C7_P_btm.n174 C7_P_btm.n173 4.60698
R55061 C7_P_btm.n178 C7_P_btm.n177 4.60698
R55062 C7_P_btm.n177 C7_P_btm.n176 4.60698
R55063 C7_P_btm.n181 C7_P_btm.n180 4.60698
R55064 C7_P_btm.n180 C7_P_btm.n179 4.60698
R55065 C7_P_btm.n184 C7_P_btm.n183 4.60698
R55066 C7_P_btm.n183 C7_P_btm.n182 4.60698
R55067 C7_P_btm.n240 C7_P_btm.n239 4.60698
R55068 C7_P_btm.n241 C7_P_btm.n240 4.60698
R55069 C7_P_btm.n247 C7_P_btm.n246 4.60698
R55070 C7_P_btm.n246 C7_P_btm.n245 4.60698
R55071 C7_P_btm.n250 C7_P_btm.n249 4.60698
R55072 C7_P_btm.n249 C7_P_btm.n248 4.60698
R55073 C7_P_btm.n105 C7_P_btm.n104 4.60698
R55074 C7_P_btm.n106 C7_P_btm.n105 4.60698
R55075 C7_P_btm.n108 C7_P_btm.n107 4.60698
R55076 C7_P_btm.n109 C7_P_btm.n108 4.60698
R55077 C7_P_btm.n95 C7_P_btm.n94 4.60698
R55078 C7_P_btm.n94 C7_P_btm.n93 4.60698
R55079 C7_P_btm.n89 C7_P_btm.n88 4.60698
R55080 C7_P_btm.n88 C7_P_btm.n86 4.60698
R55081 C7_P_btm.n80 C7_P_btm.n79 4.60698
R55082 C7_P_btm.n81 C7_P_btm.n80 4.60698
R55083 C7_P_btm.n74 C7_P_btm.n73 4.60698
R55084 C7_P_btm.n73 C7_P_btm.n72 4.60698
R55085 C7_P_btm.n68 C7_P_btm.n67 4.60698
R55086 C7_P_btm.n67 C7_P_btm.n65 4.60698
R55087 C7_P_btm.n59 C7_P_btm.n58 4.60698
R55088 C7_P_btm.n60 C7_P_btm.n59 4.60698
R55089 C7_P_btm.n53 C7_P_btm.n52 4.60698
R55090 C7_P_btm.n52 C7_P_btm.n51 4.60698
R55091 C7_P_btm.n47 C7_P_btm.n46 4.60698
R55092 C7_P_btm.n46 C7_P_btm.n44 4.60698
R55093 C7_P_btm.n39 C7_P_btm.n38 4.60698
R55094 C7_P_btm.n38 C7_P_btm.n37 4.60698
R55095 C7_P_btm.n344 C7_P_btm.t6 4.03712
R55096 C7_P_btm.n342 C7_P_btm.t23 3.98193
R55097 C7_P_btm.n338 C7_P_btm.t60 3.98193
R55098 C7_P_btm.n331 C7_P_btm.t43 3.98193
R55099 C7_P_btm.n324 C7_P_btm.t29 3.98193
R55100 C7_P_btm.n321 C7_P_btm.t134 3.98193
R55101 C7_P_btm.n310 C7_P_btm.t97 3.98193
R55102 C7_P_btm.n303 C7_P_btm.t50 3.98193
R55103 C7_P_btm.n300 C7_P_btm.t38 3.98193
R55104 C7_P_btm.n289 C7_P_btm.t71 3.98193
R55105 C7_P_btm.n282 C7_P_btm.t115 3.98193
R55106 C7_P_btm.n142 C7_P_btm.t45 3.98193
R55107 C7_P_btm.n185 C7_P_btm.t56 3.98193
R55108 C7_P_btm.n242 C7_P_btm.t48 3.98193
R55109 C7_P_btm.n244 C7_P_btm.t9 3.98193
R55110 C7_P_btm.n110 C7_P_btm.t13 3.98193
R55111 C7_P_btm.n92 C7_P_btm.t98 3.98193
R55112 C7_P_btm.n85 C7_P_btm.t101 3.98193
R55113 C7_P_btm.n82 C7_P_btm.t113 3.98193
R55114 C7_P_btm.n71 C7_P_btm.t67 3.98193
R55115 C7_P_btm.n64 C7_P_btm.t78 3.98193
R55116 C7_P_btm.n61 C7_P_btm.t90 3.98193
R55117 C7_P_btm.n50 C7_P_btm.t68 3.98193
R55118 C7_P_btm.n43 C7_P_btm.t130 3.98193
R55119 C7_P_btm.n40 C7_P_btm.t27 3.98193
R55120 C7_P_btm.n36 C7_P_btm.t36 3.98193
R55121 C7_P_btm.n45 C7_P_btm.t66 3.98193
R55122 C7_P_btm.n54 C7_P_btm.t126 3.98193
R55123 C7_P_btm.n57 C7_P_btm.t100 3.98193
R55124 C7_P_btm.n66 C7_P_btm.t87 3.98193
R55125 C7_P_btm.n75 C7_P_btm.t76 3.98193
R55126 C7_P_btm.n78 C7_P_btm.t121 3.98193
R55127 C7_P_btm.n87 C7_P_btm.t111 3.98193
R55128 C7_P_btm.n96 C7_P_btm.t35 3.98193
R55129 C7_P_btm.n21 C7_P_btm.t77 3.98193
R55130 C7_P_btm.n271 C7_P_btm.t127 3.98193
R55131 C7_P_btm.n274 C7_P_btm.t63 3.98193
R55132 C7_P_btm.n284 C7_P_btm.t128 3.98193
R55133 C7_P_btm.n293 C7_P_btm.t69 3.98193
R55134 C7_P_btm.n296 C7_P_btm.t39 3.98193
R55135 C7_P_btm.n305 C7_P_btm.t112 3.98193
R55136 C7_P_btm.n314 C7_P_btm.t10 3.98193
R55137 C7_P_btm.n317 C7_P_btm.t15 3.98193
R55138 C7_P_btm.n326 C7_P_btm.t89 3.98193
R55139 C7_P_btm.n335 C7_P_btm.t103 3.98193
R55140 C7_P_btm.n103 C7_P_btm.t107 3.92851
R55141 C7_P_btm.n102 C7_P_btm.t30 3.92851
R55142 C7_P_btm.n101 C7_P_btm.t129 3.92851
R55143 C7_P_btm.n100 C7_P_btm.t37 3.92851
R55144 C7_P_btm.n99 C7_P_btm.t65 3.92851
R55145 C7_P_btm.n251 C7_P_btm.t93 3.92851
R55146 C7_P_btm.n252 C7_P_btm.t16 3.92851
R55147 C7_P_btm.n253 C7_P_btm.t109 3.92851
R55148 C7_P_btm.n254 C7_P_btm.t57 3.92851
R55149 C7_P_btm.n255 C7_P_btm.t116 3.92851
R55150 C7_P_btm.n256 C7_P_btm.t85 3.92851
R55151 C7_P_btm.n257 C7_P_btm.t21 3.92851
R55152 C7_P_btm.n258 C7_P_btm.t91 3.92851
R55153 C7_P_btm.n259 C7_P_btm.t64 3.92851
R55154 C7_P_btm.n260 C7_P_btm.t106 3.92851
R55155 C7_P_btm.n261 C7_P_btm.t72 3.92851
R55156 C7_P_btm.n262 C7_P_btm.t114 3.92851
R55157 C7_P_btm.n263 C7_P_btm.t83 3.92851
R55158 C7_P_btm.n264 C7_P_btm.t80 3.92851
R55159 C7_P_btm.n19 C7_P_btm.t61 3.92851
R55160 C7_P_btm.n18 C7_P_btm.t95 3.92851
R55161 C7_P_btm.n17 C7_P_btm.t62 3.92851
R55162 C7_P_btm.n16 C7_P_btm.t81 3.92851
R55163 C7_P_btm.n15 C7_P_btm.t47 3.92851
R55164 C7_P_btm.n0 C7_P_btm.t2 3.57113
R55165 C7_P_btm.n0 C7_P_btm.t1 3.57113
R55166 C7_P_btm.n340 C7_P_btm.t86 1.67819
R55167 C7_P_btm.n333 C7_P_btm.t12 1.67819
R55168 C7_P_btm.n327 C7_P_btm.t54 1.67819
R55169 C7_P_btm.n319 C7_P_btm.t125 1.67819
R55170 C7_P_btm.n312 C7_P_btm.t33 1.67819
R55171 C7_P_btm.n306 C7_P_btm.t25 1.67819
R55172 C7_P_btm.n298 C7_P_btm.t58 1.67819
R55173 C7_P_btm.n291 C7_P_btm.t55 1.67819
R55174 C7_P_btm.n285 C7_P_btm.t84 1.67819
R55175 C7_P_btm.n276 C7_P_btm.t74 1.67819
R55176 C7_P_btm.n278 C7_P_btm.t102 1.67819
R55177 C7_P_btm.n266 C7_P_btm.t88 1.67819
R55178 C7_P_btm.n269 C7_P_btm.t135 1.67819
R55179 C7_P_btm.n189 C7_P_btm.t108 1.67819
R55180 C7_P_btm.n192 C7_P_btm.t14 1.67819
R55181 C7_P_btm.n195 C7_P_btm.t92 1.67819
R55182 C7_P_btm.n198 C7_P_btm.t53 1.67819
R55183 C7_P_btm.n201 C7_P_btm.t40 1.67819
R55184 C7_P_btm.n204 C7_P_btm.t44 1.67819
R55185 C7_P_btm.n207 C7_P_btm.t32 1.67819
R55186 C7_P_btm.n210 C7_P_btm.t110 1.67819
R55187 C7_P_btm.n213 C7_P_btm.t17 1.67819
R55188 C7_P_btm.n216 C7_P_btm.t132 1.67819
R55189 C7_P_btm.n219 C7_P_btm.t120 1.67819
R55190 C7_P_btm.n222 C7_P_btm.t42 1.67819
R55191 C7_P_btm.n225 C7_P_btm.t59 1.67819
R55192 C7_P_btm.n228 C7_P_btm.t34 1.67819
R55193 C7_P_btm.n231 C7_P_btm.t117 1.67819
R55194 C7_P_btm.n234 C7_P_btm.t24 1.67819
R55195 C7_P_btm.n237 C7_P_btm.t133 1.67819
R55196 C7_P_btm.n144 C7_P_btm.t18 1.67819
R55197 C7_P_btm.n147 C7_P_btm.t51 1.67819
R55198 C7_P_btm.n150 C7_P_btm.t49 1.67819
R55199 C7_P_btm.n153 C7_P_btm.t136 1.67819
R55200 C7_P_btm.n156 C7_P_btm.t28 1.67819
R55201 C7_P_btm.n159 C7_P_btm.t22 1.67819
R55202 C7_P_btm.n162 C7_P_btm.t123 1.67819
R55203 C7_P_btm.n165 C7_P_btm.t11 1.67819
R55204 C7_P_btm.n168 C7_P_btm.t96 1.67819
R55205 C7_P_btm.n171 C7_P_btm.t20 1.67819
R55206 C7_P_btm.n174 C7_P_btm.t104 1.67819
R55207 C7_P_btm.n177 C7_P_btm.t119 1.67819
R55208 C7_P_btm.n180 C7_P_btm.t46 1.67819
R55209 C7_P_btm.n183 C7_P_btm.t79 1.67819
R55210 C7_P_btm.n240 C7_P_btm.t73 1.67819
R55211 C7_P_btm.n246 C7_P_btm.t41 1.67819
R55212 C7_P_btm.n249 C7_P_btm.t70 1.67819
R55213 C7_P_btm.n105 C7_P_btm.t52 1.67819
R55214 C7_P_btm.n108 C7_P_btm.t131 1.67819
R55215 C7_P_btm.n94 C7_P_btm.t118 1.67819
R55216 C7_P_btm.n88 C7_P_btm.t19 1.67819
R55217 C7_P_btm.n80 C7_P_btm.t31 1.67819
R55218 C7_P_btm.n73 C7_P_btm.t105 1.67819
R55219 C7_P_btm.n67 C7_P_btm.t122 1.67819
R55220 C7_P_btm.n59 C7_P_btm.t26 1.67819
R55221 C7_P_btm.n52 C7_P_btm.t82 1.67819
R55222 C7_P_btm.n46 C7_P_btm.t94 1.67819
R55223 C7_P_btm.n38 C7_P_btm.t124 1.67819
R55224 C7_P_btm.n186 C7_P_btm.n185 1.05569
R55225 C7_P_btm.n142 C7_P_btm.n113 1.05569
R55226 C7_P_btm.n243 C7_P_btm.n242 1.05569
R55227 C7_P_btm.n272 C7_P_btm.n21 1.05569
R55228 C7_P_btm.n330 C7_P_btm.n5 1.0005
R55229 C7_P_btm.n330 C7_P_btm.n329 1.0005
R55230 C7_P_btm.n329 C7_P_btm.n7 1.0005
R55231 C7_P_btm.n309 C7_P_btm.n7 1.0005
R55232 C7_P_btm.n309 C7_P_btm.n308 1.0005
R55233 C7_P_btm.n308 C7_P_btm.n10 1.0005
R55234 C7_P_btm.n288 C7_P_btm.n10 1.0005
R55235 C7_P_btm.n288 C7_P_btm.n287 1.0005
R55236 C7_P_btm.n287 C7_P_btm.n13 1.0005
R55237 C7_P_btm.n22 C7_P_btm.n13 1.0005
R55238 C7_P_btm.n187 C7_P_btm.n22 1.0005
R55239 C7_P_btm.n186 C7_P_btm.n14 1.0005
R55240 C7_P_btm.n141 C7_P_btm.n114 1.0005
R55241 C7_P_btm.n140 C7_P_btm.n115 1.0005
R55242 C7_P_btm.n139 C7_P_btm.n116 1.0005
R55243 C7_P_btm.n138 C7_P_btm.n117 1.0005
R55244 C7_P_btm.n137 C7_P_btm.n118 1.0005
R55245 C7_P_btm.n136 C7_P_btm.n119 1.0005
R55246 C7_P_btm.n135 C7_P_btm.n120 1.0005
R55247 C7_P_btm.n134 C7_P_btm.n121 1.0005
R55248 C7_P_btm.n133 C7_P_btm.n122 1.0005
R55249 C7_P_btm.n132 C7_P_btm.n123 1.0005
R55250 C7_P_btm.n131 C7_P_btm.n124 1.0005
R55251 C7_P_btm.n130 C7_P_btm.n125 1.0005
R55252 C7_P_btm.n129 C7_P_btm.n126 1.0005
R55253 C7_P_btm.n128 C7_P_btm.n127 1.0005
R55254 C7_P_btm.n112 C7_P_btm.n24 1.0005
R55255 C7_P_btm.n26 C7_P_btm.n24 1.0005
R55256 C7_P_btm.n91 C7_P_btm.n26 1.0005
R55257 C7_P_btm.n91 C7_P_btm.n90 1.0005
R55258 C7_P_btm.n90 C7_P_btm.n28 1.0005
R55259 C7_P_btm.n70 C7_P_btm.n28 1.0005
R55260 C7_P_btm.n70 C7_P_btm.n69 1.0005
R55261 C7_P_btm.n69 C7_P_btm.n31 1.0005
R55262 C7_P_btm.n49 C7_P_btm.n31 1.0005
R55263 C7_P_btm.n49 C7_P_btm.n48 1.0005
R55264 C7_P_btm.n48 C7_P_btm.n34 1.0005
R55265 C7_P_btm.n35 C7_P_btm.n33 1.0005
R55266 C7_P_btm.n42 C7_P_btm.n32 1.0005
R55267 C7_P_btm.n42 C7_P_btm.n41 1.0005
R55268 C7_P_btm.n56 C7_P_btm.n55 1.0005
R55269 C7_P_btm.n55 C7_P_btm.n33 1.0005
R55270 C7_P_btm.n63 C7_P_btm.n62 1.0005
R55271 C7_P_btm.n62 C7_P_btm.n32 1.0005
R55272 C7_P_btm.n76 C7_P_btm.n30 1.0005
R55273 C7_P_btm.n56 C7_P_btm.n30 1.0005
R55274 C7_P_btm.n83 C7_P_btm.n29 1.0005
R55275 C7_P_btm.n63 C7_P_btm.n29 1.0005
R55276 C7_P_btm.n77 C7_P_btm.n27 1.0005
R55277 C7_P_btm.n77 C7_P_btm.n76 1.0005
R55278 C7_P_btm.n84 C7_P_btm.n25 1.0005
R55279 C7_P_btm.n84 C7_P_btm.n83 1.0005
R55280 C7_P_btm.n98 C7_P_btm.n97 1.0005
R55281 C7_P_btm.n97 C7_P_btm.n27 1.0005
R55282 C7_P_btm.n243 C7_P_btm.n111 1.0005
R55283 C7_P_btm.n111 C7_P_btm.n25 1.0005
R55284 C7_P_btm.n113 C7_P_btm.n23 1.0005
R55285 C7_P_btm.n98 C7_P_btm.n23 1.0005
R55286 C7_P_btm.n273 C7_P_btm.n272 1.0005
R55287 C7_P_btm.n280 C7_P_btm.n14 1.0005
R55288 C7_P_btm.n281 C7_P_btm.n280 1.0005
R55289 C7_P_btm.n273 C7_P_btm.n12 1.0005
R55290 C7_P_btm.n294 C7_P_btm.n12 1.0005
R55291 C7_P_btm.n281 C7_P_btm.n11 1.0005
R55292 C7_P_btm.n301 C7_P_btm.n11 1.0005
R55293 C7_P_btm.n295 C7_P_btm.n294 1.0005
R55294 C7_P_btm.n295 C7_P_btm.n9 1.0005
R55295 C7_P_btm.n302 C7_P_btm.n301 1.0005
R55296 C7_P_btm.n302 C7_P_btm.n8 1.0005
R55297 C7_P_btm.n315 C7_P_btm.n9 1.0005
R55298 C7_P_btm.n316 C7_P_btm.n315 1.0005
R55299 C7_P_btm.n322 C7_P_btm.n8 1.0005
R55300 C7_P_btm.n323 C7_P_btm.n322 1.0005
R55301 C7_P_btm.n316 C7_P_btm.n6 1.0005
R55302 C7_P_btm.n336 C7_P_btm.n6 1.0005
R55303 C7_P_btm.n323 C7_P_btm.n4 1.0005
R55304 C7_P_btm.n343 C7_P_btm.n4 1.0005
R55305 C7_P_btm.n337 C7_P_btm.n336 1.0005
R55306 C7_P_btm.n344 C7_P_btm.n343 1.0005
R55307 C7_P_btm.n100 C7_P_btm.n99 0.840176
R55308 C7_P_btm.n101 C7_P_btm.n100 0.840176
R55309 C7_P_btm.n102 C7_P_btm.n101 0.840176
R55310 C7_P_btm.n103 C7_P_btm.n102 0.840176
R55311 C7_P_btm.n264 C7_P_btm.n263 0.840176
R55312 C7_P_btm.n263 C7_P_btm.n262 0.840176
R55313 C7_P_btm.n262 C7_P_btm.n261 0.840176
R55314 C7_P_btm.n261 C7_P_btm.n260 0.840176
R55315 C7_P_btm.n260 C7_P_btm.n259 0.840176
R55316 C7_P_btm.n259 C7_P_btm.n258 0.840176
R55317 C7_P_btm.n258 C7_P_btm.n257 0.840176
R55318 C7_P_btm.n257 C7_P_btm.n256 0.840176
R55319 C7_P_btm.n256 C7_P_btm.n255 0.840176
R55320 C7_P_btm.n255 C7_P_btm.n254 0.840176
R55321 C7_P_btm.n254 C7_P_btm.n253 0.840176
R55322 C7_P_btm.n253 C7_P_btm.n252 0.840176
R55323 C7_P_btm.n252 C7_P_btm.n251 0.840176
R55324 C7_P_btm.n16 C7_P_btm.n15 0.840176
R55325 C7_P_btm.n17 C7_P_btm.n16 0.840176
R55326 C7_P_btm.n18 C7_P_btm.n17 0.840176
R55327 C7_P_btm.n19 C7_P_btm.n18 0.840176
R55328 C7_P_btm.n104 C7_P_btm.n103 0.732838
R55329 C7_P_btm.n265 C7_P_btm.n264 0.732838
R55330 C7_P_btm.n251 C7_P_btm.n250 0.732838
R55331 C7_P_btm.n20 C7_P_btm.n19 0.732838
R55332 C7_P_btm.n185 C7_P_btm.n184 0.679419
R55333 C7_P_btm.n143 C7_P_btm.n142 0.679419
R55334 C7_P_btm.n37 C7_P_btm.n36 0.679419
R55335 C7_P_btm.n40 C7_P_btm.n39 0.679419
R55336 C7_P_btm.n44 C7_P_btm.n43 0.679419
R55337 C7_P_btm.n47 C7_P_btm.n45 0.679419
R55338 C7_P_btm.n54 C7_P_btm.n53 0.679419
R55339 C7_P_btm.n51 C7_P_btm.n50 0.679419
R55340 C7_P_btm.n61 C7_P_btm.n60 0.679419
R55341 C7_P_btm.n58 C7_P_btm.n57 0.679419
R55342 C7_P_btm.n68 C7_P_btm.n66 0.679419
R55343 C7_P_btm.n65 C7_P_btm.n64 0.679419
R55344 C7_P_btm.n72 C7_P_btm.n71 0.679419
R55345 C7_P_btm.n75 C7_P_btm.n74 0.679419
R55346 C7_P_btm.n79 C7_P_btm.n78 0.679419
R55347 C7_P_btm.n82 C7_P_btm.n81 0.679419
R55348 C7_P_btm.n86 C7_P_btm.n85 0.679419
R55349 C7_P_btm.n89 C7_P_btm.n87 0.679419
R55350 C7_P_btm.n96 C7_P_btm.n95 0.679419
R55351 C7_P_btm.n93 C7_P_btm.n92 0.679419
R55352 C7_P_btm.n110 C7_P_btm.n109 0.679419
R55353 C7_P_btm.n245 C7_P_btm.n244 0.679419
R55354 C7_P_btm.n242 C7_P_btm.n241 0.679419
R55355 C7_P_btm.n188 C7_P_btm.n21 0.679419
R55356 C7_P_btm.n271 C7_P_btm.n270 0.679419
R55357 C7_P_btm.n275 C7_P_btm.n274 0.679419
R55358 C7_P_btm.n286 C7_P_btm.n284 0.679419
R55359 C7_P_btm.n283 C7_P_btm.n282 0.679419
R55360 C7_P_btm.n290 C7_P_btm.n289 0.679419
R55361 C7_P_btm.n293 C7_P_btm.n292 0.679419
R55362 C7_P_btm.n297 C7_P_btm.n296 0.679419
R55363 C7_P_btm.n300 C7_P_btm.n299 0.679419
R55364 C7_P_btm.n304 C7_P_btm.n303 0.679419
R55365 C7_P_btm.n307 C7_P_btm.n305 0.679419
R55366 C7_P_btm.n314 C7_P_btm.n313 0.679419
R55367 C7_P_btm.n311 C7_P_btm.n310 0.679419
R55368 C7_P_btm.n321 C7_P_btm.n320 0.679419
R55369 C7_P_btm.n318 C7_P_btm.n317 0.679419
R55370 C7_P_btm.n328 C7_P_btm.n326 0.679419
R55371 C7_P_btm.n325 C7_P_btm.n324 0.679419
R55372 C7_P_btm.n332 C7_P_btm.n331 0.679419
R55373 C7_P_btm.n335 C7_P_btm.n334 0.679419
R55374 C7_P_btm.n339 C7_P_btm.n338 0.679419
R55375 C7_P_btm.n342 C7_P_btm.n341 0.679419
R55376 C7_P_btm.n182 C7_P_btm.n181 0.6255
R55377 C7_P_btm.n179 C7_P_btm.n178 0.6255
R55378 C7_P_btm.n176 C7_P_btm.n175 0.6255
R55379 C7_P_btm.n173 C7_P_btm.n172 0.6255
R55380 C7_P_btm.n170 C7_P_btm.n169 0.6255
R55381 C7_P_btm.n167 C7_P_btm.n166 0.6255
R55382 C7_P_btm.n164 C7_P_btm.n163 0.6255
R55383 C7_P_btm.n161 C7_P_btm.n160 0.6255
R55384 C7_P_btm.n158 C7_P_btm.n157 0.6255
R55385 C7_P_btm.n155 C7_P_btm.n154 0.6255
R55386 C7_P_btm.n152 C7_P_btm.n151 0.6255
R55387 C7_P_btm.n149 C7_P_btm.n148 0.6255
R55388 C7_P_btm.n146 C7_P_btm.n145 0.6255
R55389 C7_P_btm.n107 C7_P_btm.n106 0.6255
R55390 C7_P_btm.n248 C7_P_btm.n247 0.6255
R55391 C7_P_btm.n239 C7_P_btm.n238 0.6255
R55392 C7_P_btm.n236 C7_P_btm.n235 0.6255
R55393 C7_P_btm.n233 C7_P_btm.n232 0.6255
R55394 C7_P_btm.n230 C7_P_btm.n229 0.6255
R55395 C7_P_btm.n227 C7_P_btm.n226 0.6255
R55396 C7_P_btm.n224 C7_P_btm.n223 0.6255
R55397 C7_P_btm.n221 C7_P_btm.n220 0.6255
R55398 C7_P_btm.n218 C7_P_btm.n217 0.6255
R55399 C7_P_btm.n215 C7_P_btm.n214 0.6255
R55400 C7_P_btm.n212 C7_P_btm.n211 0.6255
R55401 C7_P_btm.n209 C7_P_btm.n208 0.6255
R55402 C7_P_btm.n206 C7_P_btm.n205 0.6255
R55403 C7_P_btm.n203 C7_P_btm.n202 0.6255
R55404 C7_P_btm.n200 C7_P_btm.n199 0.6255
R55405 C7_P_btm.n197 C7_P_btm.n196 0.6255
R55406 C7_P_btm.n194 C7_P_btm.n193 0.6255
R55407 C7_P_btm.n191 C7_P_btm.n190 0.6255
R55408 C7_P_btm.n268 C7_P_btm.n267 0.6255
R55409 C7_P_btm.n279 C7_P_btm.n277 0.6255
R55410 C7_P_btm.n182 C7_P_btm.n128 0.109875
R55411 C7_P_btm.n184 C7_P_btm.n128 0.109875
R55412 C7_P_btm.n179 C7_P_btm.n129 0.109875
R55413 C7_P_btm.n181 C7_P_btm.n129 0.109875
R55414 C7_P_btm.n176 C7_P_btm.n130 0.109875
R55415 C7_P_btm.n178 C7_P_btm.n130 0.109875
R55416 C7_P_btm.n173 C7_P_btm.n131 0.109875
R55417 C7_P_btm.n175 C7_P_btm.n131 0.109875
R55418 C7_P_btm.n170 C7_P_btm.n132 0.109875
R55419 C7_P_btm.n172 C7_P_btm.n132 0.109875
R55420 C7_P_btm.n167 C7_P_btm.n133 0.109875
R55421 C7_P_btm.n169 C7_P_btm.n133 0.109875
R55422 C7_P_btm.n164 C7_P_btm.n134 0.109875
R55423 C7_P_btm.n166 C7_P_btm.n134 0.109875
R55424 C7_P_btm.n161 C7_P_btm.n135 0.109875
R55425 C7_P_btm.n163 C7_P_btm.n135 0.109875
R55426 C7_P_btm.n158 C7_P_btm.n136 0.109875
R55427 C7_P_btm.n160 C7_P_btm.n136 0.109875
R55428 C7_P_btm.n155 C7_P_btm.n137 0.109875
R55429 C7_P_btm.n157 C7_P_btm.n137 0.109875
R55430 C7_P_btm.n152 C7_P_btm.n138 0.109875
R55431 C7_P_btm.n154 C7_P_btm.n138 0.109875
R55432 C7_P_btm.n149 C7_P_btm.n139 0.109875
R55433 C7_P_btm.n151 C7_P_btm.n139 0.109875
R55434 C7_P_btm.n146 C7_P_btm.n140 0.109875
R55435 C7_P_btm.n148 C7_P_btm.n140 0.109875
R55436 C7_P_btm.n143 C7_P_btm.n141 0.109875
R55437 C7_P_btm.n145 C7_P_btm.n141 0.109875
R55438 C7_P_btm.n39 C7_P_btm.n34 0.109875
R55439 C7_P_btm.n37 C7_P_btm.n34 0.109875
R55440 C7_P_btm.n48 C7_P_btm.n44 0.109875
R55441 C7_P_btm.n48 C7_P_btm.n47 0.109875
R55442 C7_P_btm.n51 C7_P_btm.n49 0.109875
R55443 C7_P_btm.n53 C7_P_btm.n49 0.109875
R55444 C7_P_btm.n60 C7_P_btm.n31 0.109875
R55445 C7_P_btm.n58 C7_P_btm.n31 0.109875
R55446 C7_P_btm.n69 C7_P_btm.n65 0.109875
R55447 C7_P_btm.n69 C7_P_btm.n68 0.109875
R55448 C7_P_btm.n72 C7_P_btm.n70 0.109875
R55449 C7_P_btm.n74 C7_P_btm.n70 0.109875
R55450 C7_P_btm.n81 C7_P_btm.n28 0.109875
R55451 C7_P_btm.n79 C7_P_btm.n28 0.109875
R55452 C7_P_btm.n90 C7_P_btm.n86 0.109875
R55453 C7_P_btm.n90 C7_P_btm.n89 0.109875
R55454 C7_P_btm.n93 C7_P_btm.n91 0.109875
R55455 C7_P_btm.n95 C7_P_btm.n91 0.109875
R55456 C7_P_btm.n109 C7_P_btm.n26 0.109875
R55457 C7_P_btm.n107 C7_P_btm.n26 0.109875
R55458 C7_P_btm.n106 C7_P_btm.n98 0.109875
R55459 C7_P_btm.n104 C7_P_btm.n98 0.109875
R55460 C7_P_btm.n248 C7_P_btm.n23 0.109875
R55461 C7_P_btm.n250 C7_P_btm.n23 0.109875
R55462 C7_P_btm.n245 C7_P_btm.n24 0.109875
R55463 C7_P_btm.n247 C7_P_btm.n24 0.109875
R55464 C7_P_btm.n241 C7_P_btm.n112 0.109875
R55465 C7_P_btm.n239 C7_P_btm.n112 0.109875
R55466 C7_P_btm.n238 C7_P_btm.n113 0.109875
R55467 C7_P_btm.n236 C7_P_btm.n113 0.109875
R55468 C7_P_btm.n235 C7_P_btm.n114 0.109875
R55469 C7_P_btm.n233 C7_P_btm.n114 0.109875
R55470 C7_P_btm.n232 C7_P_btm.n115 0.109875
R55471 C7_P_btm.n230 C7_P_btm.n115 0.109875
R55472 C7_P_btm.n229 C7_P_btm.n116 0.109875
R55473 C7_P_btm.n227 C7_P_btm.n116 0.109875
R55474 C7_P_btm.n226 C7_P_btm.n117 0.109875
R55475 C7_P_btm.n224 C7_P_btm.n117 0.109875
R55476 C7_P_btm.n223 C7_P_btm.n118 0.109875
R55477 C7_P_btm.n221 C7_P_btm.n118 0.109875
R55478 C7_P_btm.n220 C7_P_btm.n119 0.109875
R55479 C7_P_btm.n218 C7_P_btm.n119 0.109875
R55480 C7_P_btm.n217 C7_P_btm.n120 0.109875
R55481 C7_P_btm.n215 C7_P_btm.n120 0.109875
R55482 C7_P_btm.n214 C7_P_btm.n121 0.109875
R55483 C7_P_btm.n212 C7_P_btm.n121 0.109875
R55484 C7_P_btm.n211 C7_P_btm.n122 0.109875
R55485 C7_P_btm.n209 C7_P_btm.n122 0.109875
R55486 C7_P_btm.n208 C7_P_btm.n123 0.109875
R55487 C7_P_btm.n206 C7_P_btm.n123 0.109875
R55488 C7_P_btm.n205 C7_P_btm.n124 0.109875
R55489 C7_P_btm.n203 C7_P_btm.n124 0.109875
R55490 C7_P_btm.n202 C7_P_btm.n125 0.109875
R55491 C7_P_btm.n200 C7_P_btm.n125 0.109875
R55492 C7_P_btm.n199 C7_P_btm.n126 0.109875
R55493 C7_P_btm.n197 C7_P_btm.n126 0.109875
R55494 C7_P_btm.n196 C7_P_btm.n127 0.109875
R55495 C7_P_btm.n194 C7_P_btm.n127 0.109875
R55496 C7_P_btm.n193 C7_P_btm.n186 0.109875
R55497 C7_P_btm.n191 C7_P_btm.n186 0.109875
R55498 C7_P_btm.n190 C7_P_btm.n187 0.109875
R55499 C7_P_btm.n188 C7_P_btm.n187 0.109875
R55500 C7_P_btm.n268 C7_P_btm.n22 0.109875
R55501 C7_P_btm.n270 C7_P_btm.n22 0.109875
R55502 C7_P_btm.n265 C7_P_btm.n14 0.109875
R55503 C7_P_btm.n267 C7_P_btm.n14 0.109875
R55504 C7_P_btm.n280 C7_P_btm.n20 0.109875
R55505 C7_P_btm.n280 C7_P_btm.n279 0.109875
R55506 C7_P_btm.n277 C7_P_btm.n13 0.109875
R55507 C7_P_btm.n275 C7_P_btm.n13 0.109875
R55508 C7_P_btm.n287 C7_P_btm.n283 0.109875
R55509 C7_P_btm.n287 C7_P_btm.n286 0.109875
R55510 C7_P_btm.n290 C7_P_btm.n288 0.109875
R55511 C7_P_btm.n292 C7_P_btm.n288 0.109875
R55512 C7_P_btm.n299 C7_P_btm.n10 0.109875
R55513 C7_P_btm.n297 C7_P_btm.n10 0.109875
R55514 C7_P_btm.n308 C7_P_btm.n304 0.109875
R55515 C7_P_btm.n308 C7_P_btm.n307 0.109875
R55516 C7_P_btm.n311 C7_P_btm.n309 0.109875
R55517 C7_P_btm.n313 C7_P_btm.n309 0.109875
R55518 C7_P_btm.n320 C7_P_btm.n7 0.109875
R55519 C7_P_btm.n318 C7_P_btm.n7 0.109875
R55520 C7_P_btm.n329 C7_P_btm.n325 0.109875
R55521 C7_P_btm.n329 C7_P_btm.n328 0.109875
R55522 C7_P_btm.n332 C7_P_btm.n330 0.109875
R55523 C7_P_btm.n334 C7_P_btm.n330 0.109875
R55524 C7_P_btm.n341 C7_P_btm.n5 0.109875
R55525 C7_P_btm.n339 C7_P_btm.n5 0.109875
R55526 C7_P_btm.n36 C7_P_btm.n35 0.0556875
R55527 C7_P_btm.n41 C7_P_btm.n40 0.0556875
R55528 C7_P_btm.n43 C7_P_btm.n42 0.0556875
R55529 C7_P_btm.n45 C7_P_btm.n33 0.0556875
R55530 C7_P_btm.n55 C7_P_btm.n54 0.0556875
R55531 C7_P_btm.n50 C7_P_btm.n32 0.0556875
R55532 C7_P_btm.n62 C7_P_btm.n61 0.0556875
R55533 C7_P_btm.n57 C7_P_btm.n56 0.0556875
R55534 C7_P_btm.n66 C7_P_btm.n30 0.0556875
R55535 C7_P_btm.n64 C7_P_btm.n63 0.0556875
R55536 C7_P_btm.n71 C7_P_btm.n29 0.0556875
R55537 C7_P_btm.n76 C7_P_btm.n75 0.0556875
R55538 C7_P_btm.n78 C7_P_btm.n77 0.0556875
R55539 C7_P_btm.n83 C7_P_btm.n82 0.0556875
R55540 C7_P_btm.n85 C7_P_btm.n84 0.0556875
R55541 C7_P_btm.n87 C7_P_btm.n27 0.0556875
R55542 C7_P_btm.n97 C7_P_btm.n96 0.0556875
R55543 C7_P_btm.n92 C7_P_btm.n25 0.0556875
R55544 C7_P_btm.n111 C7_P_btm.n110 0.0556875
R55545 C7_P_btm.n244 C7_P_btm.n243 0.0556875
R55546 C7_P_btm.n272 C7_P_btm.n271 0.0556875
R55547 C7_P_btm.n274 C7_P_btm.n273 0.0556875
R55548 C7_P_btm.n284 C7_P_btm.n12 0.0556875
R55549 C7_P_btm.n282 C7_P_btm.n281 0.0556875
R55550 C7_P_btm.n289 C7_P_btm.n11 0.0556875
R55551 C7_P_btm.n294 C7_P_btm.n293 0.0556875
R55552 C7_P_btm.n296 C7_P_btm.n295 0.0556875
R55553 C7_P_btm.n301 C7_P_btm.n300 0.0556875
R55554 C7_P_btm.n303 C7_P_btm.n302 0.0556875
R55555 C7_P_btm.n305 C7_P_btm.n9 0.0556875
R55556 C7_P_btm.n315 C7_P_btm.n314 0.0556875
R55557 C7_P_btm.n310 C7_P_btm.n8 0.0556875
R55558 C7_P_btm.n322 C7_P_btm.n321 0.0556875
R55559 C7_P_btm.n317 C7_P_btm.n316 0.0556875
R55560 C7_P_btm.n326 C7_P_btm.n6 0.0556875
R55561 C7_P_btm.n324 C7_P_btm.n323 0.0556875
R55562 C7_P_btm.n331 C7_P_btm.n4 0.0556875
R55563 C7_P_btm.n336 C7_P_btm.n335 0.0556875
R55564 C7_P_btm.n338 C7_P_btm.n337 0.0556875
R55565 C7_P_btm.n343 C7_P_btm.n342 0.0556875
R55566 a_20892_30659.n1 a_20892_30659.t4 868.625
R55567 a_20892_30659.n1 a_20892_30659.n0 380.32
R55568 a_20892_30659.n2 a_20892_30659.n1 185
R55569 a_20892_30659.n0 a_20892_30659.t3 26.5955
R55570 a_20892_30659.n0 a_20892_30659.t2 26.5955
R55571 a_20892_30659.n2 a_20892_30659.t0 24.9236
R55572 a_20892_30659.t1 a_20892_30659.n2 24.9236
R55573 a_n1551_45412.n2 a_n1551_45412.n0 329.507
R55574 a_n1551_45412.n6 a_n1551_45412.n5 305.616
R55575 a_n1551_45412.n9 a_n1551_45412.n8 300.118
R55576 a_n1551_45412.n2 a_n1551_45412.n1 299.834
R55577 a_n1551_45412.n10 a_n1551_45412.n9 291.81
R55578 a_n1551_45412.n3 a_n1551_45412.t10 276.464
R55579 a_n1551_45412.n5 a_n1551_45412.t12 212.081
R55580 a_n1551_45412.n4 a_n1551_45412.t11 212.081
R55581 a_n1551_45412.n6 a_n1551_45412.n3 205.322
R55582 a_n1551_45412.n3 a_n1551_45412.t13 196.131
R55583 a_n1551_45412.n5 a_n1551_45412.t9 139.78
R55584 a_n1551_45412.n4 a_n1551_45412.t8 139.78
R55585 a_n1551_45412.n5 a_n1551_45412.n4 61.346
R55586 a_n1551_45412.n9 a_n1551_45412.n7 56.2452
R55587 a_n1551_45412.n8 a_n1551_45412.t2 26.5955
R55588 a_n1551_45412.n8 a_n1551_45412.t3 26.5955
R55589 a_n1551_45412.n1 a_n1551_45412.t6 26.5955
R55590 a_n1551_45412.n1 a_n1551_45412.t7 26.5955
R55591 a_n1551_45412.n0 a_n1551_45412.t5 26.5955
R55592 a_n1551_45412.n0 a_n1551_45412.t4 26.5955
R55593 a_n1551_45412.n10 a_n1551_45412.t0 24.9236
R55594 a_n1551_45412.t1 a_n1551_45412.n10 24.9236
R55595 a_n1551_45412.n7 a_n1551_45412.n2 23.5584
R55596 a_n1551_45412.n7 a_n1551_45412.n6 10.8268
R55597 a_n1735_43236.n10 a_n1735_43236.n9 312.635
R55598 a_n1735_43236.n8 a_n1735_43236.n5 304.618
R55599 a_n1735_43236.n2 a_n1735_43236.n1 300.118
R55600 a_n1735_43236.n4 a_n1735_43236.n3 299.834
R55601 a_n1735_43236.n2 a_n1735_43236.n0 291.81
R55602 a_n1735_43236.n5 a_n1735_43236.t13 276.464
R55603 a_n1735_43236.n8 a_n1735_43236.n7 225.791
R55604 a_n1735_43236.n7 a_n1735_43236.t8 212.081
R55605 a_n1735_43236.n6 a_n1735_43236.t11 212.081
R55606 a_n1735_43236.n5 a_n1735_43236.t9 196.131
R55607 a_n1735_43236.n7 a_n1735_43236.t12 139.78
R55608 a_n1735_43236.n6 a_n1735_43236.t10 139.78
R55609 a_n1735_43236.n4 a_n1735_43236.n2 79.8031
R55610 a_n1735_43236.n7 a_n1735_43236.n6 61.346
R55611 a_n1735_43236.n3 a_n1735_43236.t2 26.5955
R55612 a_n1735_43236.n3 a_n1735_43236.t3 26.5955
R55613 a_n1735_43236.n1 a_n1735_43236.t6 26.5955
R55614 a_n1735_43236.n1 a_n1735_43236.t7 26.5955
R55615 a_n1735_43236.n10 a_n1735_43236.t1 26.5955
R55616 a_n1735_43236.t0 a_n1735_43236.n10 26.5955
R55617 a_n1735_43236.n0 a_n1735_43236.t5 24.9236
R55618 a_n1735_43236.n0 a_n1735_43236.t4 24.9236
R55619 a_n1735_43236.n9 a_n1735_43236.n4 16.8732
R55620 a_n1735_43236.n9 a_n1735_43236.n8 9.3005
R55621 a_3222_30651.n19 a_3222_30651.t16 1421.83
R55622 a_3222_30651.n9 a_3222_30651.t11 1421.83
R55623 a_3222_30651.n12 a_3222_30651.t6 1327.11
R55624 a_3222_30651.n16 a_3222_30651.t9 1327.11
R55625 a_3222_30651.n18 a_3222_30651.t17 1327.11
R55626 a_3222_30651.n8 a_3222_30651.t19 1327.11
R55627 a_3222_30651.n6 a_3222_30651.t5 1327.11
R55628 a_3222_30651.n2 a_3222_30651.t13 1327.11
R55629 a_3222_30651.n19 a_3222_30651.t20 1320.68
R55630 a_3222_30651.n17 a_3222_30651.t15 1320.68
R55631 a_3222_30651.n15 a_3222_30651.t10 1320.68
R55632 a_3222_30651.n13 a_3222_30651.t8 1320.68
R55633 a_3222_30651.n3 a_3222_30651.t12 1320.68
R55634 a_3222_30651.n5 a_3222_30651.t4 1320.68
R55635 a_3222_30651.n7 a_3222_30651.t21 1320.68
R55636 a_3222_30651.n9 a_3222_30651.t7 1320.68
R55637 a_3222_30651.n24 a_3222_30651.n0 380.32
R55638 a_3222_30651.n22 a_3222_30651.t14 260.322
R55639 a_3222_30651.n25 a_3222_30651.n24 185
R55640 a_3222_30651.n23 a_3222_30651.n22 178.451
R55641 a_3222_30651.n22 a_3222_30651.t18 175.169
R55642 a_3222_30651.n14 a_3222_30651.n13 161.701
R55643 a_3222_30651.n4 a_3222_30651.n3 161.701
R55644 a_3222_30651.n20 a_3222_30651.n19 161.3
R55645 a_3222_30651.n15 a_3222_30651.n14 161.3
R55646 a_3222_30651.n17 a_3222_30651.n11 161.3
R55647 a_3222_30651.n10 a_3222_30651.n9 161.3
R55648 a_3222_30651.n7 a_3222_30651.n1 161.3
R55649 a_3222_30651.n5 a_3222_30651.n4 161.3
R55650 a_3222_30651.n13 a_3222_30651.n12 94.7191
R55651 a_3222_30651.n15 a_3222_30651.n12 94.7191
R55652 a_3222_30651.n16 a_3222_30651.n15 94.7191
R55653 a_3222_30651.n17 a_3222_30651.n16 94.7191
R55654 a_3222_30651.n18 a_3222_30651.n17 94.7191
R55655 a_3222_30651.n19 a_3222_30651.n18 94.7191
R55656 a_3222_30651.n9 a_3222_30651.n8 94.7191
R55657 a_3222_30651.n8 a_3222_30651.n7 94.7191
R55658 a_3222_30651.n7 a_3222_30651.n6 94.7191
R55659 a_3222_30651.n6 a_3222_30651.n5 94.7191
R55660 a_3222_30651.n5 a_3222_30651.n2 94.7191
R55661 a_3222_30651.n3 a_3222_30651.n2 94.7191
R55662 a_3222_30651.n23 a_3222_30651.n21 91.881
R55663 a_3222_30651.n21 a_3222_30651.n20 43.5224
R55664 a_3222_30651.n21 a_3222_30651.n10 39.3015
R55665 a_3222_30651.n0 a_3222_30651.t3 26.5955
R55666 a_3222_30651.n0 a_3222_30651.t2 26.5955
R55667 a_3222_30651.n25 a_3222_30651.t0 24.9236
R55668 a_3222_30651.t1 a_3222_30651.n25 24.9236
R55669 a_3222_30651.n24 a_3222_30651.n23 17.7246
R55670 a_3222_30651.n14 a_3222_30651.n11 0.4005
R55671 a_3222_30651.n20 a_3222_30651.n11 0.4005
R55672 a_3222_30651.n10 a_3222_30651.n1 0.4005
R55673 a_3222_30651.n4 a_3222_30651.n1 0.4005
R55674 VCM.n60 VCM.n59 60.7943
R55675 VCM.n30 VCM.t23 47.8989
R55676 VCM.n1 VCM.t22 47.8989
R55677 VCM.n30 VCM.t45 47.4614
R55678 VCM.n31 VCM.t55 47.4614
R55679 VCM.n32 VCM.t21 47.4614
R55680 VCM.n33 VCM.t46 47.4614
R55681 VCM.n34 VCM.t26 47.4614
R55682 VCM.n37 VCM.t52 47.4614
R55683 VCM.n8 VCM.t50 47.4614
R55684 VCM.n5 VCM.t27 47.4614
R55685 VCM.n4 VCM.t47 47.4614
R55686 VCM.n3 VCM.t20 47.4614
R55687 VCM.n2 VCM.t54 47.4614
R55688 VCM.n1 VCM.t44 47.4614
R55689 VCM.n36 VCM.n35 37.5614
R55690 VCM.n7 VCM.n6 37.5614
R55691 VCM.n60 VCM.n29 35.4847
R55692 VCM.n59 VCM.t32 17.4125
R55693 VCM.n29 VCM.t37 17.4125
R55694 VCM.n40 VCM.n38 15.4323
R55695 VCM.n10 VCM.n0 15.4323
R55696 VCM.n58 VCM.n57 14.9375
R55697 VCM.n56 VCM.n55 14.9375
R55698 VCM.n54 VCM.n53 14.9375
R55699 VCM.n52 VCM.n51 14.9375
R55700 VCM.n50 VCM.n49 14.9375
R55701 VCM.n48 VCM.n47 14.9375
R55702 VCM.n46 VCM.n45 14.9375
R55703 VCM.n44 VCM.n43 14.9375
R55704 VCM.n42 VCM.n41 14.9375
R55705 VCM.n40 VCM.n39 14.9375
R55706 VCM.n28 VCM.n27 14.9375
R55707 VCM.n26 VCM.n25 14.9375
R55708 VCM.n24 VCM.n23 14.9375
R55709 VCM.n22 VCM.n21 14.9375
R55710 VCM.n20 VCM.n19 14.9375
R55711 VCM.n18 VCM.n17 14.9375
R55712 VCM.n16 VCM.n15 14.9375
R55713 VCM.n14 VCM.n13 14.9375
R55714 VCM.n12 VCM.n11 14.9375
R55715 VCM.n10 VCM.n9 14.9375
R55716 VCM.n35 VCM.t51 9.9005
R55717 VCM.n35 VCM.t24 9.9005
R55718 VCM.n6 VCM.t25 9.9005
R55719 VCM.n6 VCM.t53 9.9005
R55720 VCM.n40 VCM.n37 8.35002
R55721 VCM.n10 VCM.n8 8.35002
R55722 VCM VCM.n60 5.52202
R55723 VCM.n57 VCM.t35 2.4755
R55724 VCM.n57 VCM.t34 2.4755
R55725 VCM.n55 VCM.t33 2.4755
R55726 VCM.n55 VCM.t29 2.4755
R55727 VCM.n53 VCM.t31 2.4755
R55728 VCM.n53 VCM.t28 2.4755
R55729 VCM.n51 VCM.t30 2.4755
R55730 VCM.n51 VCM.t8 2.4755
R55731 VCM.n49 VCM.t6 2.4755
R55732 VCM.n49 VCM.t13 2.4755
R55733 VCM.n47 VCM.t15 2.4755
R55734 VCM.n47 VCM.t17 2.4755
R55735 VCM.n45 VCM.t11 2.4755
R55736 VCM.n45 VCM.t5 2.4755
R55737 VCM.n43 VCM.t4 2.4755
R55738 VCM.n43 VCM.t60 2.4755
R55739 VCM.n41 VCM.t59 2.4755
R55740 VCM.n41 VCM.t58 2.4755
R55741 VCM.n39 VCM.t61 2.4755
R55742 VCM.n39 VCM.t1 2.4755
R55743 VCM.n38 VCM.t3 2.4755
R55744 VCM.n38 VCM.t49 2.4755
R55745 VCM.n27 VCM.t36 2.4755
R55746 VCM.n27 VCM.t39 2.4755
R55747 VCM.n25 VCM.t40 2.4755
R55748 VCM.n25 VCM.t41 2.4755
R55749 VCM.n23 VCM.t38 2.4755
R55750 VCM.n23 VCM.t42 2.4755
R55751 VCM.n21 VCM.t18 2.4755
R55752 VCM.n21 VCM.t43 2.4755
R55753 VCM.n19 VCM.t14 2.4755
R55754 VCM.n19 VCM.t9 2.4755
R55755 VCM.n17 VCM.t10 2.4755
R55756 VCM.n17 VCM.t7 2.4755
R55757 VCM.n15 VCM.t12 2.4755
R55758 VCM.n15 VCM.t16 2.4755
R55759 VCM.n13 VCM.t62 2.4755
R55760 VCM.n13 VCM.t19 2.4755
R55761 VCM.n11 VCM.t56 2.4755
R55762 VCM.n11 VCM.t63 2.4755
R55763 VCM.n9 VCM.t0 2.4755
R55764 VCM.n9 VCM.t57 2.4755
R55765 VCM.n0 VCM.t48 2.4755
R55766 VCM.n0 VCM.t2 2.4755
R55767 VCM.n46 VCM.n44 0.53175
R55768 VCM.n54 VCM.n52 0.53175
R55769 VCM.n16 VCM.n14 0.53175
R55770 VCM.n24 VCM.n22 0.53175
R55771 VCM.n44 VCM.n42 0.5005
R55772 VCM.n48 VCM.n46 0.5005
R55773 VCM.n50 VCM.n48 0.5005
R55774 VCM.n52 VCM.n50 0.5005
R55775 VCM.n56 VCM.n54 0.5005
R55776 VCM.n58 VCM.n56 0.5005
R55777 VCM.n59 VCM.n58 0.5005
R55778 VCM.n14 VCM.n12 0.5005
R55779 VCM.n18 VCM.n16 0.5005
R55780 VCM.n20 VCM.n18 0.5005
R55781 VCM.n22 VCM.n20 0.5005
R55782 VCM.n26 VCM.n24 0.5005
R55783 VCM.n28 VCM.n26 0.5005
R55784 VCM.n29 VCM.n28 0.5005
R55785 VCM.n42 VCM.n40 0.495292
R55786 VCM.n12 VCM.n10 0.495292
R55787 VCM.n36 VCM.n34 0.438
R55788 VCM.n34 VCM.n33 0.438
R55789 VCM.n33 VCM.n32 0.438
R55790 VCM.n32 VCM.n31 0.438
R55791 VCM.n31 VCM.n30 0.438
R55792 VCM.n2 VCM.n1 0.438
R55793 VCM.n3 VCM.n2 0.438
R55794 VCM.n4 VCM.n3 0.438
R55795 VCM.n5 VCM.n4 0.438
R55796 VCM.n7 VCM.n5 0.438
R55797 VCM.n37 VCM.n36 0.396333
R55798 VCM.n8 VCM.n7 0.396333
R55799 C2_N_btm.n1 C2_N_btm.t8 101.621
R55800 C2_N_btm.n2 C2_N_btm.t1 98.936
R55801 C2_N_btm.n0 C2_N_btm.t7 54.9311
R55802 C2_N_btm C2_N_btm.n2 52.2505
R55803 C2_N_btm.n0 C2_N_btm.t0 47.3635
R55804 C2_N_btm C2_N_btm.n6 8.11925
R55805 C2_N_btm.n1 C2_N_btm.n0 7.71404
R55806 C2_N_btm.n2 C2_N_btm.n1 7.20883
R55807 C2_N_btm.n3 C2_N_btm.t5 4.76819
R55808 C2_N_btm.n5 C2_N_btm.t3 4.03712
R55809 C2_N_btm.n6 C2_N_btm.t6 4.03712
R55810 C2_N_btm.n4 C2_N_btm.t2 3.98193
R55811 C2_N_btm.n3 C2_N_btm.t4 3.92851
R55812 C2_N_btm.n5 C2_N_btm.n4 1.05569
R55813 C2_N_btm.n6 C2_N_btm.n5 1.0005
R55814 C2_N_btm.n4 C2_N_btm.n3 0.786757
R55815 COMP_P.n9 COMP_P.n7 267.779
R55816 COMP_P.n8 COMP_P.t9 260.322
R55817 COMP_P.n2 COMP_P.n1 244.069
R55818 COMP_P.n5 COMP_P.n3 236.589
R55819 COMP_P.n7 COMP_P.t8 230.155
R55820 COMP_P.n2 COMP_P.n0 204.893
R55821 COMP_P.n5 COMP_P.n4 200.321
R55822 COMP_P.n9 COMP_P.n8 194.517
R55823 COMP_P.n8 COMP_P.t10 175.169
R55824 COMP_P.n7 COMP_P.t11 157.856
R55825 COMP_P COMP_P.n9 30.5786
R55826 COMP_P.n6 COMP_P.n2 30.0599
R55827 COMP_P.n6 COMP_P.n5 27.5565
R55828 COMP_P.n0 COMP_P.t4 26.5955
R55829 COMP_P.n0 COMP_P.t6 26.5955
R55830 COMP_P.n1 COMP_P.t5 26.5955
R55831 COMP_P.n1 COMP_P.t7 26.5955
R55832 COMP_P.n3 COMP_P.t2 24.9236
R55833 COMP_P.n3 COMP_P.t0 24.9236
R55834 COMP_P.n4 COMP_P.t1 24.9236
R55835 COMP_P.n4 COMP_P.t3 24.9236
R55836 COMP_P COMP_P.n6 14.6286
R55837 a_n2467_30659.n1 a_n2467_30659.t6 756.547
R55838 a_n2467_30659.n7 a_n2467_30659.t7 756.231
R55839 a_n2467_30659.n6 a_n2467_30659.t4 756.226
R55840 a_n2467_30659.n5 a_n2467_30659.t9 756.226
R55841 a_n2467_30659.n4 a_n2467_30659.t8 756.226
R55842 a_n2467_30659.n3 a_n2467_30659.t11 756.226
R55843 a_n2467_30659.n2 a_n2467_30659.t10 756.226
R55844 a_n2467_30659.n1 a_n2467_30659.t5 756.226
R55845 a_n2467_30659.n8 a_n2467_30659.n0 287.752
R55846 a_n2467_30659.n9 a_n2467_30659.n8 277.568
R55847 a_n2467_30659.n8 a_n2467_30659.n7 117.487
R55848 a_n2467_30659.n0 a_n2467_30659.t2 26.5955
R55849 a_n2467_30659.n0 a_n2467_30659.t3 26.5955
R55850 a_n2467_30659.t1 a_n2467_30659.n9 24.9236
R55851 a_n2467_30659.n9 a_n2467_30659.t0 24.9236
R55852 a_n2467_30659.n2 a_n2467_30659.n1 0.3205
R55853 a_n2467_30659.n3 a_n2467_30659.n2 0.3205
R55854 a_n2467_30659.n4 a_n2467_30659.n3 0.3205
R55855 a_n2467_30659.n5 a_n2467_30659.n4 0.3205
R55856 a_n2467_30659.n6 a_n2467_30659.n5 0.3205
R55857 a_n2467_30659.n7 a_n2467_30659.n6 0.298833
R55858 a_10227_47214.n2 a_10227_47214.n0 647.148
R55859 a_10227_47214.n18 a_10227_47214.t25 408.63
R55860 a_10227_47214.n14 a_10227_47214.t34 408.63
R55861 a_10227_47214.n10 a_10227_47214.t18 408.63
R55862 a_10227_47214.n3 a_10227_47214.t28 408.63
R55863 a_10227_47214.n7 a_10227_47214.t37 408.63
R55864 a_10227_47214.n35 a_10227_47214.t41 408.63
R55865 a_10227_47214.n31 a_10227_47214.t14 408.63
R55866 a_10227_47214.n27 a_10227_47214.t45 408.63
R55867 a_10227_47214.n22 a_10227_47214.t30 408.63
R55868 a_10227_47214.n19 a_10227_47214.t21 347.577
R55869 a_10227_47214.n15 a_10227_47214.t33 347.577
R55870 a_10227_47214.n11 a_10227_47214.t20 347.577
R55871 a_10227_47214.n4 a_10227_47214.t12 347.577
R55872 a_10227_47214.n6 a_10227_47214.t22 347.577
R55873 a_10227_47214.n36 a_10227_47214.t13 347.577
R55874 a_10227_47214.n32 a_10227_47214.t42 347.577
R55875 a_10227_47214.n28 a_10227_47214.t9 347.577
R55876 a_10227_47214.n23 a_10227_47214.t39 347.577
R55877 a_10227_47214.n25 a_10227_47214.t31 261.887
R55878 a_10227_47214.n41 a_10227_47214.n40 243.627
R55879 a_10227_47214.n42 a_10227_47214.n41 200.262
R55880 a_10227_47214.n2 a_10227_47214.n1 194.441
R55881 a_10227_47214.n19 a_10227_47214.t16 193.337
R55882 a_10227_47214.n15 a_10227_47214.t11 193.337
R55883 a_10227_47214.n11 a_10227_47214.t27 193.337
R55884 a_10227_47214.n4 a_10227_47214.t40 193.337
R55885 a_10227_47214.n6 a_10227_47214.t43 193.337
R55886 a_10227_47214.n36 a_10227_47214.t10 193.337
R55887 a_10227_47214.n32 a_10227_47214.t44 193.337
R55888 a_10227_47214.n28 a_10227_47214.t26 193.337
R55889 a_10227_47214.n23 a_10227_47214.t15 193.337
R55890 a_10227_47214.n26 a_10227_47214.n25 179.504
R55891 a_10227_47214.n24 a_10227_47214.n22 167.666
R55892 a_10227_47214.n16 a_10227_47214.n14 167.663
R55893 a_10227_47214.n29 a_10227_47214.n27 167.663
R55894 a_10227_47214.n37 a_10227_47214.n35 167.605
R55895 a_10227_47214.n5 a_10227_47214.n3 167.567
R55896 a_10227_47214.n33 a_10227_47214.n31 165.179
R55897 a_10227_47214.n20 a_10227_47214.n18 165.072
R55898 a_10227_47214.n12 a_10227_47214.n10 165.072
R55899 a_10227_47214.n8 a_10227_47214.n7 165.072
R55900 a_10227_47214.n8 a_10227_47214.n6 163.007
R55901 a_10227_47214.n20 a_10227_47214.n19 163.006
R55902 a_10227_47214.n12 a_10227_47214.n11 163.006
R55903 a_10227_47214.n33 a_10227_47214.n32 162.835
R55904 a_10227_47214.n5 a_10227_47214.n4 160.512
R55905 a_10227_47214.n37 a_10227_47214.n36 160.476
R55906 a_10227_47214.n24 a_10227_47214.n23 160.415
R55907 a_10227_47214.n16 a_10227_47214.n15 160.415
R55908 a_10227_47214.n29 a_10227_47214.n28 160.415
R55909 a_10227_47214.n25 a_10227_47214.t19 155.847
R55910 a_10227_47214.n18 a_10227_47214.t36 132.282
R55911 a_10227_47214.n14 a_10227_47214.t23 132.282
R55912 a_10227_47214.n10 a_10227_47214.t29 132.282
R55913 a_10227_47214.n3 a_10227_47214.t8 132.282
R55914 a_10227_47214.n7 a_10227_47214.t38 132.282
R55915 a_10227_47214.n35 a_10227_47214.t17 132.282
R55916 a_10227_47214.n31 a_10227_47214.t24 132.282
R55917 a_10227_47214.n27 a_10227_47214.t32 132.282
R55918 a_10227_47214.n22 a_10227_47214.t35 132.282
R55919 a_10227_47214.n40 a_10227_47214.t0 40.0005
R55920 a_10227_47214.n40 a_10227_47214.t2 40.0005
R55921 a_10227_47214.t3 a_10227_47214.n42 40.0005
R55922 a_10227_47214.n42 a_10227_47214.t1 40.0005
R55923 a_10227_47214.n39 a_10227_47214.n2 32.1002
R55924 a_10227_47214.n38 a_10227_47214.n34 29.5017
R55925 a_10227_47214.n1 a_10227_47214.t7 27.5805
R55926 a_10227_47214.n1 a_10227_47214.t4 27.5805
R55927 a_10227_47214.n0 a_10227_47214.t6 27.5805
R55928 a_10227_47214.n0 a_10227_47214.t5 27.5805
R55929 a_10227_47214.n41 a_10227_47214.n39 18.4708
R55930 a_10227_47214.n34 a_10227_47214.n30 14.1049
R55931 a_10227_47214.n30 a_10227_47214.n26 11.6197
R55932 a_10227_47214.n38 a_10227_47214.n37 11.5442
R55933 a_10227_47214.n17 a_10227_47214.n13 9.88649
R55934 a_10227_47214.n39 a_10227_47214.n38 9.3005
R55935 a_10227_47214.n13 a_10227_47214.n12 8.45044
R55936 a_10227_47214.n9 a_10227_47214.n8 7.23894
R55937 a_10227_47214.n38 a_10227_47214.n21 7.08841
R55938 a_10227_47214.n13 a_10227_47214.n9 7.0527
R55939 a_10227_47214.n21 a_10227_47214.n20 6.15515
R55940 a_10227_47214.n17 a_10227_47214.n16 4.95334
R55941 a_10227_47214.n30 a_10227_47214.n29 4.54976
R55942 a_10227_47214.n34 a_10227_47214.n33 4.5005
R55943 a_10227_47214.n21 a_10227_47214.n17 4.11863
R55944 a_10227_47214.n9 a_10227_47214.n5 0.209244
R55945 a_10227_47214.n26 a_10227_47214.n24 0.0492375
R55946 a_n2810_47070.n1 a_n2810_47070.t6 756.547
R55947 a_n2810_47070.n3 a_n2810_47070.t5 756.226
R55948 a_n2810_47070.n2 a_n2810_47070.t7 756.226
R55949 a_n2810_47070.n1 a_n2810_47070.t4 756.226
R55950 a_n2810_47070.n4 a_n2810_47070.n0 287.752
R55951 a_n2810_47070.n5 a_n2810_47070.n4 277.568
R55952 a_n2810_47070.n4 a_n2810_47070.n3 119.692
R55953 a_n2810_47070.n0 a_n2810_47070.t3 26.5955
R55954 a_n2810_47070.n0 a_n2810_47070.t2 26.5955
R55955 a_n2810_47070.t1 a_n2810_47070.n5 24.9236
R55956 a_n2810_47070.n5 a_n2810_47070.t0 24.9236
R55957 a_n2810_47070.n2 a_n2810_47070.n1 0.3205
R55958 a_n2810_47070.n3 a_n2810_47070.n2 0.304667
R55959 SMPL_ON_N.n7 SMPL_ON_N.t8 260.322
R55960 SMPL_ON_N.n5 SMPL_ON_N.n3 244.069
R55961 SMPL_ON_N.n2 SMPL_ON_N.n1 236.589
R55962 SMPL_ON_N.n5 SMPL_ON_N.n4 204.893
R55963 SMPL_ON_N.n2 SMPL_ON_N.n0 200.321
R55964 SMPL_ON_N SMPL_ON_N.n7 178.226
R55965 SMPL_ON_N.n7 SMPL_ON_N.t9 175.169
R55966 SMPL_ON_N SMPL_ON_N.n6 71.3118
R55967 SMPL_ON_N.n6 SMPL_ON_N.n5 27.3803
R55968 SMPL_ON_N.n4 SMPL_ON_N.t7 26.5955
R55969 SMPL_ON_N.n4 SMPL_ON_N.t4 26.5955
R55970 SMPL_ON_N.n3 SMPL_ON_N.t6 26.5955
R55971 SMPL_ON_N.n3 SMPL_ON_N.t5 26.5955
R55972 SMPL_ON_N.n0 SMPL_ON_N.t2 24.9236
R55973 SMPL_ON_N.n0 SMPL_ON_N.t1 24.9236
R55974 SMPL_ON_N.n1 SMPL_ON_N.t0 24.9236
R55975 SMPL_ON_N.n1 SMPL_ON_N.t3 24.9236
R55976 SMPL_ON_N.n6 SMPL_ON_N.n2 24.8776
R55977 a_1343_38525.t10 a_1343_38525.n4 542.547
R55978 a_1343_38525.n7 a_1343_38525.t10 542.081
R55979 a_1343_38525.n2 a_1343_38525.n0 344.094
R55980 a_1343_38525.n2 a_1343_38525.n1 313.916
R55981 a_1343_38525.n6 a_1343_38525.t8 270.545
R55982 a_1343_38525.n12 a_1343_38525.n11 230.554
R55983 a_1343_38525.n11 a_1343_38525.n10 200.375
R55984 a_1343_38525.n3 a_1343_38525.t9 199.597
R55985 a_1343_38525.n5 a_1343_38525.t12 199.572
R55986 a_1343_38525.n3 a_1343_38525.t11 197.951
R55987 a_1343_38525.n5 a_1343_38525.t13 197.947
R55988 a_1343_38525.n0 a_1343_38525.t4 26.5955
R55989 a_1343_38525.n0 a_1343_38525.t7 26.5955
R55990 a_1343_38525.n1 a_1343_38525.t6 26.5955
R55991 a_1343_38525.n1 a_1343_38525.t5 26.5955
R55992 a_1343_38525.n10 a_1343_38525.t0 24.9236
R55993 a_1343_38525.n10 a_1343_38525.t1 24.9236
R55994 a_1343_38525.n12 a_1343_38525.t2 24.9236
R55995 a_1343_38525.t3 a_1343_38525.n12 24.9236
R55996 a_1343_38525.n9 a_1343_38525.n8 20.9036
R55997 a_1343_38525.n9 a_1343_38525.n2 9.56818
R55998 a_1343_38525.n11 a_1343_38525.n9 8.79242
R55999 a_1343_38525.n7 a_1343_38525.n6 4.16605
R56000 a_1343_38525.n6 a_1343_38525.n5 2.52511
R56001 a_1343_38525.n8 a_1343_38525.n4 1.76521
R56002 a_1343_38525.n4 a_1343_38525.n3 1.27548
R56003 a_1343_38525.n8 a_1343_38525.n7 0.473054
R56004 a_8727_47222.n20 a_8727_47222.n0 589.152
R56005 a_8727_47222.n5 a_8727_47222.t15 408.63
R56006 a_8727_47222.n2 a_8727_47222.t6 408.63
R56007 a_8727_47222.n9 a_8727_47222.t19 408.63
R56008 a_8727_47222.n4 a_8727_47222.t11 347.577
R56009 a_8727_47222.n1 a_8727_47222.t10 347.577
R56010 a_8727_47222.n10 a_8727_47222.t12 347.577
R56011 a_8727_47222.n21 a_8727_47222.n20 289.462
R56012 a_8727_47222.n17 a_8727_47222.t13 238.59
R56013 a_8727_47222.n14 a_8727_47222.t7 238.59
R56014 a_8727_47222.n16 a_8727_47222.t16 224.984
R56015 a_8727_47222.n17 a_8727_47222.t18 203.244
R56016 a_8727_47222.n14 a_8727_47222.t14 203.244
R56017 a_8727_47222.n18 a_8727_47222.n16 199.341
R56018 a_8727_47222.n4 a_8727_47222.t21 193.337
R56019 a_8727_47222.n1 a_8727_47222.t4 193.337
R56020 a_8727_47222.n10 a_8727_47222.t9 193.337
R56021 a_8727_47222.n16 a_8727_47222.t8 187.714
R56022 a_8727_47222.n15 a_8727_47222.n14 177.137
R56023 a_8727_47222.n18 a_8727_47222.n17 172.637
R56024 a_8727_47222.n3 a_8727_47222.n2 165.077
R56025 a_8727_47222.n6 a_8727_47222.n5 165.072
R56026 a_8727_47222.n6 a_8727_47222.n4 163.007
R56027 a_8727_47222.n3 a_8727_47222.n1 163
R56028 a_8727_47222.n11 a_8727_47222.n10 162.957
R56029 a_8727_47222.n12 a_8727_47222.n9 158.144
R56030 a_8727_47222.n5 a_8727_47222.t5 132.282
R56031 a_8727_47222.n2 a_8727_47222.t20 132.282
R56032 a_8727_47222.n9 a_8727_47222.t17 132.282
R56033 a_8727_47222.t1 a_8727_47222.n21 38.5719
R56034 a_8727_47222.n21 a_8727_47222.t0 38.5719
R56035 a_8727_47222.n15 a_8727_47222.n13 29.6103
R56036 a_8727_47222.n13 a_8727_47222.n12 27.7325
R56037 a_8727_47222.n0 a_8727_47222.t2 26.5955
R56038 a_8727_47222.n0 a_8727_47222.t3 26.5955
R56039 a_8727_47222.n7 a_8727_47222.n3 21.0049
R56040 a_8727_47222.n19 a_8727_47222.n18 19.8116
R56041 a_8727_47222.n8 a_8727_47222.n7 11.5527
R56042 a_8727_47222.n19 a_8727_47222.n15 10.4842
R56043 a_8727_47222.n12 a_8727_47222.n11 9.3005
R56044 a_8727_47222.n20 a_8727_47222.n19 9.3005
R56045 a_8727_47222.n7 a_8727_47222.n6 0.488944
R56046 a_8727_47222.n11 a_8727_47222.n8 0.175249
R56047 a_8727_47222.n13 a_8727_47222.n8 0.0101154
R56048 a_n1741_47596.n5 a_n1741_47596.n0 594.054
R56049 a_n1741_47596.n3 a_n1741_47596.t5 276.464
R56050 a_n1741_47596.n6 a_n1741_47596.n5 258.8
R56051 a_n1741_47596.n1 a_n1741_47596.t6 212.081
R56052 a_n1741_47596.n2 a_n1741_47596.t9 212.081
R56053 a_n1741_47596.n4 a_n1741_47596.n2 211.435
R56054 a_n1741_47596.n3 a_n1741_47596.t7 196.131
R56055 a_n1741_47596.n4 a_n1741_47596.n3 192.407
R56056 a_n1741_47596.n1 a_n1741_47596.t8 139.78
R56057 a_n1741_47596.n2 a_n1741_47596.t4 139.78
R56058 a_n1741_47596.n2 a_n1741_47596.n1 61.346
R56059 a_n1741_47596.n0 a_n1741_47596.t2 26.5955
R56060 a_n1741_47596.n0 a_n1741_47596.t3 26.5955
R56061 a_n1741_47596.n6 a_n1741_47596.t0 24.9236
R56062 a_n1741_47596.t1 a_n1741_47596.n6 24.9236
R56063 a_n1741_47596.n5 a_n1741_47596.n4 18.4905
R56064 a_n1827_44868.n8 a_n1827_44868.n7 300.118
R56065 a_n1827_44868.n5 a_n1827_44868.n4 299.834
R56066 a_n1827_44868.n10 a_n1827_44868.n9 299.834
R56067 a_n1827_44868.n8 a_n1827_44868.n6 291.81
R56068 a_n1827_44868.n0 a_n1827_44868.t9 276.464
R56069 a_n1827_44868.n3 a_n1827_44868.n2 254.654
R56070 a_n1827_44868.n2 a_n1827_44868.t10 212.081
R56071 a_n1827_44868.n1 a_n1827_44868.t11 212.081
R56072 a_n1827_44868.n3 a_n1827_44868.n0 204.424
R56073 a_n1827_44868.n0 a_n1827_44868.t8 196.131
R56074 a_n1827_44868.n2 a_n1827_44868.t13 139.78
R56075 a_n1827_44868.n1 a_n1827_44868.t12 139.78
R56076 a_n1827_44868.n9 a_n1827_44868.n8 79.8031
R56077 a_n1827_44868.n2 a_n1827_44868.n1 61.346
R56078 a_n1827_44868.n9 a_n1827_44868.n5 29.6732
R56079 a_n1827_44868.n7 a_n1827_44868.t5 26.5955
R56080 a_n1827_44868.n7 a_n1827_44868.t4 26.5955
R56081 a_n1827_44868.n4 a_n1827_44868.t6 26.5955
R56082 a_n1827_44868.n4 a_n1827_44868.t7 26.5955
R56083 a_n1827_44868.n10 a_n1827_44868.t1 26.5955
R56084 a_n1827_44868.t0 a_n1827_44868.n10 26.5955
R56085 a_n1827_44868.n6 a_n1827_44868.t2 24.9236
R56086 a_n1827_44868.n6 a_n1827_44868.t3 24.9236
R56087 a_n1827_44868.n5 a_n1827_44868.n3 10.4582
R56088 a_5142_30651.n2 a_5142_30651.t4 1421.83
R56089 a_5142_30651.n1 a_5142_30651.t5 1421.83
R56090 a_5142_30651.n2 a_5142_30651.t6 1320.68
R56091 a_5142_30651.n1 a_5142_30651.t9 1320.68
R56092 a_5142_30651.n6 a_5142_30651.n0 380.32
R56093 a_5142_30651.n4 a_5142_30651.t8 260.322
R56094 a_5142_30651.n3 a_5142_30651.n2 194.853
R56095 a_5142_30651.n3 a_5142_30651.n1 192.882
R56096 a_5142_30651.n7 a_5142_30651.n6 185
R56097 a_5142_30651.n4 a_5142_30651.t7 175.169
R56098 a_5142_30651.n5 a_5142_30651.n4 173.925
R56099 a_5142_30651.n5 a_5142_30651.n3 73.4209
R56100 a_5142_30651.n0 a_5142_30651.t2 26.5955
R56101 a_5142_30651.n0 a_5142_30651.t3 26.5955
R56102 a_5142_30651.n7 a_5142_30651.t0 24.9236
R56103 a_5142_30651.t1 a_5142_30651.n7 24.9236
R56104 a_5142_30651.n6 a_5142_30651.n5 16.8317
R56105 a_13144_47452.t4 a_13144_47452.t2 392.027
R56106 a_13144_47452.n1 a_13144_47452.t4 382.327
R56107 a_13144_47452.n2 a_13144_47452.t1 366.548
R56108 a_13144_47452.n0 a_13144_47452.t3 329.007
R56109 a_13144_47452.t0 a_13144_47452.n2 310.909
R56110 a_13144_47452.n0 a_13144_47452.t5 200.475
R56111 a_13144_47452.n1 a_13144_47452.n0 167.381
R56112 a_13144_47452.n2 a_13144_47452.n1 45.5515
R56113 a_12769_44594.n2 a_12769_44594.t7 722.096
R56114 a_12769_44594.n3 a_12769_44594.t5 722.096
R56115 a_12769_44594.n7 a_12769_44594.t1 364.055
R56116 a_12769_44594.t0 a_12769_44594.n7 292.207
R56117 a_12769_44594.n0 a_12769_44594.t9 238.59
R56118 a_12769_44594.n1 a_12769_44594.t6 230.793
R56119 a_12769_44594.n0 a_12769_44594.t3 203.244
R56120 a_12769_44594.n4 a_12769_44594.n3 181.345
R56121 a_12769_44594.n6 a_12769_44594.n0 174.696
R56122 a_12769_44594.n4 a_12769_44594.n2 168.016
R56123 a_12769_44594.n5 a_12769_44594.n1 164.367
R56124 a_12769_44594.n2 a_12769_44594.t2 162.963
R56125 a_12769_44594.n3 a_12769_44594.t4 162.963
R56126 a_12769_44594.n1 a_12769_44594.t8 158.494
R56127 a_12769_44594.n7 a_12769_44594.n6 23.4881
R56128 a_12769_44594.n5 a_12769_44594.n4 18.4277
R56129 a_12769_44594.n6 a_12769_44594.n5 4.04171
R56130 a_n237_45454.n20 a_n237_45454.n0 633.351
R56131 a_n237_45454.n9 a_n237_45454.t23 327.057
R56132 a_n237_45454.n18 a_n237_45454.t20 261.887
R56133 a_n237_45454.n16 a_n237_45454.t15 261.887
R56134 a_n237_45454.n1 a_n237_45454.t9 261.887
R56135 a_n237_45454.n13 a_n237_45454.t17 261.887
R56136 a_n237_45454.n3 a_n237_45454.t5 261.887
R56137 a_n237_45454.n5 a_n237_45454.t10 261.887
R56138 a_n237_45454.n4 a_n237_45454.t13 261.887
R56139 a_n237_45454.n2 a_n237_45454.t22 261.887
R56140 a_n237_45454.n21 a_n237_45454.n20 245.263
R56141 a_n237_45454.n9 a_n237_45454.t16 239.768
R56142 a_n237_45454.n11 a_n237_45454.t19 238.155
R56143 a_n237_45454.n17 a_n237_45454.n16 186.877
R56144 a_n237_45454.n10 a_n237_45454.n9 186.042
R56145 a_n237_45454.n7 a_n237_45454.n3 179.673
R56146 a_n237_45454.n14 a_n237_45454.n13 179.181
R56147 a_n237_45454.n8 a_n237_45454.n2 177.716
R56148 a_n237_45454.n19 a_n237_45454.n18 176.554
R56149 a_n237_45454.n12 a_n237_45454.n11 174.821
R56150 a_n237_45454.n11 a_n237_45454.t11 165.856
R56151 a_n237_45454.n6 a_n237_45454.n4 164.382
R56152 a_n237_45454.n15 a_n237_45454.n1 162.969
R56153 a_n237_45454.n6 a_n237_45454.n5 162.429
R56154 a_n237_45454.n18 a_n237_45454.t8 155.847
R56155 a_n237_45454.n16 a_n237_45454.t7 155.847
R56156 a_n237_45454.n1 a_n237_45454.t14 155.847
R56157 a_n237_45454.n13 a_n237_45454.t12 155.847
R56158 a_n237_45454.n3 a_n237_45454.t21 155.847
R56159 a_n237_45454.n5 a_n237_45454.t6 155.847
R56160 a_n237_45454.n4 a_n237_45454.t18 155.847
R56161 a_n237_45454.n2 a_n237_45454.t4 155.847
R56162 a_n237_45454.t1 a_n237_45454.n21 38.5719
R56163 a_n237_45454.n21 a_n237_45454.t0 38.5719
R56164 a_n237_45454.n20 a_n237_45454.n19 29.2773
R56165 a_n237_45454.n0 a_n237_45454.t2 26.5955
R56166 a_n237_45454.n0 a_n237_45454.t3 26.5955
R56167 a_n237_45454.n7 a_n237_45454.n6 23.4169
R56168 a_n237_45454.n14 a_n237_45454.n12 10.5403
R56169 a_n237_45454.n8 a_n237_45454.n7 10.5115
R56170 a_n237_45454.n17 a_n237_45454.n15 8.09528
R56171 a_n237_45454.n12 a_n237_45454.n10 6.44032
R56172 a_n237_45454.n15 a_n237_45454.n14 5.86314
R56173 a_n237_45454.n10 a_n237_45454.n8 4.85096
R56174 a_n237_45454.n19 a_n237_45454.n17 0.69006
R56175 a_927_42692.n3 a_927_42692.t19 334.723
R56176 a_927_42692.n7 a_927_42692.t13 267.065
R56177 a_927_42692.n4 a_927_42692.t16 256.716
R56178 a_927_42692.n2 a_927_42692.n0 248.088
R56179 a_927_42692.n16 a_927_42692.t11 241.536
R56180 a_927_42692.n14 a_927_42692.t8 238.397
R56181 a_927_42692.n13 a_927_42692.t14 231.835
R56182 a_927_42692.n8 a_927_42692.t9 221.72
R56183 a_927_42692.n9 a_927_42692.t21 221.72
R56184 a_927_42692.n2 a_927_42692.n1 208.508
R56185 a_927_42692.n3 a_927_42692.t22 206.19
R56186 a_927_42692.n14 a_927_42692.t12 195.017
R56187 a_927_42692.n19 a_927_42692.n3 187.038
R56188 a_927_42692.n11 a_927_42692.n7 185.536
R56189 a_927_42692.n17 a_927_42692.n16 178.263
R56190 a_927_42692.n16 a_927_42692.t18 169.237
R56191 a_927_42692.n11 a_927_42692.n10 168.752
R56192 a_927_42692.n6 a_927_42692.n4 164.01
R56193 a_927_42692.n6 a_927_42692.n5 163.944
R56194 a_927_42692.n15 a_927_42692.n13 163.349
R56195 a_927_42692.n15 a_927_42692.n14 162.29
R56196 a_927_42692.n4 a_927_42692.t23 161.275
R56197 a_927_42692.n13 a_927_42692.t25 157.07
R56198 a_927_42692.n8 a_927_42692.t17 149.421
R56199 a_927_42692.n9 a_927_42692.t20 149.421
R56200 a_927_42692.n7 a_927_42692.t15 148.35
R56201 a_927_42692.n23 a_927_42692.n22 137.575
R56202 a_927_42692.n5 a_927_42692.t24 137.177
R56203 a_927_42692.n5 a_927_42692.t10 121.109
R56204 a_927_42692.n22 a_927_42692.n21 99.1749
R56205 a_927_42692.n10 a_927_42692.n8 37.4894
R56206 a_927_42692.n10 a_927_42692.n9 37.4894
R56207 a_927_42692.n22 a_927_42692.n20 36.0958
R56208 a_927_42692.n0 a_927_42692.t5 26.5955
R56209 a_927_42692.n0 a_927_42692.t7 26.5955
R56210 a_927_42692.n1 a_927_42692.t6 26.5955
R56211 a_927_42692.n1 a_927_42692.t4 26.5955
R56212 a_927_42692.n21 a_927_42692.t2 24.9236
R56213 a_927_42692.n21 a_927_42692.t1 24.9236
R56214 a_927_42692.t3 a_927_42692.n23 24.9236
R56215 a_927_42692.n23 a_927_42692.t0 24.9236
R56216 a_927_42692.n20 a_927_42692.n2 17.2539
R56217 a_927_42692.n20 a_927_42692.n19 14.7145
R56218 a_927_42692.n17 a_927_42692.n15 12.6018
R56219 a_927_42692.n19 a_927_42692.n18 9.04987
R56220 a_927_42692.n12 a_927_42692.n11 8.30957
R56221 a_927_42692.n12 a_927_42692.n6 5.88649
R56222 a_927_42692.n18 a_927_42692.n12 4.55733
R56223 a_927_42692.n18 a_927_42692.n17 0.914477
R56224 a_17930_32299.n3 a_17930_32299.t4 1415.15
R56225 a_17930_32299.n2 a_17930_32299.t5 1330.32
R56226 a_17930_32299.n1 a_17930_32299.t6 1320.68
R56227 a_17930_32299.n3 a_17930_32299.t7 1320.68
R56228 a_17930_32299.n5 a_17930_32299.n0 380.32
R56229 a_17930_32299.n6 a_17930_32299.n5 185
R56230 a_17930_32299.n4 a_17930_32299.n1 161.764
R56231 a_17930_32299.n4 a_17930_32299.n3 161.3
R56232 a_17930_32299.n5 a_17930_32299.n4 119.462
R56233 a_17930_32299.n3 a_17930_32299.n2 84.8325
R56234 a_17930_32299.n2 a_17930_32299.n1 84.8325
R56235 a_17930_32299.n0 a_17930_32299.t3 26.5955
R56236 a_17930_32299.n0 a_17930_32299.t2 26.5955
R56237 a_17930_32299.n6 a_17930_32299.t0 24.9236
R56238 a_17930_32299.t1 a_17930_32299.n6 24.9236
R56239 a_20163_31459.n1 a_20163_31459.t4 604.578
R56240 a_20163_31459.n1 a_20163_31459.n0 287.752
R56241 a_20163_31459.n2 a_20163_31459.n1 277.568
R56242 a_20163_31459.n0 a_20163_31459.t2 26.5955
R56243 a_20163_31459.n0 a_20163_31459.t3 26.5955
R56244 a_20163_31459.t1 a_20163_31459.n2 24.9236
R56245 a_20163_31459.n2 a_20163_31459.t0 24.9236
R56246 C3_N_btm.n1 C3_N_btm.t1 101.516
R56247 C3_N_btm.n2 C3_N_btm.t0 100.142
R56248 C3_N_btm.n0 C3_N_btm.t12 54.9311
R56249 C3_N_btm C3_N_btm.n2 47.7713
R56250 C3_N_btm.n0 C3_N_btm.t11 47.3635
R56251 C3_N_btm.n2 C3_N_btm.n1 9.7505
R56252 C3_N_btm C3_N_btm.n10 9.213
R56253 C3_N_btm.n1 C3_N_btm.n0 7.43279
R56254 C3_N_btm.n3 C3_N_btm.t5 4.76719
R56255 C3_N_btm.n8 C3_N_btm.t4 4.03712
R56256 C3_N_btm.n9 C3_N_btm.t2 4.03712
R56257 C3_N_btm.n10 C3_N_btm.t10 4.03712
R56258 C3_N_btm.n7 C3_N_btm.t3 3.98193
R56259 C3_N_btm.n6 C3_N_btm.t6 3.92851
R56260 C3_N_btm.n5 C3_N_btm.t9 3.92851
R56261 C3_N_btm.n4 C3_N_btm.t7 3.92851
R56262 C3_N_btm.n3 C3_N_btm.t8 3.92851
R56263 C3_N_btm.n8 C3_N_btm.n7 1.05569
R56264 C3_N_btm.n9 C3_N_btm.n8 1.0005
R56265 C3_N_btm.n10 C3_N_btm.n9 1.0005
R56266 C3_N_btm.n4 C3_N_btm.n3 0.840176
R56267 C3_N_btm.n5 C3_N_btm.n4 0.840176
R56268 C3_N_btm.n6 C3_N_btm.n5 0.840176
R56269 C3_N_btm.n7 C3_N_btm.n6 0.786757
R56270 a_n2109_47596.n5 a_n2109_47596.n0 664.928
R56271 a_n2109_47596.n4 a_n2109_47596.n3 284.575
R56272 a_n2109_47596.n3 a_n2109_47596.t5 276.464
R56273 a_n2109_47596.n4 a_n2109_47596.n2 223.156
R56274 a_n2109_47596.n1 a_n2109_47596.t9 212.081
R56275 a_n2109_47596.n2 a_n2109_47596.t8 212.081
R56276 a_n2109_47596.n3 a_n2109_47596.t4 196.131
R56277 a_n2109_47596.n6 a_n2109_47596.n5 187.927
R56278 a_n2109_47596.n1 a_n2109_47596.t6 139.78
R56279 a_n2109_47596.n2 a_n2109_47596.t7 139.78
R56280 a_n2109_47596.n2 a_n2109_47596.n1 61.346
R56281 a_n2109_47596.n0 a_n2109_47596.t3 26.5955
R56282 a_n2109_47596.n0 a_n2109_47596.t2 26.5955
R56283 a_n2109_47596.n6 a_n2109_47596.t0 24.9236
R56284 a_n2109_47596.t1 a_n2109_47596.n6 24.9236
R56285 a_n2109_47596.n5 a_n2109_47596.n4 9.3005
R56286 a_13248_45956.n21 a_13248_45956.n0 589.152
R56287 a_13248_45956.t14 a_13248_45956.t7 547.874
R56288 a_13248_45956.t12 a_13248_45956.t27 395.01
R56289 a_13248_45956.n2 a_13248_45956.t8 377.241
R56290 a_13248_45956.n11 a_13248_45956.t12 333.245
R56291 a_13248_45956.n17 a_13248_45956.t13 329.902
R56292 a_13248_45956.n7 a_13248_45956.t16 322.216
R56293 a_13248_45956.n6 a_13248_45956.t22 305.267
R56294 a_13248_45956.n22 a_13248_45956.n21 289.462
R56295 a_13248_45956.n12 a_13248_45956.t6 241.536
R56296 a_13248_45956.n18 a_13248_45956.t9 230.155
R56297 a_13248_45956.n3 a_13248_45956.t20 223.327
R56298 a_13248_45956.n14 a_13248_45956.t15 212.081
R56299 a_13248_45956.n13 a_13248_45956.t19 212.081
R56300 a_13248_45956.n15 a_13248_45956.n14 200.048
R56301 a_13248_45956.n1 a_13248_45956.t10 196.549
R56302 a_13248_45956.n8 a_13248_45956.t18 194.213
R56303 a_13248_45956.n9 a_13248_45956.n5 186.18
R56304 a_13248_45956.n9 a_13248_45956.n8 182.131
R56305 a_13248_45956.n6 a_13248_45956.t26 179.823
R56306 a_13248_45956.n10 a_13248_45956.n1 177.911
R56307 a_13248_45956.n2 a_13248_45956.t5 173.996
R56308 a_13248_45956.n15 a_13248_45956.n12 170.375
R56309 a_13248_45956.n12 a_13248_45956.t4 169.237
R56310 a_13248_45956.n19 a_13248_45956.n17 165.312
R56311 a_13248_45956.n19 a_13248_45956.n18 163.605
R56312 a_13248_45956.n18 a_13248_45956.t23 157.856
R56313 a_13248_45956.n1 a_13248_45956.t21 148.35
R56314 a_13248_45956.n14 a_13248_45956.t25 139.78
R56315 a_13248_45956.n13 a_13248_45956.t17 139.78
R56316 a_13248_45956.n17 a_13248_45956.t11 132.282
R56317 a_13248_45956.n5 a_13248_45956.t24 130.27
R56318 a_13248_45956.n7 a_13248_45956.n6 126.803
R56319 a_13248_45956.n4 a_13248_45956.t14 123.43
R56320 a_13248_45956.n14 a_13248_45956.n13 61.346
R56321 a_13248_45956.n4 a_13248_45956.n3 41.3757
R56322 a_13248_45956.n22 a_13248_45956.t0 38.5719
R56323 a_13248_45956.t1 a_13248_45956.n22 38.5719
R56324 a_13248_45956.n21 a_13248_45956.n20 32.501
R56325 a_13248_45956.n0 a_13248_45956.t3 26.5955
R56326 a_13248_45956.n0 a_13248_45956.t2 26.5955
R56327 a_13248_45956.n5 a_13248_45956.n4 24.7519
R56328 a_13248_45956.n20 a_13248_45956.n19 12.1366
R56329 a_13248_45956.n16 a_13248_45956.n11 8.49363
R56330 a_13248_45956.n16 a_13248_45956.n15 7.40435
R56331 a_13248_45956.n11 a_13248_45956.n10 4.5005
R56332 a_13248_45956.n20 a_13248_45956.n16 3.56506
R56333 a_13248_45956.n10 a_13248_45956.n9 3.20792
R56334 a_13248_45956.n3 a_13248_45956.n2 1.78419
R56335 a_13248_45956.n8 a_13248_45956.n7 0.53017
R56336 a_n1067_42718.n2 a_n1067_42718.t4 471.289
R56337 a_n1067_42718.n5 a_n1067_42718.t1 366.548
R56338 a_n1067_42718.t0 a_n1067_42718.n5 307.562
R56339 a_n1067_42718.n0 a_n1067_42718.t3 256.07
R56340 a_n1067_42718.n1 a_n1067_42718.t2 239.505
R56341 a_n1067_42718.n3 a_n1067_42718.n1 200.108
R56342 a_n1067_42718.n4 a_n1067_42718.n0 196.395
R56343 a_n1067_42718.n1 a_n1067_42718.t6 167.204
R56344 a_n1067_42718.n3 a_n1067_42718.n2 162.514
R56345 a_n1067_42718.n0 a_n1067_42718.t7 150.03
R56346 a_n1067_42718.n2 a_n1067_42718.t5 148.35
R56347 a_n1067_42718.n5 a_n1067_42718.n4 24.9173
R56348 a_n1067_42718.n4 a_n1067_42718.n3 23.4989
R56349 a_n1890_42718.n1 a_n1890_42718.t4 682.793
R56350 a_n1890_42718.n1 a_n1890_42718.n0 296.139
R56351 a_n1890_42718.n2 a_n1890_42718.n1 269.182
R56352 a_n1890_42718.n0 a_n1890_42718.t3 26.5955
R56353 a_n1890_42718.n0 a_n1890_42718.t2 26.5955
R56354 a_n1890_42718.t1 a_n1890_42718.n2 24.9236
R56355 a_n1890_42718.n2 a_n1890_42718.t0 24.9236
R56356 a_1334_43494.n4 a_1334_43494.t13 334.723
R56357 a_1334_43494.n3 a_1334_43494.t8 330.12
R56358 a_1334_43494.n13 a_1334_43494.t19 267.065
R56359 a_1334_43494.n16 a_1334_43494.t18 256.728
R56360 a_1334_43494.n2 a_1334_43494.n0 248.087
R56361 a_1334_43494.n19 a_1334_43494.t14 241.536
R56362 a_1334_43494.n6 a_1334_43494.t24 238.397
R56363 a_1334_43494.n7 a_1334_43494.t25 231.835
R56364 a_1334_43494.n9 a_1334_43494.t16 221.72
R56365 a_1334_43494.n10 a_1334_43494.t11 221.72
R56366 a_1334_43494.n5 a_1334_43494.n4 211.958
R56367 a_1334_43494.n14 a_1334_43494.n13 210.103
R56368 a_1334_43494.n2 a_1334_43494.n1 208.507
R56369 a_1334_43494.n4 a_1334_43494.t21 206.19
R56370 a_1334_43494.n3 a_1334_43494.t9 201.587
R56371 a_1334_43494.n6 a_1334_43494.t26 195.017
R56372 a_1334_43494.n8 a_1334_43494.n6 189.375
R56373 a_1334_43494.n20 a_1334_43494.n19 186.225
R56374 a_1334_43494.n19 a_1334_43494.t17 169.237
R56375 a_1334_43494.n5 a_1334_43494.n3 168.578
R56376 a_1334_43494.n17 a_1334_43494.n16 168.351
R56377 a_1334_43494.n15 a_1334_43494.n11 166.288
R56378 a_1334_43494.n8 a_1334_43494.n7 163.349
R56379 a_1334_43494.n14 a_1334_43494.n12 163.024
R56380 a_1334_43494.n16 a_1334_43494.t10 161.275
R56381 a_1334_43494.n7 a_1334_43494.t23 157.07
R56382 a_1334_43494.n9 a_1334_43494.t12 149.421
R56383 a_1334_43494.n10 a_1334_43494.t22 149.421
R56384 a_1334_43494.n13 a_1334_43494.t15 148.35
R56385 a_1334_43494.n25 a_1334_43494.n24 137.576
R56386 a_1334_43494.n12 a_1334_43494.t20 137.177
R56387 a_1334_43494.n12 a_1334_43494.t27 121.109
R56388 a_1334_43494.n24 a_1334_43494.n23 99.1759
R56389 a_1334_43494.n22 a_1334_43494.n2 38.4831
R56390 a_1334_43494.n11 a_1334_43494.n9 37.4894
R56391 a_1334_43494.n11 a_1334_43494.n10 37.4894
R56392 a_1334_43494.n0 a_1334_43494.t4 26.5955
R56393 a_1334_43494.n0 a_1334_43494.t5 26.5955
R56394 a_1334_43494.n1 a_1334_43494.t6 26.5955
R56395 a_1334_43494.n1 a_1334_43494.t7 26.5955
R56396 a_1334_43494.n23 a_1334_43494.t0 24.9236
R56397 a_1334_43494.n23 a_1334_43494.t1 24.9236
R56398 a_1334_43494.n25 a_1334_43494.t2 24.9236
R56399 a_1334_43494.t3 a_1334_43494.n25 24.9236
R56400 a_1334_43494.n21 a_1334_43494.n5 18.8206
R56401 a_1334_43494.n24 a_1334_43494.n22 14.8665
R56402 a_1334_43494.n18 a_1334_43494.n8 13.013
R56403 a_1334_43494.n22 a_1334_43494.n21 9.48846
R56404 a_1334_43494.n17 a_1334_43494.n15 8.57056
R56405 a_1334_43494.n21 a_1334_43494.n20 6.09528
R56406 a_1334_43494.n18 a_1334_43494.n17 4.5005
R56407 a_1334_43494.n15 a_1334_43494.n14 3.28621
R56408 a_1334_43494.n20 a_1334_43494.n18 0.69006
R56409 a_5734_30651.n2 a_5734_30651.t5 646.679
R56410 a_5734_30651.n2 a_5734_30651.t6 642.65
R56411 a_5734_30651.n4 a_5734_30651.n0 380.32
R56412 a_5734_30651.n1 a_5734_30651.t4 260.322
R56413 a_5734_30651.n5 a_5734_30651.n4 185
R56414 a_5734_30651.n3 a_5734_30651.n1 176.254
R56415 a_5734_30651.n1 a_5734_30651.t7 175.169
R56416 a_5734_30651.n3 a_5734_30651.n2 133.279
R56417 a_5734_30651.n0 a_5734_30651.t3 26.5955
R56418 a_5734_30651.n0 a_5734_30651.t2 26.5955
R56419 a_5734_30651.n5 a_5734_30651.t0 24.9236
R56420 a_5734_30651.t1 a_5734_30651.n5 24.9236
R56421 a_5734_30651.n4 a_5734_30651.n3 21.2067
R56422 a_n690_43494.n20 a_n690_43494.n0 688.152
R56423 a_n690_43494.n17 a_n690_43494.t7 294.557
R56424 a_n690_43494.n2 a_n690_43494.t18 294.557
R56425 a_n690_43494.n12 a_n690_43494.t15 294.557
R56426 a_n690_43494.n11 a_n690_43494.t13 294.557
R56427 a_n690_43494.n8 a_n690_43494.t4 294.557
R56428 a_n690_43494.n9 a_n690_43494.t9 294.557
R56429 a_n690_43494.n6 a_n690_43494.t10 294.557
R56430 a_n690_43494.n4 a_n690_43494.t12 294.557
R56431 a_n690_43494.n3 a_n690_43494.t20 294.557
R56432 a_n690_43494.n1 a_n690_43494.t14 294.557
R56433 a_n690_43494.n17 a_n690_43494.t8 211.01
R56434 a_n690_43494.n2 a_n690_43494.t11 211.01
R56435 a_n690_43494.n12 a_n690_43494.t21 211.01
R56436 a_n690_43494.n11 a_n690_43494.t19 211.01
R56437 a_n690_43494.n8 a_n690_43494.t16 211.01
R56438 a_n690_43494.n9 a_n690_43494.t22 211.01
R56439 a_n690_43494.n6 a_n690_43494.t6 211.01
R56440 a_n690_43494.n4 a_n690_43494.t5 211.01
R56441 a_n690_43494.n3 a_n690_43494.t23 211.01
R56442 a_n690_43494.n1 a_n690_43494.t17 211.01
R56443 a_n690_43494.n21 a_n690_43494.n20 190.62
R56444 a_n690_43494.n5 a_n690_43494.n3 186.94
R56445 a_n690_43494.n10 a_n690_43494.n8 179.332
R56446 a_n690_43494.n13 a_n690_43494.n11 177.274
R56447 a_n690_43494.n16 a_n690_43494.n2 175.269
R56448 a_n690_43494.n18 a_n690_43494.n17 175.213
R56449 a_n690_43494.n19 a_n690_43494.n1 174.95
R56450 a_n690_43494.n13 a_n690_43494.n12 174.832
R56451 a_n690_43494.n7 a_n690_43494.n6 174.832
R56452 a_n690_43494.n5 a_n690_43494.n4 174.832
R56453 a_n690_43494.n10 a_n690_43494.n9 171.477
R56454 a_n690_43494.n21 a_n690_43494.t0 38.5719
R56455 a_n690_43494.t1 a_n690_43494.n21 38.5719
R56456 a_n690_43494.n0 a_n690_43494.t2 26.5955
R56457 a_n690_43494.n0 a_n690_43494.t3 26.5955
R56458 a_n690_43494.n19 a_n690_43494.n18 24.1297
R56459 a_n690_43494.n16 a_n690_43494.n15 15.0582
R56460 a_n690_43494.n15 a_n690_43494.n14 13.4758
R56461 a_n690_43494.n20 a_n690_43494.n19 9.3005
R56462 a_n690_43494.n14 a_n690_43494.n10 9.06305
R56463 a_n690_43494.n7 a_n690_43494.n5 8.09819
R56464 a_n690_43494.n14 a_n690_43494.n13 6.04682
R56465 a_n690_43494.n15 a_n690_43494.n7 3.16962
R56466 a_n690_43494.n18 a_n690_43494.n16 1.9222
R56467 a_17738_32299.n1 a_17738_32299.t5 1415.15
R56468 a_17738_32299.n1 a_17738_32299.t4 1320.68
R56469 a_17738_32299.n2 a_17738_32299.n0 296.139
R56470 a_17738_32299.n2 a_17738_32299.n1 282.541
R56471 a_17738_32299.n3 a_17738_32299.n2 269.182
R56472 a_17738_32299.n0 a_17738_32299.t2 26.5955
R56473 a_17738_32299.n0 a_17738_32299.t3 26.5955
R56474 a_17738_32299.t1 a_17738_32299.n3 24.9236
R56475 a_17738_32299.n3 a_17738_32299.t0 24.9236
R56476 a_6974_31099.n1 a_6974_31099.t5 570.641
R56477 a_6974_31099.n1 a_6974_31099.t4 568.112
R56478 a_6974_31099.n2 a_6974_31099.n0 380.32
R56479 a_6974_31099.n2 a_6974_31099.n1 200.976
R56480 a_6974_31099.n3 a_6974_31099.n2 185
R56481 a_6974_31099.n0 a_6974_31099.t2 26.5955
R56482 a_6974_31099.n0 a_6974_31099.t3 26.5955
R56483 a_6974_31099.t1 a_6974_31099.n3 24.9236
R56484 a_6974_31099.n3 a_6974_31099.t0 24.9236
R56485 a_n2661_45420.n5 a_n2661_45420.n0 664.928
R56486 a_n2661_45420.n4 a_n2661_45420.n3 321.416
R56487 a_n2661_45420.n1 a_n2661_45420.t5 276.464
R56488 a_n2661_45420.n2 a_n2661_45420.t8 212.081
R56489 a_n2661_45420.n3 a_n2661_45420.t9 212.081
R56490 a_n2661_45420.n4 a_n2661_45420.n1 202.663
R56491 a_n2661_45420.n1 a_n2661_45420.t4 196.131
R56492 a_n2661_45420.n6 a_n2661_45420.n5 187.927
R56493 a_n2661_45420.n2 a_n2661_45420.t6 139.78
R56494 a_n2661_45420.n3 a_n2661_45420.t7 139.78
R56495 a_n2661_45420.n3 a_n2661_45420.n2 61.346
R56496 a_n2661_45420.n0 a_n2661_45420.t3 26.5955
R56497 a_n2661_45420.n0 a_n2661_45420.t2 26.5955
R56498 a_n2661_45420.t1 a_n2661_45420.n6 24.9236
R56499 a_n2661_45420.n6 a_n2661_45420.t0 24.9236
R56500 a_n2661_45420.n5 a_n2661_45420.n4 14.0946
R56501 a_n2442_44894.n3 a_n2442_44894.t4 1415.15
R56502 a_n2442_44894.n2 a_n2442_44894.t7 1330.32
R56503 a_n2442_44894.n1 a_n2442_44894.t6 1320.68
R56504 a_n2442_44894.n3 a_n2442_44894.t5 1320.68
R56505 a_n2442_44894.n5 a_n2442_44894.n0 380.32
R56506 a_n2442_44894.n6 a_n2442_44894.n5 185
R56507 a_n2442_44894.n4 a_n2442_44894.n1 161.764
R56508 a_n2442_44894.n4 a_n2442_44894.n3 161.3
R56509 a_n2442_44894.n5 a_n2442_44894.n4 123.016
R56510 a_n2442_44894.n3 a_n2442_44894.n2 84.8325
R56511 a_n2442_44894.n2 a_n2442_44894.n1 84.8325
R56512 a_n2442_44894.n0 a_n2442_44894.t3 26.5955
R56513 a_n2442_44894.n0 a_n2442_44894.t2 26.5955
R56514 a_n2442_44894.n6 a_n2442_44894.t0 24.9236
R56515 a_n2442_44894.t1 a_n2442_44894.n6 24.9236
R56516 C0_dummy_N_btm.n0 C0_dummy_N_btm.t0 104.561
R56517 C0_dummy_N_btm.n0 C0_dummy_N_btm.t1 62.8375
R56518 C0_dummy_N_btm C0_dummy_N_btm.n0 48.3234
R56519 C0_dummy_N_btm C0_dummy_N_btm.n1 8.36925
R56520 C0_dummy_N_btm.n1 C0_dummy_N_btm.t2 5.03712
R56521 C0_dummy_N_btm.n1 C0_dummy_N_btm.t3 4.03712
R56522 a_n1827_45412.n2 a_n1827_45412.n0 329.507
R56523 a_n1827_45412.n4 a_n1827_45412.n3 300.118
R56524 a_n1827_45412.n2 a_n1827_45412.n1 299.834
R56525 a_n1827_45412.n5 a_n1827_45412.t11 276.464
R56526 a_n1827_45412.n10 a_n1827_45412.n9 228.13
R56527 a_n1827_45412.n8 a_n1827_45412.n7 213.678
R56528 a_n1827_45412.n7 a_n1827_45412.t9 212.081
R56529 a_n1827_45412.n6 a_n1827_45412.t8 212.081
R56530 a_n1827_45412.n5 a_n1827_45412.t10 196.131
R56531 a_n1827_45412.n8 a_n1827_45412.n5 185.81
R56532 a_n1827_45412.n7 a_n1827_45412.t13 139.78
R56533 a_n1827_45412.n6 a_n1827_45412.t12 139.78
R56534 a_n1827_45412.n4 a_n1827_45412.n2 79.8031
R56535 a_n1827_45412.n9 a_n1827_45412.n4 64.9023
R56536 a_n1827_45412.n7 a_n1827_45412.n6 61.346
R56537 a_n1827_45412.n3 a_n1827_45412.t3 26.5955
R56538 a_n1827_45412.n3 a_n1827_45412.t2 26.5955
R56539 a_n1827_45412.n1 a_n1827_45412.t5 26.5955
R56540 a_n1827_45412.n1 a_n1827_45412.t4 26.5955
R56541 a_n1827_45412.n0 a_n1827_45412.t7 26.5955
R56542 a_n1827_45412.n0 a_n1827_45412.t6 26.5955
R56543 a_n1827_45412.t1 a_n1827_45412.n10 24.9236
R56544 a_n1827_45412.n10 a_n1827_45412.t0 24.9236
R56545 a_n1827_45412.n9 a_n1827_45412.n8 17.2864
R56546 a_1429_47222.t23 a_1429_47222.t20 378.255
R56547 a_1429_47222.t15 a_1429_47222.t22 378.255
R56548 a_1429_47222.t16 a_1429_47222.t10 378.255
R56549 a_1429_47222.t9 a_1429_47222.t13 378.255
R56550 a_1429_47222.n5 a_1429_47222.t23 359.743
R56551 a_1429_47222.n4 a_1429_47222.t16 350.745
R56552 a_1429_47222.n11 a_1429_47222.t9 342.108
R56553 a_1429_47222.n4 a_1429_47222.t15 330.017
R56554 a_1429_47222.n16 a_1429_47222.n15 296.139
R56555 a_1429_47222.n17 a_1429_47222.n16 269.182
R56556 a_1429_47222.n1 a_1429_47222.t5 267.065
R56557 a_1429_47222.n0 a_1429_47222.t21 241.536
R56558 a_1429_47222.n8 a_1429_47222.t7 234.173
R56559 a_1429_47222.n3 a_1429_47222.t8 231.017
R56560 a_1429_47222.n2 a_1429_47222.t11 230.363
R56561 a_1429_47222.n14 a_1429_47222.n0 198.067
R56562 a_1429_47222.n12 a_1429_47222.t12 196.549
R56563 a_1429_47222.n10 a_1429_47222.n1 194.507
R56564 a_1429_47222.n13 a_1429_47222.n12 182.49
R56565 a_1429_47222.n9 a_1429_47222.n8 179.75
R56566 a_1429_47222.n0 a_1429_47222.t6 169.237
R56567 a_1429_47222.n6 a_1429_47222.n3 165.423
R56568 a_1429_47222.n7 a_1429_47222.n2 163.536
R56569 a_1429_47222.n8 a_1429_47222.t19 161.873
R56570 a_1429_47222.n3 a_1429_47222.t4 158.716
R56571 a_1429_47222.n2 a_1429_47222.t14 158.064
R56572 a_1429_47222.n12 a_1429_47222.t17 148.35
R56573 a_1429_47222.n1 a_1429_47222.t18 148.35
R56574 a_1429_47222.n15 a_1429_47222.t3 26.5955
R56575 a_1429_47222.n15 a_1429_47222.t2 26.5955
R56576 a_1429_47222.n17 a_1429_47222.t0 24.9236
R56577 a_1429_47222.t1 a_1429_47222.n17 24.9236
R56578 a_1429_47222.n10 a_1429_47222.n9 23.8976
R56579 a_1429_47222.n6 a_1429_47222.n5 17.1628
R56580 a_1429_47222.n7 a_1429_47222.n6 14.7203
R56581 a_1429_47222.n13 a_1429_47222.n11 13.0537
R56582 a_1429_47222.n9 a_1429_47222.n7 12.7397
R56583 a_1429_47222.n16 a_1429_47222.n14 11.8141
R56584 a_1429_47222.n14 a_1429_47222.n13 7.84305
R56585 a_1429_47222.n5 a_1429_47222.n4 5.57347
R56586 a_1429_47222.n11 a_1429_47222.n10 4.5005
R56587 C5_N_btm.n1 C5_N_btm.t36 101.204
R56588 C5_N_btm.n2 C5_N_btm.t0 98.0923
R56589 C5_N_btm C5_N_btm.n2 57.6255
R56590 C5_N_btm.n0 C5_N_btm.t37 54.9311
R56591 C5_N_btm.n0 C5_N_btm.t1 47.3635
R56592 C5_N_btm.n2 C5_N_btm.n1 8.08383
R56593 C5_N_btm C5_N_btm.n91 7.49425
R56594 C5_N_btm.n1 C5_N_btm.n0 6.87029
R56595 C5_N_btm.n12 C5_N_btm.t35 5.03712
R56596 C5_N_btm.n84 C5_N_btm.n83 4.60698
R56597 C5_N_btm.n83 C5_N_btm.n82 4.60698
R56598 C5_N_btm.n81 C5_N_btm.n80 4.60698
R56599 C5_N_btm.n80 C5_N_btm.n79 4.60698
R56600 C5_N_btm.n78 C5_N_btm.n77 4.60698
R56601 C5_N_btm.n77 C5_N_btm.n76 4.60698
R56602 C5_N_btm.n75 C5_N_btm.n74 4.60698
R56603 C5_N_btm.n74 C5_N_btm.n73 4.60698
R56604 C5_N_btm.n72 C5_N_btm.n71 4.60698
R56605 C5_N_btm.n71 C5_N_btm.n70 4.60698
R56606 C5_N_btm.n69 C5_N_btm.n68 4.60698
R56607 C5_N_btm.n68 C5_N_btm.n67 4.60698
R56608 C5_N_btm.n66 C5_N_btm.n65 4.60698
R56609 C5_N_btm.n65 C5_N_btm.n64 4.60698
R56610 C5_N_btm.n63 C5_N_btm.n62 4.60698
R56611 C5_N_btm.n62 C5_N_btm.n61 4.60698
R56612 C5_N_btm.n57 C5_N_btm.n56 4.60698
R56613 C5_N_btm.n56 C5_N_btm.n55 4.60698
R56614 C5_N_btm.n54 C5_N_btm.n53 4.60698
R56615 C5_N_btm.n53 C5_N_btm.n52 4.60698
R56616 C5_N_btm.n51 C5_N_btm.n50 4.60698
R56617 C5_N_btm.n50 C5_N_btm.n49 4.60698
R56618 C5_N_btm.n47 C5_N_btm.n46 4.60698
R56619 C5_N_btm.n48 C5_N_btm.n47 4.60698
R56620 C5_N_btm.n44 C5_N_btm.n43 4.60698
R56621 C5_N_btm.n45 C5_N_btm.n44 4.60698
R56622 C5_N_btm.n41 C5_N_btm.n40 4.60698
R56623 C5_N_btm.n42 C5_N_btm.n41 4.60698
R56624 C5_N_btm.n28 C5_N_btm.n27 4.60698
R56625 C5_N_btm.n29 C5_N_btm.n28 4.60698
R56626 C5_N_btm.n25 C5_N_btm.n24 4.60698
R56627 C5_N_btm.n26 C5_N_btm.n25 4.60698
R56628 C5_N_btm.n39 C5_N_btm.n38 4.60698
R56629 C5_N_btm.n38 C5_N_btm.n37 4.60698
R56630 C5_N_btm.n36 C5_N_btm.n35 4.60698
R56631 C5_N_btm.n35 C5_N_btm.n34 4.60698
R56632 C5_N_btm.n12 C5_N_btm.t9 4.03712
R56633 C5_N_btm.n13 C5_N_btm.t4 4.03712
R56634 C5_N_btm.n14 C5_N_btm.t8 4.03712
R56635 C5_N_btm.n15 C5_N_btm.t18 4.03712
R56636 C5_N_btm.n87 C5_N_btm.t20 4.03712
R56637 C5_N_btm.n88 C5_N_btm.t5 4.03712
R56638 C5_N_btm.n89 C5_N_btm.t31 4.03712
R56639 C5_N_btm.n90 C5_N_btm.t10 4.03712
R56640 C5_N_btm.n91 C5_N_btm.t34 4.03712
R56641 C5_N_btm.n60 C5_N_btm.t23 3.98193
R56642 C5_N_btm.n58 C5_N_btm.t14 3.98193
R56643 C5_N_btm.n30 C5_N_btm.t6 3.98193
R56644 C5_N_btm.n23 C5_N_btm.t11 3.98193
R56645 C5_N_btm.n3 C5_N_btm.t15 3.98193
R56646 C5_N_btm.n85 C5_N_btm.t24 3.98193
R56647 C5_N_btm.n83 C5_N_btm.t28 1.67819
R56648 C5_N_btm.n80 C5_N_btm.t22 1.67819
R56649 C5_N_btm.n77 C5_N_btm.t13 1.67819
R56650 C5_N_btm.n74 C5_N_btm.t32 1.67819
R56651 C5_N_btm.n71 C5_N_btm.t3 1.67819
R56652 C5_N_btm.n68 C5_N_btm.t16 1.67819
R56653 C5_N_btm.n65 C5_N_btm.t25 1.67819
R56654 C5_N_btm.n62 C5_N_btm.t7 1.67819
R56655 C5_N_btm.n56 C5_N_btm.t19 1.67819
R56656 C5_N_btm.n53 C5_N_btm.t29 1.67819
R56657 C5_N_btm.n50 C5_N_btm.t33 1.67819
R56658 C5_N_btm.n47 C5_N_btm.t26 1.67819
R56659 C5_N_btm.n44 C5_N_btm.t21 1.67819
R56660 C5_N_btm.n41 C5_N_btm.t27 1.67819
R56661 C5_N_btm.n28 C5_N_btm.t12 1.67819
R56662 C5_N_btm.n25 C5_N_btm.t17 1.67819
R56663 C5_N_btm.n38 C5_N_btm.t2 1.67819
R56664 C5_N_btm.n35 C5_N_btm.t30 1.67819
R56665 C5_N_btm.n23 C5_N_btm.n18 1.05569
R56666 C5_N_btm.n31 C5_N_btm.n30 1.05569
R56667 C5_N_btm.n86 C5_N_btm.n3 1.05569
R56668 C5_N_btm.n59 C5_N_btm.n58 1.05569
R56669 C5_N_btm.n16 C5_N_btm.n11 1.0005
R56670 C5_N_btm.n17 C5_N_btm.n10 1.0005
R56671 C5_N_btm.n18 C5_N_btm.n9 1.0005
R56672 C5_N_btm.n19 C5_N_btm.n8 1.0005
R56673 C5_N_btm.n20 C5_N_btm.n7 1.0005
R56674 C5_N_btm.n21 C5_N_btm.n20 1.0005
R56675 C5_N_btm.n22 C5_N_btm.n19 1.0005
R56676 C5_N_btm.n31 C5_N_btm.n6 1.0005
R56677 C5_N_btm.n32 C5_N_btm.n5 1.0005
R56678 C5_N_btm.n33 C5_N_btm.n4 1.0005
R56679 C5_N_btm.n13 C5_N_btm.n12 1.0005
R56680 C5_N_btm.n14 C5_N_btm.n13 1.0005
R56681 C5_N_btm.n15 C5_N_btm.n14 1.0005
R56682 C5_N_btm.n59 C5_N_btm.n15 1.0005
R56683 C5_N_btm.n87 C5_N_btm.n86 1.0005
R56684 C5_N_btm.n88 C5_N_btm.n87 1.0005
R56685 C5_N_btm.n89 C5_N_btm.n88 1.0005
R56686 C5_N_btm.n90 C5_N_btm.n89 1.0005
R56687 C5_N_btm.n91 C5_N_btm.n90 1.0005
R56688 C5_N_btm.n24 C5_N_btm.n23 0.679419
R56689 C5_N_btm.n30 C5_N_btm.n29 0.679419
R56690 C5_N_btm.n34 C5_N_btm.n3 0.679419
R56691 C5_N_btm.n58 C5_N_btm.n57 0.679419
R56692 C5_N_btm.n61 C5_N_btm.n60 0.679419
R56693 C5_N_btm.n85 C5_N_btm.n84 0.679419
R56694 C5_N_btm.n27 C5_N_btm.n26 0.6255
R56695 C5_N_btm.n37 C5_N_btm.n36 0.6255
R56696 C5_N_btm.n40 C5_N_btm.n39 0.6255
R56697 C5_N_btm.n43 C5_N_btm.n42 0.6255
R56698 C5_N_btm.n46 C5_N_btm.n45 0.6255
R56699 C5_N_btm.n49 C5_N_btm.n48 0.6255
R56700 C5_N_btm.n52 C5_N_btm.n51 0.6255
R56701 C5_N_btm.n55 C5_N_btm.n54 0.6255
R56702 C5_N_btm.n64 C5_N_btm.n63 0.6255
R56703 C5_N_btm.n67 C5_N_btm.n66 0.6255
R56704 C5_N_btm.n70 C5_N_btm.n69 0.6255
R56705 C5_N_btm.n73 C5_N_btm.n72 0.6255
R56706 C5_N_btm.n76 C5_N_btm.n75 0.6255
R56707 C5_N_btm.n79 C5_N_btm.n78 0.6255
R56708 C5_N_btm.n82 C5_N_btm.n81 0.6255
R56709 C5_N_btm.n24 C5_N_btm.n22 0.109875
R56710 C5_N_btm.n26 C5_N_btm.n22 0.109875
R56711 C5_N_btm.n27 C5_N_btm.n21 0.109875
R56712 C5_N_btm.n29 C5_N_btm.n21 0.109875
R56713 C5_N_btm.n36 C5_N_btm.n33 0.109875
R56714 C5_N_btm.n34 C5_N_btm.n33 0.109875
R56715 C5_N_btm.n39 C5_N_btm.n32 0.109875
R56716 C5_N_btm.n37 C5_N_btm.n32 0.109875
R56717 C5_N_btm.n42 C5_N_btm.n31 0.109875
R56718 C5_N_btm.n40 C5_N_btm.n31 0.109875
R56719 C5_N_btm.n45 C5_N_btm.n20 0.109875
R56720 C5_N_btm.n43 C5_N_btm.n20 0.109875
R56721 C5_N_btm.n48 C5_N_btm.n19 0.109875
R56722 C5_N_btm.n46 C5_N_btm.n19 0.109875
R56723 C5_N_btm.n51 C5_N_btm.n18 0.109875
R56724 C5_N_btm.n49 C5_N_btm.n18 0.109875
R56725 C5_N_btm.n54 C5_N_btm.n17 0.109875
R56726 C5_N_btm.n52 C5_N_btm.n17 0.109875
R56727 C5_N_btm.n57 C5_N_btm.n16 0.109875
R56728 C5_N_btm.n55 C5_N_btm.n16 0.109875
R56729 C5_N_btm.n61 C5_N_btm.n11 0.109875
R56730 C5_N_btm.n63 C5_N_btm.n11 0.109875
R56731 C5_N_btm.n64 C5_N_btm.n10 0.109875
R56732 C5_N_btm.n66 C5_N_btm.n10 0.109875
R56733 C5_N_btm.n67 C5_N_btm.n9 0.109875
R56734 C5_N_btm.n69 C5_N_btm.n9 0.109875
R56735 C5_N_btm.n70 C5_N_btm.n8 0.109875
R56736 C5_N_btm.n72 C5_N_btm.n8 0.109875
R56737 C5_N_btm.n73 C5_N_btm.n7 0.109875
R56738 C5_N_btm.n75 C5_N_btm.n7 0.109875
R56739 C5_N_btm.n76 C5_N_btm.n6 0.109875
R56740 C5_N_btm.n78 C5_N_btm.n6 0.109875
R56741 C5_N_btm.n79 C5_N_btm.n5 0.109875
R56742 C5_N_btm.n81 C5_N_btm.n5 0.109875
R56743 C5_N_btm.n82 C5_N_btm.n4 0.109875
R56744 C5_N_btm.n84 C5_N_btm.n4 0.109875
R56745 C5_N_btm.n60 C5_N_btm.n59 0.0556875
R56746 C5_N_btm.n86 C5_N_btm.n85 0.0556875
R56747 a_n2442_43262.n1 a_n2442_43262.t4 687.587
R56748 a_n2442_43262.n1 a_n2442_43262.n0 287.752
R56749 a_n2442_43262.n2 a_n2442_43262.n1 277.568
R56750 a_n2442_43262.n0 a_n2442_43262.t2 26.5955
R56751 a_n2442_43262.n0 a_n2442_43262.t3 26.5955
R56752 a_n2442_43262.t1 a_n2442_43262.n2 24.9236
R56753 a_n2442_43262.n2 a_n2442_43262.t0 24.9236
R56754 a_n1551_44324.n10 a_n1551_44324.n9 329.507
R56755 a_n1551_44324.n8 a_n1551_44324.n7 300.116
R56756 a_n1551_44324.n8 a_n1551_44324.n6 291.81
R56757 a_n1551_44324.n5 a_n1551_44324.n4 291.733
R56758 a_n1551_44324.n0 a_n1551_44324.t10 276.464
R56759 a_n1551_44324.n3 a_n1551_44324.n0 255.665
R56760 a_n1551_44324.n3 a_n1551_44324.n2 229.094
R56761 a_n1551_44324.n2 a_n1551_44324.t12 212.081
R56762 a_n1551_44324.n1 a_n1551_44324.t13 212.081
R56763 a_n1551_44324.n0 a_n1551_44324.t8 196.131
R56764 a_n1551_44324.n2 a_n1551_44324.t9 139.78
R56765 a_n1551_44324.n1 a_n1551_44324.t11 139.78
R56766 a_n1551_44324.n9 a_n1551_44324.n8 79.8031
R56767 a_n1551_44324.n2 a_n1551_44324.n1 61.346
R56768 a_n1551_44324.n4 a_n1551_44324.t7 26.5955
R56769 a_n1551_44324.n4 a_n1551_44324.t6 26.5955
R56770 a_n1551_44324.n7 a_n1551_44324.t5 26.5955
R56771 a_n1551_44324.n7 a_n1551_44324.t4 26.5955
R56772 a_n1551_44324.n10 a_n1551_44324.t1 26.5955
R56773 a_n1551_44324.t0 a_n1551_44324.n10 26.5955
R56774 a_n1551_44324.n6 a_n1551_44324.t2 24.9236
R56775 a_n1551_44324.n6 a_n1551_44324.t3 24.9236
R56776 a_n1551_44324.n5 a_n1551_44324.n3 13.363
R56777 a_n1551_44324.n9 a_n1551_44324.n5 8.10106
R56778 a_n331_42718.n1 a_n331_42718.t1 457.955
R56779 a_n331_42718.n0 a_n331_42718.t2 241.536
R56780 a_n331_42718.n1 a_n331_42718.n0 225.127
R56781 a_n331_42718.t0 a_n331_42718.n1 216.155
R56782 a_n331_42718.n0 a_n331_42718.t3 169.237
R56783 C0_dummy_P_btm.n0 C0_dummy_P_btm.t0 104.561
R56784 C0_dummy_P_btm.n0 C0_dummy_P_btm.t1 62.8375
R56785 C0_dummy_P_btm C0_dummy_P_btm.n0 48.3234
R56786 C0_dummy_P_btm C0_dummy_P_btm.n1 8.36925
R56787 C0_dummy_P_btm.n1 C0_dummy_P_btm.t3 5.03712
R56788 C0_dummy_P_btm.n1 C0_dummy_P_btm.t2 4.03712
R56789 a_n2661_45956.n5 a_n2661_45956.n4 288.598
R56790 a_n2661_45956.n2 a_n2661_45956.t6 276.464
R56791 a_n2661_45956.n6 a_n2661_45956.n5 272.353
R56792 a_n2661_45956.n3 a_n2661_45956.n1 230.446
R56793 a_n2661_45956.n0 a_n2661_45956.t9 212.081
R56794 a_n2661_45956.n1 a_n2661_45956.t8 212.081
R56795 a_n2661_45956.n2 a_n2661_45956.t4 196.131
R56796 a_n2661_45956.n3 a_n2661_45956.n2 178.031
R56797 a_n2661_45956.n0 a_n2661_45956.t7 139.78
R56798 a_n2661_45956.n1 a_n2661_45956.t5 139.78
R56799 a_n2661_45956.n1 a_n2661_45956.n0 61.346
R56800 a_n2661_45956.n5 a_n2661_45956.n3 27.3993
R56801 a_n2661_45956.n4 a_n2661_45956.t3 26.5955
R56802 a_n2661_45956.n4 a_n2661_45956.t2 26.5955
R56803 a_n2661_45956.t1 a_n2661_45956.n6 24.9236
R56804 a_n2661_45956.n6 a_n2661_45956.t0 24.9236
R56805 C1_P_btm.n2 C1_P_btm.t0 102.406
R56806 C1_P_btm.n1 C1_P_btm.t6 101.787
R56807 C1_P_btm.n0 C1_P_btm.t1 54.9098
R56808 C1_P_btm C1_P_btm.n2 47.688
R56809 C1_P_btm.n0 C1_P_btm.t5 47.3635
R56810 C1_P_btm C1_P_btm.n4 8.9005
R56811 C1_P_btm.n2 C1_P_btm.n1 8.33383
R56812 C1_P_btm.n1 C1_P_btm.n0 7.99529
R56813 C1_P_btm.n3 C1_P_btm.t3 5.03712
R56814 C1_P_btm.n3 C1_P_btm.t4 4.03712
R56815 C1_P_btm.n4 C1_P_btm.t2 4.03712
R56816 C1_P_btm.n4 C1_P_btm.n3 1.0005
R56817 a_15163_45670.n9 a_15163_45670.t1 366.548
R56818 a_15163_45670.n1 a_15163_45670.t6 327.99
R56819 a_15163_45670.t0 a_15163_45670.n9 307.562
R56820 a_15163_45670.n7 a_15163_45670.t10 241.536
R56821 a_15163_45670.n4 a_15163_45670.t4 241.536
R56822 a_15163_45670.n1 a_15163_45670.t3 199.457
R56823 a_15163_45670.n8 a_15163_45670.n7 198.03
R56824 a_15163_45670.n3 a_15163_45670.t8 196.549
R56825 a_15163_45670.n0 a_15163_45670.t2 196.549
R56826 a_15163_45670.n5 a_15163_45670.n3 185.927
R56827 a_15163_45670.n2 a_15163_45670.n1 177.088
R56828 a_15163_45670.n2 a_15163_45670.n0 169.512
R56829 a_15163_45670.n7 a_15163_45670.t9 169.237
R56830 a_15163_45670.n4 a_15163_45670.t5 169.237
R56831 a_15163_45670.n5 a_15163_45670.n4 163.046
R56832 a_15163_45670.n3 a_15163_45670.t7 148.35
R56833 a_15163_45670.n0 a_15163_45670.t11 148.35
R56834 a_15163_45670.n9 a_15163_45670.n8 53.7823
R56835 a_15163_45670.n8 a_15163_45670.n6 8.08033
R56836 a_15163_45670.n6 a_15163_45670.n5 8.05815
R56837 a_15163_45670.n6 a_15163_45670.n2 6.50726
R56838 a_n2293_46508.n5 a_n2293_46508.n0 375.949
R56839 a_n2293_46508.n3 a_n2293_46508.t8 276.464
R56840 a_n2293_46508.n4 a_n2293_46508.n2 213.32
R56841 a_n2293_46508.n1 a_n2293_46508.t6 212.081
R56842 a_n2293_46508.n2 a_n2293_46508.t5 212.081
R56843 a_n2293_46508.n4 a_n2293_46508.n3 196.172
R56844 a_n2293_46508.n3 a_n2293_46508.t4 196.131
R56845 a_n2293_46508.n6 a_n2293_46508.n5 185
R56846 a_n2293_46508.n1 a_n2293_46508.t7 139.78
R56847 a_n2293_46508.n2 a_n2293_46508.t9 139.78
R56848 a_n2293_46508.n2 a_n2293_46508.n1 61.346
R56849 a_n2293_46508.n0 a_n2293_46508.t2 26.5955
R56850 a_n2293_46508.n0 a_n2293_46508.t3 26.5955
R56851 a_n2293_46508.n6 a_n2293_46508.t0 24.9236
R56852 a_n2293_46508.t1 a_n2293_46508.n6 24.9236
R56853 a_n2293_46508.n5 a_n2293_46508.n4 23.366
R56854 C6_P_btm.n4 C6_P_btm.t0 97.811
R56855 C6_P_btm.n3 C6_P_btm.t71 68.0518
R56856 C6_P_btm C6_P_btm.n4 59.563
R56857 C6_P_btm.n2 C6_P_btm.n0 45.0311
R56858 C6_P_btm.n2 C6_P_btm.n1 37.4635
R56859 C6_P_btm.n1 C6_P_btm.t73 9.9005
R56860 C6_P_btm.n1 C6_P_btm.t72 9.9005
R56861 C6_P_btm.n0 C6_P_btm.t70 9.9005
R56862 C6_P_btm.n0 C6_P_btm.t69 9.9005
R56863 C6_P_btm.n4 C6_P_btm.n3 8.0005
R56864 C6_P_btm C6_P_btm.n187 7.213
R56865 C6_P_btm.n3 C6_P_btm.n2 6.58904
R56866 C6_P_btm.n183 C6_P_btm.t2 5.03712
R56867 C6_P_btm.n39 C6_P_btm.t3 5.03712
R56868 C6_P_btm.n36 C6_P_btm.t1 5.03712
R56869 C6_P_btm.n162 C6_P_btm.n161 4.60698
R56870 C6_P_btm.n163 C6_P_btm.n162 4.60698
R56871 C6_P_btm.n143 C6_P_btm.n142 4.60698
R56872 C6_P_btm.n144 C6_P_btm.n143 4.60698
R56873 C6_P_btm.n146 C6_P_btm.n145 4.60698
R56874 C6_P_btm.n147 C6_P_btm.n146 4.60698
R56875 C6_P_btm.n149 C6_P_btm.n148 4.60698
R56876 C6_P_btm.n150 C6_P_btm.n149 4.60698
R56877 C6_P_btm.n151 C6_P_btm.n13 4.60698
R56878 C6_P_btm.n152 C6_P_btm.n151 4.60698
R56879 C6_P_btm.n156 C6_P_btm.n155 4.60698
R56880 C6_P_btm.n157 C6_P_btm.n156 4.60698
R56881 C6_P_btm.n159 C6_P_btm.n158 4.60698
R56882 C6_P_btm.n160 C6_P_btm.n159 4.60698
R56883 C6_P_btm.n77 C6_P_btm.n76 4.60698
R56884 C6_P_btm.n76 C6_P_btm.n75 4.60698
R56885 C6_P_btm.n80 C6_P_btm.n79 4.60698
R56886 C6_P_btm.n79 C6_P_btm.n78 4.60698
R56887 C6_P_btm.n83 C6_P_btm.n82 4.60698
R56888 C6_P_btm.n82 C6_P_btm.n81 4.60698
R56889 C6_P_btm.n86 C6_P_btm.n85 4.60698
R56890 C6_P_btm.n85 C6_P_btm.n84 4.60698
R56891 C6_P_btm.n88 C6_P_btm.n87 4.60698
R56892 C6_P_btm.n89 C6_P_btm.n88 4.60698
R56893 C6_P_btm.n91 C6_P_btm.n90 4.60698
R56894 C6_P_btm.n92 C6_P_btm.n91 4.60698
R56895 C6_P_btm.n94 C6_P_btm.n93 4.60698
R56896 C6_P_btm.n95 C6_P_btm.n94 4.60698
R56897 C6_P_btm.n97 C6_P_btm.n96 4.60698
R56898 C6_P_btm.n98 C6_P_btm.n97 4.60698
R56899 C6_P_btm.n62 C6_P_btm.n61 4.60698
R56900 C6_P_btm.n61 C6_P_btm.n60 4.60698
R56901 C6_P_btm.n64 C6_P_btm.n63 4.60698
R56902 C6_P_btm.n65 C6_P_btm.n64 4.60698
R56903 C6_P_btm.n67 C6_P_btm.n66 4.60698
R56904 C6_P_btm.n68 C6_P_btm.n67 4.60698
R56905 C6_P_btm.n104 C6_P_btm.n103 4.60698
R56906 C6_P_btm.n103 C6_P_btm.n102 4.60698
R56907 C6_P_btm.n107 C6_P_btm.n106 4.60698
R56908 C6_P_btm.n106 C6_P_btm.n105 4.60698
R56909 C6_P_btm.n110 C6_P_btm.n109 4.60698
R56910 C6_P_btm.n109 C6_P_btm.n108 4.60698
R56911 C6_P_btm.n113 C6_P_btm.n112 4.60698
R56912 C6_P_btm.n112 C6_P_btm.n111 4.60698
R56913 C6_P_btm.n116 C6_P_btm.n115 4.60698
R56914 C6_P_btm.n115 C6_P_btm.n114 4.60698
R56915 C6_P_btm.n119 C6_P_btm.n118 4.60698
R56916 C6_P_btm.n118 C6_P_btm.n117 4.60698
R56917 C6_P_btm.n122 C6_P_btm.n121 4.60698
R56918 C6_P_btm.n121 C6_P_btm.n120 4.60698
R56919 C6_P_btm.n125 C6_P_btm.n124 4.60698
R56920 C6_P_btm.n124 C6_P_btm.n123 4.60698
R56921 C6_P_btm.n128 C6_P_btm.n127 4.60698
R56922 C6_P_btm.n127 C6_P_btm.n126 4.60698
R56923 C6_P_btm.n131 C6_P_btm.n130 4.60698
R56924 C6_P_btm.n130 C6_P_btm.n129 4.60698
R56925 C6_P_btm.n134 C6_P_btm.n133 4.60698
R56926 C6_P_btm.n133 C6_P_btm.n132 4.60698
R56927 C6_P_btm.n138 C6_P_btm.n137 4.60698
R56928 C6_P_btm.n137 C6_P_btm.n135 4.60698
R56929 C6_P_btm.n187 C6_P_btm.t4 4.03712
R56930 C6_P_btm.n185 C6_P_btm.t44 3.98193
R56931 C6_P_btm.n184 C6_P_btm.t34 3.98193
R56932 C6_P_btm.n180 C6_P_btm.t19 3.98193
R56933 C6_P_btm.n177 C6_P_btm.t15 3.98193
R56934 C6_P_btm.n174 C6_P_btm.t62 3.98193
R56935 C6_P_btm.n171 C6_P_btm.t58 3.98193
R56936 C6_P_btm.n166 C6_P_btm.t24 3.98193
R56937 C6_P_btm.n154 C6_P_btm.t50 3.98193
R56938 C6_P_btm.n99 C6_P_btm.t35 3.98193
R56939 C6_P_btm.n59 C6_P_btm.t42 3.98193
R56940 C6_P_btm.n55 C6_P_btm.t65 3.98193
R56941 C6_P_btm.n52 C6_P_btm.t27 3.98193
R56942 C6_P_btm.n49 C6_P_btm.t67 3.98193
R56943 C6_P_btm.n44 C6_P_btm.t18 3.98193
R56944 C6_P_btm.n41 C6_P_btm.t61 3.98193
R56945 C6_P_btm.n38 C6_P_btm.t31 3.98193
R56946 C6_P_btm.n37 C6_P_btm.t59 3.98193
R56947 C6_P_btm.n42 C6_P_btm.t36 3.98193
R56948 C6_P_btm.n45 C6_P_btm.t64 3.98193
R56949 C6_P_btm.n48 C6_P_btm.t7 3.98193
R56950 C6_P_btm.n51 C6_P_btm.t49 3.98193
R56951 C6_P_btm.n56 C6_P_btm.t38 3.98193
R56952 C6_P_btm.n69 C6_P_btm.t55 3.98193
R56953 C6_P_btm.n101 C6_P_btm.t39 3.98193
R56954 C6_P_btm.n21 C6_P_btm.t14 3.98193
R56955 C6_P_btm.n20 C6_P_btm.t11 3.98193
R56956 C6_P_btm.n136 C6_P_btm.t33 3.98193
R56957 C6_P_btm.n141 C6_P_btm.t20 3.98193
R56958 C6_P_btm.n164 C6_P_btm.t57 3.98193
R56959 C6_P_btm.n167 C6_P_btm.t60 3.98193
R56960 C6_P_btm.n170 C6_P_btm.t13 3.98193
R56961 C6_P_btm.n173 C6_P_btm.t16 3.98193
R56962 C6_P_btm.n178 C6_P_btm.t23 3.98193
R56963 C6_P_btm.n181 C6_P_btm.t29 3.98193
R56964 C6_P_btm.n162 C6_P_btm.t37 1.67819
R56965 C6_P_btm.n143 C6_P_btm.t66 1.67819
R56966 C6_P_btm.n146 C6_P_btm.t46 1.67819
R56967 C6_P_btm.n149 C6_P_btm.t68 1.67819
R56968 C6_P_btm.n151 C6_P_btm.t40 1.67819
R56969 C6_P_btm.n156 C6_P_btm.t28 1.67819
R56970 C6_P_btm.n159 C6_P_btm.t56 1.67819
R56971 C6_P_btm.n76 C6_P_btm.t52 1.67819
R56972 C6_P_btm.n79 C6_P_btm.t32 1.67819
R56973 C6_P_btm.n82 C6_P_btm.t41 1.67819
R56974 C6_P_btm.n85 C6_P_btm.t30 1.67819
R56975 C6_P_btm.n88 C6_P_btm.t47 1.67819
R56976 C6_P_btm.n91 C6_P_btm.t8 1.67819
R56977 C6_P_btm.n94 C6_P_btm.t43 1.67819
R56978 C6_P_btm.n97 C6_P_btm.t54 1.67819
R56979 C6_P_btm.n61 C6_P_btm.t6 1.67819
R56980 C6_P_btm.n64 C6_P_btm.t51 1.67819
R56981 C6_P_btm.n67 C6_P_btm.t45 1.67819
R56982 C6_P_btm.n103 C6_P_btm.t22 1.67819
R56983 C6_P_btm.n106 C6_P_btm.t25 1.67819
R56984 C6_P_btm.n109 C6_P_btm.t63 1.67819
R56985 C6_P_btm.n112 C6_P_btm.t12 1.67819
R56986 C6_P_btm.n115 C6_P_btm.t26 1.67819
R56987 C6_P_btm.n118 C6_P_btm.t17 1.67819
R56988 C6_P_btm.n121 C6_P_btm.t5 1.67819
R56989 C6_P_btm.n124 C6_P_btm.t21 1.67819
R56990 C6_P_btm.n127 C6_P_btm.t9 1.67819
R56991 C6_P_btm.n130 C6_P_btm.t48 1.67819
R56992 C6_P_btm.n133 C6_P_btm.t53 1.67819
R56993 C6_P_btm.n137 C6_P_btm.t10 1.67819
R56994 C6_P_btm.n154 C6_P_btm.n153 1.05569
R56995 C6_P_btm.n70 C6_P_btm.n69 1.05569
R56996 C6_P_btm.n22 C6_P_btm.n21 1.05569
R56997 C6_P_btm.n20 C6_P_btm.n19 1.05569
R56998 C6_P_btm.n136 C6_P_btm.n8 1.05569
R56999 C6_P_btm.n101 C6_P_btm.n100 1.05569
R57000 C6_P_btm.n140 C6_P_btm.n9 1.0005
R57001 C6_P_btm.n14 C6_P_btm.n11 1.0005
R57002 C6_P_btm.n15 C6_P_btm.n10 1.0005
R57003 C6_P_btm.n43 C6_P_btm.n36 1.0005
R57004 C6_P_btm.n40 C6_P_btm.n35 1.0005
R57005 C6_P_btm.n40 C6_P_btm.n39 1.0005
R57006 C6_P_btm.n47 C6_P_btm.n46 1.0005
R57007 C6_P_btm.n46 C6_P_btm.n43 1.0005
R57008 C6_P_btm.n53 C6_P_btm.n50 1.0005
R57009 C6_P_btm.n50 C6_P_btm.n35 1.0005
R57010 C6_P_btm.n57 C6_P_btm.n34 1.0005
R57011 C6_P_btm.n47 C6_P_btm.n34 1.0005
R57012 C6_P_btm.n54 C6_P_btm.n28 1.0005
R57013 C6_P_btm.n54 C6_P_btm.n53 1.0005
R57014 C6_P_btm.n58 C6_P_btm.n29 1.0005
R57015 C6_P_btm.n58 C6_P_btm.n57 1.0005
R57016 C6_P_btm.n33 C6_P_btm.n30 1.0005
R57017 C6_P_btm.n32 C6_P_btm.n31 1.0005
R57018 C6_P_btm.n29 C6_P_btm.n27 1.0005
R57019 C6_P_btm.n30 C6_P_btm.n26 1.0005
R57020 C6_P_btm.n31 C6_P_btm.n25 1.0005
R57021 C6_P_btm.n70 C6_P_btm.n24 1.0005
R57022 C6_P_btm.n71 C6_P_btm.n23 1.0005
R57023 C6_P_btm.n72 C6_P_btm.n22 1.0005
R57024 C6_P_btm.n73 C6_P_btm.n19 1.0005
R57025 C6_P_btm.n74 C6_P_btm.n18 1.0005
R57026 C6_P_btm.n153 C6_P_btm.n12 1.0005
R57027 C6_P_btm.n17 C6_P_btm.n14 1.0005
R57028 C6_P_btm.n16 C6_P_btm.n15 1.0005
R57029 C6_P_btm.n140 C6_P_btm.n139 1.0005
R57030 C6_P_btm.n100 C6_P_btm.n28 1.0005
R57031 C6_P_btm.n165 C6_P_btm.n8 1.0005
R57032 C6_P_btm.n168 C6_P_btm.n165 1.0005
R57033 C6_P_btm.n9 C6_P_btm.n7 1.0005
R57034 C6_P_btm.n172 C6_P_btm.n7 1.0005
R57035 C6_P_btm.n169 C6_P_btm.n168 1.0005
R57036 C6_P_btm.n169 C6_P_btm.n6 1.0005
R57037 C6_P_btm.n175 C6_P_btm.n172 1.0005
R57038 C6_P_btm.n176 C6_P_btm.n175 1.0005
R57039 C6_P_btm.n179 C6_P_btm.n6 1.0005
R57040 C6_P_btm.n182 C6_P_btm.n179 1.0005
R57041 C6_P_btm.n176 C6_P_btm.n5 1.0005
R57042 C6_P_btm.n186 C6_P_btm.n5 1.0005
R57043 C6_P_btm.n183 C6_P_btm.n182 1.0005
R57044 C6_P_btm.n187 C6_P_btm.n186 1.0005
R57045 C6_P_btm.n38 C6_P_btm.n37 0.733338
R57046 C6_P_btm.n42 C6_P_btm.n41 0.733338
R57047 C6_P_btm.n45 C6_P_btm.n44 0.733338
R57048 C6_P_btm.n49 C6_P_btm.n48 0.733338
R57049 C6_P_btm.n52 C6_P_btm.n51 0.733338
R57050 C6_P_btm.n56 C6_P_btm.n55 0.733338
R57051 C6_P_btm.n21 C6_P_btm.n20 0.733338
R57052 C6_P_btm.n167 C6_P_btm.n166 0.733338
R57053 C6_P_btm.n171 C6_P_btm.n170 0.733338
R57054 C6_P_btm.n174 C6_P_btm.n173 0.733338
R57055 C6_P_btm.n178 C6_P_btm.n177 0.733338
R57056 C6_P_btm.n181 C6_P_btm.n180 0.733338
R57057 C6_P_btm.n185 C6_P_btm.n184 0.733338
R57058 C6_P_btm.n155 C6_P_btm.n154 0.679419
R57059 C6_P_btm.n69 C6_P_btm.n68 0.679419
R57060 C6_P_btm.n60 C6_P_btm.n59 0.679419
R57061 C6_P_btm.n138 C6_P_btm.n136 0.679419
R57062 C6_P_btm.n102 C6_P_btm.n101 0.679419
R57063 C6_P_btm.n99 C6_P_btm.n98 0.679419
R57064 C6_P_btm.n142 C6_P_btm.n141 0.679419
R57065 C6_P_btm.n164 C6_P_btm.n163 0.679419
R57066 C6_P_btm.n161 C6_P_btm.n160 0.6255
R57067 C6_P_btm.n158 C6_P_btm.n157 0.6255
R57068 C6_P_btm.n66 C6_P_btm.n65 0.6255
R57069 C6_P_btm.n63 C6_P_btm.n62 0.6255
R57070 C6_P_btm.n135 C6_P_btm.n134 0.6255
R57071 C6_P_btm.n132 C6_P_btm.n131 0.6255
R57072 C6_P_btm.n129 C6_P_btm.n128 0.6255
R57073 C6_P_btm.n126 C6_P_btm.n125 0.6255
R57074 C6_P_btm.n123 C6_P_btm.n122 0.6255
R57075 C6_P_btm.n120 C6_P_btm.n119 0.6255
R57076 C6_P_btm.n117 C6_P_btm.n116 0.6255
R57077 C6_P_btm.n114 C6_P_btm.n113 0.6255
R57078 C6_P_btm.n111 C6_P_btm.n110 0.6255
R57079 C6_P_btm.n108 C6_P_btm.n107 0.6255
R57080 C6_P_btm.n105 C6_P_btm.n104 0.6255
R57081 C6_P_btm.n96 C6_P_btm.n95 0.6255
R57082 C6_P_btm.n93 C6_P_btm.n92 0.6255
R57083 C6_P_btm.n90 C6_P_btm.n89 0.6255
R57084 C6_P_btm.n87 C6_P_btm.n86 0.6255
R57085 C6_P_btm.n84 C6_P_btm.n83 0.6255
R57086 C6_P_btm.n81 C6_P_btm.n80 0.6255
R57087 C6_P_btm.n78 C6_P_btm.n77 0.6255
R57088 C6_P_btm.n75 C6_P_btm.n13 0.6255
R57089 C6_P_btm.n152 C6_P_btm.n150 0.6255
R57090 C6_P_btm.n148 C6_P_btm.n147 0.6255
R57091 C6_P_btm.n145 C6_P_btm.n144 0.6255
R57092 C6_P_btm.n158 C6_P_btm.n10 0.109875
R57093 C6_P_btm.n160 C6_P_btm.n10 0.109875
R57094 C6_P_btm.n155 C6_P_btm.n11 0.109875
R57095 C6_P_btm.n157 C6_P_btm.n11 0.109875
R57096 C6_P_btm.n66 C6_P_btm.n32 0.109875
R57097 C6_P_btm.n68 C6_P_btm.n32 0.109875
R57098 C6_P_btm.n63 C6_P_btm.n33 0.109875
R57099 C6_P_btm.n65 C6_P_btm.n33 0.109875
R57100 C6_P_btm.n60 C6_P_btm.n58 0.109875
R57101 C6_P_btm.n62 C6_P_btm.n58 0.109875
R57102 C6_P_btm.n139 C6_P_btm.n135 0.109875
R57103 C6_P_btm.n139 C6_P_btm.n138 0.109875
R57104 C6_P_btm.n132 C6_P_btm.n16 0.109875
R57105 C6_P_btm.n134 C6_P_btm.n16 0.109875
R57106 C6_P_btm.n129 C6_P_btm.n17 0.109875
R57107 C6_P_btm.n131 C6_P_btm.n17 0.109875
R57108 C6_P_btm.n126 C6_P_btm.n12 0.109875
R57109 C6_P_btm.n128 C6_P_btm.n12 0.109875
R57110 C6_P_btm.n123 C6_P_btm.n18 0.109875
R57111 C6_P_btm.n125 C6_P_btm.n18 0.109875
R57112 C6_P_btm.n120 C6_P_btm.n19 0.109875
R57113 C6_P_btm.n122 C6_P_btm.n19 0.109875
R57114 C6_P_btm.n117 C6_P_btm.n22 0.109875
R57115 C6_P_btm.n119 C6_P_btm.n22 0.109875
R57116 C6_P_btm.n114 C6_P_btm.n23 0.109875
R57117 C6_P_btm.n116 C6_P_btm.n23 0.109875
R57118 C6_P_btm.n111 C6_P_btm.n24 0.109875
R57119 C6_P_btm.n113 C6_P_btm.n24 0.109875
R57120 C6_P_btm.n108 C6_P_btm.n25 0.109875
R57121 C6_P_btm.n110 C6_P_btm.n25 0.109875
R57122 C6_P_btm.n105 C6_P_btm.n26 0.109875
R57123 C6_P_btm.n107 C6_P_btm.n26 0.109875
R57124 C6_P_btm.n102 C6_P_btm.n27 0.109875
R57125 C6_P_btm.n104 C6_P_btm.n27 0.109875
R57126 C6_P_btm.n98 C6_P_btm.n29 0.109875
R57127 C6_P_btm.n96 C6_P_btm.n29 0.109875
R57128 C6_P_btm.n95 C6_P_btm.n30 0.109875
R57129 C6_P_btm.n93 C6_P_btm.n30 0.109875
R57130 C6_P_btm.n92 C6_P_btm.n31 0.109875
R57131 C6_P_btm.n90 C6_P_btm.n31 0.109875
R57132 C6_P_btm.n89 C6_P_btm.n70 0.109875
R57133 C6_P_btm.n87 C6_P_btm.n70 0.109875
R57134 C6_P_btm.n86 C6_P_btm.n71 0.109875
R57135 C6_P_btm.n84 C6_P_btm.n71 0.109875
R57136 C6_P_btm.n83 C6_P_btm.n72 0.109875
R57137 C6_P_btm.n81 C6_P_btm.n72 0.109875
R57138 C6_P_btm.n80 C6_P_btm.n73 0.109875
R57139 C6_P_btm.n78 C6_P_btm.n73 0.109875
R57140 C6_P_btm.n77 C6_P_btm.n74 0.109875
R57141 C6_P_btm.n75 C6_P_btm.n74 0.109875
R57142 C6_P_btm.n153 C6_P_btm.n13 0.109875
R57143 C6_P_btm.n153 C6_P_btm.n152 0.109875
R57144 C6_P_btm.n150 C6_P_btm.n14 0.109875
R57145 C6_P_btm.n148 C6_P_btm.n14 0.109875
R57146 C6_P_btm.n147 C6_P_btm.n15 0.109875
R57147 C6_P_btm.n145 C6_P_btm.n15 0.109875
R57148 C6_P_btm.n144 C6_P_btm.n140 0.109875
R57149 C6_P_btm.n142 C6_P_btm.n140 0.109875
R57150 C6_P_btm.n161 C6_P_btm.n9 0.109875
R57151 C6_P_btm.n163 C6_P_btm.n9 0.109875
R57152 C6_P_btm.n37 C6_P_btm.n36 0.0556875
R57153 C6_P_btm.n39 C6_P_btm.n38 0.0556875
R57154 C6_P_btm.n41 C6_P_btm.n40 0.0556875
R57155 C6_P_btm.n43 C6_P_btm.n42 0.0556875
R57156 C6_P_btm.n46 C6_P_btm.n45 0.0556875
R57157 C6_P_btm.n44 C6_P_btm.n35 0.0556875
R57158 C6_P_btm.n50 C6_P_btm.n49 0.0556875
R57159 C6_P_btm.n48 C6_P_btm.n47 0.0556875
R57160 C6_P_btm.n51 C6_P_btm.n34 0.0556875
R57161 C6_P_btm.n53 C6_P_btm.n52 0.0556875
R57162 C6_P_btm.n55 C6_P_btm.n54 0.0556875
R57163 C6_P_btm.n57 C6_P_btm.n56 0.0556875
R57164 C6_P_btm.n59 C6_P_btm.n28 0.0556875
R57165 C6_P_btm.n100 C6_P_btm.n99 0.0556875
R57166 C6_P_btm.n141 C6_P_btm.n8 0.0556875
R57167 C6_P_btm.n165 C6_P_btm.n164 0.0556875
R57168 C6_P_btm.n166 C6_P_btm.n7 0.0556875
R57169 C6_P_btm.n168 C6_P_btm.n167 0.0556875
R57170 C6_P_btm.n170 C6_P_btm.n169 0.0556875
R57171 C6_P_btm.n172 C6_P_btm.n171 0.0556875
R57172 C6_P_btm.n175 C6_P_btm.n174 0.0556875
R57173 C6_P_btm.n173 C6_P_btm.n6 0.0556875
R57174 C6_P_btm.n179 C6_P_btm.n178 0.0556875
R57175 C6_P_btm.n177 C6_P_btm.n176 0.0556875
R57176 C6_P_btm.n180 C6_P_btm.n5 0.0556875
R57177 C6_P_btm.n182 C6_P_btm.n181 0.0556875
R57178 C6_P_btm.n184 C6_P_btm.n183 0.0556875
R57179 C6_P_btm.n186 C6_P_btm.n185 0.0556875
R57180 EN_VIN_BSTR_N.n20 EN_VIN_BSTR_N.t21 1559.46
R57181 EN_VIN_BSTR_N.n19 EN_VIN_BSTR_N.t22 1415.15
R57182 EN_VIN_BSTR_N.n19 EN_VIN_BSTR_N.t11 1320.68
R57183 EN_VIN_BSTR_N.n4 EN_VIN_BSTR_N.t9 748.122
R57184 EN_VIN_BSTR_N.n4 EN_VIN_BSTR_N.t17 678.014
R57185 EN_VIN_BSTR_N.n11 EN_VIN_BSTR_N.t7 605.802
R57186 EN_VIN_BSTR_N.n10 EN_VIN_BSTR_N.t12 444.502
R57187 EN_VIN_BSTR_N.n5 EN_VIN_BSTR_N.t19 398.577
R57188 EN_VIN_BSTR_N.n9 EN_VIN_BSTR_N.t15 382.812
R57189 EN_VIN_BSTR_N.n17 EN_VIN_BSTR_N.t16 381.798
R57190 EN_VIN_BSTR_N.n9 EN_VIN_BSTR_N.t18 381.793
R57191 EN_VIN_BSTR_N.n16 EN_VIN_BSTR_N.t23 381.788
R57192 EN_VIN_BSTR_N.n15 EN_VIN_BSTR_N.t10 381.413
R57193 EN_VIN_BSTR_N.n14 EN_VIN_BSTR_N.t20 381.413
R57194 EN_VIN_BSTR_N.n13 EN_VIN_BSTR_N.t14 381.413
R57195 EN_VIN_BSTR_N.n12 EN_VIN_BSTR_N.t13 381.413
R57196 EN_VIN_BSTR_N.n10 EN_VIN_BSTR_N.t8 356.68
R57197 EN_VIN_BSTR_N.n5 EN_VIN_BSTR_N.n4 176.418
R57198 EN_VIN_BSTR_N.n11 EN_VIN_BSTR_N.n10 161.768
R57199 EN_VIN_BSTR_N.n20 EN_VIN_BSTR_N.n19 161.3
R57200 EN_VIN_BSTR_N.n7 EN_VIN_BSTR_N.n2 56.3527
R57201 EN_VIN_BSTR_N.n6 EN_VIN_BSTR_N.n3 56.3527
R57202 EN_VIN_BSTR_N.n21 EN_VIN_BSTR_N.n18 28.2777
R57203 EN_VIN_BSTR_N.n0 EN_VIN_BSTR_N.t4 24.8246
R57204 EN_VIN_BSTR_N.n0 EN_VIN_BSTR_N.t6 24.1869
R57205 EN_VIN_BSTR_N.n1 EN_VIN_BSTR_N.t5 24.1612
R57206 EN_VIN_BSTR_N EN_VIN_BSTR_N.n21 22.2703
R57207 EN_VIN_BSTR_N EN_VIN_BSTR_N.n8 8.3965
R57208 EN_VIN_BSTR_N.n3 EN_VIN_BSTR_N.t1 8.12675
R57209 EN_VIN_BSTR_N.n3 EN_VIN_BSTR_N.t2 8.12675
R57210 EN_VIN_BSTR_N.n2 EN_VIN_BSTR_N.t0 8.12675
R57211 EN_VIN_BSTR_N.n2 EN_VIN_BSTR_N.t3 8.12675
R57212 EN_VIN_BSTR_N.n21 EN_VIN_BSTR_N.n20 4.51508
R57213 EN_VIN_BSTR_N.n6 EN_VIN_BSTR_N.n5 2.39112
R57214 EN_VIN_BSTR_N.n1 EN_VIN_BSTR_N.n0 0.989971
R57215 EN_VIN_BSTR_N.n17 EN_VIN_BSTR_N.n16 0.9005
R57216 EN_VIN_BSTR_N.n8 EN_VIN_BSTR_N.n7 0.888337
R57217 EN_VIN_BSTR_N.n18 EN_VIN_BSTR_N.n17 0.7005
R57218 EN_VIN_BSTR_N.n13 EN_VIN_BSTR_N.n12 0.512318
R57219 EN_VIN_BSTR_N.n14 EN_VIN_BSTR_N.n13 0.512318
R57220 EN_VIN_BSTR_N.n15 EN_VIN_BSTR_N.n14 0.512318
R57221 EN_VIN_BSTR_N.n7 EN_VIN_BSTR_N.n6 0.462038
R57222 EN_VIN_BSTR_N.n18 EN_VIN_BSTR_N.n9 0.3755
R57223 EN_VIN_BSTR_N.n12 EN_VIN_BSTR_N.n11 0.267318
R57224 EN_VIN_BSTR_N.n16 EN_VIN_BSTR_N.n15 0.138909
R57225 EN_VIN_BSTR_N.n8 EN_VIN_BSTR_N.n1 0.003
R57226 VIN_N.n1 VIN_N.t0 92.1604
R57227 VIN_N.n3 VIN_N.t11 91.0227
R57228 VIN_N.n7 VIN_N.t3 90.7102
R57229 VIN_N.n6 VIN_N.t2 90.7102
R57230 VIN_N.n5 VIN_N.t12 90.7102
R57231 VIN_N.n4 VIN_N.t10 90.7102
R57232 VIN_N.n1 VIN_N.t13 90.6265
R57233 VIN_N.n2 VIN_N.t1 90.6219
R57234 VIN_N.n10 VIN_N.t8 47.4586
R57235 VIN_N.n9 VIN_N.n8 37.5586
R57236 VIN_N.n14 VIN_N.n12 32.094
R57237 VIN_N.n13 VIN_N.t15 25.3459
R57238 VIN_N.n13 VIN_N.t14 25.1227
R57239 VIN_N.n14 VIN_N.n13 17.3942
R57240 VIN_N.n12 VIN_N.t4 16.5266
R57241 VIN_N.n11 VIN_N.n0 14.0516
R57242 VIN_N.n11 VIN_N.n10 11.2899
R57243 VIN_N VIN_N.n14 10.1221
R57244 VIN_N.n8 VIN_N.t7 9.9005
R57245 VIN_N.n8 VIN_N.t9 9.9005
R57246 VIN_N.n0 VIN_N.t5 2.4755
R57247 VIN_N.n0 VIN_N.t6 2.4755
R57248 VIN_N.n2 VIN_N.n1 1.6255
R57249 VIN_N.n3 VIN_N.n2 1.2505
R57250 VIN_N.n9 VIN_N.n7 0.8755
R57251 VIN_N.n5 VIN_N.n4 0.563
R57252 VIN_N.n6 VIN_N.n5 0.563
R57253 VIN_N.n7 VIN_N.n6 0.563
R57254 VIN_N.n10 VIN_N.n9 0.453625
R57255 VIN_N.n12 VIN_N.n11 0.438
R57256 VIN_N.n4 VIN_N.n3 0.2505
R57257 a_7754_40130.t11 a_7754_40130.n24 578.173
R57258 a_7754_40130.n6 a_7754_40130.t12 578.173
R57259 a_7754_40130.n7 a_7754_40130.t12 578.173
R57260 a_7754_40130.n25 a_7754_40130.t11 577.779
R57261 a_7754_40130.t9 a_7754_40130.n0 577.749
R57262 a_7754_40130.n24 a_7754_40130.t9 577.749
R57263 a_7754_40130.t13 a_7754_40130.n22 577.749
R57264 a_7754_40130.n23 a_7754_40130.t13 577.749
R57265 a_7754_40130.n21 a_7754_40130.t4 577.749
R57266 a_7754_40130.t4 a_7754_40130.n1 577.749
R57267 a_7754_40130.n20 a_7754_40130.t14 577.749
R57268 a_7754_40130.t14 a_7754_40130.n19 577.749
R57269 a_7754_40130.t8 a_7754_40130.n2 577.749
R57270 a_7754_40130.n18 a_7754_40130.t8 577.749
R57271 a_7754_40130.n14 a_7754_40130.t1 577.749
R57272 a_7754_40130.t1 a_7754_40130.n3 577.749
R57273 a_7754_40130.n13 a_7754_40130.t10 577.749
R57274 a_7754_40130.t10 a_7754_40130.n12 577.749
R57275 a_7754_40130.t15 a_7754_40130.n4 577.749
R57276 a_7754_40130.n11 a_7754_40130.t15 577.749
R57277 a_7754_40130.t5 a_7754_40130.n9 577.749
R57278 a_7754_40130.n10 a_7754_40130.t5 577.749
R57279 a_7754_40130.n8 a_7754_40130.t7 577.749
R57280 a_7754_40130.t7 a_7754_40130.n5 577.749
R57281 a_7754_40130.n7 a_7754_40130.t6 577.749
R57282 a_7754_40130.t6 a_7754_40130.n6 577.749
R57283 a_7754_40130.n26 a_7754_40130.t3 233.501
R57284 a_7754_40130.t0 a_7754_40130.n26 48.462
R57285 a_7754_40130.n16 a_7754_40130.t2 29.4286
R57286 a_7754_40130.n26 a_7754_40130.n25 9.38245
R57287 a_7754_40130.n17 a_7754_40130.n16 2.29004
R57288 a_7754_40130.n16 a_7754_40130.n15 2.27754
R57289 a_7754_40130.n6 a_7754_40130.n5 0.4255
R57290 a_7754_40130.n10 a_7754_40130.n5 0.4255
R57291 a_7754_40130.n11 a_7754_40130.n10 0.4255
R57292 a_7754_40130.n12 a_7754_40130.n11 0.4255
R57293 a_7754_40130.n12 a_7754_40130.n3 0.4255
R57294 a_7754_40130.n19 a_7754_40130.n18 0.4255
R57295 a_7754_40130.n19 a_7754_40130.n1 0.4255
R57296 a_7754_40130.n23 a_7754_40130.n1 0.4255
R57297 a_7754_40130.n24 a_7754_40130.n23 0.4255
R57298 a_7754_40130.n8 a_7754_40130.n7 0.4255
R57299 a_7754_40130.n9 a_7754_40130.n8 0.4255
R57300 a_7754_40130.n9 a_7754_40130.n4 0.4255
R57301 a_7754_40130.n13 a_7754_40130.n4 0.4255
R57302 a_7754_40130.n14 a_7754_40130.n13 0.4255
R57303 a_7754_40130.n20 a_7754_40130.n2 0.4255
R57304 a_7754_40130.n21 a_7754_40130.n20 0.4255
R57305 a_7754_40130.n22 a_7754_40130.n21 0.4255
R57306 a_7754_40130.n22 a_7754_40130.n0 0.4255
R57307 a_7754_40130.n25 a_7754_40130.n0 0.395812
R57308 a_7754_40130.n18 a_7754_40130.n17 0.303625
R57309 a_7754_40130.n15 a_7754_40130.n2 0.303625
R57310 a_7754_40130.n17 a_7754_40130.n3 0.122375
R57311 a_7754_40130.n15 a_7754_40130.n14 0.122375
R57312 a_11206_38545.n2 a_11206_38545.n1 225.84
R57313 a_11206_38545.n0 a_11206_38545.t3 39.2429
R57314 a_11206_38545.n0 a_11206_38545.t2 34.125
R57315 a_11206_38545.n1 a_11206_38545.t1 34.125
R57316 a_11206_38545.n2 a_11206_38545.t4 28.5655
R57317 a_11206_38545.t0 a_11206_38545.n2 28.5655
R57318 a_11206_38545.n1 a_11206_38545.n0 0.563
R57319 a_n1827_44324.n5 a_n1827_44324.n0 664.928
R57320 a_n1827_44324.n4 a_n1827_44324.n1 278.68
R57321 a_n1827_44324.n1 a_n1827_44324.t9 276.464
R57322 a_n1827_44324.n4 a_n1827_44324.n3 237.296
R57323 a_n1827_44324.n3 a_n1827_44324.t6 212.081
R57324 a_n1827_44324.n2 a_n1827_44324.t5 212.081
R57325 a_n1827_44324.n1 a_n1827_44324.t7 196.131
R57326 a_n1827_44324.n6 a_n1827_44324.n5 187.927
R57327 a_n1827_44324.n3 a_n1827_44324.t8 139.78
R57328 a_n1827_44324.n2 a_n1827_44324.t4 139.78
R57329 a_n1827_44324.n3 a_n1827_44324.n2 61.346
R57330 a_n1827_44324.n0 a_n1827_44324.t3 26.5955
R57331 a_n1827_44324.n0 a_n1827_44324.t2 26.5955
R57332 a_n1827_44324.t1 a_n1827_44324.n6 24.9236
R57333 a_n1827_44324.n6 a_n1827_44324.t0 24.9236
R57334 a_n1827_44324.n5 a_n1827_44324.n4 9.3005
R57335 a_2755_43494.n20 a_2755_43494.n19 287.752
R57336 a_2755_43494.n21 a_2755_43494.n20 277.568
R57337 a_2755_43494.n16 a_2755_43494.t10 239.505
R57338 a_2755_43494.n2 a_2755_43494.t16 239.505
R57339 a_2755_43494.n3 a_2755_43494.t13 239.505
R57340 a_2755_43494.n11 a_2755_43494.t20 239.505
R57341 a_2755_43494.n8 a_2755_43494.t8 239.505
R57342 a_2755_43494.n6 a_2755_43494.t23 239.505
R57343 a_2755_43494.n5 a_2755_43494.t19 239.505
R57344 a_2755_43494.n1 a_2755_43494.t22 239.505
R57345 a_2755_43494.n0 a_2755_43494.t21 239.505
R57346 a_2755_43494.n4 a_2755_43494.t18 231.017
R57347 a_2755_43494.n7 a_2755_43494.n5 194.73
R57348 a_2755_43494.n12 a_2755_43494.n11 190.78
R57349 a_2755_43494.n18 a_2755_43494.n0 187.512
R57350 a_2755_43494.n7 a_2755_43494.n6 175.958
R57351 a_2755_43494.n9 a_2755_43494.n8 175.66
R57352 a_2755_43494.n15 a_2755_43494.n1 175.088
R57353 a_2755_43494.n10 a_2755_43494.n4 172.714
R57354 a_2755_43494.n14 a_2755_43494.n2 169.702
R57355 a_2755_43494.n13 a_2755_43494.n3 169.702
R57356 a_2755_43494.n17 a_2755_43494.n16 169.514
R57357 a_2755_43494.n16 a_2755_43494.t9 167.204
R57358 a_2755_43494.n2 a_2755_43494.t11 167.204
R57359 a_2755_43494.n3 a_2755_43494.t4 167.204
R57360 a_2755_43494.n11 a_2755_43494.t14 167.204
R57361 a_2755_43494.n8 a_2755_43494.t5 167.204
R57362 a_2755_43494.n6 a_2755_43494.t7 167.204
R57363 a_2755_43494.n5 a_2755_43494.t6 167.204
R57364 a_2755_43494.n1 a_2755_43494.t17 167.204
R57365 a_2755_43494.n0 a_2755_43494.t15 167.204
R57366 a_2755_43494.n4 a_2755_43494.t12 158.716
R57367 a_2755_43494.n20 a_2755_43494.n18 36.091
R57368 a_2755_43494.n19 a_2755_43494.t2 26.5955
R57369 a_2755_43494.n19 a_2755_43494.t3 26.5955
R57370 a_2755_43494.n15 a_2755_43494.n14 25.2423
R57371 a_2755_43494.n21 a_2755_43494.t0 24.9236
R57372 a_2755_43494.t1 a_2755_43494.n21 24.9236
R57373 a_2755_43494.n13 a_2755_43494.n12 19.6956
R57374 a_2755_43494.n17 a_2755_43494.n15 17.5799
R57375 a_2755_43494.n10 a_2755_43494.n9 16.2615
R57376 a_2755_43494.n9 a_2755_43494.n7 7.80678
R57377 a_2755_43494.n18 a_2755_43494.n17 3.81896
R57378 a_2755_43494.n14 a_2755_43494.n13 3.69693
R57379 a_2755_43494.n12 a_2755_43494.n10 2.2972
R57380 a_1847_45528.n4 a_1847_45528.t23 334.723
R57381 a_1847_45528.n15 a_1847_45528.t21 256.716
R57382 a_1847_45528.n3 a_1847_45528.n1 248.087
R57383 a_1847_45528.n5 a_1847_45528.t14 241.536
R57384 a_1847_45528.n11 a_1847_45528.t24 241.536
R57385 a_1847_45528.n9 a_1847_45528.t27 238.397
R57386 a_1847_45528.n16 a_1847_45528.t22 231.835
R57387 a_1847_45528.n6 a_1847_45528.t18 221.72
R57388 a_1847_45528.n7 a_1847_45528.t8 221.72
R57389 a_1847_45528.n3 a_1847_45528.n2 208.507
R57390 a_1847_45528.n4 a_1847_45528.t10 206.19
R57391 a_1847_45528.n10 a_1847_45528.t9 206.19
R57392 a_1847_45528.n9 a_1847_45528.t16 195.017
R57393 a_1847_45528.n19 a_1847_45528.n9 176.345
R57394 a_1847_45528.n21 a_1847_45528.n5 173.359
R57395 a_1847_45528.n14 a_1847_45528.n10 170.994
R57396 a_1847_45528.n5 a_1847_45528.t11 169.237
R57397 a_1847_45528.n11 a_1847_45528.t13 169.237
R57398 a_1847_45528.n20 a_1847_45528.n8 166.288
R57399 a_1847_45528.n17 a_1847_45528.n15 164.831
R57400 a_1847_45528.n13 a_1847_45528.n12 164.379
R57401 a_1847_45528.n17 a_1847_45528.n16 163.643
R57402 a_1847_45528.n22 a_1847_45528.n4 162.752
R57403 a_1847_45528.n13 a_1847_45528.n11 162.286
R57404 a_1847_45528.n15 a_1847_45528.t25 161.275
R57405 a_1847_45528.n16 a_1847_45528.t26 157.07
R57406 a_1847_45528.n6 a_1847_45528.t15 149.421
R57407 a_1847_45528.n7 a_1847_45528.t19 149.421
R57408 a_1847_45528.n10 a_1847_45528.t17 148.35
R57409 a_1847_45528.n24 a_1847_45528.n0 137.576
R57410 a_1847_45528.n12 a_1847_45528.t20 137.177
R57411 a_1847_45528.n12 a_1847_45528.t12 121.109
R57412 a_1847_45528.n25 a_1847_45528.n24 99.1759
R57413 a_1847_45528.n8 a_1847_45528.n6 37.4894
R57414 a_1847_45528.n8 a_1847_45528.n7 37.4894
R57415 a_1847_45528.n24 a_1847_45528.n23 36.0958
R57416 a_1847_45528.n1 a_1847_45528.t4 26.5955
R57417 a_1847_45528.n1 a_1847_45528.t5 26.5955
R57418 a_1847_45528.n2 a_1847_45528.t7 26.5955
R57419 a_1847_45528.n2 a_1847_45528.t6 26.5955
R57420 a_1847_45528.n0 a_1847_45528.t1 24.9236
R57421 a_1847_45528.n0 a_1847_45528.t0 24.9236
R57422 a_1847_45528.t3 a_1847_45528.n25 24.9236
R57423 a_1847_45528.n25 a_1847_45528.t2 24.9236
R57424 a_1847_45528.n23 a_1847_45528.n22 20.9461
R57425 a_1847_45528.n23 a_1847_45528.n3 17.2539
R57426 a_1847_45528.n18 a_1847_45528.n17 12.0032
R57427 a_1847_45528.n14 a_1847_45528.n13 10.154
R57428 a_1847_45528.n22 a_1847_45528.n21 9.63099
R57429 a_1847_45528.n18 a_1847_45528.n14 5.02935
R57430 a_1847_45528.n19 a_1847_45528.n18 4.5005
R57431 a_1847_45528.n20 a_1847_45528.n19 4.04171
R57432 a_1847_45528.n21 a_1847_45528.n20 1.64336
R57433 a_4000_42718.n2 a_4000_42718.t7 581.006
R57434 a_4000_42718.n2 a_4000_42718.t6 579.977
R57435 a_4000_42718.n4 a_4000_42718.n0 380.32
R57436 a_4000_42718.n1 a_4000_42718.t4 260.322
R57437 a_4000_42718.n5 a_4000_42718.n4 185
R57438 a_4000_42718.n1 a_4000_42718.t5 175.169
R57439 a_4000_42718.n3 a_4000_42718.n1 170.712
R57440 a_4000_42718.n3 a_4000_42718.n2 107.648
R57441 a_4000_42718.n0 a_4000_42718.t3 26.5955
R57442 a_4000_42718.n0 a_4000_42718.t2 26.5955
R57443 a_4000_42718.t1 a_4000_42718.n5 24.9236
R57444 a_4000_42718.n5 a_4000_42718.t0 24.9236
R57445 a_4000_42718.n4 a_4000_42718.n3 21.8317
R57446 C3_P_btm.n1 C3_P_btm.t1 101.516
R57447 C3_P_btm.n2 C3_P_btm.t0 100.142
R57448 C3_P_btm.n0 C3_P_btm.t2 54.9311
R57449 C3_P_btm C3_P_btm.n2 47.8026
R57450 C3_P_btm.n0 C3_P_btm.t12 47.3635
R57451 C3_P_btm.n2 C3_P_btm.n1 9.7505
R57452 C3_P_btm C3_P_btm.n10 9.18175
R57453 C3_P_btm.n1 C3_P_btm.n0 7.43279
R57454 C3_P_btm.n3 C3_P_btm.t6 4.76719
R57455 C3_P_btm.n8 C3_P_btm.t8 4.03712
R57456 C3_P_btm.n9 C3_P_btm.t7 4.03712
R57457 C3_P_btm.n10 C3_P_btm.t3 4.03712
R57458 C3_P_btm.n7 C3_P_btm.t11 3.98193
R57459 C3_P_btm.n6 C3_P_btm.t4 3.92851
R57460 C3_P_btm.n5 C3_P_btm.t9 3.92851
R57461 C3_P_btm.n4 C3_P_btm.t10 3.92851
R57462 C3_P_btm.n3 C3_P_btm.t5 3.92851
R57463 C3_P_btm.n8 C3_P_btm.n7 1.05569
R57464 C3_P_btm.n9 C3_P_btm.n8 1.0005
R57465 C3_P_btm.n10 C3_P_btm.n9 1.0005
R57466 C3_P_btm.n4 C3_P_btm.n3 0.840176
R57467 C3_P_btm.n5 C3_P_btm.n4 0.840176
R57468 C3_P_btm.n6 C3_P_btm.n5 0.840176
R57469 C3_P_btm.n7 C3_P_btm.n6 0.786757
R57470 a_2587_44868.n29 a_2587_44868.t18 722.096
R57471 a_2587_44868.n6 a_2587_44868.t20 722.096
R57472 a_2587_44868.n24 a_2587_44868.t26 722.096
R57473 a_2587_44868.n18 a_2587_44868.t9 722.096
R57474 a_2587_44868.n19 a_2587_44868.t12 722.096
R57475 a_2587_44868.n20 a_2587_44868.t19 722.096
R57476 a_2587_44868.n16 a_2587_44868.t13 722.096
R57477 a_2587_44868.n27 a_2587_44868.t11 722.096
R57478 a_2587_44868.n2 a_2587_44868.n0 647.148
R57479 a_2587_44868.n5 a_2587_44868.t14 231.017
R57480 a_2587_44868.n8 a_2587_44868.t31 212.081
R57481 a_2587_44868.n10 a_2587_44868.t30 212.081
R57482 a_2587_44868.n12 a_2587_44868.t32 212.081
R57483 a_2587_44868.n13 a_2587_44868.t24 212.081
R57484 a_2587_44868.n4 a_2587_44868.n3 200.262
R57485 a_2587_44868.n2 a_2587_44868.n1 194.441
R57486 a_2587_44868.n33 a_2587_44868.n32 185
R57487 a_2587_44868.n30 a_2587_44868.n29 182.946
R57488 a_2587_44868.n21 a_2587_44868.n20 180.119
R57489 a_2587_44868.n31 a_2587_44868.n5 179.516
R57490 a_2587_44868.n22 a_2587_44868.n18 178.042
R57491 a_2587_44868.n28 a_2587_44868.n27 174.41
R57492 a_2587_44868.n17 a_2587_44868.n16 172.516
R57493 a_2587_44868.n15 a_2587_44868.n14 170.945
R57494 a_2587_44868.n26 a_2587_44868.n6 169.314
R57495 a_2587_44868.n25 a_2587_44868.n24 168.016
R57496 a_2587_44868.n21 a_2587_44868.n19 168.016
R57497 a_2587_44868.n29 a_2587_44868.t29 162.963
R57498 a_2587_44868.n6 a_2587_44868.t16 162.963
R57499 a_2587_44868.n24 a_2587_44868.t17 162.963
R57500 a_2587_44868.n18 a_2587_44868.t23 162.963
R57501 a_2587_44868.n19 a_2587_44868.t10 162.963
R57502 a_2587_44868.n20 a_2587_44868.t27 162.963
R57503 a_2587_44868.n16 a_2587_44868.t21 162.963
R57504 a_2587_44868.n27 a_2587_44868.t22 162.963
R57505 a_2587_44868.n5 a_2587_44868.t25 158.716
R57506 a_2587_44868.n11 a_2587_44868.n7 152
R57507 a_2587_44868.n8 a_2587_44868.t28 139.78
R57508 a_2587_44868.n10 a_2587_44868.t8 139.78
R57509 a_2587_44868.n12 a_2587_44868.t15 139.78
R57510 a_2587_44868.n13 a_2587_44868.t33 139.78
R57511 a_2587_44868.n9 a_2587_44868.n7 101.177
R57512 a_2587_44868.n32 a_2587_44868.n4 58.6278
R57513 a_2587_44868.n4 a_2587_44868.n2 50.5705
R57514 a_2587_44868.n10 a_2587_44868.n9 42.8185
R57515 a_2587_44868.n3 a_2587_44868.t0 40.0005
R57516 a_2587_44868.n3 a_2587_44868.t2 40.0005
R57517 a_2587_44868.n33 a_2587_44868.t1 40.0005
R57518 a_2587_44868.t3 a_2587_44868.n33 40.0005
R57519 a_2587_44868.n31 a_2587_44868.n30 35.6186
R57520 a_2587_44868.n11 a_2587_44868.n10 30.6732
R57521 a_2587_44868.n12 a_2587_44868.n11 30.6732
R57522 a_2587_44868.n14 a_2587_44868.n12 30.6732
R57523 a_2587_44868.n14 a_2587_44868.n13 30.6732
R57524 a_2587_44868.n1 a_2587_44868.t7 27.5805
R57525 a_2587_44868.n1 a_2587_44868.t6 27.5805
R57526 a_2587_44868.n0 a_2587_44868.t4 27.5805
R57527 a_2587_44868.n0 a_2587_44868.t5 27.5805
R57528 a_2587_44868.n32 a_2587_44868.n31 23.5699
R57529 a_2587_44868.n30 a_2587_44868.n28 18.5335
R57530 a_2587_44868.n17 a_2587_44868.n15 16.3858
R57531 a_2587_44868.n9 a_2587_44868.n8 16.0782
R57532 a_2587_44868.n28 a_2587_44868.n26 15.8102
R57533 a_2587_44868.n25 a_2587_44868.n23 14.6258
R57534 a_2587_44868.n23 a_2587_44868.n22 8.40127
R57535 a_2587_44868.n22 a_2587_44868.n21 6.93233
R57536 a_2587_44868.n26 a_2587_44868.n25 2.58681
R57537 a_2587_44868.n15 a_2587_44868.n7 2.5605
R57538 a_2587_44868.n23 a_2587_44868.n17 2.12876
R57539 a_1203_42692.n28 a_1203_42692.n26 252.931
R57540 a_1203_42692.n23 a_1203_42692.t17 230.363
R57541 a_1203_42692.n19 a_1203_42692.t15 230.363
R57542 a_1203_42692.n17 a_1203_42692.t8 230.363
R57543 a_1203_42692.n15 a_1203_42692.t28 230.363
R57544 a_1203_42692.n13 a_1203_42692.t33 230.363
R57545 a_1203_42692.n11 a_1203_42692.t27 230.363
R57546 a_1203_42692.n8 a_1203_42692.t13 230.363
R57547 a_1203_42692.n5 a_1203_42692.t29 230.363
R57548 a_1203_42692.n2 a_1203_42692.t11 230.363
R57549 a_1203_42692.n1 a_1203_42692.t20 230.363
R57550 a_1203_42692.n21 a_1203_42692.t16 230.363
R57551 a_1203_42692.n6 a_1203_42692.n4 213.519
R57552 a_1203_42692.n3 a_1203_42692.t14 212.081
R57553 a_1203_42692.n4 a_1203_42692.t18 212.081
R57554 a_1203_42692.n28 a_1203_42692.n27 208.507
R57555 a_1203_42692.n9 a_1203_42692.n8 176.423
R57556 a_1203_42692.n12 a_1203_42692.n11 168.143
R57557 a_1203_42692.n24 a_1203_42692.n23 167.849
R57558 a_1203_42692.n22 a_1203_42692.n21 166.998
R57559 a_1203_42692.n16 a_1203_42692.n15 166.421
R57560 a_1203_42692.n6 a_1203_42692.n5 164.536
R57561 a_1203_42692.n7 a_1203_42692.n2 163.536
R57562 a_1203_42692.n10 a_1203_42692.n1 163.536
R57563 a_1203_42692.n20 a_1203_42692.n19 163.349
R57564 a_1203_42692.n18 a_1203_42692.n17 163.349
R57565 a_1203_42692.n14 a_1203_42692.n13 163.349
R57566 a_1203_42692.n23 a_1203_42692.t22 158.064
R57567 a_1203_42692.n19 a_1203_42692.t9 158.064
R57568 a_1203_42692.n17 a_1203_42692.t23 158.064
R57569 a_1203_42692.n15 a_1203_42692.t31 158.064
R57570 a_1203_42692.n13 a_1203_42692.t12 158.064
R57571 a_1203_42692.n11 a_1203_42692.t25 158.064
R57572 a_1203_42692.n8 a_1203_42692.t21 158.064
R57573 a_1203_42692.n5 a_1203_42692.t10 158.064
R57574 a_1203_42692.n2 a_1203_42692.t26 158.064
R57575 a_1203_42692.n1 a_1203_42692.t30 158.064
R57576 a_1203_42692.n21 a_1203_42692.t24 158.064
R57577 a_1203_42692.n3 a_1203_42692.t32 139.78
R57578 a_1203_42692.n4 a_1203_42692.t19 139.78
R57579 a_1203_42692.n30 a_1203_42692.n29 99.1759
R57580 a_1203_42692.n25 a_1203_42692.n0 91.5647
R57581 a_1203_42692.n29 a_1203_42692.n28 78.4622
R57582 a_1203_42692.n4 a_1203_42692.n3 61.346
R57583 a_1203_42692.n29 a_1203_42692.n25 46.0117
R57584 a_1203_42692.n25 a_1203_42692.n24 34.6867
R57585 a_1203_42692.n26 a_1203_42692.t6 26.5955
R57586 a_1203_42692.n26 a_1203_42692.t7 26.5955
R57587 a_1203_42692.n27 a_1203_42692.t4 26.5955
R57588 a_1203_42692.n27 a_1203_42692.t5 26.5955
R57589 a_1203_42692.n0 a_1203_42692.t2 24.9236
R57590 a_1203_42692.n0 a_1203_42692.t1 24.9236
R57591 a_1203_42692.n30 a_1203_42692.t0 24.9236
R57592 a_1203_42692.t3 a_1203_42692.n30 24.9236
R57593 a_1203_42692.n20 a_1203_42692.n18 21.2089
R57594 a_1203_42692.n14 a_1203_42692.n12 15.918
R57595 a_1203_42692.n12 a_1203_42692.n10 12.5636
R57596 a_1203_42692.n18 a_1203_42692.n16 12.417
R57597 a_1203_42692.n10 a_1203_42692.n9 11.4346
R57598 a_1203_42692.n7 a_1203_42692.n6 8.58978
R57599 a_1203_42692.n22 a_1203_42692.n20 8.28892
R57600 a_1203_42692.n24 a_1203_42692.n22 7.38649
R57601 a_1203_42692.n9 a_1203_42692.n7 4.86314
R57602 a_1203_42692.n16 a_1203_42692.n14 4.32038
R57603 a_14766_45596.n9 a_14766_45596.t1 366.548
R57604 a_14766_45596.t0 a_14766_45596.n9 307.562
R57605 a_14766_45596.n1 a_14766_45596.t9 293.969
R57606 a_14766_45596.n3 a_14766_45596.t2 241.536
R57607 a_14766_45596.n0 a_14766_45596.t8 231.017
R57608 a_14766_45596.n2 a_14766_45596.t3 222.018
R57609 a_14766_45596.n5 a_14766_45596.t6 186.03
R57610 a_14766_45596.n4 a_14766_45596.n3 182.418
R57611 a_14766_45596.n3 a_14766_45596.t5 169.237
R57612 a_14766_45596.n6 a_14766_45596.n5 168.034
R57613 a_14766_45596.n7 a_14766_45596.n1 164.066
R57614 a_14766_45596.n8 a_14766_45596.n0 162.952
R57615 a_14766_45596.n0 a_14766_45596.t11 158.716
R57616 a_14766_45596.n2 a_14766_45596.t7 140.064
R57617 a_14766_45596.n1 a_14766_45596.t4 138.338
R57618 a_14766_45596.n5 a_14766_45596.t10 137.829
R57619 a_14766_45596.n4 a_14766_45596.n2 91.5532
R57620 a_14766_45596.n9 a_14766_45596.n8 50.1195
R57621 a_14766_45596.n8 a_14766_45596.n7 13.0516
R57622 a_14766_45596.n7 a_14766_45596.n6 7.22577
R57623 a_14766_45596.n6 a_14766_45596.n4 4.57742
R57624 a_21020_30659.n1 a_21020_30659.t4 756.514
R57625 a_21020_30659.n1 a_21020_30659.t5 756.239
R57626 a_21020_30659.n2 a_21020_30659.n0 380.32
R57627 a_21020_30659.n3 a_21020_30659.n2 185
R57628 a_21020_30659.n2 a_21020_30659.n1 112.513
R57629 a_21020_30659.n0 a_21020_30659.t3 26.5955
R57630 a_21020_30659.n0 a_21020_30659.t2 26.5955
R57631 a_21020_30659.t1 a_21020_30659.n3 24.9236
R57632 a_21020_30659.n3 a_21020_30659.t0 24.9236
R57633 a_18314_32299.n9 a_18314_32299.t4 1415.15
R57634 a_18314_32299.n8 a_18314_32299.t6 1330.32
R57635 a_18314_32299.n6 a_18314_32299.t7 1330.32
R57636 a_18314_32299.n2 a_18314_32299.t9 1330.32
R57637 a_18314_32299.n3 a_18314_32299.t5 1320.68
R57638 a_18314_32299.n5 a_18314_32299.t8 1320.68
R57639 a_18314_32299.n7 a_18314_32299.t10 1320.68
R57640 a_18314_32299.n9 a_18314_32299.t11 1320.68
R57641 a_18314_32299.n11 a_18314_32299.n0 287.752
R57642 a_18314_32299.n12 a_18314_32299.n11 277.568
R57643 a_18314_32299.n4 a_18314_32299.n3 161.78
R57644 a_18314_32299.n5 a_18314_32299.n4 161.3
R57645 a_18314_32299.n7 a_18314_32299.n1 161.3
R57646 a_18314_32299.n10 a_18314_32299.n9 161.3
R57647 a_18314_32299.n11 a_18314_32299.n10 127.082
R57648 a_18314_32299.n9 a_18314_32299.n8 84.8325
R57649 a_18314_32299.n8 a_18314_32299.n7 84.8325
R57650 a_18314_32299.n7 a_18314_32299.n6 84.8325
R57651 a_18314_32299.n6 a_18314_32299.n5 84.8325
R57652 a_18314_32299.n5 a_18314_32299.n2 84.8325
R57653 a_18314_32299.n3 a_18314_32299.n2 84.8325
R57654 a_18314_32299.n0 a_18314_32299.t3 26.5955
R57655 a_18314_32299.n0 a_18314_32299.t2 26.5955
R57656 a_18314_32299.t1 a_18314_32299.n12 24.9236
R57657 a_18314_32299.n12 a_18314_32299.t0 24.9236
R57658 a_18314_32299.n4 a_18314_32299.n1 0.4805
R57659 a_18314_32299.n10 a_18314_32299.n1 0.4655
R57660 EN_VIN_BSTR_P.n20 EN_VIN_BSTR_P.t16 1559.46
R57661 EN_VIN_BSTR_P.n19 EN_VIN_BSTR_P.t9 1415.15
R57662 EN_VIN_BSTR_P.n19 EN_VIN_BSTR_P.t8 1320.68
R57663 EN_VIN_BSTR_P.n2 EN_VIN_BSTR_P.t19 748.122
R57664 EN_VIN_BSTR_P.n2 EN_VIN_BSTR_P.t7 678.014
R57665 EN_VIN_BSTR_P.n11 EN_VIN_BSTR_P.t12 605.802
R57666 EN_VIN_BSTR_P.n10 EN_VIN_BSTR_P.t15 444.502
R57667 EN_VIN_BSTR_P.n3 EN_VIN_BSTR_P.t18 398.575
R57668 EN_VIN_BSTR_P.n9 EN_VIN_BSTR_P.t17 382.812
R57669 EN_VIN_BSTR_P.n17 EN_VIN_BSTR_P.t21 381.798
R57670 EN_VIN_BSTR_P.n9 EN_VIN_BSTR_P.t23 381.793
R57671 EN_VIN_BSTR_P.n16 EN_VIN_BSTR_P.t10 381.788
R57672 EN_VIN_BSTR_P.n15 EN_VIN_BSTR_P.t22 381.413
R57673 EN_VIN_BSTR_P.n14 EN_VIN_BSTR_P.t14 381.413
R57674 EN_VIN_BSTR_P.n13 EN_VIN_BSTR_P.t20 381.413
R57675 EN_VIN_BSTR_P.n12 EN_VIN_BSTR_P.t11 381.413
R57676 EN_VIN_BSTR_P.n10 EN_VIN_BSTR_P.t13 356.68
R57677 EN_VIN_BSTR_P.n3 EN_VIN_BSTR_P.n2 176.421
R57678 EN_VIN_BSTR_P.n11 EN_VIN_BSTR_P.n10 161.768
R57679 EN_VIN_BSTR_P.n20 EN_VIN_BSTR_P.n19 161.3
R57680 EN_VIN_BSTR_P.n4 EN_VIN_BSTR_P.n1 56.3527
R57681 EN_VIN_BSTR_P.n5 EN_VIN_BSTR_P.n0 56.3527
R57682 EN_VIN_BSTR_P.n21 EN_VIN_BSTR_P.n18 28.2777
R57683 EN_VIN_BSTR_P.n6 EN_VIN_BSTR_P.t0 24.8256
R57684 EN_VIN_BSTR_P.n6 EN_VIN_BSTR_P.t2 24.1869
R57685 EN_VIN_BSTR_P.n7 EN_VIN_BSTR_P.t1 24.1612
R57686 EN_VIN_BSTR_P EN_VIN_BSTR_P.n21 22.3265
R57687 EN_VIN_BSTR_P EN_VIN_BSTR_P.n8 8.34025
R57688 EN_VIN_BSTR_P.n1 EN_VIN_BSTR_P.t5 8.12675
R57689 EN_VIN_BSTR_P.n1 EN_VIN_BSTR_P.t6 8.12675
R57690 EN_VIN_BSTR_P.n0 EN_VIN_BSTR_P.t4 8.12675
R57691 EN_VIN_BSTR_P.n0 EN_VIN_BSTR_P.t3 8.12675
R57692 EN_VIN_BSTR_P.n21 EN_VIN_BSTR_P.n20 4.51508
R57693 EN_VIN_BSTR_P.n4 EN_VIN_BSTR_P.n3 2.39112
R57694 EN_VIN_BSTR_P.n7 EN_VIN_BSTR_P.n6 0.989971
R57695 EN_VIN_BSTR_P.n17 EN_VIN_BSTR_P.n16 0.9005
R57696 EN_VIN_BSTR_P.n8 EN_VIN_BSTR_P.n5 0.888337
R57697 EN_VIN_BSTR_P.n18 EN_VIN_BSTR_P.n17 0.7005
R57698 EN_VIN_BSTR_P.n13 EN_VIN_BSTR_P.n12 0.512318
R57699 EN_VIN_BSTR_P.n14 EN_VIN_BSTR_P.n13 0.512318
R57700 EN_VIN_BSTR_P.n15 EN_VIN_BSTR_P.n14 0.512318
R57701 EN_VIN_BSTR_P.n5 EN_VIN_BSTR_P.n4 0.462038
R57702 EN_VIN_BSTR_P.n18 EN_VIN_BSTR_P.n9 0.3755
R57703 EN_VIN_BSTR_P.n12 EN_VIN_BSTR_P.n11 0.267318
R57704 EN_VIN_BSTR_P.n16 EN_VIN_BSTR_P.n15 0.138909
R57705 EN_VIN_BSTR_P.n8 EN_VIN_BSTR_P.n7 0.003
R57706 a_n2293_47044.n5 a_n2293_47044.n0 664.928
R57707 a_n2293_47044.n3 a_n2293_47044.t6 276.464
R57708 a_n2293_47044.n4 a_n2293_47044.n2 219.061
R57709 a_n2293_47044.n1 a_n2293_47044.t8 212.081
R57710 a_n2293_47044.n2 a_n2293_47044.t5 212.081
R57711 a_n2293_47044.n4 a_n2293_47044.n3 204.071
R57712 a_n2293_47044.n3 a_n2293_47044.t7 196.131
R57713 a_n2293_47044.n6 a_n2293_47044.n5 187.927
R57714 a_n2293_47044.n1 a_n2293_47044.t4 139.78
R57715 a_n2293_47044.n2 a_n2293_47044.t9 139.78
R57716 a_n2293_47044.n2 a_n2293_47044.n1 61.346
R57717 a_n2293_47044.n0 a_n2293_47044.t2 26.5955
R57718 a_n2293_47044.n0 a_n2293_47044.t3 26.5955
R57719 a_n2293_47044.t1 a_n2293_47044.n6 24.9236
R57720 a_n2293_47044.n6 a_n2293_47044.t0 24.9236
R57721 a_n2293_47044.n5 a_n2293_47044.n4 9.3005
R57722 a_n2103_45412.n4 a_n2103_45412.n3 335.238
R57723 a_n2103_45412.n10 a_n2103_45412.n9 300.118
R57724 a_n2103_45412.n6 a_n2103_45412.n5 299.834
R57725 a_n2103_45412.n8 a_n2103_45412.n7 299.834
R57726 a_n2103_45412.n9 a_n2103_45412.n0 291.81
R57727 a_n2103_45412.n1 a_n2103_45412.t9 276.464
R57728 a_n2103_45412.n3 a_n2103_45412.t8 212.081
R57729 a_n2103_45412.n2 a_n2103_45412.t13 212.081
R57730 a_n2103_45412.n4 a_n2103_45412.n1 196.959
R57731 a_n2103_45412.n1 a_n2103_45412.t11 196.131
R57732 a_n2103_45412.n3 a_n2103_45412.t12 139.78
R57733 a_n2103_45412.n2 a_n2103_45412.t10 139.78
R57734 a_n2103_45412.n9 a_n2103_45412.n8 79.8031
R57735 a_n2103_45412.n3 a_n2103_45412.n2 61.346
R57736 a_n2103_45412.n8 a_n2103_45412.n6 29.6732
R57737 a_n2103_45412.n7 a_n2103_45412.t5 26.5955
R57738 a_n2103_45412.n7 a_n2103_45412.t4 26.5955
R57739 a_n2103_45412.n5 a_n2103_45412.t6 26.5955
R57740 a_n2103_45412.n5 a_n2103_45412.t7 26.5955
R57741 a_n2103_45412.n10 a_n2103_45412.t0 26.5955
R57742 a_n2103_45412.t1 a_n2103_45412.n10 26.5955
R57743 a_n2103_45412.n0 a_n2103_45412.t2 24.9236
R57744 a_n2103_45412.n0 a_n2103_45412.t3 24.9236
R57745 a_n2103_45412.n6 a_n2103_45412.n4 10.2702
R57746 DEBUG_MUX[2].n0 DEBUG_MUX[2].t0 260.322
R57747 DEBUG_MUX[2].n0 DEBUG_MUX[2].t1 175.169
R57748 DEBUG_MUX[2] DEBUG_MUX[2].n0 169.506
R57749 a_n1732_35090.n3 a_n1732_35090.t11 749.612
R57750 a_n1732_35090.n9 a_n1732_35090.t14 748.122
R57751 a_n1732_35090.n7 a_n1732_35090.t8 748.122
R57752 a_n1732_35090.n3 a_n1732_35090.t13 684.441
R57753 a_n1732_35090.n5 a_n1732_35090.t9 684.441
R57754 a_n1732_35090.n4 a_n1732_35090.t10 684.441
R57755 a_n1732_35090.n9 a_n1732_35090.t15 678.014
R57756 a_n1732_35090.n7 a_n1732_35090.t12 678.014
R57757 a_n1732_35090.n13 a_n1732_35090.n12 244.069
R57758 a_n1732_35090.n2 a_n1732_35090.n0 236.589
R57759 a_n1732_35090.n14 a_n1732_35090.n13 204.892
R57760 a_n1732_35090.n2 a_n1732_35090.n1 200.321
R57761 a_n1732_35090.n8 a_n1732_35090.n7 163.538
R57762 a_n1732_35090.n10 a_n1732_35090.n9 163.538
R57763 a_n1732_35090.n6 a_n1732_35090.n5 161.512
R57764 a_n1732_35090.n6 a_n1732_35090.n3 161.488
R57765 a_n1732_35090.n4 a_n1732_35090.n3 65.1723
R57766 a_n1732_35090.n5 a_n1732_35090.n4 65.1723
R57767 a_n1732_35090.n11 a_n1732_35090.n2 26.8022
R57768 a_n1732_35090.n12 a_n1732_35090.t6 26.5955
R57769 a_n1732_35090.n12 a_n1732_35090.t1 26.5955
R57770 a_n1732_35090.n14 a_n1732_35090.t7 26.5955
R57771 a_n1732_35090.t0 a_n1732_35090.n14 26.5955
R57772 a_n1732_35090.n13 a_n1732_35090.n11 25.4552
R57773 a_n1732_35090.n0 a_n1732_35090.t2 24.9236
R57774 a_n1732_35090.n0 a_n1732_35090.t3 24.9236
R57775 a_n1732_35090.n1 a_n1732_35090.t4 24.9236
R57776 a_n1732_35090.n1 a_n1732_35090.t5 24.9236
R57777 a_n1732_35090.n8 a_n1732_35090.n6 7.9226
R57778 a_n1732_35090.n11 a_n1732_35090.n10 5.92878
R57779 a_n1732_35090.n10 a_n1732_35090.n8 2.47042
R57780 a_11455_44576.n18 a_11455_44576.t8 334.723
R57781 a_11455_44576.n10 a_11455_44576.t19 334.723
R57782 a_11455_44576.n9 a_11455_44576.t11 267.065
R57783 a_11455_44576.n8 a_11455_44576.t14 256.728
R57784 a_11455_44576.n2 a_11455_44576.n0 248.088
R57785 a_11455_44576.n7 a_11455_44576.t20 241.536
R57786 a_11455_44576.n11 a_11455_44576.t13 238.397
R57787 a_11455_44576.n3 a_11455_44576.t18 231.835
R57788 a_11455_44576.n4 a_11455_44576.t27 221.72
R57789 a_11455_44576.n5 a_11455_44576.t16 221.72
R57790 a_11455_44576.n2 a_11455_44576.n1 208.508
R57791 a_11455_44576.n18 a_11455_44576.t10 206.19
R57792 a_11455_44576.n10 a_11455_44576.t26 206.19
R57793 a_11455_44576.n20 a_11455_44576.n6 196.22
R57794 a_11455_44576.n11 a_11455_44576.t22 195.017
R57795 a_11455_44576.n12 a_11455_44576.n10 176.965
R57796 a_11455_44576.n12 a_11455_44576.n11 173.276
R57797 a_11455_44576.n17 a_11455_44576.n7 173.008
R57798 a_11455_44576.n7 a_11455_44576.t25 169.237
R57799 a_11455_44576.n13 a_11455_44576.n9 167.695
R57800 a_11455_44576.n15 a_11455_44576.n14 167.337
R57801 a_11455_44576.n21 a_11455_44576.n3 166.361
R57802 a_11455_44576.n16 a_11455_44576.n8 165.121
R57803 a_11455_44576.n19 a_11455_44576.n18 163.689
R57804 a_11455_44576.n8 a_11455_44576.t21 161.275
R57805 a_11455_44576.n3 a_11455_44576.t23 157.07
R57806 a_11455_44576.n4 a_11455_44576.t9 149.421
R57807 a_11455_44576.n5 a_11455_44576.t15 149.421
R57808 a_11455_44576.n9 a_11455_44576.t17 148.35
R57809 a_11455_44576.n25 a_11455_44576.n24 137.575
R57810 a_11455_44576.n14 a_11455_44576.t24 137.177
R57811 a_11455_44576.n14 a_11455_44576.t12 121.109
R57812 a_11455_44576.n24 a_11455_44576.n23 99.1749
R57813 a_11455_44576.n22 a_11455_44576.n2 38.4831
R57814 a_11455_44576.n6 a_11455_44576.n4 37.4894
R57815 a_11455_44576.n6 a_11455_44576.n5 37.4894
R57816 a_11455_44576.n0 a_11455_44576.t5 26.5955
R57817 a_11455_44576.n0 a_11455_44576.t6 26.5955
R57818 a_11455_44576.n1 a_11455_44576.t7 26.5955
R57819 a_11455_44576.n1 a_11455_44576.t4 26.5955
R57820 a_11455_44576.n23 a_11455_44576.t1 24.9236
R57821 a_11455_44576.n23 a_11455_44576.t2 24.9236
R57822 a_11455_44576.n25 a_11455_44576.t0 24.9236
R57823 a_11455_44576.t3 a_11455_44576.n25 24.9236
R57824 a_11455_44576.n24 a_11455_44576.n22 14.8665
R57825 a_11455_44576.n21 a_11455_44576.n20 13.1985
R57826 a_11455_44576.n15 a_11455_44576.n13 11.6063
R57827 a_11455_44576.n16 a_11455_44576.n15 9.52935
R57828 a_11455_44576.n22 a_11455_44576.n21 9.3005
R57829 a_11455_44576.n20 a_11455_44576.n19 5.20533
R57830 a_11455_44576.n19 a_11455_44576.n17 3.83532
R57831 a_11455_44576.n17 a_11455_44576.n16 1.98814
R57832 a_11455_44576.n13 a_11455_44576.n12 0.755995
R57833 a_3990_30651.n19 a_3990_30651.t20 1421.83
R57834 a_3990_30651.n9 a_3990_30651.t8 1421.83
R57835 a_3990_30651.n12 a_3990_30651.t12 1327.11
R57836 a_3990_30651.n16 a_3990_30651.t10 1327.11
R57837 a_3990_30651.n18 a_3990_30651.t15 1327.11
R57838 a_3990_30651.n8 a_3990_30651.t14 1327.11
R57839 a_3990_30651.n6 a_3990_30651.t19 1327.11
R57840 a_3990_30651.n2 a_3990_30651.t5 1327.11
R57841 a_3990_30651.n19 a_3990_30651.t9 1320.68
R57842 a_3990_30651.n17 a_3990_30651.t7 1320.68
R57843 a_3990_30651.n15 a_3990_30651.t18 1320.68
R57844 a_3990_30651.n13 a_3990_30651.t21 1320.68
R57845 a_3990_30651.n3 a_3990_30651.t4 1320.68
R57846 a_3990_30651.n5 a_3990_30651.t11 1320.68
R57847 a_3990_30651.n7 a_3990_30651.t16 1320.68
R57848 a_3990_30651.n9 a_3990_30651.t6 1320.68
R57849 a_3990_30651.n24 a_3990_30651.n0 296.139
R57850 a_3990_30651.n25 a_3990_30651.n24 269.182
R57851 a_3990_30651.n22 a_3990_30651.t13 260.322
R57852 a_3990_30651.n22 a_3990_30651.t17 175.169
R57853 a_3990_30651.n23 a_3990_30651.n22 174.507
R57854 a_3990_30651.n14 a_3990_30651.n13 161.701
R57855 a_3990_30651.n4 a_3990_30651.n3 161.701
R57856 a_3990_30651.n20 a_3990_30651.n19 161.3
R57857 a_3990_30651.n15 a_3990_30651.n14 161.3
R57858 a_3990_30651.n17 a_3990_30651.n11 161.3
R57859 a_3990_30651.n10 a_3990_30651.n9 161.3
R57860 a_3990_30651.n7 a_3990_30651.n1 161.3
R57861 a_3990_30651.n5 a_3990_30651.n4 161.3
R57862 a_3990_30651.n13 a_3990_30651.n12 94.7191
R57863 a_3990_30651.n15 a_3990_30651.n12 94.7191
R57864 a_3990_30651.n16 a_3990_30651.n15 94.7191
R57865 a_3990_30651.n17 a_3990_30651.n16 94.7191
R57866 a_3990_30651.n18 a_3990_30651.n17 94.7191
R57867 a_3990_30651.n19 a_3990_30651.n18 94.7191
R57868 a_3990_30651.n9 a_3990_30651.n8 94.7191
R57869 a_3990_30651.n8 a_3990_30651.n7 94.7191
R57870 a_3990_30651.n7 a_3990_30651.n6 94.7191
R57871 a_3990_30651.n6 a_3990_30651.n5 94.7191
R57872 a_3990_30651.n5 a_3990_30651.n2 94.7191
R57873 a_3990_30651.n3 a_3990_30651.n2 94.7191
R57874 a_3990_30651.n23 a_3990_30651.n21 81.2143
R57875 a_3990_30651.n21 a_3990_30651.n20 39.6536
R57876 a_3990_30651.n21 a_3990_30651.n10 36.1828
R57877 a_3990_30651.n0 a_3990_30651.t3 26.5955
R57878 a_3990_30651.n0 a_3990_30651.t2 26.5955
R57879 a_3990_30651.n25 a_3990_30651.t0 24.9236
R57880 a_3990_30651.t1 a_3990_30651.n25 24.9236
R57881 a_3990_30651.n24 a_3990_30651.n23 22.2526
R57882 a_3990_30651.n14 a_3990_30651.n11 0.4005
R57883 a_3990_30651.n20 a_3990_30651.n11 0.4005
R57884 a_3990_30651.n10 a_3990_30651.n1 0.4005
R57885 a_3990_30651.n4 a_3990_30651.n1 0.4005
R57886 a_1736_39043.n1 a_1736_39043.t5 440.13
R57887 a_1736_39043.t0 a_1736_39043.n4 239.113
R57888 a_1736_39043.n0 a_1736_39043.t3 230.576
R57889 a_1736_39043.n1 a_1736_39043.t4 192.331
R57890 a_1736_39043.n2 a_1736_39043.n0 169.999
R57891 a_1736_39043.n0 a_1736_39043.t6 158.275
R57892 a_1736_39043.n3 a_1736_39043.t1 85.6451
R57893 a_1736_39043.n4 a_1736_39043.t2 61.169
R57894 a_1736_39043.n3 a_1736_39043.n2 5.84425
R57895 a_1736_39043.n2 a_1736_39043.n1 4.5005
R57896 a_1736_39043.n4 a_1736_39043.n3 1.59495
R57897 a_135_43540.n2 a_135_43540.n1 647.148
R57898 a_135_43540.n5 a_135_43540.t20 408.63
R57899 a_135_43540.n13 a_135_43540.t25 408.63
R57900 a_135_43540.n9 a_135_43540.t45 408.63
R57901 a_135_43540.n19 a_135_43540.t13 408.63
R57902 a_135_43540.n22 a_135_43540.t34 408.63
R57903 a_135_43540.n25 a_135_43540.t35 408.63
R57904 a_135_43540.n28 a_135_43540.t32 408.63
R57905 a_135_43540.n16 a_135_43540.t8 408.63
R57906 a_135_43540.n35 a_135_43540.t14 408.63
R57907 a_135_43540.n6 a_135_43540.t11 408.63
R57908 a_135_43540.n41 a_135_43540.t29 347.577
R57909 a_135_43540.n12 a_135_43540.t39 347.577
R57910 a_135_43540.n10 a_135_43540.t28 347.577
R57911 a_135_43540.n20 a_135_43540.t41 347.577
R57912 a_135_43540.n23 a_135_43540.t10 347.577
R57913 a_135_43540.n26 a_135_43540.t46 347.577
R57914 a_135_43540.n29 a_135_43540.t23 347.577
R57915 a_135_43540.n17 a_135_43540.t19 347.577
R57916 a_135_43540.n36 a_135_43540.t15 347.577
R57917 a_135_43540.n7 a_135_43540.t31 347.577
R57918 a_135_43540.n4 a_135_43540.n3 243.627
R57919 a_135_43540.n2 a_135_43540.n0 194.441
R57920 a_135_43540.n41 a_135_43540.t26 193.337
R57921 a_135_43540.n12 a_135_43540.t9 193.337
R57922 a_135_43540.n10 a_135_43540.t40 193.337
R57923 a_135_43540.n20 a_135_43540.t17 193.337
R57924 a_135_43540.n23 a_135_43540.t44 193.337
R57925 a_135_43540.n26 a_135_43540.t38 193.337
R57926 a_135_43540.n29 a_135_43540.t30 193.337
R57927 a_135_43540.n17 a_135_43540.t37 193.337
R57928 a_135_43540.n36 a_135_43540.t22 193.337
R57929 a_135_43540.n7 a_135_43540.t18 193.337
R57930 a_135_43540.n45 a_135_43540.n44 185
R57931 a_135_43540.n11 a_135_43540.n9 167.666
R57932 a_135_43540.n21 a_135_43540.n19 167.666
R57933 a_135_43540.n27 a_135_43540.n25 167.666
R57934 a_135_43540.n8 a_135_43540.n6 167.666
R57935 a_135_43540.n30 a_135_43540.n28 167.663
R57936 a_135_43540.n37 a_135_43540.n35 167.663
R57937 a_135_43540.n18 a_135_43540.n16 167.601
R57938 a_135_43540.n43 a_135_43540.n5 167.567
R57939 a_135_43540.n14 a_135_43540.n13 165.524
R57940 a_135_43540.n24 a_135_43540.n22 165.072
R57941 a_135_43540.n24 a_135_43540.n23 163.006
R57942 a_135_43540.n14 a_135_43540.n12 162.424
R57943 a_135_43540.n18 a_135_43540.n17 160.476
R57944 a_135_43540.n42 a_135_43540.n41 160.415
R57945 a_135_43540.n11 a_135_43540.n10 160.415
R57946 a_135_43540.n21 a_135_43540.n20 160.415
R57947 a_135_43540.n27 a_135_43540.n26 160.415
R57948 a_135_43540.n8 a_135_43540.n7 160.415
R57949 a_135_43540.n30 a_135_43540.n29 160.415
R57950 a_135_43540.n37 a_135_43540.n36 160.415
R57951 a_135_43540.n5 a_135_43540.t12 132.282
R57952 a_135_43540.n13 a_135_43540.t33 132.282
R57953 a_135_43540.n9 a_135_43540.t21 132.282
R57954 a_135_43540.n19 a_135_43540.t24 132.282
R57955 a_135_43540.n22 a_135_43540.t36 132.282
R57956 a_135_43540.n25 a_135_43540.t16 132.282
R57957 a_135_43540.n28 a_135_43540.t42 132.282
R57958 a_135_43540.n16 a_135_43540.t43 132.282
R57959 a_135_43540.n35 a_135_43540.t27 132.282
R57960 a_135_43540.n6 a_135_43540.t47 132.282
R57961 a_135_43540.n4 a_135_43540.n2 50.5705
R57962 a_135_43540.n3 a_135_43540.t1 40.0005
R57963 a_135_43540.n3 a_135_43540.t2 40.0005
R57964 a_135_43540.n45 a_135_43540.t0 40.0005
R57965 a_135_43540.t3 a_135_43540.n45 40.0005
R57966 a_135_43540.n0 a_135_43540.t5 27.5805
R57967 a_135_43540.n0 a_135_43540.t7 27.5805
R57968 a_135_43540.n1 a_135_43540.t4 27.5805
R57969 a_135_43540.n1 a_135_43540.t6 27.5805
R57970 a_135_43540.n42 a_135_43540.n40 24.8474
R57971 a_135_43540.n44 a_135_43540.n43 20.0436
R57972 a_135_43540.n38 a_135_43540.n34 18.8287
R57973 a_135_43540.n44 a_135_43540.n4 15.262
R57974 a_135_43540.n33 a_135_43540.n32 14.8865
R57975 a_135_43540.n15 a_135_43540.n11 14.4351
R57976 a_135_43540.n31 a_135_43540.n27 13.2577
R57977 a_135_43540.n39 a_135_43540.n38 13.1245
R57978 a_135_43540.n33 a_135_43540.n21 9.33666
R57979 a_135_43540.n32 a_135_43540.n24 8.0068
R57980 a_135_43540.n40 a_135_43540.n39 6.49707
R57981 a_135_43540.n15 a_135_43540.n14 4.5005
R57982 a_135_43540.n34 a_135_43540.n33 4.5005
R57983 a_135_43540.n39 a_135_43540.n15 2.30064
R57984 a_135_43540.n32 a_135_43540.n31 0.572959
R57985 a_135_43540.n34 a_135_43540.n18 0.443874
R57986 a_135_43540.n43 a_135_43540.n42 0.0989262
R57987 a_135_43540.n31 a_135_43540.n30 0.0497651
R57988 a_135_43540.n40 a_135_43540.n8 0.0491212
R57989 a_135_43540.n38 a_135_43540.n37 0.0482664
R57990 a_134_42718.n2 a_134_42718.t5 586.74
R57991 a_134_42718.n2 a_134_42718.t6 586.269
R57992 a_134_42718.n4 a_134_42718.n0 380.32
R57993 a_134_42718.n1 a_134_42718.t7 260.322
R57994 a_134_42718.n5 a_134_42718.n4 185
R57995 a_134_42718.n1 a_134_42718.t4 175.169
R57996 a_134_42718.n3 a_134_42718.n1 173.109
R57997 a_134_42718.n3 a_134_42718.n2 130.141
R57998 a_134_42718.n0 a_134_42718.t2 26.5955
R57999 a_134_42718.n0 a_134_42718.t3 26.5955
R58000 a_134_42718.n5 a_134_42718.t0 24.9236
R58001 a_134_42718.t1 a_134_42718.n5 24.9236
R58002 a_134_42718.n4 a_134_42718.n3 21.2221
R58003 a_n2810_44350.n1 a_n2810_44350.t5 1415.15
R58004 a_n2810_44350.n1 a_n2810_44350.t4 1320.68
R58005 a_n2810_44350.n2 a_n2810_44350.n0 296.139
R58006 a_n2810_44350.n2 a_n2810_44350.n1 283.193
R58007 a_n2810_44350.n3 a_n2810_44350.n2 269.182
R58008 a_n2810_44350.n0 a_n2810_44350.t3 26.5955
R58009 a_n2810_44350.n0 a_n2810_44350.t2 26.5955
R58010 a_n2810_44350.t1 a_n2810_44350.n3 24.9236
R58011 a_n2810_44350.n3 a_n2810_44350.t0 24.9236
R58012 DATA[3].n3 DATA[3].n2 647.148
R58013 DATA[3].n5 DATA[3].n4 200.262
R58014 DATA[3].n3 DATA[3].n1 194.441
R58015 DATA[3].n6 DATA[3].n0 185
R58016 DATA[3].n6 DATA[3].n5 58.6278
R58017 DATA[3].n5 DATA[3].n3 50.5705
R58018 DATA[3].n0 DATA[3].t0 40.0005
R58019 DATA[3].n0 DATA[3].t3 40.0005
R58020 DATA[3].n4 DATA[3].t1 40.0005
R58021 DATA[3].n4 DATA[3].t2 40.0005
R58022 DATA[3].n1 DATA[3].t6 27.5805
R58023 DATA[3].n1 DATA[3].t5 27.5805
R58024 DATA[3].n2 DATA[3].t7 27.5805
R58025 DATA[3].n2 DATA[3].t4 27.5805
R58026 DATA[3] DATA[3].n6 18.089
R58027 C0_N_btm.n1 C0_N_btm.t0 101.944
R58028 C0_N_btm.n2 C0_N_btm.t1 99.4985
R58029 C0_N_btm.n0 C0_N_btm.t5 54.9098
R58030 C0_N_btm C0_N_btm.n2 49.2505
R58031 C0_N_btm.n0 C0_N_btm.t2 47.3635
R58032 C0_N_btm C0_N_btm.n3 8.68175
R58033 C0_N_btm.n1 C0_N_btm.n0 8.27654
R58034 C0_N_btm.n2 C0_N_btm.n1 6.33383
R58035 C0_N_btm.n3 C0_N_btm.t3 5.03712
R58036 C0_N_btm.n3 C0_N_btm.t4 4.03712
R58037 a_n2293_45420.n5 a_n2293_45420.n0 664.928
R58038 a_n2293_45420.n1 a_n2293_45420.t5 276.464
R58039 a_n2293_45420.n4 a_n2293_45420.n3 222.924
R58040 a_n2293_45420.n2 a_n2293_45420.t8 212.081
R58041 a_n2293_45420.n3 a_n2293_45420.t4 212.081
R58042 a_n2293_45420.n4 a_n2293_45420.n1 196.593
R58043 a_n2293_45420.n1 a_n2293_45420.t7 196.131
R58044 a_n2293_45420.n6 a_n2293_45420.n5 187.927
R58045 a_n2293_45420.n2 a_n2293_45420.t6 139.78
R58046 a_n2293_45420.n3 a_n2293_45420.t9 139.78
R58047 a_n2293_45420.n3 a_n2293_45420.n2 61.346
R58048 a_n2293_45420.n0 a_n2293_45420.t2 26.5955
R58049 a_n2293_45420.n0 a_n2293_45420.t3 26.5955
R58050 a_n2293_45420.n6 a_n2293_45420.t0 24.9236
R58051 a_n2293_45420.t1 a_n2293_45420.n6 24.9236
R58052 a_n2293_45420.n5 a_n2293_45420.n4 19.08
R58053 a_14297_32299.n1 a_14297_32299.t4 674.803
R58054 a_14297_32299.n1 a_14297_32299.n0 380.32
R58055 a_14297_32299.n2 a_14297_32299.n1 185
R58056 a_14297_32299.n0 a_14297_32299.t3 26.5955
R58057 a_14297_32299.n0 a_14297_32299.t2 26.5955
R58058 a_14297_32299.t1 a_14297_32299.n2 24.9236
R58059 a_14297_32299.n2 a_14297_32299.t0 24.9236
R58060 EN_COMP.n4 EN_COMP.n2 380.32
R58061 EN_COMP.n5 EN_COMP.n1 292.096
R58062 EN_COMP.n0 EN_COMP.t4 235.763
R58063 EN_COMP.n1 EN_COMP.t5 230.155
R58064 EN_COMP.n4 EN_COMP.n3 185
R58065 EN_COMP EN_COMP.n0 167.787
R58066 EN_COMP.n0 EN_COMP.t6 163.464
R58067 EN_COMP.n1 EN_COMP.t7 157.856
R58068 EN_COMP.n5 EN_COMP.n4 39.7555
R58069 EN_COMP EN_COMP.n5 29.8078
R58070 EN_COMP.n2 EN_COMP.t2 26.5955
R58071 EN_COMP.n2 EN_COMP.t3 26.5955
R58072 EN_COMP.n3 EN_COMP.t0 24.9236
R58073 EN_COMP.n3 EN_COMP.t1 24.9236
R58074 C5_P_btm.n1 C5_P_btm.t0 101.204
R58075 C5_P_btm.n2 C5_P_btm.t1 98.0923
R58076 C5_P_btm C5_P_btm.n2 57.563
R58077 C5_P_btm.n0 C5_P_btm.t37 54.9311
R58078 C5_P_btm.n0 C5_P_btm.t2 47.3635
R58079 C5_P_btm.n2 C5_P_btm.n1 8.08383
R58080 C5_P_btm C5_P_btm.n91 7.55675
R58081 C5_P_btm.n1 C5_P_btm.n0 6.87029
R58082 C5_P_btm.n55 C5_P_btm.t3 5.03712
R58083 C5_P_btm.n83 C5_P_btm.n82 4.60698
R58084 C5_P_btm.n84 C5_P_btm.n83 4.60698
R58085 C5_P_btm.n80 C5_P_btm.n79 4.60698
R58086 C5_P_btm.n81 C5_P_btm.n80 4.60698
R58087 C5_P_btm.n77 C5_P_btm.n76 4.60698
R58088 C5_P_btm.n78 C5_P_btm.n77 4.60698
R58089 C5_P_btm.n74 C5_P_btm.n73 4.60698
R58090 C5_P_btm.n75 C5_P_btm.n74 4.60698
R58091 C5_P_btm.n71 C5_P_btm.n70 4.60698
R58092 C5_P_btm.n72 C5_P_btm.n71 4.60698
R58093 C5_P_btm.n68 C5_P_btm.n67 4.60698
R58094 C5_P_btm.n69 C5_P_btm.n68 4.60698
R58095 C5_P_btm.n65 C5_P_btm.n64 4.60698
R58096 C5_P_btm.n66 C5_P_btm.n65 4.60698
R58097 C5_P_btm.n62 C5_P_btm.n61 4.60698
R58098 C5_P_btm.n63 C5_P_btm.n62 4.60698
R58099 C5_P_btm.n52 C5_P_btm.n51 4.60698
R58100 C5_P_btm.n53 C5_P_btm.n52 4.60698
R58101 C5_P_btm.n49 C5_P_btm.n48 4.60698
R58102 C5_P_btm.n50 C5_P_btm.n49 4.60698
R58103 C5_P_btm.n46 C5_P_btm.n45 4.60698
R58104 C5_P_btm.n47 C5_P_btm.n46 4.60698
R58105 C5_P_btm.n43 C5_P_btm.n42 4.60698
R58106 C5_P_btm.n44 C5_P_btm.n43 4.60698
R58107 C5_P_btm.n40 C5_P_btm.n39 4.60698
R58108 C5_P_btm.n41 C5_P_btm.n40 4.60698
R58109 C5_P_btm.n37 C5_P_btm.n36 4.60698
R58110 C5_P_btm.n38 C5_P_btm.n37 4.60698
R58111 C5_P_btm.n25 C5_P_btm.n24 4.60698
R58112 C5_P_btm.n24 C5_P_btm.n23 4.60698
R58113 C5_P_btm.n22 C5_P_btm.n21 4.60698
R58114 C5_P_btm.n21 C5_P_btm.n20 4.60698
R58115 C5_P_btm.n34 C5_P_btm.n33 4.60698
R58116 C5_P_btm.n35 C5_P_btm.n34 4.60698
R58117 C5_P_btm.n31 C5_P_btm.n30 4.60698
R58118 C5_P_btm.n32 C5_P_btm.n31 4.60698
R58119 C5_P_btm.n55 C5_P_btm.t16 4.03712
R58120 C5_P_btm.n56 C5_P_btm.t32 4.03712
R58121 C5_P_btm.n57 C5_P_btm.t28 4.03712
R58122 C5_P_btm.n58 C5_P_btm.t7 4.03712
R58123 C5_P_btm.n87 C5_P_btm.t10 4.03712
R58124 C5_P_btm.n88 C5_P_btm.t29 4.03712
R58125 C5_P_btm.n89 C5_P_btm.t33 4.03712
R58126 C5_P_btm.n90 C5_P_btm.t8 4.03712
R58127 C5_P_btm.n91 C5_P_btm.t4 4.03712
R58128 C5_P_btm.n85 C5_P_btm.t23 3.98193
R58129 C5_P_btm.n60 C5_P_btm.t22 3.98193
R58130 C5_P_btm.n54 C5_P_btm.t36 3.98193
R58131 C5_P_btm.n19 C5_P_btm.t12 3.98193
R58132 C5_P_btm.n26 C5_P_btm.t17 3.98193
R58133 C5_P_btm.n3 C5_P_btm.t19 3.98193
R58134 C5_P_btm.n83 C5_P_btm.t24 1.67819
R58135 C5_P_btm.n80 C5_P_btm.t21 1.67819
R58136 C5_P_btm.n77 C5_P_btm.t14 1.67819
R58137 C5_P_btm.n74 C5_P_btm.t34 1.67819
R58138 C5_P_btm.n71 C5_P_btm.t25 1.67819
R58139 C5_P_btm.n68 C5_P_btm.t31 1.67819
R58140 C5_P_btm.n65 C5_P_btm.t11 1.67819
R58141 C5_P_btm.n62 C5_P_btm.t6 1.67819
R58142 C5_P_btm.n52 C5_P_btm.t5 1.67819
R58143 C5_P_btm.n49 C5_P_btm.t20 1.67819
R58144 C5_P_btm.n46 C5_P_btm.t27 1.67819
R58145 C5_P_btm.n43 C5_P_btm.t26 1.67819
R58146 C5_P_btm.n40 C5_P_btm.t30 1.67819
R58147 C5_P_btm.n37 C5_P_btm.t9 1.67819
R58148 C5_P_btm.n24 C5_P_btm.t15 1.67819
R58149 C5_P_btm.n21 C5_P_btm.t18 1.67819
R58150 C5_P_btm.n34 C5_P_btm.t35 1.67819
R58151 C5_P_btm.n31 C5_P_btm.t13 1.67819
R58152 C5_P_btm.n19 C5_P_btm.n14 1.05569
R58153 C5_P_btm.n27 C5_P_btm.n26 1.05569
R58154 C5_P_btm.n86 C5_P_btm.n3 1.05569
R58155 C5_P_btm.n59 C5_P_btm.n54 1.05569
R58156 C5_P_btm.n56 C5_P_btm.n55 1.0005
R58157 C5_P_btm.n57 C5_P_btm.n56 1.0005
R58158 C5_P_btm.n58 C5_P_btm.n57 1.0005
R58159 C5_P_btm.n12 C5_P_btm.n11 1.0005
R58160 C5_P_btm.n13 C5_P_btm.n10 1.0005
R58161 C5_P_btm.n14 C5_P_btm.n9 1.0005
R58162 C5_P_btm.n15 C5_P_btm.n8 1.0005
R58163 C5_P_btm.n16 C5_P_btm.n7 1.0005
R58164 C5_P_btm.n17 C5_P_btm.n16 1.0005
R58165 C5_P_btm.n18 C5_P_btm.n15 1.0005
R58166 C5_P_btm.n27 C5_P_btm.n6 1.0005
R58167 C5_P_btm.n28 C5_P_btm.n5 1.0005
R58168 C5_P_btm.n29 C5_P_btm.n4 1.0005
R58169 C5_P_btm.n59 C5_P_btm.n58 1.0005
R58170 C5_P_btm.n87 C5_P_btm.n86 1.0005
R58171 C5_P_btm.n88 C5_P_btm.n87 1.0005
R58172 C5_P_btm.n89 C5_P_btm.n88 1.0005
R58173 C5_P_btm.n90 C5_P_btm.n89 1.0005
R58174 C5_P_btm.n91 C5_P_btm.n90 1.0005
R58175 C5_P_btm.n20 C5_P_btm.n19 0.679419
R58176 C5_P_btm.n26 C5_P_btm.n25 0.679419
R58177 C5_P_btm.n30 C5_P_btm.n3 0.679419
R58178 C5_P_btm.n54 C5_P_btm.n53 0.679419
R58179 C5_P_btm.n61 C5_P_btm.n60 0.679419
R58180 C5_P_btm.n85 C5_P_btm.n84 0.679419
R58181 C5_P_btm.n23 C5_P_btm.n22 0.6255
R58182 C5_P_btm.n33 C5_P_btm.n32 0.6255
R58183 C5_P_btm.n36 C5_P_btm.n35 0.6255
R58184 C5_P_btm.n39 C5_P_btm.n38 0.6255
R58185 C5_P_btm.n42 C5_P_btm.n41 0.6255
R58186 C5_P_btm.n45 C5_P_btm.n44 0.6255
R58187 C5_P_btm.n48 C5_P_btm.n47 0.6255
R58188 C5_P_btm.n51 C5_P_btm.n50 0.6255
R58189 C5_P_btm.n64 C5_P_btm.n63 0.6255
R58190 C5_P_btm.n67 C5_P_btm.n66 0.6255
R58191 C5_P_btm.n70 C5_P_btm.n69 0.6255
R58192 C5_P_btm.n73 C5_P_btm.n72 0.6255
R58193 C5_P_btm.n76 C5_P_btm.n75 0.6255
R58194 C5_P_btm.n79 C5_P_btm.n78 0.6255
R58195 C5_P_btm.n82 C5_P_btm.n81 0.6255
R58196 C5_P_btm.n20 C5_P_btm.n18 0.109875
R58197 C5_P_btm.n22 C5_P_btm.n18 0.109875
R58198 C5_P_btm.n23 C5_P_btm.n17 0.109875
R58199 C5_P_btm.n25 C5_P_btm.n17 0.109875
R58200 C5_P_btm.n32 C5_P_btm.n29 0.109875
R58201 C5_P_btm.n30 C5_P_btm.n29 0.109875
R58202 C5_P_btm.n35 C5_P_btm.n28 0.109875
R58203 C5_P_btm.n33 C5_P_btm.n28 0.109875
R58204 C5_P_btm.n38 C5_P_btm.n27 0.109875
R58205 C5_P_btm.n36 C5_P_btm.n27 0.109875
R58206 C5_P_btm.n41 C5_P_btm.n16 0.109875
R58207 C5_P_btm.n39 C5_P_btm.n16 0.109875
R58208 C5_P_btm.n44 C5_P_btm.n15 0.109875
R58209 C5_P_btm.n42 C5_P_btm.n15 0.109875
R58210 C5_P_btm.n47 C5_P_btm.n14 0.109875
R58211 C5_P_btm.n45 C5_P_btm.n14 0.109875
R58212 C5_P_btm.n50 C5_P_btm.n13 0.109875
R58213 C5_P_btm.n48 C5_P_btm.n13 0.109875
R58214 C5_P_btm.n53 C5_P_btm.n12 0.109875
R58215 C5_P_btm.n51 C5_P_btm.n12 0.109875
R58216 C5_P_btm.n61 C5_P_btm.n11 0.109875
R58217 C5_P_btm.n63 C5_P_btm.n11 0.109875
R58218 C5_P_btm.n64 C5_P_btm.n10 0.109875
R58219 C5_P_btm.n66 C5_P_btm.n10 0.109875
R58220 C5_P_btm.n67 C5_P_btm.n9 0.109875
R58221 C5_P_btm.n69 C5_P_btm.n9 0.109875
R58222 C5_P_btm.n70 C5_P_btm.n8 0.109875
R58223 C5_P_btm.n72 C5_P_btm.n8 0.109875
R58224 C5_P_btm.n73 C5_P_btm.n7 0.109875
R58225 C5_P_btm.n75 C5_P_btm.n7 0.109875
R58226 C5_P_btm.n76 C5_P_btm.n6 0.109875
R58227 C5_P_btm.n78 C5_P_btm.n6 0.109875
R58228 C5_P_btm.n79 C5_P_btm.n5 0.109875
R58229 C5_P_btm.n81 C5_P_btm.n5 0.109875
R58230 C5_P_btm.n82 C5_P_btm.n4 0.109875
R58231 C5_P_btm.n84 C5_P_btm.n4 0.109875
R58232 C5_P_btm.n60 C5_P_btm.n59 0.0556875
R58233 C5_P_btm.n86 C5_P_btm.n85 0.0556875
R58234 a_885_44868.n28 a_885_44868.n26 459.668
R58235 a_885_44868.n32 a_885_44868.n31 433.394
R58236 a_885_44868.n25 a_885_44868.n24 433.394
R58237 a_885_44868.n10 a_885_44868.n9 433.394
R58238 a_885_44868.n16 a_885_44868.n14 433.394
R58239 a_885_44868.n13 a_885_44868.n12 433.394
R58240 a_885_44868.n30 a_885_44868.t31 329.902
R58241 a_885_44868.n23 a_885_44868.t21 329.902
R58242 a_885_44868.n27 a_885_44868.t26 329.902
R58243 a_885_44868.n8 a_885_44868.t28 329.902
R58244 a_885_44868.n15 a_885_44868.t36 329.902
R58245 a_885_44868.n11 a_885_44868.t15 329.902
R58246 a_885_44868.n31 a_885_44868.t30 272.062
R58247 a_885_44868.n24 a_885_44868.t23 272.062
R58248 a_885_44868.n26 a_885_44868.t13 272.062
R58249 a_885_44868.n9 a_885_44868.t17 272.062
R58250 a_885_44868.n14 a_885_44868.t14 272.062
R58251 a_885_44868.n12 a_885_44868.t33 272.062
R58252 a_885_44868.n5 a_885_44868.n4 256.103
R58253 a_885_44868.n2 a_885_44868.n0 241.847
R58254 a_885_44868.n17 a_885_44868.t35 241.536
R58255 a_885_44868.n31 a_885_44868.t27 206.19
R58256 a_885_44868.n24 a_885_44868.t39 206.19
R58257 a_885_44868.n26 a_885_44868.t32 206.19
R58258 a_885_44868.n21 a_885_44868.t18 206.19
R58259 a_885_44868.n9 a_885_44868.t20 206.19
R58260 a_885_44868.n14 a_885_44868.t12 206.19
R58261 a_885_44868.n12 a_885_44868.t38 206.19
R58262 a_885_44868.n37 a_885_44868.n36 205.28
R58263 a_885_44868.n5 a_885_44868.n3 202.095
R58264 a_885_44868.n35 a_885_44868.n7 190.911
R58265 a_885_44868.n2 a_885_44868.n1 185
R58266 a_885_44868.n32 a_885_44868.n30 178.274
R58267 a_885_44868.n25 a_885_44868.n23 178.274
R58268 a_885_44868.n10 a_885_44868.n8 178.274
R58269 a_885_44868.n16 a_885_44868.n15 178.274
R58270 a_885_44868.n13 a_885_44868.n11 178.274
R58271 a_885_44868.n22 a_885_44868.n21 169.674
R58272 a_885_44868.n17 a_885_44868.t24 169.237
R58273 a_885_44868.n18 a_885_44868.n17 167.368
R58274 a_885_44868.n28 a_885_44868.n27 152
R58275 a_885_44868.n30 a_885_44868.t19 148.35
R58276 a_885_44868.n23 a_885_44868.t29 148.35
R58277 a_885_44868.n27 a_885_44868.t16 148.35
R58278 a_885_44868.n8 a_885_44868.t34 148.35
R58279 a_885_44868.n15 a_885_44868.t25 148.35
R58280 a_885_44868.n11 a_885_44868.t22 148.35
R58281 a_885_44868.n21 a_885_44868.t37 142.344
R58282 a_885_44868.n36 a_885_44868.n35 52.7703
R58283 a_885_44868.n36 a_885_44868.n6 37.2711
R58284 a_885_44868.n6 a_885_44868.n2 28.2251
R58285 a_885_44868.n7 a_885_44868.t1 26.5955
R58286 a_885_44868.n7 a_885_44868.t2 26.5955
R58287 a_885_44868.n3 a_885_44868.t9 26.5955
R58288 a_885_44868.n3 a_885_44868.t11 26.5955
R58289 a_885_44868.n4 a_885_44868.t8 26.5955
R58290 a_885_44868.n4 a_885_44868.t10 26.5955
R58291 a_885_44868.n37 a_885_44868.t0 26.5955
R58292 a_885_44868.t3 a_885_44868.n37 26.5955
R58293 a_885_44868.n1 a_885_44868.t7 24.9236
R58294 a_885_44868.n1 a_885_44868.t5 24.9236
R58295 a_885_44868.n0 a_885_44868.t6 24.9236
R58296 a_885_44868.n0 a_885_44868.t4 24.9236
R58297 a_885_44868.n18 a_885_44868.n16 23.8283
R58298 a_885_44868.n29 a_885_44868.n25 22.7306
R58299 a_885_44868.n29 a_885_44868.n28 21.9529
R58300 a_885_44868.n35 a_885_44868.n34 19.2755
R58301 a_885_44868.n34 a_885_44868.n22 15.576
R58302 a_885_44868.n6 a_885_44868.n5 13.5534
R58303 a_885_44868.n34 a_885_44868.n33 13.1186
R58304 a_885_44868.n19 a_885_44868.n13 12.0589
R58305 a_885_44868.n22 a_885_44868.n20 11.2268
R58306 a_885_44868.n33 a_885_44868.n29 10.1901
R58307 a_885_44868.n33 a_885_44868.n32 9.3005
R58308 a_885_44868.n20 a_885_44868.n10 9.3005
R58309 a_885_44868.n19 a_885_44868.n18 8.9222
R58310 a_885_44868.n20 a_885_44868.n19 1.52676
R58311 a_12651_44576.n9 a_12651_44576.t25 334.723
R58312 a_12651_44576.n12 a_12651_44576.t8 323.342
R58313 a_12651_44576.n8 a_12651_44576.t18 267.065
R58314 a_12651_44576.n13 a_12651_44576.t14 256.728
R58315 a_12651_44576.n2 a_12651_44576.n0 248.088
R58316 a_12651_44576.n7 a_12651_44576.t12 241.536
R58317 a_12651_44576.n6 a_12651_44576.t23 238.397
R58318 a_12651_44576.n20 a_12651_44576.t15 231.835
R58319 a_12651_44576.n3 a_12651_44576.t21 221.72
R58320 a_12651_44576.n4 a_12651_44576.t16 221.72
R58321 a_12651_44576.n2 a_12651_44576.n1 208.508
R58322 a_12651_44576.n9 a_12651_44576.t10 206.19
R58323 a_12651_44576.n6 a_12651_44576.t24 195.017
R58324 a_12651_44576.n12 a_12651_44576.t22 194.809
R58325 a_12651_44576.n16 a_12651_44576.n8 191.333
R58326 a_12651_44576.n19 a_12651_44576.n5 191.22
R58327 a_12651_44576.n14 a_12651_44576.n12 179.601
R58328 a_12651_44576.n18 a_12651_44576.n6 174.286
R58329 a_12651_44576.n17 a_12651_44576.n7 174.073
R58330 a_12651_44576.n21 a_12651_44576.n20 173.446
R58331 a_12651_44576.n7 a_12651_44576.t19 169.237
R58332 a_12651_44576.n11 a_12651_44576.n9 168.62
R58333 a_12651_44576.n11 a_12651_44576.n10 162.837
R58334 a_12651_44576.n14 a_12651_44576.n13 162.464
R58335 a_12651_44576.n13 a_12651_44576.t27 161.275
R58336 a_12651_44576.n20 a_12651_44576.t20 157.07
R58337 a_12651_44576.n3 a_12651_44576.t26 149.421
R58338 a_12651_44576.n4 a_12651_44576.t11 149.421
R58339 a_12651_44576.n8 a_12651_44576.t9 148.35
R58340 a_12651_44576.n25 a_12651_44576.n24 137.575
R58341 a_12651_44576.n10 a_12651_44576.t17 137.177
R58342 a_12651_44576.n10 a_12651_44576.t13 121.109
R58343 a_12651_44576.n24 a_12651_44576.n23 99.1749
R58344 a_12651_44576.n22 a_12651_44576.n2 38.4831
R58345 a_12651_44576.n5 a_12651_44576.n3 37.4894
R58346 a_12651_44576.n5 a_12651_44576.n4 37.4894
R58347 a_12651_44576.n0 a_12651_44576.t7 26.5955
R58348 a_12651_44576.n0 a_12651_44576.t5 26.5955
R58349 a_12651_44576.n1 a_12651_44576.t6 26.5955
R58350 a_12651_44576.n1 a_12651_44576.t4 26.5955
R58351 a_12651_44576.n23 a_12651_44576.t2 24.9236
R58352 a_12651_44576.n23 a_12651_44576.t1 24.9236
R58353 a_12651_44576.t3 a_12651_44576.n25 24.9236
R58354 a_12651_44576.n25 a_12651_44576.t0 24.9236
R58355 a_12651_44576.n16 a_12651_44576.n15 23.1942
R58356 a_12651_44576.n15 a_12651_44576.n11 15.1985
R58357 a_12651_44576.n22 a_12651_44576.n21 14.916
R58358 a_12651_44576.n24 a_12651_44576.n22 14.8665
R58359 a_12651_44576.n17 a_12651_44576.n16 8.72028
R58360 a_12651_44576.n19 a_12651_44576.n18 6.61314
R58361 a_12651_44576.n15 a_12651_44576.n14 4.5005
R58362 a_12651_44576.n21 a_12651_44576.n19 3.51149
R58363 a_12651_44576.n18 a_12651_44576.n17 1.98814
R58364 a_n2810_43806.n1 a_n2810_43806.t4 444.502
R58365 a_n2810_43806.n1 a_n2810_43806.t5 356.68
R58366 a_n2810_43806.n2 a_n2810_43806.n1 296.587
R58367 a_n2810_43806.n2 a_n2810_43806.n0 296.139
R58368 a_n2810_43806.n3 a_n2810_43806.n2 269.182
R58369 a_n2810_43806.n0 a_n2810_43806.t3 26.5955
R58370 a_n2810_43806.n0 a_n2810_43806.t2 26.5955
R58371 a_n2810_43806.n3 a_n2810_43806.t0 24.9236
R58372 a_n2810_43806.t1 a_n2810_43806.n3 24.9236
R58373 a_n2103_44868.n9 a_n2103_44868.n8 300.118
R58374 a_n2103_44868.n5 a_n2103_44868.n4 299.834
R58375 a_n2103_44868.n7 a_n2103_44868.n6 299.834
R58376 a_n2103_44868.n10 a_n2103_44868.n9 291.81
R58377 a_n2103_44868.n0 a_n2103_44868.t12 276.464
R58378 a_n2103_44868.n3 a_n2103_44868.n2 228.173
R58379 a_n2103_44868.n2 a_n2103_44868.t10 212.081
R58380 a_n2103_44868.n1 a_n2103_44868.t13 212.081
R58381 a_n2103_44868.n3 a_n2103_44868.n0 208.881
R58382 a_n2103_44868.n0 a_n2103_44868.t9 196.131
R58383 a_n2103_44868.n2 a_n2103_44868.t11 139.78
R58384 a_n2103_44868.n1 a_n2103_44868.t8 139.78
R58385 a_n2103_44868.n9 a_n2103_44868.n7 79.8031
R58386 a_n2103_44868.n2 a_n2103_44868.n1 61.346
R58387 a_n2103_44868.n7 a_n2103_44868.n5 29.6732
R58388 a_n2103_44868.n8 a_n2103_44868.t2 26.5955
R58389 a_n2103_44868.n8 a_n2103_44868.t3 26.5955
R58390 a_n2103_44868.n6 a_n2103_44868.t6 26.5955
R58391 a_n2103_44868.n6 a_n2103_44868.t7 26.5955
R58392 a_n2103_44868.n4 a_n2103_44868.t4 26.5955
R58393 a_n2103_44868.n4 a_n2103_44868.t5 26.5955
R58394 a_n2103_44868.n10 a_n2103_44868.t0 24.9236
R58395 a_n2103_44868.t1 a_n2103_44868.n10 24.9236
R58396 a_n2103_44868.n5 a_n2103_44868.n3 10.2702
R58397 a_5840_42718.n2 a_5840_42718.t4 581.59
R58398 a_5840_42718.n2 a_5840_42718.t6 579.811
R58399 a_5840_42718.n4 a_5840_42718.n0 380.32
R58400 a_5840_42718.n1 a_5840_42718.t5 260.322
R58401 a_5840_42718.n5 a_5840_42718.n4 185
R58402 a_5840_42718.n1 a_5840_42718.t7 175.169
R58403 a_5840_42718.n3 a_5840_42718.n1 170.444
R58404 a_5840_42718.n3 a_5840_42718.n2 116.037
R58405 a_5840_42718.n0 a_5840_42718.t2 26.5955
R58406 a_5840_42718.n0 a_5840_42718.t3 26.5955
R58407 a_5840_42718.n5 a_5840_42718.t0 24.9236
R58408 a_5840_42718.t1 a_5840_42718.n5 24.9236
R58409 a_5840_42718.n4 a_5840_42718.n3 21.5639
R58410 a_15549_47044.n5 a_15549_47044.t10 241.536
R58411 a_15549_47044.n0 a_15549_47044.t11 231.017
R58412 a_15549_47044.n6 a_15549_47044.t3 229.184
R58413 a_15549_47044.n9 a_15549_47044.t1 217.506
R58414 a_15549_47044.n4 a_15549_47044.n3 216.15
R58415 a_15549_47044.n1 a_15549_47044.t5 212.081
R58416 a_15549_47044.n2 a_15549_47044.t9 212.081
R58417 a_15549_47044.n10 a_15549_47044.n9 181.583
R58418 a_15549_47044.n7 a_15549_47044.n6 181.071
R58419 a_15549_47044.n4 a_15549_47044.n0 174.13
R58420 a_15549_47044.n7 a_15549_47044.n5 169.44
R58421 a_15549_47044.n5 a_15549_47044.t6 169.237
R58422 a_15549_47044.n0 a_15549_47044.t8 158.716
R58423 a_15549_47044.n6 a_15549_47044.t4 156.883
R58424 a_15549_47044.n1 a_15549_47044.t12 139.78
R58425 a_15549_47044.n2 a_15549_47044.t7 139.78
R58426 a_15549_47044.n8 a_15549_47044.n7 31.8605
R58427 a_15549_47044.n3 a_15549_47044.n1 31.4035
R58428 a_15549_47044.n3 a_15549_47044.n2 31.4035
R58429 a_15549_47044.t0 a_15549_47044.n10 24.9236
R58430 a_15549_47044.n10 a_15549_47044.t2 24.9236
R58431 a_15549_47044.n9 a_15549_47044.n8 18.9814
R58432 a_15549_47044.n8 a_15549_47044.n4 7.37154
R58433 a_n2293_45956.n5 a_n2293_45956.n0 664.928
R58434 a_n2293_45956.n3 a_n2293_45956.t6 276.464
R58435 a_n2293_45956.n4 a_n2293_45956.n2 236.279
R58436 a_n2293_45956.n4 a_n2293_45956.n3 215.228
R58437 a_n2293_45956.n1 a_n2293_45956.t7 212.081
R58438 a_n2293_45956.n2 a_n2293_45956.t5 212.081
R58439 a_n2293_45956.n3 a_n2293_45956.t4 196.131
R58440 a_n2293_45956.n6 a_n2293_45956.n5 187.927
R58441 a_n2293_45956.n1 a_n2293_45956.t9 139.78
R58442 a_n2293_45956.n2 a_n2293_45956.t8 139.78
R58443 a_n2293_45956.n2 a_n2293_45956.n1 61.346
R58444 a_n2293_45956.n0 a_n2293_45956.t3 26.5955
R58445 a_n2293_45956.n0 a_n2293_45956.t2 26.5955
R58446 a_n2293_45956.t1 a_n2293_45956.n6 24.9236
R58447 a_n2293_45956.n6 a_n2293_45956.t0 24.9236
R58448 a_n2293_45956.n5 a_n2293_45956.n4 9.3005
R58449 a_14601_32299.n1 a_14601_32299.t5 444.502
R58450 a_14601_32299.n1 a_14601_32299.t4 356.68
R58451 a_14601_32299.n2 a_14601_32299.n1 303.603
R58452 a_14601_32299.n2 a_14601_32299.n0 287.752
R58453 a_14601_32299.n3 a_14601_32299.n2 277.568
R58454 a_14601_32299.n0 a_14601_32299.t2 26.5955
R58455 a_14601_32299.n0 a_14601_32299.t3 26.5955
R58456 a_14601_32299.n3 a_14601_32299.t0 24.9236
R58457 a_14601_32299.t1 a_14601_32299.n3 24.9236
R58458 C4_N_btm.n1 C4_N_btm.t0 101.361
R58459 C4_N_btm.n2 C4_N_btm.t2 98.3735
R58460 C4_N_btm.n0 C4_N_btm.t1 54.9311
R58461 C4_N_btm C4_N_btm.n2 54.563
R58462 C4_N_btm.n0 C4_N_btm.t3 47.3635
R58463 C4_N_btm.n2 C4_N_btm.n1 8.08383
R58464 C4_N_btm C4_N_btm.n22 7.74425
R58465 C4_N_btm.n1 C4_N_btm.n0 7.15154
R58466 C4_N_btm.n4 C4_N_btm.t22 5.03712
R58467 C4_N_btm.n18 C4_N_btm.t20 5.03712
R58468 C4_N_btm.n4 C4_N_btm.t10 4.03712
R58469 C4_N_btm.n5 C4_N_btm.t5 4.03712
R58470 C4_N_btm.n6 C4_N_btm.t14 4.03712
R58471 C4_N_btm.n15 C4_N_btm.t13 4.03712
R58472 C4_N_btm.n22 C4_N_btm.t21 4.03712
R58473 C4_N_btm.n20 C4_N_btm.t6 3.98193
R58474 C4_N_btm.n14 C4_N_btm.t15 3.98193
R58475 C4_N_btm.n7 C4_N_btm.t17 3.98193
R58476 C4_N_btm.n3 C4_N_btm.t9 3.98193
R58477 C4_N_btm.n16 C4_N_btm.t12 3.98193
R58478 C4_N_btm.n19 C4_N_btm.t16 3.98193
R58479 C4_N_btm.n13 C4_N_btm.t4 3.92851
R58480 C4_N_btm.n12 C4_N_btm.t8 3.92851
R58481 C4_N_btm.n11 C4_N_btm.t19 3.92851
R58482 C4_N_btm.n10 C4_N_btm.t7 3.92851
R58483 C4_N_btm.n9 C4_N_btm.t18 3.92851
R58484 C4_N_btm.n8 C4_N_btm.t11 3.92851
R58485 C4_N_btm.n7 C4_N_btm.n6 1.05569
R58486 C4_N_btm.n15 C4_N_btm.n14 1.05569
R58487 C4_N_btm.n21 C4_N_btm.n3 1.05569
R58488 C4_N_btm.n5 C4_N_btm.n4 1.0005
R58489 C4_N_btm.n6 C4_N_btm.n5 1.0005
R58490 C4_N_btm.n17 C4_N_btm.n15 1.0005
R58491 C4_N_btm.n18 C4_N_btm.n17 1.0005
R58492 C4_N_btm.n22 C4_N_btm.n21 1.0005
R58493 C4_N_btm.n9 C4_N_btm.n8 0.840176
R58494 C4_N_btm.n10 C4_N_btm.n9 0.840176
R58495 C4_N_btm.n11 C4_N_btm.n10 0.840176
R58496 C4_N_btm.n12 C4_N_btm.n11 0.840176
R58497 C4_N_btm.n13 C4_N_btm.n12 0.840176
R58498 C4_N_btm.n8 C4_N_btm.n7 0.786757
R58499 C4_N_btm.n14 C4_N_btm.n13 0.786757
R58500 C4_N_btm.n16 C4_N_btm.n3 0.733338
R58501 C4_N_btm.n20 C4_N_btm.n19 0.733338
R58502 C4_N_btm.n17 C4_N_btm.n16 0.0556875
R58503 C4_N_btm.n19 C4_N_btm.n18 0.0556875
R58504 C4_N_btm.n21 C4_N_btm.n20 0.0556875
R58505 a_21276_30659.n1 a_21276_30659.t7 756.547
R58506 a_21276_30659.n3 a_21276_30659.t5 756.226
R58507 a_21276_30659.n1 a_21276_30659.t6 756.226
R58508 a_21276_30659.n2 a_21276_30659.t4 756.226
R58509 a_21276_30659.n4 a_21276_30659.n0 287.752
R58510 a_21276_30659.n5 a_21276_30659.n4 277.568
R58511 a_21276_30659.n4 a_21276_30659.n3 119.04
R58512 a_21276_30659.n0 a_21276_30659.t3 26.5955
R58513 a_21276_30659.n0 a_21276_30659.t2 26.5955
R58514 a_21276_30659.n5 a_21276_30659.t0 24.9236
R58515 a_21276_30659.t1 a_21276_30659.n5 24.9236
R58516 a_21276_30659.n2 a_21276_30659.n1 0.3205
R58517 a_21276_30659.n3 a_21276_30659.n2 0.304667
R58518 a_n2442_44350.n1 a_n2442_44350.t4 1692.18
R58519 a_n2442_44350.n1 a_n2442_44350.n0 287.752
R58520 a_n2442_44350.n2 a_n2442_44350.n1 277.568
R58521 a_n2442_44350.n0 a_n2442_44350.t2 26.5955
R58522 a_n2442_44350.n0 a_n2442_44350.t3 26.5955
R58523 a_n2442_44350.n2 a_n2442_44350.t0 24.9236
R58524 a_n2442_44350.t1 a_n2442_44350.n2 24.9236
R58525 C1_N_btm.n2 C1_N_btm.t0 102.406
R58526 C1_N_btm.n1 C1_N_btm.t5 101.787
R58527 C1_N_btm.n0 C1_N_btm.t4 54.9098
R58528 C1_N_btm C1_N_btm.n2 47.6567
R58529 C1_N_btm.n0 C1_N_btm.t6 47.3635
R58530 C1_N_btm C1_N_btm.n4 8.93175
R58531 C1_N_btm.n2 C1_N_btm.n1 8.33383
R58532 C1_N_btm.n1 C1_N_btm.n0 7.99529
R58533 C1_N_btm.n3 C1_N_btm.t2 5.03712
R58534 C1_N_btm.n3 C1_N_btm.t1 4.03712
R58535 C1_N_btm.n4 C1_N_btm.t3 4.03712
R58536 C1_N_btm.n4 C1_N_btm.n3 1.0005
R58537 a_13667_32299.n1 a_13667_32299.t4 676.463
R58538 a_13667_32299.n1 a_13667_32299.n0 380.32
R58539 a_13667_32299.n2 a_13667_32299.n1 185
R58540 a_13667_32299.n0 a_13667_32299.t2 26.5955
R58541 a_13667_32299.n0 a_13667_32299.t3 26.5955
R58542 a_13667_32299.t1 a_13667_32299.n2 24.9236
R58543 a_13667_32299.n2 a_13667_32299.t0 24.9236
R58544 a_7557_43236.n4 a_7557_43236.t12 330.12
R58545 a_7557_43236.n3 a_7557_43236.t23 310.457
R58546 a_7557_43236.n12 a_7557_43236.t8 267.065
R58547 a_7557_43236.n8 a_7557_43236.t9 256.726
R58548 a_7557_43236.n2 a_7557_43236.n0 248.088
R58549 a_7557_43236.n7 a_7557_43236.t25 241.536
R58550 a_7557_43236.n14 a_7557_43236.t20 238.397
R58551 a_7557_43236.n6 a_7557_43236.t15 231.835
R58552 a_7557_43236.n16 a_7557_43236.t16 221.72
R58553 a_7557_43236.n17 a_7557_43236.t10 221.72
R58554 a_7557_43236.n3 a_7557_43236.t11 220.484
R58555 a_7557_43236.n2 a_7557_43236.n1 208.508
R58556 a_7557_43236.n4 a_7557_43236.t18 201.587
R58557 a_7557_43236.n9 a_7557_43236.n8 200.221
R58558 a_7557_43236.n5 a_7557_43236.n4 197.452
R58559 a_7557_43236.n14 a_7557_43236.t24 195.017
R58560 a_7557_43236.n13 a_7557_43236.n12 185.349
R58561 a_7557_43236.n13 a_7557_43236.n11 182.62
R58562 a_7557_43236.n15 a_7557_43236.n14 179.73
R58563 a_7557_43236.n5 a_7557_43236.n3 178.505
R58564 a_7557_43236.n9 a_7557_43236.n7 173.312
R58565 a_7557_43236.n7 a_7557_43236.t26 169.237
R58566 a_7557_43236.n10 a_7557_43236.n6 168.323
R58567 a_7557_43236.n19 a_7557_43236.n18 166.101
R58568 a_7557_43236.n8 a_7557_43236.t14 161.275
R58569 a_7557_43236.n6 a_7557_43236.t17 157.07
R58570 a_7557_43236.n16 a_7557_43236.t21 149.421
R58571 a_7557_43236.n17 a_7557_43236.t27 149.421
R58572 a_7557_43236.n12 a_7557_43236.t22 148.35
R58573 a_7557_43236.n25 a_7557_43236.n24 137.575
R58574 a_7557_43236.n11 a_7557_43236.t19 137.177
R58575 a_7557_43236.n11 a_7557_43236.t13 121.109
R58576 a_7557_43236.n24 a_7557_43236.n23 99.1749
R58577 a_7557_43236.n18 a_7557_43236.n16 37.4894
R58578 a_7557_43236.n18 a_7557_43236.n17 37.4894
R58579 a_7557_43236.n24 a_7557_43236.n22 36.0958
R58580 a_7557_43236.n0 a_7557_43236.t5 26.5955
R58581 a_7557_43236.n0 a_7557_43236.t7 26.5955
R58582 a_7557_43236.n1 a_7557_43236.t6 26.5955
R58583 a_7557_43236.n1 a_7557_43236.t4 26.5955
R58584 a_7557_43236.n23 a_7557_43236.t1 24.9236
R58585 a_7557_43236.n23 a_7557_43236.t0 24.9236
R58586 a_7557_43236.t3 a_7557_43236.n25 24.9236
R58587 a_7557_43236.n25 a_7557_43236.t2 24.9236
R58588 a_7557_43236.n21 a_7557_43236.n5 17.4128
R58589 a_7557_43236.n22 a_7557_43236.n2 17.2539
R58590 a_7557_43236.n21 a_7557_43236.n20 10.1339
R58591 a_7557_43236.n22 a_7557_43236.n21 9.3005
R58592 a_7557_43236.n19 a_7557_43236.n15 8.65705
R58593 a_7557_43236.n10 a_7557_43236.n9 8.13099
R58594 a_7557_43236.n15 a_7557_43236.n13 7.8509
R58595 a_7557_43236.n20 a_7557_43236.n19 6.7972
R58596 a_7557_43236.n20 a_7557_43236.n10 1.98814
R58597 a_7029_44350.n2 a_7029_44350.t1 275.784
R58598 a_7029_44350.t0 a_7029_44350.n1 272.971
R58599 a_7029_44350.t0 a_7029_44350.n2 258.846
R58600 a_7029_44350.n0 a_7029_44350.t3 241.536
R58601 a_7029_44350.n1 a_7029_44350.n0 215.407
R58602 a_7029_44350.n0 a_7029_44350.t2 169.237
R58603 a_7029_44350.n2 a_7029_44350.n1 7.90638
R58604 RST_Z.n0 RST_Z.t3 751.299
R58605 RST_Z.n0 RST_Z.t5 403.308
R58606 RST_Z.n3 RST_Z.t0 260.322
R58607 RST_Z.n1 RST_Z.t1 230.576
R58608 RST_Z.n3 RST_Z.t2 175.169
R58609 RST_Z RST_Z.n3 171.174
R58610 RST_Z.n2 RST_Z.n1 167.165
R58611 RST_Z RST_Z.n2 163.993
R58612 RST_Z.n1 RST_Z.t4 158.275
R58613 RST_Z.n2 RST_Z.n0 36.9629
R58614 a_20647_31459.n1 a_20647_31459.t4 594.891
R58615 a_20647_31459.n1 a_20647_31459.n0 380.32
R58616 a_20647_31459.n2 a_20647_31459.n1 185
R58617 a_20647_31459.n0 a_20647_31459.t3 26.5955
R58618 a_20647_31459.n0 a_20647_31459.t2 26.5955
R58619 a_20647_31459.n2 a_20647_31459.t0 24.9236
R58620 a_20647_31459.t1 a_20647_31459.n2 24.9236
R58621 a_1581_43806.n13 a_1581_43806.t21 334.723
R58622 a_1581_43806.n6 a_1581_43806.t11 310.457
R58623 a_1581_43806.n10 a_1581_43806.t12 293.969
R58624 a_1581_43806.n4 a_1581_43806.t14 267.065
R58625 a_1581_43806.n8 a_1581_43806.t18 256.07
R58626 a_1581_43806.n3 a_1581_43806.n1 248.087
R58627 a_1581_43806.n7 a_1581_43806.t13 241.536
R58628 a_1581_43806.n5 a_1581_43806.t19 241.536
R58629 a_1581_43806.n6 a_1581_43806.t15 220.484
R58630 a_1581_43806.n3 a_1581_43806.n2 208.507
R58631 a_1581_43806.n13 a_1581_43806.t17 206.19
R58632 a_1581_43806.n16 a_1581_43806.n4 190.459
R58633 a_1581_43806.n12 a_1581_43806.n6 189.552
R58634 a_1581_43806.n14 a_1581_43806.n13 189.034
R58635 a_1581_43806.n9 a_1581_43806.n8 187.738
R58636 a_1581_43806.n9 a_1581_43806.n7 173.924
R58637 a_1581_43806.n15 a_1581_43806.n5 171.444
R58638 a_1581_43806.n7 a_1581_43806.t16 169.237
R58639 a_1581_43806.n5 a_1581_43806.t9 169.237
R58640 a_1581_43806.n11 a_1581_43806.n10 164.583
R58641 a_1581_43806.n8 a_1581_43806.t10 150.03
R58642 a_1581_43806.n4 a_1581_43806.t8 148.35
R58643 a_1581_43806.n10 a_1581_43806.t20 138.338
R58644 a_1581_43806.n18 a_1581_43806.n0 137.576
R58645 a_1581_43806.n19 a_1581_43806.n18 99.1759
R58646 a_1581_43806.n15 a_1581_43806.n14 50.3303
R58647 a_1581_43806.n12 a_1581_43806.n11 28.4153
R58648 a_1581_43806.n17 a_1581_43806.n3 27.8685
R58649 a_1581_43806.n1 a_1581_43806.t7 26.5955
R58650 a_1581_43806.n1 a_1581_43806.t4 26.5955
R58651 a_1581_43806.n2 a_1581_43806.t5 26.5955
R58652 a_1581_43806.n2 a_1581_43806.t6 26.5955
R58653 a_1581_43806.n18 a_1581_43806.n17 25.4811
R58654 a_1581_43806.n0 a_1581_43806.t2 24.9236
R58655 a_1581_43806.n0 a_1581_43806.t1 24.9236
R58656 a_1581_43806.t3 a_1581_43806.n19 24.9236
R58657 a_1581_43806.n19 a_1581_43806.t0 24.9236
R58658 a_1581_43806.n11 a_1581_43806.n9 24.5259
R58659 a_1581_43806.n17 a_1581_43806.n16 17.7502
R58660 a_1581_43806.n16 a_1581_43806.n15 7.75649
R58661 a_1581_43806.n14 a_1581_43806.n12 6.18061
R58662 a_2424_46794.n11 a_2424_46794.t1 427.791
R58663 a_2424_46794.n7 a_2424_46794.t8 414.432
R58664 a_2424_46794.n7 a_2424_46794.t2 300.349
R58665 a_2424_46794.n1 a_2424_46794.t10 268.135
R58666 a_2424_46794.n8 a_2424_46794.t9 256.07
R58667 a_2424_46794.n2 a_2424_46794.t11 221.72
R58668 a_2424_46794.t0 a_2424_46794.n11 209.923
R58669 a_2424_46794.n4 a_2424_46794.t5 206.547
R58670 a_2424_46794.n0 a_2424_46794.t4 196.549
R58671 a_2424_46794.n9 a_2424_46794.n8 181.849
R58672 a_2424_46794.n6 a_2424_46794.n0 177.244
R58673 a_2424_46794.n5 a_2424_46794.n1 175.041
R58674 a_2424_46794.n5 a_2424_46794.n4 152
R58675 a_2424_46794.n8 a_2424_46794.t7 150.03
R58676 a_2424_46794.n3 a_2424_46794.t3 149.421
R58677 a_2424_46794.n0 a_2424_46794.t6 148.35
R58678 a_2424_46794.n9 a_2424_46794.n7 127.868
R58679 a_2424_46794.n6 a_2424_46794.n5 46.7605
R58680 a_2424_46794.n2 a_2424_46794.n1 28.5635
R58681 a_2424_46794.n10 a_2424_46794.n9 20.0009
R58682 a_2424_46794.n3 a_2424_46794.n2 17.8524
R58683 a_2424_46794.n4 a_2424_46794.n3 17.8524
R58684 a_2424_46794.n11 a_2424_46794.n10 15.324
R58685 a_2424_46794.n10 a_2424_46794.n6 10.7804
R58686 a_5923_31099.n2 a_5923_31099.t5 582.686
R58687 a_5923_31099.n2 a_5923_31099.t7 579.407
R58688 a_5923_31099.n4 a_5923_31099.n0 380.32
R58689 a_5923_31099.n1 a_5923_31099.t6 260.322
R58690 a_5923_31099.n5 a_5923_31099.n4 185
R58691 a_5923_31099.n1 a_5923_31099.t4 175.169
R58692 a_5923_31099.n3 a_5923_31099.n1 169.41
R58693 a_5923_31099.n3 a_5923_31099.n2 125.022
R58694 a_5923_31099.n0 a_5923_31099.t2 26.5955
R58695 a_5923_31099.n0 a_5923_31099.t3 26.5955
R58696 a_5923_31099.t1 a_5923_31099.n5 24.9236
R58697 a_5923_31099.n5 a_5923_31099.t0 24.9236
R58698 a_5923_31099.n4 a_5923_31099.n3 20.8769
R58699 a_n4515_30659.n0 a_n4515_30659.t17 756.547
R58700 a_n4515_30659.n14 a_n4515_30659.t16 756.226
R58701 a_n4515_30659.n13 a_n4515_30659.t8 756.226
R58702 a_n4515_30659.n12 a_n4515_30659.t10 756.226
R58703 a_n4515_30659.n11 a_n4515_30659.t9 756.226
R58704 a_n4515_30659.n10 a_n4515_30659.t15 756.226
R58705 a_n4515_30659.n9 a_n4515_30659.t13 756.226
R58706 a_n4515_30659.n8 a_n4515_30659.t7 756.226
R58707 a_n4515_30659.n7 a_n4515_30659.t4 756.226
R58708 a_n4515_30659.n6 a_n4515_30659.t11 756.226
R58709 a_n4515_30659.n5 a_n4515_30659.t6 756.226
R58710 a_n4515_30659.n4 a_n4515_30659.t18 756.226
R58711 a_n4515_30659.n3 a_n4515_30659.t14 756.226
R58712 a_n4515_30659.n2 a_n4515_30659.t12 756.226
R58713 a_n4515_30659.n1 a_n4515_30659.t5 756.226
R58714 a_n4515_30659.n0 a_n4515_30659.t19 756.226
R58715 a_n4515_30659.n16 a_n4515_30659.n15 380.32
R58716 a_n4515_30659.n17 a_n4515_30659.n16 185
R58717 a_n4515_30659.n16 a_n4515_30659.n14 107.011
R58718 a_n4515_30659.n15 a_n4515_30659.t2 26.5955
R58719 a_n4515_30659.n15 a_n4515_30659.t3 26.5955
R58720 a_n4515_30659.n17 a_n4515_30659.t0 24.9236
R58721 a_n4515_30659.t1 a_n4515_30659.n17 24.9236
R58722 a_n4515_30659.n1 a_n4515_30659.n0 0.3205
R58723 a_n4515_30659.n2 a_n4515_30659.n1 0.3205
R58724 a_n4515_30659.n3 a_n4515_30659.n2 0.3205
R58725 a_n4515_30659.n4 a_n4515_30659.n3 0.3205
R58726 a_n4515_30659.n5 a_n4515_30659.n4 0.3205
R58727 a_n4515_30659.n6 a_n4515_30659.n5 0.3205
R58728 a_n4515_30659.n7 a_n4515_30659.n6 0.3205
R58729 a_n4515_30659.n8 a_n4515_30659.n7 0.3205
R58730 a_n4515_30659.n9 a_n4515_30659.n8 0.3205
R58731 a_n4515_30659.n10 a_n4515_30659.n9 0.3205
R58732 a_n4515_30659.n11 a_n4515_30659.n10 0.3205
R58733 a_n4515_30659.n12 a_n4515_30659.n11 0.3205
R58734 a_n4515_30659.n13 a_n4515_30659.n12 0.3205
R58735 a_n4515_30659.n14 a_n4515_30659.n13 0.303833
R58736 DATA[5].n3 DATA[5].n2 647.148
R58737 DATA[5].n5 DATA[5].n4 200.262
R58738 DATA[5].n3 DATA[5].n1 194.441
R58739 DATA[5].n6 DATA[5].n0 185
R58740 DATA[5].n6 DATA[5].n5 58.6278
R58741 DATA[5].n5 DATA[5].n3 50.5705
R58742 DATA[5].n0 DATA[5].t0 40.0005
R58743 DATA[5].n0 DATA[5].t2 40.0005
R58744 DATA[5].n4 DATA[5].t3 40.0005
R58745 DATA[5].n4 DATA[5].t1 40.0005
R58746 DATA[5].n1 DATA[5].t6 27.5805
R58747 DATA[5].n1 DATA[5].t5 27.5805
R58748 DATA[5].n2 DATA[5].t7 27.5805
R58749 DATA[5].n2 DATA[5].t4 27.5805
R58750 DATA[5] DATA[5].n6 15.6247
R58751 a_3754_38470.n3 a_3754_38470.t9 542.561
R58752 a_3754_38470.n1 a_3754_38470.t8 542.561
R58753 a_3754_38470.n0 a_3754_38470.t10 542.561
R58754 a_3754_38470.n6 a_3754_38470.t7 542.545
R58755 a_3754_38470.n3 a_3754_38470.t4 542.081
R58756 a_3754_38470.n5 a_3754_38470.t5 542.081
R58757 a_3754_38470.n1 a_3754_38470.t3 542.081
R58758 a_3754_38470.n0 a_3754_38470.t6 542.081
R58759 a_3754_38470.t0 a_3754_38470.n8 100.382
R58760 a_3754_38470.n8 a_3754_38470.t1 44.988
R58761 a_3754_38470.n7 a_3754_38470.t2 44.0791
R58762 a_3754_38470.n8 a_3754_38470.n7 18.1307
R58763 a_3754_38470.n7 a_3754_38470.n6 2.16717
R58764 a_3754_38470.n4 a_3754_38470.n2 1.438
R58765 a_3754_38470.n4 a_3754_38470.n3 0.703
R58766 a_3754_38470.n2 a_3754_38470.n0 0.588
R58767 a_3754_38470.n2 a_3754_38470.n1 0.463
R58768 a_3754_38470.n5 a_3754_38470.n4 0.348
R58769 a_3754_38470.n6 a_3754_38470.n5 0.0155
R58770 a_17564_32305.n1 a_17564_32305.t4 1688.87
R58771 a_17564_32305.n1 a_17564_32305.n0 287.752
R58772 a_17564_32305.n2 a_17564_32305.n1 277.568
R58773 a_17564_32305.n0 a_17564_32305.t2 26.5955
R58774 a_17564_32305.n0 a_17564_32305.t3 26.5955
R58775 a_17564_32305.n2 a_17564_32305.t0 24.9236
R58776 a_17564_32305.t1 a_17564_32305.n2 24.9236
R58777 a_4830_43958.n15 a_4830_43958.n0 659.109
R58778 a_4830_43958.n9 a_4830_43958.t7 294.557
R58779 a_4830_43958.n7 a_4830_43958.t9 294.557
R58780 a_4830_43958.n5 a_4830_43958.t12 294.557
R58781 a_4830_43958.n4 a_4830_43958.t10 294.557
R58782 a_4830_43958.n1 a_4830_43958.t14 260.322
R58783 a_4830_43958.n3 a_4830_43958.t4 224.984
R58784 a_4830_43958.n13 a_4830_43958.t17 224.984
R58785 a_4830_43958.n16 a_4830_43958.n15 219.663
R58786 a_4830_43958.n9 a_4830_43958.t11 211.01
R58787 a_4830_43958.n7 a_4830_43958.t15 211.01
R58788 a_4830_43958.n5 a_4830_43958.t6 211.01
R58789 a_4830_43958.n4 a_4830_43958.t16 211.01
R58790 a_4830_43958.n3 a_4830_43958.t8 187.714
R58791 a_4830_43958.n13 a_4830_43958.t18 187.714
R58792 a_4830_43958.n6 a_4830_43958.n4 186.798
R58793 a_4830_43958.n8 a_4830_43958.n7 185.786
R58794 a_4830_43958.n14 a_4830_43958.n13 181.548
R58795 a_4830_43958.n11 a_4830_43958.n3 181.03
R58796 a_4830_43958.n10 a_4830_43958.n9 179.332
R58797 a_4830_43958.n1 a_4830_43958.t5 175.169
R58798 a_4830_43958.n2 a_4830_43958.n1 164.45
R58799 a_4830_43958.n6 a_4830_43958.n5 162.398
R58800 a_4830_43958.n2 a_4830_43958.t13 59.3472
R58801 a_4830_43958.t1 a_4830_43958.n16 38.5719
R58802 a_4830_43958.n16 a_4830_43958.t0 38.5719
R58803 a_4830_43958.n0 a_4830_43958.t2 26.5955
R58804 a_4830_43958.n0 a_4830_43958.t3 26.5955
R58805 a_4830_43958.n12 a_4830_43958.n2 14.6118
R58806 a_4830_43958.n15 a_4830_43958.n14 14.0946
R58807 a_4830_43958.n8 a_4830_43958.n6 10.7764
R58808 a_4830_43958.n11 a_4830_43958.n10 7.66376
R58809 a_4830_43958.n10 a_4830_43958.n8 4.72577
R58810 a_4830_43958.n14 a_4830_43958.n12 3.48639
R58811 a_4830_43958.n12 a_4830_43958.n11 1.58127
R58812 C4_P_btm.n1 C4_P_btm.t22 101.361
R58813 C4_P_btm.n2 C4_P_btm.t2 98.3735
R58814 C4_P_btm.n0 C4_P_btm.t0 54.9311
R58815 C4_P_btm C4_P_btm.n2 54.563
R58816 C4_P_btm.n0 C4_P_btm.t1 47.3635
R58817 C4_P_btm.n2 C4_P_btm.n1 8.08383
R58818 C4_P_btm C4_P_btm.n22 7.74425
R58819 C4_P_btm.n1 C4_P_btm.n0 7.15154
R58820 C4_P_btm.n18 C4_P_btm.t5 5.03712
R58821 C4_P_btm.n4 C4_P_btm.t3 5.03712
R58822 C4_P_btm.n4 C4_P_btm.t13 4.03712
R58823 C4_P_btm.n5 C4_P_btm.t14 4.03712
R58824 C4_P_btm.n6 C4_P_btm.t12 4.03712
R58825 C4_P_btm.n15 C4_P_btm.t11 4.03712
R58826 C4_P_btm.n22 C4_P_btm.t4 4.03712
R58827 C4_P_btm.n20 C4_P_btm.t16 3.98193
R58828 C4_P_btm.n14 C4_P_btm.t7 3.98193
R58829 C4_P_btm.n7 C4_P_btm.t6 3.98193
R58830 C4_P_btm.n3 C4_P_btm.t8 3.98193
R58831 C4_P_btm.n16 C4_P_btm.t10 3.98193
R58832 C4_P_btm.n19 C4_P_btm.t18 3.98193
R58833 C4_P_btm.n13 C4_P_btm.t19 3.92851
R58834 C4_P_btm.n12 C4_P_btm.t9 3.92851
R58835 C4_P_btm.n11 C4_P_btm.t21 3.92851
R58836 C4_P_btm.n10 C4_P_btm.t17 3.92851
R58837 C4_P_btm.n9 C4_P_btm.t20 3.92851
R58838 C4_P_btm.n8 C4_P_btm.t15 3.92851
R58839 C4_P_btm.n7 C4_P_btm.n6 1.05569
R58840 C4_P_btm.n15 C4_P_btm.n14 1.05569
R58841 C4_P_btm.n21 C4_P_btm.n3 1.05569
R58842 C4_P_btm.n5 C4_P_btm.n4 1.0005
R58843 C4_P_btm.n6 C4_P_btm.n5 1.0005
R58844 C4_P_btm.n17 C4_P_btm.n15 1.0005
R58845 C4_P_btm.n18 C4_P_btm.n17 1.0005
R58846 C4_P_btm.n22 C4_P_btm.n21 1.0005
R58847 C4_P_btm.n9 C4_P_btm.n8 0.840176
R58848 C4_P_btm.n10 C4_P_btm.n9 0.840176
R58849 C4_P_btm.n11 C4_P_btm.n10 0.840176
R58850 C4_P_btm.n12 C4_P_btm.n11 0.840176
R58851 C4_P_btm.n13 C4_P_btm.n12 0.840176
R58852 C4_P_btm.n8 C4_P_btm.n7 0.786757
R58853 C4_P_btm.n14 C4_P_btm.n13 0.786757
R58854 C4_P_btm.n16 C4_P_btm.n3 0.733338
R58855 C4_P_btm.n20 C4_P_btm.n19 0.733338
R58856 C4_P_btm.n17 C4_P_btm.n16 0.0556875
R58857 C4_P_btm.n19 C4_P_btm.n18 0.0556875
R58858 C4_P_btm.n21 C4_P_btm.n20 0.0556875
R58859 VIN_P.n1 VIN_P.t3 92.1604
R58860 VIN_P.n3 VIN_P.t0 91.0227
R58861 VIN_P.n7 VIN_P.t5 90.7102
R58862 VIN_P.n6 VIN_P.t2 90.7102
R58863 VIN_P.n5 VIN_P.t1 90.7102
R58864 VIN_P.n4 VIN_P.t7 90.7102
R58865 VIN_P.n1 VIN_P.t4 90.6265
R58866 VIN_P.n2 VIN_P.t6 90.6219
R58867 VIN_P.n10 VIN_P.t11 47.4586
R58868 VIN_P.n9 VIN_P.n8 37.5586
R58869 VIN_P.n14 VIN_P.n12 32.094
R58870 VIN_P.n13 VIN_P.t14 25.3459
R58871 VIN_P.n13 VIN_P.t13 25.1217
R58872 VIN_P.n14 VIN_P.n13 17.3942
R58873 VIN_P.n12 VIN_P.t8 16.5266
R58874 VIN_P.n11 VIN_P.n0 14.0516
R58875 VIN_P.n11 VIN_P.n10 11.2899
R58876 VIN_P VIN_P.n14 10.1163
R58877 VIN_P.n8 VIN_P.t15 9.9005
R58878 VIN_P.n8 VIN_P.t10 9.9005
R58879 VIN_P.n0 VIN_P.t12 2.4755
R58880 VIN_P.n0 VIN_P.t9 2.4755
R58881 VIN_P.n2 VIN_P.n1 1.6255
R58882 VIN_P.n3 VIN_P.n2 1.2505
R58883 VIN_P.n9 VIN_P.n7 0.8755
R58884 VIN_P.n5 VIN_P.n4 0.563
R58885 VIN_P.n6 VIN_P.n5 0.563
R58886 VIN_P.n7 VIN_P.n6 0.563
R58887 VIN_P.n10 VIN_P.n9 0.453625
R58888 VIN_P.n12 VIN_P.n11 0.438
R58889 VIN_P.n4 VIN_P.n3 0.2505
R58890 CAL_P.n5 CAL_P.n4 601.067
R58891 CAL_P.n5 CAL_P.t1 251.581
R58892 CAL_P CAL_P.t6 137
R58893 CAL_P.n4 CAL_P.t0 77.3934
R58894 CAL_P.n4 CAL_P.t2 77.3934
R58895 CAL_P.n1 CAL_P.t4 36.3712
R58896 CAL_P.t5 CAL_P.n0 36.2721
R58897 CAL_P.n2 CAL_P.t4 35.5162
R58898 CAL_P.n3 CAL_P.t5 35.4454
R58899 CAL_P.n2 CAL_P.t3 31.2287
R58900 CAL_P.t3 CAL_P.n1 31.2287
R58901 CAL_P CAL_P.n6 25.3442
R58902 CAL_P.n6 CAL_P.n5 8.34425
R58903 CAL_P.n6 CAL_P.n3 7.5005
R58904 CAL_P.n6 CAL_P.n0 5.95883
R58905 CAL_P.n1 CAL_P.n0 0.0713333
R58906 CAL_P.n3 CAL_P.n2 0.0713333
R58907 a_n2497_42870.n3 a_n2497_42870.n2 291.312
R58908 a_n2497_42870.n6 a_n2497_42870.n0 273.32
R58909 a_n2497_42870.n1 a_n2497_42870.t9 238.59
R58910 a_n2497_42870.n3 a_n2497_42870.n1 220.887
R58911 a_n2497_42870.n1 a_n2497_42870.t8 203.244
R58912 a_n2497_42870.n7 a_n2497_42870.n6 190.726
R58913 a_n2497_42870.n5 a_n2497_42870.n4 96.3105
R58914 a_n2497_42870.n6 a_n2497_42870.n5 47.8
R58915 a_n2497_42870.n5 a_n2497_42870.n3 45.4744
R58916 a_n2497_42870.n2 a_n2497_42870.t5 27.5805
R58917 a_n2497_42870.n2 a_n2497_42870.t4 27.5805
R58918 a_n2497_42870.n0 a_n2497_42870.t2 25.8467
R58919 a_n2497_42870.n0 a_n2497_42870.t3 25.8467
R58920 a_n2497_42870.n4 a_n2497_42870.t6 25.8467
R58921 a_n2497_42870.n4 a_n2497_42870.t7 25.8467
R58922 a_n2497_42870.n7 a_n2497_42870.t0 25.8467
R58923 a_n2497_42870.t1 a_n2497_42870.n7 25.8467
R58924 a_19679_31459.n1 a_19679_31459.t4 595.367
R58925 a_19679_31459.n1 a_19679_31459.n0 380.32
R58926 a_19679_31459.n2 a_19679_31459.n1 185
R58927 a_19679_31459.n0 a_19679_31459.t2 26.5955
R58928 a_19679_31459.n0 a_19679_31459.t3 26.5955
R58929 a_19679_31459.t1 a_19679_31459.n2 24.9236
R58930 a_19679_31459.n2 a_19679_31459.t0 24.9236
R58931 a_18394_35068.n3 a_18394_35068.t11 749.612
R58932 a_18394_35068.n9 a_18394_35068.t14 748.122
R58933 a_18394_35068.n7 a_18394_35068.t9 748.122
R58934 a_18394_35068.n5 a_18394_35068.t8 684.441
R58935 a_18394_35068.n3 a_18394_35068.t10 684.441
R58936 a_18394_35068.n4 a_18394_35068.t13 684.441
R58937 a_18394_35068.n9 a_18394_35068.t15 678.014
R58938 a_18394_35068.n7 a_18394_35068.t12 678.014
R58939 a_18394_35068.n14 a_18394_35068.n13 244.067
R58940 a_18394_35068.n2 a_18394_35068.n0 236.589
R58941 a_18394_35068.n13 a_18394_35068.n12 204.893
R58942 a_18394_35068.n2 a_18394_35068.n1 200.321
R58943 a_18394_35068.n8 a_18394_35068.n7 163.538
R58944 a_18394_35068.n10 a_18394_35068.n9 163.538
R58945 a_18394_35068.n6 a_18394_35068.n5 161.513
R58946 a_18394_35068.n6 a_18394_35068.n3 161.487
R58947 a_18394_35068.n5 a_18394_35068.n4 65.1723
R58948 a_18394_35068.n4 a_18394_35068.n3 65.1723
R58949 a_18394_35068.n11 a_18394_35068.n2 26.8022
R58950 a_18394_35068.n12 a_18394_35068.t3 26.5955
R58951 a_18394_35068.n12 a_18394_35068.t6 26.5955
R58952 a_18394_35068.n14 a_18394_35068.t5 26.5955
R58953 a_18394_35068.t0 a_18394_35068.n14 26.5955
R58954 a_18394_35068.n13 a_18394_35068.n11 25.4552
R58955 a_18394_35068.n0 a_18394_35068.t7 24.9236
R58956 a_18394_35068.n0 a_18394_35068.t4 24.9236
R58957 a_18394_35068.n1 a_18394_35068.t2 24.9236
R58958 a_18394_35068.n1 a_18394_35068.t1 24.9236
R58959 a_18394_35068.n8 a_18394_35068.n6 7.92231
R58960 a_18394_35068.n11 a_18394_35068.n10 5.93105
R58961 a_18394_35068.n10 a_18394_35068.n8 2.47042
R58962 SMPL.n2 SMPL.n1 647.148
R58963 SMPL.n5 SMPL.n3 243.627
R58964 SMPL.n19 SMPL.t23 212.081
R58965 SMPL.n21 SMPL.t9 212.081
R58966 SMPL.n23 SMPL.t22 212.081
R58967 SMPL.n17 SMPL.t12 212.081
R58968 SMPL.n7 SMPL.t17 212.081
R58969 SMPL.n13 SMPL.t8 212.081
R58970 SMPL.n11 SMPL.t14 212.081
R58971 SMPL.n9 SMPL.t19 212.081
R58972 SMPL.n5 SMPL.n4 200.262
R58973 SMPL.n26 SMPL.n17 194.47
R58974 SMPL.n16 SMPL.n7 194.47
R58975 SMPL.n2 SMPL.n0 194.441
R58976 SMPL.n20 SMPL.n18 173.505
R58977 SMPL.n10 SMPL.n8 173.505
R58978 SMPL.n27 SMPL.n16 162.155
R58979 SMPL.n25 SMPL.n24 152
R58980 SMPL.n22 SMPL.n18 152
R58981 SMPL.n12 SMPL.n8 152
R58982 SMPL.n15 SMPL.n14 152
R58983 SMPL.n19 SMPL.t18 139.78
R58984 SMPL.n21 SMPL.t21 139.78
R58985 SMPL.n23 SMPL.t13 139.78
R58986 SMPL.n17 SMPL.t15 139.78
R58987 SMPL.n7 SMPL.t20 139.78
R58988 SMPL.n13 SMPL.t16 139.78
R58989 SMPL.n11 SMPL.t11 139.78
R58990 SMPL.n9 SMPL.t10 139.78
R58991 SMPL.n6 SMPL.n2 42.8458
R58992 SMPL.n3 SMPL.t0 40.0005
R58993 SMPL.n3 SMPL.t1 40.0005
R58994 SMPL.n4 SMPL.t2 40.0005
R58995 SMPL.n4 SMPL.t3 40.0005
R58996 SMPL.n27 SMPL.n26 39.6921
R58997 SMPL.n20 SMPL.n19 30.6732
R58998 SMPL.n21 SMPL.n20 30.6732
R58999 SMPL.n22 SMPL.n21 30.6732
R59000 SMPL.n23 SMPL.n22 30.6732
R59001 SMPL.n24 SMPL.n23 30.6732
R59002 SMPL.n24 SMPL.n17 30.6732
R59003 SMPL.n14 SMPL.n7 30.6732
R59004 SMPL.n14 SMPL.n13 30.6732
R59005 SMPL.n13 SMPL.n12 30.6732
R59006 SMPL.n12 SMPL.n11 30.6732
R59007 SMPL.n11 SMPL.n10 30.6732
R59008 SMPL.n10 SMPL.n9 30.6732
R59009 SMPL.n0 SMPL.t6 27.5805
R59010 SMPL.n0 SMPL.t5 27.5805
R59011 SMPL.n1 SMPL.t7 27.5805
R59012 SMPL.n1 SMPL.t4 27.5805
R59013 SMPL.n25 SMPL.n18 21.5045
R59014 SMPL.n15 SMPL.n8 21.5045
R59015 SMPL SMPL.n6 18.7273
R59016 SMPL.n26 SMPL.n25 8.08129
R59017 SMPL.n16 SMPL.n15 8.08128
R59018 SMPL.n6 SMPL.n5 7.72512
R59019 SMPL SMPL.n27 4.64857
R59020 a_6485_44582.t12 a_6485_44582.t14 378.255
R59021 a_6485_44582.n5 a_6485_44582.t12 362.913
R59022 a_6485_44582.n4 a_6485_44582.t27 334.723
R59023 a_6485_44582.n11 a_6485_44582.t10 323.342
R59024 a_6485_44582.n10 a_6485_44582.t9 256.726
R59025 a_6485_44582.n3 a_6485_44582.n1 248.087
R59026 a_6485_44582.n19 a_6485_44582.t19 241.536
R59027 a_6485_44582.n15 a_6485_44582.t26 238.397
R59028 a_6485_44582.n18 a_6485_44582.t8 231.835
R59029 a_6485_44582.n6 a_6485_44582.t18 221.72
R59030 a_6485_44582.n7 a_6485_44582.t20 221.72
R59031 a_6485_44582.n3 a_6485_44582.n2 208.507
R59032 a_6485_44582.n4 a_6485_44582.t13 206.19
R59033 a_6485_44582.n15 a_6485_44582.t16 195.017
R59034 a_6485_44582.n11 a_6485_44582.t24 194.809
R59035 a_6485_44582.n5 a_6485_44582.n4 188.506
R59036 a_6485_44582.n20 a_6485_44582.n19 184.362
R59037 a_6485_44582.n12 a_6485_44582.n11 182.215
R59038 a_6485_44582.n12 a_6485_44582.n10 175.758
R59039 a_6485_44582.n19 a_6485_44582.t11 169.237
R59040 a_6485_44582.n20 a_6485_44582.n18 168.621
R59041 a_6485_44582.n9 a_6485_44582.n8 166.101
R59042 a_6485_44582.n14 a_6485_44582.n13 162.837
R59043 a_6485_44582.n16 a_6485_44582.n15 161.981
R59044 a_6485_44582.n10 a_6485_44582.t15 161.275
R59045 a_6485_44582.n18 a_6485_44582.t23 157.07
R59046 a_6485_44582.n6 a_6485_44582.t25 149.421
R59047 a_6485_44582.n7 a_6485_44582.t17 149.421
R59048 a_6485_44582.n23 a_6485_44582.n0 137.576
R59049 a_6485_44582.n13 a_6485_44582.t22 137.177
R59050 a_6485_44582.n13 a_6485_44582.t21 121.109
R59051 a_6485_44582.n24 a_6485_44582.n23 99.1759
R59052 a_6485_44582.n22 a_6485_44582.n3 38.4831
R59053 a_6485_44582.n8 a_6485_44582.n6 37.4894
R59054 a_6485_44582.n8 a_6485_44582.n7 37.4894
R59055 a_6485_44582.n1 a_6485_44582.t7 26.5955
R59056 a_6485_44582.n1 a_6485_44582.t4 26.5955
R59057 a_6485_44582.n2 a_6485_44582.t6 26.5955
R59058 a_6485_44582.n2 a_6485_44582.t5 26.5955
R59059 a_6485_44582.n0 a_6485_44582.t0 24.9236
R59060 a_6485_44582.n0 a_6485_44582.t1 24.9236
R59061 a_6485_44582.n24 a_6485_44582.t2 24.9236
R59062 a_6485_44582.t3 a_6485_44582.n24 24.9236
R59063 a_6485_44582.n16 a_6485_44582.n14 17.4485
R59064 a_6485_44582.n23 a_6485_44582.n22 14.8665
R59065 a_6485_44582.n9 a_6485_44582.n5 12.4702
R59066 a_6485_44582.n21 a_6485_44582.n17 10.131
R59067 a_6485_44582.n22 a_6485_44582.n21 9.3005
R59068 a_6485_44582.n17 a_6485_44582.n16 7.48535
R59069 a_6485_44582.n17 a_6485_44582.n9 6.7972
R59070 a_6485_44582.n21 a_6485_44582.n20 6.68663
R59071 a_6485_44582.n14 a_6485_44582.n12 2.19246
R59072 a_5700_37509.n8 a_5700_37509.t17 120.882
R59073 a_5700_37509.n9 a_5700_37509.t16 120.57
R59074 a_5700_37509.n8 a_5700_37509.n7 104.317
R59075 a_5700_37509.n17 a_5700_37509.n16 39.965
R59076 a_5700_37509.n2 a_5700_37509.n0 39.792
R59077 a_5700_37509.n12 a_5700_37509.n11 39.6681
R59078 a_5700_37509.n14 a_5700_37509.n13 39.6681
R59079 a_5700_37509.n16 a_5700_37509.n15 39.6681
R59080 a_5700_37509.n6 a_5700_37509.n5 39.4951
R59081 a_5700_37509.n4 a_5700_37509.n3 39.4951
R59082 a_5700_37509.n2 a_5700_37509.n1 39.4951
R59083 a_5700_37509.n7 a_5700_37509.t18 16.253
R59084 a_5700_37509.n7 a_5700_37509.t19 16.253
R59085 a_5700_37509.n12 a_5700_37509.n10 14.9015
R59086 a_5700_37509.n10 a_5700_37509.n9 14.0786
R59087 a_5700_37509.n11 a_5700_37509.t8 4.76133
R59088 a_5700_37509.n11 a_5700_37509.t10 4.76133
R59089 a_5700_37509.n13 a_5700_37509.t14 4.76133
R59090 a_5700_37509.n13 a_5700_37509.t0 4.76133
R59091 a_5700_37509.n15 a_5700_37509.t6 4.76133
R59092 a_5700_37509.n15 a_5700_37509.t7 4.76133
R59093 a_5700_37509.n5 a_5700_37509.t9 4.76133
R59094 a_5700_37509.n5 a_5700_37509.t1 4.76133
R59095 a_5700_37509.n3 a_5700_37509.t4 4.76133
R59096 a_5700_37509.n3 a_5700_37509.t13 4.76133
R59097 a_5700_37509.n1 a_5700_37509.t3 4.76133
R59098 a_5700_37509.n1 a_5700_37509.t12 4.76133
R59099 a_5700_37509.n0 a_5700_37509.t5 4.76133
R59100 a_5700_37509.n0 a_5700_37509.t11 4.76133
R59101 a_5700_37509.n17 a_5700_37509.t2 4.76133
R59102 a_5700_37509.t15 a_5700_37509.n17 4.76133
R59103 a_5700_37509.n10 a_5700_37509.n6 1.96925
R59104 a_5700_37509.n4 a_5700_37509.n2 0.313
R59105 a_5700_37509.n6 a_5700_37509.n4 0.313
R59106 a_5700_37509.n16 a_5700_37509.n14 0.313
R59107 a_5700_37509.n14 a_5700_37509.n12 0.313
R59108 a_5700_37509.n9 a_5700_37509.n8 0.297375
R59109 CLK_DATA.n5 CLK_DATA.n4 647.148
R59110 CLK_DATA.n2 CLK_DATA.n0 243.627
R59111 CLK_DATA.n2 CLK_DATA.n1 200.262
R59112 CLK_DATA.n5 CLK_DATA.n3 194.441
R59113 CLK_DATA.n6 CLK_DATA.n5 42.8458
R59114 CLK_DATA.n0 CLK_DATA.t1 40.0005
R59115 CLK_DATA.n0 CLK_DATA.t2 40.0005
R59116 CLK_DATA.n1 CLK_DATA.t0 40.0005
R59117 CLK_DATA.n1 CLK_DATA.t3 40.0005
R59118 CLK_DATA.n3 CLK_DATA.t7 27.5805
R59119 CLK_DATA.n3 CLK_DATA.t5 27.5805
R59120 CLK_DATA.n4 CLK_DATA.t6 27.5805
R59121 CLK_DATA.n4 CLK_DATA.t4 27.5805
R59122 CLK_DATA CLK_DATA.n6 15.0398
R59123 CLK_DATA.n6 CLK_DATA.n2 7.72512
R59124 a_n2497_47846.n0 a_n2497_47846.t6 241.536
R59125 a_n2497_47846.n1 a_n2497_47846.t7 238.59
R59126 a_n2497_47846.n2 a_n2497_47846.t3 230.793
R59127 a_n2497_47846.n5 a_n2497_47846.t1 223.441
R59128 a_n2497_47846.n3 a_n2497_47846.n1 207.612
R59129 a_n2497_47846.n1 a_n2497_47846.t4 203.244
R59130 a_n2497_47846.n3 a_n2497_47846.n2 178.3
R59131 a_n2497_47846.n4 a_n2497_47846.n0 177.918
R59132 a_n2497_47846.n6 a_n2497_47846.n5 175.649
R59133 a_n2497_47846.n0 a_n2497_47846.t5 169.237
R59134 a_n2497_47846.n2 a_n2497_47846.t8 158.494
R59135 a_n2497_47846.t0 a_n2497_47846.n6 24.9236
R59136 a_n2497_47846.n6 a_n2497_47846.t2 24.9236
R59137 a_n2497_47846.n5 a_n2497_47846.n4 13.7724
R59138 a_n2497_47846.n4 a_n2497_47846.n3 2.34819
R59139 a_n1925_47044.n5 a_n1925_47044.n0 664.928
R59140 a_n1925_47044.n3 a_n1925_47044.t7 276.464
R59141 a_n1925_47044.n4 a_n1925_47044.n2 221.514
R59142 a_n1925_47044.n1 a_n1925_47044.t4 212.081
R59143 a_n1925_47044.n2 a_n1925_47044.t8 212.081
R59144 a_n1925_47044.n3 a_n1925_47044.t9 196.131
R59145 a_n1925_47044.n4 a_n1925_47044.n3 190.56
R59146 a_n1925_47044.n6 a_n1925_47044.n5 187.927
R59147 a_n1925_47044.n1 a_n1925_47044.t5 139.78
R59148 a_n1925_47044.n2 a_n1925_47044.t6 139.78
R59149 a_n1925_47044.n2 a_n1925_47044.n1 61.346
R59150 a_n1925_47044.n0 a_n1925_47044.t3 26.5955
R59151 a_n1925_47044.n0 a_n1925_47044.t2 26.5955
R59152 a_n1925_47044.t1 a_n1925_47044.n6 24.9236
R59153 a_n1925_47044.n6 a_n1925_47044.t0 24.9236
R59154 a_n1925_47044.n5 a_n1925_47044.n4 18.428
R59155 a_n99_45438.n0 a_n99_45438.t3 471.289
R59156 a_n99_45438.t0 a_n99_45438.n3 349.469
R59157 a_n99_45438.n3 a_n99_45438.t1 338.243
R59158 a_n99_45438.n1 a_n99_45438.t2 224.984
R59159 a_n99_45438.n2 a_n99_45438.n0 213.208
R59160 a_n99_45438.n2 a_n99_45438.n1 189.421
R59161 a_n99_45438.n1 a_n99_45438.t4 187.714
R59162 a_n99_45438.n0 a_n99_45438.t5 148.35
R59163 a_n99_45438.n3 a_n99_45438.n2 18.6721
R59164 a_5334_30651.n2 a_5334_30651.t6 1615.23
R59165 a_5334_30651.n2 a_5334_30651.t7 1614.01
R59166 a_5334_30651.n4 a_5334_30651.n0 380.32
R59167 a_5334_30651.n1 a_5334_30651.t4 260.322
R59168 a_5334_30651.n5 a_5334_30651.n4 185
R59169 a_5334_30651.n3 a_5334_30651.n1 175.222
R59170 a_5334_30651.n1 a_5334_30651.t5 175.169
R59171 a_5334_30651.n3 a_5334_30651.n2 79.9157
R59172 a_5334_30651.n0 a_5334_30651.t2 26.5955
R59173 a_5334_30651.n0 a_5334_30651.t3 26.5955
R59174 a_5334_30651.n5 a_5334_30651.t0 24.9236
R59175 a_5334_30651.t1 a_5334_30651.n5 24.9236
R59176 a_5334_30651.n4 a_5334_30651.n3 18.3786
R59177 a_10114_45276.t2 a_10114_45276.t4 378.255
R59178 a_10114_45276.t6 a_10114_45276.t10 378.255
R59179 a_10114_45276.t3 a_10114_45276.t7 378.255
R59180 a_10114_45276.t9 a_10114_45276.t11 378.255
R59181 a_10114_45276.n1 a_10114_45276.t6 374.745
R59182 a_10114_45276.n5 a_10114_45276.t1 366.548
R59183 a_10114_45276.n2 a_10114_45276.t3 351.127
R59184 a_10114_45276.n4 a_10114_45276.t9 327.175
R59185 a_10114_45276.n1 a_10114_45276.t2 325.223
R59186 a_10114_45276.t0 a_10114_45276.n5 307.562
R59187 a_10114_45276.n0 a_10114_45276.t8 241.536
R59188 a_10114_45276.n3 a_10114_45276.n0 180.82
R59189 a_10114_45276.n0 a_10114_45276.t5 169.237
R59190 a_10114_45276.n5 a_10114_45276.n4 16.7712
R59191 a_10114_45276.n3 a_10114_45276.n2 13.3741
R59192 a_10114_45276.n2 a_10114_45276.n1 9.72319
R59193 a_10114_45276.n4 a_10114_45276.n3 3.41413
R59194 a_21788_30659.n0 a_21788_30659.t6 756.547
R59195 a_21788_30659.n6 a_21788_30659.t5 756.231
R59196 a_21788_30659.n0 a_21788_30659.t10 756.226
R59197 a_21788_30659.n1 a_21788_30659.t8 756.226
R59198 a_21788_30659.n2 a_21788_30659.t9 756.226
R59199 a_21788_30659.n3 a_21788_30659.t4 756.226
R59200 a_21788_30659.n4 a_21788_30659.t11 756.226
R59201 a_21788_30659.n5 a_21788_30659.t7 756.226
R59202 a_21788_30659.n8 a_21788_30659.n7 380.32
R59203 a_21788_30659.n9 a_21788_30659.n8 185
R59204 a_21788_30659.n8 a_21788_30659.n6 106.856
R59205 a_21788_30659.n7 a_21788_30659.t3 26.5955
R59206 a_21788_30659.n7 a_21788_30659.t2 26.5955
R59207 a_21788_30659.t1 a_21788_30659.n9 24.9236
R59208 a_21788_30659.n9 a_21788_30659.t0 24.9236
R59209 a_21788_30659.n5 a_21788_30659.n4 0.3205
R59210 a_21788_30659.n4 a_21788_30659.n3 0.3205
R59211 a_21788_30659.n3 a_21788_30659.n2 0.3205
R59212 a_21788_30659.n2 a_21788_30659.n1 0.3205
R59213 a_21788_30659.n1 a_21788_30659.n0 0.3205
R59214 a_21788_30659.n6 a_21788_30659.n5 0.298833
R59215 a_20405_31459.n1 a_20405_31459.t4 602.967
R59216 a_20405_31459.n1 a_20405_31459.n0 287.752
R59217 a_20405_31459.n2 a_20405_31459.n1 277.568
R59218 a_20405_31459.n0 a_20405_31459.t3 26.5955
R59219 a_20405_31459.n0 a_20405_31459.t2 26.5955
R59220 a_20405_31459.n2 a_20405_31459.t0 24.9236
R59221 a_20405_31459.t1 a_20405_31459.n2 24.9236
R59222 DATA[4].n3 DATA[4].n2 647.148
R59223 DATA[4].n5 DATA[4].n4 200.262
R59224 DATA[4].n3 DATA[4].n1 194.441
R59225 DATA[4].n6 DATA[4].n0 185
R59226 DATA[4].n6 DATA[4].n5 58.6278
R59227 DATA[4].n5 DATA[4].n3 50.5705
R59228 DATA[4].n0 DATA[4].t0 40.0005
R59229 DATA[4].n0 DATA[4].t2 40.0005
R59230 DATA[4].n4 DATA[4].t3 40.0005
R59231 DATA[4].n4 DATA[4].t1 40.0005
R59232 DATA[4].n1 DATA[4].t6 27.5805
R59233 DATA[4].n1 DATA[4].t5 27.5805
R59234 DATA[4].n2 DATA[4].t7 27.5805
R59235 DATA[4].n2 DATA[4].t4 27.5805
R59236 DATA[4] DATA[4].n6 15.6247
R59237 a_n2810_46526.n1 a_n2810_46526.t4 871.097
R59238 a_n2810_46526.n1 a_n2810_46526.n0 380.32
R59239 a_n2810_46526.n2 a_n2810_46526.n1 185
R59240 a_n2810_46526.n0 a_n2810_46526.t2 26.5955
R59241 a_n2810_46526.n0 a_n2810_46526.t3 26.5955
R59242 a_n2810_46526.t1 a_n2810_46526.n2 24.9236
R59243 a_n2810_46526.n2 a_n2810_46526.t0 24.9236
R59244 COMP_N.n7 COMP_N.t9 260.322
R59245 COMP_N.n5 COMP_N.n3 244.069
R59246 COMP_N.n2 COMP_N.n0 236.589
R59247 COMP_N COMP_N.n7 230.381
R59248 COMP_N.n5 COMP_N.n4 204.893
R59249 COMP_N.n2 COMP_N.n1 200.321
R59250 COMP_N.n7 COMP_N.t8 175.169
R59251 COMP_N.n6 COMP_N.n5 29.5768
R59252 COMP_N.n6 COMP_N.n2 28.0395
R59253 COMP_N.n4 COMP_N.t5 26.5955
R59254 COMP_N.n4 COMP_N.t6 26.5955
R59255 COMP_N.n3 COMP_N.t4 26.5955
R59256 COMP_N.n3 COMP_N.t7 26.5955
R59257 COMP_N.n0 COMP_N.t1 24.9236
R59258 COMP_N.n0 COMP_N.t0 24.9236
R59259 COMP_N.n1 COMP_N.t3 24.9236
R59260 COMP_N.n1 COMP_N.t2 24.9236
R59261 COMP_N COMP_N.n6 14.5974
R59262 VDAC_Pi VDAC_Pi.t9 388.01
R59263 VDAC_Pi.n3 VDAC_Pi.t10 234.685
R59264 VDAC_Pi.n2 VDAC_Pi.n0 104.316
R59265 VDAC_Pi.n2 VDAC_Pi.n1 104.019
R59266 VDAC_Pi.n3 VDAC_Pi.t8 50.2666
R59267 VDAC_Pi.n8 VDAC_Pi.n7 37.3277
R59268 VDAC_Pi.n6 VDAC_Pi.n5 37.3277
R59269 VDAC_Pi.n1 VDAC_Pi.t7 16.253
R59270 VDAC_Pi.n1 VDAC_Pi.t5 16.253
R59271 VDAC_Pi.n0 VDAC_Pi.t4 16.253
R59272 VDAC_Pi.n0 VDAC_Pi.t6 16.253
R59273 VDAC_Pi VDAC_Pi.n8 14.5151
R59274 VDAC_Pi.n7 VDAC_Pi.t2 9.9005
R59275 VDAC_Pi.n7 VDAC_Pi.t3 9.9005
R59276 VDAC_Pi.n5 VDAC_Pi.t0 9.9005
R59277 VDAC_Pi.n5 VDAC_Pi.t1 9.9005
R59278 VDAC_Pi.n4 VDAC_Pi.n3 6.15675
R59279 VDAC_Pi.n4 VDAC_Pi.n2 1.46925
R59280 VDAC_Pi.n6 VDAC_Pi.n4 0.359875
R59281 VDAC_Pi.n8 VDAC_Pi.n6 0.297375
R59282 a_13458_32299.n1 a_13458_32299.t4 689.486
R59283 a_13458_32299.n1 a_13458_32299.n0 287.752
R59284 a_13458_32299.n2 a_13458_32299.n1 277.568
R59285 a_13458_32299.n0 a_13458_32299.t2 26.5955
R59286 a_13458_32299.n0 a_13458_32299.t3 26.5955
R59287 a_13458_32299.t1 a_13458_32299.n2 24.9236
R59288 a_13458_32299.n2 a_13458_32299.t0 24.9236
R59289 a_1412_46794.n11 a_1412_46794.t1 427.791
R59290 a_1412_46794.n8 a_1412_46794.t10 414.432
R59291 a_1412_46794.n8 a_1412_46794.t9 300.349
R59292 a_1412_46794.n2 a_1412_46794.t5 268.135
R59293 a_1412_46794.n0 a_1412_46794.t6 256.07
R59294 a_1412_46794.n3 a_1412_46794.t4 221.72
R59295 a_1412_46794.t0 a_1412_46794.n11 209.923
R59296 a_1412_46794.n5 a_1412_46794.t8 206.547
R59297 a_1412_46794.n1 a_1412_46794.t11 196.549
R59298 a_1412_46794.n10 a_1412_46794.n0 191.082
R59299 a_1412_46794.n7 a_1412_46794.n1 177.958
R59300 a_1412_46794.n6 a_1412_46794.n2 175.041
R59301 a_1412_46794.n6 a_1412_46794.n5 152
R59302 a_1412_46794.n0 a_1412_46794.t3 150.03
R59303 a_1412_46794.n4 a_1412_46794.t2 149.421
R59304 a_1412_46794.n1 a_1412_46794.t7 148.35
R59305 a_1412_46794.n7 a_1412_46794.n6 47.2963
R59306 a_1412_46794.n3 a_1412_46794.n2 28.5635
R59307 a_1412_46794.n9 a_1412_46794.n8 27.3955
R59308 a_1412_46794.n11 a_1412_46794.n10 20.1181
R59309 a_1412_46794.n4 a_1412_46794.n3 17.8524
R59310 a_1412_46794.n5 a_1412_46794.n4 17.8524
R59311 a_1412_46794.n9 a_1412_46794.n7 3.95019
R59312 a_1412_46794.n10 a_1412_46794.n9 0.914477
R59313 a_1736_39587.n0 a_1736_39587.t6 440.495
R59314 a_1736_39587.n4 a_1736_39587.t2 239.103
R59315 a_1736_39587.n1 a_1736_39587.t3 230.576
R59316 a_1736_39587.n0 a_1736_39587.t5 191.952
R59317 a_1736_39587.n2 a_1736_39587.n1 174.163
R59318 a_1736_39587.n1 a_1736_39587.t4 158.275
R59319 a_1736_39587.n3 a_1736_39587.t1 85.1701
R59320 a_1736_39587.t0 a_1736_39587.n4 61.169
R59321 a_1736_39587.n2 a_1736_39587.n0 5.84425
R59322 a_1736_39587.n3 a_1736_39587.n2 4.5005
R59323 a_1736_39587.n4 a_1736_39587.n3 2.04495
R59324 DATA[0].n5 DATA[0].n4 647.148
R59325 DATA[0].n2 DATA[0].n0 243.627
R59326 DATA[0].n2 DATA[0].n1 200.262
R59327 DATA[0].n5 DATA[0].n3 194.441
R59328 DATA[0].n6 DATA[0].n5 42.8458
R59329 DATA[0].n0 DATA[0].t2 40.0005
R59330 DATA[0].n0 DATA[0].t0 40.0005
R59331 DATA[0].n1 DATA[0].t1 40.0005
R59332 DATA[0].n1 DATA[0].t3 40.0005
R59333 DATA[0].n3 DATA[0].t4 27.5805
R59334 DATA[0].n3 DATA[0].t5 27.5805
R59335 DATA[0].n4 DATA[0].t7 27.5805
R59336 DATA[0].n4 DATA[0].t6 27.5805
R59337 DATA[0] DATA[0].n6 14.7904
R59338 DATA[0].n6 DATA[0].n2 7.72512
R59339 a_13878_32299.n1 a_13878_32299.t4 686.933
R59340 a_13878_32299.n1 a_13878_32299.n0 287.752
R59341 a_13878_32299.n2 a_13878_32299.n1 277.568
R59342 a_13878_32299.n0 a_13878_32299.t3 26.5955
R59343 a_13878_32299.n0 a_13878_32299.t2 26.5955
R59344 a_13878_32299.n2 a_13878_32299.t0 24.9236
R59345 a_13878_32299.t1 a_13878_32299.n2 24.9236
R59346 a_5542_30651.n3 a_5542_30651.t4 444.502
R59347 a_5542_30651.n2 a_5542_30651.t6 444.502
R59348 a_5542_30651.n6 a_5542_30651.n0 380.32
R59349 a_5542_30651.n3 a_5542_30651.t9 356.68
R59350 a_5542_30651.n2 a_5542_30651.t5 356.68
R59351 a_5542_30651.n1 a_5542_30651.t8 260.322
R59352 a_5542_30651.n4 a_5542_30651.n2 202.673
R59353 a_5542_30651.n4 a_5542_30651.n3 197.893
R59354 a_5542_30651.n7 a_5542_30651.n6 185
R59355 a_5542_30651.n1 a_5542_30651.t7 175.169
R59356 a_5542_30651.n5 a_5542_30651.n1 171.319
R59357 a_5542_30651.n5 a_5542_30651.n4 141.487
R59358 a_5542_30651.n0 a_5542_30651.t3 26.5955
R59359 a_5542_30651.n0 a_5542_30651.t2 26.5955
R59360 a_5542_30651.n7 a_5542_30651.t0 24.9236
R59361 a_5542_30651.t1 a_5542_30651.n7 24.9236
R59362 a_5542_30651.n6 a_5542_30651.n5 21.2067
R59363 a_1651_47044.n1 a_1651_47044.t1 457.955
R59364 a_1651_47044.n1 a_1651_47044.n0 288.253
R59365 a_1651_47044.n0 a_1651_47044.t3 239.505
R59366 a_1651_47044.t0 a_1651_47044.n1 216.155
R59367 a_1651_47044.n0 a_1651_47044.t2 167.204
R59368 a_n2103_43780.n8 a_n2103_43780.n7 300.118
R59369 a_n2103_43780.n5 a_n2103_43780.n4 299.834
R59370 a_n2103_43780.n10 a_n2103_43780.n9 299.834
R59371 a_n2103_43780.n8 a_n2103_43780.n6 291.81
R59372 a_n2103_43780.n3 a_n2103_43780.n0 283.969
R59373 a_n2103_43780.n0 a_n2103_43780.t11 276.464
R59374 a_n2103_43780.n3 a_n2103_43780.n2 251.452
R59375 a_n2103_43780.n2 a_n2103_43780.t8 212.081
R59376 a_n2103_43780.n1 a_n2103_43780.t10 212.081
R59377 a_n2103_43780.n0 a_n2103_43780.t13 196.131
R59378 a_n2103_43780.n2 a_n2103_43780.t9 139.78
R59379 a_n2103_43780.n1 a_n2103_43780.t12 139.78
R59380 a_n2103_43780.n9 a_n2103_43780.n8 79.8031
R59381 a_n2103_43780.n2 a_n2103_43780.n1 61.346
R59382 a_n2103_43780.n9 a_n2103_43780.n5 29.6732
R59383 a_n2103_43780.n7 a_n2103_43780.t6 26.5955
R59384 a_n2103_43780.n7 a_n2103_43780.t7 26.5955
R59385 a_n2103_43780.n4 a_n2103_43780.t2 26.5955
R59386 a_n2103_43780.n4 a_n2103_43780.t3 26.5955
R59387 a_n2103_43780.n10 a_n2103_43780.t0 26.5955
R59388 a_n2103_43780.t1 a_n2103_43780.n10 26.5955
R59389 a_n2103_43780.n6 a_n2103_43780.t4 24.9236
R59390 a_n2103_43780.n6 a_n2103_43780.t5 24.9236
R59391 a_n2103_43780.n5 a_n2103_43780.n3 14.7702
R59392 DATA[2].n3 DATA[2].n2 647.148
R59393 DATA[2].n5 DATA[2].n4 200.262
R59394 DATA[2].n3 DATA[2].n1 194.441
R59395 DATA[2].n6 DATA[2].n0 185
R59396 DATA[2].n6 DATA[2].n5 58.6278
R59397 DATA[2].n5 DATA[2].n3 50.5705
R59398 DATA[2].n0 DATA[2].t0 40.0005
R59399 DATA[2].n0 DATA[2].t3 40.0005
R59400 DATA[2].n4 DATA[2].t1 40.0005
R59401 DATA[2].n4 DATA[2].t2 40.0005
R59402 DATA[2].n1 DATA[2].t4 27.5805
R59403 DATA[2].n1 DATA[2].t7 27.5805
R59404 DATA[2].n2 DATA[2].t6 27.5805
R59405 DATA[2].n2 DATA[2].t5 27.5805
R59406 DATA[2] DATA[2].n6 15.6247
R59407 CLK.n0 CLK.t0 260.322
R59408 CLK.n0 CLK.t1 175.169
R59409 CLK CLK.n0 169.487
R59410 a_n2661_47044.n5 a_n2661_47044.n0 664.928
R59411 a_n2661_47044.n1 a_n2661_47044.t6 276.464
R59412 a_n2661_47044.n4 a_n2661_47044.n1 256.538
R59413 a_n2661_47044.n4 a_n2661_47044.n3 218.405
R59414 a_n2661_47044.n2 a_n2661_47044.t9 212.081
R59415 a_n2661_47044.n3 a_n2661_47044.t8 212.081
R59416 a_n2661_47044.n1 a_n2661_47044.t7 196.131
R59417 a_n2661_47044.n6 a_n2661_47044.n5 187.927
R59418 a_n2661_47044.n2 a_n2661_47044.t4 139.78
R59419 a_n2661_47044.n3 a_n2661_47044.t5 139.78
R59420 a_n2661_47044.n3 a_n2661_47044.n2 61.346
R59421 a_n2661_47044.n0 a_n2661_47044.t2 26.5955
R59422 a_n2661_47044.n0 a_n2661_47044.t3 26.5955
R59423 a_n2661_47044.t1 a_n2661_47044.n6 24.9236
R59424 a_n2661_47044.n6 a_n2661_47044.t0 24.9236
R59425 a_n2661_47044.n5 a_n2661_47044.n4 14.0946
R59426 a_n2442_45982.n1 a_n2442_45982.t4 595.52
R59427 a_n2442_45982.n1 a_n2442_45982.n0 380.32
R59428 a_n2442_45982.n2 a_n2442_45982.n1 185
R59429 a_n2442_45982.n0 a_n2442_45982.t2 26.5955
R59430 a_n2442_45982.n0 a_n2442_45982.t3 26.5955
R59431 a_n2442_45982.n2 a_n2442_45982.t0 24.9236
R59432 a_n2442_45982.t1 a_n2442_45982.n2 24.9236
R59433 a_n2810_43262.n1 a_n2810_43262.t4 677.35
R59434 a_n2810_43262.n1 a_n2810_43262.n0 380.32
R59435 a_n2810_43262.n2 a_n2810_43262.n1 185
R59436 a_n2810_43262.n0 a_n2810_43262.t3 26.5955
R59437 a_n2810_43262.n0 a_n2810_43262.t2 26.5955
R59438 a_n2810_43262.n2 a_n2810_43262.t0 24.9236
R59439 a_n2810_43262.t1 a_n2810_43262.n2 24.9236
R59440 a_14409_32299.n1 a_14409_32299.t4 738.654
R59441 a_14409_32299.n1 a_14409_32299.n0 380.32
R59442 a_14409_32299.n2 a_14409_32299.n1 185
R59443 a_14409_32299.n0 a_14409_32299.t3 26.5955
R59444 a_14409_32299.n0 a_14409_32299.t2 26.5955
R59445 a_14409_32299.t1 a_14409_32299.n2 24.9236
R59446 a_14409_32299.n2 a_14409_32299.t0 24.9236
R59447 C2_P_btm.n1 C2_P_btm.t0 101.621
R59448 C2_P_btm.n2 C2_P_btm.t2 98.936
R59449 C2_P_btm.n0 C2_P_btm.t3 54.9311
R59450 C2_P_btm C2_P_btm.n2 52.0317
R59451 C2_P_btm.n0 C2_P_btm.t1 47.3635
R59452 C2_P_btm C2_P_btm.n6 8.338
R59453 C2_P_btm.n1 C2_P_btm.n0 7.71404
R59454 C2_P_btm.n2 C2_P_btm.n1 7.20883
R59455 C2_P_btm.n3 C2_P_btm.t5 4.76819
R59456 C2_P_btm.n5 C2_P_btm.t6 4.03712
R59457 C2_P_btm.n6 C2_P_btm.t4 4.03712
R59458 C2_P_btm.n4 C2_P_btm.t8 3.98193
R59459 C2_P_btm.n3 C2_P_btm.t7 3.92851
R59460 C2_P_btm.n5 C2_P_btm.n4 1.05569
R59461 C2_P_btm.n6 C2_P_btm.n5 1.0005
R59462 C2_P_btm.n4 C2_P_btm.n3 0.786757
R59463 a_n2103_44324.n5 a_n2103_44324.n0 664.928
R59464 a_n2103_44324.n1 a_n2103_44324.t7 276.464
R59465 a_n2103_44324.n4 a_n2103_44324.n3 224.893
R59466 a_n2103_44324.n3 a_n2103_44324.t8 212.081
R59467 a_n2103_44324.n2 a_n2103_44324.t6 212.081
R59468 a_n2103_44324.n1 a_n2103_44324.t4 196.131
R59469 a_n2103_44324.n4 a_n2103_44324.n1 195.061
R59470 a_n2103_44324.n6 a_n2103_44324.n5 187.927
R59471 a_n2103_44324.n3 a_n2103_44324.t9 139.78
R59472 a_n2103_44324.n2 a_n2103_44324.t5 139.78
R59473 a_n2103_44324.n3 a_n2103_44324.n2 61.346
R59474 a_n2103_44324.n0 a_n2103_44324.t3 26.5955
R59475 a_n2103_44324.n0 a_n2103_44324.t2 26.5955
R59476 a_n2103_44324.t1 a_n2103_44324.n6 24.9236
R59477 a_n2103_44324.n6 a_n2103_44324.t0 24.9236
R59478 a_n2103_44324.n5 a_n2103_44324.n4 9.3005
R59479 a_n2810_45982.n1 a_n2810_45982.t4 597.014
R59480 a_n2810_45982.n1 a_n2810_45982.n0 296.139
R59481 a_n2810_45982.n2 a_n2810_45982.n1 269.182
R59482 a_n2810_45982.n0 a_n2810_45982.t3 26.5955
R59483 a_n2810_45982.n0 a_n2810_45982.t2 26.5955
R59484 a_n2810_45982.t1 a_n2810_45982.n2 24.9236
R59485 a_n2810_45982.n2 a_n2810_45982.t0 24.9236
R59486 a_n2442_46526.n1 a_n2442_46526.t4 606.707
R59487 a_n2442_46526.n1 a_n2442_46526.n0 287.752
R59488 a_n2442_46526.n2 a_n2442_46526.n1 277.568
R59489 a_n2442_46526.n0 a_n2442_46526.t2 26.5955
R59490 a_n2442_46526.n0 a_n2442_46526.t3 26.5955
R59491 a_n2442_46526.n2 a_n2442_46526.t0 24.9236
R59492 a_n2442_46526.t1 a_n2442_46526.n2 24.9236
R59493 a_n1890_47614.n1 a_n1890_47614.t5 756.514
R59494 a_n1890_47614.n1 a_n1890_47614.t4 756.239
R59495 a_n1890_47614.n2 a_n1890_47614.n0 287.752
R59496 a_n1890_47614.n3 a_n1890_47614.n2 277.568
R59497 a_n1890_47614.n2 a_n1890_47614.n1 122.615
R59498 a_n1890_47614.n0 a_n1890_47614.t3 26.5955
R59499 a_n1890_47614.n0 a_n1890_47614.t2 26.5955
R59500 a_n1890_47614.t1 a_n1890_47614.n3 24.9236
R59501 a_n1890_47614.n3 a_n1890_47614.t0 24.9236
R59502 a_n1435_47614.n1 a_n1435_47614.t1 366.548
R59503 a_n1435_47614.t0 a_n1435_47614.n1 310.909
R59504 a_n1435_47614.n0 a_n1435_47614.t3 241.536
R59505 a_n1435_47614.n1 a_n1435_47614.n0 240.081
R59506 a_n1435_47614.n0 a_n1435_47614.t2 169.237
R59507 a_4338_37500.t0 a_4338_37500.n4 258.05
R59508 a_4338_37500.n4 a_4338_37500.n3 53.4434
R59509 a_4338_37500.n1 a_4338_37500.t4 47.8126
R59510 a_4338_37500.n2 a_4338_37500.t1 47.5157
R59511 a_4338_37500.n1 a_4338_37500.n0 37.6157
R59512 a_4338_37500.n3 a_4338_37500.t5 10.4216
R59513 a_4338_37500.n3 a_4338_37500.t6 10.4216
R59514 a_4338_37500.n0 a_4338_37500.t2 9.9005
R59515 a_4338_37500.n0 a_4338_37500.t3 9.9005
R59516 a_4338_37500.n4 a_4338_37500.n2 2.8755
R59517 a_4338_37500.n2 a_4338_37500.n1 0.313
R59518 DEBUG_OUT.n5 DEBUG_OUT.n4 647.148
R59519 DEBUG_OUT.n2 DEBUG_OUT.n0 243.627
R59520 DEBUG_OUT.n2 DEBUG_OUT.n1 200.262
R59521 DEBUG_OUT.n5 DEBUG_OUT.n3 194.441
R59522 DEBUG_OUT.n6 DEBUG_OUT.n5 42.8458
R59523 DEBUG_OUT.n0 DEBUG_OUT.t1 40.0005
R59524 DEBUG_OUT.n0 DEBUG_OUT.t0 40.0005
R59525 DEBUG_OUT.n1 DEBUG_OUT.t3 40.0005
R59526 DEBUG_OUT.n1 DEBUG_OUT.t2 40.0005
R59527 DEBUG_OUT.n3 DEBUG_OUT.t7 27.5805
R59528 DEBUG_OUT.n3 DEBUG_OUT.t4 27.5805
R59529 DEBUG_OUT.n4 DEBUG_OUT.t6 27.5805
R59530 DEBUG_OUT.n4 DEBUG_OUT.t5 27.5805
R59531 DEBUG_OUT DEBUG_OUT.n6 17.1381
R59532 DEBUG_OUT.n6 DEBUG_OUT.n2 7.72512
R59533 a_2252_42718.n2 a_2252_42718.t7 580.423
R59534 a_2252_42718.n2 a_2252_42718.t4 580.144
R59535 a_2252_42718.n4 a_2252_42718.n0 380.32
R59536 a_2252_42718.n1 a_2252_42718.t5 260.322
R59537 a_2252_42718.n5 a_2252_42718.n4 185
R59538 a_2252_42718.n3 a_2252_42718.n1 176.272
R59539 a_2252_42718.n1 a_2252_42718.t6 175.169
R59540 a_2252_42718.n3 a_2252_42718.n2 123.112
R59541 a_2252_42718.n0 a_2252_42718.t2 26.5955
R59542 a_2252_42718.n0 a_2252_42718.t3 26.5955
R59543 a_2252_42718.t1 a_2252_42718.n5 24.9236
R59544 a_2252_42718.n5 a_2252_42718.t0 24.9236
R59545 a_2252_42718.n4 a_2252_42718.n3 22.2424
R59546 a_19921_31459.n1 a_19921_31459.t4 594.867
R59547 a_19921_31459.n1 a_19921_31459.n0 380.32
R59548 a_19921_31459.n2 a_19921_31459.n1 185
R59549 a_19921_31459.n0 a_19921_31459.t3 26.5955
R59550 a_19921_31459.n0 a_19921_31459.t2 26.5955
R59551 a_19921_31459.t1 a_19921_31459.n2 24.9236
R59552 a_19921_31459.n2 a_19921_31459.t0 24.9236
R59553 DEBUG_MUX[1].n0 DEBUG_MUX[1].t0 224.984
R59554 DEBUG_MUX[1].n0 DEBUG_MUX[1].t1 187.714
R59555 DEBUG_MUX[1] DEBUG_MUX[1].n0 180.094
R59556 a_n2442_45438.n1 a_n2442_45438.t4 608.11
R59557 a_n2442_45438.n1 a_n2442_45438.n0 287.752
R59558 a_n2442_45438.n2 a_n2442_45438.n1 277.568
R59559 a_n2442_45438.n0 a_n2442_45438.t2 26.5955
R59560 a_n2442_45438.n0 a_n2442_45438.t3 26.5955
R59561 a_n2442_45438.n2 a_n2442_45438.t0 24.9236
R59562 a_n2442_45438.t1 a_n2442_45438.n2 24.9236
R59563 w_11534_34010.n51 w_11534_34010.n10 27635.6
R59564 w_11534_34010.n50 w_11534_34010.n9 14784.7
R59565 w_11534_34010.n53 w_11534_34010.n9 14784.7
R59566 w_11534_34010.n53 w_11534_34010.n8 14784.7
R59567 w_11534_34010.n17 w_11534_34010.n8 11195.3
R59568 w_11534_34010.n28 w_11534_34010.n20 3017.65
R59569 w_11534_34010.n28 w_11534_34010.n19 3017.65
R59570 w_11534_34010.n30 w_11534_34010.n19 3017.65
R59571 w_11534_34010.n16 w_11534_34010.n15 1757.65
R59572 w_11534_34010.n17 w_11534_34010.n11 1757.65
R59573 w_11534_34010.n50 w_11534_34010.n11 1711.76
R59574 w_11534_34010.n54 w_11534_34010.n7 1577.04
R59575 w_11534_34010.n55 w_11534_34010.n6 1373.85
R59576 w_11534_34010.n30 w_11534_34010.n16 1080
R59577 w_11534_34010.n49 w_11534_34010.n48 936.562
R59578 w_11534_34010.t8 w_11534_34010.n34 905.04
R59579 w_11534_34010.n35 w_11534_34010.t8 812.54
R59580 w_11534_34010.n53 w_11534_34010.t10 724.569
R59581 w_11534_34010.t13 w_11534_34010.n51 717.962
R59582 w_11534_34010.n52 w_11534_34010.t13 668.146
R59583 w_11534_34010.t10 w_11534_34010.n52 668.146
R59584 w_11534_34010.n13 w_11534_34010.n12 621.929
R59585 w_11534_34010.n12 w_11534_34010.n6 572.236
R59586 w_11534_34010.n34 w_11534_34010.n16 557.648
R59587 w_11534_34010.n34 w_11534_34010.n17 557.648
R59588 w_11534_34010.n36 w_11534_34010.n15 557.648
R59589 w_11534_34010.n36 w_11534_34010.n11 557.648
R59590 w_11534_34010.n48 w_11534_34010.n7 497.269
R59591 w_11534_34010.n27 w_11534_34010.n26 298.877
R59592 w_11534_34010.n23 w_11534_34010.n18 280.202
R59593 w_11534_34010.n25 w_11534_34010.n24 277.776
R59594 w_11534_34010.n39 w_11534_34010.t9 228.215
R59595 w_11534_34010.n55 w_11534_34010.n54 195.883
R59596 w_11534_34010.n47 w_11534_34010.n13 187.482
R59597 w_11534_34010.n32 w_11534_34010.n14 187.482
R59598 w_11534_34010.n49 w_11534_34010.n47 182.589
R59599 w_11534_34010.t0 w_11534_34010.n19 137.529
R59600 w_11534_34010.n32 w_11534_34010.n31 115.201
R59601 w_11534_34010.n35 w_11534_34010.n10 103.859
R59602 w_11534_34010.n37 w_11534_34010.n36 92.5005
R59603 w_11534_34010.n36 w_11534_34010.n35 92.5005
R59604 w_11534_34010.n34 w_11534_34010.n33 92.5005
R59605 w_11534_34010.t6 w_11534_34010.n10 75.2024
R59606 w_11534_34010.t4 w_11534_34010.t0 73.6677
R59607 w_11534_34010.t2 w_11534_34010.t6 73.6677
R59608 w_11534_34010.n68 w_11534_34010.t1 65.4041
R59609 w_11534_34010.n66 w_11534_34010.t7 62.5643
R59610 w_11534_34010.n5 w_11534_34010.t17 61.7296
R59611 w_11534_34010.n44 w_11534_34010.t14 61.7296
R59612 w_11534_34010.n59 w_11534_34010.t12 61.7296
R59613 w_11534_34010.n62 w_11534_34010.t15 61.7296
R59614 w_11534_34010.n20 w_11534_34010.n15 60.0005
R59615 w_11534_34010.n37 w_11534_34010.n14 59.4829
R59616 w_11534_34010.n47 w_11534_34010.n37 59.4829
R59617 w_11534_34010.n33 w_11534_34010.n32 59.4829
R59618 w_11534_34010.n33 w_11534_34010.n13 59.4829
R59619 w_11534_34010.n69 w_11534_34010.n68 56.8163
R59620 w_11534_34010.n43 w_11534_34010.n42 54.1123
R59621 w_11534_34010.n61 w_11534_34010.n60 54.1123
R59622 w_11534_34010.n29 w_11534_34010.t4 36.8341
R59623 w_11534_34010.n29 w_11534_34010.t2 36.8341
R59624 w_11534_34010.n31 w_11534_34010.n30 26.4291
R59625 w_11534_34010.n30 w_11534_34010.n29 26.4291
R59626 w_11534_34010.n28 w_11534_34010.n27 26.4291
R59627 w_11534_34010.n29 w_11534_34010.n28 26.4291
R59628 w_11534_34010.n24 w_11534_34010.n23 20.4805
R59629 w_11534_34010.n31 w_11534_34010.n18 16.9417
R59630 w_11534_34010.n38 w_11534_34010.n2 15.2505
R59631 w_11534_34010.n26 w_11534_34010.n20 13.2148
R59632 w_11534_34010.n20 w_11534_34010.n10 13.2148
R59633 w_11534_34010.n24 w_11534_34010.n19 13.2148
R59634 w_11534_34010.n27 w_11534_34010.n25 8.2968
R59635 w_11534_34010.t5 w_11534_34010.n69 8.12675
R59636 w_11534_34010.n69 w_11534_34010.t3 8.12675
R59637 w_11534_34010.t14 w_11534_34010.n43 7.61783
R59638 w_11534_34010.n43 w_11534_34010.t16 7.61783
R59639 w_11534_34010.t15 w_11534_34010.n61 7.61783
R59640 w_11534_34010.n61 w_11534_34010.t11 7.61783
R59641 w_11534_34010.n54 w_11534_34010.n53 6.60764
R59642 w_11534_34010.n50 w_11534_34010.n49 6.60764
R59643 w_11534_34010.n51 w_11534_34010.n50 6.60764
R59644 w_11534_34010.n58 w_11534_34010.n3 6.41545
R59645 w_11534_34010.n26 w_11534_34010.n14 6.4005
R59646 w_11534_34010.n57 w_11534_34010.n4 6.37679
R59647 w_11534_34010.n68 w_11534_34010.n67 2.72081
R59648 w_11534_34010.n63 w_11534_34010.n3 2.50761
R59649 w_11534_34010.n40 w_11534_34010.n4 2.12421
R59650 w_11534_34010.n9 w_11534_34010.n7 2.03347
R59651 w_11534_34010.n52 w_11534_34010.n9 2.03347
R59652 w_11534_34010.n8 w_11534_34010.n6 2.03347
R59653 w_11534_34010.n52 w_11534_34010.n8 2.03347
R59654 w_11534_34010.n25 w_11534_34010.n1 1.5505
R59655 w_11534_34010.n21 w_11534_34010.n18 1.5505
R59656 w_11534_34010.n22 w_11534_34010.n1 1.26012
R59657 w_11534_34010.n23 w_11534_34010.n22 1.03383
R59658 w_11534_34010.n47 w_11534_34010.n46 1.03383
R59659 w_11534_34010.n56 w_11534_34010.n55 1.03383
R59660 w_11534_34010.n66 w_11534_34010.n65 1.00774
R59661 w_11534_34010.n22 w_11534_34010.n21 0.937356
R59662 w_11534_34010.n62 w_11534_34010.n60 0.891526
R59663 w_11534_34010.n60 w_11534_34010.n59 0.891526
R59664 w_11534_34010.n44 w_11534_34010.n42 0.891526
R59665 w_11534_34010.n42 w_11534_34010.n5 0.891526
R59666 w_11534_34010.n58 w_11534_34010.n57 0.741479
R59667 w_11534_34010.n65 w_11534_34010.n1 0.543562
R59668 w_11534_34010.n40 w_11534_34010.n0 0.494823
R59669 w_11534_34010.n21 w_11534_34010.n0 0.44251
R59670 w_11534_34010.n67 w_11534_34010.n0 0.428803
R59671 w_11534_34010.n64 w_11534_34010.n2 0.286876
R59672 w_11534_34010.n64 w_11534_34010.n63 0.260999
R59673 w_11534_34010.n41 w_11534_34010.n40 0.253077
R59674 w_11534_34010.n48 w_11534_34010.n3 0.227329
R59675 w_11534_34010.n12 w_11534_34010.n4 0.227329
R59676 w_11534_34010.n65 w_11534_34010.n64 0.192353
R59677 w_11534_34010.n45 w_11534_34010.n2 0.178335
R59678 w_11534_34010.n39 w_11534_34010.n38 0.0711522
R59679 w_11534_34010.n45 w_11534_34010.n41 0.0700876
R59680 w_11534_34010.n67 w_11534_34010.n66 0.057539
R59681 w_11534_34010.n59 w_11534_34010.n58 0.035465
R59682 w_11534_34010.n56 w_11534_34010.n5 0.0340082
R59683 w_11534_34010.n63 w_11534_34010.n62 0.0330567
R59684 w_11534_34010.n45 w_11534_34010.n44 0.0325513
R59685 w_11534_34010.n41 w_11534_34010.n39 0.0303913
R59686 w_11534_34010.n46 w_11534_34010.n38 0.0136119
R59687 w_11534_34010.n57 w_11534_34010.n56 0.00195688
R59688 w_11534_34010.n46 w_11534_34010.n45 0.0016655
R59689 DEBUG_MUX[0].n0 DEBUG_MUX[0].t1 224.984
R59690 DEBUG_MUX[0].n0 DEBUG_MUX[0].t0 187.714
R59691 DEBUG_MUX[0] DEBUG_MUX[0].n0 178.951
R59692 a_6104_45706.n11 a_6104_45706.t1 427.791
R59693 a_6104_45706.n7 a_6104_45706.t11 414.432
R59694 a_6104_45706.n7 a_6104_45706.t5 300.349
R59695 a_6104_45706.n1 a_6104_45706.t4 268.135
R59696 a_6104_45706.n8 a_6104_45706.t3 256.07
R59697 a_6104_45706.n2 a_6104_45706.t7 221.72
R59698 a_6104_45706.t0 a_6104_45706.n11 209.923
R59699 a_6104_45706.n4 a_6104_45706.t2 206.547
R59700 a_6104_45706.n0 a_6104_45706.t6 196.549
R59701 a_6104_45706.n9 a_6104_45706.n8 181.852
R59702 a_6104_45706.n5 a_6104_45706.n1 175.041
R59703 a_6104_45706.n6 a_6104_45706.n0 172.947
R59704 a_6104_45706.n5 a_6104_45706.n4 152
R59705 a_6104_45706.n8 a_6104_45706.t8 150.03
R59706 a_6104_45706.n3 a_6104_45706.t9 149.421
R59707 a_6104_45706.n0 a_6104_45706.t10 148.35
R59708 a_6104_45706.n6 a_6104_45706.n5 47.0546
R59709 a_6104_45706.n9 a_6104_45706.n7 33.4218
R59710 a_6104_45706.n2 a_6104_45706.n1 28.5635
R59711 a_6104_45706.n11 a_6104_45706.n10 19.824
R59712 a_6104_45706.n3 a_6104_45706.n2 17.8524
R59713 a_6104_45706.n4 a_6104_45706.n3 17.8524
R59714 a_6104_45706.n10 a_6104_45706.n9 5.45754
R59715 a_6104_45706.n10 a_6104_45706.n6 3.20792
R59716 CAL_N.n6 CAL_N.n5 600.547
R59717 CAL_N.n6 CAL_N.t1 260.075
R59718 CAL_N CAL_N.t3 138.526
R59719 CAL_N.n5 CAL_N.t0 77.3934
R59720 CAL_N.n5 CAL_N.t2 77.3934
R59721 CAL_N.n1 CAL_N.t4 36.3712
R59722 CAL_N.n2 CAL_N.t4 36.3712
R59723 CAL_N.n3 CAL_N.t5 36.2721
R59724 CAL_N.t5 CAL_N.n0 36.2721
R59725 CAL_N.n2 CAL_N.t6 31.2287
R59726 CAL_N.t6 CAL_N.n1 31.2287
R59727 CAL_N CAL_N.n7 29.3678
R59728 CAL_N.n7 CAL_N.n6 10.1411
R59729 CAL_N.n4 CAL_N.n0 8.938
R59730 CAL_N.n4 CAL_N.n3 4.5005
R59731 CAL_N.n1 CAL_N.n0 0.0713333
R59732 CAL_N.n3 CAL_N.n2 0.0713333
R59733 CAL_N.n7 CAL_N.n4 0.0213333
R59734 a_4758_30651.n7 a_4758_30651.t11 1421.83
R59735 a_4758_30651.n1 a_4758_30651.t9 1421.83
R59736 a_4758_30651.n6 a_4758_30651.t4 1327.11
R59737 a_4758_30651.n2 a_4758_30651.t7 1327.11
R59738 a_4758_30651.n7 a_4758_30651.t13 1320.68
R59739 a_4758_30651.n5 a_4758_30651.t6 1320.68
R59740 a_4758_30651.n3 a_4758_30651.t10 1320.68
R59741 a_4758_30651.n1 a_4758_30651.t8 1320.68
R59742 a_4758_30651.n12 a_4758_30651.n0 380.32
R59743 a_4758_30651.n10 a_4758_30651.t5 260.322
R59744 a_4758_30651.n13 a_4758_30651.n12 185
R59745 a_4758_30651.n10 a_4758_30651.t12 175.169
R59746 a_4758_30651.n11 a_4758_30651.n10 173.97
R59747 a_4758_30651.n8 a_4758_30651.n5 161.698
R59748 a_4758_30651.n4 a_4758_30651.n3 161.698
R59749 a_4758_30651.n8 a_4758_30651.n7 161.303
R59750 a_4758_30651.n4 a_4758_30651.n1 161.303
R59751 a_4758_30651.n6 a_4758_30651.n5 94.7191
R59752 a_4758_30651.n7 a_4758_30651.n6 94.7191
R59753 a_4758_30651.n2 a_4758_30651.n1 94.7191
R59754 a_4758_30651.n3 a_4758_30651.n2 94.7191
R59755 a_4758_30651.n11 a_4758_30651.n9 84.88
R59756 a_4758_30651.n9 a_4758_30651.n8 35.787
R59757 a_4758_30651.n9 a_4758_30651.n4 33.0661
R59758 a_4758_30651.n0 a_4758_30651.t3 26.5955
R59759 a_4758_30651.n0 a_4758_30651.t2 26.5955
R59760 a_4758_30651.t1 a_4758_30651.n13 24.9236
R59761 a_4758_30651.n13 a_4758_30651.t0 24.9236
R59762 a_4758_30651.n12 a_4758_30651.n11 16.8764
R59763 a_11730_34132.n17 a_11730_34132.n16 21.0497
R59764 a_11730_34132.n16 a_11730_34132.n15 20.1816
R59765 a_11730_34132.t6 a_11730_34132.n1 10.7351
R59766 a_11730_34132.n12 a_11730_34132.t6 10.7351
R59767 a_11730_34132.t4 a_11730_34132.n5 10.7351
R59768 a_11730_34132.n6 a_11730_34132.t4 10.7351
R59769 a_11730_34132.n5 a_11730_34132.t7 10.7351
R59770 a_11730_34132.t7 a_11730_34132.n3 10.7351
R59771 a_11730_34132.n12 a_11730_34132.t5 10.7351
R59772 a_11730_34132.t5 a_11730_34132.n0 10.7351
R59773 a_11730_34132.n16 a_11730_34132.n14 8.273
R59774 a_11730_34132.n13 a_11730_34132.n1 6.92882
R59775 a_11730_34132.n14 a_11730_34132.n0 6.39
R59776 a_11730_34132.n10 a_11730_34132.n1 5.96919
R59777 a_11730_34132.n7 a_11730_34132.n6 5.82288
R59778 a_11730_34132.n6 a_11730_34132.n4 5.7297
R59779 a_11730_34132.n4 a_11730_34132.n3 5.57478
R59780 a_11730_34132.n15 a_11730_34132.t2 4.9505
R59781 a_11730_34132.n15 a_11730_34132.t3 4.9505
R59782 a_11730_34132.n17 a_11730_34132.t0 4.9505
R59783 a_11730_34132.t1 a_11730_34132.n17 4.9505
R59784 a_11730_34132.n13 a_11730_34132.n12 3.29339
R59785 a_11730_34132.n8 a_11730_34132.n7 3.27354
R59786 a_11730_34132.n10 a_11730_34132.n9 3.26815
R59787 a_11730_34132.n9 a_11730_34132.n8 3.08438
R59788 a_11730_34132.n5 a_11730_34132.n4 2.93843
R59789 a_11730_34132.n9 a_11730_34132.n0 2.59618
R59790 a_11730_34132.n8 a_11730_34132.n3 2.38498
R59791 a_11730_34132.n7 a_11730_34132.n2 2.24345
R59792 a_11730_34132.n11 a_11730_34132.n10 2.23748
R59793 a_11730_34132.n11 a_11730_34132.n2 1.16457
R59794 a_11730_34132.n12 a_11730_34132.n11 0.786485
R59795 a_11730_34132.n5 a_11730_34132.n2 0.739126
R59796 a_11730_34132.n14 a_11730_34132.n13 0.34925
R59797 a_n2810_45438.n1 a_n2810_45438.t4 597.876
R59798 a_n2810_45438.n1 a_n2810_45438.n0 380.32
R59799 a_n2810_45438.n2 a_n2810_45438.n1 185
R59800 a_n2810_45438.n0 a_n2810_45438.t3 26.5955
R59801 a_n2810_45438.n0 a_n2810_45438.t2 26.5955
R59802 a_n2810_45438.t1 a_n2810_45438.n2 24.9236
R59803 a_n2810_45438.n2 a_n2810_45438.t0 24.9236
R59804 DATA[1].n5 DATA[1].n4 647.148
R59805 DATA[1].n2 DATA[1].n0 243.627
R59806 DATA[1].n2 DATA[1].n1 200.262
R59807 DATA[1].n5 DATA[1].n3 194.441
R59808 DATA[1].n6 DATA[1].n5 42.8458
R59809 DATA[1].n0 DATA[1].t2 40.0005
R59810 DATA[1].n0 DATA[1].t1 40.0005
R59811 DATA[1].n1 DATA[1].t0 40.0005
R59812 DATA[1].n1 DATA[1].t3 40.0005
R59813 DATA[1].n3 DATA[1].t6 27.5805
R59814 DATA[1].n3 DATA[1].t5 27.5805
R59815 DATA[1].n4 DATA[1].t4 27.5805
R59816 DATA[1].n4 DATA[1].t7 27.5805
R59817 DATA[1] DATA[1].n6 15.5175
R59818 DATA[1].n6 DATA[1].n2 7.72512
R59819 EN_OFFSET_CAL.n0 EN_OFFSET_CAL.t1 260.322
R59820 EN_OFFSET_CAL.n0 EN_OFFSET_CAL.t0 175.169
R59821 EN_OFFSET_CAL EN_OFFSET_CAL.n0 168.62
R59822 a_10199_47846.n1 a_10199_47846.t1 381.774
R59823 a_10199_47846.n0 a_10199_47846.t3 238.59
R59824 a_10199_47846.n1 a_10199_47846.n0 206.989
R59825 a_10199_47846.n0 a_10199_47846.t2 203.244
R59826 a_10199_47846.t0 a_10199_47846.n1 185.649
R59827 a_n2074_43262.n1 a_n2074_43262.t4 685.83
R59828 a_n2074_43262.n1 a_n2074_43262.n0 287.752
R59829 a_n2074_43262.n2 a_n2074_43262.n1 277.568
R59830 a_n2074_43262.n0 a_n2074_43262.t2 26.5955
R59831 a_n2074_43262.n0 a_n2074_43262.t3 26.5955
R59832 a_n2074_43262.n2 a_n2074_43262.t0 24.9236
R59833 a_n2074_43262.t1 a_n2074_43262.n2 24.9236
R59834 a_n2109_42692.t0 a_n2109_42692.n3 392.767
R59835 a_n2109_42692.n1 a_n2109_42692.t5 276.464
R59836 a_n2109_42692.n2 a_n2109_42692.n1 212.656
R59837 a_n2109_42692.n2 a_n2109_42692.t1 209.923
R59838 a_n2109_42692.n1 a_n2109_42692.t4 196.131
R59839 a_n2109_42692.n3 a_n2109_42692.n0 192.906
R59840 a_n2109_42692.n3 a_n2109_42692.n2 66.3848
R59841 a_n2109_42692.n0 a_n2109_42692.t2 24.9236
R59842 a_n2109_42692.n0 a_n2109_42692.t3 24.9236
R59843 START.n0 START.t0 260.322
R59844 START.n0 START.t1 175.169
R59845 START START.n0 168.62
R59846 a_n2074_47070.n1 a_n2074_47070.t4 599.491
R59847 a_n2074_47070.n1 a_n2074_47070.n0 380.32
R59848 a_n2074_47070.n2 a_n2074_47070.n1 185
R59849 a_n2074_47070.n0 a_n2074_47070.t2 26.5955
R59850 a_n2074_47070.n0 a_n2074_47070.t3 26.5955
R59851 a_n2074_47070.n2 a_n2074_47070.t0 24.9236
R59852 a_n2074_47070.t1 a_n2074_47070.n2 24.9236
R59853 a_19437_31459.n1 a_19437_31459.t4 604.801
R59854 a_19437_31459.n1 a_19437_31459.n0 287.752
R59855 a_19437_31459.n2 a_19437_31459.n1 277.568
R59856 a_19437_31459.n0 a_19437_31459.t2 26.5955
R59857 a_19437_31459.n0 a_19437_31459.t3 26.5955
R59858 a_19437_31459.t1 a_19437_31459.n2 24.9236
R59859 a_19437_31459.n2 a_19437_31459.t0 24.9236
R59860 a_14087_32299.n1 a_14087_32299.t4 684.321
R59861 a_14087_32299.n1 a_14087_32299.n0 287.752
R59862 a_14087_32299.n2 a_14087_32299.n1 277.568
R59863 a_14087_32299.n0 a_14087_32299.t2 26.5955
R59864 a_14087_32299.n0 a_14087_32299.t3 26.5955
R59865 a_14087_32299.n2 a_14087_32299.t0 24.9236
R59866 a_14087_32299.t1 a_14087_32299.n2 24.9236
R59867 C0_P_btm.n1 C0_P_btm.t0 101.944
R59868 C0_P_btm.n2 C0_P_btm.t1 99.4985
R59869 C0_P_btm.n0 C0_P_btm.t5 54.9098
R59870 C0_P_btm C0_P_btm.n2 49.2817
R59871 C0_P_btm.n0 C0_P_btm.t2 47.3635
R59872 C0_P_btm C0_P_btm.n3 8.6505
R59873 C0_P_btm.n1 C0_P_btm.n0 8.27654
R59874 C0_P_btm.n2 C0_P_btm.n1 6.33383
R59875 C0_P_btm.n3 C0_P_btm.t4 5.03712
R59876 C0_P_btm.n3 C0_P_btm.t3 4.03712
R59877 DEBUG_MUX[3].n0 DEBUG_MUX[3].t0 260.322
R59878 DEBUG_MUX[3].n0 DEBUG_MUX[3].t1 175.169
R59879 DEBUG_MUX[3] DEBUG_MUX[3].n0 169.877
R59880 a_n2442_43806.n1 a_n2442_43806.t4 742.208
R59881 a_n2442_43806.n1 a_n2442_43806.n0 380.32
R59882 a_n2442_43806.n2 a_n2442_43806.n1 185
R59883 a_n2442_43806.n0 a_n2442_43806.t2 26.5955
R59884 a_n2442_43806.n0 a_n2442_43806.t3 26.5955
R59885 a_n2442_43806.n2 a_n2442_43806.t0 24.9236
R59886 a_n2442_43806.t1 a_n2442_43806.n2 24.9236
C0 a_n685_43268# a_n169_43640# 0.105914f
C1 a_n519_43268# a_49_43236# 0.175891f
C2 a_3165_45982# a_3882_44324# 0.203371f
C3 a_10428_47338# a_10554_47436# 0.174625f
C4 a_10467_47212# a_10623_47307# 0.105766f
C5 a_15437_47044# a_15329_47044# 0.146948f
C6 a_n2288_47588# VDD 0.2896f
C7 a_4005_46500# VDD 0.205629f
C8 C5_N_btm VIN_N 0.502107f
C9 VDD DEBUG_OUT 0.391267f
C10 C3_N_btm VCM 0.716273f
C11 C4_N_btm VREF 0.98728f
C12 a_171_44019# VDD 0.467266f
C13 a_n1741_42692# a_n1920_42692# 0.176311f
C14 a_2043_43958# VDD 0.207559f
C15 a_13635_43566# VDD 0.453505f
C16 COMP_N a_1239_39043# 0.38801f
C17 a_5655_43780# a_6091_43780# 0.343552f
C18 a_14219_47070# VDD 0.216184f
C19 VDAC_N RST_Z 0.154233f
C20 a_3179_44403# a_3576_44364# 0.156867f
C21 a_4908_45956# a_6235_46124# 0.240532f
C22 a_18404_46526# VDD 0.134504f
C23 a_n133_43806# a_33_43806# 0.613203f
C24 a_8192_44874# VDD 1.04201f
C25 a_11427_43566# a_11252_43640# 0.234322f
C26 a_4322_46134# a_9179_44592# 0.148969f
C27 a_10447_44403# VDD 0.210712f
C28 a_17073_44056# VDD 0.267697f
C29 a_13023_42718# VDD 0.227979f
C30 a_9973_46526# VDD 0.494675f
C31 a_22959_44894# VDD 0.304443f
C32 a_10428_47338# a_10623_47307# 0.214221f
C33 a_3437_46532# VDD 0.279044f
C34 C4_N_btm VIN_N 0.502665f
C35 VDD DATA[5] 0.333656f
C36 C2_N_btm VCM 0.716172f
C37 C3_N_btm VREF 0.984942f
C38 a_10596_44324# a_10447_44403# 0.167531f
C39 a_10251_45454# a_14635_44324# 0.119134f
C40 a_948_43806# VDD 0.274505f
C41 a_12895_43640# VDD 0.198729f
C42 a_5655_43780# a_5351_43806# 0.152354f
C43 a_12896_47044# VDD 0.13999f
C44 VDAC_N VDD 4.59312f
C45 a_14950_43958# a_17715_44356# 0.35843f
C46 a_14853_45438# a_14953_45554# 0.167615f
C47 a_n2472_47044# VDD 0.293473f
C48 a_22733_47833# DEBUG_MUX[3] 0.200886f
C49 a_12833_42718# VDD 0.219881f
C50 a_10251_45454# a_16128_46134# 0.11558f
C51 a_18971_44654# a_18796_44728# 0.234322f
C52 a_n685_43268# a_n519_43268# 0.571005f
C53 a_2075_42870# a_2075_42718# 0.175451f
C54 a_3165_45982# a_3179_44403# 0.109673f
C55 a_10428_47338# a_10467_47212# 0.71995f
C56 a_n2833_47874# VDD 0.451564f
C57 a_3575_46697# VDD 0.666774f
C58 C3_N_btm VIN_N 0.455092f
C59 VDD DATA[4] 0.337633f
C60 C1_N_btm VCM 0.716121f
C61 C2_N_btm VREF 0.987884f
C62 a_16555_46616# a_16651_46500# 0.197934f
C63 a_10251_45454# a_16085_45982# 0.131882f
C64 a_1123_43780# VDD 0.462684f
C65 a_13113_43236# VDD 0.205187f
C66 a_5655_43780# a_5569_44048# 0.159469f
C67 a_11795_47044# VDD 0.409409f
C68 a_6886_37412# VDD 0.235486f
C69 a_4908_45956# a_5655_43780# 0.439759f
C70 SMPL_ON_N VIN_N 0.547248f
C71 a_8530_39574# a_3726_37500# 1.35509f
C72 a_10251_45454# a_15079_46134# 0.403004f
C73 a_11788_46134# a_13181_45982# 0.165846f
C74 a_15437_47044# a_15005_47222# 0.166981f
C75 a_4061_47044# a_4035_45609# 0.353032f
C76 a_3271_46532# VDD 0.49936f
C77 C2_N_btm VIN_N 0.502448f
C78 VDD DATA[3] 0.336359f
C79 C0_N_btm VCM 0.718136f
C80 C1_N_btm VREF 0.98698f
C81 a_n381_43433# a_n264_43628# 0.174251f
C82 a_636_42870# VDD 1.14989f
C83 a_383_43806# VDD 0.202202f
C84 a_12545_43268# VDD 0.245652f
C85 a_12684_45276# a_12287_44894# 0.159788f
C86 VDAC_N C10_N_btm 0.246383p
C87 a_22959_46534# VDD 0.308733f
C88 a_3470_45982# a_3165_45982# 0.137217f
C89 a_8055_45491# VDD 0.208706f
C90 a_10337_43268# a_11252_43640# 0.118759f
C91 VDAC_Ni a_6886_37412# 0.178275f
C92 a_7754_38470# a_3726_37500# 0.124796f
C93 a_11788_46134# a_13151_45956# 0.221092f
C94 a_22591_44894# VDD 0.283244f
C95 a_10150_47322# a_10467_47212# 0.102355f
C96 a_22400_42718# a_22465_38541# 0.231082f
C97 a_2645_46824# VDD 0.24457f
C98 C1_N_btm VIN_N 0.392375f
C99 VDD DATA[2] 0.332136f
C100 C0_dummy_N_btm VCM 0.311452f
C101 C0_N_btm VREF 0.444099f
C102 a_9159_43262# a_9898_44350# 0.170162f
C103 a_16291_44914# a_16555_46616# 0.111975f
C104 a_9343_45982# VDD 0.349695f
C105 a_601_44048# VDD 0.203312f
C106 EN_COMP a_1177_38525# 0.206071f
C107 a_12379_43268# VDD 0.441245f
C108 a_5655_43780# a_4835_43806# 0.296644f
C109 VDAC_N C9_N_btm 0.123396p
C110 a_n2293_43780# a_n2472_43780# 0.160389f
C111 a_10245_46532# a_10684_45670# 0.143941f
C112 a_3320_46134# a_3165_45982# 0.11586f
C113 a_10905_43236# a_10687_43640# 0.209641f
C114 COMP_N a_n501_42718# 0.194808f
C115 a_n2840_47044# VDD 0.306455f
C116 a_7754_38470# a_8530_39574# 0.143675f
C117 a_7851_46526# VDD 0.132317f
C118 a_17881_44356# a_18796_44728# 0.125324f
C119 a_15443_44582# a_15415_44350# 0.115039f
C120 a_19371_46579# a_19566_45670# 0.159295f
C121 a_22399_44894# VDD 0.462845f
C122 a_10150_47322# a_10428_47338# 0.118759f
C123 a_22775_42718# a_22465_38541# 0.330544f
C124 a_16475_45412# a_19566_45670# 0.160735f
C125 a_82_45670# VDD 1.17785f
C126 C0_N_btm VIN_N 0.529701f
C127 VDD DATA[1] 0.39041f
C128 C0_dummy_P_btm VCM 0.311452f
C129 a_10251_45454# a_15328_46134# 0.251056f
C130 a_16291_46758# a_16555_46616# 0.143485f
C131 a_16703_45982# a_16750_46134# 0.133906f
C132 a_8192_44874# a_8423_42718# 0.109681f
C133 a_8379_46134# VDD 0.140803f
C134 a_829_45221# VDD 0.193132f
C135 a_11788_46134# a_15468_45412# 0.121364f
C136 a_33_43806# VDD 0.415714f
C137 COMP_P a_1239_39587# 0.388739f
C138 a_11252_43640# VDD 0.275864f
C139 a_3726_37500# RST_Z 1.60318f
C140 a_10768_47436# VDD 0.132346f
C141 EN_VIN_BSTR_P a_n283_35174# 0.653211f
C142 VDAC_N C8_N_btm 61.725304f
C143 a_4908_45956# a_4700_46134# 0.188459f
C144 a_22223_46534# VDD 0.261133f
C145 a_3320_46134# a_3470_45982# 0.188181f
C146 a_10337_43268# a_10687_43640# 0.210642f
C147 a_10171_43268# a_11252_43640# 0.102355f
C148 a_13715_43780# a_16211_44582# 0.116158f
C149 a_10251_45454# a_15033_46526# 0.164515f
C150 a_17715_44356# a_18796_44728# 0.101963f
C151 a_18449_44324# a_18231_44728# 0.209641f
C152 a_22123_44894# VDD 0.407453f
C153 a_9517_46539# a_4908_45956# 0.383809f
C154 a_15133_43582# VDD 0.34574f
C155 C0_dummy_N_btm VIN_N 0.544204f
C156 VDD DATA[0] 0.3263f
C157 C0_P_btm VCM 0.718136f
C158 a_16291_46758# a_16291_44914# 0.220146f
C159 a_7552_46134# VDD 0.102045f
C160 a_n2293_43780# VDD 0.403439f
C161 a_n133_43806# VDD 0.506506f
C162 COMP_P a_22465_38541# 0.104544f
C163 a_11427_43566# VDD 0.455634f
C164 a_18689_45412# a_18803_47070# 0.213721f
C165 a_8530_39574# RST_Z 0.431385f
C166 VDAC_N C7_N_btm 30.8477f
C167 a_3726_37500# VDD 0.341303f
C168 a_3328_44324# a_3179_44403# 0.167531f
C169 a_10337_43268# a_10905_43236# 0.169363f
C170 a_10415_47846# a_9517_46539# 0.110775f
C171 a_15579_44172# VDD 0.132044f
C172 a_12427_42883# VDD 0.234353f
C173 a_13715_43780# a_15443_44582# 0.135399f
C174 a_17881_44356# a_18231_44728# 0.219399f
C175 a_3165_45982# a_3328_44324# 0.158757f
C176 a_22223_42718# a_22400_42718# 0.15592f
C177 a_12436_44868# a_12287_44894# 0.167531f
C178 VDD CLK_DATA 0.39166f
C179 a_1633_46824# VDD 0.213582f
C180 C1_P_btm VCM 0.716121f
C181 C0_P_btm VREF 0.444099f
C182 a_1387_45670# a_1659_45528# 0.13675f
C183 a_n2073_43806# VDD 0.354314f
C184 COMP_P a_22400_42718# 0.670553f
C185 a_10687_43640# VDD 0.198322f
C186 a_10901_42718# a_11183_42718# 0.201276f
C187 a_5419_47258# a_7227_46532# 0.250363f
C188 a_10251_45454# a_18803_47070# 0.295253f
C189 VDAC_N C6_N_btm 15.443401f
C190 a_8530_39574# VDD 0.346613f
C191 a_19566_45670# VDD 1.23228f
C192 a_10171_43268# a_10687_43640# 0.113784f
C193 COMP_P COMP_N 2.94856f
C194 a_11599_42883# VDD 0.254299f
C195 VDAC_Ni a_3726_37500# 1.5261f
C196 a_21629_47833# DEBUG_MUX[2] 0.222638f
C197 a_17715_44356# a_18231_44728# 0.11066f
C198 a_17881_44356# a_18449_44324# 0.17523f
C199 a_18247_46348# VDD 0.142103f
C200 a_14301_44035# a_14647_43494# 0.110063f
C201 a_9947_47044# a_10150_47322# 0.233657f
C202 a_571_46830# a_396_46904# 0.233657f
C203 C0_dummy_P_btm VIN_P 0.544204f
C204 VDD START 0.17687f
C205 C1_P_btm VREF 0.98698f
C206 C2_P_btm VCM 0.716172f
C207 a_22399_44894# a_22591_43958# 0.179992f
C208 a_6536_46348# VDD 0.142103f
C209 a_n2661_44332# a_n2293_44332# 0.216462f
C210 a_10905_43236# VDD 0.202023f
C211 a_5419_47258# a_6631_44582# 0.174501f
C212 a_18530_47070# a_18803_47070# 0.119431f
C213 VDAC_N C5_N_btm 7.727f
C214 a_7754_38470# VDD 0.302129f
C215 a_14635_44324# a_14545_44569# 0.185796f
C216 a_4908_45956# a_3165_45982# 0.310241f
C217 a_19371_46579# VDD 0.207529f
C218 a_10475_43433# a_10337_43268# 0.268976f
C219 a_9863_47874# a_9517_46539# 0.189169f
C220 COMP_P a_n1237_42718# 0.203614f
C221 a_17242_43806# VDD 0.201255f
C222 a_16475_45412# VDD 1.3744f
C223 a_11183_42718# VDD 0.225197f
C224 a_13715_43780# a_14133_43780# 0.266891f
C225 a_14573_47070# a_14757_45982# 0.254785f
C226 a_13003_43262# VDD 0.132317f
C227 C0_P_btm VIN_P 0.529701f
C228 VDD CLK 0.105075f
C229 a_396_46904# VDD 0.271327f
C230 C2_P_btm VREF 0.987884f
C231 C3_P_btm VCM 0.716273f
C232 a_11671_44019# a_11788_43806# 0.168541f
C233 a_16211_43780# a_16036_43806# 0.233657f
C234 a_6091_43780# a_5916_43806# 0.234322f
C235 a_10383_46697# a_10389_45438# 0.229511f
C236 a_2471_45046# VDD 0.217381f
C237 a_n2472_43780# VDD 0.27693f
C238 a_10337_43268# VDD 0.265635f
C239 a_17927_46195# a_18803_47070# 0.222028f
C240 a_n1586_35608# EN_VIN_BSTR_P 0.573165f
C241 VDAC_N C4_N_btm 3.90019f
C242 a_7760_45956# a_7981_45956# 0.101174f
C243 a_2687_45956# a_2512_45982# 0.233657f
C244 a_10171_43268# a_10337_43268# 0.735812f
C245 a_18879_45956# a_18704_45982# 0.233657f
C246 a_16036_43806# VDD 0.275246f
C247 a_16102_47044# VDD 0.251224f
C248 a_20159_47588# DEBUG_MUX[1] 0.228771f
C249 a_10901_42718# VDD 0.218725f
C250 a_17531_44894# a_17613_44894# 0.104085f
C251 a_17715_44356# a_17881_44356# 0.631599f
C252 a_18704_45982# VDD 0.293808f
C253 C3_P_btm VREF 0.984942f
C254 C1_P_btm VIN_P 0.392375f
C255 VDD RST_Z 1.26375f
C256 a_571_46830# VDD 0.335928f
C257 C4_P_btm VCM 0.716447f
C258 a_22399_44894# a_22031_44350# 0.287357f
C259 a_1663_45046# VDD 0.126255f
C260 a_10475_43433# VDD 0.531064f
C261 a_4035_45609# a_4322_46134# 0.154572f
C262 VDAC_N C3_N_btm 1.94557f
C263 a_7760_45956# a_7648_46134# 0.138043f
C264 a_15309_45438# a_11788_46134# 0.31466f
C265 a_4355_45438# VDD 0.132363f
C266 a_10171_43268# a_10475_43433# 0.172073f
C267 a_11299_47832# a_11507_47833# 0.136826f
C268 a_16211_43780# VDD 0.340832f
C269 a_7754_38636# a_7754_38470# 0.296258f
C270 a_18879_45956# VDD 0.35014f
C271 a_11788_46134# a_12121_45956# 0.222183f
C272 a_14757_47614# a_17927_46195# 0.127112f
C273 a_9943_45046# a_10215_44874# 0.13675f
C274 a_n519_46532# a_396_46904# 0.118423f
C275 a_n169_46904# VDD 0.213194f
C276 C4_P_btm VREF 0.98728f
C277 C2_P_btm VIN_P 0.502448f
C278 C5_P_btm VCM 0.719982f
C279 a_15192_46500# a_15309_45438# 0.124211f
C280 a_4993_47044# a_5536_44324# 0.136984f
C281 a_9349_46539# a_11415_45670# 0.102555f
C282 a_n2840_43780# VDD 0.302192f
C283 EN_COMP a_22465_38541# 0.54769f
C284 a_10171_43268# VDD 0.410111f
C285 a_4993_47044# a_6126_46642# 0.253663f
C286 VDAC_N C2_N_btm 1.04092f
C287 a_10596_44324# VDD 0.147006f
C288 a_15471_43806# VDD 0.199842f
C289 a_18135_47588# DEBUG_MUX[0] 0.230748f
C290 a_10069_42968# VDD 0.187255f
C291 a_18139_45982# VDD 0.2037f
C292 a_9943_45046# a_9304_43494# 0.102478f
C293 a_49_46500# a_n169_46904# 0.209641f
C294 a_n685_46532# a_396_46904# 0.102325f
C295 a_49_46500# VDD 0.218504f
C296 C5_P_btm VREF 0.987144f
C297 C3_P_btm VIN_P 0.455092f
C298 C6_P_btm VCM 0.877162f
C299 a_15192_46500# a_14757_45982# 0.12237f
C300 a_15121_43806# a_16036_43806# 0.118759f
C301 a_14757_43806# a_15376_43806# 0.159668f
C302 a_5001_43806# a_5916_43806# 0.118759f
C303 a_9349_46539# a_11017_45736# 0.170736f
C304 a_n2293_44868# VDD 0.309186f
C305 EN_COMP a_22400_42718# 0.407136f
C306 a_9637_43560# VDD 0.162425f
C307 a_4993_47044# a_5784_44364# 0.195031f
C308 VDAC_N C1_N_btm 0.562089f
C309 VDAC_Ni VDD 0.288547f
C310 a_1597_45982# a_2512_45982# 0.123255f
C311 a_17789_45982# a_18704_45982# 0.125324f
C312 a_5382_44582# a_5387_44403# 0.159139f
C313 a_9159_43262# VDD 0.447395f
C314 a_11143_47588# a_11299_47832# 0.414032f
C315 EN_COMP COMP_N 0.989098f
C316 a_15689_44048# VDD 0.204426f
C317 a_5663_45982# a_8055_45491# 0.173284f
C318 a_18357_46224# VDD 0.20998f
C319 a_10475_43433# a_9987_42968# 0.117754f
C320 a_n519_46532# a_n169_46904# 0.21686f
C321 a_n519_46532# VDD 0.286105f
C322 C6_P_btm VREF 1.41944f
C323 C4_P_btm VIN_P 0.502665f
C324 C10_N_btm VDD 2.40649f
C325 C7_P_btm VCM 1.58335f
C326 a_5569_44048# a_5351_43806# 0.209641f
C327 a_4835_43806# a_5916_43806# 0.102355f
C328 a_15689_44048# a_15471_43806# 0.209641f
C329 a_14955_43806# a_16036_43806# 0.102355f
C330 a_9349_46539# a_10389_45438# 0.351201f
C331 a_1209_47588# a_380_47222# 1.21533f
C332 SMPL a_22400_42718# 0.204987f
C333 VDAC_P C0_dummy_P_btm 0.297092f
C334 VDAC_N C0_N_btm 0.324396f
C335 a_n2038_35608# a_n1586_35608# 0.150796f
C336 a_10383_46697# a_10500_46892# 0.161235f
C337 a_2165_46224# a_1947_45982# 0.209641f
C338 a_17623_45982# a_18704_45982# 0.102325f
C339 a_18357_46224# a_18139_45982# 0.209641f
C340 a_9266_44350# VDD 0.208519f
C341 SMPL COMP_N 1.49521f
C342 a_15121_43806# VDD 0.342131f
C343 a_16335_47614# EN_OFFSET_CAL 0.194785f
C344 a_9987_42968# VDD 0.209595f
C345 a_17789_45982# VDD 0.577933f
C346 a_4322_46134# a_13469_44894# 0.287601f
C347 a_17531_44894# VDD 0.347961f
C348 a_2627_42718# a_2655_42870# 0.114056f
C349 a_n685_46532# VDD 0.483837f
C350 a_n519_46532# a_49_46500# 0.181217f
C351 a_n685_46532# a_n169_46904# 0.110532f
C352 C7_P_btm VREF 1.818f
C353 C5_P_btm VIN_P 0.502107f
C354 C9_N_btm VDD 0.345685f
C355 C8_P_btm VCM 2.61094f
C356 a_n381_43433# a_n519_43268# 0.322013f
C357 a_14470_46526# a_14757_45982# 0.10142f
C358 a_5001_43806# a_5351_43806# 0.21686f
C359 a_15121_43806# a_15471_43806# 0.218335f
C360 a_n2472_44868# VDD 0.276925f
C361 a_5655_43780# a_7020_44894# 0.212984f
C362 a_22591_43958# VDD 0.541259f
C363 a_7347_43494# VDD 0.250386f
C364 a_9987_42968# a_10069_42968# 0.171361f
C365 VDAC_N C0_dummy_N_btm 0.297444f
C366 VDAC_P C0_P_btm 0.324235f
C367 a_13469_44894# a_13561_44350# 0.113832f
C368 a_2134_44324# a_1736_43276# 0.109218f
C369 a_1431_45982# a_2512_45982# 0.102325f
C370 a_1597_45982# a_1947_45982# 0.207548f
C371 a_16475_45412# a_16824_45276# 0.948484f
C372 a_17789_45982# a_18139_45982# 0.220803f
C373 a_9335_44324# VDD 0.208486f
C374 EN_COMP COMP_P 10.149f
C375 a_14955_43806# VDD 0.452787f
C376 a_15437_47044# VDD 0.450409f
C377 a_22465_38541# a_22609_38842# 0.20695f
C378 a_9343_42718# VDD 0.262366f
C379 a_17623_45982# VDD 0.497466f
C380 a_9159_43262# a_9208_43494# 0.134846f
C381 a_12101_44048# VDD 0.209467f
C382 C8_P_btm VREF 3.6701f
C383 C6_P_btm VIN_P 0.391979f
C384 C9_P_btm VCM 6.06251f
C385 C8_N_btm VDD 0.19922f
C386 a_n381_43433# a_n685_43268# 0.146405f
C387 a_15121_43806# a_15689_44048# 0.171935f
C388 a_14955_43806# a_15471_43806# 0.103167f
C389 a_5001_43806# a_5569_44048# 0.181217f
C390 a_4835_43806# a_5351_43806# 0.110532f
C391 a_5655_43780# a_7195_44868# 0.270075f
C392 a_6519_43494# VDD 0.275264f
C393 a_n2472_44868# a_n2293_44868# 0.16963f
C394 a_18133_47235# a_14950_43958# 0.110384f
C395 a_16475_45412# a_12127_46744# 0.174033f
C396 a_n381_46697# a_n264_46892# 0.183714f
C397 VDAC_P C1_P_btm 0.561606f
C398 a_10079_46532# a_9973_46526# 0.12616f
C399 a_1597_45982# a_2165_46224# 0.173341f
C400 a_17623_45982# a_18139_45982# 0.107257f
C401 a_17789_45982# a_18357_46224# 0.177993f
C402 a_9140_44466# VDD 0.251279f
C403 SMPL COMP_P 6.57089f
C404 a_14757_43806# VDD 0.436695f
C405 a_22959_47622# VDD 0.243049f
C406 a_8423_42718# VDD 0.259801f
C407 a_7208_47044# a_19566_45670# 0.38243f
C408 a_6631_44582# a_7195_44868# 0.122363f
C409 a_8204_45412# a_8055_45491# 0.167531f
C410 a_11533_43806# VDD 0.391061f
C411 a_10795_43262# VDD 0.132284f
C412 a_n685_46532# a_n519_46532# 0.855623f
C413 a_n2472_46500# VDD 0.246993f
C414 C9_P_btm VREF 7.3695f
C415 C9_N_btm C10_N_btm 37.7035f
C416 C7_P_btm VIN_P 1.52459f
C417 C10_P_btm VCM 10.237201f
C418 C7_N_btm VDD 0.121904f
C419 a_5129_45956# VDD 0.157327f
C420 a_n2840_44868# VDD 0.302192f
C421 a_5655_43780# a_6455_44894# 0.181356f
C422 a_22031_44350# VDD 0.686954f
C423 a_4352_43640# VDD 0.293164f
C424 a_12747_47070# a_4908_45956# 0.107387f
C425 VDAC_P C2_P_btm 1.04676f
C426 a_16475_45412# a_15187_44868# 0.129899f
C427 a_15321_46526# VDD 0.200994f
C428 a_10844_44364# a_10414_43780# 0.126432f
C429 a_1431_45982# a_1947_45982# 0.110816f
C430 a_546_43100# a_468_42870# 0.205474f
C431 a_9179_44592# VDD 0.412686f
C432 a_7208_47044# a_19371_46579# 0.10194f
C433 a_12427_46758# VDD 0.145798f
C434 a_16824_45276# VDD 1.12472f
C435 a_284_47222# a_380_47222# 0.318297f
C436 a_16475_45412# a_7208_47044# 0.491615f
C437 a_11367_43806# VDD 0.401891f
C438 C10_P_btm VREF 14.776899f
C439 C8_N_btm C10_N_btm 0.607425f
C440 C8_P_btm VIN_P 0.907769f
C441 C6_N_btm VDD 0.210613f
C442 a_9140_44466# a_9159_43262# 0.556033f
C443 a_9335_44324# a_9266_44350# 0.209641f
C444 a_4279_46232# VDD 0.26765f
C445 a_14955_43806# a_15121_43806# 0.600991f
C446 a_4835_43806# a_5001_43806# 0.859504f
C447 a_5655_43780# a_6673_45136# 0.163603f
C448 a_18339_44350# VDD 0.142103f
C449 a_4527_43566# VDD 0.469304f
C450 VDAC_P C3_P_btm 1.95121f
C451 a_7760_45956# a_7552_46134# 0.230725f
C452 a_4908_45956# a_13266_45412# 0.204235f
C453 a_546_43100# a_1387_42883# 0.107644f
C454 a_1735_46195# a_1597_45982# 0.204866f
C455 a_17623_45982# a_17789_45982# 0.696827f
C456 a_8862_44482# VDD 0.279653f
C457 a_22733_47833# VDD 0.195741f
C458 a_3754_38802# VDAC_Ni 0.301032f
C459 a_15113_47222# a_15033_46526# 0.178543f
C460 a_12127_46744# VDD 0.585067f
C461 a_16427_44894# VDD 0.216111f
C462 a_8848_44868# a_8699_44894# 0.167531f
C463 a_n2840_46500# VDD 0.295278f
C464 C8_N_btm C9_N_btm 29.4361f
C465 C7_N_btm C10_N_btm 0.521459f
C466 C9_P_btm VIN_P 1.8284f
C467 C5_N_btm VDD 0.267489f
C468 a_9140_44466# a_9266_44350# 0.175128f
C469 a_9179_44592# a_9159_43262# 0.443401f
C470 a_13930_46842# a_14658_46526# 0.139577f
C471 a_14757_43806# a_15121_43806# 0.210823f
C472 a_82_45670# a_1339_43315# 0.122923f
C473 a_3787_43640# VDD 0.203412f
C474 a_15329_47044# a_15155_47070# 0.134825f
C475 a_7429_47044# VDD 0.158509f
C476 VDAC_P C4_P_btm 3.89919f
C477 a_9349_46539# a_9973_46526# 0.250164f
C478 a_1431_45982# a_1597_45982# 0.578623f
C479 a_8659_44324# VDD 0.356233f
C480 a_22223_47622# VDD 0.221814f
C481 VDAC_Pi a_6886_37412# 0.259481f
C482 a_22465_38541# a_22469_39973# 0.576946f
C483 a_10251_45454# a_16291_44914# 0.263779f
C484 a_11971_46500# VDD 0.304646f
C485 a_12379_44350# a_12461_44350# 0.171361f
C486 a_15187_44868# VDD 0.293409f
C487 a_6631_44582# a_6105_44894# 0.148911f
C488 a_18495_44868# VDD 0.211979f
C489 a_284_47222# a_85_47070# 0.24192f
C490 C7_N_btm C9_N_btm 0.206278f
C491 C6_N_btm C10_N_btm 0.317819f
C492 C10_P_btm VIN_P 3.66108f
C493 C4_N_btm VDD 0.265463f
C494 a_9140_44466# a_9335_44324# 0.209838f
C495 a_13930_46842# a_14470_46526# 0.166823f
C496 a_n2293_43244# a_n2472_43236# 0.174724f
C497 a_14757_43806# a_14955_43806# 0.188893f
C498 a_4005_43236# VDD 0.210988f
C499 a_10251_45454# a_14573_47070# 0.1252f
C500 a_7208_47044# VDD 1.01153f
C501 VDAC_P C5_P_btm 7.72615f
C502 a_1431_45982# a_1735_46195# 0.16027f
C503 a_546_43100# a_283_42692# 0.168785f
C504 a_7415_44466# VDD 0.127937f
C505 SMPL_ON_N RST_Z 2.26371f
C506 a_7556_42692# VDD 0.302278f
C507 a_7754_38968# a_7754_38636# 0.296258f
C508 a_11160_46904# VDD 0.278301f
C509 a_11533_43806# a_12101_44048# 0.171279f
C510 a_18319_44868# VDD 0.149767f
C511 a_21847_43806# a_21855_42718# 0.175524f
C512 a_9416_43530# VDD 0.28296f
C513 a_n193_47098# a_85_47070# 0.114867f
C514 a_n447_47044# a_n381_46697# 0.111762f
C515 C7_N_btm C8_N_btm 23.997501f
C516 C6_N_btm C9_N_btm 0.155878f
C517 C5_N_btm C10_N_btm 0.236062f
C518 a_20064_35138# VIN_N 0.367112f
C519 C3_N_btm VDD 0.26836f
C520 a_9179_44592# a_9335_44324# 0.107415f
C521 a_4322_46134# a_5655_43780# 0.448326f
C522 a_22031_45438# VDD 0.559647f
C523 a_5655_43780# a_5939_44894# 0.424145f
C524 a_656_45670# a_1387_45670# 0.118752f
C525 a_3437_43268# VDD 0.57711f
C526 a_n2661_44332# a_n2293_43244# 0.258627f
C527 a_5663_45982# VDD 0.99076f
C528 VDAC_P C6_P_btm 15.442699f
C529 a_4322_46134# a_3897_45444# 0.362676f
C530 a_14301_44035# VDD 0.220852f
C531 SMPL EN_COMP 0.545493f
C532 SMPL_ON_N VDD 0.502078f
C533 a_14757_47614# DEBUG_MUX[0] 0.229213f
C534 a_22465_38541# a_22545_39429# 0.253407f
C535 a_22400_42718# a_22821_39429# 0.136508f
C536 a_4322_46134# a_6631_44582# 0.250916f
C537 a_5382_44582# a_6126_46642# 0.170931f
C538 a_11335_46830# VDD 0.350821f
C539 a_11183_44350# a_11265_44350# 0.171361f
C540 a_11692_46134# a_11788_46134# 0.318454f
C541 a_17951_44868# VDD 0.224205f
C542 a_n193_47098# a_n194_47222# 0.119456f
C543 a_19037_42718# a_22223_42718# 0.178055f
C544 a_22959_47070# VDD 0.304494f
C545 C6_N_btm C8_N_btm 0.162414f
C546 C4_N_btm C10_N_btm 0.273376f
C547 C5_N_btm C9_N_btm 0.146663f
C548 EN_VIN_BSTR_N VCM 0.927905f
C549 C2_N_btm VDD 0.268945f
C550 a_9179_44592# a_9140_44466# 0.713769f
C551 a_n2661_43244# a_n2840_43236# 0.173451f
C552 a_9416_43530# a_9637_43560# 0.120571f
C553 a_656_45670# a_989_45736# 0.372162f
C554 a_20049_43262# a_22400_42718# 0.159114f
C555 a_3165_43262# VDD 0.335194f
C556 VDAC_P C7_P_btm 30.8471f
C557 a_13937_46602# VDD 0.256195f
C558 a_4322_46134# a_3731_45444# 0.3462f
C559 a_14077_44133# VDD 0.169924f
C560 a_n2288_42692# EN_COMP 0.157259f
C561 a_6631_42883# VDD 0.271567f
C562 a_22465_38541# a_22521_39947# 0.902378f
C563 a_21997_47833# VDD 0.192536f
C564 a_5382_44582# a_5784_44364# 0.670665f
C565 a_10595_46904# VDD 0.198947f
C566 a_15121_46232# VDD 0.168461f
C567 a_11367_43806# a_11533_43806# 0.630208f
C568 a_5784_44364# a_6243_45107# 0.326315f
C569 a_14204_44350# VDD 0.879903f
C570 a_n447_47044# a_n194_47222# 0.574208f
C571 C4_N_btm C9_N_btm 0.148287f
C572 C3_N_btm C10_N_btm 0.1871f
C573 C5_N_btm C8_N_btm 0.144827f
C574 C6_N_btm C7_N_btm 20.7485f
C575 C1_N_btm VDD 0.264503f
C576 a_8862_44482# a_9140_44466# 0.118759f
C577 a_10251_45454# a_11788_46134# 0.627384f
C578 a_3733_46348# VDD 0.145475f
C579 a_9416_43530# a_9208_43494# 0.186647f
C580 a_656_45670# a_361_45438# 0.107954f
C581 a_20049_43262# a_22775_42718# 0.238362f
C582 a_3271_43268# VDD 0.426871f
C583 a_7760_45956# VDD 0.371008f
C584 VDAC_P C8_P_btm 61.725f
C585 a_13373_46526# VDD 0.201758f
C586 a_15415_44350# a_15489_43268# 0.228886f
C587 a_4527_43566# a_4352_43640# 0.234322f
C588 a_4322_46134# a_4651_44350# 0.156906f
C589 a_7311_47614# a_7595_47614# 0.231974f
C590 a_14331_44133# VDD 0.104917f
C591 a_21629_47833# VDD 0.215165f
C592 VDAC_Pi a_3726_37500# 1.17174f
C593 a_5663_42718# VDD 0.26306f
C594 a_16703_45982# a_16291_44914# 0.174189f
C595 a_10813_46500# VDD 0.202305f
C596 a_15037_46232# VDD 0.151766f
C597 a_16576_44868# VDD 0.147876f
C598 EN_VIN_BSTR_N VIN_N 1.41696f
C599 C4_N_btm C8_N_btm 0.144911f
C600 C3_N_btm C9_N_btm 0.135794f
C601 C2_N_btm C10_N_btm 0.193308f
C602 C5_N_btm C7_N_btm 0.151868f
C603 C0_N_btm VDD 1.02806f
C604 a_8862_44482# a_9179_44592# 0.102355f
C605 a_13457_46892# a_14470_46526# 0.334357f
C606 a_2535_45670# VDD 0.13797f
C607 a_17763_44868# VDD 0.581382f
C608 a_560_45670# a_361_45438# 0.213677f
C609 a_6951_47070# a_6635_47044# 0.182065f
C610 a_16335_47614# a_16475_45412# 0.11032f
C611 a_14950_43958# a_15323_43268# 0.275453f
C612 a_2627_43262# VDD 0.260323f
C613 a_10251_45454# a_4908_45956# 0.883755f
C614 VDAC_P C9_P_btm 0.123395p
C615 a_22400_42718# VCM 0.19149f
C616 a_13207_46526# VDD 0.12327f
C617 a_8204_45412# VDD 0.123752f
C618 a_15415_44350# a_15323_43268# 0.23249f
C619 a_n2833_42692# SMPL 0.329111f
C620 a_12438_45412# a_12684_45276# 0.129687f
C621 a_22465_38541# a_22459_39581# 0.985539f
C622 a_20159_47588# VDD 0.268731f
C623 a_16427_44894# a_16824_45276# 0.155594f
C624 a_10245_46532# VDD 0.497144f
C625 a_22087_43244# a_22223_43494# 0.183402f
C626 a_16074_45046# VDD 0.125126f
C627 a_7493_43262# VDD 0.188359f
C628 a_22591_47070# VDD 0.310468f
C629 C3_N_btm C8_N_btm 0.13458f
C630 C2_N_btm C9_N_btm 0.140712f
C631 C1_N_btm C10_N_btm 0.182095f
C632 C5_N_btm C6_N_btm 18.5121f
C633 C4_N_btm C7_N_btm 0.145744f
C634 EN_VIN_BSTR_P VCM 0.929333f
C635 a_83_45776# a_361_45438# 0.112535f
C636 a_560_45670# a_656_45670# 0.31839f
C637 a_15589_44350# VDD 0.17658f
C638 a_1339_43315# VDD 0.222943f
C639 VDAC_P C10_P_btm 0.246383p
C640 a_22400_42718# VREF 0.106195f
C641 a_22609_38842# a_22609_38426# 0.32625f
C642 a_7705_45736# VDD 0.16212f
C643 a_22223_43494# a_22223_43270# 0.208338f
C644 a_6951_47070# a_7311_47614# 0.138795f
C645 a_14950_43958# a_17623_43806# 0.287893f
C646 COMP_N VREF 0.128449f
C647 a_22465_38541# a_22521_40491# 0.214039f
C648 a_22400_42718# a_22459_39581# 0.242947f
C649 a_18135_47588# VDD 0.271165f
C650 a_4791_42883# VDD 0.262948f
C651 a_10383_46697# VDD 0.440105f
C652 a_15323_44894# VDD 0.225458f
C653 a_6665_43262# VDD 0.193494f
C654 C2_N_btm C8_N_btm 0.139221f
C655 C1_N_btm C9_N_btm 0.130686f
C656 C0_N_btm C10_N_btm 0.230054f
C657 C4_N_btm C6_N_btm 0.14422f
C658 C3_N_btm C7_N_btm 0.13519f
C659 a_17531_44894# a_18136_44716# 0.157914f
C660 a_8659_44324# a_8862_44482# 0.233657f
C661 a_13457_46892# a_13930_46842# 0.201865f
C662 a_n61_43262# VDD 0.157273f
C663 a_7754_39632# VDD 0.205733f
C664 a_4833_47320# VDD 0.203491f
C665 CAL_P a_22609_38426# 0.205305f
C666 a_22031_45438# a_22031_44350# 0.117355f
C667 a_11971_46500# a_12127_46744# 0.238033f
C668 a_16921_46364# VDD 0.725714f
C669 a_6985_45438# VDD 0.31619f
C670 a_3437_43268# a_4352_43640# 0.124988f
C671 a_4733_44350# VDD 0.190838f
C672 a_14950_43958# a_17515_43806# 0.200434f
C673 a_21197_42718# a_21303_42718# 0.110402f
C674 a_7754_39964# a_7754_38470# 0.241119f
C675 a_22400_42718# a_22521_40491# 0.681186f
C676 a_16335_47614# VDD 0.21551f
C677 COMP_P VCM 0.117667f
C678 a_3754_39134# a_3754_38802# 0.296258f
C679 a_4239_42883# VDD 0.232406f
C680 a_10079_46532# VDD 0.391023f
C681 a_16750_46134# VDD 0.180108f
C682 a_14635_44324# VDD 0.533893f
C683 a_7851_44172# VDD 0.142103f
C684 a_4993_47044# a_5749_47222# 0.720518f
C685 a_7208_47044# a_12127_46744# 0.140403f
C686 C0_P_btm VDD 1.02806f
C687 C1_N_btm C8_N_btm 0.12931f
C688 C0_N_btm C9_N_btm 0.144582f
C689 C0_dummy_N_btm C10_N_btm 0.397081f
C690 C4_N_btm C5_N_btm 16.137598f
C691 C3_N_btm C6_N_btm 0.13406f
C692 C2_N_btm C7_N_btm 0.138838f
C693 a_15605_45438# VDD 0.198957f
C694 a_5839_47070# a_5749_47222# 0.109471f
C695 a_4035_45609# VDD 0.486983f
C696 a_16128_46134# VDD 0.343744f
C697 a_7372_45670# VDD 0.825228f
C698 a_4005_43236# a_3787_43640# 0.209641f
C699 a_22087_43244# a_21908_43236# 0.188236f
C700 a_22223_43494# a_21719_43244# 0.125271f
C701 a_7208_47044# a_7429_47044# 0.15357f
C702 a_15871_47614# VDD 0.149325f
C703 COMP_P VREF 0.415113f
C704 a_3823_42718# VDD 0.228325f
C705 a_9547_46565# VDD 0.100025f
C706 a_16085_45982# VDD 0.43763f
C707 a_4993_47044# a_5419_47258# 0.43668f
C708 C1_P_btm VDD 0.264503f
C709 EN_VIN_BSTR_P VIN_P 1.41696f
C710 C3_N_btm C5_N_btm 0.135784f
C711 C0_N_btm C8_N_btm 0.146681f
C712 C0_dummy_N_btm C9_N_btm 0.112646f
C713 C2_N_btm C6_N_btm 0.137649f
C714 C1_N_btm C7_N_btm 0.128768f
C715 a_7016_46231# a_6954_46348# 0.157972f
C716 a_7347_43494# a_7493_43262# 0.171361f
C717 VDAC_Pi VDD 0.591846f
C718 a_7754_39964# RST_Z 0.843939f
C719 a_15079_46134# VDD 0.577649f
C720 a_3271_43268# a_4352_43640# 0.102325f
C721 a_3437_43268# a_3787_43640# 0.229804f
C722 a_12127_46744# a_17951_44868# 0.232417f
C723 a_21197_42718# a_21027_42718# 0.109088f
C724 a_15691_47614# VDD 0.178828f
C725 a_22465_38541# a_22521_41035# 0.132396f
C726 a_22400_42718# a_22469_41061# 0.954898f
C727 a_7754_39300# a_7754_38968# 0.296258f
C728 a_3541_42718# VDD 0.240932f
C729 a_18319_44868# a_18495_44868# 0.185422f
C730 a_14204_44350# a_16824_45276# 0.209609f
C731 a_12684_45276# a_12683_43433# 0.388974f
C732 a_15582_45982# a_15309_45438# 0.126444f
C733 a_9293_46565# VDD 0.174771f
C734 a_14955_45982# VDD 0.205018f
C735 a_10414_43780# VDD 0.282341f
C736 a_4993_47044# a_5089_47044# 0.163078f
C737 C2_P_btm VDD 0.268945f
C738 C2_N_btm C5_N_btm 0.138263f
C739 C3_N_btm C4_N_btm 7.944839f
C740 C1_N_btm C6_N_btm 0.127984f
C741 C0_dummy_N_btm C8_N_btm 0.237239f
C742 C0_N_btm C7_N_btm 0.141209f
C743 a_10475_43433# a_10592_43628# 0.159936f
C744 a_22469_39973# a_22609_38426# 0.490939f
C745 a_7754_39964# VDD 0.848281f
C746 a_1387_44582# a_1659_44440# 0.13675f
C747 a_6707_45776# VDD 0.19755f
C748 a_3437_43268# a_4005_43236# 0.186387f
C749 a_6491_44716# VDD 0.402085f
C750 a_5839_47070# a_5847_47614# 0.218998f
C751 a_15139_47730# VDD 0.14187f
C752 a_5663_45982# a_7208_47044# 0.291725f
C753 a_22400_42718# a_22521_41035# 0.133592f
C754 VDAC_Pi VDAC_Ni 3.18068f
C755 a_9349_46539# VDD 1.08305f
C756 a_636_42870# a_468_42870# 0.105626f
C757 a_9863_43958# VDD 0.212536f
C758 a_22223_47070# VDD 0.283428f
C759 C3_P_btm VDD 0.26836f
C760 C2_N_btm C4_N_btm 7.37802f
C761 C1_N_btm C5_N_btm 0.127667f
C762 C0_N_btm C6_N_btm 0.139432f
C763 C0_dummy_N_btm C7_N_btm 0.12244f
C764 a_7309_44466# a_7415_44466# 0.13675f
C765 a_2055_46348# VDD 0.134504f
C766 a_6519_43494# a_6665_43262# 0.171361f
C767 a_11335_46830# a_11160_46904# 0.233657f
C768 a_7208_47044# a_19168_45758# 0.141853f
C769 a_6325_45736# VDD 0.162248f
C770 a_3271_43268# a_3787_43640# 0.110532f
C771 a_5387_44403# VDD 0.214403f
C772 a_11991_44172# VDD 0.137588f
C773 a_7760_45956# a_7429_47044# 0.144147f
C774 a_2801_42968# VDD 0.175227f
C775 a_7754_39964# VDAC_Ni 0.207118f
C776 a_16576_44868# a_16427_44894# 0.167531f
C777 a_8308_46904# VDD 0.280609f
C778 a_1736_43276# a_2627_42718# 0.54596f
C779 a_15328_46134# VDD 0.31481f
C780 a_12127_46744# a_17763_44868# 0.119021f
C781 a_13469_44894# VDD 0.210271f
C782 a_9343_43806# VDD 0.272524f
C783 a_4704_47044# a_5089_47044# 0.126169f
C784 C4_P_btm VDD 0.265463f
C785 a_n1586_35608# VIN_P 0.367112f
C786 C1_N_btm C4_N_btm 0.128431f
C787 C0_N_btm C5_N_btm 0.138379f
C788 C2_N_btm C3_N_btm 5.69083f
C789 C0_dummy_N_btm C6_N_btm 0.122824f
C790 a_82_45670# a_1488_43236# 0.155815f
C791 a_20283_43262# a_20383_42718# 0.174404f
C792 a_n2293_44332# a_n2472_44324# 0.169554f
C793 a_22469_39973# a_22609_38842# 0.198764f
C794 a_15033_46526# VDD 0.522104f
C795 a_636_42870# a_571_43566# 0.114052f
C796 a_5419_47258# a_7842_44868# 0.264389f
C797 a_3165_43262# a_3437_43268# 0.235263f
C798 a_5139_44019# VDD 0.443187f
C799 a_8483_46830# VDD 0.369728f
C800 a_636_42870# a_428_42724# 0.124528f
C801 a_8308_43806# VDD 0.299225f
C802 COMP_P a_22521_41035# 0.201896f
C803 C5_P_btm VDD 0.267489f
C804 C0_N_btm C4_N_btm 0.138615f
C805 C0_dummy_N_btm C5_N_btm 0.117097f
C806 C1_N_btm C3_N_btm 7.588649f
C807 a_7016_46231# VDD 0.439585f
C808 a_14077_44133# a_14301_44035# 0.101354f
C809 a_15415_44350# a_15744_43628# 0.160322f
C810 a_22959_45446# VDD 0.29903f
C811 a_21540_43236# a_21719_43244# 0.175513f
C812 a_13819_44350# VDD 0.190131f
C813 a_21997_47833# SMPL_ON_N 0.198659f
C814 a_n1429_43262# VDD 0.474044f
C815 a_10251_45454# a_18689_45412# 0.156506f
C816 a_22521_39947# a_22609_38426# 0.333805f
C817 VDAC_N EN_VIN_BSTR_N 0.33104f
C818 a_18803_47070# a_18822_46526# 0.157972f
C819 a_3271_43268# a_3437_43268# 0.901096f
C820 a_19566_45670# a_18970_45412# 0.118887f
C821 a_13536_43780# VDD 0.238143f
C822 a_11248_47319# a_11186_47436# 0.15568f
C823 a_2655_42870# VDD 0.203565f
C824 EN_COMP VREF 0.436981f
C825 SMPL VCM 0.415258f
C826 a_7743_46904# VDD 0.195871f
C827 a_14819_44582# a_15091_44440# 0.13675f
C828 a_14382_46348# VDD 0.287972f
C829 a_19520_46500# a_19371_46579# 0.167531f
C830 a_n105_46195# a_361_45438# 0.22352f
C831 a_8483_43780# VDD 0.494804f
C832 a_19037_42718# a_19187_42718# 0.14775f
C833 a_8969_43582# VDD 0.462725f
C834 EN_COMP a_22459_39581# 0.415926f
C835 a_18803_47070# VDD 0.324953f
C836 C6_P_btm VDD 0.210613f
C837 C0_N_btm C3_N_btm 0.409922f
C838 C1_N_btm C2_N_btm 5.10246f
C839 C0_dummy_N_btm C4_N_btm 0.116511f
C840 a_3575_46697# a_4061_45956# 0.112953f
C841 a_13427_46756# a_13457_46892# 0.345508f
C842 a_6322_46348# VDD 0.205536f
C843 a_14331_44133# a_14301_44035# 0.191278f
C844 a_15139_47730# a_15437_47044# 0.100719f
C845 a_12461_44350# VDD 0.193651f
C846 a_n1741_42692# VDD 0.428519f
C847 a_n2661_44332# a_n2840_44324# 0.180301f
C848 VDAC_P EN_VIN_BSTR_P 0.328367f
C849 a_n2661_43244# a_n2293_43244# 0.385024f
C850 a_10245_46532# a_11160_46904# 0.117156f
C851 a_4812_45816# VDD 0.278927f
C852 a_3271_43268# a_3165_43262# 0.396956f
C853 a_4091_47070# a_4651_47614# 0.223504f
C854 a_12448_43806# VDD 0.276211f
C855 SMPL VREF 1.00301f
C856 a_2075_42718# VDD 0.289476f
C857 a_7961_46500# VDD 0.201518f
C858 a_14819_44582# a_14133_43780# 0.100092f
C859 a_14194_46348# VDD 0.237618f
C860 a_11059_45956# a_10884_45982# 0.233657f
C861 a_12287_44894# VDD 0.217102f
C862 a_7743_43806# VDD 0.196098f
C863 SMPL_ON_P a_n2038_35608# 0.39925f
C864 a_18445_42718# a_19187_42718# 0.171185f
C865 a_7735_42692# VDD 0.4525f
C866 EN_COMP a_22521_40491# 0.260972f
C867 C7_P_btm VDD 0.121904f
C868 C0_N_btm C2_N_btm 0.698837f
C869 a_6391_46219# VDD 0.203777f
C870 a_22455_45420# VDD 0.357155f
C871 a_11265_44350# VDD 0.190422f
C872 a_19633_43262# a_21303_42718# 0.17018f
C873 a_713_47044# VDD 0.151418f
C874 a_22521_39947# a_22609_38842# 0.23688f
C875 a_22459_39581# a_22609_38426# 0.172129f
C876 a_10813_46500# a_10595_46904# 0.209641f
C877 a_847_45956# a_672_45982# 0.233657f
C878 a_9159_43262# a_8969_43582# 0.129265f
C879 a_380_47222# a_1663_45046# 0.100635f
C880 a_4987_45742# VDD 0.348231f
C881 a_2627_43262# a_3165_43262# 0.119318f
C882 a_12623_43780# VDD 0.462939f
C883 a_15187_44868# a_14635_44324# 0.521291f
C884 a_14757_47614# VDD 0.399746f
C885 a_3754_39466# a_3754_39134# 0.296258f
C886 a_7393_46532# VDD 0.265637f
C887 a_14545_44569# a_14133_43780# 0.13311f
C888 a_5663_45982# a_7705_45736# 0.120128f
C889 a_21719_43244# a_20049_43262# 0.325829f
C890 a_7961_44048# VDD 0.203316f
C891 a_18445_42718# a_19037_42718# 0.133606f
C892 C8_P_btm VDD 0.19922f
C893 C0_N_btm C1_N_btm 11.1057f
C894 C0_dummy_N_btm C2_N_btm 6.84965f
C895 a_6235_46124# VDD 0.419878f
C896 a_22276_45412# VDD 0.300131f
C897 a_4091_47070# a_4061_47044# 0.102717f
C898 a_17927_46195# a_10251_45454# 0.187385f
C899 a_380_47222# VDD 0.911834f
C900 a_2684_37794# VDD 0.286898f
C901 a_22521_40491# a_22609_38426# 0.234448f
C902 a_10245_46532# a_10595_46904# 0.218763f
C903 a_10079_46532# a_11160_46904# 0.102355f
C904 a_19520_46500# VDD 0.142917f
C905 a_4908_45956# a_10111_45776# 0.127495f
C906 a_4247_45816# VDD 0.192118f
C907 a_11883_43806# VDD 0.20547f
C908 a_9551_47203# VDD 1.22917f
C909 a_2113_38308# VDAC_Ni 0.315941f
C910 a_7503_45982# VDD 0.450342f
C911 a_13661_46298# VDD 0.256644f
C912 a_5663_45982# a_6985_45438# 0.128862f
C913 a_16475_45412# a_16287_45744# 0.202881f
C914 a_7393_43806# VDD 0.581175f
C915 a_7372_45670# a_7415_44466# 0.100399f
C916 C9_P_btm VDD 0.345685f
C917 C0_dummy_N_btm C1_N_btm 1.25238f
C918 a_6196_46250# VDD 0.504321f
C919 a_18970_45412# VDD 0.299714f
C920 a_17927_46195# a_18530_47070# 0.233767f
C921 a_n381_46697# VDD 0.376622f
C922 a_1177_38525# VDD 0.373545f
C923 a_22459_39581# a_22609_38842# 0.12318f
C924 a_10245_46532# a_10813_46500# 0.171912f
C925 a_18190_46526# VDD 0.204312f
C926 a_4465_45412# VDD 0.208076f
C927 a_8969_43582# a_9343_42718# 0.166198f
C928 a_7754_39632# a_7754_39300# 0.296258f
C929 a_7227_46532# VDD 0.455412f
C930 a_9969_45982# a_10884_45982# 0.117156f
C931 a_7319_43262# VDD 0.442693f
C932 a_18759_42746# a_19037_42718# 0.112562f
C933 a_18361_47320# VDD 0.195068f
C934 C10_P_btm VDD 2.40649f
C935 C0_dummy_N_btm C0_N_btm 7.84944f
C936 a_5655_43780# VDD 1.41441f
C937 a_18282_45670# VDD 0.138595f
C938 a_9480_44350# VDD 0.1325f
C939 a_10251_45454# a_19003_43262# 0.24035f
C940 a_1488_43236# VDD 0.15221f
C941 a_85_47070# VDD 0.220213f
C942 a_2112_39137# VDD 0.284849f
C943 a_22521_40491# a_22609_38842# 0.1922f
C944 a_22469_41061# a_22609_38426# 0.130478f
C945 a_10079_46532# a_10595_46904# 0.104565f
C946 a_18259_46500# VDD 0.194344f
C947 a_n105_46195# a_12_45982# 0.161376f
C948 a_n243_45982# a_672_45982# 0.125324f
C949 a_3897_45444# VDD 0.248869f
C950 a_2343_47070# a_2351_47614# 0.224073f
C951 SMPL_ON_P SMPL 2.4279f
C952 a_11415_45670# a_11687_45528# 0.13675f
C953 a_468_42870# VDD 0.232854f
C954 a_6631_44582# VDD 1.4778f
C955 a_4035_45609# a_4152_45804# 0.170785f
C956 a_9803_45982# a_10884_45982# 0.102325f
C957 a_10537_46224# a_10319_45982# 0.209641f
C958 a_9304_43494# VDD 0.785062f
C959 a_19771_43600# a_20049_43262# 0.112563f
C960 a_7227_43806# VDD 0.493915f
C961 a_6243_45107# a_6360_44894# 0.157972f
C962 a_14950_43958# VDD 0.93129f
C963 a_21789_35634# VDD 0.523706f
C964 a_5918_46234# VDD 0.276687f
C965 a_3699_43780# a_3524_43806# 0.234322f
C966 a_16287_45744# VDD 0.229588f
C967 a_15415_44350# VDD 0.460063f
C968 a_2343_47070# a_2167_46526# 0.113725f
C969 a_10251_45454# a_18766_43236# 0.204361f
C970 a_396_43640# VDD 0.28022f
C971 a_n381_46697# a_n519_46532# 0.220835f
C972 a_n194_47222# VDD 1.24745f
C973 a_22545_39429# a_22821_39429# 0.235701f
C974 a_22521_39947# a_22469_39973# 1.02751f
C975 a_10383_46697# a_10245_46532# 0.281236f
C976 a_18064_46642# VDD 0.31723f
C977 a_325_46224# a_107_45982# 0.209641f
C978 a_11533_43806# a_12448_43806# 0.118423f
C979 a_3731_45444# VDD 0.443046f
C980 a_5536_44324# VDD 0.177079f
C981 a_5655_43780# a_9159_43262# 0.278672f
C982 a_1387_42883# VDD 0.248037f
C983 a_6126_46642# VDD 0.203339f
C984 a_5663_45982# a_6707_45776# 0.153585f
C985 a_9863_43958# a_9416_43530# 0.110214f
C986 a_9969_45982# a_10319_45982# 0.21686f
C987 a_5473_43582# VDD 0.523711f
C988 a_16671_47320# VDD 0.242615f
C989 a_20064_35138# VDD 0.317561f
C990 C3_P_btm C3_N_btm 1.60138f
C991 a_7208_47044# a_15328_46134# 0.42513f
C992 a_5715_45956# VDD 0.34439f
C993 a_9304_43494# a_9637_43560# 0.23339f
C994 a_2627_42718# a_2864_43806# 0.158041f
C995 a_16111_45412# VDD 0.145141f
C996 a_18766_43236# a_21197_42718# 0.127506f
C997 a_22959_44358# VDD 0.298068f
C998 a_571_43566# VDD 0.343528f
C999 a_n381_46697# a_n685_46532# 0.281644f
C1000 a_12896_47044# a_4908_45956# 0.12667f
C1001 a_4993_47044# a_5382_44582# 0.516895f
C1002 a_5089_47044# a_4322_46134# 0.150419f
C1003 a_5419_47258# a_5441_46500# 0.130857f
C1004 a_11248_47319# VDD 0.629645f
C1005 a_22521_39947# a_22821_39429# 0.112629f
C1006 a_1239_39043# VDD 0.507578f
C1007 a_10079_46532# a_10245_46532# 0.696021f
C1008 a_7503_45982# a_7648_46892# 0.159135f
C1009 a_18103_46768# VDD 0.4118f
C1010 a_n243_45982# a_107_45982# 0.219633f
C1011 a_n409_45982# a_672_45982# 0.102355f
C1012 a_12101_44048# a_11883_43806# 0.209641f
C1013 a_11367_43806# a_12448_43806# 0.102355f
C1014 a_2151_45670# VDD 0.442092f
C1015 a_14955_45982# a_15121_46232# 0.143754f
C1016 a_4651_44350# VDD 0.181788f
C1017 a_5655_43780# a_9266_44350# 0.175191f
C1018 a_428_42724# VDD 0.115396f
C1019 a_14635_44324# a_16074_45046# 0.14815f
C1020 a_5784_44364# VDD 1.43891f
C1021 a_13151_45956# VDD 0.31891f
C1022 a_9803_45982# a_10319_45982# 0.110532f
C1023 a_9969_45982# a_10537_46224# 0.181217f
C1024 a_4322_46134# a_12931_44894# 0.184319f
C1025 a_3895_43262# VDD 0.142104f
C1026 a_7195_44868# a_7020_44894# 0.233657f
C1027 a_19320_35138# VDD 0.322581f
C1028 a_4700_46134# VDD 0.105613f
C1029 a_9304_43494# a_9208_43494# 0.319593f
C1030 a_13715_43780# VDD 0.53776f
C1031 a_7319_43262# a_7347_43494# 0.13713f
C1032 a_19003_43262# a_19191_43262# 0.141213f
C1033 a_22223_44358# VDD 0.274783f
C1034 a_n169_43640# VDD 0.221249f
C1035 a_4993_47044# a_4322_46134# 0.281041f
C1036 a_15582_45982# a_10251_45454# 0.131925f
C1037 a_10554_47436# VDD 0.197831f
C1038 a_22521_39947# a_22545_39429# 0.27533f
C1039 a_22459_39581# a_22469_39973# 0.351623f
C1040 a_10079_46532# a_10383_46697# 0.162368f
C1041 a_17786_46658# VDD 0.278159f
C1042 a_n243_45982# a_325_46224# 0.175891f
C1043 a_n2073_43806# a_n2104_43236# 0.221106f
C1044 a_11533_43806# a_11883_43806# 0.218541f
C1045 a_3882_44324# VDD 0.287827f
C1046 a_5655_43780# a_9335_44324# 0.160674f
C1047 a_9517_46539# VDD 0.322084f
C1048 a_283_42692# VDD 0.260222f
C1049 a_9863_47874# DEBUG_OUT 0.329921f
C1050 a_14635_44324# a_15323_44894# 0.200592f
C1051 a_3575_46697# a_3692_46892# 0.159828f
C1052 a_13097_46348# VDD 0.201758f
C1053 a_14950_43958# a_17531_44894# 0.202365f
C1054 a_4322_46134# a_12436_44868# 0.172027f
C1055 a_7372_45670# a_7705_45736# 0.205648f
C1056 a_15962_47320# VDD 0.184829f
C1057 C0_P_btm C0_dummy_P_btm 7.84944f
C1058 a_2609_43806# a_3524_43806# 0.125324f
C1059 a_16921_46364# a_16750_46134# 0.162771f
C1060 a_15468_45412# VDD 0.17431f
C1061 a_21755_44350# VDD 0.45549f
C1062 a_49_43236# VDD 0.221845f
C1063 a_12896_47044# a_12747_47070# 0.167531f
C1064 CAL_N a_22609_38842# 0.204621f
C1065 a_10623_47307# VDD 0.194685f
C1066 a_5663_45982# a_7016_46231# 0.121894f
C1067 a_17583_46500# VDD 0.358374f
C1068 a_n409_45982# a_107_45982# 0.110816f
C1069 a_11367_43806# a_11883_43806# 0.10279f
C1070 a_3576_44364# VDD 1.40038f
C1071 a_999_47846# a_1209_47588# 0.146768f
C1072 a_14950_43958# a_14955_43806# 0.445935f
C1073 VDAC_Pi a_3754_39466# 0.308867f
C1074 a_14587_47614# START 0.190445f
C1075 a_12684_45276# a_13991_42883# 0.108494f
C1076 a_12931_46348# VDD 0.125433f
C1077 a_9803_45982# a_9969_45982# 0.882077f
C1078 a_7372_45670# a_6985_45438# 0.13458f
C1079 a_16475_45412# a_16291_44914# 0.121519f
C1080 EN_VIN_BSTR_N VDD 1.32068f
C1081 C1_P_btm C0_dummy_P_btm 1.25238f
C1082 a_4061_45956# VDD 0.195732f
C1083 a_3177_44048# a_2959_43806# 0.209641f
C1084 a_14953_45554# VDD 0.196549f
C1085 a_18796_44728# VDD 0.307716f
C1086 a_n519_43268# VDD 0.536784f
C1087 a_16561_45982# a_16703_45982# 0.775861f
C1088 a_22459_39581# a_22545_39429# 0.121283f
C1089 a_22521_40491# a_22821_39429# 0.131339f
C1090 CAL_N CAL_P 6.10044f
C1091 a_1239_39587# VDD 0.529955f
C1092 a_10467_47212# VDD 0.441934f
C1093 a_16651_46500# VDD 0.130905f
C1094 a_n105_46195# a_n243_45982# 0.214791f
C1095 a_82_45670# a_1736_43276# 0.132129f
C1096 a_3179_44403# VDD 0.265862f
C1097 a_14950_43958# a_14757_43806# 0.246268f
C1098 a_7735_42692# a_7556_42692# 0.169093f
C1099 a_5655_43780# a_9179_44592# 0.325147f
C1100 a_104_42692# VDD 0.276761f
C1101 a_7595_47614# DATA[5] 0.355242f
C1102 a_13715_43780# a_15121_43806# 0.414724f
C1103 a_3895_46526# VDD 0.132317f
C1104 a_8699_44894# VDD 0.262208f
C1105 a_21197_42718# a_19633_43262# 0.27574f
C1106 a_7276_45670# a_6985_45438# 0.217735f
C1107 a_1115_47044# a_1431_47070# 0.133144f
C1108 a_6105_44894# a_7020_44894# 0.118759f
C1109 C2_P_btm C0_dummy_P_btm 6.84965f
C1110 C1_P_btm C0_P_btm 11.1057f
C1111 a_3165_45982# VDD 0.760484f
C1112 a_2609_43806# a_2959_43806# 0.222782f
C1113 a_2443_43806# a_3524_43806# 0.102355f
C1114 a_16128_46134# a_16085_45982# 0.120717f
C1115 a_14853_45438# VDD 0.16923f
C1116 a_18971_44654# VDD 0.549305f
C1117 a_n685_43268# VDD 0.479888f
C1118 a_22469_41061# a_22469_39973# 0.604831f
C1119 a_22465_38541# VDD 1.31228f
C1120 a_10428_47338# VDD 0.248002f
C1121 a_22400_42718# RST_Z 0.26468f
C1122 a_16555_46616# VDD 0.279439f
C1123 a_n409_45982# a_n243_45982# 0.584389f
C1124 a_82_45670# a_2134_44324# 0.202213f
C1125 a_663_47874# a_999_47846# 0.254397f
C1126 a_18093_43262# a_18348_43262# 0.114664f
C1127 a_5655_43780# a_8862_44482# 0.22079f
C1128 a_n501_42718# VDD 0.27866f
C1129 a_12887_47833# CLK 0.215051f
C1130 a_7754_39964# a_7754_39632# 0.296522f
C1131 a_636_42870# a_768_44670# 0.147971f
C1132 a_7208_47044# a_19520_46500# 0.130221f
C1133 a_13715_43780# a_14955_43806# 0.434352f
C1134 VREF VCM 19.8663f
C1135 a_15079_46134# a_16128_46134# 0.212032f
C1136 a_5419_47258# a_8192_44874# 0.120113f
C1137 a_12684_45276# a_12833_42718# 0.110804f
C1138 a_12127_46744# a_18282_45670# 0.145381f
C1139 a_14950_43958# a_16824_45276# 0.331169f
C1140 a_7276_45670# a_7372_45670# 0.322481f
C1141 a_6707_45776# a_6985_45438# 0.112567f
C1142 a_5459_44172# VDD 0.13244f
C1143 a_9551_47203# a_7208_47044# 0.207554f
C1144 a_2709_43262# VDD 0.190016f
C1145 a_6673_45136# a_6455_44894# 0.209641f
C1146 EN_VIN_BSTR_N C10_N_btm 0.320716f
C1147 a_n283_35174# VDD 0.295224f
C1148 C2_P_btm C0_P_btm 0.698837f
C1149 a_82_45670# a_1597_45982# 0.168419f
C1150 a_3470_45982# VDD 0.13294f
C1151 a_22399_44894# a_22959_43806# 0.179691f
C1152 a_2609_43806# a_3177_44048# 0.180299f
C1153 a_18231_44728# VDD 0.200102f
C1154 a_15691_47614# a_15871_47614# 0.185422f
C1155 a_n2104_43236# VDD 0.285703f
C1156 a_3541_42718# a_3823_42718# 0.213334f
C1157 a_22521_41035# a_22469_39973# 0.380006f
C1158 a_22521_40491# a_22521_39947# 0.457858f
C1159 a_22400_42718# VDD 0.564661f
C1160 a_5663_45982# a_6235_46124# 0.278198f
C1161 a_16291_44914# VDD 1.84595f
C1162 a_n409_45982# a_n105_46195# 0.165925f
C1163 a_7208_47044# a_18970_45412# 0.230461f
C1164 a_10251_45454# a_10111_45776# 0.152168f
C1165 a_9973_46526# a_10224_45982# 0.15794f
C1166 a_19633_43262# a_20049_43262# 0.334778f
C1167 a_5655_43780# a_8659_44324# 0.270599f
C1168 a_14587_47614# VDD 0.264721f
C1169 COMP_N VDD 1.7049f
C1170 a_14950_43958# a_12127_46744# 0.950188f
C1171 a_13715_43780# a_14757_43806# 0.10314f
C1172 VIN_N VCM 1.69426f
C1173 a_12379_44350# a_12683_43433# 0.11018f
C1174 a_6105_44894# a_6455_44894# 0.218541f
C1175 a_5939_44894# a_7020_44894# 0.102355f
C1176 a_14573_47070# VDD 0.316031f
C1177 EN_VIN_BSTR_N C9_N_btm 0.226586f
C1178 C2_P_btm C1_P_btm 5.10246f
C1179 C3_P_btm C0_P_btm 0.409922f
C1180 C4_P_btm C0_dummy_P_btm 0.116511f
C1181 EN_VIN_BSTR_P VDD 0.92857f
C1182 a_82_45670# a_1735_46195# 0.198691f
C1183 a_3320_46134# VDD 0.273551f
C1184 a_2443_43806# a_2959_43806# 0.104514f
C1185 a_15079_46134# a_14955_45982# 0.153663f
C1186 a_18449_44324# VDD 0.205113f
C1187 a_10251_45454# a_14647_43494# 0.15515f
C1188 a_n2472_43236# VDD 0.289269f
C1189 a_10150_47322# VDD 0.279005f
C1190 a_22775_42718# VDD 0.425541f
C1191 a_n172_44582# a_1387_44582# 0.106794f
C1192 a_5663_45982# a_6196_46250# 0.305381f
C1193 a_9349_46539# a_9547_46565# 0.36083f
C1194 a_16291_46758# VDD 0.207388f
C1195 a_n2293_44332# VDD 0.473468f
C1196 a_11507_47833# RST_Z 0.208697f
C1197 a_12887_47833# VDD 0.234784f
C1198 a_n1237_42718# VDD 0.206895f
C1199 VIN_P VCM 1.69434f
C1200 VIN_N VREF 2.15636f
C1201 a_5916_43806# VDD 0.284617f
C1202 a_6105_44894# a_6673_45136# 0.171912f
C1203 C3_P_btm C1_P_btm 7.588649f
C1204 C4_P_btm C0_P_btm 0.138615f
C1205 C5_P_btm C0_dummy_P_btm 0.117097f
C1206 a_82_45670# a_1431_45982# 0.150693f
C1207 a_2512_45982# VDD 0.296164f
C1208 a_2627_42718# a_2609_43806# 0.271694f
C1209 a_16579_43566# a_16404_43640# 0.234322f
C1210 a_6631_44582# a_7415_44466# 0.293733f
C1211 a_17881_44356# VDD 0.568453f
C1212 a_n2840_43236# VDD 0.292205f
C1213 a_9947_47044# VDD 0.346007f
C1214 a_15582_45982# a_15879_47320# 0.133998f
C1215 a_22223_42718# VDD 0.290006f
C1216 a_22469_41061# a_22521_39947# 0.65678f
C1217 a_22521_40491# a_22459_39581# 0.129251f
C1218 a_5663_45982# a_5655_43780# 0.222017f
C1219 a_9349_46539# a_9293_46565# 0.202007f
C1220 a_15309_45438# VDD 0.199747f
C1221 a_21755_44350# a_22031_44350# 0.164707f
C1222 a_82_45670# a_361_45438# 0.388322f
C1223 a_n2661_44332# VDD 0.500568f
C1224 a_15328_46134# a_16085_45982# 0.144398f
C1225 a_11299_47832# RST_Z 0.165956f
C1226 a_11507_47833# VDD 0.245864f
C1227 a_5847_47614# DATA[4] 0.354723f
C1228 COMP_P VDD 1.12332f
C1229 VIN_P VREF 3.95249f
C1230 a_9304_43494# a_9416_43530# 0.229048f
C1231 a_5419_47258# a_8055_45491# 0.117119f
C1232 a_12121_45956# VDD 0.234975f
C1233 a_10684_45670# a_11017_45736# 0.20918f
C1234 a_18766_43236# a_19633_43262# 0.789069f
C1235 a_6091_43780# VDD 0.478158f
C1236 a_16513_42718# a_16703_42718# 0.23663f
C1237 a_5939_44894# a_6455_44894# 0.102974f
C1238 EN_VIN_BSTR_N C7_N_btm 0.115875f
C1239 a_22469_41061# VCM 0.151816f
C1240 C3_P_btm C2_P_btm 5.69083f
C1241 C5_P_btm C0_P_btm 0.138379f
C1242 C4_P_btm C1_P_btm 0.128431f
C1243 C6_P_btm C0_dummy_P_btm 0.122824f
C1244 a_7208_47044# a_13181_45982# 0.683409f
C1245 a_2687_45956# VDD 0.356034f
C1246 a_2443_43806# a_2609_43806# 0.682512f
C1247 a_15079_46134# a_15328_46134# 0.167707f
C1248 a_17715_44356# VDD 0.444367f
C1249 a_15691_47436# a_15879_47320# 0.141213f
C1250 a_9395_47044# VDD 0.321529f
C1251 a_22521_41035# a_22521_39947# 0.365591f
C1252 a_n60_44618# a_161_44648# 0.135748f
C1253 a_n172_44582# a_570_44324# 0.280446f
C1254 a_14757_45982# VDD 0.432514f
C1255 a_82_45670# a_656_45670# 0.2145f
C1256 a_n2661_44868# VDD 0.647169f
C1257 a_15328_46134# a_14955_45982# 0.126962f
C1258 a_3328_44324# VDD 0.14565f
C1259 a_n1085_47874# a_n749_47846# 0.224669f
C1260 a_11299_47832# VDD 0.149784f
C1261 SMPL_ON_N a_21789_35634# 0.39925f
C1262 a_11788_46134# VDD 0.844546f
C1263 a_10684_45670# a_10389_45438# 0.134085f
C1264 a_5351_43806# VDD 0.21035f
C1265 a_6243_45107# a_6105_44894# 0.211344f
C1266 EN_VIN_BSTR_N C6_N_btm 0.118916f
C1267 C6_P_btm C0_P_btm 0.139432f
C1268 C5_P_btm C1_P_btm 0.127667f
C1269 C4_P_btm C2_P_btm 7.37802f
C1270 C7_P_btm C0_dummy_P_btm 0.12244f
C1271 a_n1586_35608# VDD 0.373377f
C1272 a_1947_45982# VDD 0.194091f
C1273 a_2443_43806# a_2627_42718# 0.14367f
C1274 a_16670_44324# VDD 0.348099f
C1275 a_8391_47044# VDD 0.426657f
C1276 a_21855_42718# VDD 0.254469f
C1277 a_22469_41061# a_22459_39581# 0.245891f
C1278 a_n172_44582# a_161_44648# 0.231693f
C1279 a_22031_45438# a_22959_44358# 0.17985f
C1280 a_15192_46500# VDD 0.184577f
C1281 a_5663_45982# a_5715_45956# 0.114408f
C1282 a_7208_47044# a_13715_43780# 0.188721f
C1283 a_1736_43276# VDD 1.98805f
C1284 a_n2661_44868# a_n2293_44868# 0.191136f
C1285 a_11143_47588# VDD 0.236935f
C1286 a_n1552_42692# VDD 0.236103f
C1287 a_11183_44350# a_11671_44019# 0.113951f
C1288 a_18879_43780# a_18704_43806# 0.234322f
C1289 a_10684_45670# a_10588_45670# 0.319682f
C1290 a_15187_44868# a_15468_45412# 0.105091f
C1291 a_5569_44048# VDD 0.205813f
C1292 a_5939_44894# a_6105_44894# 0.575906f
C1293 a_4908_45956# VDD 0.91969f
C1294 EN_VIN_BSTR_N C5_N_btm 0.115337f
C1295 CAL_N VCM 1.57021f
C1296 C6_P_btm C1_P_btm 0.127984f
C1297 C7_P_btm C0_P_btm 0.141209f
C1298 C4_P_btm C3_P_btm 7.944839f
C1299 C5_P_btm C2_P_btm 0.138263f
C1300 C8_P_btm C0_dummy_P_btm 0.237239f
C1301 a_n2038_35608# VDD 0.522811f
C1302 a_17531_44894# a_17881_44356# 0.223452f
C1303 a_2165_46224# VDD 0.208745f
C1304 a_15489_43268# a_16404_43640# 0.118759f
C1305 a_n749_47846# a_n447_47044# 0.104387f
C1306 a_16211_44582# VDD 0.201859f
C1307 a_15329_47044# a_15879_47320# 0.13383f
C1308 a_7839_47222# VDD 0.218287f
C1309 a_22521_41035# a_22459_39581# 1.41583f
C1310 a_n172_44582# a_n60_44618# 0.264935f
C1311 a_14658_46526# VDD 0.282433f
C1312 a_82_45670# a_83_45776# 0.124413f
C1313 a_2134_44324# VDD 0.353194f
C1314 a_10415_47846# VDD 0.208411f
C1315 a_4651_47614# DATA[3] 0.348453f
C1316 a_3754_39964# VDAC_Pi 0.296508f
C1317 a_4322_46134# a_5382_44582# 0.272648f
C1318 a_5001_43806# VDD 0.273682f
C1319 a_5939_44894# a_6243_45107# 0.16171f
C1320 EN_VIN_BSTR_N C4_N_btm 0.116925f
C1321 C6_P_btm C2_P_btm 0.137649f
C1322 C7_P_btm C1_P_btm 0.128768f
C1323 C8_P_btm C0_P_btm 0.146681f
C1324 C5_P_btm C3_P_btm 0.135784f
C1325 C9_P_btm C0_dummy_P_btm 0.112646f
C1326 a_17531_44894# a_17715_44356# 0.215128f
C1327 a_1597_45982# VDD 0.361411f
C1328 a_15323_43268# a_16404_43640# 0.102355f
C1329 a_16057_43236# a_15839_43640# 0.209641f
C1330 a_15443_44582# VDD 0.180102f
C1331 a_22959_43806# VDD 0.304494f
C1332 a_5784_44364# a_6631_42883# 0.109681f
C1333 a_21303_42718# VDD 0.234525f
C1334 a_n268_44582# a_n60_44618# 0.18948f
C1335 a_22031_45438# a_21755_44350# 0.138756f
C1336 a_14470_46526# VDD 0.197468f
C1337 a_8483_46830# a_8308_46904# 0.233657f
C1338 a_12683_43433# a_12545_43268# 0.217668f
C1339 a_1387_45670# VDD 0.128707f
C1340 a_1488_43236# a_1339_43315# 0.167531f
C1341 a_5473_43582# a_5663_42718# 0.175134f
C1342 SMPL_ON_P VIN_P 0.537806f
C1343 a_n1920_42692# VDD 0.289765f
C1344 a_2113_38308# VDAC_Pi 0.170908f
C1345 a_5441_46500# a_5382_44582# 0.161119f
C1346 a_13561_44350# a_13725_44350# 0.146896f
C1347 a_4835_43806# VDD 0.438935f
C1348 a_13715_43780# a_14204_44350# 0.364696f
C1349 a_12747_47070# VDD 0.228651f
C1350 VDAC_P VCM 9.97461f
C1351 EN_VIN_BSTR_N C3_N_btm 0.100325f
C1352 C6_P_btm C3_P_btm 0.13406f
C1353 C7_P_btm C2_P_btm 0.138838f
C1354 C5_P_btm C4_P_btm 16.137598f
C1355 C9_P_btm C0_P_btm 0.144582f
C1356 C8_P_btm C1_P_btm 0.12931f
C1357 C10_P_btm C0_dummy_P_btm 0.397081f
C1358 a_12127_46744# a_16291_44914# 0.752857f
C1359 a_1735_46195# VDD 0.433052f
C1360 a_15489_43268# a_15839_43640# 0.21686f
C1361 a_2655_42870# a_2801_42968# 0.171361f
C1362 a_15221_47044# a_15582_45982# 0.200706f
C1363 a_3726_37500# CAL_P 0.102027f
C1364 a_n268_44582# a_n172_44582# 0.318161f
C1365 a_12683_43433# a_12379_43268# 0.314205f
C1366 a_989_45736# VDD 0.141508f
C1367 a_9973_46526# a_9969_45982# 0.261632f
C1368 a_2535_45670# a_2151_45670# 0.114727f
C1369 SMPL_ON_P a_n1605_47614# 0.197768f
C1370 a_9863_47874# VDD 0.369394f
C1371 EN_COMP VDD 1.0311f
C1372 a_2684_37794# VDAC_Pi 0.133177f
C1373 SMPL RST_Z 0.667857f
C1374 a_n2293_43780# a_n2661_43780# 0.168132f
C1375 a_171_44019# a_546_43100# 0.255712f
C1376 a_5441_46500# a_4322_46134# 0.107082f
C1377 a_19566_45670# a_19555_42718# 0.109084f
C1378 a_17789_43806# a_18704_43806# 0.118759f
C1379 a_17515_43806# a_18044_43806# 0.157595f
C1380 a_2075_42870# VDD 0.434186f
C1381 EN_VIN_BSTR_N C2_N_btm 0.118072f
C1382 C6_P_btm C4_P_btm 0.14422f
C1383 C7_P_btm C3_P_btm 0.13519f
C1384 C9_P_btm C1_P_btm 0.130686f
C1385 C8_P_btm C2_P_btm 0.139221f
C1386 C10_P_btm C0_P_btm 0.230054f
C1387 a_1431_45982# VDD 0.39929f
C1388 a_13266_45412# VDD 0.339343f
C1389 a_16291_44914# a_15187_44868# 0.219325f
C1390 a_15323_43268# a_15839_43640# 0.107482f
C1391 a_15489_43268# a_16057_43236# 0.181217f
C1392 a_16291_44914# a_18495_44868# 0.236508f
C1393 a_14133_43780# VDD 0.731541f
C1394 a_22591_43806# VDD 0.279529f
C1395 a_6635_47044# VDD 0.242658f
C1396 a_22521_41035# a_22469_41061# 1.99154f
C1397 a_21027_42718# VDD 0.260436f
C1398 a_361_45438# VDD 0.206258f
C1399 a_9973_46526# a_9803_45982# 0.161044f
C1400 a_n2661_44868# a_n2840_44868# 0.180889f
C1401 a_10588_45670# a_10389_45438# 0.206051f
C1402 a_2351_47614# DATA[2] 0.352341f
C1403 a_7595_47614# VDD 0.411688f
C1404 SMPL VDD 1.99499f
C1405 a_n2293_43780# a_n2293_43244# 0.279555f
C1406 a_7208_47044# a_16291_44914# 0.238558f
C1407 a_4035_45609# a_3897_45444# 0.230321f
C1408 a_18357_44048# a_18139_43806# 0.209641f
C1409 a_17623_43806# a_18704_43806# 0.102355f
C1410 a_8483_43780# a_8308_43806# 0.234322f
C1411 a_7319_43262# a_7648_43806# 0.158898f
C1412 VDAC_N VCM 9.97552f
C1413 EN_VIN_BSTR_N C1_N_btm 0.110046f
C1414 C6_P_btm C5_P_btm 18.5121f
C1415 C7_P_btm C4_P_btm 0.145744f
C1416 C9_P_btm C2_P_btm 0.140712f
C1417 C8_P_btm C3_P_btm 0.13458f
C1418 C10_P_btm C1_P_btm 0.182095f
C1419 a_12684_45276# VDD 1.66726f
C1420 a_6631_44582# a_7372_45670# 0.11084f
C1421 a_22223_43494# VDD 0.3214f
C1422 a_5749_47222# VDD 0.420798f
C1423 a_7393_46532# a_8308_46904# 0.118423f
C1424 a_656_45670# VDD 0.67087f
C1425 a_10111_45776# a_10389_45438# 0.110359f
C1426 a_7311_47614# VDD 0.284832f
C1427 a_n2288_42692# VDD 0.285197f
C1428 a_4527_46830# a_4322_46134# 0.392881f
C1429 a_n2293_43244# a_n2073_43806# 0.207813f
C1430 a_4035_45609# a_3731_45444# 0.3262f
C1431 a_10427_46348# VDD 0.132317f
C1432 a_17789_43806# a_18139_43806# 0.216297f
C1433 a_6563_45260# VDD 0.142103f
C1434 a_22959_43270# VDD 0.301579f
C1435 EN_VIN_BSTR_N C0_N_btm 0.12803f
C1436 C7_P_btm C5_P_btm 0.151868f
C1437 C9_P_btm C3_P_btm 0.135794f
C1438 C8_P_btm C4_P_btm 0.144911f
C1439 C10_P_btm C2_P_btm 0.193308f
C1440 VDAC_P VIN_P 0.239029f
C1441 a_16824_45276# a_16670_44324# 0.120875f
C1442 a_4651_44350# a_4733_44350# 0.171361f
C1443 a_4908_45956# a_5129_45956# 0.159289f
C1444 a_12438_45412# VDD 0.301165f
C1445 a_15323_43268# a_15489_43268# 0.894542f
C1446 a_22087_43244# VDD 0.319982f
C1447 a_15221_47044# a_15329_47044# 0.959048f
C1448 a_5419_47258# VDD 0.7238f
C1449 a_20383_42718# VDD 0.292509f
C1450 a_7961_46500# a_7743_46904# 0.209641f
C1451 a_9947_47044# a_7208_47044# 0.119479f
C1452 a_6951_47070# VDD 0.642794f
C1453 a_n2833_42692# VDD 0.445057f
C1454 a_171_44019# a_n60_44618# 0.111907f
C1455 a_636_42870# a_546_43100# 0.412608f
C1456 a_n60_44618# a_2043_43958# 0.109407f
C1457 a_17789_43806# a_18357_44048# 0.181217f
C1458 a_17623_43806# a_18139_43806# 0.110532f
C1459 a_22223_43270# VDD 0.223567f
C1460 C9_P_btm C4_P_btm 0.148287f
C1461 C8_P_btm C5_P_btm 0.144827f
C1462 C7_P_btm C6_P_btm 20.7485f
C1463 CAL_P RST_Z 0.551822f
C1464 VDAC_N VIN_N 0.240454f
C1465 a_22609_38842# VDD 0.317066f
C1466 C10_P_btm C3_P_btm 0.1871f
C1467 a_7208_47044# a_12121_45956# 0.133182f
C1468 a_6235_46124# a_7016_46231# 0.169139f
C1469 a_6391_46219# a_6322_46348# 0.209641f
C1470 a_3165_45982# a_2535_45670# 0.261028f
C1471 a_3576_44364# a_4791_42883# 0.109162f
C1472 a_6631_44582# a_6491_44716# 0.144307f
C1473 a_16291_44914# a_14204_44350# 0.368966f
C1474 a_21847_43806# VDD 0.417955f
C1475 a_15113_47222# a_15329_47044# 0.119807f
C1476 a_5089_47044# VDD 0.195754f
C1477 a_19555_42718# VDD 0.261178f
C1478 a_7393_46532# a_7743_46904# 0.21686f
C1479 a_7227_46532# a_8308_46904# 0.102325f
C1480 a_22591_43958# a_22591_43806# 0.213024f
C1481 a_83_45776# VDD 0.200318f
C1482 a_n381_43433# VDD 0.829526f
C1483 a_13654_46032# a_14382_46348# 0.14396f
C1484 a_16475_45412# a_10251_45454# 0.112019f
C1485 a_5847_47614# VDD 0.41489f
C1486 a_636_42870# a_570_44324# 0.209407f
C1487 a_4527_46830# a_4352_46904# 0.234322f
C1488 a_7393_43806# a_8308_43806# 0.125324f
C1489 a_12931_44894# VDD 0.405145f
C1490 a_4987_45742# a_4812_45816# 0.233657f
C1491 a_3067_44172# VDD 0.142196f
C1492 a_16475_45412# a_19037_42718# 0.137012f
C1493 a_21908_43236# VDD 0.224212f
C1494 a_5655_43780# a_9343_43806# 0.209102f
C1495 C10_P_btm C4_P_btm 0.273376f
C1496 CAL_P VDD 22.6485f
C1497 C8_P_btm C6_P_btm 0.162414f
C1498 C9_P_btm C5_P_btm 0.146663f
C1499 a_7208_47044# a_11788_46134# 0.196149f
C1500 a_215_46348# VDD 0.144089f
C1501 a_12623_43780# a_12448_43806# 0.234322f
C1502 a_6196_46250# a_7016_46231# 0.221177f
C1503 a_2627_43262# a_2709_43262# 0.171361f
C1504 a_15468_45412# a_15605_45438# 0.126609f
C1505 a_15113_47222# a_15221_47044# 0.106465f
C1506 a_9517_46539# a_9547_46565# 0.228665f
C1507 a_4993_47044# VDD 0.909253f
C1508 a_7393_46532# a_7961_46500# 0.181217f
C1509 a_n377_45776# VDD 0.218781f
C1510 a_16291_44914# a_17763_44868# 0.264924f
C1511 a_n2661_43780# VDD 0.824738f
C1512 a_13654_46032# a_14194_46348# 0.17174f
C1513 a_5839_47070# VDD 0.497065f
C1514 a_n2661_43780# a_n2840_43780# 0.180219f
C1515 a_18689_45412# a_18879_45956# 0.117588f
C1516 a_11692_46134# VDD 0.100434f
C1517 a_7961_44048# a_7743_43806# 0.209641f
C1518 a_17623_43806# a_17789_43806# 0.856458f
C1519 a_12436_44868# VDD 0.103776f
C1520 a_21719_43244# VDD 0.496877f
C1521 a_16475_45412# a_18445_42718# 0.631062f
C1522 a_5655_43780# a_8308_43806# 0.254973f
C1523 a_18689_45412# VDD 0.8396f
C1524 C10_P_btm C5_P_btm 0.236062f
C1525 C8_P_btm C7_P_btm 23.997501f
C1526 C9_P_btm C6_P_btm 0.155878f
C1527 a_5536_44324# a_5387_44403# 0.167531f
C1528 a_6235_46124# a_6391_46219# 0.108815f
C1529 a_3320_46134# a_2535_45670# 0.102168f
C1530 a_6196_46250# a_6322_46348# 0.170582f
C1531 a_22276_45412# a_22455_45420# 0.180033f
C1532 a_15005_47222# a_15221_47044# 0.134523f
C1533 a_9517_46539# a_9293_46565# 0.1014f
C1534 a_19187_42718# VDD 0.213892f
C1535 a_7227_46532# a_7743_46904# 0.110532f
C1536 a_n2293_43244# VDD 0.563734f
C1537 a_380_47222# a_713_47044# 0.229444f
C1538 a_663_47874# DATA[1] 0.332128f
C1539 a_2684_37794# a_2113_38308# 0.468006f
C1540 a_4651_47614# VDD 0.463603f
C1541 a_636_42870# a_n60_44618# 0.270172f
C1542 a_n61_46526# VDD 0.144346f
C1543 a_17927_46195# a_18044_45982# 0.170138f
C1544 a_10884_45982# VDD 0.27228f
C1545 a_7393_43806# a_7743_43806# 0.229804f
C1546 a_7227_43806# a_8308_43806# 0.102355f
C1547 a_17515_43806# a_17789_43806# 0.302154f
C1548 a_7648_46134# a_7981_45956# 0.374822f
C1549 a_9943_45046# VDD 0.135644f
C1550 a_21540_43236# VDD 0.310006f
C1551 a_5655_43780# a_8483_43780# 0.397656f
C1552 a_10251_45454# VDD 1.54728f
C1553 C10_P_btm C6_P_btm 0.317819f
C1554 C9_P_btm C7_P_btm 0.206278f
C1555 a_672_45982# VDD 0.289648f
C1556 a_6196_46250# a_6391_46219# 0.222728f
C1557 a_5655_43780# a_6322_46348# 0.164709f
C1558 a_5784_44364# a_5387_44403# 0.159011f
C1559 a_12683_43433# VDD 0.434946f
C1560 a_15005_47222# a_15113_47222# 0.126434f
C1561 a_5663_45982# a_4908_45956# 0.124459f
C1562 a_9517_46539# a_9349_46539# 0.140592f
C1563 a_4704_47044# VDD 0.151144f
C1564 a_19037_42718# VDD 0.952658f
C1565 a_7503_45982# a_7393_46532# 0.266197f
C1566 a_n2472_45412# VDD 0.278172f
C1567 a_13661_46298# a_13654_46032# 0.124623f
C1568 a_n2661_43244# VDD 0.625982f
C1569 a_7000_47222# a_7208_47044# 0.188009f
C1570 a_4091_47070# VDD 0.926413f
C1571 a_636_42870# a_n172_44582# 0.14881f
C1572 a_3437_46532# a_4352_46904# 0.118759f
C1573 a_4908_45956# a_11335_46830# 0.11327f
C1574 a_7503_45982# a_6235_46124# 0.107145f
C1575 a_16291_44914# a_16921_46364# 0.1497f
C1576 a_11059_45956# VDD 0.340432f
C1577 a_7393_43806# a_7961_44048# 0.186387f
C1578 a_17515_43806# a_17623_43806# 0.378676f
C1579 a_8848_44868# VDD 0.141781f
C1580 a_3897_45444# a_4812_45816# 0.117156f
C1581 a_21197_42718# VDD 0.460612f
C1582 a_16475_45412# a_18759_42746# 0.191677f
C1583 a_5655_43780# a_7743_43806# 0.190047f
C1584 a_18530_47070# VDD 0.189054f
C1585 C10_P_btm C7_P_btm 0.521459f
C1586 a_22469_39973# VDD 0.361538f
C1587 C9_P_btm C8_P_btm 29.4361f
C1588 a_4651_44350# a_5139_44019# 0.113805f
C1589 a_847_45956# VDD 0.351674f
C1590 a_5655_43780# a_6391_46219# 0.154841f
C1591 a_6196_46250# a_6235_46124# 0.748414f
C1592 a_22031_44350# a_22959_43270# 0.180946f
C1593 a_3165_43262# a_3692_43628# 0.157662f
C1594 a_18445_42718# VDD 0.23244f
C1595 a_4061_47044# VDD 0.77553f
C1596 a_7227_46532# a_7393_46532# 0.883799f
C1597 a_18803_47070# a_18064_46642# 0.206294f
C1598 a_13427_46756# VDD 0.33754f
C1599 a_85_47070# a_713_47044# 0.104406f
C1600 a_2112_39137# a_2113_38308# 0.479143f
C1601 a_20283_43262# VDD 0.547443f
C1602 a_2351_47614# VDD 0.471111f
C1603 a_4005_46500# a_3787_46904# 0.209641f
C1604 a_n60_44618# a_33_43806# 0.307709f
C1605 a_10319_45982# VDD 0.192921f
C1606 a_7227_43806# a_7743_43806# 0.107482f
C1607 a_8379_46134# a_8651_45962# 0.13675f
C1608 a_7842_44868# VDD 0.23726f
C1609 a_4465_45412# a_4247_45816# 0.209641f
C1610 a_3731_45444# a_4812_45816# 0.102355f
C1611 a_3524_43806# VDD 0.295638f
C1612 a_19771_43600# VDD 0.216005f
C1613 a_5655_43780# a_7961_44048# 0.182764f
C1614 C10_P_btm C8_P_btm 0.607425f
C1615 a_22821_39429# VDD 0.432227f
C1616 a_17927_46195# VDD 0.482821f
C1617 EN_VIN_BSTR_P C0_P_btm 0.12803f
C1618 a_171_44019# a_288_43806# 0.170113f
C1619 a_107_45982# VDD 0.217937f
C1620 a_5655_43780# a_6235_46124# 0.304838f
C1621 a_13635_43566# a_13460_43640# 0.234322f
C1622 a_2167_46526# VDD 0.344304f
C1623 a_7227_46532# a_7503_45982# 0.168793f
C1624 a_18803_47070# a_18103_46768# 0.16233f
C1625 a_n2840_45412# VDD 0.289706f
C1626 a_13181_45982# a_14194_46348# 0.334357f
C1627 a_7839_47222# a_7760_45956# 0.110662f
C1628 a_n1085_47874# DATA[0] 0.333089f
C1629 a_20049_43262# VDD 1.34355f
C1630 a_2343_47070# VDD 0.502619f
C1631 a_3437_46532# a_3787_46904# 0.21686f
C1632 a_3271_46532# a_4352_46904# 0.102325f
C1633 a_13715_43780# a_13536_43780# 0.166329f
C1634 a_10447_44403# a_10844_44364# 0.155736f
C1635 a_16291_46758# a_16128_46134# 0.10013f
C1636 a_10537_46224# VDD 0.203945f
C1637 a_7319_43262# a_7393_43806# 0.220737f
C1638 a_10251_45454# a_17531_44894# 0.295391f
C1639 a_7020_44894# VDD 0.276426f
C1640 a_3897_45444# a_4247_45816# 0.206912f
C1641 a_3699_43780# VDD 0.493074f
C1642 a_19191_43262# VDD 0.184093f
C1643 C10_P_btm C9_P_btm 37.7035f
C1644 a_22545_39429# VDD 0.537013f
C1645 a_18133_47235# VDD 0.196538f
C1646 EN_VIN_BSTR_P C1_P_btm 0.110046f
C1647 a_325_46224# VDD 0.207826f
C1648 a_5918_46234# a_6235_46124# 0.102355f
C1649 a_11671_44019# VDD 0.629986f
C1650 VDAC_N VDAC_P 4.87144f
C1651 a_18759_42746# VDD 0.19724f
C1652 a_1431_47070# VDD 0.53748f
C1653 a_14573_47070# a_15079_46134# 0.107326f
C1654 a_13181_45982# a_13654_46032# 0.202937f
C1655 a_1387_44582# VDD 0.126597f
C1656 a_n194_47222# a_380_47222# 0.468641f
C1657 a_85_47070# a_n381_46697# 0.241069f
C1658 a_19274_43262# VDD 0.199134f
C1659 a_1209_47588# VDD 0.639113f
C1660 a_3437_46532# a_4005_46500# 0.181217f
C1661 a_10251_45454# a_17623_45982# 0.231468f
C1662 a_18259_46500# a_18190_46526# 0.209641f
C1663 a_1736_43276# a_1339_43315# 0.162652f
C1664 a_9969_45982# VDD 0.256145f
C1665 a_14133_43780# a_14301_44035# 0.136023f
C1666 a_7227_43806# a_7393_43806# 0.895425f
C1667 a_7195_44868# VDD 0.342003f
C1668 a_3897_45444# a_4465_45412# 0.17072f
C1669 a_3731_45444# a_4247_45816# 0.105988f
C1670 a_2959_43806# VDD 0.205367f
C1671 a_19003_43262# VDD 0.239804f
C1672 a_22521_39947# VDD 0.916455f
C1673 a_16703_45982# VDD 0.290362f
C1674 EN_VIN_BSTR_P C2_P_btm 0.118072f
C1675 a_n243_45982# VDD 0.600462f
C1676 a_5918_46234# a_6196_46250# 0.118759f
C1677 a_12683_43433# a_12800_43628# 0.168655f
C1678 SMPL_ON_N SMPL 2.53207f
C1679 a_18247_44172# VDD 0.132018f
C1680 a_546_43100# VDD 1.08464f
C1681 a_6631_44582# a_7319_43262# 0.102133f
C1682 a_999_47846# VDD 0.272872f
C1683 a_18348_43262# VDD 0.349722f
C1684 a_4908_45956# a_10383_46697# 0.172393f
C1685 a_3271_46532# a_3787_46904# 0.110532f
C1686 VDD VCM 8.287621f
C1687 a_6631_44582# a_5655_43780# 0.168237f
C1688 a_17927_46195# a_17789_45982# 0.613603f
C1689 a_13930_46842# a_13937_46602# 0.123819f
C1690 a_18064_46642# a_18190_46526# 0.170692f
C1691 a_9803_45982# VDD 0.458214f
C1692 a_14133_43780# a_14077_44133# 0.201055f
C1693 a_7227_43806# a_7319_43262# 0.169707f
C1694 a_6455_44894# VDD 0.199934f
C1695 a_3177_44048# VDD 0.210412f
C1696 a_18766_43236# VDD 0.391919f
C1697 a_12833_42718# a_13023_42718# 0.23961f
C1698 a_5655_43780# a_7227_43806# 0.537358f
C1699 a_16561_45982# VDD 0.374051f
C1700 EN_VIN_BSTR_P C3_P_btm 0.100325f
C1701 a_12127_46744# a_13457_46892# 0.692198f
C1702 a_n105_46195# VDD 0.393384f
C1703 a_5918_46234# a_5655_43780# 0.213109f
C1704 a_1736_43276# a_4239_42883# 0.108491f
C1705 a_12545_43268# a_13460_43640# 0.118759f
C1706 a_17671_42883# VDD 0.260436f
C1707 a_10684_45670# VDD 1.22514f
C1708 a_15443_44582# a_15589_44350# 0.171361f
C1709 a_570_44324# VDD 0.264111f
C1710 a_663_47874# VDD 0.432093f
C1711 SMPL_ON_P CLK_DATA 0.263144f
C1712 a_16102_47044# a_15582_45982# 0.122441f
C1713 a_5419_47258# a_5663_45982# 0.499285f
C1714 a_18093_43262# VDD 0.314927f
C1715 a_4908_45956# a_10079_46532# 0.36296f
C1716 a_3575_46697# a_3437_46532# 0.267414f
C1717 VDD VREF 9.84717f
C1718 a_17927_46195# a_17623_45982# 0.495626f
C1719 a_18064_46642# a_18259_46500# 0.206455f
C1720 a_14133_43780# a_14331_44133# 0.336679f
C1721 a_6673_45136# VDD 0.205844f
C1722 a_3731_45444# a_3897_45444# 0.72184f
C1723 a_2609_43806# VDD 0.552297f
C1724 a_16404_43640# VDD 0.279068f
C1725 a_636_42870# a_171_44019# 0.484794f
C1726 a_15879_47320# VDD 0.174839f
C1727 a_22459_39581# VDD 0.66988f
C1728 EN_VIN_BSTR_P C4_P_btm 0.116925f
C1729 a_636_42870# a_2043_43958# 0.121904f
C1730 a_n409_45982# VDD 0.457491f
C1731 a_1123_43780# a_948_43806# 0.234322f
C1732 a_5715_45956# a_5655_43780# 0.268513f
C1733 a_12379_43268# a_13460_43640# 0.102355f
C1734 a_13113_43236# a_12895_43640# 0.209641f
C1735 a_14950_43958# a_15415_44350# 0.108851f
C1736 a_14819_44582# VDD 0.126669f
C1737 a_9517_46539# a_9551_47203# 0.101174f
C1738 a_15133_43582# a_15008_42692# 0.176313f
C1739 a_20107_43806# VDD 0.459402f
C1740 a_1115_47044# VDD 0.238782f
C1741 a_16703_42718# VDD 0.236187f
C1742 a_10703_46526# VDD 0.142103f
C1743 a_5139_44019# a_5256_43806# 0.169472f
C1744 a_22959_45982# VDD 0.304443f
C1745 a_161_44648# VDD 0.179912f
C1746 a_8055_45491# a_8192_44874# 0.155836f
C1747 a_n749_47846# VDD 0.72849f
C1748 a_3271_46532# a_3437_46532# 0.880442f
C1749 a_10251_45454# a_12127_46744# 0.144261f
C1750 C10_N_btm VCM 10.2371f
C1751 VDD VIN_N 0.942438f
C1752 a_18103_46768# a_18259_46500# 0.105995f
C1753 a_5784_44364# a_5655_43780# 0.315575f
C1754 a_8379_46134# a_7648_46134# 0.121305f
C1755 a_6105_44894# VDD 0.510895f
C1756 a_2627_42718# VDD 0.585643f
C1757 a_16579_43566# VDD 0.464827f
C1758 a_15582_45982# VDD 0.428744f
C1759 a_22521_40491# VDD 1.05499f
C1760 EN_VIN_BSTR_P C5_P_btm 0.115337f
C1761 a_20064_35138# a_21789_35634# 0.150796f
C1762 a_7208_47044# a_11692_46134# 0.189453f
C1763 a_5715_45956# a_5918_46234# 0.233657f
C1764 a_1736_43276# a_3541_42718# 0.148428f
C1765 a_11415_45670# VDD 0.124265f
C1766 a_12545_43268# a_12895_43640# 0.20669f
C1767 a_14545_44569# VDD 0.204155f
C1768 a_18704_43806# VDD 0.272876f
C1769 a_428_42724# a_468_42870# 0.167531f
C1770 a_16111_45412# a_16287_45744# 0.185422f
C1771 a_7208_47044# a_18689_45412# 0.195542f
C1772 a_8530_39574# CAL_N 0.644218f
C1773 a_16513_42718# VDD 0.231163f
C1774 a_14950_43958# a_18103_46768# 0.50225f
C1775 a_571_43566# a_396_43640# 0.233657f
C1776 a_n60_44618# VDD 1.22676f
C1777 a_n1085_47874# VDD 0.41946f
C1778 a_5419_47258# a_7760_45956# 0.111363f
C1779 a_5382_44582# VDD 1.12495f
C1780 a_3271_46532# a_3575_46697# 0.169167f
C1781 C9_N_btm VCM 6.06251f
C1782 C10_N_btm VREF 14.776899f
C1783 VDD VIN_P 0.955108f
C1784 a_18103_46768# a_18064_46642# 0.576869f
C1785 a_7552_46134# a_7648_46134# 0.318706f
C1786 a_6243_45107# VDD 0.494612f
C1787 a_2443_43806# VDD 0.424358f
C1788 a_15839_43640# VDD 0.196785f
C1789 a_2471_45046# a_2617_45144# 0.171361f
C1790 a_15691_47436# VDD 0.243142f
C1791 EN_VIN_BSTR_P C6_P_btm 0.118916f
C1792 a_171_44019# a_33_43806# 0.758807f
C1793 a_11671_44019# a_11533_43806# 0.298912f
C1794 a_11017_45736# VDD 0.1384f
C1795 a_12379_43268# a_12895_43640# 0.102946f
C1796 a_12545_43268# a_13113_43236# 0.17072f
C1797 a_13725_44350# VDD 0.163289f
C1798 a_18879_43780# VDD 0.455477f
C1799 a_n193_47098# VDD 0.226328f
C1800 a_13151_45956# a_13181_45982# 0.342055f
C1801 a_n172_44582# VDD 0.737777f
C1802 a_n1605_47614# VDD 0.200166f
C1803 a_19633_43262# VDD 0.480707f
C1804 a_4908_45956# a_9349_46539# 0.209972f
C1805 a_4322_46134# VDD 1.82629f
C1806 VDD DEBUG_MUX[3] 0.126156f
C1807 C10_N_btm VIN_N 3.66108f
C1808 C8_N_btm VCM 2.61094f
C1809 C9_N_btm VREF 7.36949f
C1810 a_5419_47258# a_8204_45412# 0.153533f
C1811 a_17786_46658# a_18064_46642# 0.118759f
C1812 a_5939_44894# VDD 0.447912f
C1813 a_10844_44364# a_12427_42883# 0.109681f
C1814 a_n1429_43262# COMP_P 0.159541f
C1815 a_16057_43236# VDD 0.205742f
C1816 a_22469_41061# VDD 0.563604f
C1817 EN_VIN_BSTR_P C7_P_btm 0.115875f
C1818 a_171_44019# a_n133_43806# 0.617619f
C1819 a_14635_44324# a_14133_43780# 0.122967f
C1820 a_12427_46758# a_12699_46616# 0.13675f
C1821 a_n2472_45956# VDD 0.258378f
C1822 a_33_43806# a_948_43806# 0.11703f
C1823 a_11671_44019# a_11367_43806# 0.118652f
C1824 a_10389_45438# VDD 0.198302f
C1825 a_13561_44350# VDD 0.166885f
C1826 a_14587_47614# a_14757_47614# 0.108611f
C1827 a_18139_43806# VDD 0.192513f
C1828 a_n447_47044# VDD 0.425307f
C1829 a_15831_42883# VDD 0.270165f
C1830 a_22591_45982# VDD 0.292485f
C1831 a_n268_44582# VDD 0.148506f
C1832 SMPL_ON_P VDD 1.06867f
C1833 a_5441_46500# VDD 0.543353f
C1834 C9_N_btm VIN_N 1.8284f
C1835 C7_N_btm VCM 1.58335f
C1836 VDD DEBUG_MUX[2] 0.101099f
C1837 C8_N_btm VREF 3.6701f
C1838 a_17786_46658# a_18103_46768# 0.102355f
C1839 a_10251_45454# a_17951_44868# 0.194121f
C1840 a_2617_45144# VDD 0.192625f
C1841 a_15489_43268# VDD 0.25388f
C1842 a_15329_47044# VDD 0.166961f
C1843 a_22521_41035# VDD 0.802597f
C1844 a_601_44048# a_383_43806# 0.209641f
C1845 a_n133_43806# a_948_43806# 0.102325f
C1846 a_14757_45982# a_14382_46348# 0.141114f
C1847 a_12379_43268# a_12545_43268# 0.573172f
C1848 a_13023_44716# VDD 0.399413f
C1849 a_18357_44048# VDD 0.20366f
C1850 a_283_42692# a_428_42724# 0.113515f
C1851 a_n519_43268# a_396_43640# 0.125324f
C1852 a_n2472_44324# VDD 0.268754f
C1853 a_4352_46904# VDD 0.280034f
C1854 C8_N_btm VIN_N 0.907769f
C1855 C6_N_btm VCM 0.877241f
C1856 C7_N_btm VREF 1.818f
C1857 a_14658_46526# a_15033_46526# 0.131018f
C1858 a_17242_43806# a_17515_43806# 0.118466f
C1859 a_n1429_43262# a_n1552_42692# 0.186492f
C1860 a_15323_43268# VDD 0.397912f
C1861 a_15221_47044# VDD 0.14964f
C1862 EN_VIN_BSTR_N a_20064_35138# 0.573165f
C1863 CAL_N VDD 26.421099f
C1864 EN_VIN_BSTR_P C9_P_btm 0.226586f
C1865 a_12427_46758# a_10684_45670# 0.100381f
C1866 a_n2840_45956# VDD 0.302566f
C1867 a_33_43806# a_383_43806# 0.216095f
C1868 a_16824_45276# a_17671_42883# 0.109681f
C1869 a_18689_45412# a_17763_44868# 0.100343f
C1870 a_10111_45776# VDD 0.210601f
C1871 a_5663_45982# a_7842_44868# 0.126374f
C1872 a_12379_44350# VDD 0.265901f
C1873 a_12887_47833# a_9551_47203# 0.108584f
C1874 a_17789_43806# VDD 0.249687f
C1875 a_15008_42692# VDD 0.293782f
C1876 a_3726_37500# a_6886_37412# 0.702909f
C1877 a_5139_44019# a_5001_43806# 0.308636f
C1878 a_21755_44350# a_22223_44358# 0.173482f
C1879 a_n685_43268# a_396_43640# 0.101963f
C1880 a_49_43236# a_n169_43640# 0.209641f
C1881 a_16291_44914# a_18282_45670# 0.221561f
C1882 a_n2840_44324# VDD 0.289706f
C1883 a_10467_47212# a_11248_47319# 0.157453f
C1884 a_15437_47044# a_15691_47436# 0.259284f
C1885 a_10623_47307# a_10554_47436# 0.209641f
C1886 a_n1920_47588# VDD 0.230743f
C1887 a_n2833_47874# CLK_DATA 0.33085f
C1888 a_4527_46830# VDD 0.462001f
C1889 C7_N_btm VIN_N 1.52459f
C1890 C5_N_btm VCM 0.719982f
C1891 C6_N_btm VREF 1.41944f
C1892 a_17583_46500# a_17786_46658# 0.233657f
C1893 a_7981_45956# VDD 0.156459f
C1894 a_491_44172# VDD 0.132148f
C1895 a_14647_43494# VDD 0.20962f
C1896 a_1663_45046# a_1935_44874# 0.13675f
C1897 a_2471_45046# a_171_44019# 0.119778f
C1898 a_15113_47222# VDD 0.170889f
C1899 EN_VIN_BSTR_N a_19320_35138# 0.653211f
C1900 VDAC_P RST_Z 0.158793f
C1901 EN_VIN_BSTR_P C10_P_btm 0.320716f
C1902 a_3576_44364# a_3882_44324# 0.128115f
C1903 a_6243_45107# a_6519_43494# 0.109781f
C1904 a_n133_43806# a_383_43806# 0.105995f
C1905 a_33_43806# a_601_44048# 0.17072f
C1906 a_1735_46195# a_1852_45982# 0.157972f
C1907 a_10251_45454# a_17763_44868# 0.347443f
C1908 a_11183_44350# VDD 0.212579f
C1909 a_17623_43806# VDD 0.402554f
C1910 a_n2104_47044# VDD 0.29454f
C1911 a_7754_38470# VDAC_N 0.110573f
C1912 a_8530_39574# a_6886_37412# 0.616015f
C1913 a_22123_44894# a_22591_44894# 0.179973f
C1914 a_5139_44019# a_4835_43806# 0.213794f
C1915 a_n519_43268# a_n169_43640# 0.219633f
C1916 a_10428_47338# a_11248_47319# 0.202821f
C1917 a_15947_43262# VDD 0.132317f
C1918 a_3787_46904# VDD 0.195983f
C1919 C6_N_btm VIN_N 0.391985f
C1920 C4_N_btm VCM 0.716447f
C1921 C5_N_btm VREF 0.987144f
C1922 a_16291_44914# a_18064_46642# 0.130967f
C1923 a_7648_46134# VDD 0.74622f
C1924 a_9551_47203# a_9395_47044# 0.232491f
C1925 a_13460_43640# VDD 0.278505f
C1926 a_5655_43780# a_5916_43806# 0.229916f
C1927 a_15005_47222# VDD 0.390929f
C1928 VDAC_P VDD 5.16188f
C1929 a_3165_45982# a_4700_46134# 0.100857f
C1930 a_8850_45412# VDD 0.342392f
C1931 a_10844_44364# VDD 0.814057f
C1932 a_104_42692# a_283_42692# 0.176024f
C1933 a_17515_43806# VDD 0.324214f
C1934 a_13991_42883# VDD 0.278333f
C1935 a_7754_38470# a_6886_37412# 0.180842f
C1936 a_22123_44894# a_22399_44894# 0.138665f
C1937 VCM VSS 22.07842f
C1938 VREF VSS 17.869415f
C1939 VIN_N VSS 17.048048f
C1940 VIN_P VSS 16.52358f
C1941 DEBUG_MUX[3] VSS 0.520798f
C1942 DEBUG_MUX[2] VSS 0.396995f
C1943 DEBUG_MUX[1] VSS 0.41791f
C1944 DEBUG_MUX[0] VSS 0.457552f
C1945 EN_OFFSET_CAL VSS 0.425939f
C1946 DEBUG_OUT VSS 0.613768f
C1947 DATA[5] VSS 0.684062f
C1948 DATA[4] VSS 0.671412f
C1949 DATA[3] VSS 1.12992f
C1950 DATA[2] VSS 0.7311f
C1951 DATA[1] VSS 0.70246f
C1952 DATA[0] VSS 0.502377f
C1953 CLK_DATA VSS 0.417892f
C1954 START VSS 0.499328f
C1955 CLK VSS 0.516784f
C1956 RST_Z VSS 15.835025f
C1957 VDD VSS 0.696667p
C1958 C10_N_btm VSS 0.276046p
C1959 C9_N_btm VSS 0.120738p
C1960 C8_N_btm VSS 63.980186f
C1961 C7_N_btm VSS 35.240353f
C1962 C6_N_btm VSS 20.613462f
C1963 C5_N_btm VSS 13.73659f
C1964 C4_N_btm VSS 11.615809f
C1965 C3_N_btm VSS 9.62813f
C1966 C2_N_btm VSS 9.169419f
C1967 C1_N_btm VSS 8.6589f
C1968 C0_N_btm VSS 9.241811f
C1969 C0_dummy_N_btm VSS 8.066401f
C1970 C0_dummy_P_btm VSS 8.047689f
C1971 C0_P_btm VSS 9.274731f
C1972 C1_P_btm VSS 8.695661f
C1973 C2_P_btm VSS 9.18044f
C1974 C3_P_btm VSS 9.64071f
C1975 C4_P_btm VSS 11.60488f
C1976 C5_P_btm VSS 13.73231f
C1977 C6_P_btm VSS 20.60929f
C1978 C7_P_btm VSS 35.236233f
C1979 C8_P_btm VSS 63.976162f
C1980 C9_P_btm VSS 0.120729p
C1981 C10_P_btm VSS 0.276064p
C1982 a_21789_35634# VSS 0.737759f
C1983 a_20064_35138# VSS 1.74491f
C1984 a_19320_35138# VSS 1.696f
C1985 EN_VIN_BSTR_N VSS 10.286273f
C1986 a_n283_35174# VSS 1.73472f
C1987 EN_VIN_BSTR_P VSS 10.516015f
C1988 a_n1586_35608# VSS 1.7452f
C1989 a_n2038_35608# VSS 0.738209f
C1990 a_22609_38426# VSS 0.48998f
C1991 a_22609_38842# VSS 0.519727f
C1992 CAL_P VSS 11.382667f
C1993 a_22469_39973# VSS 2.78847f
C1994 a_22821_39429# VSS 0.551882f
C1995 a_22545_39429# VSS 0.354928f
C1996 a_22521_39947# VSS 1.85573f
C1997 a_22459_39581# VSS 2.1545f
C1998 a_22521_40491# VSS 1.21462f
C1999 a_22469_41061# VSS 1.7314f
C2000 a_22521_41035# VSS 1.84244f
C2001 CAL_N VSS 9.044225f
C2002 VDAC_P VSS 80.75824f
C2003 VDAC_N VSS 81.33162f
C2004 a_6886_37412# VSS 3.84703f
C2005 a_3726_37500# VSS 4.50043f
C2006 a_8530_39574# VSS 2.76322f
C2007 a_7754_38470# VSS 3.24669f
C2008 VDAC_Ni VSS 3.07659f
C2009 a_7754_38636# VSS 0.353706f
C2010 a_3754_38802# VSS 0.390074f
C2011 a_7754_38968# VSS 0.330037f
C2012 a_3754_39134# VSS 0.401983f
C2013 a_7754_39300# VSS 0.330682f
C2014 a_3754_39466# VSS 0.401172f
C2015 a_7754_39632# VSS 0.340942f
C2016 VDAC_Pi VSS 3.946915f
C2017 a_7754_39964# VSS 2.62481f
C2018 a_3754_39964# VSS 0.671366f
C2019 a_2113_38308# VSS 2.64406f
C2020 a_2684_37794# VSS 0.414596f
C2021 a_1177_38525# VSS 0.64211f
C2022 a_2112_39137# VSS 0.414253f
C2023 a_1239_39043# VSS 0.613805f
C2024 a_1239_39587# VSS 0.634479f
C2025 a_22465_38541# VSS 1.85672f
C2026 a_22400_42718# VSS 2.20472f
C2027 a_22775_42718# VSS 0.598102f
C2028 a_22223_42718# VSS 0.35376f
C2029 a_21855_42718# VSS 0.330415f
C2030 a_21303_42718# VSS 0.305065f
C2031 a_21027_42718# VSS 0.254456f
C2032 a_20383_42718# VSS 0.381474f
C2033 a_19555_42718# VSS 0.264139f
C2034 a_19187_42718# VSS 0.295422f
C2035 a_19037_42718# VSS 0.556866f
C2036 a_18445_42718# VSS 0.354312f
C2037 a_18759_42746# VSS 0.236318f
C2038 a_17671_42883# VSS 0.275069f
C2039 a_16703_42718# VSS 0.354618f
C2040 a_16513_42718# VSS 0.313719f
C2041 a_15831_42883# VSS 0.26686f
C2042 a_15008_42692# VSS 0.358583f
C2043 a_13991_42883# VSS 0.268554f
C2044 a_13023_42718# VSS 0.356024f
C2045 a_12833_42718# VSS 0.316542f
C2046 a_12427_42883# VSS 0.253f
C2047 a_11599_42883# VSS 0.260716f
C2048 a_11183_42718# VSS 0.326381f
C2049 a_10901_42718# VSS 0.351974f
C2050 a_9987_42968# VSS 0.369438f
C2051 a_9343_42718# VSS 0.336174f
C2052 a_8423_42718# VSS 0.292932f
C2053 a_7556_42692# VSS 0.362489f
C2054 a_6631_42883# VSS 0.268954f
C2055 a_5663_42718# VSS 0.373241f
C2056 a_4791_42883# VSS 0.269936f
C2057 a_4239_42883# VSS 0.243224f
C2058 a_3823_42718# VSS 0.328502f
C2059 a_3541_42718# VSS 0.318534f
C2060 a_2655_42870# VSS 0.375651f
C2061 a_2075_42718# VSS 0.349289f
C2062 a_468_42870# VSS 0.274851f
C2063 a_1387_42883# VSS 0.260413f
C2064 a_428_42724# VSS 0.411807f
C2065 a_283_42692# VSS 0.480504f
C2066 a_104_42692# VSS 0.324311f
C2067 a_n501_42718# VSS 0.276955f
C2068 COMP_N VSS 4.32737f
C2069 a_n1237_42718# VSS 0.254079f
C2070 COMP_P VSS 6.21892f
C2071 a_n1552_42692# VSS 0.309339f
C2072 a_n1920_42692# VSS 0.34902f
C2073 EN_COMP VSS 6.90846f
C2074 SMPL VSS 11.695511f
C2075 a_n2288_42692# VSS 0.351055f
C2076 a_n2833_42692# VSS 0.607654f
C2077 a_20283_43262# VSS 0.368993f
C2078 a_20049_43262# VSS 0.577664f
C2079 a_19633_43262# VSS 0.492249f
C2080 a_18541_43582# VSS 0.262572f
C2081 a_15133_43582# VSS 0.403353f
C2082 a_8969_43582# VSS 0.586904f
C2083 a_7735_42692# VSS 0.573616f
C2084 a_5473_43582# VSS 0.396943f
C2085 a_2075_42870# VSS 0.345465f
C2086 a_22959_43270# VSS 0.340508f
C2087 a_22223_43270# VSS 0.301232f
C2088 a_21908_43236# VSS 0.301841f
C2089 a_21719_43244# VSS 0.422943f
C2090 a_21540_43236# VSS 0.340463f
C2091 a_21197_42718# VSS 0.334383f
C2092 a_19771_43600# VSS 0.221721f
C2093 a_19191_43262# VSS 0.366256f
C2094 a_19003_43262# VSS 0.217513f
C2095 a_18766_43236# VSS 1.80153f
C2096 a_16404_43640# VSS 0.265567f
C2097 a_16579_43566# VSS 0.80329f
C2098 a_15839_43640# VSS 0.263388f
C2099 a_16057_43236# VSS 0.18191f
C2100 a_15489_43268# VSS 0.296553f
C2101 a_15323_43268# VSS 0.568054f
C2102 a_14647_43494# VSS 0.261364f
C2103 a_13460_43640# VSS 0.265959f
C2104 a_13635_43566# VSS 0.791232f
C2105 a_12895_43640# VSS 0.264457f
C2106 a_13113_43236# VSS 0.180143f
C2107 a_12545_43268# VSS 0.311807f
C2108 a_12379_43268# VSS 0.548002f
C2109 a_11252_43640# VSS 0.260731f
C2110 a_11427_43566# VSS 0.784536f
C2111 a_10687_43640# VSS 0.267689f
C2112 a_10905_43236# VSS 0.184446f
C2113 a_10337_43268# VSS 0.305311f
C2114 a_10475_43433# VSS 0.297015f
C2115 a_10171_43268# VSS 0.645859f
C2116 a_9637_43560# VSS 0.298551f
C2117 a_9208_43494# VSS 0.250621f
C2118 a_7347_43494# VSS 0.371409f
C2119 a_6519_43494# VSS 0.369749f
C2120 a_4352_43640# VSS 0.26331f
C2121 a_4527_43566# VSS 0.79431f
C2122 a_3787_43640# VSS 0.255739f
C2123 a_4005_43236# VSS 0.178849f
C2124 a_3437_43268# VSS 0.2947f
C2125 a_3165_43262# VSS 0.41398f
C2126 a_3271_43268# VSS 0.523979f
C2127 a_2627_43262# VSS 0.371717f
C2128 a_1339_43315# VSS 0.240943f
C2129 a_n1429_43262# VSS 0.349868f
C2130 a_n1741_42692# VSS 0.34585f
C2131 a_1488_43236# VSS 0.432387f
C2132 a_396_43640# VSS 0.269395f
C2133 a_571_43566# VSS 0.503099f
C2134 a_n169_43640# VSS 0.257052f
C2135 a_49_43236# VSS 0.183041f
C2136 a_n519_43268# VSS 0.301512f
C2137 a_n685_43268# VSS 0.567194f
C2138 a_n2104_43236# VSS 0.332519f
C2139 a_n2472_43236# VSS 0.333624f
C2140 a_n2840_43236# VSS 0.3411f
C2141 a_22959_43806# VSS 0.345335f
C2142 a_22591_43806# VSS 0.324913f
C2143 a_22223_43494# VSS 0.523101f
C2144 a_22087_43244# VSS 0.467296f
C2145 a_21847_43806# VSS 0.498815f
C2146 a_20107_43806# VSS 0.654308f
C2147 a_18704_43806# VSS 0.256559f
C2148 a_18879_43780# VSS 0.768734f
C2149 a_18139_43806# VSS 0.254459f
C2150 a_18357_44048# VSS 0.179724f
C2151 a_17789_43806# VSS 0.292062f
C2152 a_17623_43806# VSS 0.582502f
C2153 a_17515_43806# VSS 0.262832f
C2154 a_17242_43806# VSS 0.268821f
C2155 a_16036_43806# VSS 0.260052f
C2156 a_16211_43780# VSS 0.493477f
C2157 a_15471_43806# VSS 0.254196f
C2158 a_15689_44048# VSS 0.175874f
C2159 a_15121_43806# VSS 0.298131f
C2160 a_14955_43806# VSS 0.5491f
C2161 a_14757_43806# VSS 0.606408f
C2162 a_14301_44035# VSS 0.669876f
C2163 a_14077_44133# VSS 0.283524f
C2164 a_14331_44133# VSS 0.268784f
C2165 a_10612_43806# VSS 0.18415f
C2166 a_10362_43806# VSS 0.260002f
C2167 a_13536_43780# VSS 0.307058f
C2168 a_12448_43806# VSS 0.257604f
C2169 a_12623_43780# VSS 0.758145f
C2170 a_11883_43806# VSS 0.265551f
C2171 a_12101_44048# VSS 0.174512f
C2172 a_11533_43806# VSS 0.297036f
C2173 a_11367_43806# VSS 0.51972f
C2174 a_9416_43530# VSS 0.636336f
C2175 a_10414_43780# VSS 0.306684f
C2176 a_9863_43958# VSS 0.242658f
C2177 a_9343_43806# VSS 0.31883f
C2178 a_8308_43806# VSS 0.265008f
C2179 a_8483_43780# VSS 0.759819f
C2180 a_7743_43806# VSS 0.280127f
C2181 a_7961_44048# VSS 0.195871f
C2182 a_7393_43806# VSS 0.306016f
C2183 a_7319_43262# VSS 0.401189f
C2184 a_7227_43806# VSS 0.554242f
C2185 a_5916_43806# VSS 0.264628f
C2186 a_6091_43780# VSS 0.777418f
C2187 a_5351_43806# VSS 0.250116f
C2188 a_5569_44048# VSS 0.17997f
C2189 a_5001_43806# VSS 0.289424f
C2190 a_4835_43806# VSS 0.523822f
C2191 a_3524_43806# VSS 0.259361f
C2192 a_3699_43780# VSS 0.759715f
C2193 a_2959_43806# VSS 0.255603f
C2194 a_3177_44048# VSS 0.179433f
C2195 a_2609_43806# VSS 0.297852f
C2196 a_2627_42718# VSS 0.364833f
C2197 a_2443_43806# VSS 0.526629f
C2198 a_2043_43958# VSS 0.23333f
C2199 a_948_43806# VSS 0.261292f
C2200 a_1123_43780# VSS 0.768791f
C2201 a_383_43806# VSS 0.26443f
C2202 a_601_44048# VSS 0.189664f
C2203 a_33_43806# VSS 0.300862f
C2204 a_n133_43806# VSS 0.559871f
C2205 a_n2073_43806# VSS 0.504203f
C2206 a_n2472_43780# VSS 0.323815f
C2207 a_n2840_43780# VSS 0.327636f
C2208 a_22591_43958# VSS 0.332056f
C2209 a_22031_44350# VSS 0.64304f
C2210 a_16868_44670# VSS 0.179613f
C2211 a_16618_44670# VSS 0.255869f
C2212 a_15415_44350# VSS 0.591199f
C2213 a_22959_44358# VSS 0.341461f
C2214 a_22223_44358# VSS 0.330214f
C2215 a_21755_44350# VSS 0.362345f
C2216 a_18796_44728# VSS 0.268f
C2217 a_18971_44654# VSS 0.769803f
C2218 a_18231_44728# VSS 0.262514f
C2219 a_18449_44324# VSS 0.184533f
C2220 a_17881_44356# VSS 0.294994f
C2221 a_17715_44356# VSS 0.589315f
C2222 a_16670_44324# VSS 0.341243f
C2223 a_16211_44582# VSS 0.236534f
C2224 a_15443_44582# VSS 0.356077f
C2225 a_15091_44440# VSS 0.20859f
C2226 a_14133_43780# VSS 0.458275f
C2227 a_12683_43433# VSS 0.29982f
C2228 a_11671_44019# VSS 0.357116f
C2229 a_14819_44582# VSS 0.328746f
C2230 a_14545_44569# VSS 0.216724f
C2231 a_13725_44350# VSS 0.320205f
C2232 a_13561_44350# VSS 0.198639f
C2233 a_13023_44716# VSS 0.239821f
C2234 a_12379_44350# VSS 0.355519f
C2235 a_11183_44350# VSS 0.372184f
C2236 a_10844_44364# VSS 1.32199f
C2237 a_10447_44403# VSS 0.216951f
C2238 a_10596_44324# VSS 0.407912f
C2239 a_9159_43262# VSS 0.643188f
C2240 a_9266_44350# VSS 0.181586f
C2241 a_9335_44324# VSS 0.253997f
C2242 a_9140_44466# VSS 0.296807f
C2243 a_9179_44592# VSS 0.505851f
C2244 a_8862_44482# VSS 0.260283f
C2245 a_8659_44324# VSS 0.479122f
C2246 a_7415_44466# VSS 0.340276f
C2247 a_7309_44466# VSS 0.211621f
C2248 a_6491_44716# VSS 0.273533f
C2249 a_5387_44403# VSS 0.232413f
C2250 a_5139_44019# VSS 0.259754f
C2251 a_4080_44670# VSS 0.165523f
C2252 a_3830_44670# VSS 0.247727f
C2253 a_5536_44324# VSS 0.463872f
C2254 a_4651_44350# VSS 0.357207f
C2255 a_3882_44324# VSS 0.320037f
C2256 a_3576_44364# VSS 0.466897f
C2257 a_3179_44403# VSS 0.25695f
C2258 a_2332_44670# VSS 0.172554f
C2259 a_2082_44670# VSS 0.26684f
C2260 a_3328_44324# VSS 0.375262f
C2261 a_1736_43276# VSS 0.515198f
C2262 a_2134_44324# VSS 0.379805f
C2263 a_1659_44440# VSS 0.208782f
C2264 a_768_44670# VSS 0.181655f
C2265 a_518_44670# VSS 0.276019f
C2266 a_n381_43433# VSS 0.414791f
C2267 a_n2661_43780# VSS 0.452594f
C2268 a_n2293_43244# VSS 0.467621f
C2269 a_n2661_43244# VSS 0.559552f
C2270 a_1387_44582# VSS 0.332858f
C2271 a_546_43100# VSS 0.486528f
C2272 a_570_44324# VSS 0.308737f
C2273 a_161_44648# VSS 0.265599f
C2274 a_n60_44618# VSS 0.349173f
C2275 a_n172_44582# VSS 0.35074f
C2276 a_n268_44582# VSS 0.279143f
C2277 a_n2472_44324# VSS 0.331111f
C2278 a_n2840_44324# VSS 0.344855f
C2279 a_22959_44894# VSS 0.34535f
C2280 a_22591_44894# VSS 0.332786f
C2281 a_22399_44894# VSS 0.732543f
C2282 a_22123_44894# VSS 0.480559f
C2283 a_17613_44894# VSS 0.158531f
C2284 a_17531_44894# VSS 0.608913f
C2285 a_16824_45276# VSS 0.6536f
C2286 a_16427_44894# VSS 0.237297f
C2287 a_18495_44868# VSS 0.237293f
C2288 a_18319_44868# VSS 0.205156f
C2289 a_17951_44868# VSS 0.29118f
C2290 a_14204_44350# VSS 0.313448f
C2291 a_16576_44868# VSS 0.498937f
C2292 a_16074_45046# VSS 0.201908f
C2293 a_15323_44894# VSS 0.316044f
C2294 a_14635_44324# VSS 0.669251f
C2295 a_13469_44894# VSS 0.685781f
C2296 a_12287_44894# VSS 0.230752f
C2297 a_10215_44874# VSS 0.220224f
C2298 a_9304_43494# VSS 0.508582f
C2299 a_8699_44894# VSS 0.278238f
C2300 a_4703_44894# VSS 0.548619f
C2301 a_12931_44894# VSS 0.253016f
C2302 a_12436_44868# VSS 0.377707f
C2303 a_9943_45046# VSS 0.346523f
C2304 a_8848_44868# VSS 0.485694f
C2305 a_7842_44868# VSS 0.457431f
C2306 a_7020_44894# VSS 0.260397f
C2307 a_7195_44868# VSS 0.477363f
C2308 a_6455_44894# VSS 0.25686f
C2309 a_6673_45136# VSS 0.179477f
C2310 a_6105_44894# VSS 0.291282f
C2311 a_6243_45107# VSS 0.68028f
C2312 a_5939_44894# VSS 0.53906f
C2313 a_1935_44874# VSS 0.222352f
C2314 a_171_44019# VSS 0.969035f
C2315 a_636_42870# VSS 1.40743f
C2316 a_829_45221# VSS 0.328058f
C2317 a_n2293_43780# VSS 0.639185f
C2318 a_2471_45046# VSS 0.402687f
C2319 a_1663_45046# VSS 0.326509f
C2320 a_1083_45221# VSS 0.250946f
C2321 a_n2293_44868# VSS 0.347509f
C2322 a_n2472_44868# VSS 0.327725f
C2323 a_n2840_44868# VSS 0.327636f
C2324 a_22031_45438# VSS 0.930131f
C2325 a_19168_45758# VSS 0.177937f
C2326 a_18918_45758# VSS 0.274194f
C2327 a_17763_44868# VSS 0.293429f
C2328 a_22959_45446# VSS 0.3401f
C2329 a_22455_45420# VSS 0.459866f
C2330 a_22276_45412# VSS 0.347816f
C2331 a_18970_45412# VSS 0.386247f
C2332 a_18282_45670# VSS 0.229276f
C2333 a_16287_45744# VSS 0.229345f
C2334 a_16111_45412# VSS 0.20415f
C2335 a_13715_43780# VSS 0.754805f
C2336 a_15468_45412# VSS 0.394591f
C2337 a_14953_45554# VSS 0.227427f
C2338 a_14853_45438# VSS 0.198465f
C2339 a_13464_45758# VSS 0.166022f
C2340 a_13214_45758# VSS 0.245637f
C2341 a_12636_45758# VSS 0.165382f
C2342 a_12386_45758# VSS 0.267556f
C2343 a_13266_45412# VSS 0.368563f
C2344 a_12684_45276# VSS 0.517472f
C2345 a_12438_45412# VSS 0.287693f
C2346 a_11687_45528# VSS 0.220936f
C2347 a_9048_45758# VSS 0.165362f
C2348 a_8798_45758# VSS 0.249659f
C2349 a_11415_45670# VSS 0.33983f
C2350 a_11017_45736# VSS 0.286225f
C2351 a_10389_45438# VSS 0.304638f
C2352 a_10588_45670# VSS 0.271373f
C2353 a_10111_45776# VSS 0.244251f
C2354 a_8850_45412# VSS 0.379236f
C2355 a_8192_44874# VSS 0.728202f
C2356 a_8055_45491# VSS 0.220165f
C2357 a_2301_45758# VSS 0.208812f
C2358 a_8204_45412# VSS 0.392056f
C2359 a_7705_45736# VSS 0.2777f
C2360 a_6985_45438# VSS 0.354444f
C2361 a_7372_45670# VSS 0.483497f
C2362 a_7276_45670# VSS 0.263703f
C2363 a_6707_45776# VSS 0.221264f
C2364 a_6325_45736# VSS 0.280745f
C2365 a_5896_45670# VSS 0.261734f
C2366 a_4812_45816# VSS 0.260026f
C2367 a_4987_45742# VSS 0.47633f
C2368 a_4247_45816# VSS 0.260931f
C2369 a_4465_45412# VSS 0.179989f
C2370 a_3897_45444# VSS 0.300352f
C2371 a_3731_45444# VSS 0.571277f
C2372 a_2151_45670# VSS 0.304299f
C2373 a_1659_45528# VSS 0.213768f
C2374 a_n2293_44332# VSS 0.920405f
C2375 a_n2661_44332# VSS 0.471405f
C2376 a_n2661_44868# VSS 0.354678f
C2377 a_1387_45670# VSS 0.336507f
C2378 a_989_45736# VSS 0.276345f
C2379 a_361_45438# VSS 0.318362f
C2380 a_656_45670# VSS 0.307407f
C2381 a_560_45670# VSS 0.274896f
C2382 a_83_45776# VSS 0.230216f
C2383 a_n377_45776# VSS 0.261823f
C2384 a_n2472_45412# VSS 0.326765f
C2385 a_n2840_45412# VSS 0.340687f
C2386 a_22959_45982# VSS 0.34535f
C2387 a_22591_45982# VSS 0.364526f
C2388 a_16177_45982# VSS 0.200794f
C2389 a_13738_46032# VSS 0.110759f
C2390 a_13572_46032# VSS 0.239084f
C2391 a_12931_45982# VSS 0.25841f
C2392 a_18704_45982# VSS 0.265234f
C2393 a_18879_45956# VSS 0.515938f
C2394 a_18139_45982# VSS 0.258912f
C2395 a_18357_46224# VSS 0.178783f
C2396 a_17789_45982# VSS 0.291971f
C2397 a_17623_45982# VSS 0.543076f
C2398 a_15187_44868# VSS 1.6572f
C2399 a_16750_46134# VSS 0.329655f
C2400 a_16085_45982# VSS 0.248665f
C2401 a_14955_45982# VSS 0.532416f
C2402 a_15328_46134# VSS 0.580212f
C2403 a_14382_46348# VSS 0.315272f
C2404 a_14194_46348# VSS 0.2215f
C2405 a_13151_45956# VSS 0.388876f
C2406 a_12121_45956# VSS 0.341096f
C2407 a_11788_46134# VSS 1.52216f
C2408 a_11692_46134# VSS 0.260658f
C2409 a_10884_45982# VSS 0.258645f
C2410 a_11059_45956# VSS 0.475832f
C2411 a_10319_45982# VSS 0.258264f
C2412 a_10537_46224# VSS 0.178741f
C2413 a_9969_45982# VSS 0.293075f
C2414 a_9803_45982# VSS 0.546136f
C2415 a_8651_45962# VSS 0.218146f
C2416 a_7981_45956# VSS 0.275743f
C2417 a_7648_46134# VSS 0.287601f
C2418 a_9343_45982# VSS 0.346088f
C2419 a_8379_46134# VSS 0.32098f
C2420 a_7552_46134# VSS 0.24601f
C2421 a_5129_45956# VSS 0.285091f
C2422 a_2535_45670# VSS 0.672209f
C2423 a_7016_46231# VSS 0.478472f
C2424 a_6322_46348# VSS 0.180083f
C2425 a_6391_46219# VSS 0.256321f
C2426 a_6235_46124# VSS 0.503906f
C2427 a_6196_46250# VSS 0.290175f
C2428 a_5655_43780# VSS 3.16689f
C2429 a_5918_46234# VSS 0.259525f
C2430 a_5715_45956# VSS 0.479674f
C2431 a_4700_46134# VSS 0.26664f
C2432 a_4061_45956# VSS 0.285185f
C2433 a_3165_45982# VSS 1.05287f
C2434 a_3470_45982# VSS 0.292857f
C2435 a_3320_46134# VSS 0.208094f
C2436 a_2512_45982# VSS 0.253039f
C2437 a_2687_45956# VSS 0.486421f
C2438 a_1947_45982# VSS 0.264771f
C2439 a_2165_46224# VSS 0.185513f
C2440 a_1597_45982# VSS 0.302033f
C2441 a_1735_46195# VSS 0.705483f
C2442 a_1431_45982# VSS 0.551523f
C2443 a_672_45982# VSS 0.283236f
C2444 a_847_45956# VSS 0.480253f
C2445 a_107_45982# VSS 0.267162f
C2446 a_325_46224# VSS 0.191551f
C2447 a_n243_45982# VSS 0.319397f
C2448 a_n105_46195# VSS 0.812722f
C2449 a_n409_45982# VSS 0.691293f
C2450 a_n2472_45956# VSS 0.34647f
C2451 a_n2840_45956# VSS 0.344757f
C2452 a_22959_46534# VSS 0.345334f
C2453 a_22223_46534# VSS 0.379678f
C2454 a_19566_45670# VSS 1.14128f
C2455 a_19371_46579# VSS 0.244045f
C2456 a_16921_46364# VSS 0.256092f
C2457 a_16128_46134# VSS 0.18552f
C2458 a_15079_46134# VSS 0.271292f
C2459 a_15033_46526# VSS 0.223394f
C2460 a_19520_46500# VSS 0.459581f
C2461 a_18190_46526# VSS 0.179726f
C2462 a_18259_46500# VSS 0.259381f
C2463 a_18064_46642# VSS 0.291431f
C2464 a_18103_46768# VSS 0.515254f
C2465 a_17786_46658# VSS 0.265919f
C2466 a_17583_46500# VSS 0.503241f
C2467 a_16651_46500# VSS 0.228426f
C2468 a_16555_46616# VSS 0.17847f
C2469 a_16291_44914# VSS 1.49632f
C2470 a_16291_46758# VSS 0.320944f
C2471 a_15309_45438# VSS 0.453309f
C2472 a_14757_45982# VSS 0.228174f
C2473 a_15192_46500# VSS 0.343602f
C2474 a_14658_46526# VSS 0.309789f
C2475 a_14470_46526# VSS 0.234916f
C2476 a_14014_46842# VSS 0.110542f
C2477 a_13848_46842# VSS 0.239079f
C2478 a_13207_46892# VSS 0.255986f
C2479 a_13427_46756# VSS 0.38761f
C2480 a_12699_46616# VSS 0.215405f
C2481 a_10684_45670# VSS 0.451513f
C2482 a_9973_46526# VSS 0.255725f
C2483 a_12427_46758# VSS 0.324097f
C2484 a_12127_46744# VSS 3.27347f
C2485 a_11971_46500# VSS 0.338384f
C2486 a_11160_46904# VSS 0.260214f
C2487 a_11335_46830# VSS 0.481209f
C2488 a_10595_46904# VSS 0.258541f
C2489 a_10813_46500# VSS 0.174521f
C2490 a_10245_46532# VSS 0.291905f
C2491 a_10383_46697# VSS 0.47335f
C2492 a_10079_46532# VSS 0.502368f
C2493 a_9547_46565# VSS 0.242569f
C2494 a_9293_46565# VSS 0.296391f
C2495 a_9349_46539# VSS 0.388872f
C2496 a_8308_46904# VSS 0.264268f
C2497 a_8483_46830# VSS 0.491437f
C2498 a_7743_46904# VSS 0.261039f
C2499 a_7961_46500# VSS 0.18117f
C2500 a_7393_46532# VSS 0.299652f
C2501 a_7503_45982# VSS 0.26104f
C2502 a_7227_46532# VSS 0.546522f
C2503 a_6631_44582# VSS 1.64026f
C2504 a_6126_46642# VSS 0.402949f
C2505 a_5784_44364# VSS 0.591f
C2506 a_5626_46846# VSS 0.208297f
C2507 a_5382_44582# VSS 0.838724f
C2508 a_4322_46134# VSS 4.55741f
C2509 a_5441_46500# VSS 0.237953f
C2510 a_4352_46904# VSS 0.263214f
C2511 a_4527_46830# VSS 0.765866f
C2512 a_3787_46904# VSS 0.260402f
C2513 a_4005_46500# VSS 0.183581f
C2514 a_3437_46532# VSS 0.285237f
C2515 a_3575_46697# VSS 0.299332f
C2516 a_3271_46532# VSS 0.534342f
C2517 a_2645_46824# VSS 0.333326f
C2518 a_82_45670# VSS 0.994669f
C2519 a_2216_46758# VSS 0.269229f
C2520 a_1633_46824# VSS 0.308239f
C2521 a_1204_46758# VSS 0.263734f
C2522 a_396_46904# VSS 0.279108f
C2523 a_571_46830# VSS 0.499186f
C2524 a_n169_46904# VSS 0.259048f
C2525 a_49_46500# VSS 0.183309f
C2526 a_n519_46532# VSS 0.307889f
C2527 a_n685_46532# VSS 0.609657f
C2528 a_n2472_46500# VSS 0.342754f
C2529 a_n2840_46500# VSS 0.340313f
C2530 a_22959_47070# VSS 0.345439f
C2531 a_22591_47070# VSS 0.33284f
C2532 a_22223_47070# VSS 0.33659f
C2533 a_18803_47070# VSS 0.379517f
C2534 a_15155_47070# VSS 0.315028f
C2535 a_14950_43958# VSS 3.22761f
C2536 a_14573_47070# VSS 0.359955f
C2537 a_4908_45956# VSS 3.33493f
C2538 a_12747_47070# VSS 0.262856f
C2539 a_18689_45412# VSS 0.89418f
C2540 a_10251_45454# VSS 5.03531f
C2541 a_18530_47070# VSS 0.286339f
C2542 a_17927_46195# VSS 0.779881f
C2543 a_18133_47235# VSS 0.25425f
C2544 a_16703_45982# VSS 0.408993f
C2545 a_16561_45982# VSS 0.406143f
C2546 a_15879_47320# VSS 0.36634f
C2547 a_15582_45982# VSS 0.283825f
C2548 a_15691_47436# VSS 0.209316f
C2549 a_15329_47044# VSS 0.901189f
C2550 a_15221_47044# VSS 0.342975f
C2551 a_15113_47222# VSS 0.27905f
C2552 a_15005_47222# VSS 0.141613f
C2553 a_14219_47070# VSS 0.259428f
C2554 a_12896_47044# VSS 0.491832f
C2555 a_11795_47044# VSS 0.658686f
C2556 a_7429_47044# VSS 0.280959f
C2557 a_7208_47044# VSS 7.02295f
C2558 a_5663_45982# VSS 1.32924f
C2559 a_7760_45956# VSS 0.45426f
C2560 a_4035_45609# VSS 0.774799f
C2561 a_713_47044# VSS 0.291731f
C2562 a_380_47222# VSS 0.450989f
C2563 a_n381_46697# VSS 0.822009f
C2564 a_85_47070# VSS 0.472461f
C2565 a_n194_47222# VSS 0.532579f
C2566 a_11248_47319# VSS 0.316376f
C2567 a_10554_47436# VSS 0.187856f
C2568 a_10623_47307# VSS 0.257645f
C2569 a_10467_47212# VSS 0.520916f
C2570 a_10428_47338# VSS 0.293186f
C2571 a_10150_47322# VSS 0.261818f
C2572 a_9947_47044# VSS 0.48295f
C2573 a_9395_47044# VSS 0.376159f
C2574 a_8391_47044# VSS 0.674785f
C2575 a_7839_47222# VSS 0.239015f
C2576 a_7000_47222# VSS 0.264125f
C2577 a_6635_47044# VSS 0.326716f
C2578 a_5749_47222# VSS 0.626402f
C2579 a_5419_47258# VSS 2.20741f
C2580 a_5089_47044# VSS 0.533395f
C2581 a_4993_47044# VSS 0.919136f
C2582 a_4704_47044# VSS 0.350951f
C2583 a_4061_47044# VSS 0.571551f
C2584 a_2167_46526# VSS 0.571922f
C2585 a_1431_47070# VSS 0.72581f
C2586 a_1115_47044# VSS 0.298278f
C2587 a_284_47222# VSS 0.288394f
C2588 a_n193_47098# VSS 0.270684f
C2589 a_n447_47044# VSS 1.02649f
C2590 a_n2104_47044# VSS 0.343495f
C2591 a_n2472_47044# VSS 0.323981f
C2592 a_n2840_47044# VSS 0.328049f
C2593 a_16475_45412# VSS 2.6694f
C2594 a_16102_47044# VSS 0.206374f
C2595 a_15437_47044# VSS 0.377093f
C2596 a_22959_47622# VSS 0.314903f
C2597 a_22733_47833# VSS 0.22632f
C2598 a_22223_47622# VSS 0.32008f
C2599 SMPL_ON_N VSS 8.374041f
C2600 a_21997_47833# VSS 0.235531f
C2601 a_21629_47833# VSS 0.23347f
C2602 a_20159_47588# VSS 0.408589f
C2603 a_18135_47588# VSS 0.376962f
C2604 a_16335_47614# VSS 0.232001f
C2605 a_15871_47614# VSS 0.212431f
C2606 a_15691_47614# VSS 0.228455f
C2607 a_15139_47730# VSS 0.33154f
C2608 a_14757_47614# VSS 2.84195f
C2609 a_9551_47203# VSS 0.319997f
C2610 a_9517_46539# VSS 0.903198f
C2611 a_14587_47614# VSS 0.265543f
C2612 a_12887_47833# VSS 0.275787f
C2613 a_11507_47833# VSS 0.261094f
C2614 a_11299_47832# VSS 0.328275f
C2615 a_11143_47588# VSS 0.31161f
C2616 a_10415_47846# VSS 0.25088f
C2617 a_9863_47874# VSS 0.552881f
C2618 a_7595_47614# VSS 0.587796f
C2619 a_7311_47614# VSS 0.341037f
C2620 a_6951_47070# VSS 0.407912f
C2621 a_5847_47614# VSS 0.630493f
C2622 a_5839_47070# VSS 0.366337f
C2623 a_4651_47614# VSS 0.613894f
C2624 a_4091_47070# VSS 0.377596f
C2625 a_2351_47614# VSS 0.649511f
C2626 a_2343_47070# VSS 0.389243f
C2627 a_1209_47588# VSS 0.568213f
C2628 a_999_47846# VSS 0.423662f
C2629 a_663_47874# VSS 0.659011f
C2630 a_n749_47846# VSS 0.506925f
C2631 a_n1085_47874# VSS 0.684414f
C2632 a_n1605_47614# VSS 0.239738f
C2633 SMPL_ON_P VSS 7.6046f
C2634 a_n1920_47588# VSS 0.310464f
C2635 a_n2288_47588# VSS 0.34713f
C2636 a_n2833_47874# VSS 0.602779f
C2637 a_n2442_43806.n0 VSS 0.197962f
C2638 a_n2442_43806.t4 VSS 2.36492f
C2639 a_n2442_43806.n1 VSS 19.0336f
C2640 C0_P_btm.t0 VSS 1.37053f
C2641 C0_P_btm.t5 VSS 0.408265f
C2642 C0_P_btm.t2 VSS 0.275201f
C2643 C0_P_btm.n0 VSS 2.21668f
C2644 C0_P_btm.n1 VSS 3.36018f
C2645 C0_P_btm.t1 VSS 0.19597f
C2646 C0_P_btm.n2 VSS 3.88706f
C2647 C0_P_btm.t4 VSS 1.2515f
C2648 C0_P_btm.t3 VSS 1.18437f
C2649 C0_P_btm.n3 VSS 1.08249f
C2650 a_14087_32299.n0 VSS 0.126869f
C2651 a_14087_32299.t4 VSS 2.59395f
C2652 a_14087_32299.n1 VSS 18.8173f
C2653 a_14087_32299.n2 VSS 0.152641f
C2654 a_19437_31459.n0 VSS 0.121988f
C2655 a_19437_31459.t4 VSS 3.06749f
C2656 a_19437_31459.n1 VSS 15.062501f
C2657 a_19437_31459.n2 VSS 0.146769f
C2658 a_n2074_47070.n0 VSS 0.179596f
C2659 a_n2074_47070.t4 VSS 2.90799f
C2660 a_n2074_47070.n1 VSS 15.137099f
C2661 a_n2109_42692.n1 VSS 2.15062f
C2662 a_n2109_42692.n2 VSS 10.7108f
C2663 a_n2109_42692.n3 VSS 0.302295f
C2664 a_n2109_42692.t0 VSS 0.215183f
C2665 a_n2074_43262.n0 VSS 0.122763f
C2666 a_n2074_43262.t4 VSS 2.5595f
C2667 a_n2074_43262.n1 VSS 18.6676f
C2668 a_n2074_43262.n2 VSS 0.1477f
C2669 a_10199_47846.t1 VSS 0.125574f
C2670 a_10199_47846.n0 VSS 0.279876f
C2671 a_10199_47846.n1 VSS 1.91682f
C2672 a_10199_47846.t0 VSS 0.103245f
C2673 a_n2810_45438.t4 VSS 2.91575f
C2674 a_n2810_45438.n0 VSS 0.184889f
C2675 a_n2810_45438.n1 VSS 15.115901f
C2676 a_11730_34132.n0 VSS 1.72361f
C2677 a_11730_34132.n1 VSS 1.7928f
C2678 a_11730_34132.t6 VSS 4.75589f
C2679 a_11730_34132.n2 VSS 0.393499f
C2680 a_11730_34132.n3 VSS 1.67051f
C2681 a_11730_34132.n4 VSS 0.532613f
C2682 a_11730_34132.t7 VSS 4.75589f
C2683 a_11730_34132.n5 VSS 3.7477f
C2684 a_11730_34132.t4 VSS 4.75589f
C2685 a_11730_34132.n6 VSS 1.72657f
C2686 a_11730_34132.n7 VSS 0.438123f
C2687 a_11730_34132.n8 VSS 0.171855f
C2688 a_11730_34132.n9 VSS 0.172177f
C2689 a_11730_34132.n10 VSS 0.441755f
C2690 a_11730_34132.n11 VSS 0.397556f
C2691 a_11730_34132.t5 VSS 4.75589f
C2692 a_11730_34132.n12 VSS 3.76147f
C2693 a_11730_34132.n13 VSS 0.435659f
C2694 a_11730_34132.n14 VSS 0.442094f
C2695 a_11730_34132.n16 VSS 0.512191f
C2696 a_4758_30651.n0 VSS 0.124511f
C2697 a_4758_30651.t8 VSS 0.546341f
C2698 a_4758_30651.t9 VSS 0.562631f
C2699 a_4758_30651.n1 VSS 0.496254f
C2700 a_4758_30651.t10 VSS 0.546341f
C2701 a_4758_30651.t7 VSS 0.547263f
C2702 a_4758_30651.n2 VSS 0.251135f
C2703 a_4758_30651.n3 VSS 0.270041f
C2704 a_4758_30651.n4 VSS 1.71278f
C2705 a_4758_30651.t6 VSS 0.546341f
C2706 a_4758_30651.n5 VSS 0.270041f
C2707 a_4758_30651.t13 VSS 0.546341f
C2708 a_4758_30651.t4 VSS 0.547263f
C2709 a_4758_30651.n6 VSS 0.251135f
C2710 a_4758_30651.t11 VSS 0.562631f
C2711 a_4758_30651.n7 VSS 0.496254f
C2712 a_4758_30651.n8 VSS 1.85692f
C2713 a_4758_30651.n9 VSS 7.53757f
C2714 a_4758_30651.n10 VSS 0.155346f
C2715 a_4758_30651.n11 VSS 4.2424f
C2716 a_4758_30651.n12 VSS 0.334792f
C2717 CAL_N.n0 VSS 2.22732f
C2718 CAL_N.t4 VSS 6.16073f
C2719 CAL_N.n1 VSS 4.30995f
C2720 CAL_N.t6 VSS 5.48889f
C2721 CAL_N.n2 VSS 4.30902f
C2722 CAL_N.t5 VSS 6.14892f
C2723 CAL_N.n3 VSS 2.15694f
C2724 CAL_N.n4 VSS 0.211393f
C2725 CAL_N.n6 VSS 0.412662f
C2726 CAL_N.n7 VSS 0.435954f
C2727 CAL_N.t3 VSS 0.121809f
C2728 a_6104_45706.n6 VSS 0.409845f
C2729 a_6104_45706.n7 VSS 0.807806f
C2730 a_6104_45706.n9 VSS 4.707911f
C2731 a_6104_45706.n10 VSS 0.293066f
C2732 a_6104_45706.n11 VSS 0.152853f
C2733 w_11534_34010.n3 VSS 0.568392f
C2734 w_11534_34010.n4 VSS 0.540037f
C2735 w_11534_34010.n5 VSS 1.1728f
C2736 w_11534_34010.n6 VSS 0.148417f
C2737 w_11534_34010.n7 VSS 0.1697f
C2738 w_11534_34010.n8 VSS 0.211327f
C2739 w_11534_34010.n9 VSS 0.240728f
C2740 w_11534_34010.n10 VSS 0.45959f
C2741 w_11534_34010.n17 VSS 0.109775f
C2742 w_11534_34010.n19 VSS 0.302685f
C2743 w_11534_34010.t0 VSS 0.296285f
C2744 w_11534_34010.t4 VSS 0.150361f
C2745 w_11534_34010.n22 VSS 0.140807f
C2746 w_11534_34010.t6 VSS 0.20257f
C2747 w_11534_34010.t2 VSS 0.150361f
C2748 w_11534_34010.n29 VSS 0.100241f
C2749 w_11534_34010.t8 VSS 0.149521f
C2750 w_11534_34010.n40 VSS 0.174293f
C2751 w_11534_34010.n42 VSS 2.23079f
C2752 w_11534_34010.n44 VSS 1.17099f
C2753 w_11534_34010.n48 VSS 0.138908f
C2754 w_11534_34010.n50 VSS 0.134774f
C2755 w_11534_34010.n51 VSS 3.24248f
C2756 w_11534_34010.t13 VSS 5.81627f
C2757 w_11534_34010.n52 VSS 5.60723f
C2758 w_11534_34010.t10 VSS 5.84551f
C2759 w_11534_34010.n53 VSS 3.4195f
C2760 w_11534_34010.n54 VSS 0.136143f
C2761 w_11534_34010.n55 VSS 0.122267f
C2762 w_11534_34010.n57 VSS 0.495855f
C2763 w_11534_34010.n58 VSS 0.53986f
C2764 w_11534_34010.n59 VSS 1.17461f
C2765 w_11534_34010.n60 VSS 2.23079f
C2766 w_11534_34010.n62 VSS 1.1722f
C2767 w_11534_34010.n63 VSS 0.259475f
C2768 w_11534_34010.n65 VSS 0.113577f
C2769 w_11534_34010.n66 VSS 0.147261f
C2770 w_11534_34010.n68 VSS 0.262162f
C2771 a_n2442_45438.n0 VSS 0.120694f
C2772 a_n2442_45438.t4 VSS 3.09965f
C2773 a_n2442_45438.n1 VSS 14.7354f
C2774 a_n2442_45438.n2 VSS 0.145211f
C2775 a_19921_31459.n0 VSS 0.180578f
C2776 a_19921_31459.t4 VSS 2.80592f
C2777 a_19921_31459.n1 VSS 15.3367f
C2778 a_2252_42718.n0 VSS 0.145352f
C2779 a_2252_42718.n1 VSS 0.217481f
C2780 a_2252_42718.t7 VSS 0.319526f
C2781 a_2252_42718.t4 VSS 0.317625f
C2782 a_2252_42718.n2 VSS 15.062099f
C2783 a_2252_42718.n3 VSS 9.41684f
C2784 a_2252_42718.n4 VSS 0.475932f
C2785 a_4338_37500.n1 VSS 0.347491f
C2786 a_4338_37500.n2 VSS 0.476562f
C2787 a_4338_37500.n3 VSS 0.110266f
C2788 a_4338_37500.n4 VSS 1.30834f
C2789 a_n1435_47614.n0 VSS 0.277643f
C2790 a_n1435_47614.n1 VSS 1.62141f
C2791 a_n1435_47614.t0 VSS 0.105249f
C2792 a_n1890_47614.t5 VSS 1.57442f
C2793 a_n1890_47614.t4 VSS 1.57421f
C2794 a_n1890_47614.n1 VSS 8.4357f
C2795 a_n1890_47614.n2 VSS 6.25719f
C2796 a_n1890_47614.n3 VSS 0.111953f
C2797 a_n2442_46526.n0 VSS 0.12126f
C2798 a_n2442_46526.t4 VSS 3.1053f
C2799 a_n2442_46526.n1 VSS 14.827499f
C2800 a_n2442_46526.n2 VSS 0.145892f
C2801 a_n2810_45982.n0 VSS 0.126961f
C2802 a_n2810_45982.t4 VSS 2.92111f
C2803 a_n2810_45982.n1 VSS 15.0069f
C2804 a_n2810_45982.n2 VSS 0.14024f
C2805 a_n2103_44324.n1 VSS 0.459725f
C2806 a_n2103_44324.n3 VSS 0.320096f
C2807 a_n2103_44324.n4 VSS 7.029871f
C2808 C2_P_btm.t0 VSS 1.43551f
C2809 C2_P_btm.t3 VSS 0.436024f
C2810 C2_P_btm.t1 VSS 0.292486f
C2811 C2_P_btm.n0 VSS 2.30503f
C2812 C2_P_btm.n1 VSS 3.53635f
C2813 C2_P_btm.t2 VSS 0.199791f
C2814 C2_P_btm.n2 VSS 4.28972f
C2815 C2_P_btm.t5 VSS 1.29119f
C2816 C2_P_btm.t7 VSS 1.25457f
C2817 C2_P_btm.n3 VSS 0.416387f
C2818 C2_P_btm.t8 VSS 1.25665f
C2819 C2_P_btm.n4 VSS 0.394884f
C2820 C2_P_btm.t6 VSS 1.25876f
C2821 C2_P_btm.n5 VSS 0.44674f
C2822 C2_P_btm.t4 VSS 1.25876f
C2823 C2_P_btm.n6 VSS 0.815094f
C2824 a_14409_32299.n0 VSS 0.194736f
C2825 a_14409_32299.t4 VSS 2.25864f
C2826 a_14409_32299.n1 VSS 19.2481f
C2827 a_n2810_43262.t4 VSS 2.50052f
C2828 a_n2810_43262.n0 VSS 0.200941f
C2829 a_n2810_43262.n1 VSS 18.8905f
C2830 a_n2442_45982.n0 VSS 0.177304f
C2831 a_n2442_45982.t4 VSS 2.77325f
C2832 a_n2442_45982.n1 VSS 15.177599f
C2833 a_n2661_47044.n1 VSS 1.0299f
C2834 a_n2661_47044.n3 VSS 0.434649f
C2835 a_n2661_47044.n4 VSS 10.0283f
C2836 a_n2661_47044.n5 VSS 0.154833f
C2837 a_n2103_43780.n0 VSS 1.86657f
C2838 a_n2103_43780.n2 VSS 0.51593f
C2839 a_n2103_43780.n3 VSS 9.9264f
C2840 a_n2103_43780.n5 VSS 0.144493f
C2841 a_n2103_43780.n8 VSS 0.315298f
C2842 a_n2103_43780.n9 VSS 0.175706f
C2843 a_1651_47044.n0 VSS 0.445914f
C2844 a_1651_47044.n1 VSS 1.68331f
C2845 a_5542_30651.n0 VSS 0.106151f
C2846 a_5542_30651.n1 VSS 0.129987f
C2847 a_5542_30651.t5 VSS 0.112023f
C2848 a_5542_30651.t6 VSS 0.128813f
C2849 a_5542_30651.n2 VSS 0.512283f
C2850 a_5542_30651.t9 VSS 0.112023f
C2851 a_5542_30651.t4 VSS 0.128813f
C2852 a_5542_30651.n3 VSS 0.443957f
C2853 a_5542_30651.n4 VSS 11.8132f
C2854 a_5542_30651.n5 VSS 7.3358f
C2855 a_5542_30651.n6 VSS 0.324865f
C2856 a_13878_32299.n0 VSS 0.120711f
C2857 a_13878_32299.t4 VSS 2.57761f
C2858 a_13878_32299.n1 VSS 19.057402f
C2859 a_13878_32299.n2 VSS 0.145232f
C2860 a_1736_39587.t6 VSS 0.129045f
C2861 a_1736_39587.n0 VSS 0.790958f
C2862 a_1736_39587.n2 VSS 0.582262f
C2863 a_1736_39587.n3 VSS 0.316293f
C2864 a_1736_39587.n4 VSS 0.599955f
C2865 a_1736_39587.t0 VSS 0.313767f
C2866 a_1412_46794.n7 VSS 0.225487f
C2867 a_1412_46794.n8 VSS 0.45839f
C2868 a_1412_46794.n9 VSS 1.28872f
C2869 a_1412_46794.n10 VSS 0.205105f
C2870 a_13458_32299.t4 VSS 1.54944f
C2871 a_13458_32299.n1 VSS 11.3788f
C2872 VDAC_Pi.n2 VSS 0.665943f
C2873 VDAC_Pi.t8 VSS 0.180328f
C2874 VDAC_Pi.t10 VSS 0.150409f
C2875 VDAC_Pi.n3 VSS 2.14996f
C2876 VDAC_Pi.n4 VSS 0.329095f
C2877 VDAC_Pi.n5 VSS 0.109636f
C2878 VDAC_Pi.n6 VSS 0.242751f
C2879 VDAC_Pi.n7 VSS 0.109636f
C2880 VDAC_Pi.n8 VSS 0.442463f
C2881 COMP_N.n2 VSS 0.118121f
C2882 COMP_N.n5 VSS 0.159963f
C2883 COMP_N.n7 VSS 0.361261f
C2884 a_n2810_46526.t4 VSS 3.15421f
C2885 a_n2810_46526.n0 VSS 0.174614f
C2886 a_n2810_46526.n1 VSS 14.903501f
C2887 a_20405_31459.n0 VSS 0.123019f
C2888 a_20405_31459.t4 VSS 3.06767f
C2889 a_20405_31459.n1 VSS 15.058401f
C2890 a_20405_31459.n2 VSS 0.148008f
C2891 a_21788_30659.t5 VSS 0.833111f
C2892 a_21788_30659.t6 VSS 0.833239f
C2893 a_21788_30659.t10 VSS 0.83311f
C2894 a_21788_30659.n0 VSS 0.618066f
C2895 a_21788_30659.t8 VSS 0.83311f
C2896 a_21788_30659.n1 VSS 0.313199f
C2897 a_21788_30659.t9 VSS 0.83311f
C2898 a_21788_30659.n2 VSS 0.313199f
C2899 a_21788_30659.t4 VSS 0.83311f
C2900 a_21788_30659.n3 VSS 0.313199f
C2901 a_21788_30659.t11 VSS 0.83311f
C2902 a_21788_30659.n4 VSS 0.313199f
C2903 a_21788_30659.t7 VSS 0.83311f
C2904 a_21788_30659.n5 VSS 0.312158f
C2905 a_21788_30659.n6 VSS 3.71193f
C2906 a_21788_30659.n8 VSS 3.25297f
C2907 a_10114_45276.t3 VSS 0.102759f
C2908 a_10114_45276.t6 VSS 0.118353f
C2909 a_10114_45276.n1 VSS 1.22735f
C2910 a_10114_45276.n2 VSS 1.03928f
C2911 a_10114_45276.n3 VSS 0.533351f
C2912 a_10114_45276.n4 VSS 0.530824f
C2913 a_10114_45276.n5 VSS 0.180914f
C2914 a_5334_30651.n0 VSS 0.147836f
C2915 a_5334_30651.n1 VSS 0.206752f
C2916 a_5334_30651.t7 VSS 0.74063f
C2917 a_5334_30651.t6 VSS 0.743566f
C2918 a_5334_30651.n2 VSS 12.2363f
C2919 a_5334_30651.n3 VSS 6.94436f
C2920 a_5334_30651.n4 VSS 0.429467f
C2921 a_n99_45438.t1 VSS 0.136698f
C2922 a_n99_45438.n0 VSS 0.267231f
C2923 a_n99_45438.n1 VSS 0.102263f
C2924 a_n99_45438.n2 VSS 2.60765f
C2925 a_n99_45438.n3 VSS 0.29179f
C2926 a_n1925_47044.n2 VSS 0.694322f
C2927 a_n1925_47044.n3 VSS 0.364295f
C2928 a_n1925_47044.n4 VSS 17.524601f
C2929 a_n1925_47044.n5 VSS 0.203479f
C2930 a_n2497_47846.n1 VSS 0.204789f
C2931 a_n2497_47846.n3 VSS 1.52811f
C2932 a_n2497_47846.n4 VSS 0.177733f
C2933 a_n2497_47846.n5 VSS 0.127513f
C2934 a_5700_37509.t2 VSS 0.231968f
C2935 a_5700_37509.t5 VSS 0.231968f
C2936 a_5700_37509.t11 VSS 0.231968f
C2937 a_5700_37509.n0 VSS 0.462462f
C2938 a_5700_37509.t3 VSS 0.231968f
C2939 a_5700_37509.t12 VSS 0.231968f
C2940 a_5700_37509.n1 VSS 0.462027f
C2941 a_5700_37509.n2 VSS 0.180212f
C2942 a_5700_37509.t4 VSS 0.231968f
C2943 a_5700_37509.t13 VSS 0.231968f
C2944 a_5700_37509.n3 VSS 0.462027f
C2945 a_5700_37509.n4 VSS 0.127652f
C2946 a_5700_37509.t9 VSS 0.231968f
C2947 a_5700_37509.t1 VSS 0.231968f
C2948 a_5700_37509.n5 VSS 0.462027f
C2949 a_5700_37509.n6 VSS 0.692908f
C2950 a_5700_37509.t17 VSS 0.321046f
C2951 a_5700_37509.n7 VSS 0.200876f
C2952 a_5700_37509.n8 VSS 1.25965f
C2953 a_5700_37509.t16 VSS 0.319458f
C2954 a_5700_37509.n9 VSS 1.6989f
C2955 a_5700_37509.n10 VSS 3.49156f
C2956 a_5700_37509.t8 VSS 0.231968f
C2957 a_5700_37509.t10 VSS 0.231968f
C2958 a_5700_37509.n11 VSS 0.556177f
C2959 a_5700_37509.n12 VSS 1.34054f
C2960 a_5700_37509.t14 VSS 0.231968f
C2961 a_5700_37509.t0 VSS 0.231968f
C2962 a_5700_37509.n13 VSS 0.556177f
C2963 a_5700_37509.n14 VSS 0.827046f
C2964 a_5700_37509.t6 VSS 0.231968f
C2965 a_5700_37509.t7 VSS 0.231968f
C2966 a_5700_37509.n15 VSS 0.556177f
C2967 a_5700_37509.n16 VSS 1.57381f
C2968 a_5700_37509.n17 VSS 0.561806f
C2969 a_5700_37509.t15 VSS 0.231968f
C2970 a_6485_44582.n3 VSS 0.165972f
C2971 a_6485_44582.n5 VSS 1.01727f
C2972 a_6485_44582.n9 VSS 0.188689f
C2973 a_6485_44582.n12 VSS 0.393769f
C2974 a_6485_44582.n14 VSS 0.323069f
C2975 a_6485_44582.n16 VSS 0.292858f
C2976 a_6485_44582.n17 VSS 0.297837f
C2977 a_6485_44582.n20 VSS 0.496931f
C2978 a_6485_44582.n21 VSS 0.145879f
C2979 a_6485_44582.n23 VSS 0.107495f
C2980 SMPL.n2 VSS 0.178963f
C2981 SMPL.n5 VSS 0.116156f
C2982 SMPL.n6 VSS 0.166503f
C2983 SMPL.n16 VSS 4.62672f
C2984 SMPL.n26 VSS 1.38122f
C2985 SMPL.n27 VSS 5.50488f
C2986 a_18394_35068.n6 VSS 0.222907f
C2987 a_18394_35068.n8 VSS 0.354753f
C2988 a_18394_35068.n10 VSS 0.232182f
C2989 a_18394_35068.n13 VSS 0.11498f
C2990 a_19679_31459.t4 VSS 2.86393f
C2991 a_19679_31459.n0 VSS 0.184629f
C2992 a_19679_31459.n1 VSS 15.3684f
C2993 a_n2497_42870.n1 VSS 1.55473f
C2994 a_n2497_42870.n3 VSS 8.8673f
C2995 a_n2497_42870.n5 VSS 0.109195f
C2996 a_n2497_42870.n6 VSS 0.127284f
C2997 CAL_P.n0 VSS 1.91718f
C2998 CAL_P.t4 VSS 5.40604f
C2999 CAL_P.n1 VSS 3.80814f
C3000 CAL_P.t3 VSS 4.85086f
C3001 CAL_P.n2 VSS 3.90725f
C3002 CAL_P.t5 VSS 5.3968f
C3003 CAL_P.n3 VSS 2.03587f
C3004 CAL_P.n5 VSS 0.341488f
C3005 CAL_P.n6 VSS 0.539035f
C3006 CAL_P.t6 VSS 0.104492f
C3007 VIN_P.n0 VSS 0.249602f
C3008 VIN_P.n1 VSS 0.101674f
C3009 VIN_P.n9 VSS 0.105296f
C3010 VIN_P.n10 VSS 0.396356f
C3011 VIN_P.n11 VSS 0.467332f
C3012 VIN_P.t8 VSS 0.32821f
C3013 VIN_P.n12 VSS 0.781954f
C3014 VIN_P.t14 VSS 0.130802f
C3015 VIN_P.t13 VSS 0.12923f
C3016 VIN_P.n13 VSS 0.691453f
C3017 VIN_P.n14 VSS 2.29913f
C3018 C4_P_btm.t22 VSS 1.04503f
C3019 C4_P_btm.t1 VSS 0.216174f
C3020 C4_P_btm.t0 VSS 0.322262f
C3021 C4_P_btm.n0 VSS 1.66162f
C3022 C4_P_btm.n1 VSS 2.58914f
C3023 C4_P_btm.t2 VSS 0.141684f
C3024 C4_P_btm.n2 VSS 3.26208f
C3025 C4_P_btm.t8 VSS 0.92878f
C3026 C4_P_btm.n3 VSS 0.289222f
C3027 C4_P_btm.t18 VSS 0.92878f
C3028 C4_P_btm.t6 VSS 0.92878f
C3029 C4_P_btm.t3 VSS 0.96551f
C3030 C4_P_btm.t13 VSS 0.930343f
C3031 C4_P_btm.n4 VSS 0.464144f
C3032 C4_P_btm.t14 VSS 0.930343f
C3033 C4_P_btm.n5 VSS 0.322189f
C3034 C4_P_btm.t12 VSS 0.930343f
C3035 C4_P_btm.n6 VSS 0.330183f
C3036 C4_P_btm.n7 VSS 0.291856f
C3037 C4_P_btm.t15 VSS 0.927241f
C3038 C4_P_btm.n8 VSS 0.181129f
C3039 C4_P_btm.t20 VSS 0.927241f
C3040 C4_P_btm.n9 VSS 0.183763f
C3041 C4_P_btm.t17 VSS 0.927241f
C3042 C4_P_btm.n10 VSS 0.183763f
C3043 C4_P_btm.t21 VSS 0.927241f
C3044 C4_P_btm.n11 VSS 0.183763f
C3045 C4_P_btm.t9 VSS 0.927241f
C3046 C4_P_btm.n12 VSS 0.183763f
C3047 C4_P_btm.t19 VSS 0.927241f
C3048 C4_P_btm.n13 VSS 0.181129f
C3049 C4_P_btm.t7 VSS 0.92878f
C3050 C4_P_btm.n14 VSS 0.291856f
C3051 C4_P_btm.t11 VSS 0.930343f
C3052 C4_P_btm.n15 VSS 0.330183f
C3053 C4_P_btm.t10 VSS 0.92878f
C3054 C4_P_btm.n16 VSS 0.144381f
C3055 C4_P_btm.n17 VSS 0.209446f
C3056 C4_P_btm.t5 VSS 0.96551f
C3057 C4_P_btm.n18 VSS 0.351401f
C3058 C4_P_btm.n19 VSS 0.144381f
C3059 C4_P_btm.t16 VSS 0.92878f
C3060 C4_P_btm.n20 VSS 0.144381f
C3061 C4_P_btm.n21 VSS 0.217439f
C3062 C4_P_btm.t4 VSS 0.930343f
C3063 C4_P_btm.n22 VSS 0.575857f
C3064 a_4830_43958.t13 VSS 0.146639f
C3065 a_4830_43958.n2 VSS 0.987904f
C3066 a_4830_43958.n6 VSS 0.571077f
C3067 a_4830_43958.n8 VSS 0.486754f
C3068 a_4830_43958.n10 VSS 0.250992f
C3069 a_4830_43958.n11 VSS 0.622546f
C3070 a_4830_43958.n12 VSS 2.32045f
C3071 a_4830_43958.n14 VSS 0.26518f
C3072 a_4830_43958.n15 VSS 0.15367f
C3073 a_17564_32305.n0 VSS 0.112651f
C3074 a_17564_32305.t4 VSS 1.5128f
C3075 a_17564_32305.n1 VSS 15.853201f
C3076 a_17564_32305.n2 VSS 0.135534f
C3077 a_3754_38470.t1 VSS 0.367463f
C3078 a_3754_38470.n7 VSS 0.413441f
C3079 a_3754_38470.n8 VSS 0.933763f
C3080 a_n4515_30659.t17 VSS 0.550271f
C3081 a_n4515_30659.t19 VSS 0.550187f
C3082 a_n4515_30659.n0 VSS 0.406366f
C3083 a_n4515_30659.t5 VSS 0.550187f
C3084 a_n4515_30659.n1 VSS 0.206837f
C3085 a_n4515_30659.t12 VSS 0.550187f
C3086 a_n4515_30659.n2 VSS 0.206837f
C3087 a_n4515_30659.t14 VSS 0.550187f
C3088 a_n4515_30659.n3 VSS 0.206837f
C3089 a_n4515_30659.t18 VSS 0.550187f
C3090 a_n4515_30659.n4 VSS 0.206837f
C3091 a_n4515_30659.t6 VSS 0.550187f
C3092 a_n4515_30659.n5 VSS 0.206837f
C3093 a_n4515_30659.t11 VSS 0.550187f
C3094 a_n4515_30659.n6 VSS 0.206837f
C3095 a_n4515_30659.t4 VSS 0.550187f
C3096 a_n4515_30659.n7 VSS 0.206837f
C3097 a_n4515_30659.t7 VSS 0.550187f
C3098 a_n4515_30659.n8 VSS 0.206837f
C3099 a_n4515_30659.t13 VSS 0.550187f
C3100 a_n4515_30659.n9 VSS 0.206837f
C3101 a_n4515_30659.t15 VSS 0.550187f
C3102 a_n4515_30659.n10 VSS 0.206837f
C3103 a_n4515_30659.t9 VSS 0.550187f
C3104 a_n4515_30659.n11 VSS 0.206837f
C3105 a_n4515_30659.t10 VSS 0.550187f
C3106 a_n4515_30659.n12 VSS 0.206837f
C3107 a_n4515_30659.t8 VSS 0.550187f
C3108 a_n4515_30659.n13 VSS 0.20644f
C3109 a_n4515_30659.t16 VSS 0.550187f
C3110 a_n4515_30659.n14 VSS 2.44131f
C3111 a_n4515_30659.n16 VSS 1.83721f
C3112 a_5923_31099.n0 VSS 0.175913f
C3113 a_5923_31099.n1 VSS 0.199678f
C3114 a_5923_31099.t5 VSS 0.418293f
C3115 a_5923_31099.t7 VSS 0.389978f
C3116 a_5923_31099.n2 VSS 18.837599f
C3117 a_5923_31099.n3 VSS 10.578799f
C3118 a_5923_31099.n4 VSS 0.482005f
C3119 a_2424_46794.n6 VSS 0.356538f
C3120 a_2424_46794.n7 VSS 0.382728f
C3121 a_2424_46794.n9 VSS 1.57222f
C3122 a_2424_46794.n10 VSS 0.421737f
C3123 a_2424_46794.n11 VSS 0.109442f
C3124 a_1581_43806.n3 VSS 0.157021f
C3125 a_1581_43806.n9 VSS 0.81903f
C3126 a_1581_43806.n11 VSS 0.817122f
C3127 a_1581_43806.n12 VSS 0.816734f
C3128 a_1581_43806.n14 VSS 1.11042f
C3129 a_1581_43806.n15 VSS 1.17561f
C3130 a_1581_43806.n16 VSS 0.515292f
C3131 a_1581_43806.n17 VSS 0.105467f
C3132 a_1581_43806.n18 VSS 0.125105f
C3133 a_20647_31459.n0 VSS 0.174685f
C3134 a_20647_31459.t4 VSS 2.75242f
C3135 a_20647_31459.n1 VSS 15.4051f
C3136 RST_Z.t3 VSS 0.196434f
C3137 RST_Z.n0 VSS 1.74464f
C3138 RST_Z.n2 VSS 4.42662f
C3139 a_7029_44350.n0 VSS 0.61374f
C3140 a_7029_44350.n1 VSS 4.57868f
C3141 a_7029_44350.t1 VSS 0.140414f
C3142 a_7029_44350.n2 VSS 0.222062f
C3143 a_7557_43236.n5 VSS 0.521582f
C3144 a_7557_43236.n9 VSS 0.443597f
C3145 a_7557_43236.n13 VSS 0.360554f
C3146 a_7557_43236.n15 VSS 0.162092f
C3147 a_7557_43236.n19 VSS 0.101391f
C3148 a_7557_43236.n20 VSS 0.126076f
C3149 a_7557_43236.n21 VSS 0.264767f
C3150 a_13667_32299.n0 VSS 0.188178f
C3151 a_13667_32299.t4 VSS 2.35257f
C3152 a_13667_32299.n1 VSS 19.370802f
C3153 C1_N_btm.t5 VSS 1.55202f
C3154 C1_N_btm.t4 VSS 0.465838f
C3155 C1_N_btm.t6 VSS 0.31401f
C3156 C1_N_btm.n0 VSS 2.49999f
C3157 C1_N_btm.n1 VSS 3.88666f
C3158 C1_N_btm.t0 VSS 0.280658f
C3159 C1_N_btm.n2 VSS 4.85761f
C3160 C1_N_btm.t2 VSS 1.42799f
C3161 C1_N_btm.t1 VSS 1.35139f
C3162 C1_N_btm.n3 VSS 0.777183f
C3163 C1_N_btm.t3 VSS 1.35139f
C3164 C1_N_btm.n4 VSS 0.954486f
C3165 a_n2442_44350.n0 VSS 0.111988f
C3166 a_n2442_44350.t4 VSS 1.52924f
C3167 a_n2442_44350.n1 VSS 15.639299f
C3168 a_n2442_44350.n2 VSS 0.134737f
C3169 a_21276_30659.t7 VSS 1.29613f
C3170 a_21276_30659.t6 VSS 1.29593f
C3171 a_21276_30659.n1 VSS 0.960004f
C3172 a_21276_30659.t4 VSS 1.29593f
C3173 a_21276_30659.n2 VSS 0.486232f
C3174 a_21276_30659.t5 VSS 1.29593f
C3175 a_21276_30659.n3 VSS 6.15273f
C3176 a_21276_30659.n4 VSS 4.422009f
C3177 C4_N_btm.t0 VSS 1.04503f
C3178 C4_N_btm.t1 VSS 0.322262f
C3179 C4_N_btm.t3 VSS 0.216174f
C3180 C4_N_btm.n0 VSS 1.66162f
C3181 C4_N_btm.n1 VSS 2.58914f
C3182 C4_N_btm.t2 VSS 0.141684f
C3183 C4_N_btm.n2 VSS 3.26208f
C3184 C4_N_btm.t9 VSS 0.92878f
C3185 C4_N_btm.n3 VSS 0.289222f
C3186 C4_N_btm.t16 VSS 0.92878f
C3187 C4_N_btm.t20 VSS 0.96551f
C3188 C4_N_btm.t22 VSS 0.96551f
C3189 C4_N_btm.t10 VSS 0.930343f
C3190 C4_N_btm.n4 VSS 0.464144f
C3191 C4_N_btm.t5 VSS 0.930343f
C3192 C4_N_btm.n5 VSS 0.322189f
C3193 C4_N_btm.t14 VSS 0.930343f
C3194 C4_N_btm.n6 VSS 0.330183f
C3195 C4_N_btm.t17 VSS 0.92878f
C3196 C4_N_btm.n7 VSS 0.291856f
C3197 C4_N_btm.t11 VSS 0.927241f
C3198 C4_N_btm.n8 VSS 0.181129f
C3199 C4_N_btm.t18 VSS 0.927241f
C3200 C4_N_btm.n9 VSS 0.183763f
C3201 C4_N_btm.t7 VSS 0.927241f
C3202 C4_N_btm.n10 VSS 0.183763f
C3203 C4_N_btm.t19 VSS 0.927241f
C3204 C4_N_btm.n11 VSS 0.183763f
C3205 C4_N_btm.t8 VSS 0.927241f
C3206 C4_N_btm.n12 VSS 0.183763f
C3207 C4_N_btm.t4 VSS 0.927241f
C3208 C4_N_btm.n13 VSS 0.181129f
C3209 C4_N_btm.t15 VSS 0.92878f
C3210 C4_N_btm.n14 VSS 0.291856f
C3211 C4_N_btm.t13 VSS 0.930343f
C3212 C4_N_btm.n15 VSS 0.330183f
C3213 C4_N_btm.t12 VSS 0.92878f
C3214 C4_N_btm.n16 VSS 0.144381f
C3215 C4_N_btm.n17 VSS 0.209446f
C3216 C4_N_btm.n18 VSS 0.351401f
C3217 C4_N_btm.n19 VSS 0.144381f
C3218 C4_N_btm.t6 VSS 0.92878f
C3219 C4_N_btm.n20 VSS 0.144381f
C3220 C4_N_btm.n21 VSS 0.217439f
C3221 C4_N_btm.t21 VSS 0.930343f
C3222 C4_N_btm.n22 VSS 0.575857f
C3223 a_14601_32299.n0 VSS 0.105763f
C3224 a_14601_32299.t4 VSS 0.167391f
C3225 a_14601_32299.t5 VSS 0.19248f
C3226 a_14601_32299.n1 VSS 4.683259f
C3227 a_14601_32299.n2 VSS 13.4494f
C3228 a_14601_32299.n3 VSS 0.127248f
C3229 a_n2293_45956.n2 VSS 1.27513f
C3230 a_n2293_45956.n3 VSS 0.371302f
C3231 a_n2293_45956.n4 VSS 13.1905f
C3232 a_n2293_45956.n5 VSS 0.127379f
C3233 a_15549_47044.n4 VSS 1.46657f
C3234 a_15549_47044.n6 VSS 0.120859f
C3235 a_15549_47044.n7 VSS 1.1789f
C3236 a_15549_47044.n8 VSS 0.768485f
C3237 a_15549_47044.n9 VSS 0.180739f
C3238 a_5840_42718.n0 VSS 0.163756f
C3239 a_5840_42718.n1 VSS 0.193658f
C3240 a_5840_42718.t4 VSS 0.38234f
C3241 a_5840_42718.t6 VSS 0.367953f
C3242 a_5840_42718.n2 VSS 16.9332f
C3243 a_5840_42718.n3 VSS 9.36375f
C3244 a_5840_42718.n4 VSS 0.506496f
C3245 a_n2103_44868.n0 VSS 0.352076f
C3246 a_n2103_44868.n2 VSS 0.964184f
C3247 a_n2103_44868.n3 VSS 11.976f
C3248 a_n2103_44868.n7 VSS 0.131656f
C3249 a_n2103_44868.n9 VSS 0.236252f
C3250 a_n2810_43806.n0 VSS 0.114759f
C3251 a_n2810_43806.t5 VSS 0.177594f
C3252 a_n2810_43806.t4 VSS 0.204212f
C3253 a_n2810_43806.n1 VSS 4.52432f
C3254 a_n2810_43806.n2 VSS 13.2673f
C3255 a_n2810_43806.n3 VSS 0.126762f
C3256 a_12651_44576.n2 VSS 0.148391f
C3257 a_12651_44576.n11 VSS 0.32195f
C3258 a_12651_44576.n14 VSS 0.146408f
C3259 a_12651_44576.n15 VSS 0.531274f
C3260 a_12651_44576.n16 VSS 0.452312f
C3261 a_12651_44576.n17 VSS 0.231256f
C3262 a_12651_44576.n18 VSS 0.322683f
C3263 a_12651_44576.n19 VSS 0.174153f
C3264 a_12651_44576.n21 VSS 0.362223f
C3265 a_885_44868.n5 VSS 0.174669f
C3266 a_885_44868.n9 VSS 0.116255f
C3267 a_885_44868.n10 VSS 0.164069f
C3268 a_885_44868.n12 VSS 0.116255f
C3269 a_885_44868.n13 VSS 0.181619f
C3270 a_885_44868.n14 VSS 0.116255f
C3271 a_885_44868.n16 VSS 0.346154f
C3272 a_885_44868.n18 VSS 0.805002f
C3273 a_885_44868.n19 VSS 0.229704f
C3274 a_885_44868.n20 VSS 0.228704f
C3275 a_885_44868.n22 VSS 0.490384f
C3276 a_885_44868.n24 VSS 0.116255f
C3277 a_885_44868.n25 VSS 0.304753f
C3278 a_885_44868.n26 VSS 0.124688f
C3279 a_885_44868.n28 VSS 0.190286f
C3280 a_885_44868.n29 VSS 0.591596f
C3281 a_885_44868.n31 VSS 0.116255f
C3282 a_885_44868.n32 VSS 0.164069f
C3283 a_885_44868.n33 VSS 0.328087f
C3284 a_885_44868.n34 VSS 0.463013f
C3285 a_885_44868.n36 VSS 0.122667f
C3286 C5_P_btm.t0 VSS 0.800169f
C3287 C5_P_btm.t37 VSS 0.248689f
C3288 C5_P_btm.t2 VSS 0.166821f
C3289 C5_P_btm.n0 VSS 1.26557f
C3290 C5_P_btm.n1 VSS 1.978f
C3291 C5_P_btm.t1 VSS 0.107115f
C3292 C5_P_btm.n2 VSS 2.60859f
C3293 C5_P_btm.t19 VSS 0.716737f
C3294 C5_P_btm.n3 VSS 0.218419f
C3295 C5_P_btm.t36 VSS 0.716737f
C3296 C5_P_btm.n14 VSS 0.131769f
C3297 C5_P_btm.n15 VSS 0.1256f
C3298 C5_P_btm.n16 VSS 0.1256f
C3299 C5_P_btm.t12 VSS 0.716737f
C3300 C5_P_btm.n19 VSS 0.218419f
C3301 C5_P_btm.t18 VSS 0.646259f
C3302 C5_P_btm.n21 VSS 0.120948f
C3303 C5_P_btm.t15 VSS 0.646259f
C3304 C5_P_btm.n24 VSS 0.120948f
C3305 C5_P_btm.t17 VSS 0.716737f
C3306 C5_P_btm.n26 VSS 0.218419f
C3307 C5_P_btm.n27 VSS 0.131769f
C3308 C5_P_btm.t13 VSS 0.646259f
C3309 C5_P_btm.n31 VSS 0.120948f
C3310 C5_P_btm.t35 VSS 0.646259f
C3311 C5_P_btm.n34 VSS 0.120948f
C3312 C5_P_btm.t9 VSS 0.646259f
C3313 C5_P_btm.n37 VSS 0.120948f
C3314 C5_P_btm.t30 VSS 0.646259f
C3315 C5_P_btm.n40 VSS 0.120948f
C3316 C5_P_btm.t26 VSS 0.646259f
C3317 C5_P_btm.n43 VSS 0.120948f
C3318 C5_P_btm.t27 VSS 0.646259f
C3319 C5_P_btm.n46 VSS 0.120948f
C3320 C5_P_btm.t20 VSS 0.646259f
C3321 C5_P_btm.n49 VSS 0.120948f
C3322 C5_P_btm.t5 VSS 0.646259f
C3323 C5_P_btm.n52 VSS 0.120948f
C3324 C5_P_btm.n54 VSS 0.218419f
C3325 C5_P_btm.t3 VSS 0.745082f
C3326 C5_P_btm.t16 VSS 0.717943f
C3327 C5_P_btm.n55 VSS 0.358179f
C3328 C5_P_btm.t32 VSS 0.717943f
C3329 C5_P_btm.n56 VSS 0.248633f
C3330 C5_P_btm.t28 VSS 0.717943f
C3331 C5_P_btm.n57 VSS 0.248633f
C3332 C5_P_btm.t7 VSS 0.717943f
C3333 C5_P_btm.n58 VSS 0.248633f
C3334 C5_P_btm.n59 VSS 0.167798f
C3335 C5_P_btm.t22 VSS 0.716737f
C3336 C5_P_btm.n60 VSS 0.106646f
C3337 C5_P_btm.t6 VSS 0.646259f
C3338 C5_P_btm.n62 VSS 0.120948f
C3339 C5_P_btm.t11 VSS 0.646259f
C3340 C5_P_btm.n65 VSS 0.120948f
C3341 C5_P_btm.t31 VSS 0.646259f
C3342 C5_P_btm.n68 VSS 0.120948f
C3343 C5_P_btm.t25 VSS 0.646259f
C3344 C5_P_btm.n71 VSS 0.120948f
C3345 C5_P_btm.t34 VSS 0.646259f
C3346 C5_P_btm.n74 VSS 0.120948f
C3347 C5_P_btm.t14 VSS 0.646259f
C3348 C5_P_btm.n77 VSS 0.120948f
C3349 C5_P_btm.t21 VSS 0.646259f
C3350 C5_P_btm.n80 VSS 0.120948f
C3351 C5_P_btm.t24 VSS 0.646259f
C3352 C5_P_btm.n83 VSS 0.120948f
C3353 C5_P_btm.t23 VSS 0.716737f
C3354 C5_P_btm.n85 VSS 0.106646f
C3355 C5_P_btm.n86 VSS 0.167798f
C3356 C5_P_btm.t10 VSS 0.717943f
C3357 C5_P_btm.n87 VSS 0.248633f
C3358 C5_P_btm.t29 VSS 0.717943f
C3359 C5_P_btm.n88 VSS 0.248633f
C3360 C5_P_btm.t33 VSS 0.717943f
C3361 C5_P_btm.n89 VSS 0.248633f
C3362 C5_P_btm.t8 VSS 0.717943f
C3363 C5_P_btm.n90 VSS 0.248633f
C3364 C5_P_btm.t4 VSS 0.717943f
C3365 C5_P_btm.n91 VSS 0.429614f
C3366 EN_COMP.n1 VSS 1.9035f
C3367 EN_COMP.n4 VSS 0.731672f
C3368 EN_COMP.n5 VSS 9.23273f
C3369 a_14297_32299.t4 VSS 2.41824f
C3370 a_14297_32299.n0 VSS 0.198795f
C3371 a_14297_32299.n1 VSS 18.978199f
C3372 a_n2293_45420.n1 VSS 0.199643f
C3373 a_n2293_45420.n3 VSS 0.79461f
C3374 a_n2293_45420.n4 VSS 13.5659f
C3375 a_n2293_45420.n5 VSS 0.218521f
C3376 C0_N_btm.t0 VSS 1.37053f
C3377 C0_N_btm.t5 VSS 0.408265f
C3378 C0_N_btm.t2 VSS 0.275201f
C3379 C0_N_btm.n0 VSS 2.21668f
C3380 C0_N_btm.n1 VSS 3.36018f
C3381 C0_N_btm.t1 VSS 0.19597f
C3382 C0_N_btm.n2 VSS 3.88487f
C3383 C0_N_btm.t3 VSS 1.2515f
C3384 C0_N_btm.t4 VSS 1.18437f
C3385 C0_N_btm.n3 VSS 1.08331f
C3386 a_n2810_44350.n0 VSS 0.118527f
C3387 a_n2810_44350.t4 VSS 0.762664f
C3388 a_n2810_44350.t5 VSS 0.784531f
C3389 a_n2810_44350.n1 VSS 4.45898f
C3390 a_n2810_44350.n2 VSS 13.053201f
C3391 a_n2810_44350.n3 VSS 0.130925f
C3392 a_134_42718.n0 VSS 0.135553f
C3393 a_134_42718.n1 VSS 0.172873f
C3394 a_134_42718.t6 VSS 0.28866f
C3395 a_134_42718.t5 VSS 0.291541f
C3396 a_134_42718.n2 VSS 14.2708f
C3397 a_134_42718.n3 VSS 9.24833f
C3398 a_134_42718.n4 VSS 0.470382f
C3399 a_135_43540.n8 VSS 0.110143f
C3400 a_135_43540.n11 VSS 0.176325f
C3401 a_135_43540.n14 VSS 0.120668f
C3402 a_135_43540.n15 VSS 0.124919f
C3403 a_135_43540.n18 VSS 0.116768f
C3404 a_135_43540.n21 VSS 0.161146f
C3405 a_135_43540.n24 VSS 0.174329f
C3406 a_135_43540.n27 VSS 0.172026f
C3407 a_135_43540.n30 VSS 0.110068f
C3408 a_135_43540.n32 VSS 0.134284f
C3409 a_135_43540.n33 VSS 0.155871f
C3410 a_135_43540.n34 VSS 0.134306f
C3411 a_135_43540.n37 VSS 0.109841f
C3412 a_135_43540.n38 VSS 0.210749f
C3413 a_135_43540.n39 VSS 0.105947f
C3414 a_135_43540.n40 VSS 0.305114f
C3415 a_135_43540.n42 VSS 0.29532f
C3416 a_135_43540.n43 VSS 0.1315f
C3417 a_1736_39043.t5 VSS 0.129773f
C3418 a_1736_39043.n1 VSS 0.793746f
C3419 a_1736_39043.n2 VSS 0.356005f
C3420 a_1736_39043.n3 VSS 0.354214f
C3421 a_1736_39043.t2 VSS 0.31643f
C3422 a_1736_39043.n4 VSS 0.586153f
C3423 a_3990_30651.n1 VSS 0.162922f
C3424 a_3990_30651.t6 VSS 0.424791f
C3425 a_3990_30651.t8 VSS 0.437457f
C3426 a_3990_30651.t14 VSS 0.425508f
C3427 a_3990_30651.t16 VSS 0.424791f
C3428 a_3990_30651.t19 VSS 0.425508f
C3429 a_3990_30651.t11 VSS 0.424791f
C3430 a_3990_30651.t5 VSS 0.425508f
C3431 a_3990_30651.n2 VSS 0.195263f
C3432 a_3990_30651.t4 VSS 0.424791f
C3433 a_3990_30651.n3 VSS 0.209972f
C3434 a_3990_30651.n4 VSS 0.280384f
C3435 a_3990_30651.n5 VSS 0.218432f
C3436 a_3990_30651.n6 VSS 0.195263f
C3437 a_3990_30651.n7 VSS 0.218432f
C3438 a_3990_30651.n8 VSS 0.195263f
C3439 a_3990_30651.n9 VSS 0.385847f
C3440 a_3990_30651.n10 VSS 1.36362f
C3441 a_3990_30651.n11 VSS 0.162922f
C3442 a_3990_30651.t9 VSS 0.424791f
C3443 a_3990_30651.t15 VSS 0.425508f
C3444 a_3990_30651.t7 VSS 0.424791f
C3445 a_3990_30651.t10 VSS 0.425508f
C3446 a_3990_30651.t18 VSS 0.424791f
C3447 a_3990_30651.t12 VSS 0.425508f
C3448 a_3990_30651.n12 VSS 0.195263f
C3449 a_3990_30651.t21 VSS 0.424791f
C3450 a_3990_30651.n13 VSS 0.209972f
C3451 a_3990_30651.n14 VSS 0.280384f
C3452 a_3990_30651.n15 VSS 0.218432f
C3453 a_3990_30651.n16 VSS 0.195263f
C3454 a_3990_30651.n17 VSS 0.218432f
C3455 a_3990_30651.n18 VSS 0.195263f
C3456 a_3990_30651.t20 VSS 0.437457f
C3457 a_3990_30651.n19 VSS 0.385847f
C3458 a_3990_30651.n20 VSS 1.50787f
C3459 a_3990_30651.n21 VSS 6.13436f
C3460 a_3990_30651.n22 VSS 0.118412f
C3461 a_3990_30651.n23 VSS 4.22249f
C3462 a_3990_30651.n24 VSS 0.376512f
C3463 a_11455_44576.n2 VSS 0.116887f
C3464 a_11455_44576.n12 VSS 0.239269f
C3465 a_11455_44576.n13 VSS 0.166537f
C3466 a_11455_44576.n15 VSS 0.252357f
C3467 a_11455_44576.n16 VSS 0.162404f
C3468 a_11455_44576.n17 VSS 0.108874f
C3469 a_11455_44576.n19 VSS 0.144912f
C3470 a_11455_44576.n20 VSS 0.347761f
C3471 a_11455_44576.n21 VSS 0.246469f
C3472 a_n1732_35090.n6 VSS 0.223004f
C3473 a_n1732_35090.n8 VSS 0.354792f
C3474 a_n1732_35090.n10 VSS 0.232088f
C3475 a_n1732_35090.n13 VSS 0.11498f
C3476 a_n2103_45412.n1 VSS 0.279597f
C3477 a_n2103_45412.n3 VSS 2.06353f
C3478 a_n2103_45412.n4 VSS 9.063901f
C3479 a_n2103_45412.n6 VSS 0.124191f
C3480 a_n2103_45412.n8 VSS 0.165552f
C3481 a_n2103_45412.n9 VSS 0.297076f
C3482 a_n2293_47044.n2 VSS 0.1953f
C3483 a_n2293_47044.n3 VSS 1.06479f
C3484 a_n2293_47044.n4 VSS 12.1792f
C3485 a_n2293_47044.n5 VSS 0.126855f
C3486 EN_VIN_BSTR_P.n3 VSS 0.302094f
C3487 EN_VIN_BSTR_P.t1 VSS 0.107284f
C3488 EN_VIN_BSTR_P.t0 VSS 0.110779f
C3489 EN_VIN_BSTR_P.t2 VSS 0.107415f
C3490 EN_VIN_BSTR_P.n6 VSS 0.284789f
C3491 EN_VIN_BSTR_P.n7 VSS 0.170171f
C3492 EN_VIN_BSTR_P.n8 VSS 0.15757f
C3493 EN_VIN_BSTR_P.n9 VSS 0.114651f
C3494 EN_VIN_BSTR_P.n18 VSS 0.351313f
C3495 EN_VIN_BSTR_P.n21 VSS 0.488964f
C3496 a_18314_32299.n1 VSS 0.167814f
C3497 a_18314_32299.t11 VSS 0.513501f
C3498 a_18314_32299.t4 VSS 0.528224f
C3499 a_18314_32299.t6 VSS 0.514801f
C3500 a_18314_32299.t10 VSS 0.513501f
C3501 a_18314_32299.t7 VSS 0.514801f
C3502 a_18314_32299.t8 VSS 0.513501f
C3503 a_18314_32299.t9 VSS 0.514801f
C3504 a_18314_32299.n2 VSS 0.246764f
C3505 a_18314_32299.t5 VSS 0.513501f
C3506 a_18314_32299.n3 VSS 0.25509f
C3507 a_18314_32299.n4 VSS 0.297596f
C3508 a_18314_32299.n5 VSS 0.266526f
C3509 a_18314_32299.n6 VSS 0.246764f
C3510 a_18314_32299.n7 VSS 0.266526f
C3511 a_18314_32299.n8 VSS 0.246764f
C3512 a_18314_32299.n9 VSS 0.477018f
C3513 a_18314_32299.n10 VSS 6.29784f
C3514 a_18314_32299.n11 VSS 5.40405f
C3515 a_21020_30659.n0 VSS 0.145982f
C3516 a_21020_30659.t5 VSS 1.64675f
C3517 a_21020_30659.t4 VSS 1.64697f
C3518 a_21020_30659.n1 VSS 8.14992f
C3519 a_21020_30659.n2 VSS 6.48659f
C3520 a_14766_45596.n1 VSS 0.135045f
C3521 a_14766_45596.n2 VSS 0.169983f
C3522 a_14766_45596.n4 VSS 0.768458f
C3523 a_14766_45596.n6 VSS 0.443285f
C3524 a_14766_45596.n7 VSS 0.348791f
C3525 a_14766_45596.n8 VSS 1.16104f
C3526 a_14766_45596.n9 VSS 0.755026f
C3527 a_1203_42692.n6 VSS 0.565577f
C3528 a_1203_42692.n7 VSS 0.231614f
C3529 a_1203_42692.n9 VSS 0.421798f
C3530 a_1203_42692.n10 VSS 0.358609f
C3531 a_1203_42692.n12 VSS 0.307134f
C3532 a_1203_42692.n14 VSS 0.303515f
C3533 a_1203_42692.n16 VSS 0.274587f
C3534 a_1203_42692.n18 VSS 0.462268f
C3535 a_1203_42692.n20 VSS 0.301331f
C3536 a_1203_42692.n22 VSS 0.29346f
C3537 a_1203_42692.n24 VSS 0.508659f
C3538 a_1203_42692.n25 VSS 0.181426f
C3539 a_1203_42692.n28 VSS 0.131245f
C3540 a_2587_44868.n2 VSS 0.171835f
C3541 a_2587_44868.n4 VSS 0.133805f
C3542 a_2587_44868.n17 VSS 0.258017f
C3543 a_2587_44868.n21 VSS 0.327028f
C3544 a_2587_44868.n22 VSS 0.884245f
C3545 a_2587_44868.n23 VSS 0.712002f
C3546 a_2587_44868.n25 VSS 0.380054f
C3547 a_2587_44868.n26 VSS 0.736337f
C3548 a_2587_44868.n28 VSS 1.34541f
C3549 a_2587_44868.n30 VSS 1.32246f
C3550 a_2587_44868.n31 VSS 1.01568f
C3551 a_2587_44868.n32 VSS 0.177342f
C3552 C3_P_btm.t1 VSS 0.973133f
C3553 C3_P_btm.t2 VSS 0.297776f
C3554 C3_P_btm.t12 VSS 0.199749f
C3555 C3_P_btm.n0 VSS 1.55495f
C3556 C3_P_btm.n1 VSS 2.46584f
C3557 C3_P_btm.t0 VSS 0.151676f
C3558 C3_P_btm.n2 VSS 2.91699f
C3559 C3_P_btm.t11 VSS 0.858208f
C3560 C3_P_btm.t6 VSS 0.881786f
C3561 C3_P_btm.t5 VSS 0.856786f
C3562 C3_P_btm.n3 VSS 0.286809f
C3563 C3_P_btm.t10 VSS 0.856786f
C3564 C3_P_btm.n4 VSS 0.1698f
C3565 C3_P_btm.t9 VSS 0.856786f
C3566 C3_P_btm.n5 VSS 0.1698f
C3567 C3_P_btm.t4 VSS 0.856786f
C3568 C3_P_btm.n6 VSS 0.167366f
C3569 C3_P_btm.n7 VSS 0.26968f
C3570 C3_P_btm.t8 VSS 0.859652f
C3571 C3_P_btm.n8 VSS 0.305094f
C3572 C3_P_btm.t7 VSS 0.859652f
C3573 C3_P_btm.n9 VSS 0.297708f
C3574 C3_P_btm.t3 VSS 0.859652f
C3575 C3_P_btm.n10 VSS 0.624475f
C3576 a_4000_42718.n0 VSS 0.120726f
C3577 a_4000_42718.n1 VSS 0.14354f
C3578 a_4000_42718.t7 VSS 0.27359f
C3579 a_4000_42718.t6 VSS 0.267611f
C3580 a_4000_42718.n2 VSS 11.856799f
C3581 a_4000_42718.n3 VSS 6.47446f
C3582 a_4000_42718.n4 VSS 0.376629f
C3583 a_1847_45528.n13 VSS 0.198756f
C3584 a_1847_45528.n14 VSS 0.227493f
C3585 a_1847_45528.n17 VSS 0.180802f
C3586 a_1847_45528.n18 VSS 0.211478f
C3587 a_1847_45528.n19 VSS 0.127044f
C3588 a_1847_45528.n20 VSS 0.107728f
C3589 a_1847_45528.n21 VSS 0.187819f
C3590 a_1847_45528.n22 VSS 0.254942f
C3591 a_2755_43494.n7 VSS 0.554667f
C3592 a_2755_43494.n9 VSS 0.457027f
C3593 a_2755_43494.n10 VSS 0.468326f
C3594 a_2755_43494.n12 VSS 0.423555f
C3595 a_2755_43494.n13 VSS 0.451138f
C3596 a_2755_43494.n14 VSS 0.441349f
C3597 a_2755_43494.n15 VSS 0.625472f
C3598 a_2755_43494.n17 VSS 0.396877f
C3599 a_2755_43494.n18 VSS 0.451015f
C3600 a_2755_43494.n20 VSS 0.210066f
C3601 a_n1827_44324.n1 VSS 1.95629f
C3602 a_n1827_44324.n3 VSS 0.435098f
C3603 a_n1827_44324.n4 VSS 9.722321f
C3604 a_n1827_44324.n5 VSS 0.177895f
C3605 a_11206_38545.t3 VSS 1.21993f
C3606 a_11206_38545.t2 VSS 1.02548f
C3607 a_11206_38545.n0 VSS 2.85069f
C3608 a_11206_38545.t1 VSS 1.02548f
C3609 a_11206_38545.n1 VSS 2.55854f
C3610 a_11206_38545.n2 VSS 0.157657f
C3611 a_7754_40130.n0 VSS 0.22704f
C3612 a_7754_40130.n1 VSS 0.230022f
C3613 a_7754_40130.n2 VSS 0.21778f
C3614 a_7754_40130.n3 VSS 0.199574f
C3615 a_7754_40130.n4 VSS 0.230022f
C3616 a_7754_40130.n5 VSS 0.230022f
C3617 a_7754_40130.t12 VSS 0.441623f
C3618 a_7754_40130.n6 VSS 0.436037f
C3619 a_7754_40130.t6 VSS 0.44132f
C3620 a_7754_40130.n7 VSS 0.436037f
C3621 a_7754_40130.t7 VSS 0.44132f
C3622 a_7754_40130.n8 VSS 0.230022f
C3623 a_7754_40130.n9 VSS 0.230022f
C3624 a_7754_40130.t5 VSS 0.44132f
C3625 a_7754_40130.n10 VSS 0.230022f
C3626 a_7754_40130.t15 VSS 0.44132f
C3627 a_7754_40130.n11 VSS 0.230022f
C3628 a_7754_40130.n12 VSS 0.230022f
C3629 a_7754_40130.t10 VSS 0.44132f
C3630 a_7754_40130.n13 VSS 0.230022f
C3631 a_7754_40130.t1 VSS 0.44132f
C3632 a_7754_40130.n14 VSS 0.199574f
C3633 a_7754_40130.n15 VSS 0.11668f
C3634 a_7754_40130.t2 VSS 0.33407f
C3635 a_7754_40130.n16 VSS 0.396147f
C3636 a_7754_40130.n17 VSS 0.116902f
C3637 a_7754_40130.t8 VSS 0.44132f
C3638 a_7754_40130.n18 VSS 0.21778f
C3639 a_7754_40130.n19 VSS 0.230022f
C3640 a_7754_40130.t14 VSS 0.44132f
C3641 a_7754_40130.n20 VSS 0.230022f
C3642 a_7754_40130.t4 VSS 0.44132f
C3643 a_7754_40130.n21 VSS 0.230022f
C3644 a_7754_40130.n22 VSS 0.230022f
C3645 a_7754_40130.t13 VSS 0.44132f
C3646 a_7754_40130.n23 VSS 0.230022f
C3647 a_7754_40130.t9 VSS 0.44132f
C3648 a_7754_40130.n24 VSS 0.434782f
C3649 a_7754_40130.t11 VSS 0.441479f
C3650 a_7754_40130.n25 VSS 0.361405f
C3651 a_7754_40130.n26 VSS 0.926274f
C3652 VIN_N.n0 VSS 0.191386f
C3653 VIN_N.n10 VSS 0.303912f
C3654 VIN_N.n11 VSS 0.358334f
C3655 VIN_N.t4 VSS 0.25166f
C3656 VIN_N.n12 VSS 0.599576f
C3657 VIN_N.t15 VSS 0.100295f
C3658 VIN_N.n13 VSS 0.530178f
C3659 VIN_N.n14 VSS 1.76056f
C3660 EN_VIN_BSTR_N.t4 VSS 0.110775f
C3661 EN_VIN_BSTR_N.t6 VSS 0.107415f
C3662 EN_VIN_BSTR_N.n0 VSS 0.284793f
C3663 EN_VIN_BSTR_N.t5 VSS 0.107284f
C3664 EN_VIN_BSTR_N.n1 VSS 0.170171f
C3665 EN_VIN_BSTR_N.n5 VSS 0.302093f
C3666 EN_VIN_BSTR_N.n8 VSS 0.158258f
C3667 EN_VIN_BSTR_N.n9 VSS 0.114651f
C3668 EN_VIN_BSTR_N.n18 VSS 0.351313f
C3669 EN_VIN_BSTR_N.n21 VSS 0.488519f
C3670 C6_P_btm.t71 VSS 1.04079f
C3671 C6_P_btm.n0 VSS 0.153224f
C3672 C6_P_btm.n2 VSS 0.837749f
C3673 C6_P_btm.n3 VSS 1.30605f
C3674 C6_P_btm.n4 VSS 1.89867f
C3675 C6_P_btm.n5 VSS 0.115577f
C3676 C6_P_btm.n6 VSS 0.115577f
C3677 C6_P_btm.n7 VSS 0.115577f
C3678 C6_P_btm.t13 VSS 0.512523f
C3679 C6_P_btm.n8 VSS 0.119988f
C3680 C6_P_btm.t11 VSS 0.512523f
C3681 C6_P_btm.n20 VSS 0.159599f
C3682 C6_P_btm.t14 VSS 0.512523f
C3683 C6_P_btm.n21 VSS 0.159599f
C3684 C6_P_btm.t39 VSS 0.512523f
C3685 C6_P_btm.n28 VSS 0.115577f
C3686 C6_P_btm.n34 VSS 0.115577f
C3687 C6_P_btm.n35 VSS 0.115577f
C3688 C6_P_btm.t7 VSS 0.512523f
C3689 C6_P_btm.t1 VSS 0.532791f
C3690 C6_P_btm.n36 VSS 0.193911f
C3691 C6_P_btm.t3 VSS 0.532791f
C3692 C6_P_btm.t59 VSS 0.512523f
C3693 C6_P_btm.t31 VSS 0.512523f
C3694 C6_P_btm.n39 VSS 0.193911f
C3695 C6_P_btm.n40 VSS 0.115577f
C3696 C6_P_btm.t61 VSS 0.512523f
C3697 C6_P_btm.t36 VSS 0.512523f
C3698 C6_P_btm.n43 VSS 0.115577f
C3699 C6_P_btm.t18 VSS 0.512523f
C3700 C6_P_btm.t64 VSS 0.512523f
C3701 C6_P_btm.n46 VSS 0.115577f
C3702 C6_P_btm.n47 VSS 0.115577f
C3703 C6_P_btm.t67 VSS 0.512523f
C3704 C6_P_btm.n50 VSS 0.115577f
C3705 C6_P_btm.t49 VSS 0.512523f
C3706 C6_P_btm.t27 VSS 0.512523f
C3707 C6_P_btm.n53 VSS 0.115577f
C3708 C6_P_btm.n54 VSS 0.115577f
C3709 C6_P_btm.t65 VSS 0.512523f
C3710 C6_P_btm.t38 VSS 0.512523f
C3711 C6_P_btm.n57 VSS 0.115577f
C3712 C6_P_btm.t42 VSS 0.512523f
C3713 C6_P_btm.t6 VSS 0.462125f
C3714 C6_P_btm.t51 VSS 0.462125f
C3715 C6_P_btm.t45 VSS 0.462125f
C3716 C6_P_btm.t55 VSS 0.512523f
C3717 C6_P_btm.n69 VSS 0.109928f
C3718 C6_P_btm.t52 VSS 0.462125f
C3719 C6_P_btm.t32 VSS 0.462125f
C3720 C6_P_btm.t41 VSS 0.462125f
C3721 C6_P_btm.t30 VSS 0.462125f
C3722 C6_P_btm.t47 VSS 0.462125f
C3723 C6_P_btm.t8 VSS 0.462125f
C3724 C6_P_btm.t43 VSS 0.462125f
C3725 C6_P_btm.t54 VSS 0.462125f
C3726 C6_P_btm.t35 VSS 0.512523f
C3727 C6_P_btm.n100 VSS 0.119988f
C3728 C6_P_btm.n101 VSS 0.156187f
C3729 C6_P_btm.t22 VSS 0.462125f
C3730 C6_P_btm.t25 VSS 0.462125f
C3731 C6_P_btm.t63 VSS 0.462125f
C3732 C6_P_btm.t12 VSS 0.462125f
C3733 C6_P_btm.t26 VSS 0.462125f
C3734 C6_P_btm.t17 VSS 0.462125f
C3735 C6_P_btm.t5 VSS 0.462125f
C3736 C6_P_btm.t21 VSS 0.462125f
C3737 C6_P_btm.t9 VSS 0.462125f
C3738 C6_P_btm.t48 VSS 0.462125f
C3739 C6_P_btm.t53 VSS 0.462125f
C3740 C6_P_btm.t33 VSS 0.512523f
C3741 C6_P_btm.n136 VSS 0.156187f
C3742 C6_P_btm.t10 VSS 0.462125f
C3743 C6_P_btm.t20 VSS 0.512523f
C3744 C6_P_btm.t66 VSS 0.462125f
C3745 C6_P_btm.t46 VSS 0.462125f
C3746 C6_P_btm.t68 VSS 0.462125f
C3747 C6_P_btm.t40 VSS 0.462125f
C3748 C6_P_btm.t50 VSS 0.512523f
C3749 C6_P_btm.n154 VSS 0.109928f
C3750 C6_P_btm.t28 VSS 0.462125f
C3751 C6_P_btm.t56 VSS 0.462125f
C3752 C6_P_btm.t37 VSS 0.462125f
C3753 C6_P_btm.t57 VSS 0.512523f
C3754 C6_P_btm.n165 VSS 0.115577f
C3755 C6_P_btm.t24 VSS 0.512523f
C3756 C6_P_btm.t60 VSS 0.512523f
C3757 C6_P_btm.n168 VSS 0.115577f
C3758 C6_P_btm.n169 VSS 0.115577f
C3759 C6_P_btm.t58 VSS 0.512523f
C3760 C6_P_btm.n172 VSS 0.115577f
C3761 C6_P_btm.t16 VSS 0.512523f
C3762 C6_P_btm.t62 VSS 0.512523f
C3763 C6_P_btm.n175 VSS 0.115577f
C3764 C6_P_btm.n176 VSS 0.115577f
C3765 C6_P_btm.t15 VSS 0.512523f
C3766 C6_P_btm.t23 VSS 0.512523f
C3767 C6_P_btm.n179 VSS 0.115577f
C3768 C6_P_btm.t19 VSS 0.512523f
C3769 C6_P_btm.t29 VSS 0.512523f
C3770 C6_P_btm.n182 VSS 0.115577f
C3771 C6_P_btm.t2 VSS 0.532791f
C3772 C6_P_btm.n183 VSS 0.193911f
C3773 C6_P_btm.t34 VSS 0.512523f
C3774 C6_P_btm.t44 VSS 0.512523f
C3775 C6_P_btm.n186 VSS 0.115577f
C3776 C6_P_btm.t4 VSS 0.513385f
C3777 C6_P_btm.n187 VSS 0.294937f
C3778 a_n2293_46508.n2 VSS 0.232868f
C3779 a_n2293_46508.n3 VSS 0.529763f
C3780 a_n2293_46508.n4 VSS 10.2622f
C3781 a_n2293_46508.n5 VSS 0.151929f
C3782 a_15163_45670.n1 VSS 0.107375f
C3783 a_15163_45670.n2 VSS 0.502258f
C3784 a_15163_45670.n5 VSS 0.786688f
C3785 a_15163_45670.n6 VSS 0.403102f
C3786 a_15163_45670.n8 VSS 1.87357f
C3787 a_15163_45670.n9 VSS 0.805266f
C3788 C1_P_btm.t6 VSS 1.55202f
C3789 C1_P_btm.t1 VSS 0.465838f
C3790 C1_P_btm.t5 VSS 0.31401f
C3791 C1_P_btm.n0 VSS 2.49999f
C3792 C1_P_btm.n1 VSS 3.88666f
C3793 C1_P_btm.t0 VSS 0.280658f
C3794 C1_P_btm.n2 VSS 4.86011f
C3795 C1_P_btm.t3 VSS 1.42799f
C3796 C1_P_btm.t4 VSS 1.35139f
C3797 C1_P_btm.n3 VSS 0.777183f
C3798 C1_P_btm.t2 VSS 1.35139f
C3799 C1_P_btm.n4 VSS 0.953534f
C3800 a_n2661_45956.n1 VSS 0.304656f
C3801 a_n2661_45956.n3 VSS 5.2003f
C3802 C0_dummy_P_btm.t1 VSS 0.577719f
C3803 C0_dummy_P_btm.t0 VSS 0.306925f
C3804 C0_dummy_P_btm.n0 VSS 6.05197f
C3805 C0_dummy_P_btm.t3 VSS 1.34954f
C3806 C0_dummy_P_btm.t2 VSS 1.27716f
C3807 C0_dummy_P_btm.n1 VSS 1.14f
C3808 a_n331_42718.n0 VSS 0.347058f
C3809 a_n331_42718.n1 VSS 2.40082f
C3810 a_n1551_44324.n0 VSS 0.737729f
C3811 a_n1551_44324.n2 VSS 0.525416f
C3812 a_n1551_44324.n3 VSS 8.14518f
C3813 a_n1551_44324.n8 VSS 0.192233f
C3814 a_n1551_44324.n9 VSS 0.139712f
C3815 a_n2442_43262.n0 VSS 0.131505f
C3816 a_n2442_43262.t4 VSS 2.72527f
C3817 a_n2442_43262.n1 VSS 18.4681f
C3818 a_n2442_43262.n2 VSS 0.158219f
C3819 C5_N_btm.t36 VSS 0.800169f
C3820 C5_N_btm.t37 VSS 0.248689f
C3821 C5_N_btm.t1 VSS 0.166821f
C3822 C5_N_btm.n0 VSS 1.26557f
C3823 C5_N_btm.n1 VSS 1.978f
C3824 C5_N_btm.t0 VSS 0.107115f
C3825 C5_N_btm.n2 VSS 2.61124f
C3826 C5_N_btm.t15 VSS 0.716738f
C3827 C5_N_btm.n3 VSS 0.218419f
C3828 C5_N_btm.t35 VSS 0.745082f
C3829 C5_N_btm.t9 VSS 0.717943f
C3830 C5_N_btm.n12 VSS 0.358179f
C3831 C5_N_btm.t4 VSS 0.717943f
C3832 C5_N_btm.n13 VSS 0.248633f
C3833 C5_N_btm.t8 VSS 0.717943f
C3834 C5_N_btm.n14 VSS 0.248633f
C3835 C5_N_btm.t18 VSS 0.717943f
C3836 C5_N_btm.n15 VSS 0.248633f
C3837 C5_N_btm.n18 VSS 0.131769f
C3838 C5_N_btm.n19 VSS 0.1256f
C3839 C5_N_btm.n20 VSS 0.1256f
C3840 C5_N_btm.t11 VSS 0.716738f
C3841 C5_N_btm.n23 VSS 0.218419f
C3842 C5_N_btm.t17 VSS 0.646259f
C3843 C5_N_btm.n25 VSS 0.120948f
C3844 C5_N_btm.t12 VSS 0.646259f
C3845 C5_N_btm.n28 VSS 0.120948f
C3846 C5_N_btm.t6 VSS 0.716738f
C3847 C5_N_btm.n30 VSS 0.218419f
C3848 C5_N_btm.n31 VSS 0.131769f
C3849 C5_N_btm.t30 VSS 0.646259f
C3850 C5_N_btm.n35 VSS 0.120948f
C3851 C5_N_btm.t2 VSS 0.646259f
C3852 C5_N_btm.n38 VSS 0.120948f
C3853 C5_N_btm.t27 VSS 0.646259f
C3854 C5_N_btm.n41 VSS 0.120948f
C3855 C5_N_btm.t21 VSS 0.646259f
C3856 C5_N_btm.n44 VSS 0.120948f
C3857 C5_N_btm.t26 VSS 0.646259f
C3858 C5_N_btm.n47 VSS 0.120948f
C3859 C5_N_btm.t33 VSS 0.646259f
C3860 C5_N_btm.n50 VSS 0.120948f
C3861 C5_N_btm.t29 VSS 0.646259f
C3862 C5_N_btm.n53 VSS 0.120948f
C3863 C5_N_btm.t19 VSS 0.646259f
C3864 C5_N_btm.n56 VSS 0.120948f
C3865 C5_N_btm.t14 VSS 0.716738f
C3866 C5_N_btm.n58 VSS 0.218419f
C3867 C5_N_btm.n59 VSS 0.167798f
C3868 C5_N_btm.t23 VSS 0.716738f
C3869 C5_N_btm.n60 VSS 0.106646f
C3870 C5_N_btm.t7 VSS 0.646259f
C3871 C5_N_btm.n62 VSS 0.120948f
C3872 C5_N_btm.t25 VSS 0.646259f
C3873 C5_N_btm.n65 VSS 0.120948f
C3874 C5_N_btm.t16 VSS 0.646259f
C3875 C5_N_btm.n68 VSS 0.120948f
C3876 C5_N_btm.t3 VSS 0.646259f
C3877 C5_N_btm.n71 VSS 0.120948f
C3878 C5_N_btm.t32 VSS 0.646259f
C3879 C5_N_btm.n74 VSS 0.120948f
C3880 C5_N_btm.t13 VSS 0.646259f
C3881 C5_N_btm.n77 VSS 0.120948f
C3882 C5_N_btm.t22 VSS 0.646259f
C3883 C5_N_btm.n80 VSS 0.120948f
C3884 C5_N_btm.t28 VSS 0.646259f
C3885 C5_N_btm.n83 VSS 0.120948f
C3886 C5_N_btm.t24 VSS 0.716738f
C3887 C5_N_btm.n85 VSS 0.106646f
C3888 C5_N_btm.n86 VSS 0.167798f
C3889 C5_N_btm.t20 VSS 0.717943f
C3890 C5_N_btm.n87 VSS 0.248633f
C3891 C5_N_btm.t5 VSS 0.717943f
C3892 C5_N_btm.n88 VSS 0.248633f
C3893 C5_N_btm.t31 VSS 0.717943f
C3894 C5_N_btm.n89 VSS 0.248633f
C3895 C5_N_btm.t10 VSS 0.717943f
C3896 C5_N_btm.n90 VSS 0.248633f
C3897 C5_N_btm.t34 VSS 0.717943f
C3898 C5_N_btm.n91 VSS 0.42878f
C3899 a_1429_47222.n4 VSS 0.722854f
C3900 a_1429_47222.n5 VSS 0.454134f
C3901 a_1429_47222.n6 VSS 0.737681f
C3902 a_1429_47222.n7 VSS 0.533327f
C3903 a_1429_47222.n9 VSS 0.647926f
C3904 a_1429_47222.n10 VSS 0.482077f
C3905 a_1429_47222.n11 VSS 2.4563f
C3906 a_1429_47222.n13 VSS 2.81848f
C3907 a_1429_47222.n14 VSS 0.233935f
C3908 a_1429_47222.n16 VSS 0.129052f
C3909 a_n1827_45412.n2 VSS 0.178962f
C3910 a_n1827_45412.n4 VSS 0.110851f
C3911 a_n1827_45412.n5 VSS 0.192129f
C3912 a_n1827_45412.n7 VSS 0.261843f
C3913 a_n1827_45412.n8 VSS 10.9405f
C3914 a_n1827_45412.n9 VSS 0.115092f
C3915 C0_dummy_N_btm.t1 VSS 0.577719f
C3916 C0_dummy_N_btm.t0 VSS 0.306925f
C3917 C0_dummy_N_btm.n0 VSS 6.05197f
C3918 C0_dummy_N_btm.t2 VSS 1.34954f
C3919 C0_dummy_N_btm.t3 VSS 1.27716f
C3920 C0_dummy_N_btm.n1 VSS 1.14f
C3921 a_n2442_44894.n0 VSS 0.151634f
C3922 a_n2442_44894.t6 VSS 0.665356f
C3923 a_n2442_44894.n1 VSS 0.330494f
C3924 a_n2442_44894.t5 VSS 0.665356f
C3925 a_n2442_44894.t7 VSS 0.667041f
C3926 a_n2442_44894.n2 VSS 0.319738f
C3927 a_n2442_44894.t4 VSS 0.684433f
C3928 a_n2442_44894.n3 VSS 0.618085f
C3929 a_n2442_44894.n4 VSS 7.86205f
C3930 a_n2442_44894.n5 VSS 6.70337f
C3931 a_n2661_45420.n0 VSS 0.101218f
C3932 a_n2661_45420.n1 VSS 0.467687f
C3933 a_n2661_45420.n2 VSS 0.116647f
C3934 a_n2661_45420.n3 VSS 2.40249f
C3935 a_n2661_45420.n4 VSS 12.2254f
C3936 a_n2661_45420.n5 VSS 0.256162f
C3937 a_6974_31099.n0 VSS 0.163252f
C3938 a_6974_31099.t5 VSS 0.32074f
C3939 a_6974_31099.t4 VSS 0.304506f
C3940 a_6974_31099.n1 VSS 20.5883f
C3941 a_6974_31099.n2 VSS 11.573f
C3942 a_17738_32299.n0 VSS 0.119963f
C3943 a_17738_32299.t4 VSS 0.7719f
C3944 a_17738_32299.t5 VSS 0.794031f
C3945 a_17738_32299.n1 VSS 4.47819f
C3946 a_17738_32299.n2 VSS 13.1099f
C3947 a_17738_32299.n3 VSS 0.13251f
C3948 a_n690_43494.n5 VSS 0.380534f
C3949 a_n690_43494.n7 VSS 0.235566f
C3950 a_n690_43494.n10 VSS 0.683813f
C3951 a_n690_43494.n13 VSS 0.399617f
C3952 a_n690_43494.n14 VSS 0.605733f
C3953 a_n690_43494.n15 VSS 0.344626f
C3954 a_n690_43494.n16 VSS 0.188742f
C3955 a_n690_43494.n18 VSS 0.557222f
C3956 a_n690_43494.n19 VSS 0.482174f
C3957 a_n690_43494.n20 VSS 0.143238f
C3958 a_5734_30651.n0 VSS 0.176734f
C3959 a_5734_30651.n1 VSS 0.261761f
C3960 a_5734_30651.t5 VSS 0.448749f
C3961 a_5734_30651.t6 VSS 0.416504f
C3962 a_5734_30651.n2 VSS 19.8088f
C3963 a_5734_30651.n3 VSS 12.2269f
C3964 a_5734_30651.n4 VSS 0.540878f
C3965 a_1334_43494.n2 VSS 0.113293f
C3966 a_1334_43494.n4 VSS 0.14913f
C3967 a_1334_43494.n5 VSS 1.16186f
C3968 a_1334_43494.n8 VSS 0.308226f
C3969 a_1334_43494.n14 VSS 0.335874f
C3970 a_1334_43494.n15 VSS 0.133657f
C3971 a_1334_43494.n17 VSS 0.143015f
C3972 a_1334_43494.n20 VSS 0.261348f
C3973 a_1334_43494.n21 VSS 0.318262f
C3974 a_n1890_42718.n0 VSS 0.134362f
C3975 a_n1890_42718.t4 VSS 2.60255f
C3976 a_n1890_42718.n1 VSS 19.398f
C3977 a_n1890_42718.n2 VSS 0.148416f
C3978 a_n1067_42718.n3 VSS 1.60892f
C3979 a_n1067_42718.n4 VSS 2.18924f
C3980 a_13248_45956.n1 VSS 0.104336f
C3981 a_13248_45956.n3 VSS 0.129402f
C3982 a_13248_45956.n4 VSS 0.154871f
C3983 a_13248_45956.n5 VSS 0.121541f
C3984 a_13248_45956.n6 VSS 0.147965f
C3985 a_13248_45956.n7 VSS 0.147737f
C3986 a_13248_45956.n9 VSS 0.992564f
C3987 a_13248_45956.n10 VSS 0.817192f
C3988 a_13248_45956.t12 VSS 0.108653f
C3989 a_13248_45956.n11 VSS 0.503519f
C3990 a_13248_45956.n14 VSS 0.147422f
C3991 a_13248_45956.n15 VSS 0.938815f
C3992 a_13248_45956.n16 VSS 0.59511f
C3993 a_13248_45956.n18 VSS 0.115731f
C3994 a_13248_45956.n19 VSS 0.506844f
C3995 a_13248_45956.n20 VSS 1.30958f
C3996 a_13248_45956.n21 VSS 0.678824f
C3997 a_13248_45956.n22 VSS 0.100437f
C3998 a_n2109_47596.n2 VSS 0.160501f
C3999 a_n2109_47596.n3 VSS 1.27695f
C4000 a_n2109_47596.n4 VSS 5.48402f
C4001 a_n2109_47596.n5 VSS 0.108264f
C4002 C3_N_btm.t1 VSS 0.973133f
C4003 C3_N_btm.t12 VSS 0.297776f
C4004 C3_N_btm.t11 VSS 0.199749f
C4005 C3_N_btm.n0 VSS 1.55495f
C4006 C3_N_btm.n1 VSS 2.46584f
C4007 C3_N_btm.t0 VSS 0.151676f
C4008 C3_N_btm.n2 VSS 2.91541f
C4009 C3_N_btm.t5 VSS 0.881786f
C4010 C3_N_btm.t8 VSS 0.856786f
C4011 C3_N_btm.n3 VSS 0.286809f
C4012 C3_N_btm.t7 VSS 0.856786f
C4013 C3_N_btm.n4 VSS 0.1698f
C4014 C3_N_btm.t9 VSS 0.856786f
C4015 C3_N_btm.n5 VSS 0.1698f
C4016 C3_N_btm.t6 VSS 0.856786f
C4017 C3_N_btm.n6 VSS 0.167366f
C4018 C3_N_btm.t3 VSS 0.858208f
C4019 C3_N_btm.n7 VSS 0.26968f
C4020 C3_N_btm.t4 VSS 0.859652f
C4021 C3_N_btm.n8 VSS 0.305094f
C4022 C3_N_btm.t2 VSS 0.859652f
C4023 C3_N_btm.n9 VSS 0.297708f
C4024 C3_N_btm.t10 VSS 0.859652f
C4025 C3_N_btm.n10 VSS 0.625101f
C4026 a_20163_31459.n0 VSS 0.115994f
C4027 a_20163_31459.t4 VSS 2.97226f
C4028 a_20163_31459.n1 VSS 15.180901f
C4029 a_20163_31459.n2 VSS 0.139556f
C4030 a_17930_32299.n0 VSS 0.150407f
C4031 a_17930_32299.t6 VSS 0.659973f
C4032 a_17930_32299.n1 VSS 0.32782f
C4033 a_17930_32299.t7 VSS 0.659973f
C4034 a_17930_32299.t4 VSS 0.678895f
C4035 a_17930_32299.t5 VSS 0.661643f
C4036 a_17930_32299.n2 VSS 0.317151f
C4037 a_17930_32299.n3 VSS 0.613084f
C4038 a_17930_32299.n4 VSS 7.70741f
C4039 a_17930_32299.n5 VSS 7.09307f
C4040 a_927_42692.n2 VSS 0.141353f
C4041 a_927_42692.n3 VSS 0.248719f
C4042 a_927_42692.n6 VSS 0.179207f
C4043 a_927_42692.n11 VSS 0.341072f
C4044 a_927_42692.n12 VSS 0.20517f
C4045 a_927_42692.n15 VSS 0.313237f
C4046 a_927_42692.n17 VSS 0.268358f
C4047 a_927_42692.n18 VSS 0.666784f
C4048 a_927_42692.n19 VSS 3.73743f
C4049 a_927_42692.n22 VSS 0.137671f
C4050 a_n237_45454.n6 VSS 0.196257f
C4051 a_n237_45454.n7 VSS 0.461232f
C4052 a_n237_45454.n8 VSS 0.343416f
C4053 a_n237_45454.n10 VSS 0.746842f
C4054 a_n237_45454.n12 VSS 0.194552f
C4055 a_n237_45454.n14 VSS 0.346494f
C4056 a_n237_45454.n15 VSS 0.181208f
C4057 a_n237_45454.n17 VSS 0.439651f
C4058 a_n237_45454.n19 VSS 0.334063f
C4059 a_n237_45454.n20 VSS 0.190893f
C4060 a_12769_44594.n4 VSS 0.99504f
C4061 a_12769_44594.n5 VSS 0.579981f
C4062 a_12769_44594.n6 VSS 0.887905f
C4063 a_12769_44594.n7 VSS 0.257805f
C4064 a_13144_47452.n1 VSS 1.56368f
C4065 a_13144_47452.n2 VSS 0.550354f
C4066 a_5142_30651.n0 VSS 0.15291f
C4067 a_5142_30651.t9 VSS 0.670955f
C4068 a_5142_30651.t5 VSS 0.69096f
C4069 a_5142_30651.n1 VSS 0.880057f
C4070 a_5142_30651.t6 VSS 0.670955f
C4071 a_5142_30651.t4 VSS 0.69096f
C4072 a_5142_30651.n2 VSS 0.91668f
C4073 a_5142_30651.n3 VSS 11.391201f
C4074 a_5142_30651.n4 VSS 0.190644f
C4075 a_5142_30651.n5 VSS 5.77119f
C4076 a_5142_30651.n6 VSS 0.410339f
C4077 a_n1827_44868.n0 VSS 0.754372f
C4078 a_n1827_44868.n2 VSS 0.364566f
C4079 a_n1827_44868.n3 VSS 6.65089f
C4080 a_n1827_44868.n8 VSS 0.176972f
C4081 a_n1741_47596.n2 VSS 0.234377f
C4082 a_n1741_47596.n3 VSS 0.441704f
C4083 a_n1741_47596.n4 VSS 15.5836f
C4084 a_n1741_47596.n5 VSS 0.163879f
C4085 a_8727_47222.n3 VSS 0.35005f
C4086 a_8727_47222.n6 VSS 0.214407f
C4087 a_8727_47222.n7 VSS 0.338557f
C4088 a_8727_47222.n11 VSS 0.170752f
C4089 a_8727_47222.n13 VSS 0.52113f
C4090 a_8727_47222.n15 VSS 1.03517f
C4091 a_8727_47222.n18 VSS 1.02782f
C4092 a_8727_47222.n19 VSS 0.520454f
C4093 a_8727_47222.n20 VSS 0.111269f
C4094 a_1343_38525.n2 VSS 0.120195f
C4095 a_1343_38525.n3 VSS 0.545196f
C4096 a_1343_38525.n4 VSS 0.243609f
C4097 a_1343_38525.n5 VSS 0.658075f
C4098 a_1343_38525.n6 VSS 0.300753f
C4099 a_1343_38525.n7 VSS 0.261686f
C4100 a_1343_38525.n8 VSS 0.321183f
C4101 a_1343_38525.n9 VSS 0.121769f
C4102 SMPL_ON_N.n2 VSS 0.27022f
C4103 SMPL_ON_N.n3 VSS 0.105922f
C4104 SMPL_ON_N.n5 VSS 0.367767f
C4105 SMPL_ON_N.n6 VSS 3.62083f
C4106 SMPL_ON_N.n7 VSS 0.183946f
C4107 a_n2810_47070.t6 VSS 1.29695f
C4108 a_n2810_47070.t4 VSS 1.29675f
C4109 a_n2810_47070.n1 VSS 0.960609f
C4110 a_n2810_47070.t7 VSS 1.29675f
C4111 a_n2810_47070.n2 VSS 0.486539f
C4112 a_n2810_47070.t5 VSS 1.29675f
C4113 a_n2810_47070.n3 VSS 6.19402f
C4114 a_n2810_47070.n4 VSS 4.47635f
C4115 a_10227_47214.n5 VSS 0.106688f
C4116 a_10227_47214.n8 VSS 0.153814f
C4117 a_10227_47214.n12 VSS 0.148081f
C4118 a_10227_47214.n13 VSS 0.114575f
C4119 a_10227_47214.n16 VSS 0.117815f
C4120 a_10227_47214.n17 VSS 0.102965f
C4121 a_10227_47214.n20 VSS 0.126569f
C4122 a_10227_47214.n26 VSS 0.190543f
C4123 a_10227_47214.n29 VSS 0.108219f
C4124 a_10227_47214.n30 VSS 0.12477f
C4125 a_10227_47214.n33 VSS 0.107478f
C4126 a_10227_47214.n34 VSS 0.540932f
C4127 a_10227_47214.n37 VSS 0.137574f
C4128 a_10227_47214.n38 VSS 0.307666f
C4129 a_n2467_30659.t6 VSS 0.836236f
C4130 a_n2467_30659.t5 VSS 0.836106f
C4131 a_n2467_30659.n1 VSS 0.620289f
C4132 a_n2467_30659.t10 VSS 0.836106f
C4133 a_n2467_30659.n2 VSS 0.314326f
C4134 a_n2467_30659.t11 VSS 0.836106f
C4135 a_n2467_30659.n3 VSS 0.314326f
C4136 a_n2467_30659.t8 VSS 0.836106f
C4137 a_n2467_30659.n4 VSS 0.314326f
C4138 a_n2467_30659.t9 VSS 0.836106f
C4139 a_n2467_30659.n5 VSS 0.314326f
C4140 a_n2467_30659.t4 VSS 0.836106f
C4141 a_n2467_30659.n6 VSS 0.313281f
C4142 a_n2467_30659.t7 VSS 0.836108f
C4143 a_n2467_30659.n7 VSS 3.98617f
C4144 a_n2467_30659.n8 VSS 2.94358f
C4145 COMP_P.n1 VSS 0.132565f
C4146 COMP_P.n2 VSS 0.462534f
C4147 COMP_P.n5 VSS 0.340041f
C4148 COMP_P.n6 VSS 0.174925f
C4149 COMP_P.n7 VSS 2.29879f
C4150 COMP_P.n8 VSS 0.378195f
C4151 COMP_P.n9 VSS 13.4253f
C4152 C2_N_btm.t8 VSS 1.43552f
C4153 C2_N_btm.t7 VSS 0.436024f
C4154 C2_N_btm.t0 VSS 0.292486f
C4155 C2_N_btm.n0 VSS 2.30503f
C4156 C2_N_btm.n1 VSS 3.53635f
C4157 C2_N_btm.t1 VSS 0.199791f
C4158 C2_N_btm.n2 VSS 4.30601f
C4159 C2_N_btm.t5 VSS 1.29119f
C4160 C2_N_btm.t4 VSS 1.25457f
C4161 C2_N_btm.n3 VSS 0.416387f
C4162 C2_N_btm.t2 VSS 1.25665f
C4163 C2_N_btm.n4 VSS 0.394884f
C4164 C2_N_btm.t3 VSS 1.25876f
C4165 C2_N_btm.n5 VSS 0.44674f
C4166 C2_N_btm.t6 VSS 1.25876f
C4167 C2_N_btm.n6 VSS 0.809132f
C4168 VCM.t48 VSS 0.193436f
C4169 VCM.t2 VSS 0.193436f
C4170 VCM.n0 VSS 0.802861f
C4171 VCM.t22 VSS 0.184424f
C4172 VCM.t44 VSS 0.181802f
C4173 VCM.n1 VSS 0.604443f
C4174 VCM.t54 VSS 0.181802f
C4175 VCM.n2 VSS 0.320018f
C4176 VCM.t20 VSS 0.181802f
C4177 VCM.n3 VSS 0.320018f
C4178 VCM.t47 VSS 0.181802f
C4179 VCM.n4 VSS 0.320018f
C4180 VCM.t27 VSS 0.181802f
C4181 VCM.n5 VSS 0.320018f
C4182 VCM.n6 VSS 0.131979f
C4183 VCM.n7 VSS 0.28045f
C4184 VCM.t50 VSS 0.181802f
C4185 VCM.n8 VSS 0.774244f
C4186 VCM.t0 VSS 0.193436f
C4187 VCM.t57 VSS 0.193436f
C4188 VCM.n9 VSS 0.783937f
C4189 VCM.n10 VSS 1.60249f
C4190 VCM.t56 VSS 0.193436f
C4191 VCM.t63 VSS 0.193436f
C4192 VCM.n11 VSS 0.783937f
C4193 VCM.n12 VSS 0.609248f
C4194 VCM.t62 VSS 0.193436f
C4195 VCM.t19 VSS 0.193436f
C4196 VCM.n13 VSS 0.783937f
C4197 VCM.n14 VSS 0.610914f
C4198 VCM.t12 VSS 0.193436f
C4199 VCM.t16 VSS 0.193436f
C4200 VCM.n15 VSS 0.783937f
C4201 VCM.n16 VSS 0.610914f
C4202 VCM.t10 VSS 0.193436f
C4203 VCM.t7 VSS 0.193436f
C4204 VCM.n17 VSS 0.783937f
C4205 VCM.n18 VSS 0.609449f
C4206 VCM.t14 VSS 0.193436f
C4207 VCM.t9 VSS 0.193436f
C4208 VCM.n19 VSS 0.783937f
C4209 VCM.n20 VSS 0.609449f
C4210 VCM.t18 VSS 0.193436f
C4211 VCM.t43 VSS 0.193436f
C4212 VCM.n21 VSS 0.783937f
C4213 VCM.n22 VSS 0.610914f
C4214 VCM.t38 VSS 0.193436f
C4215 VCM.t42 VSS 0.193436f
C4216 VCM.n23 VSS 0.783937f
C4217 VCM.n24 VSS 0.610914f
C4218 VCM.t40 VSS 0.193436f
C4219 VCM.t41 VSS 0.193436f
C4220 VCM.n25 VSS 0.783937f
C4221 VCM.n26 VSS 0.609449f
C4222 VCM.t36 VSS 0.193436f
C4223 VCM.t39 VSS 0.193436f
C4224 VCM.n27 VSS 0.783937f
C4225 VCM.n28 VSS 0.609449f
C4226 VCM.t37 VSS 0.991655f
C4227 VCM.n29 VSS 2.66959f
C4228 VCM.t23 VSS 0.184424f
C4229 VCM.t45 VSS 0.181802f
C4230 VCM.n30 VSS 0.604443f
C4231 VCM.t55 VSS 0.181802f
C4232 VCM.n31 VSS 0.320018f
C4233 VCM.t21 VSS 0.181802f
C4234 VCM.n32 VSS 0.320018f
C4235 VCM.t46 VSS 0.181802f
C4236 VCM.n33 VSS 0.320018f
C4237 VCM.t26 VSS 0.181802f
C4238 VCM.n34 VSS 0.320018f
C4239 VCM.n35 VSS 0.131979f
C4240 VCM.n36 VSS 0.28045f
C4241 VCM.t52 VSS 0.181802f
C4242 VCM.n37 VSS 0.774244f
C4243 VCM.t3 VSS 0.193436f
C4244 VCM.t49 VSS 0.193436f
C4245 VCM.n38 VSS 0.802861f
C4246 VCM.t61 VSS 0.193436f
C4247 VCM.t1 VSS 0.193436f
C4248 VCM.n39 VSS 0.783937f
C4249 VCM.n40 VSS 1.60249f
C4250 VCM.t59 VSS 0.193436f
C4251 VCM.t58 VSS 0.193436f
C4252 VCM.n41 VSS 0.783937f
C4253 VCM.n42 VSS 0.609248f
C4254 VCM.t4 VSS 0.193436f
C4255 VCM.t60 VSS 0.193436f
C4256 VCM.n43 VSS 0.783937f
C4257 VCM.n44 VSS 0.610914f
C4258 VCM.t11 VSS 0.193436f
C4259 VCM.t5 VSS 0.193436f
C4260 VCM.n45 VSS 0.783937f
C4261 VCM.n46 VSS 0.610914f
C4262 VCM.t15 VSS 0.193436f
C4263 VCM.t17 VSS 0.193436f
C4264 VCM.n47 VSS 0.783937f
C4265 VCM.n48 VSS 0.609449f
C4266 VCM.t6 VSS 0.193436f
C4267 VCM.t13 VSS 0.193436f
C4268 VCM.n49 VSS 0.783937f
C4269 VCM.n50 VSS 0.609449f
C4270 VCM.t30 VSS 0.193436f
C4271 VCM.t8 VSS 0.193436f
C4272 VCM.n51 VSS 0.783937f
C4273 VCM.n52 VSS 0.610914f
C4274 VCM.t31 VSS 0.193436f
C4275 VCM.t28 VSS 0.193436f
C4276 VCM.n53 VSS 0.783937f
C4277 VCM.n54 VSS 0.610914f
C4278 VCM.t33 VSS 0.193436f
C4279 VCM.t29 VSS 0.193436f
C4280 VCM.n55 VSS 0.783937f
C4281 VCM.n56 VSS 0.609449f
C4282 VCM.t35 VSS 0.193436f
C4283 VCM.t34 VSS 0.193436f
C4284 VCM.n57 VSS 0.783937f
C4285 VCM.n58 VSS 0.609449f
C4286 VCM.t32 VSS 0.991655f
C4287 VCM.n59 VSS 9.33799f
C4288 VCM.n60 VSS 21.565f
C4289 a_3222_30651.n1 VSS 0.103491f
C4290 a_3222_30651.t7 VSS 0.269835f
C4291 a_3222_30651.t11 VSS 0.27788f
C4292 a_3222_30651.t19 VSS 0.27029f
C4293 a_3222_30651.t21 VSS 0.269835f
C4294 a_3222_30651.t5 VSS 0.27029f
C4295 a_3222_30651.t4 VSS 0.269835f
C4296 a_3222_30651.t13 VSS 0.27029f
C4297 a_3222_30651.n2 VSS 0.124034f
C4298 a_3222_30651.t12 VSS 0.269835f
C4299 a_3222_30651.n3 VSS 0.133387f
C4300 a_3222_30651.n4 VSS 0.181739f
C4301 a_3222_30651.n5 VSS 0.138752f
C4302 a_3222_30651.n6 VSS 0.124034f
C4303 a_3222_30651.n7 VSS 0.138752f
C4304 a_3222_30651.n8 VSS 0.124034f
C4305 a_3222_30651.n9 VSS 0.245096f
C4306 a_3222_30651.n10 VSS 0.959896f
C4307 a_3222_30651.n11 VSS 0.103491f
C4308 a_3222_30651.t20 VSS 0.269835f
C4309 a_3222_30651.t17 VSS 0.27029f
C4310 a_3222_30651.t15 VSS 0.269835f
C4311 a_3222_30651.t9 VSS 0.27029f
C4312 a_3222_30651.t10 VSS 0.269835f
C4313 a_3222_30651.t6 VSS 0.27029f
C4314 a_3222_30651.n12 VSS 0.124034f
C4315 a_3222_30651.t8 VSS 0.269835f
C4316 a_3222_30651.n13 VSS 0.133387f
C4317 a_3222_30651.n14 VSS 0.181739f
C4318 a_3222_30651.n15 VSS 0.138752f
C4319 a_3222_30651.n16 VSS 0.124034f
C4320 a_3222_30651.n17 VSS 0.138752f
C4321 a_3222_30651.n18 VSS 0.124034f
C4322 a_3222_30651.t16 VSS 0.27788f
C4323 a_3222_30651.n19 VSS 0.245096f
C4324 a_3222_30651.n20 VSS 1.07208f
C4325 a_3222_30651.n21 VSS 4.381741f
C4326 a_3222_30651.n23 VSS 3.05082f
C4327 a_3222_30651.n24 VSS 0.172287f
C4328 a_n1735_43236.n2 VSS 0.176989f
C4329 a_n1735_43236.n5 VSS 1.29891f
C4330 a_n1735_43236.n7 VSS 0.160601f
C4331 a_n1735_43236.n8 VSS 5.20978f
C4332 a_n1551_45412.n2 VSS 0.314529f
C4333 a_n1551_45412.n3 VSS 1.02212f
C4334 a_n1551_45412.n4 VSS 0.100678f
C4335 a_n1551_45412.n5 VSS 1.78137f
C4336 a_n1551_45412.n6 VSS 14.6307f
C4337 a_n1551_45412.n9 VSS 0.357721f
C4338 a_n1551_45412.n10 VSS 0.11205f
C4339 a_20892_30659.t4 VSS 3.10232f
C4340 a_20892_30659.n0 VSS 0.173492f
C4341 a_20892_30659.n1 VSS 15.058199f
C4342 C7_P_btm.n0 VSS 0.507967f
C4343 C7_P_btm.t137 VSS 0.60976f
C4344 C7_P_btm.n1 VSS 1.13336f
C4345 C7_P_btm.t138 VSS 0.613007f
C4346 C7_P_btm.n2 VSS 0.606693f
C4347 C7_P_btm.t0 VSS 0.115562f
C4348 C7_P_btm.n3 VSS 1.49629f
C4349 C7_P_btm.t7 VSS 0.401902f
C4350 C7_P_btm.n5 VSS 0.12684f
C4351 C7_P_btm.t15 VSS 0.386613f
C4352 C7_P_btm.t39 VSS 0.386613f
C4353 C7_P_btm.t75 VSS 0.397234f
C4354 C7_P_btm.t47 VSS 0.385972f
C4355 C7_P_btm.n15 VSS 0.129204f
C4356 C7_P_btm.t81 VSS 0.385972f
C4357 C7_P_btm.t62 VSS 0.385972f
C4358 C7_P_btm.t95 VSS 0.385972f
C4359 C7_P_btm.t61 VSS 0.385972f
C4360 C7_P_btm.t63 VSS 0.386613f
C4361 C7_P_btm.t77 VSS 0.386613f
C4362 C7_P_btm.n21 VSS 0.117817f
C4363 C7_P_btm.t121 VSS 0.386613f
C4364 C7_P_btm.t100 VSS 0.386613f
C4365 C7_P_btm.t3 VSS 0.401902f
C4366 C7_P_btm.n34 VSS 0.12684f
C4367 C7_P_btm.t4 VSS 0.401902f
C4368 C7_P_btm.t8 VSS 0.401902f
C4369 C7_P_btm.n35 VSS 0.146274f
C4370 C7_P_btm.t36 VSS 0.386613f
C4371 C7_P_btm.t124 VSS 0.348597f
C4372 C7_P_btm.t27 VSS 0.386613f
C4373 C7_P_btm.n41 VSS 0.146274f
C4374 C7_P_btm.t130 VSS 0.386613f
C4375 C7_P_btm.t66 VSS 0.386613f
C4376 C7_P_btm.t94 VSS 0.348597f
C4377 C7_P_btm.t68 VSS 0.386613f
C4378 C7_P_btm.t82 VSS 0.348597f
C4379 C7_P_btm.t126 VSS 0.386613f
C4380 C7_P_btm.t26 VSS 0.348597f
C4381 C7_P_btm.t90 VSS 0.386613f
C4382 C7_P_btm.t78 VSS 0.386613f
C4383 C7_P_btm.t87 VSS 0.386613f
C4384 C7_P_btm.t122 VSS 0.348597f
C4385 C7_P_btm.t67 VSS 0.386613f
C4386 C7_P_btm.t105 VSS 0.348597f
C4387 C7_P_btm.t76 VSS 0.386613f
C4388 C7_P_btm.t31 VSS 0.348597f
C4389 C7_P_btm.t113 VSS 0.386613f
C4390 C7_P_btm.t101 VSS 0.386613f
C4391 C7_P_btm.t111 VSS 0.386613f
C4392 C7_P_btm.t19 VSS 0.348597f
C4393 C7_P_btm.t98 VSS 0.386613f
C4394 C7_P_btm.t118 VSS 0.348597f
C4395 C7_P_btm.t35 VSS 0.386613f
C4396 C7_P_btm.t99 VSS 0.397234f
C4397 C7_P_btm.t65 VSS 0.385972f
C4398 C7_P_btm.n99 VSS 0.129204f
C4399 C7_P_btm.t37 VSS 0.385972f
C4400 C7_P_btm.t129 VSS 0.385972f
C4401 C7_P_btm.t30 VSS 0.385972f
C4402 C7_P_btm.t107 VSS 0.385972f
C4403 C7_P_btm.t52 VSS 0.348597f
C4404 C7_P_btm.t131 VSS 0.348597f
C4405 C7_P_btm.t13 VSS 0.386613f
C4406 C7_P_btm.t48 VSS 0.386613f
C4407 C7_P_btm.t45 VSS 0.386613f
C4408 C7_P_btm.n142 VSS 0.117817f
C4409 C7_P_btm.t18 VSS 0.348597f
C4410 C7_P_btm.t51 VSS 0.348597f
C4411 C7_P_btm.t49 VSS 0.348597f
C4412 C7_P_btm.t136 VSS 0.348597f
C4413 C7_P_btm.t28 VSS 0.348597f
C4414 C7_P_btm.t22 VSS 0.348597f
C4415 C7_P_btm.t123 VSS 0.348597f
C4416 C7_P_btm.t11 VSS 0.348597f
C4417 C7_P_btm.t96 VSS 0.348597f
C4418 C7_P_btm.t20 VSS 0.348597f
C4419 C7_P_btm.t104 VSS 0.348597f
C4420 C7_P_btm.t119 VSS 0.348597f
C4421 C7_P_btm.t46 VSS 0.348597f
C4422 C7_P_btm.t79 VSS 0.348597f
C4423 C7_P_btm.t56 VSS 0.386613f
C4424 C7_P_btm.n185 VSS 0.117817f
C4425 C7_P_btm.t108 VSS 0.348597f
C4426 C7_P_btm.t14 VSS 0.348597f
C4427 C7_P_btm.t92 VSS 0.348597f
C4428 C7_P_btm.t53 VSS 0.348597f
C4429 C7_P_btm.t40 VSS 0.348597f
C4430 C7_P_btm.t44 VSS 0.348597f
C4431 C7_P_btm.t32 VSS 0.348597f
C4432 C7_P_btm.t110 VSS 0.348597f
C4433 C7_P_btm.t17 VSS 0.348597f
C4434 C7_P_btm.t132 VSS 0.348597f
C4435 C7_P_btm.t120 VSS 0.348597f
C4436 C7_P_btm.t42 VSS 0.348597f
C4437 C7_P_btm.t59 VSS 0.348597f
C4438 C7_P_btm.t34 VSS 0.348597f
C4439 C7_P_btm.t117 VSS 0.348597f
C4440 C7_P_btm.t24 VSS 0.348597f
C4441 C7_P_btm.t133 VSS 0.348597f
C4442 C7_P_btm.t73 VSS 0.348597f
C4443 C7_P_btm.n242 VSS 0.117817f
C4444 C7_P_btm.t9 VSS 0.386613f
C4445 C7_P_btm.t41 VSS 0.348597f
C4446 C7_P_btm.t70 VSS 0.348597f
C4447 C7_P_btm.t93 VSS 0.385972f
C4448 C7_P_btm.t16 VSS 0.385972f
C4449 C7_P_btm.t109 VSS 0.385972f
C4450 C7_P_btm.t57 VSS 0.385972f
C4451 C7_P_btm.t116 VSS 0.385972f
C4452 C7_P_btm.t85 VSS 0.385972f
C4453 C7_P_btm.t21 VSS 0.385972f
C4454 C7_P_btm.t91 VSS 0.385972f
C4455 C7_P_btm.t64 VSS 0.385972f
C4456 C7_P_btm.t106 VSS 0.385972f
C4457 C7_P_btm.t72 VSS 0.385972f
C4458 C7_P_btm.t114 VSS 0.385972f
C4459 C7_P_btm.t83 VSS 0.385972f
C4460 C7_P_btm.t80 VSS 0.385972f
C4461 C7_P_btm.t88 VSS 0.348597f
C4462 C7_P_btm.t135 VSS 0.348597f
C4463 C7_P_btm.t127 VSS 0.386613f
C4464 C7_P_btm.t74 VSS 0.348597f
C4465 C7_P_btm.t102 VSS 0.348597f
C4466 C7_P_btm.t115 VSS 0.386613f
C4467 C7_P_btm.t128 VSS 0.386613f
C4468 C7_P_btm.t84 VSS 0.348597f
C4469 C7_P_btm.t71 VSS 0.386613f
C4470 C7_P_btm.t55 VSS 0.348597f
C4471 C7_P_btm.t69 VSS 0.386613f
C4472 C7_P_btm.t58 VSS 0.348597f
C4473 C7_P_btm.t38 VSS 0.386613f
C4474 C7_P_btm.t50 VSS 0.386613f
C4475 C7_P_btm.t112 VSS 0.386613f
C4476 C7_P_btm.t25 VSS 0.348597f
C4477 C7_P_btm.t97 VSS 0.386613f
C4478 C7_P_btm.t33 VSS 0.348597f
C4479 C7_P_btm.t10 VSS 0.386613f
C4480 C7_P_btm.t125 VSS 0.348597f
C4481 C7_P_btm.t134 VSS 0.386613f
C4482 C7_P_btm.t29 VSS 0.386613f
C4483 C7_P_btm.t89 VSS 0.386613f
C4484 C7_P_btm.t54 VSS 0.348597f
C4485 C7_P_btm.t43 VSS 0.386613f
C4486 C7_P_btm.t12 VSS 0.348597f
C4487 C7_P_btm.t103 VSS 0.386613f
C4488 C7_P_btm.t5 VSS 0.401902f
C4489 C7_P_btm.n337 VSS 0.146274f
C4490 C7_P_btm.t60 VSS 0.386613f
C4491 C7_P_btm.t86 VSS 0.348597f
C4492 C7_P_btm.t23 VSS 0.386613f
C4493 C7_P_btm.t6 VSS 0.387263f
C4494 C7_P_btm.n344 VSS 0.2137f
C4495 C7_N_btm.n0 VSS 0.507968f
C4496 C7_N_btm.t137 VSS 0.60976f
C4497 C7_N_btm.n1 VSS 1.13336f
C4498 C7_N_btm.t138 VSS 0.613007f
C4499 C7_N_btm.n2 VSS 0.606693f
C4500 C7_N_btm.t2 VSS 0.115562f
C4501 C7_N_btm.n3 VSS 1.49414f
C4502 C7_N_btm.t135 VSS 0.401902f
C4503 C7_N_btm.n5 VSS 0.12684f
C4504 C7_N_btm.t85 VSS 0.386613f
C4505 C7_N_btm.t134 VSS 0.401902f
C4506 C7_N_btm.t23 VSS 0.386613f
C4507 C7_N_btm.t42 VSS 0.386613f
C4508 C7_N_btm.t61 VSS 0.397234f
C4509 C7_N_btm.t43 VSS 0.385972f
C4510 C7_N_btm.n15 VSS 0.129204f
C4511 C7_N_btm.t33 VSS 0.385972f
C4512 C7_N_btm.t52 VSS 0.385972f
C4513 C7_N_btm.t18 VSS 0.385972f
C4514 C7_N_btm.t107 VSS 0.385972f
C4515 C7_N_btm.t97 VSS 0.386613f
C4516 C7_N_btm.t67 VSS 0.386613f
C4517 C7_N_btm.n21 VSS 0.117817f
C4518 C7_N_btm.t84 VSS 0.386613f
C4519 C7_N_btm.t101 VSS 0.386613f
C4520 C7_N_btm.t136 VSS 0.401902f
C4521 C7_N_btm.n34 VSS 0.12684f
C4522 C7_N_btm.t132 VSS 0.401902f
C4523 C7_N_btm.t122 VSS 0.386613f
C4524 C7_N_btm.t131 VSS 0.401902f
C4525 C7_N_btm.n35 VSS 0.146274f
C4526 C7_N_btm.t78 VSS 0.348597f
C4527 C7_N_btm.t49 VSS 0.386613f
C4528 C7_N_btm.n41 VSS 0.146274f
C4529 C7_N_btm.t98 VSS 0.386613f
C4530 C7_N_btm.t4 VSS 0.386613f
C4531 C7_N_btm.t36 VSS 0.348597f
C4532 C7_N_btm.t114 VSS 0.386613f
C4533 C7_N_btm.t56 VSS 0.348597f
C4534 C7_N_btm.t19 VSS 0.386613f
C4535 C7_N_btm.t120 VSS 0.348597f
C4536 C7_N_btm.t95 VSS 0.386613f
C4537 C7_N_btm.t103 VSS 0.386613f
C4538 C7_N_btm.t41 VSS 0.386613f
C4539 C7_N_btm.t14 VSS 0.348597f
C4540 C7_N_btm.t3 VSS 0.386613f
C4541 C7_N_btm.t26 VSS 0.348597f
C4542 C7_N_btm.t127 VSS 0.386613f
C4543 C7_N_btm.t106 VSS 0.348597f
C4544 C7_N_btm.t74 VSS 0.386613f
C4545 C7_N_btm.t87 VSS 0.386613f
C4546 C7_N_btm.t93 VSS 0.386613f
C4547 C7_N_btm.t8 VSS 0.348597f
C4548 C7_N_btm.t50 VSS 0.386613f
C4549 C7_N_btm.t79 VSS 0.348597f
C4550 C7_N_btm.t124 VSS 0.386613f
C4551 C7_N_btm.t22 VSS 0.397234f
C4552 C7_N_btm.t118 VSS 0.385972f
C4553 C7_N_btm.n99 VSS 0.129204f
C4554 C7_N_btm.t75 VSS 0.385972f
C4555 C7_N_btm.t123 VSS 0.385972f
C4556 C7_N_btm.t69 VSS 0.385972f
C4557 C7_N_btm.t28 VSS 0.385972f
C4558 C7_N_btm.t130 VSS 0.348597f
C4559 C7_N_btm.t90 VSS 0.348597f
C4560 C7_N_btm.t58 VSS 0.386613f
C4561 C7_N_btm.t125 VSS 0.386613f
C4562 C7_N_btm.n142 VSS 0.117817f
C4563 C7_N_btm.t7 VSS 0.348597f
C4564 C7_N_btm.t82 VSS 0.348597f
C4565 C7_N_btm.t21 VSS 0.348597f
C4566 C7_N_btm.t128 VSS 0.348597f
C4567 C7_N_btm.t27 VSS 0.348597f
C4568 C7_N_btm.t76 VSS 0.348597f
C4569 C7_N_btm.t45 VSS 0.348597f
C4570 C7_N_btm.t65 VSS 0.348597f
C4571 C7_N_btm.t102 VSS 0.348597f
C4572 C7_N_btm.t20 VSS 0.348597f
C4573 C7_N_btm.t109 VSS 0.348597f
C4574 C7_N_btm.t113 VSS 0.348597f
C4575 C7_N_btm.t59 VSS 0.348597f
C4576 C7_N_btm.t91 VSS 0.348597f
C4577 C7_N_btm.t119 VSS 0.386613f
C4578 C7_N_btm.n185 VSS 0.117817f
C4579 C7_N_btm.t92 VSS 0.348597f
C4580 C7_N_btm.t44 VSS 0.348597f
C4581 C7_N_btm.t80 VSS 0.348597f
C4582 C7_N_btm.t9 VSS 0.348597f
C4583 C7_N_btm.t13 VSS 0.348597f
C4584 C7_N_btm.t99 VSS 0.348597f
C4585 C7_N_btm.t5 VSS 0.348597f
C4586 C7_N_btm.t94 VSS 0.348597f
C4587 C7_N_btm.t46 VSS 0.348597f
C4588 C7_N_btm.t30 VSS 0.348597f
C4589 C7_N_btm.t116 VSS 0.348597f
C4590 C7_N_btm.t15 VSS 0.348597f
C4591 C7_N_btm.t51 VSS 0.348597f
C4592 C7_N_btm.t10 VSS 0.348597f
C4593 C7_N_btm.t39 VSS 0.348597f
C4594 C7_N_btm.t48 VSS 0.348597f
C4595 C7_N_btm.t32 VSS 0.348597f
C4596 C7_N_btm.t62 VSS 0.348597f
C4597 C7_N_btm.t54 VSS 0.386613f
C4598 C7_N_btm.n242 VSS 0.117817f
C4599 C7_N_btm.t68 VSS 0.386613f
C4600 C7_N_btm.t100 VSS 0.348597f
C4601 C7_N_btm.t73 VSS 0.348597f
C4602 C7_N_btm.t121 VSS 0.385972f
C4603 C7_N_btm.t81 VSS 0.385972f
C4604 C7_N_btm.t57 VSS 0.385972f
C4605 C7_N_btm.t88 VSS 0.385972f
C4606 C7_N_btm.t63 VSS 0.385972f
C4607 C7_N_btm.t34 VSS 0.385972f
C4608 C7_N_btm.t71 VSS 0.385972f
C4609 C7_N_btm.t117 VSS 0.385972f
C4610 C7_N_btm.t55 VSS 0.385972f
C4611 C7_N_btm.t112 VSS 0.385972f
C4612 C7_N_btm.t16 VSS 0.385972f
C4613 C7_N_btm.t129 VSS 0.385972f
C4614 C7_N_btm.t31 VSS 0.385972f
C4615 C7_N_btm.t24 VSS 0.385972f
C4616 C7_N_btm.t37 VSS 0.348597f
C4617 C7_N_btm.t6 VSS 0.348597f
C4618 C7_N_btm.t105 VSS 0.386613f
C4619 C7_N_btm.t115 VSS 0.348597f
C4620 C7_N_btm.t83 VSS 0.348597f
C4621 C7_N_btm.t12 VSS 0.386613f
C4622 C7_N_btm.t86 VSS 0.386613f
C4623 C7_N_btm.t110 VSS 0.348597f
C4624 C7_N_btm.t60 VSS 0.386613f
C4625 C7_N_btm.t29 VSS 0.348597f
C4626 C7_N_btm.t72 VSS 0.386613f
C4627 C7_N_btm.t17 VSS 0.348597f
C4628 C7_N_btm.t53 VSS 0.386613f
C4629 C7_N_btm.t89 VSS 0.386613f
C4630 C7_N_btm.t35 VSS 0.386613f
C4631 C7_N_btm.t64 VSS 0.348597f
C4632 C7_N_btm.t77 VSS 0.386613f
C4633 C7_N_btm.t111 VSS 0.348597f
C4634 C7_N_btm.t25 VSS 0.386613f
C4635 C7_N_btm.t40 VSS 0.348597f
C4636 C7_N_btm.t66 VSS 0.386613f
C4637 C7_N_btm.t104 VSS 0.386613f
C4638 C7_N_btm.t126 VSS 0.386613f
C4639 C7_N_btm.t38 VSS 0.348597f
C4640 C7_N_btm.t96 VSS 0.386613f
C4641 C7_N_btm.t70 VSS 0.348597f
C4642 C7_N_btm.t47 VSS 0.386613f
C4643 C7_N_btm.n337 VSS 0.146274f
C4644 C7_N_btm.t108 VSS 0.348597f
C4645 C7_N_btm.t11 VSS 0.386613f
C4646 C7_N_btm.t133 VSS 0.387263f
C4647 C7_N_btm.n344 VSS 0.214334f
C4648 a_13273_44868.n9 VSS 0.431905f
C4649 a_13273_44868.n11 VSS 0.101145f
C4650 a_13273_44868.n14 VSS 0.215217f
C4651 a_13273_44868.n16 VSS 0.202755f
C4652 a_13273_44868.n17 VSS 0.127109f
C4653 a_13273_44868.n18 VSS 0.174362f
C4654 a_13273_44868.n23 VSS 0.253846f
C4655 a_13273_44868.n24 VSS 0.180845f
C4656 C8_N_btm.n0 VSS 0.220789f
C4657 C8_N_btm.n1 VSS 0.214012f
C4658 C8_N_btm.n2 VSS 0.853964f
C4659 C8_N_btm.n3 VSS 0.399375f
C4660 C8_N_btm.n4 VSS 0.566193f
C4661 C8_N_btm.n5 VSS 0.402318f
C4662 C8_N_btm.n6 VSS 0.437265f
C4663 C8_N_btm.n8 VSS 1.2599f
C4664 C8_N_btm.t270 VSS 0.325831f
C4665 C8_N_btm.n10 VSS 0.102832f
C4666 C8_N_btm.t263 VSS 0.325831f
C4667 C8_N_btm.n11 VSS 0.102832f
C4668 C8_N_btm.t269 VSS 0.325831f
C4669 C8_N_btm.n12 VSS 0.102832f
C4670 C8_N_btm.t124 VSS 0.313436f
C4671 C8_N_btm.t271 VSS 0.325831f
C4672 C8_N_btm.t240 VSS 0.313436f
C4673 C8_N_btm.t197 VSS 0.313436f
C4674 C8_N_btm.t39 VSS 0.313436f
C4675 C8_N_btm.t63 VSS 0.282615f
C4676 C8_N_btm.t32 VSS 0.282615f
C4677 C8_N_btm.t150 VSS 0.313436f
C4678 C8_N_btm.t144 VSS 0.313436f
C4679 C8_N_btm.t57 VSS 0.282615f
C4680 C8_N_btm.t199 VSS 0.282615f
C4681 C8_N_btm.t111 VSS 0.313436f
C4682 C8_N_btm.t244 VSS 0.282615f
C4683 C8_N_btm.t153 VSS 0.282615f
C4684 C8_N_btm.t217 VSS 0.282615f
C4685 C8_N_btm.t139 VSS 0.282615f
C4686 C8_N_btm.t204 VSS 0.313436f
C4687 C8_N_btm.t164 VSS 0.313436f
C4688 C8_N_btm.t214 VSS 0.313436f
C4689 C8_N_btm.t52 VSS 0.313436f
C4690 C8_N_btm.t184 VSS 0.282615f
C4691 C8_N_btm.t27 VSS 0.282615f
C4692 C8_N_btm.t213 VSS 0.313436f
C4693 C8_N_btm.t89 VSS 0.313436f
C4694 C8_N_btm.t231 VSS 0.282615f
C4695 C8_N_btm.t25 VSS 0.282615f
C4696 C8_N_btm.t264 VSS 0.325831f
C4697 C8_N_btm.n156 VSS 0.118588f
C4698 C8_N_btm.t268 VSS 0.325831f
C4699 C8_N_btm.t265 VSS 0.325831f
C4700 C8_N_btm.n159 VSS 0.102832f
C4701 C8_N_btm.t262 VSS 0.325831f
C4702 C8_N_btm.n160 VSS 0.102832f
C4703 C8_N_btm.t99 VSS 0.313436f
C4704 C8_N_btm.t171 VSS 0.282615f
C4705 C8_N_btm.t116 VSS 0.282615f
C4706 C8_N_btm.t138 VSS 0.313436f
C4707 C8_N_btm.t267 VSS 0.325831f
C4708 C8_N_btm.n169 VSS 0.118588f
C4709 C8_N_btm.t202 VSS 0.282615f
C4710 C8_N_btm.n173 VSS 0.102832f
C4711 C8_N_btm.t117 VSS 0.313436f
C4712 C8_N_btm.t108 VSS 0.282615f
C4713 C8_N_btm.t253 VSS 0.282615f
C4714 C8_N_btm.t82 VSS 0.282615f
C4715 C8_N_btm.t148 VSS 0.313436f
C4716 C8_N_btm.t180 VSS 0.313436f
C4717 C8_N_btm.t104 VSS 0.282615f
C4718 C8_N_btm.t55 VSS 0.282615f
C4719 C8_N_btm.t129 VSS 0.282615f
C4720 C8_N_btm.t77 VSS 0.313436f
C4721 C8_N_btm.t51 VSS 0.282615f
C4722 C8_N_btm.t19 VSS 0.313436f
C4723 C8_N_btm.t70 VSS 0.282615f
C4724 C8_N_btm.t245 VSS 0.282615f
C4725 C8_N_btm.t46 VSS 0.282615f
C4726 C8_N_btm.t110 VSS 0.313436f
C4727 C8_N_btm.t132 VSS 0.313436f
C4728 C8_N_btm.t66 VSS 0.282615f
C4729 C8_N_btm.t16 VSS 0.282615f
C4730 C8_N_btm.t95 VSS 0.282615f
C4731 C8_N_btm.t40 VSS 0.313436f
C4732 C8_N_btm.t13 VSS 0.282615f
C4733 C8_N_btm.t189 VSS 0.313436f
C4734 C8_N_btm.t33 VSS 0.282615f
C4735 C8_N_btm.t212 VSS 0.282615f
C4736 C8_N_btm.t26 VSS 0.282615f
C4737 C8_N_btm.t72 VSS 0.313436f
C4738 C8_N_btm.t34 VSS 0.313436f
C4739 C8_N_btm.t135 VSS 0.282615f
C4740 C8_N_btm.t198 VSS 0.282615f
C4741 C8_N_btm.t14 VSS 0.313436f
C4742 C8_N_btm.t7 VSS 0.313436f
C4743 C8_N_btm.t174 VSS 0.282615f
C4744 C8_N_btm.t119 VSS 0.282615f
C4745 C8_N_btm.t206 VSS 0.282615f
C4746 C8_N_btm.t140 VSS 0.313436f
C4747 C8_N_btm.t232 VSS 0.282615f
C4748 C8_N_btm.t193 VSS 0.313436f
C4749 C8_N_btm.t223 VSS 0.282615f
C4750 C8_N_btm.t162 VSS 0.282615f
C4751 C8_N_btm.t226 VSS 0.282615f
C4752 C8_N_btm.t209 VSS 0.313436f
C4753 C8_N_btm.t127 VSS 0.282615f
C4754 C8_N_btm.t75 VSS 0.282615f
C4755 C8_N_btm.t157 VSS 0.282615f
C4756 C8_N_btm.t100 VSS 0.313436f
C4757 C8_N_btm.t256 VSS 0.313436f
C4758 C8_N_btm.t190 VSS 0.282615f
C4759 C8_N_btm.t250 VSS 0.282615f
C4760 C8_N_btm.t185 VSS 0.282615f
C4761 C8_N_btm.t98 VSS 0.282615f
C4762 C8_N_btm.t152 VSS 0.282615f
C4763 C8_N_btm.t234 VSS 0.313436f
C4764 C8_N_btm.t73 VSS 0.313436f
C4765 C8_N_btm.t149 VSS 0.313436f
C4766 C8_N_btm.t230 VSS 0.313436f
C4767 C8_N_btm.t187 VSS 0.313436f
C4768 C8_N_btm.t200 VSS 0.282615f
C4769 C8_N_btm.t114 VSS 0.282615f
C4770 C8_N_btm.t169 VSS 0.282615f
C4771 C8_N_btm.t258 VSS 0.282615f
C4772 C8_N_btm.t155 VSS 0.282615f
C4773 C8_N_btm.t219 VSS 0.282615f
C4774 C8_N_btm.t126 VSS 0.282615f
C4775 C8_N_btm.t207 VSS 0.282615f
C4776 C8_N_btm.t94 VSS 0.282615f
C4777 C8_N_btm.t178 VSS 0.282615f
C4778 C8_N_btm.t259 VSS 0.282615f
C4779 C8_N_btm.t160 VSS 0.282615f
C4780 C8_N_btm.t224 VSS 0.282615f
C4781 C8_N_btm.t31 VSS 0.282615f
C4782 C8_N_btm.t211 VSS 0.282615f
C4783 C8_N_btm.t23 VSS 0.282615f
C4784 C8_N_btm.t59 VSS 0.282615f
C4785 C8_N_btm.t218 VSS 0.282615f
C4786 C8_N_btm.t50 VSS 0.282615f
C4787 C8_N_btm.t229 VSS 0.282615f
C4788 C8_N_btm.t35 VSS 0.282615f
C4789 C8_N_btm.t88 VSS 0.282615f
C4790 C8_N_btm.t21 VSS 0.282615f
C4791 C8_N_btm.t83 VSS 0.282615f
C4792 C8_N_btm.t136 VSS 0.282615f
C4793 C8_N_btm.t60 VSS 0.282615f
C4794 C8_N_btm.t113 VSS 0.282615f
C4795 C8_N_btm.t254 VSS 0.313436f
C4796 C8_N_btm.t29 VSS 0.282615f
C4797 C8_N_btm.t238 VSS 0.282615f
C4798 C8_N_btm.t56 VSS 0.282615f
C4799 C8_N_btm.t246 VSS 0.282615f
C4800 C8_N_btm.t93 VSS 0.282615f
C4801 C8_N_btm.t133 VSS 0.282615f
C4802 C8_N_btm.t210 VSS 0.282615f
C4803 C8_N_btm.t130 VSS 0.282615f
C4804 C8_N_btm.t222 VSS 0.282615f
C4805 C8_N_btm.t158 VSS 0.282615f
C4806 C8_N_btm.t237 VSS 0.282615f
C4807 C8_N_btm.t173 VSS 0.282615f
C4808 C8_N_btm.t118 VSS 0.282615f
C4809 C8_N_btm.t205 VSS 0.282615f
C4810 C8_N_btm.t125 VSS 0.282615f
C4811 C8_N_btm.t74 VSS 0.282615f
C4812 C8_N_btm.t154 VSS 0.282615f
C4813 C8_N_btm.t87 VSS 0.282615f
C4814 C8_N_btm.t168 VSS 0.282615f
C4815 C8_N_btm.t112 VSS 0.282615f
C4816 C8_N_btm.t49 VSS 0.282615f
C4817 C8_N_btm.t252 VSS 0.282615f
C4818 C8_N_btm.t71 VSS 0.282615f
C4819 C8_N_btm.t20 VSS 0.282615f
C4820 C8_N_btm.t81 VSS 0.282615f
C4821 C8_N_btm.t30 VSS 0.282615f
C4822 C8_N_btm.t107 VSS 0.282615f
C4823 C8_N_btm.t43 VSS 0.282615f
C4824 C8_N_btm.t9 VSS 0.313436f
C4825 C8_N_btm.t122 VSS 0.282615f
C4826 C8_N_btm.t53 VSS 0.313436f
C4827 C8_N_btm.t102 VSS 0.282615f
C4828 C8_N_btm.t176 VSS 0.282615f
C4829 C8_N_btm.t92 VSS 0.282615f
C4830 C8_N_btm.t142 VSS 0.282615f
C4831 C8_N_btm.t78 VSS 0.282615f
C4832 C8_N_btm.t131 VSS 0.282615f
C4833 C8_N_btm.t195 VSS 0.282615f
C4834 C8_N_btm.t106 VSS 0.282615f
C4835 C8_N_btm.t182 VSS 0.282615f
C4836 C8_N_btm.t8 VSS 0.282615f
C4837 C8_N_btm.t147 VSS 0.282615f
C4838 C8_N_btm.t228 VSS 0.282615f
C4839 C8_N_btm.t134 VSS 0.282615f
C4840 C8_N_btm.t196 VSS 0.282615f
C4841 C8_N_btm.t243 VSS 0.282615f
C4842 C8_N_btm.t183 VSS 0.282615f
C4843 C8_N_btm.t11 VSS 0.282615f
C4844 C8_N_btm.t37 VSS 0.282615f
C4845 C8_N_btm.t233 VSS 0.282615f
C4846 C8_N_btm.t121 VSS 0.282615f
C4847 C8_N_btm.t203 VSS 0.282615f
C4848 C8_N_btm.t15 VSS 0.282615f
C4849 C8_N_btm.t64 VSS 0.282615f
C4850 C8_N_btm.t186 VSS 0.282615f
C4851 C8_N_btm.t62 VSS 0.282615f
C4852 C8_N_btm.t161 VSS 0.282615f
C4853 C8_N_btm.t38 VSS 0.282615f
C4854 C8_N_btm.t91 VSS 0.282615f
C4855 C8_N_btm.t159 VSS 0.313436f
C4856 C8_N_btm.t261 VSS 0.313436f
C4857 C8_N_btm.t68 VSS 0.282615f
C4858 C8_N_btm.t18 VSS 0.282615f
C4859 C8_N_btm.t96 VSS 0.282615f
C4860 C8_N_btm.t42 VSS 0.282615f
C4861 C8_N_btm.t235 VSS 0.282615f
C4862 C8_N_btm.t44 VSS 0.282615f
C4863 C8_N_btm.t97 VSS 0.282615f
C4864 C8_N_btm.t179 VSS 0.282615f
C4865 C8_N_btm.t41 VSS 0.282615f
C4866 C8_N_btm.t208 VSS 0.282615f
C4867 C8_N_btm.t17 VSS 0.282615f
C4868 C8_N_btm.t220 VSS 0.282615f
C4869 C8_N_btm.t156 VSS 0.282615f
C4870 C8_N_btm.t6 VSS 0.282615f
C4871 C8_N_btm.t170 VSS 0.282615f
C4872 C8_N_btm.t115 VSS 0.282615f
C4873 C8_N_btm.t201 VSS 0.282615f
C4874 C8_N_btm.t123 VSS 0.282615f
C4875 C8_N_btm.t216 VSS 0.282615f
C4876 C8_N_btm.t151 VSS 0.282615f
C4877 C8_N_btm.t86 VSS 0.282615f
C4878 C8_N_btm.t166 VSS 0.282615f
C4879 C8_N_btm.t109 VSS 0.282615f
C4880 C8_N_btm.t120 VSS 0.282615f
C4881 C8_N_btm.t249 VSS 0.282615f
C4882 C8_N_btm.t69 VSS 0.282615f
C4883 C8_N_btm.t146 VSS 0.282615f
C4884 C8_N_btm.t80 VSS 0.282615f
C4885 C8_N_btm.t28 VSS 0.313436f
C4886 C8_N_btm.t167 VSS 0.282615f
C4887 C8_N_btm.t90 VSS 0.313436f
C4888 C8_N_btm.t141 VSS 0.282615f
C4889 C8_N_btm.t221 VSS 0.282615f
C4890 C8_N_btm.t128 VSS 0.282615f
C4891 C8_N_btm.t192 VSS 0.313436f
C4892 C8_N_btm.t24 VSS 0.313436f
C4893 C8_N_btm.t227 VSS 0.282615f
C4894 C8_N_btm.t48 VSS 0.282615f
C4895 C8_N_btm.t239 VSS 0.282615f
C4896 C8_N_btm.t181 VSS 0.313436f
C4897 C8_N_btm.t215 VSS 0.282615f
C4898 C8_N_btm.t260 VSS 0.313436f
C4899 C8_N_btm.t191 VSS 0.282615f
C4900 C8_N_btm.t103 VSS 0.282615f
C4901 C8_N_btm.t175 VSS 0.282615f
C4902 C8_N_btm.t12 VSS 0.313436f
C4903 C8_N_btm.t61 VSS 0.313436f
C4904 C8_N_btm.t58 VSS 0.282615f
C4905 C8_N_btm.t85 VSS 0.282615f
C4906 C8_N_btm.t22 VSS 0.282615f
C4907 C8_N_btm.t225 VSS 0.313436f
C4908 C8_N_btm.t177 VSS 0.282615f
C4909 C8_N_btm.t242 VSS 0.313436f
C4910 C8_N_btm.t79 VSS 0.282615f
C4911 C8_N_btm.t145 VSS 0.282615f
C4912 C8_N_btm.t67 VSS 0.282615f
C4913 C8_N_btm.t248 VSS 0.313436f
C4914 C8_N_btm.t163 VSS 0.313436f
C4915 C8_N_btm.t101 VSS 0.282615f
C4916 C8_N_btm.t54 VSS 0.282615f
C4917 C8_N_btm.t76 VSS 0.313436f
C4918 C8_N_btm.t257 VSS 0.313436f
C4919 C8_N_btm.t47 VSS 0.282615f
C4920 C8_N_btm.t251 VSS 0.282615f
C4921 C8_N_btm.t241 VSS 0.282615f
C4922 C8_N_btm.t10 VSS 0.313436f
C4923 C8_N_btm.t36 VSS 0.282615f
C4924 C8_N_btm.t65 VSS 0.313436f
C4925 C8_N_btm.t247 VSS 0.282615f
C4926 C8_N_btm.t194 VSS 0.282615f
C4927 C8_N_btm.t105 VSS 0.282615f
C4928 C8_N_btm.t137 VSS 0.313436f
C4929 C8_N_btm.t84 VSS 0.282615f
C4930 C8_N_btm.t165 VSS 0.282615f
C4931 C8_N_btm.t255 VSS 0.282615f
C4932 C8_N_btm.t45 VSS 0.313436f
C4933 C8_N_btm.n890 VSS 0.118588f
C4934 C8_N_btm.t188 VSS 0.282615f
C4935 C8_N_btm.t143 VSS 0.282615f
C4936 C8_N_btm.t172 VSS 0.282615f
C4937 C8_N_btm.t236 VSS 0.313436f
C4938 C8_N_btm.t266 VSS 0.313964f
C4939 C8_N_btm.n903 VSS 0.165959f
C4940 a_10259_42870.n5 VSS 0.436003f
C4941 a_10259_42870.n10 VSS 0.253785f
C4942 a_10259_42870.n11 VSS 0.202454f
C4943 a_10259_42870.n17 VSS 0.205104f
C4944 a_10259_42870.n18 VSS 0.351774f
C4945 a_10259_42870.n20 VSS 0.104957f
C4946 a_10259_42870.n21 VSS 0.177234f
C4947 VDAC_Ni.n2 VSS 0.429559f
C4948 VDAC_Ni.t0 VSS 0.106007f
C4949 VDAC_Ni.n3 VSS 1.2327f
C4950 VDAC_Ni.n4 VSS 0.242952f
C4951 VDAC_Ni.n6 VSS 0.158267f
C4952 VDAC_Ni.n8 VSS 0.163297f
C4953 a_n1459_43236.n0 VSS 2.78033f
C4954 a_n1459_43236.n1 VSS 0.111416f
C4955 a_n1459_43236.n2 VSS 0.220076f
C4956 a_n1459_43236.n3 VSS 10.9698f
C4957 a_n1459_43236.n4 VSS 0.124002f
C4958 a_n1459_43236.n6 VSS 0.342464f
C4959 a_n1459_43236.n7 VSS 0.162913f
C4960 a_n1459_43236.n9 VSS 0.387885f
C4961 a_n1459_43236.n10 VSS 0.103904f
C4962 a_15730_45670.n6 VSS 0.172245f
C4963 a_15730_45670.n8 VSS 0.128032f
C4964 a_15730_45670.n16 VSS 0.190406f
C4965 a_15730_45670.n17 VSS 0.321765f
C4966 a_15730_45670.n18 VSS 0.147661f
C4967 a_15730_45670.n20 VSS 0.208515f
C4968 a_15730_45670.n21 VSS 0.259855f
C4969 a_15730_45670.n22 VSS 0.253425f
C4970 SMPL_ON_P.n0 VSS 0.180672f
C4971 SMPL_ON_P.n3 VSS 0.2207f
C4972 SMPL_ON_P.n6 VSS 0.30037f
C4973 SMPL_ON_P.n7 VSS 2.96463f
C4974 a_9096_45276.n1 VSS 1.15668f
C4975 a_9096_45276.n2 VSS 0.479071f
C4976 a_1053_45123.n6 VSS 0.132476f
C4977 a_1053_45123.n8 VSS 0.128824f
C4978 a_1053_45123.n9 VSS 0.143785f
C4979 a_1053_45123.n10 VSS 1.29444f
C4980 a_13524_46832.n7 VSS 0.106961f
C4981 a_13524_46832.n8 VSS 0.393722f
C4982 a_13524_46832.n10 VSS 0.529261f
C4983 a_13524_46832.n11 VSS 0.206118f
C4984 a_13524_46832.n14 VSS 0.275443f
C4985 a_13524_46832.n15 VSS 0.322357f
C4986 a_13524_46832.n16 VSS 0.502786f
C4987 a_13524_46832.n17 VSS 0.232768f
C4988 a_n53_44363.n4 VSS 0.192414f
C4989 a_n53_44363.n7 VSS 0.160362f
C4990 a_n53_44363.n9 VSS 0.263905f
C4991 a_n53_44363.n11 VSS 0.157696f
C4992 a_n53_44363.n13 VSS 0.161656f
C4993 a_n53_44363.n15 VSS 0.244119f
C4994 a_n53_44363.n17 VSS 0.220309f
C4995 VREF.t6 VSS 0.378661f
C4996 VREF.t73 VSS 0.373633f
C4997 VREF.n0 VSS 1.05072f
C4998 VREF.t70 VSS 0.373633f
C4999 VREF.n1 VSS 0.543604f
C5000 VREF.t22 VSS 0.373633f
C5001 VREF.n2 VSS 0.543604f
C5002 VREF.t72 VSS 0.373633f
C5003 VREF.n3 VSS 0.542031f
C5004 VREF.t5 VSS 0.373633f
C5005 VREF.n4 VSS 0.542031f
C5006 VREF.t69 VSS 0.182453f
C5007 VREF.t21 VSS 0.182453f
C5008 VREF.n5 VSS 0.45929f
C5009 VREF.n6 VSS 0.557667f
C5010 VREF.t20 VSS 0.182453f
C5011 VREF.t2 VSS 0.182453f
C5012 VREF.n7 VSS 0.45929f
C5013 VREF.n8 VSS 0.560813f
C5014 VREF.t0 VSS 0.182453f
C5015 VREF.t3 VSS 0.182453f
C5016 VREF.n9 VSS 0.45929f
C5017 VREF.n10 VSS 0.55924f
C5018 VREF.t1 VSS 0.182453f
C5019 VREF.t13 VSS 0.182453f
C5020 VREF.n11 VSS 0.45929f
C5021 VREF.n12 VSS 0.55924f
C5022 VREF.t12 VSS 0.182453f
C5023 VREF.t17 VSS 0.182453f
C5024 VREF.n13 VSS 0.45929f
C5025 VREF.n14 VSS 0.560813f
C5026 VREF.t18 VSS 0.182453f
C5027 VREF.t15 VSS 0.182453f
C5028 VREF.n15 VSS 0.45929f
C5029 VREF.n16 VSS 0.55924f
C5030 VREF.t16 VSS 0.182453f
C5031 VREF.t11 VSS 0.182453f
C5032 VREF.n17 VSS 0.45929f
C5033 VREF.n18 VSS 0.55924f
C5034 VREF.t14 VSS 0.182453f
C5035 VREF.t66 VSS 0.182453f
C5036 VREF.n19 VSS 0.45929f
C5037 VREF.n20 VSS 0.55924f
C5038 VREF.t68 VSS 0.182453f
C5039 VREF.t54 VSS 0.182453f
C5040 VREF.n21 VSS 0.45929f
C5041 VREF.n22 VSS 0.55924f
C5042 VREF.t61 VSS 0.182453f
C5043 VREF.t63 VSS 0.182453f
C5044 VREF.n23 VSS 0.45929f
C5045 VREF.n24 VSS 0.560813f
C5046 VREF.t67 VSS 0.182453f
C5047 VREF.t55 VSS 0.182453f
C5048 VREF.n25 VSS 0.45929f
C5049 VREF.n26 VSS 0.55924f
C5050 VREF.t60 VSS 0.182453f
C5051 VREF.t53 VSS 0.182453f
C5052 VREF.n27 VSS 0.45929f
C5053 VREF.n28 VSS 0.55924f
C5054 VREF.t56 VSS 0.182453f
C5055 VREF.t62 VSS 0.182453f
C5056 VREF.n29 VSS 0.45929f
C5057 VREF.n30 VSS 0.55924f
C5058 VREF.t64 VSS 0.182453f
C5059 VREF.t58 VSS 0.182453f
C5060 VREF.n31 VSS 0.45929f
C5061 VREF.n32 VSS 0.55924f
C5062 VREF.t59 VSS 0.182453f
C5063 VREF.t57 VSS 0.182453f
C5064 VREF.n33 VSS 0.45929f
C5065 VREF.n34 VSS 0.560813f
C5066 VREF.t65 VSS 0.757234f
C5067 VREF.n35 VSS 2.26063f
C5068 VREF.t4 VSS 0.378661f
C5069 VREF.t51 VSS 0.373633f
C5070 VREF.n36 VSS 1.05072f
C5071 VREF.t71 VSS 0.373633f
C5072 VREF.n37 VSS 0.543604f
C5073 VREF.t10 VSS 0.373633f
C5074 VREF.n38 VSS 0.543604f
C5075 VREF.t7 VSS 0.373633f
C5076 VREF.n39 VSS 0.542031f
C5077 VREF.t52 VSS 0.373633f
C5078 VREF.n40 VSS 0.542031f
C5079 VREF.t8 VSS 0.182453f
C5080 VREF.t19 VSS 0.182453f
C5081 VREF.n41 VSS 0.45929f
C5082 VREF.n42 VSS 0.557667f
C5083 VREF.t50 VSS 0.182453f
C5084 VREF.t9 VSS 0.182453f
C5085 VREF.n43 VSS 0.45929f
C5086 VREF.n44 VSS 0.560813f
C5087 VREF.t47 VSS 0.182453f
C5088 VREF.t49 VSS 0.182453f
C5089 VREF.n45 VSS 0.45929f
C5090 VREF.n46 VSS 0.55924f
C5091 VREF.t25 VSS 0.182453f
C5092 VREF.t48 VSS 0.182453f
C5093 VREF.n47 VSS 0.45929f
C5094 VREF.n48 VSS 0.55924f
C5095 VREF.t27 VSS 0.182453f
C5096 VREF.t29 VSS 0.182453f
C5097 VREF.n49 VSS 0.45929f
C5098 VREF.n50 VSS 0.560813f
C5099 VREF.t23 VSS 0.182453f
C5100 VREF.t28 VSS 0.182453f
C5101 VREF.n51 VSS 0.45929f
C5102 VREF.n52 VSS 0.55924f
C5103 VREF.t26 VSS 0.182453f
C5104 VREF.t30 VSS 0.182453f
C5105 VREF.n53 VSS 0.45929f
C5106 VREF.n54 VSS 0.55924f
C5107 VREF.t32 VSS 0.182453f
C5108 VREF.t24 VSS 0.182453f
C5109 VREF.n55 VSS 0.45929f
C5110 VREF.n56 VSS 0.55924f
C5111 VREF.t37 VSS 0.182453f
C5112 VREF.t45 VSS 0.182453f
C5113 VREF.n57 VSS 0.45929f
C5114 VREF.n58 VSS 0.55924f
C5115 VREF.t31 VSS 0.182453f
C5116 VREF.t34 VSS 0.182453f
C5117 VREF.n59 VSS 0.45929f
C5118 VREF.n60 VSS 0.560813f
C5119 VREF.t40 VSS 0.182453f
C5120 VREF.t36 VSS 0.182453f
C5121 VREF.n61 VSS 0.45929f
C5122 VREF.n62 VSS 0.55924f
C5123 VREF.t43 VSS 0.182453f
C5124 VREF.t44 VSS 0.182453f
C5125 VREF.n63 VSS 0.45929f
C5126 VREF.n64 VSS 0.55924f
C5127 VREF.t42 VSS 0.182453f
C5128 VREF.t39 VSS 0.182453f
C5129 VREF.n65 VSS 0.45929f
C5130 VREF.n66 VSS 0.55924f
C5131 VREF.t38 VSS 0.182453f
C5132 VREF.t35 VSS 0.182453f
C5133 VREF.n67 VSS 0.45929f
C5134 VREF.n68 VSS 0.55924f
C5135 VREF.t41 VSS 0.182453f
C5136 VREF.t46 VSS 0.182453f
C5137 VREF.n69 VSS 0.45929f
C5138 VREF.n70 VSS 0.560813f
C5139 VREF.t33 VSS 0.757234f
C5140 VREF.n71 VSS 12.9035f
C5141 VREF.n72 VSS 16.917599f
C5142 a_22812_30659.t5 VSS 0.55181f
C5143 a_22812_30659.t9 VSS 0.551895f
C5144 a_22812_30659.t17 VSS 0.55181f
C5145 a_22812_30659.n0 VSS 0.407565f
C5146 a_22812_30659.t10 VSS 0.55181f
C5147 a_22812_30659.n1 VSS 0.207448f
C5148 a_22812_30659.t16 VSS 0.55181f
C5149 a_22812_30659.n2 VSS 0.207448f
C5150 a_22812_30659.t6 VSS 0.55181f
C5151 a_22812_30659.n3 VSS 0.207448f
C5152 a_22812_30659.t8 VSS 0.55181f
C5153 a_22812_30659.n4 VSS 0.207448f
C5154 a_22812_30659.t4 VSS 0.55181f
C5155 a_22812_30659.n5 VSS 0.207448f
C5156 a_22812_30659.t12 VSS 0.55181f
C5157 a_22812_30659.n6 VSS 0.207448f
C5158 a_22812_30659.t18 VSS 0.55181f
C5159 a_22812_30659.n7 VSS 0.207448f
C5160 a_22812_30659.t14 VSS 0.55181f
C5161 a_22812_30659.n8 VSS 0.207448f
C5162 a_22812_30659.t19 VSS 0.55181f
C5163 a_22812_30659.n9 VSS 0.207448f
C5164 a_22812_30659.t15 VSS 0.55181f
C5165 a_22812_30659.n10 VSS 0.207448f
C5166 a_22812_30659.t11 VSS 0.55181f
C5167 a_22812_30659.n11 VSS 0.207448f
C5168 a_22812_30659.t7 VSS 0.55181f
C5169 a_22812_30659.n12 VSS 0.207448f
C5170 a_22812_30659.t13 VSS 0.55181f
C5171 a_22812_30659.n13 VSS 0.20705f
C5172 a_22812_30659.n14 VSS 2.38139f
C5173 a_22812_30659.n16 VSS 1.86166f
C5174 w_1375_34946.n7 VSS 0.109775f
C5175 w_1375_34946.n9 VSS 0.45959f
C5176 w_1375_34946.n14 VSS 0.113467f
C5177 w_1375_34946.n15 VSS 0.147261f
C5178 w_1375_34946.n17 VSS 0.262162f
C5179 w_1375_34946.n19 VSS 0.540375f
C5180 w_1375_34946.n20 VSS 1.17135f
C5181 w_1375_34946.n21 VSS 2.23079f
C5182 w_1375_34946.n23 VSS 1.1728f
C5183 w_1375_34946.n24 VSS 0.148446f
C5184 w_1375_34946.n25 VSS 1.17425f
C5185 w_1375_34946.n27 VSS 2.23079f
C5186 w_1375_34946.n28 VSS 1.17255f
C5187 w_1375_34946.n30 VSS 0.259044f
C5188 w_1375_34946.n31 VSS 0.568321f
C5189 w_1375_34946.n32 VSS 0.138906f
C5190 w_1375_34946.n33 VSS 0.169733f
C5191 w_1375_34946.n34 VSS 0.211327f
C5192 w_1375_34946.n35 VSS 0.240728f
C5193 w_1375_34946.n36 VSS 0.134774f
C5194 w_1375_34946.n37 VSS 3.24247f
C5195 w_1375_34946.t5 VSS 5.81627f
C5196 w_1375_34946.n38 VSS 5.60723f
C5197 w_1375_34946.t2 VSS 5.84551f
C5198 w_1375_34946.n39 VSS 3.4195f
C5199 w_1375_34946.n40 VSS 0.136143f
C5200 w_1375_34946.n41 VSS 0.122267f
C5201 w_1375_34946.n43 VSS 0.496373f
C5202 w_1375_34946.n44 VSS 0.540045f
C5203 w_1375_34946.n45 VSS 0.174252f
C5204 w_1375_34946.n48 VSS 0.302685f
C5205 w_1375_34946.t14 VSS 0.202569f
C5206 w_1375_34946.t16 VSS 0.150361f
C5207 w_1375_34946.t10 VSS 0.296285f
C5208 w_1375_34946.t12 VSS 0.150361f
C5209 w_1375_34946.n49 VSS 0.100241f
C5210 w_1375_34946.n54 VSS 0.140862f
C5211 w_1375_34946.t0 VSS 0.149521f
C5212 a_n1123_35174.n1 VSS 1.72358f
C5213 a_n1123_35174.n2 VSS 1.7928f
C5214 a_n1123_35174.n3 VSS 0.393605f
C5215 a_n1123_35174.n4 VSS 0.438125f
C5216 a_n1123_35174.n5 VSS 0.532591f
C5217 a_n1123_35174.n6 VSS 1.72657f
C5218 a_n1123_35174.t6 VSS 4.75589f
C5219 a_n1123_35174.n7 VSS 3.74793f
C5220 a_n1123_35174.t4 VSS 4.75589f
C5221 a_n1123_35174.n8 VSS 1.67055f
C5222 a_n1123_35174.n9 VSS 0.17189f
C5223 a_n1123_35174.n10 VSS 0.172136f
C5224 a_n1123_35174.n11 VSS 0.441752f
C5225 a_n1123_35174.n12 VSS 0.397456f
C5226 a_n1123_35174.t5 VSS 4.75589f
C5227 a_n1123_35174.t7 VSS 4.75589f
C5228 a_n1123_35174.n13 VSS 3.7613f
C5229 a_n1123_35174.n14 VSS 0.435629f
C5230 a_n1123_35174.n15 VSS 0.44208f
C5231 a_n1123_35174.n16 VSS 0.512191f
C5232 C9_P_btm.n0 VSS 0.189504f
C5233 C9_P_btm.n1 VSS 0.183284f
C5234 C9_P_btm.n2 VSS 0.576048f
C5235 C9_P_btm.n3 VSS 0.183284f
C5236 C9_P_btm.n4 VSS 0.295064f
C5237 C9_P_btm.n5 VSS 0.183284f
C5238 C9_P_btm.n6 VSS 0.467877f
C5239 C9_P_btm.n7 VSS 0.27827f
C5240 C9_P_btm.n8 VSS 0.271863f
C5241 C9_P_btm.n9 VSS 0.442689f
C5242 C9_P_btm.n10 VSS 0.26427f
C5243 C9_P_btm.t4 VSS 0.414648f
C5244 C9_P_btm.n11 VSS 0.330821f
C5245 C9_P_btm.n12 VSS 0.281049f
C5246 C9_P_btm.n13 VSS 0.274975f
C5247 C9_P_btm.n14 VSS 0.447511f
C5248 C9_P_btm.n15 VSS 1.10449f
C5249 C9_P_btm.t18 VSS 0.279048f
C5250 C9_P_btm.t16 VSS 0.279048f
C5251 C9_P_btm.t17 VSS 0.279048f
C5252 C9_P_btm.t21 VSS 0.279048f
C5253 C9_P_btm.t351 VSS 0.268433f
C5254 C9_P_btm.t117 VSS 0.268433f
C5255 C9_P_btm.t231 VSS 0.268433f
C5256 C9_P_btm.t252 VSS 0.242037f
C5257 C9_P_btm.t492 VSS 0.242037f
C5258 C9_P_btm.t96 VSS 0.242037f
C5259 C9_P_btm.t410 VSS 0.268433f
C5260 C9_P_btm.t304 VSS 0.268433f
C5261 C9_P_btm.t163 VSS 0.242037f
C5262 C9_P_btm.t63 VSS 0.242037f
C5263 C9_P_btm.t179 VSS 0.242037f
C5264 C9_P_btm.t302 VSS 0.268433f
C5265 C9_P_btm.t384 VSS 0.268433f
C5266 C9_P_btm.t105 VSS 0.242037f
C5267 C9_P_btm.t154 VSS 0.242037f
C5268 C9_P_btm.t520 VSS 0.242037f
C5269 C9_P_btm.t201 VSS 0.268433f
C5270 C9_P_btm.t473 VSS 0.268433f
C5271 C9_P_btm.t447 VSS 0.242037f
C5272 C9_P_btm.t217 VSS 0.242037f
C5273 C9_P_btm.t327 VSS 0.242037f
C5274 C9_P_btm.t194 VSS 0.268433f
C5275 C9_P_btm.t138 VSS 0.268433f
C5276 C9_P_btm.t527 VSS 0.268433f
C5277 C9_P_btm.t443 VSS 0.268433f
C5278 C9_P_btm.t371 VSS 0.242037f
C5279 C9_P_btm.t452 VSS 0.242037f
C5280 C9_P_btm.t353 VSS 0.242037f
C5281 C9_P_btm.t496 VSS 0.242037f
C5282 C9_P_btm.t158 VSS 0.242037f
C5283 C9_P_btm.t438 VSS 0.242037f
C5284 C9_P_btm.t74 VSS 0.242037f
C5285 C9_P_btm.t414 VSS 0.242037f
C5286 C9_P_btm.t49 VSS 0.242037f
C5287 C9_P_btm.t386 VSS 0.242037f
C5288 C9_P_btm.t504 VSS 0.242037f
C5289 C9_P_btm.t224 VSS 0.242037f
C5290 C9_P_btm.t445 VSS 0.242037f
C5291 C9_P_btm.t79 VSS 0.242037f
C5292 C9_P_btm.t192 VSS 0.242037f
C5293 C9_P_btm.t229 VSS 0.242037f
C5294 C9_P_btm.t169 VSS 0.242037f
C5295 C9_P_btm.t55 VSS 0.242037f
C5296 C9_P_btm.t258 VSS 0.242037f
C5297 C9_P_btm.t350 VSS 0.242037f
C5298 C9_P_btm.t84 VSS 0.242037f
C5299 C9_P_btm.t531 VSS 0.242037f
C5300 C9_P_btm.t294 VSS 0.242037f
C5301 C9_P_btm.t174 VSS 0.242037f
C5302 C9_P_btm.t275 VSS 0.242037f
C5303 C9_P_btm.t122 VSS 0.242037f
C5304 C9_P_btm.t249 VSS 0.242037f
C5305 C9_P_btm.t357 VSS 0.242037f
C5306 C9_P_btm.t214 VSS 0.242037f
C5307 C9_P_btm.t348 VSS 0.242037f
C5308 C9_P_btm.t466 VSS 0.242037f
C5309 C9_P_btm.t296 VSS 0.242037f
C5310 C9_P_btm.t412 VSS 0.242037f
C5311 C9_P_btm.t48 VSS 0.242037f
C5312 C9_P_btm.t382 VSS 0.242037f
C5313 C9_P_btm.t503 VSS 0.242037f
C5314 C9_P_btm.t360 VSS 0.242037f
C5315 C9_P_btm.t477 VSS 0.242037f
C5316 C9_P_btm.t78 VSS 0.242037f
C5317 C9_P_btm.t321 VSS 0.268433f
C5318 C9_P_btm.t185 VSS 0.268433f
C5319 C9_P_btm.t97 VSS 0.242037f
C5320 C9_P_btm.t204 VSS 0.242037f
C5321 C9_P_btm.t103 VSS 0.242037f
C5322 C9_P_btm.t237 VSS 0.242037f
C5323 C9_P_btm.t127 VSS 0.242037f
C5324 C9_P_btm.t262 VSS 0.242037f
C5325 C9_P_btm.t178 VSS 0.242037f
C5326 C9_P_btm.t40 VSS 0.242037f
C5327 C9_P_btm.t435 VSS 0.242037f
C5328 C9_P_btm.t89 VSS 0.242037f
C5329 C9_P_btm.t460 VSS 0.242037f
C5330 C9_P_btm.t120 VSS 0.242037f
C5331 C9_P_btm.t118 VSS 0.242037f
C5332 C9_P_btm.t369 VSS 0.242037f
C5333 C9_P_btm.t26 VSS 0.268433f
C5334 C9_P_btm.t148 VSS 0.242037f
C5335 C9_P_btm.t248 VSS 0.242037f
C5336 C9_P_btm.t137 VSS 0.242037f
C5337 C9_P_btm.t292 VSS 0.242037f
C5338 C9_P_btm.t367 VSS 0.242037f
C5339 C9_P_btm.t209 VSS 0.242037f
C5340 C9_P_btm.t319 VSS 0.242037f
C5341 C9_P_btm.t454 VSS 0.242037f
C5342 C9_P_btm.t291 VSS 0.242037f
C5343 C9_P_btm.t407 VSS 0.242037f
C5344 C9_P_btm.t271 VSS 0.242037f
C5345 C9_P_btm.t376 VSS 0.242037f
C5346 C9_P_btm.t498 VSS 0.242037f
C5347 C9_P_btm.t325 VSS 0.242037f
C5348 C9_P_btm.t469 VSS 0.242037f
C5349 C9_P_btm.t75 VSS 0.242037f
C5350 C9_P_btm.t415 VSS 0.242037f
C5351 C9_P_btm.t50 VSS 0.242037f
C5352 C9_P_btm.t387 VSS 0.242037f
C5353 C9_P_btm.t505 VSS 0.242037f
C5354 C9_P_btm.t131 VSS 0.242037f
C5355 C9_P_btm.t478 VSS 0.242037f
C5356 C9_P_btm.t80 VSS 0.242037f
C5357 C9_P_btm.t523 VSS 0.242037f
C5358 C9_P_btm.t112 VSS 0.242037f
C5359 C9_P_btm.t170 VSS 0.242037f
C5360 C9_P_btm.t189 VSS 0.242037f
C5361 C9_P_btm.t141 VSS 0.242037f
C5362 C9_P_btm.t377 VSS 0.242037f
C5363 C9_P_btm.t235 VSS 0.242037f
C5364 C9_P_btm.t261 VSS 0.242037f
C5365 C9_P_btm.t338 VSS 0.242037f
C5366 C9_P_btm.t525 VSS 0.242037f
C5367 C9_P_btm.t290 VSS 0.242037f
C5368 C9_P_btm.t427 VSS 0.242037f
C5369 C9_P_btm.t269 VSS 0.242037f
C5370 C9_P_btm.t375 VSS 0.242037f
C5371 C9_P_btm.t397 VSS 0.242037f
C5372 C9_P_btm.t349 VSS 0.242037f
C5373 C9_P_btm.t467 VSS 0.242037f
C5374 C9_P_btm.t494 VSS 0.268433f
C5375 C9_P_btm.t123 VSS 0.242037f
C5376 C9_P_btm.t529 VSS 0.242037f
C5377 C9_P_btm.t406 VSS 0.242037f
C5378 C9_P_btm.t33 VSS 0.242037f
C5379 C9_P_btm.t430 VSS 0.242037f
C5380 C9_P_btm.t87 VSS 0.242037f
C5381 C9_P_btm.t457 VSS 0.242037f
C5382 C9_P_btm.t340 VSS 0.242037f
C5383 C9_P_btm.t54 VSS 0.242037f
C5384 C9_P_btm.t395 VSS 0.242037f
C5385 C9_P_btm.t535 VSS 0.242037f
C5386 C9_P_btm.t402 VSS 0.242037f
C5387 C9_P_btm.t287 VSS 0.242037f
C5388 C9_P_btm.t171 VSS 0.242037f
C5389 C9_P_btm.t316 VSS 0.242037f
C5390 C9_P_btm.t207 VSS 0.242037f
C5391 C9_P_btm.t337 VSS 0.242037f
C5392 C9_P_btm.t257 VSS 0.242037f
C5393 C9_P_btm.t135 VSS 0.242037f
C5394 C9_P_btm.t284 VSS 0.242037f
C5395 C9_P_btm.t166 VSS 0.242037f
C5396 C9_P_btm.t93 VSS 0.242037f
C5397 C9_P_btm.t203 VSS 0.242037f
C5398 C9_P_btm.t77 VSS 0.242037f
C5399 C9_P_btm.t234 VSS 0.242037f
C5400 C9_P_btm.t126 VSS 0.242037f
C5401 C9_P_btm.t501 VSS 0.242037f
C5402 C9_P_btm.t159 VSS 0.242037f
C5403 C9_P_btm.t36 VSS 0.242037f
C5404 C9_P_btm.t434 VSS 0.242037f
C5405 C9_P_btm.t64 VSS 0.242037f
C5406 C9_P_btm.t459 VSS 0.242037f
C5407 C9_P_btm.t513 VSS 0.242037f
C5408 C9_P_btm.t488 VSS 0.242037f
C5409 C9_P_btm.t368 VSS 0.242037f
C5410 C9_P_btm.t515 VSS 0.242037f
C5411 C9_P_btm.t396 VSS 0.242037f
C5412 C9_P_btm.t285 VSS 0.242037f
C5413 C9_P_btm.t300 VSS 0.242037f
C5414 C9_P_btm.t448 VSS 0.242037f
C5415 C9_P_btm.t313 VSS 0.268433f
C5416 C9_P_btm.t536 VSS 0.242037f
C5417 C9_P_btm.t151 VSS 0.268433f
C5418 C9_P_btm.t276 VSS 0.242037f
C5419 C9_P_btm.t380 VSS 0.242037f
C5420 C9_P_btm.t308 VSS 0.242037f
C5421 C9_P_btm.t419 VSS 0.242037f
C5422 C9_P_btm.t221 VSS 0.242037f
C5423 C9_P_btm.t391 VSS 0.242037f
C5424 C9_P_btm.t518 VSS 0.242037f
C5425 C9_P_btm.t142 VSS 0.242037f
C5426 C9_P_btm.t485 VSS 0.242037f
C5427 C9_P_btm.t85 VSS 0.242037f
C5428 C9_P_btm.t450 VSS 0.242037f
C5429 C9_P_btm.t58 VSS 0.242037f
C5430 C9_P_btm.t175 VSS 0.242037f
C5431 C9_P_btm.t46 VSS 0.242037f
C5432 C9_P_btm.t150 VSS 0.242037f
C5433 C9_P_btm.t250 VSS 0.242037f
C5434 C9_P_btm.t91 VSS 0.242037f
C5435 C9_P_btm.t223 VSS 0.242037f
C5436 C9_P_btm.t67 VSS 0.242037f
C5437 C9_P_btm.t181 VSS 0.242037f
C5438 C9_P_btm.t305 VSS 0.242037f
C5439 C9_P_btm.t162 VSS 0.242037f
C5440 C9_P_btm.t255 VSS 0.242037f
C5441 C9_P_btm.t364 VSS 0.242037f
C5442 C9_P_btm.t241 VSS 0.242037f
C5443 C9_P_btm.t334 VSS 0.242037f
C5444 C9_P_btm.t188 VSS 0.242037f
C5445 C9_P_btm.t312 VSS 0.242037f
C5446 C9_P_btm.t423 VSS 0.242037f
C5447 C9_P_btm.t281 VSS 0.242037f
C5448 C9_P_btm.t418 VSS 0.242037f
C5449 C9_P_btm.t116 VSS 0.242037f
C5450 C9_P_btm.t366 VSS 0.242037f
C5451 C9_P_btm.t484 VSS 0.242037f
C5452 C9_P_btm.t242 VSS 0.242037f
C5453 C9_P_btm.t449 VSS 0.242037f
C5454 C9_P_btm.t57 VSS 0.242037f
C5455 C9_P_btm.t425 VSS 0.242037f
C5456 C9_P_btm.t29 VSS 0.242037f
C5457 C9_P_btm.t147 VSS 0.242037f
C5458 C9_P_btm.t31 VSS 0.268433f
C5459 C9_P_btm.t301 VSS 0.268433f
C5460 C9_P_btm.t86 VSS 0.268433f
C5461 C9_P_btm.t451 VSS 0.268433f
C5462 C9_P_btm.t53 VSS 0.268433f
C5463 C9_P_btm.t426 VSS 0.242037f
C5464 C9_P_btm.t28 VSS 0.242037f
C5465 C9_P_btm.t152 VSS 0.242037f
C5466 C9_P_btm.t168 VSS 0.268433f
C5467 C9_P_btm.t210 VSS 0.268433f
C5468 C9_P_btm.t139 VSS 0.242037f
C5469 C9_P_btm.t298 VSS 0.242037f
C5470 C9_P_btm.t342 VSS 0.242037f
C5471 C9_P_btm.t82 VSS 0.268433f
C5472 C9_P_btm.t144 VSS 0.268433f
C5473 C9_P_btm.t243 VSS 0.242037f
C5474 C9_P_btm.t172 VSS 0.242037f
C5475 C9_P_btm.t270 VSS 0.242037f
C5476 C9_P_btm.t508 VSS 0.268433f
C5477 C9_P_btm.t399 VSS 0.268433f
C5478 C9_P_btm.t483 VSS 0.242037f
C5479 C9_P_btm.t83 VSS 0.242037f
C5480 C9_P_btm.t197 VSS 0.242037f
C5481 C9_P_btm.t19 VSS 0.279048f
C5482 C9_P_btm.t421 VSS 0.268433f
C5483 C9_P_btm.t14 VSS 0.279048f
C5484 C9_P_btm.t20 VSS 0.279048f
C5485 C9_P_btm.t15 VSS 0.279048f
C5486 C9_P_btm.t486 VSS 0.268433f
C5487 C9_P_btm.t393 VSS 0.242037f
C5488 C9_P_btm.t39 VSS 0.242037f
C5489 C9_P_btm.t299 VSS 0.242037f
C5490 C9_P_btm.t24 VSS 0.279048f
C5491 C9_P_btm.t13 VSS 0.279048f
C5492 C9_P_btm.n1046 VSS 0.101561f
C5493 C9_P_btm.t306 VSS 0.268433f
C5494 C9_P_btm.t444 VSS 0.242037f
C5495 C9_P_btm.t330 VSS 0.242037f
C5496 C9_P_btm.t230 VSS 0.242037f
C5497 C9_P_btm.t361 VSS 0.242037f
C5498 C9_P_btm.t251 VSS 0.268433f
C5499 C9_P_btm.n1061 VSS 0.101561f
C5500 C9_P_btm.t244 VSS 0.242037f
C5501 C9_P_btm.t372 VSS 0.268433f
C5502 C9_P_btm.t491 VSS 0.242037f
C5503 C9_P_btm.t343 VSS 0.242037f
C5504 C9_P_btm.t463 VSS 0.242037f
C5505 C9_P_btm.t69 VSS 0.242037f
C5506 C9_P_btm.t436 VSS 0.268433f
C5507 C9_P_btm.t114 VSS 0.268433f
C5508 C9_P_btm.t253 VSS 0.242037f
C5509 C9_P_btm.t133 VSS 0.242037f
C5510 C9_P_btm.t45 VSS 0.242037f
C5511 C9_P_btm.t164 VSS 0.242037f
C5512 C9_P_btm.t51 VSS 0.268433f
C5513 C9_P_btm.t239 VSS 0.242037f
C5514 C9_P_btm.t455 VSS 0.268433f
C5515 C9_P_btm.t61 VSS 0.242037f
C5516 C9_P_btm.t428 VSS 0.242037f
C5517 C9_P_btm.t32 VSS 0.242037f
C5518 C9_P_btm.t156 VSS 0.242037f
C5519 C9_P_btm.t288 VSS 0.268433f
C5520 C9_P_btm.t519 VSS 0.268433f
C5521 C9_P_btm.t314 VSS 0.242037f
C5522 C9_P_btm.t206 VSS 0.242037f
C5523 C9_P_btm.t113 VSS 0.242037f
C5524 C9_P_btm.t246 VSS 0.242037f
C5525 C9_P_btm.t129 VSS 0.268433f
C5526 C9_P_btm.t195 VSS 0.242037f
C5527 C9_P_btm.t502 VSS 0.268433f
C5528 C9_P_btm.t356 VSS 0.242037f
C5529 C9_P_btm.t219 VSS 0.242037f
C5530 C9_P_btm.t328 VSS 0.242037f
C5531 C9_P_btm.t441 VSS 0.242037f
C5532 C9_P_btm.t303 VSS 0.268433f
C5533 C9_P_btm.t528 VSS 0.268433f
C5534 C9_P_btm.t392 VSS 0.242037f
C5535 C9_P_btm.t282 VSS 0.242037f
C5536 C9_P_btm.t183 VSS 0.242037f
C5537 C9_P_btm.t309 VSS 0.242037f
C5538 C9_P_btm.t200 VSS 0.268433f
C5539 C9_P_btm.t263 VSS 0.242037f
C5540 C9_P_btm.t322 VSS 0.268433f
C5541 C9_P_btm.t437 VSS 0.242037f
C5542 C9_P_btm.t297 VSS 0.242037f
C5543 C9_P_btm.t413 VSS 0.242037f
C5544 C9_P_btm.t37 VSS 0.242037f
C5545 C9_P_btm.t383 VSS 0.268433f
C5546 C9_P_btm.t335 VSS 0.268433f
C5547 C9_P_btm.t482 VSS 0.242037f
C5548 C9_P_btm.t365 VSS 0.242037f
C5549 C9_P_btm.t526 VSS 0.242037f
C5550 C9_P_btm.t389 VSS 0.242037f
C5551 C9_P_btm.t279 VSS 0.268433f
C5552 C9_P_btm.t59 VSS 0.242037f
C5553 C9_P_btm.t409 VSS 0.268433f
C5554 C9_P_btm.t30 VSS 0.242037f
C5555 C9_P_btm.t378 VSS 0.242037f
C5556 C9_P_btm.t510 VSS 0.242037f
C5557 C9_P_btm.t107 VSS 0.242037f
C5558 C9_P_btm.t472 VSS 0.268433f
C5559 C9_P_btm.t420 VSS 0.268433f
C5560 C9_P_btm.t228 VSS 0.242037f
C5561 C9_P_btm.t446 VSS 0.242037f
C5562 C9_P_btm.t331 VSS 0.242037f
C5563 C9_P_btm.t481 VSS 0.242037f
C5564 C9_P_btm.t363 VSS 0.268433f
C5565 C9_P_btm.t145 VSS 0.242037f
C5566 C9_P_btm.t521 VSS 0.242037f
C5567 C9_P_btm.t500 VSS 0.242037f
C5568 C9_P_btm.t216 VSS 0.242037f
C5569 C9_P_btm.t47 VSS 0.268433f
C5570 C9_P_btm.t182 VSS 0.242037f
C5571 C9_P_btm.t72 VSS 0.242037f
C5572 C9_P_btm.t465 VSS 0.242037f
C5573 C9_P_btm.t98 VSS 0.242037f
C5574 C9_P_btm.t493 VSS 0.242037f
C5575 C9_P_btm.t155 VSS 0.242037f
C5576 C9_P_btm.t245 VSS 0.242037f
C5577 C9_P_btm.t403 VSS 0.242037f
C5578 C9_P_btm.t60 VSS 0.242037f
C5579 C9_P_btm.t453 VSS 0.242037f
C5580 C9_P_btm.t317 VSS 0.242037f
C5581 C9_P_btm.t464 VSS 0.242037f
C5582 C9_P_btm.t346 VSS 0.242037f
C5583 C9_P_btm.t212 VSS 0.242037f
C5584 C9_P_btm.t374 VSS 0.242037f
C5585 C9_P_btm.t265 VSS 0.242037f
C5586 C9_P_btm.t401 VSS 0.242037f
C5587 C9_P_btm.t286 VSS 0.242037f
C5588 C9_P_btm.t191 VSS 0.268433f
C5589 C9_P_btm.t220 VSS 0.268433f
C5590 C9_P_btm.t532 VSS 0.242037f
C5591 C9_P_btm.t134 VSS 0.242037f
C5592 C9_P_btm.t283 VSS 0.242037f
C5593 C9_P_btm.t184 VSS 0.242037f
C5594 C9_P_btm.t56 VSS 0.242037f
C5595 C9_P_btm.t202 VSS 0.242037f
C5596 C9_P_btm.t99 VSS 0.242037f
C5597 C9_P_btm.t495 VSS 0.242037f
C5598 C9_P_btm.t125 VSS 0.242037f
C5599 C9_P_btm.t70 VSS 0.242037f
C5600 C9_P_btm.t176 VSS 0.242037f
C5601 C9_P_btm.t35 VSS 0.242037f
C5602 C9_P_btm.t431 VSS 0.242037f
C5603 C9_P_btm.t247 VSS 0.242037f
C5604 C9_P_btm.t400 VSS 0.242037f
C5605 C9_P_btm.t38 VSS 0.242037f
C5606 C9_P_btm.t149 VSS 0.242037f
C5607 C9_P_btm.t489 VSS 0.242037f
C5608 C9_P_btm.t92 VSS 0.242037f
C5609 C9_P_btm.t222 VSS 0.242037f
C5610 C9_P_btm.t66 VSS 0.242037f
C5611 C9_P_btm.t180 VSS 0.242037f
C5612 C9_P_btm.t43 VSS 0.242037f
C5613 C9_P_btm.t161 VSS 0.242037f
C5614 C9_P_btm.t522 VSS 0.242037f
C5615 C9_P_btm.t110 VSS 0.242037f
C5616 C9_P_btm.t240 VSS 0.242037f
C5617 C9_P_btm.t333 VSS 0.242037f
C5618 C9_P_btm.t187 VSS 0.242037f
C5619 C9_P_btm.t311 VSS 0.242037f
C5620 C9_P_btm.t167 VSS 0.242037f
C5621 C9_P_btm.t534 VSS 0.242037f
C5622 C9_P_btm.t394 VSS 0.242037f
C5623 C9_P_btm.t267 VSS 0.242037f
C5624 C9_P_btm.t339 VSS 0.242037f
C5625 C9_P_btm.t456 VSS 0.242037f
C5626 C9_P_btm.t318 VSS 0.242037f
C5627 C9_P_btm.t429 VSS 0.242037f
C5628 C9_P_btm.t273 VSS 0.242037f
C5629 C9_P_btm.t405 VSS 0.242037f
C5630 C9_P_btm.t324 VSS 0.242037f
C5631 C9_P_btm.t370 VSS 0.242037f
C5632 C9_P_btm.t517 VSS 0.242037f
C5633 C9_P_btm.t121 VSS 0.242037f
C5634 C9_P_btm.t461 VSS 0.242037f
C5635 C9_P_btm.t65 VSS 0.242037f
C5636 C9_P_btm.t198 VSS 0.242037f
C5637 C9_P_btm.t41 VSS 0.242037f
C5638 C9_P_btm.t160 VSS 0.242037f
C5639 C9_P_btm.t25 VSS 0.242037f
C5640 C9_P_btm.t128 VSS 0.242037f
C5641 C9_P_btm.t238 VSS 0.242037f
C5642 C9_P_btm.t104 VSS 0.268433f
C5643 C9_P_btm.t115 VSS 0.268433f
C5644 C9_P_btm.t524 VSS 0.242037f
C5645 C9_P_btm.t81 VSS 0.242037f
C5646 C9_P_btm.t480 VSS 0.242037f
C5647 C9_P_btm.t227 VSS 0.242037f
C5648 C9_P_btm.t506 VSS 0.242037f
C5649 C9_P_btm.t165 VSS 0.242037f
C5650 C9_P_btm.t52 VSS 0.242037f
C5651 C9_P_btm.t416 VSS 0.242037f
C5652 C9_P_btm.t76 VSS 0.242037f
C5653 C9_P_btm.t470 VSS 0.242037f
C5654 C9_P_btm.t326 VSS 0.242037f
C5655 C9_P_btm.t476 VSS 0.242037f
C5656 C9_P_btm.t359 VSS 0.242037f
C5657 C9_P_btm.t226 VSS 0.242037f
C5658 C9_P_btm.t381 VSS 0.242037f
C5659 C9_P_btm.t277 VSS 0.242037f
C5660 C9_P_btm.t411 VSS 0.242037f
C5661 C9_P_btm.t295 VSS 0.242037f
C5662 C9_P_btm.t533 VSS 0.242037f
C5663 C9_P_btm.t347 VSS 0.242037f
C5664 C9_P_btm.t213 VSS 0.242037f
C5665 C9_P_btm.t268 VSS 0.242037f
C5666 C9_P_btm.t266 VSS 0.242037f
C5667 C9_P_btm.t143 VSS 0.242037f
C5668 C9_P_btm.t289 VSS 0.242037f
C5669 C9_P_btm.t193 VSS 0.242037f
C5670 C9_P_btm.t236 VSS 0.242037f
C5671 C9_P_btm.t208 VSS 0.242037f
C5672 C9_P_btm.t232 VSS 0.242037f
C5673 C9_P_btm.t507 VSS 0.242037f
C5674 C9_P_btm.t136 VSS 0.242037f
C5675 C9_P_btm.t94 VSS 0.242037f
C5676 C9_P_btm.t186 VSS 0.242037f
C5677 C9_P_btm.t100 VSS 0.242037f
C5678 C9_P_btm.t439 VSS 0.242037f
C5679 C9_P_btm.t106 VSS 0.242037f
C5680 C9_P_btm.t471 VSS 0.242037f
C5681 C9_P_btm.t355 VSS 0.242037f
C5682 C9_P_btm.t68 VSS 0.242037f
C5683 C9_P_btm.t462 VSS 0.242037f
C5684 C9_P_btm.t320 VSS 0.268433f
C5685 C9_P_btm.t146 VSS 0.242037f
C5686 C9_P_btm.t280 VSS 0.268433f
C5687 C9_P_btm.t417 VSS 0.242037f
C5688 C9_P_btm.t109 VSS 0.242037f
C5689 C9_P_btm.t341 VSS 0.242037f
C5690 C9_P_btm.t458 VSS 0.242037f
C5691 C9_P_btm.t88 VSS 0.242037f
C5692 C9_P_btm.t140 VSS 0.268433f
C5693 C9_P_btm.t509 VSS 0.242037f
C5694 C9_P_btm.t390 VSS 0.242037f
C5695 C9_P_btm.t205 VSS 0.242037f
C5696 C9_P_btm.t111 VSS 0.242037f
C5697 C9_P_btm.t474 VSS 0.268433f
C5698 C9_P_btm.t332 VSS 0.242037f
C5699 C9_P_btm.t385 VSS 0.268433f
C5700 C9_P_btm.t34 VSS 0.242037f
C5701 C9_P_btm.t130 VSS 0.242037f
C5702 C9_P_btm.t264 VSS 0.242037f
C5703 C9_P_btm.t373 VSS 0.242037f
C5704 C9_P_btm.t102 VSS 0.268433f
C5705 C9_P_btm.t259 VSS 0.268433f
C5706 C9_P_btm.t422 VSS 0.242037f
C5707 C9_P_btm.t310 VSS 0.242037f
C5708 C9_P_btm.t307 VSS 0.242037f
C5709 C9_P_btm.t199 VSS 0.242037f
C5710 C9_P_btm.t71 VSS 0.268433f
C5711 C9_P_btm.t440 VSS 0.242037f
C5712 C9_P_btm.t497 VSS 0.268433f
C5713 C9_P_btm.t124 VSS 0.242037f
C5714 C9_P_btm.t233 VSS 0.242037f
C5715 C9_P_btm.t196 VSS 0.242037f
C5716 C9_P_btm.t293 VSS 0.242037f
C5717 C9_P_btm.t432 VSS 0.268433f
C5718 C9_P_btm.t530 VSS 0.268433f
C5719 C9_P_btm.t132 VSS 0.242037f
C5720 C9_P_btm.t42 VSS 0.242037f
C5721 C9_P_btm.t475 VSS 0.242037f
C5722 C9_P_btm.t358 VSS 0.242037f
C5723 C9_P_btm.t225 VSS 0.268433f
C5724 C9_P_btm.t44 VSS 0.242037f
C5725 C9_P_btm.t90 VSS 0.268433f
C5726 C9_P_btm.t218 VSS 0.242037f
C5727 C9_P_btm.t329 VSS 0.242037f
C5728 C9_P_btm.t254 VSS 0.242037f
C5729 C9_P_btm.t211 VSS 0.242037f
C5730 C9_P_btm.t345 VSS 0.268433f
C5731 C9_P_btm.t190 VSS 0.268433f
C5732 C9_P_btm.t108 VSS 0.242037f
C5733 C9_P_btm.t442 VSS 0.242037f
C5734 C9_P_btm.t73 VSS 0.242037f
C5735 C9_P_btm.t468 VSS 0.242037f
C5736 C9_P_btm.t323 VSS 0.268433f
C5737 C9_P_btm.t153 VSS 0.242037f
C5738 C9_P_btm.t512 VSS 0.268433f
C5739 C9_P_btm.t379 VSS 0.242037f
C5740 C9_P_btm.t511 VSS 0.242037f
C5741 C9_P_btm.t315 VSS 0.242037f
C5742 C9_P_btm.t424 VSS 0.242037f
C5743 C9_P_btm.t514 VSS 0.268433f
C5744 C9_P_btm.t487 VSS 0.268433f
C5745 C9_P_btm.t352 VSS 0.242037f
C5746 C9_P_btm.t408 VSS 0.242037f
C5747 C9_P_btm.t516 VSS 0.242037f
C5748 C9_P_btm.t157 VSS 0.268433f
C5749 C9_P_btm.t119 VSS 0.268433f
C5750 C9_P_btm.t479 VSS 0.242037f
C5751 C9_P_btm.t362 VSS 0.242037f
C5752 C9_P_btm.t177 VSS 0.242037f
C5753 C9_P_btm.t62 VSS 0.242037f
C5754 C9_P_btm.t433 VSS 0.268433f
C5755 C9_P_btm.t499 VSS 0.242037f
C5756 C9_P_btm.t344 VSS 0.268433f
C5757 C9_P_btm.t490 VSS 0.242037f
C5758 C9_P_btm.t95 VSS 0.242037f
C5759 C9_P_btm.t256 VSS 0.242037f
C5760 C9_P_btm.t336 VSS 0.242037f
C5761 C9_P_btm.t101 VSS 0.268433f
C5762 C9_P_btm.t388 VSS 0.242037f
C5763 C9_P_btm.t278 VSS 0.242037f
C5764 C9_P_btm.t274 VSS 0.242037f
C5765 C9_P_btm.t173 VSS 0.242037f
C5766 C9_P_btm.t27 VSS 0.268433f
C5767 C9_P_btm.t22 VSS 0.279048f
C5768 C9_P_btm.n1870 VSS 0.101561f
C5769 C9_P_btm.t272 VSS 0.268433f
C5770 C9_P_btm.t404 VSS 0.242037f
C5771 C9_P_btm.t260 VSS 0.242037f
C5772 C9_P_btm.t398 VSS 0.242037f
C5773 C9_P_btm.t215 VSS 0.242037f
C5774 C9_P_btm.t354 VSS 0.268433f
C5775 C9_P_btm.t23 VSS 0.268885f
C5776 C9_P_btm.n1886 VSS 0.135994f
C5777 C9_N_btm.n0 VSS 0.189503f
C5778 C9_N_btm.n1 VSS 0.183283f
C5779 C9_N_btm.n2 VSS 0.576045f
C5780 C9_N_btm.n3 VSS 0.183283f
C5781 C9_N_btm.n4 VSS 0.295062f
C5782 C9_N_btm.n5 VSS 0.183283f
C5783 C9_N_btm.n6 VSS 0.467875f
C5784 C9_N_btm.n7 VSS 0.278269f
C5785 C9_N_btm.n8 VSS 0.271861f
C5786 C9_N_btm.n9 VSS 0.442686f
C5787 C9_N_btm.n10 VSS 0.264268f
C5788 C9_N_btm.t4 VSS 0.414646f
C5789 C9_N_btm.n11 VSS 0.33082f
C5790 C9_N_btm.n12 VSS 0.281048f
C5791 C9_N_btm.n13 VSS 0.274973f
C5792 C9_N_btm.n14 VSS 0.447509f
C5793 C9_N_btm.n15 VSS 1.104f
C5794 C9_N_btm.t530 VSS 0.279047f
C5795 C9_N_btm.t532 VSS 0.279047f
C5796 C9_N_btm.t533 VSS 0.279047f
C5797 C9_N_btm.t536 VSS 0.279047f
C5798 C9_N_btm.t91 VSS 0.268432f
C5799 C9_N_btm.t526 VSS 0.279047f
C5800 C9_N_btm.t264 VSS 0.268432f
C5801 C9_N_btm.t372 VSS 0.268432f
C5802 C9_N_btm.t51 VSS 0.268432f
C5803 C9_N_btm.t94 VSS 0.242036f
C5804 C9_N_btm.t331 VSS 0.242036f
C5805 C9_N_btm.t440 VSS 0.242036f
C5806 C9_N_btm.t476 VSS 0.268432f
C5807 C9_N_btm.t488 VSS 0.268432f
C5808 C9_N_btm.t211 VSS 0.242036f
C5809 C9_N_btm.t508 VSS 0.242036f
C5810 C9_N_btm.t364 VSS 0.242036f
C5811 C9_N_btm.t116 VSS 0.268432f
C5812 C9_N_btm.t419 VSS 0.268432f
C5813 C9_N_btm.t319 VSS 0.242036f
C5814 C9_N_btm.t170 VSS 0.242036f
C5815 C9_N_btm.t274 VSS 0.242036f
C5816 C9_N_btm.t177 VSS 0.268432f
C5817 C9_N_btm.t335 VSS 0.268432f
C5818 C9_N_btm.t426 VSS 0.242036f
C5819 C9_N_btm.t74 VSS 0.242036f
C5820 C9_N_btm.t517 VSS 0.242036f
C5821 C9_N_btm.t337 VSS 0.268432f
C5822 C9_N_btm.t43 VSS 0.268432f
C5823 C9_N_btm.t128 VSS 0.268432f
C5824 C9_N_btm.t192 VSS 0.268432f
C5825 C9_N_btm.t97 VSS 0.242036f
C5826 C9_N_btm.t225 VSS 0.242036f
C5827 C9_N_btm.t333 VSS 0.242036f
C5828 C9_N_btm.t436 VSS 0.268432f
C5829 C9_N_btm.t487 VSS 0.268432f
C5830 C9_N_btm.t414 VSS 0.242036f
C5831 C9_N_btm.t50 VSS 0.242036f
C5832 C9_N_btm.t108 VSS 0.242036f
C5833 C9_N_btm.t22 VSS 0.268432f
C5834 C9_N_btm.t48 VSS 0.268432f
C5835 C9_N_btm.t484 VSS 0.242036f
C5836 C9_N_btm.t79 VSS 0.242036f
C5837 C9_N_btm.t197 VSS 0.242036f
C5838 C9_N_btm.t76 VSS 0.268432f
C5839 C9_N_btm.t137 VSS 0.268432f
C5840 C9_N_btm.t47 VSS 0.242036f
C5841 C9_N_btm.t175 VSS 0.242036f
C5842 C9_N_btm.t278 VSS 0.242036f
C5843 C9_N_btm.t527 VSS 0.279047f
C5844 C9_N_btm.t171 VSS 0.268432f
C5845 C9_N_btm.t534 VSS 0.279047f
C5846 C9_N_btm.t525 VSS 0.279047f
C5847 C9_N_btm.t535 VSS 0.279047f
C5848 C9_N_btm.t528 VSS 0.279047f
C5849 C9_N_btm.t227 VSS 0.268432f
C5850 C9_N_btm.t135 VSS 0.242036f
C5851 C9_N_btm.t518 VSS 0.242036f
C5852 C9_N_btm.t367 VSS 0.242036f
C5853 C9_N_btm.t531 VSS 0.279047f
C5854 C9_N_btm.n333 VSS 0.10156f
C5855 C9_N_btm.t397 VSS 0.268432f
C5856 C9_N_btm.t64 VSS 0.242036f
C5857 C9_N_btm.t431 VSS 0.242036f
C5858 C9_N_btm.t318 VSS 0.242036f
C5859 C9_N_btm.t452 VSS 0.242036f
C5860 C9_N_btm.t346 VSS 0.268432f
C5861 C9_N_btm.n348 VSS 0.10156f
C5862 C9_N_btm.t275 VSS 0.242036f
C5863 C9_N_btm.t215 VSS 0.268432f
C5864 C9_N_btm.t326 VSS 0.242036f
C5865 C9_N_btm.t188 VSS 0.242036f
C5866 C9_N_btm.t150 VSS 0.242036f
C5867 C9_N_btm.t412 VSS 0.242036f
C5868 C9_N_btm.t270 VSS 0.268432f
C5869 C9_N_btm.t85 VSS 0.268432f
C5870 C9_N_btm.t234 VSS 0.242036f
C5871 C9_N_btm.t243 VSS 0.242036f
C5872 C9_N_btm.t400 VSS 0.242036f
C5873 C9_N_btm.t144 VSS 0.242036f
C5874 C9_N_btm.t28 VSS 0.268432f
C5875 C9_N_btm.t519 VSS 0.242036f
C5876 C9_N_btm.t127 VSS 0.268432f
C5877 C9_N_btm.t314 VSS 0.242036f
C5878 C9_N_btm.t95 VSS 0.242036f
C5879 C9_N_btm.t221 VSS 0.242036f
C5880 C9_N_btm.t330 VSS 0.242036f
C5881 C9_N_btm.t511 VSS 0.268432f
C5882 C9_N_btm.t361 VSS 0.268432f
C5883 C9_N_btm.t149 VSS 0.242036f
C5884 C9_N_btm.t32 VSS 0.242036f
C5885 C9_N_btm.t446 VSS 0.242036f
C5886 C9_N_btm.t240 VSS 0.242036f
C5887 C9_N_btm.t470 VSS 0.268432f
C5888 C9_N_btm.t104 VSS 0.242036f
C5889 C9_N_btm.t349 VSS 0.268432f
C5890 C9_N_btm.t457 VSS 0.242036f
C5891 C9_N_btm.t321 VSS 0.242036f
C5892 C9_N_btm.t434 VSS 0.242036f
C5893 C9_N_btm.t14 VSS 0.242036f
C5894 C9_N_btm.t402 VSS 0.268432f
C5895 C9_N_btm.t450 VSS 0.268432f
C5896 C9_N_btm.t65 VSS 0.242036f
C5897 C9_N_btm.t475 VSS 0.242036f
C5898 C9_N_btm.t368 VSS 0.242036f
C5899 C9_N_btm.t498 VSS 0.242036f
C5900 C9_N_btm.t389 VSS 0.268432f
C5901 C9_N_btm.t53 VSS 0.242036f
C5902 C9_N_btm.t260 VSS 0.268432f
C5903 C9_N_btm.t375 VSS 0.242036f
C5904 C9_N_btm.t235 VSS 0.242036f
C5905 C9_N_btm.t353 VSS 0.242036f
C5906 C9_N_btm.t460 VSS 0.242036f
C5907 C9_N_btm.t323 VSS 0.268432f
C5908 C9_N_btm.t369 VSS 0.268432f
C5909 C9_N_btm.t506 VSS 0.242036f
C5910 C9_N_btm.t392 VSS 0.242036f
C5911 C9_N_btm.t279 VSS 0.242036f
C5912 C9_N_btm.t425 VSS 0.242036f
C5913 C9_N_btm.t311 VSS 0.268432f
C5914 C9_N_btm.t500 VSS 0.242036f
C5915 C9_N_btm.t183 VSS 0.268432f
C5916 C9_N_btm.t295 VSS 0.242036f
C5917 C9_N_btm.t151 VSS 0.242036f
C5918 C9_N_btm.t265 VSS 0.242036f
C5919 C9_N_btm.t378 VSS 0.242036f
C5920 C9_N_btm.t244 VSS 0.268432f
C5921 C9_N_btm.t101 VSS 0.268432f
C5922 C9_N_btm.t282 VSS 0.268432f
C5923 C9_N_btm.t428 VSS 0.242036f
C5924 C9_N_btm.t317 VSS 0.242036f
C5925 C9_N_btm.t199 VSS 0.242036f
C5926 C9_N_btm.t343 VSS 0.242036f
C5927 C9_N_btm.t229 VSS 0.268432f
C5928 C9_N_btm.t169 VSS 0.242036f
C5929 C9_N_btm.t16 VSS 0.242036f
C5930 C9_N_btm.t134 VSS 0.242036f
C5931 C9_N_btm.t514 VSS 0.242036f
C5932 C9_N_btm.t158 VSS 0.268432f
C5933 C9_N_btm.t302 VSS 0.242036f
C5934 C9_N_btm.t507 VSS 0.242036f
C5935 C9_N_btm.t516 VSS 0.242036f
C5936 C9_N_btm.t213 VSS 0.242036f
C5937 C9_N_btm.t88 VSS 0.242036f
C5938 C9_N_btm.t524 VSS 0.242036f
C5939 C9_N_btm.t289 VSS 0.242036f
C5940 C9_N_btm.t398 VSS 0.242036f
C5941 C9_N_btm.t181 VSS 0.242036f
C5942 C9_N_btm.t109 VSS 0.242036f
C5943 C9_N_btm.t443 VSS 0.242036f
C5944 C9_N_btm.t62 VSS 0.242036f
C5945 C9_N_btm.t474 VSS 0.242036f
C5946 C9_N_btm.t340 VSS 0.242036f
C5947 C9_N_btm.t497 VSS 0.242036f
C5948 C9_N_btm.t388 VSS 0.242036f
C5949 C9_N_btm.t435 VSS 0.242036f
C5950 C9_N_btm.t421 VSS 0.242036f
C5951 C9_N_btm.t309 VSS 0.268432f
C5952 C9_N_btm.t223 VSS 0.268432f
C5953 C9_N_btm.t383 VSS 0.242036f
C5954 C9_N_btm.t499 VSS 0.242036f
C5955 C9_N_btm.t411 VSS 0.242036f
C5956 C9_N_btm.t304 VSS 0.242036f
C5957 C9_N_btm.t161 VSS 0.242036f
C5958 C9_N_btm.t325 VSS 0.242036f
C5959 C9_N_btm.t214 VSS 0.242036f
C5960 C9_N_btm.t90 VSS 0.242036f
C5961 C9_N_btm.t241 VSS 0.242036f
C5962 C9_N_btm.t356 VSS 0.242036f
C5963 C9_N_btm.t291 VSS 0.242036f
C5964 C9_N_btm.t148 VSS 0.242036f
C5965 C9_N_btm.t31 VSS 0.242036f
C5966 C9_N_btm.t247 VSS 0.242036f
C5967 C9_N_btm.t303 VSS 0.242036f
C5968 C9_N_btm.t410 VSS 0.242036f
C5969 C9_N_btm.t24 VSS 0.242036f
C5970 C9_N_btm.t382 VSS 0.242036f
C5971 C9_N_btm.t486 VSS 0.242036f
C5972 C9_N_btm.t105 VSS 0.242036f
C5973 C9_N_btm.t466 VSS 0.242036f
C5974 C9_N_btm.t54 VSS 0.242036f
C5975 C9_N_btm.t441 VSS 0.242036f
C5976 C9_N_btm.t503 VSS 0.242036f
C5977 C9_N_btm.t143 VSS 0.242036f
C5978 C9_N_btm.t496 VSS 0.242036f
C5979 C9_N_btm.t236 VSS 0.242036f
C5980 C9_N_btm.t233 VSS 0.242036f
C5981 C9_N_btm.t61 VSS 0.242036f
C5982 C9_N_btm.t207 VSS 0.242036f
C5983 C9_N_btm.t37 VSS 0.242036f
C5984 C9_N_btm.t154 VSS 0.242036f
C5985 C9_N_btm.t297 VSS 0.242036f
C5986 C9_N_btm.t126 VSS 0.242036f
C5987 C9_N_btm.t253 VSS 0.242036f
C5988 C9_N_btm.t359 VSS 0.242036f
C5989 C9_N_btm.t220 VSS 0.242036f
C5990 C9_N_btm.t329 VSS 0.242036f
C5991 C9_N_btm.t166 VSS 0.242036f
C5992 C9_N_btm.t307 VSS 0.242036f
C5993 C9_N_btm.t416 VSS 0.242036f
C5994 C9_N_btm.t269 VSS 0.242036f
C5995 C9_N_btm.t406 VSS 0.242036f
C5996 C9_N_btm.t18 VSS 0.242036f
C5997 C9_N_btm.t362 VSS 0.242036f
C5998 C9_N_btm.t464 VSS 0.242036f
C5999 C9_N_btm.t78 VSS 0.242036f
C6000 C9_N_btm.t439 VSS 0.242036f
C6001 C9_N_btm.t120 VSS 0.242036f
C6002 C9_N_btm.t418 VSS 0.242036f
C6003 C9_N_btm.t254 VSS 0.242036f
C6004 C9_N_btm.t117 VSS 0.242036f
C6005 C9_N_btm.t492 VSS 0.268432f
C6006 C9_N_btm.t224 VSS 0.268432f
C6007 C9_N_btm.t133 VSS 0.268432f
C6008 C9_N_btm.t100 VSS 0.268432f
C6009 C9_N_btm.t467 VSS 0.242036f
C6010 C9_N_btm.t427 VSS 0.242036f
C6011 C9_N_btm.t267 VSS 0.242036f
C6012 C9_N_btm.t156 VSS 0.242036f
C6013 C9_N_btm.t26 VSS 0.242036f
C6014 C9_N_btm.t96 VSS 0.242036f
C6015 C9_N_btm.t288 VSS 0.242036f
C6016 C9_N_btm.t71 VSS 0.242036f
C6017 C9_N_btm.t513 VSS 0.242036f
C6018 C9_N_btm.t42 VSS 0.242036f
C6019 C9_N_btm.t168 VSS 0.242036f
C6020 C9_N_btm.t273 VSS 0.242036f
C6021 C9_N_btm.t102 VSS 0.242036f
C6022 C9_N_btm.t512 VSS 0.242036f
C6023 C9_N_btm.t365 VSS 0.242036f
C6024 C9_N_btm.t521 VSS 0.242036f
C6025 C9_N_btm.t338 VSS 0.242036f
C6026 C9_N_btm.t176 VSS 0.242036f
C6027 C9_N_btm.t280 VSS 0.242036f
C6028 C9_N_btm.t424 VSS 0.242036f
C6029 C9_N_btm.t256 VSS 0.242036f
C6030 C9_N_btm.t371 VSS 0.242036f
C6031 C9_N_btm.t477 VSS 0.242036f
C6032 C9_N_btm.t347 VSS 0.242036f
C6033 C9_N_btm.t455 VSS 0.242036f
C6034 C9_N_btm.t292 VSS 0.242036f
C6035 C9_N_btm.t432 VSS 0.242036f
C6036 C9_N_btm.t262 VSS 0.242036f
C6037 C9_N_btm.t393 VSS 0.242036f
C6038 C9_N_btm.t344 VSS 0.242036f
C6039 C9_N_btm.t124 VSS 0.242036f
C6040 C9_N_btm.t478 VSS 0.242036f
C6041 C9_N_btm.t69 VSS 0.242036f
C6042 C9_N_btm.t218 VSS 0.242036f
C6043 C9_N_btm.t40 VSS 0.242036f
C6044 C9_N_btm.t164 VSS 0.242036f
C6045 C9_N_btm.t13 VSS 0.242036f
C6046 C9_N_btm.t131 VSS 0.242036f
C6047 C9_N_btm.t249 VSS 0.242036f
C6048 C9_N_btm.t350 VSS 0.268432f
C6049 C9_N_btm.t208 VSS 0.242036f
C6050 C9_N_btm.t373 VSS 0.242036f
C6051 C9_N_btm.t257 VSS 0.242036f
C6052 C9_N_btm.t395 VSS 0.242036f
C6053 C9_N_btm.t284 VSS 0.242036f
C6054 C9_N_btm.t178 VSS 0.242036f
C6055 C9_N_btm.t342 VSS 0.242036f
C6056 C9_N_btm.t200 VSS 0.242036f
C6057 C9_N_btm.t81 VSS 0.242036f
C6058 C9_N_btm.t520 VSS 0.242036f
C6059 C9_N_btm.t106 VSS 0.242036f
C6060 C9_N_btm.t276 VSS 0.242036f
C6061 C9_N_btm.t172 VSS 0.242036f
C6062 C9_N_btm.t46 VSS 0.242036f
C6063 C9_N_btm.t193 VSS 0.268432f
C6064 C9_N_btm.t272 VSS 0.242036f
C6065 C9_N_btm.t385 VSS 0.242036f
C6066 C9_N_btm.t300 VSS 0.242036f
C6067 C9_N_btm.t407 VSS 0.242036f
C6068 C9_N_btm.t20 VSS 0.242036f
C6069 C9_N_btm.t380 VSS 0.242036f
C6070 C9_N_btm.t485 VSS 0.242036f
C6071 C9_N_btm.t103 VSS 0.242036f
C6072 C9_N_btm.t463 VSS 0.242036f
C6073 C9_N_btm.t52 VSS 0.242036f
C6074 C9_N_btm.t438 VSS 0.242036f
C6075 C9_N_btm.t113 VSS 0.242036f
C6076 C9_N_btm.t140 VSS 0.242036f
C6077 C9_N_btm.t493 VSS 0.242036f
C6078 C9_N_btm.t115 VSS 0.242036f
C6079 C9_N_btm.t232 VSS 0.242036f
C6080 C9_N_btm.t502 VSS 0.242036f
C6081 C9_N_btm.t205 VSS 0.242036f
C6082 C9_N_btm.t34 VSS 0.242036f
C6083 C9_N_btm.t152 VSS 0.242036f
C6084 C9_N_btm.t294 VSS 0.242036f
C6085 C9_N_btm.t122 VSS 0.242036f
C6086 C9_N_btm.t250 VSS 0.242036f
C6087 C9_N_btm.t358 VSS 0.242036f
C6088 C9_N_btm.t216 VSS 0.242036f
C6089 C9_N_btm.t327 VSS 0.242036f
C6090 C9_N_btm.t163 VSS 0.242036f
C6091 C9_N_btm.t305 VSS 0.242036f
C6092 C9_N_btm.t415 VSS 0.242036f
C6093 C9_N_btm.t266 VSS 0.242036f
C6094 C9_N_btm.t404 VSS 0.242036f
C6095 C9_N_btm.t515 VSS 0.242036f
C6096 C9_N_btm.t360 VSS 0.242036f
C6097 C9_N_btm.t462 VSS 0.242036f
C6098 C9_N_btm.t77 VSS 0.242036f
C6099 C9_N_btm.t437 VSS 0.242036f
C6100 C9_N_btm.t56 VSS 0.242036f
C6101 C9_N_btm.t417 VSS 0.242036f
C6102 C9_N_btm.t121 VSS 0.242036f
C6103 C9_N_btm.t111 VSS 0.242036f
C6104 C9_N_btm.t489 VSS 0.268432f
C6105 C9_N_btm.t155 VSS 0.268432f
C6106 C9_N_btm.t299 VSS 0.242036f
C6107 C9_N_btm.t186 VSS 0.242036f
C6108 C9_N_btm.t63 VSS 0.242036f
C6109 C9_N_btm.t209 VSS 0.242036f
C6110 C9_N_btm.t84 VSS 0.242036f
C6111 C9_N_btm.t258 VSS 0.242036f
C6112 C9_N_btm.t239 VSS 0.242036f
C6113 C9_N_btm.t405 VSS 0.242036f
C6114 C9_N_btm.t179 VSS 0.242036f
C6115 C9_N_btm.t55 VSS 0.242036f
C6116 C9_N_btm.t442 VSS 0.242036f
C6117 C9_N_btm.t59 VSS 0.242036f
C6118 C9_N_btm.t472 VSS 0.242036f
C6119 C9_N_btm.t339 VSS 0.242036f
C6120 C9_N_btm.t494 VSS 0.242036f
C6121 C9_N_btm.t386 VSS 0.242036f
C6122 C9_N_btm.t483 VSS 0.242036f
C6123 C9_N_btm.t420 VSS 0.242036f
C6124 C9_N_btm.t308 VSS 0.242036f
C6125 C9_N_btm.t465 VSS 0.242036f
C6126 C9_N_btm.t332 VSS 0.242036f
C6127 C9_N_btm.t222 VSS 0.242036f
C6128 C9_N_btm.t381 VSS 0.242036f
C6129 C9_N_btm.t355 VSS 0.242036f
C6130 C9_N_btm.t409 VSS 0.242036f
C6131 C9_N_btm.t301 VSS 0.242036f
C6132 C9_N_btm.t160 VSS 0.242036f
C6133 C9_N_btm.t324 VSS 0.242036f
C6134 C9_N_btm.t212 VSS 0.242036f
C6135 C9_N_btm.t87 VSS 0.242036f
C6136 C9_N_btm.t238 VSS 0.242036f
C6137 C9_N_btm.t246 VSS 0.242036f
C6138 C9_N_btm.t287 VSS 0.242036f
C6139 C9_N_btm.t147 VSS 0.242036f
C6140 C9_N_btm.t30 VSS 0.242036f
C6141 C9_N_btm.t202 VSS 0.242036f
C6142 C9_N_btm.t112 VSS 0.242036f
C6143 C9_N_btm.t468 VSS 0.242036f
C6144 C9_N_btm.t136 VSS 0.242036f
C6145 C9_N_btm.t21 VSS 0.242036f
C6146 C9_N_btm.t408 VSS 0.268432f
C6147 C9_N_btm.t363 VSS 0.242036f
C6148 C9_N_btm.t194 VSS 0.268432f
C6149 C9_N_btm.t334 VSS 0.242036f
C6150 C9_N_btm.t444 VSS 0.242036f
C6151 C9_N_btm.t387 VSS 0.242036f
C6152 C9_N_btm.t495 VSS 0.242036f
C6153 C9_N_btm.t118 VSS 0.242036f
C6154 C9_N_btm.t473 VSS 0.242036f
C6155 C9_N_btm.t60 VSS 0.242036f
C6156 C9_N_btm.t206 VSS 0.242036f
C6157 C9_N_btm.t36 VSS 0.242036f
C6158 C9_N_btm.t153 VSS 0.242036f
C6159 C9_N_btm.t298 VSS 0.242036f
C6160 C9_N_btm.t125 VSS 0.242036f
C6161 C9_N_btm.t251 VSS 0.242036f
C6162 C9_N_btm.t70 VSS 0.242036f
C6163 C9_N_btm.t219 VSS 0.242036f
C6164 C9_N_btm.t328 VSS 0.242036f
C6165 C9_N_btm.t165 VSS 0.242036f
C6166 C9_N_btm.t306 VSS 0.242036f
C6167 C9_N_btm.t132 VSS 0.242036f
C6168 C9_N_btm.t510 VSS 0.242036f
C6169 C9_N_btm.t384 VSS 0.242036f
C6170 C9_N_btm.t226 VSS 0.242036f
C6171 C9_N_btm.t336 VSS 0.242036f
C6172 C9_N_btm.t445 VSS 0.242036f
C6173 C9_N_btm.t310 VSS 0.242036f
C6174 C9_N_btm.t423 VSS 0.242036f
C6175 C9_N_btm.t523 VSS 0.242036f
C6176 C9_N_btm.t390 VSS 0.242036f
C6177 C9_N_btm.t187 VSS 0.242036f
C6178 C9_N_btm.t366 VSS 0.242036f
C6179 C9_N_btm.t490 VSS 0.242036f
C6180 C9_N_btm.t83 VSS 0.242036f
C6181 C9_N_btm.t448 VSS 0.242036f
C6182 C9_N_btm.t35 VSS 0.242036f
C6183 C9_N_btm.t184 VSS 0.242036f
C6184 C9_N_btm.t354 VSS 0.242036f
C6185 C9_N_btm.t123 VSS 0.242036f
C6186 C9_N_btm.t19 VSS 0.242036f
C6187 C9_N_btm.t93 VSS 0.242036f
C6188 C9_N_btm.t217 VSS 0.242036f
C6189 C9_N_btm.t67 VSS 0.268432f
C6190 C9_N_btm.t23 VSS 0.268432f
C6191 C9_N_btm.t173 VSS 0.242036f
C6192 C9_N_btm.t45 VSS 0.242036f
C6193 C9_N_btm.t461 VSS 0.242036f
C6194 C9_N_btm.t73 VSS 0.242036f
C6195 C9_N_btm.t480 VSS 0.242036f
C6196 C9_N_btm.t130 VSS 0.242036f
C6197 C9_N_btm.t58 VSS 0.242036f
C6198 C9_N_btm.t399 VSS 0.242036f
C6199 C9_N_btm.t39 VSS 0.242036f
C6200 C9_N_btm.t453 VSS 0.242036f
C6201 C9_N_btm.t320 VSS 0.242036f
C6202 C9_N_btm.t459 VSS 0.242036f
C6203 C9_N_btm.t351 VSS 0.242036f
C6204 C9_N_btm.t210 VSS 0.242036f
C6205 C9_N_btm.t374 VSS 0.242036f
C6206 C9_N_btm.t259 VSS 0.242036f
C6207 C9_N_btm.t396 VSS 0.242036f
C6208 C9_N_btm.t285 VSS 0.242036f
C6209 C9_N_btm.t180 VSS 0.242036f
C6210 C9_N_btm.t345 VSS 0.242036f
C6211 C9_N_btm.t201 VSS 0.242036f
C6212 C9_N_btm.t82 VSS 0.242036f
C6213 C9_N_btm.t522 VSS 0.242036f
C6214 C9_N_btm.t107 VSS 0.242036f
C6215 C9_N_btm.t277 VSS 0.242036f
C6216 C9_N_btm.t174 VSS 0.242036f
C6217 C9_N_btm.t49 VSS 0.242036f
C6218 C9_N_btm.t195 VSS 0.242036f
C6219 C9_N_btm.t75 VSS 0.242036f
C6220 C9_N_btm.t482 VSS 0.242036f
C6221 C9_N_btm.t99 VSS 0.242036f
C6222 C9_N_btm.t505 VSS 0.242036f
C6223 C9_N_btm.t162 VSS 0.242036f
C6224 C9_N_btm.t504 VSS 0.242036f
C6225 C9_N_btm.t433 VSS 0.242036f
C6226 C9_N_btm.t68 VSS 0.242036f
C6227 C9_N_btm.t456 VSS 0.242036f
C6228 C9_N_btm.t348 VSS 0.242036f
C6229 C9_N_btm.t255 VSS 0.242036f
C6230 C9_N_btm.t139 VSS 0.242036f
C6231 C9_N_btm.t57 VSS 0.268432f
C6232 C9_N_btm.t471 VSS 0.242036f
C6233 C9_N_btm.t80 VSS 0.268432f
C6234 C9_N_btm.t228 VSS 0.242036f
C6235 C9_N_btm.t341 VSS 0.242036f
C6236 C9_N_btm.t469 VSS 0.242036f
C6237 C9_N_btm.t119 VSS 0.242036f
C6238 C9_N_btm.t204 VSS 0.242036f
C6239 C9_N_btm.t159 VSS 0.268432f
C6240 C9_N_btm.t167 VSS 0.242036f
C6241 C9_N_btm.t429 VSS 0.242036f
C6242 C9_N_btm.t145 VSS 0.242036f
C6243 C9_N_btm.t29 VSS 0.242036f
C6244 C9_N_btm.t422 VSS 0.268432f
C6245 C9_N_btm.t312 VSS 0.242036f
C6246 C9_N_btm.t491 VSS 0.268432f
C6247 C9_N_btm.t114 VSS 0.242036f
C6248 C9_N_btm.t231 VSS 0.242036f
C6249 C9_N_btm.t248 VSS 0.242036f
C6250 C9_N_btm.t142 VSS 0.242036f
C6251 C9_N_btm.t283 VSS 0.268432f
C6252 C9_N_btm.t245 VSS 0.268432f
C6253 C9_N_btm.t92 VSS 0.242036f
C6254 C9_N_btm.t189 VSS 0.242036f
C6255 C9_N_btm.t38 VSS 0.242036f
C6256 C9_N_btm.t449 VSS 0.242036f
C6257 C9_N_btm.t315 VSS 0.268432f
C6258 C9_N_btm.t203 VSS 0.242036f
C6259 C9_N_btm.t391 VSS 0.268432f
C6260 C9_N_btm.t379 VSS 0.242036f
C6261 C9_N_btm.t501 VSS 0.242036f
C6262 C9_N_btm.t110 VSS 0.242036f
C6263 C9_N_btm.t230 VSS 0.242036f
C6264 C9_N_btm.t370 VSS 0.268432f
C6265 C9_N_btm.t17 VSS 0.268432f
C6266 C9_N_btm.t403 VSS 0.242036f
C6267 C9_N_btm.t296 VSS 0.242036f
C6268 C9_N_btm.t394 VSS 0.242036f
C6269 C9_N_btm.t281 VSS 0.242036f
C6270 C9_N_btm.t141 VSS 0.268432f
C6271 C9_N_btm.t86 VSS 0.242036f
C6272 C9_N_btm.t286 VSS 0.268432f
C6273 C9_N_btm.t430 VSS 0.242036f
C6274 C9_N_btm.t146 VSS 0.242036f
C6275 C9_N_btm.t198 VSS 0.242036f
C6276 C9_N_btm.t316 VSS 0.242036f
C6277 C9_N_btm.t451 VSS 0.268432f
C6278 C9_N_btm.t98 VSS 0.268432f
C6279 C9_N_btm.t481 VSS 0.242036f
C6280 C9_N_btm.t377 VSS 0.242036f
C6281 C9_N_btm.t293 VSS 0.242036f
C6282 C9_N_btm.t182 VSS 0.242036f
C6283 C9_N_btm.t33 VSS 0.268432f
C6284 C9_N_btm.t190 VSS 0.242036f
C6285 C9_N_btm.t252 VSS 0.268432f
C6286 C9_N_btm.t261 VSS 0.242036f
C6287 C9_N_btm.t376 VSS 0.242036f
C6288 C9_N_btm.t27 VSS 0.242036f
C6289 C9_N_btm.t89 VSS 0.242036f
C6290 C9_N_btm.t237 VSS 0.268432f
C6291 C9_N_btm.t322 VSS 0.268432f
C6292 C9_N_btm.t15 VSS 0.242036f
C6293 C9_N_btm.t413 VSS 0.242036f
C6294 C9_N_btm.t25 VSS 0.242036f
C6295 C9_N_btm.t138 VSS 0.268432f
C6296 C9_N_btm.t191 VSS 0.268432f
C6297 C9_N_btm.t44 VSS 0.242036f
C6298 C9_N_btm.t458 VSS 0.242036f
C6299 C9_N_btm.t509 VSS 0.242036f
C6300 C9_N_btm.t66 VSS 0.242036f
C6301 C9_N_btm.t454 VSS 0.268432f
C6302 C9_N_btm.t401 VSS 0.242036f
C6303 C9_N_btm.t263 VSS 0.268432f
C6304 C9_N_btm.t157 VSS 0.242036f
C6305 C9_N_btm.t268 VSS 0.242036f
C6306 C9_N_btm.t290 VSS 0.242036f
C6307 C9_N_btm.t185 VSS 0.242036f
C6308 C9_N_btm.t271 VSS 0.268432f
C6309 C9_N_btm.t129 VSS 0.242036f
C6310 C9_N_btm.t41 VSS 0.242036f
C6311 C9_N_btm.t72 VSS 0.242036f
C6312 C9_N_btm.t479 VSS 0.242036f
C6313 C9_N_btm.t352 VSS 0.268432f
C6314 C9_N_btm.n1870 VSS 0.10156f
C6315 C9_N_btm.t242 VSS 0.242036f
C6316 C9_N_btm.t357 VSS 0.242036f
C6317 C9_N_btm.t196 VSS 0.242036f
C6318 C9_N_btm.t313 VSS 0.242036f
C6319 C9_N_btm.t447 VSS 0.268432f
C6320 C9_N_btm.t529 VSS 0.268883f
C6321 C9_N_btm.n1886 VSS 0.136138f
C6322 C8_P_btm.n0 VSS 0.214011f
C6323 C8_P_btm.n1 VSS 0.220788f
C6324 C8_P_btm.n2 VSS 0.853963f
C6325 C8_P_btm.n3 VSS 0.399375f
C6326 C8_P_btm.n4 VSS 0.566192f
C6327 C8_P_btm.n5 VSS 0.402318f
C6328 C8_P_btm.n6 VSS 0.437264f
C6329 C8_P_btm.n8 VSS 1.26048f
C6330 C8_P_btm.t12 VSS 0.325831f
C6331 C8_P_btm.n10 VSS 0.102832f
C6332 C8_P_btm.t17 VSS 0.325831f
C6333 C8_P_btm.n11 VSS 0.102832f
C6334 C8_P_btm.t8 VSS 0.325831f
C6335 C8_P_btm.n12 VSS 0.102832f
C6336 C8_P_btm.t95 VSS 0.313436f
C6337 C8_P_btm.t32 VSS 0.313436f
C6338 C8_P_btm.t127 VSS 0.313436f
C6339 C8_P_btm.t154 VSS 0.282615f
C6340 C8_P_btm.t74 VSS 0.282615f
C6341 C8_P_btm.t71 VSS 0.313436f
C6342 C8_P_btm.t170 VSS 0.313436f
C6343 C8_P_btm.t200 VSS 0.282615f
C6344 C8_P_btm.t175 VSS 0.282615f
C6345 C8_P_btm.t122 VSS 0.313436f
C6346 C8_P_btm.t242 VSS 0.282615f
C6347 C8_P_btm.t153 VSS 0.282615f
C6348 C8_P_btm.t214 VSS 0.282615f
C6349 C8_P_btm.t142 VSS 0.282615f
C6350 C8_P_btm.t202 VSS 0.313436f
C6351 C8_P_btm.t150 VSS 0.313436f
C6352 C8_P_btm.t104 VSS 0.313436f
C6353 C8_P_btm.t84 VSS 0.313436f
C6354 C8_P_btm.t110 VSS 0.313436f
C6355 C8_P_btm.t109 VSS 0.282615f
C6356 C8_P_btm.t199 VSS 0.282615f
C6357 C8_P_btm.t47 VSS 0.282615f
C6358 C8_P_btm.t182 VSS 0.282615f
C6359 C8_P_btm.t243 VSS 0.282615f
C6360 C8_P_btm.t36 VSS 0.282615f
C6361 C8_P_btm.t216 VSS 0.282615f
C6362 C8_P_btm.t192 VSS 0.282615f
C6363 C8_P_btm.t78 VSS 0.282615f
C6364 C8_P_btm.t20 VSS 0.282615f
C6365 C8_P_btm.t65 VSS 0.282615f
C6366 C8_P_btm.t247 VSS 0.282615f
C6367 C8_P_btm.t43 VSS 0.282615f
C6368 C8_P_btm.t116 VSS 0.282615f
C6369 C8_P_btm.t30 VSS 0.282615f
C6370 C8_P_btm.t83 VSS 0.282615f
C6371 C8_P_btm.t137 VSS 0.282615f
C6372 C8_P_btm.t70 VSS 0.282615f
C6373 C8_P_btm.t260 VSS 0.282615f
C6374 C8_P_btm.t56 VSS 0.282615f
C6375 C8_P_btm.t129 VSS 0.282615f
C6376 C8_P_btm.t167 VSS 0.282615f
C6377 C8_P_btm.t97 VSS 0.282615f
C6378 C8_P_btm.t164 VSS 0.282615f
C6379 C8_P_btm.t226 VSS 0.282615f
C6380 C8_P_btm.t139 VSS 0.282615f
C6381 C8_P_btm.t197 VSS 0.282615f
C6382 C8_P_btm.t261 VSS 0.313436f
C6383 C8_P_btm.t26 VSS 0.282615f
C6384 C8_P_btm.t232 VSS 0.282615f
C6385 C8_P_btm.t176 VSS 0.282615f
C6386 C8_P_btm.t111 VSS 0.282615f
C6387 C8_P_btm.t184 VSS 0.282615f
C6388 C8_P_btm.t23 VSS 0.282615f
C6389 C8_P_btm.t204 VSS 0.282615f
C6390 C8_P_btm.t266 VSS 0.282615f
C6391 C8_P_btm.t217 VSS 0.282615f
C6392 C8_P_btm.t156 VSS 0.282615f
C6393 C8_P_btm.t230 VSS 0.282615f
C6394 C8_P_btm.t171 VSS 0.282615f
C6395 C8_P_btm.t190 VSS 0.282615f
C6396 C8_P_btm.t201 VSS 0.282615f
C6397 C8_P_btm.t262 VSS 0.282615f
C6398 C8_P_btm.t72 VSS 0.282615f
C6399 C8_P_btm.t151 VSS 0.282615f
C6400 C8_P_btm.t85 VSS 0.282615f
C6401 C8_P_btm.t165 VSS 0.282615f
C6402 C8_P_btm.t119 VSS 0.282615f
C6403 C8_P_btm.t49 VSS 0.282615f
C6404 C8_P_btm.t121 VSS 0.282615f
C6405 C8_P_btm.t68 VSS 0.282615f
C6406 C8_P_btm.t25 VSS 0.282615f
C6407 C8_P_btm.t80 VSS 0.282615f
C6408 C8_P_btm.t27 VSS 0.282615f
C6409 C8_P_btm.t113 VSS 0.282615f
C6410 C8_P_btm.t40 VSS 0.282615f
C6411 C8_P_btm.t244 VSS 0.313436f
C6412 C8_P_btm.t212 VSS 0.282615f
C6413 C8_P_btm.t177 VSS 0.313436f
C6414 C8_P_btm.t237 VSS 0.282615f
C6415 C8_P_btm.t52 VSS 0.282615f
C6416 C8_P_btm.t223 VSS 0.282615f
C6417 C8_P_btm.t54 VSS 0.282615f
C6418 C8_P_btm.t210 VSS 0.282615f
C6419 C8_P_btm.t55 VSS 0.282615f
C6420 C8_P_btm.t59 VSS 0.282615f
C6421 C8_P_btm.t240 VSS 0.282615f
C6422 C8_P_btm.t105 VSS 0.282615f
C6423 C8_P_btm.t269 VSS 0.282615f
C6424 C8_P_btm.t118 VSS 0.282615f
C6425 C8_P_btm.t89 VSS 0.282615f
C6426 C8_P_btm.t255 VSS 0.282615f
C6427 C8_P_btm.t62 VSS 0.282615f
C6428 C8_P_btm.t272 VSS 0.282615f
C6429 C8_P_btm.t130 VSS 0.282615f
C6430 C8_P_btm.t107 VSS 0.282615f
C6431 C8_P_btm.t160 VSS 0.282615f
C6432 C8_P_btm.t94 VSS 0.282615f
C6433 C8_P_btm.t147 VSS 0.282615f
C6434 C8_P_btm.t66 VSS 0.282615f
C6435 C8_P_btm.t273 VSS 0.282615f
C6436 C8_P_btm.t194 VSS 0.282615f
C6437 C8_P_btm.t252 VSS 0.282615f
C6438 C8_P_btm.t189 VSS 0.282615f
C6439 C8_P_btm.t48 VSS 0.282615f
C6440 C8_P_btm.t161 VSS 0.282615f
C6441 C8_P_btm.t222 VSS 0.282615f
C6442 C8_P_btm.t31 VSS 0.313436f
C6443 C8_P_btm.t41 VSS 0.313436f
C6444 C8_P_btm.t50 VSS 0.313436f
C6445 C8_P_btm.t141 VSS 0.313436f
C6446 C8_P_btm.t51 VSS 0.282615f
C6447 C8_P_btm.t73 VSS 0.282615f
C6448 C8_P_btm.t93 VSS 0.313436f
C6449 C8_P_btm.t99 VSS 0.313436f
C6450 C8_P_btm.t238 VSS 0.282615f
C6451 C8_P_btm.t34 VSS 0.282615f
C6452 C8_P_btm.t16 VSS 0.325831f
C6453 C8_P_btm.n503 VSS 0.118587f
C6454 C8_P_btm.t10 VSS 0.325831f
C6455 C8_P_btm.t13 VSS 0.325831f
C6456 C8_P_btm.n506 VSS 0.102832f
C6457 C8_P_btm.t11 VSS 0.325831f
C6458 C8_P_btm.n507 VSS 0.102832f
C6459 C8_P_btm.t211 VSS 0.313436f
C6460 C8_P_btm.t136 VSS 0.282615f
C6461 C8_P_btm.t81 VSS 0.282615f
C6462 C8_P_btm.t14 VSS 0.325831f
C6463 C8_P_btm.n516 VSS 0.118587f
C6464 C8_P_btm.t115 VSS 0.313436f
C6465 C8_P_btm.t163 VSS 0.282615f
C6466 C8_P_btm.n520 VSS 0.102832f
C6467 C8_P_btm.t198 VSS 0.313436f
C6468 C8_P_btm.t96 VSS 0.282615f
C6469 C8_P_btm.t169 VSS 0.282615f
C6470 C8_P_btm.t229 VSS 0.282615f
C6471 C8_P_btm.t37 VSS 0.313436f
C6472 C8_P_btm.t38 VSS 0.313436f
C6473 C8_P_btm.t206 VSS 0.282615f
C6474 C8_P_btm.t144 VSS 0.282615f
C6475 C8_P_btm.t235 VSS 0.282615f
C6476 C8_P_btm.t173 VSS 0.313436f
C6477 C8_P_btm.t58 VSS 0.282615f
C6478 C8_P_btm.t241 VSS 0.313436f
C6479 C8_P_btm.t35 VSS 0.282615f
C6480 C8_P_btm.t213 VSS 0.282615f
C6481 C8_P_btm.t18 VSS 0.282615f
C6482 C8_P_btm.t77 VSS 0.313436f
C6483 C8_P_btm.t234 VSS 0.313436f
C6484 C8_P_btm.t248 VSS 0.282615f
C6485 C8_P_btm.t187 VSS 0.282615f
C6486 C8_P_btm.t22 VSS 0.282615f
C6487 C8_P_btm.t218 VSS 0.313436f
C6488 C8_P_btm.t100 VSS 0.282615f
C6489 C8_P_btm.t102 VSS 0.313436f
C6490 C8_P_btm.t76 VSS 0.282615f
C6491 C8_P_btm.t24 VSS 0.282615f
C6492 C8_P_btm.t114 VSS 0.282615f
C6493 C8_P_btm.t246 VSS 0.313436f
C6494 C8_P_btm.t158 VSS 0.313436f
C6495 C8_P_btm.t57 VSS 0.282615f
C6496 C8_P_btm.t168 VSS 0.282615f
C6497 C8_P_btm.t181 VSS 0.313436f
C6498 C8_P_btm.t209 VSS 0.313436f
C6499 C8_P_btm.t134 VSS 0.282615f
C6500 C8_P_btm.t79 VSS 0.282615f
C6501 C8_P_btm.t162 VSS 0.282615f
C6502 C8_P_btm.t112 VSS 0.313436f
C6503 C8_P_btm.t140 VSS 0.282615f
C6504 C8_P_btm.t60 VSS 0.313436f
C6505 C8_P_btm.t233 VSS 0.282615f
C6506 C8_P_btm.t268 VSS 0.282615f
C6507 C8_P_btm.t91 VSS 0.282615f
C6508 C8_P_btm.t257 VSS 0.313436f
C6509 C8_P_btm.t178 VSS 0.282615f
C6510 C8_P_btm.t120 VSS 0.282615f
C6511 C8_P_btm.t208 VSS 0.282615f
C6512 C8_P_btm.t146 VSS 0.313436f
C6513 C8_P_btm.t126 VSS 0.313436f
C6514 C8_P_btm.t253 VSS 0.282615f
C6515 C8_P_btm.t258 VSS 0.282615f
C6516 C8_P_btm.t180 VSS 0.282615f
C6517 C8_P_btm.t98 VSS 0.282615f
C6518 C8_P_btm.t152 VSS 0.282615f
C6519 C8_P_btm.t227 VSS 0.313436f
C6520 C8_P_btm.t191 VSS 0.313436f
C6521 C8_P_btm.t250 VSS 0.282615f
C6522 C8_P_btm.t186 VSS 0.282615f
C6523 C8_P_btm.t21 VSS 0.282615f
C6524 C8_P_btm.t215 VSS 0.282615f
C6525 C8_P_btm.t143 VSS 0.282615f
C6526 C8_P_btm.t219 VSS 0.282615f
C6527 C8_P_btm.t157 VSS 0.282615f
C6528 C8_P_btm.t90 VSS 0.282615f
C6529 C8_P_btm.t172 VSS 0.282615f
C6530 C8_P_btm.t221 VSS 0.282615f
C6531 C8_P_btm.t185 VSS 0.282615f
C6532 C8_P_btm.t265 VSS 0.282615f
C6533 C8_P_btm.t75 VSS 0.282615f
C6534 C8_P_btm.t155 VSS 0.282615f
C6535 C8_P_btm.t87 VSS 0.282615f
C6536 C8_P_btm.t33 VSS 0.282615f
C6537 C8_P_btm.t128 VSS 0.282615f
C6538 C8_P_btm.t53 VSS 0.282615f
C6539 C8_P_btm.t124 VSS 0.282615f
C6540 C8_P_btm.t69 VSS 0.282615f
C6541 C8_P_btm.t271 VSS 0.282615f
C6542 C8_P_btm.t82 VSS 0.282615f
C6543 C8_P_btm.t29 VSS 0.282615f
C6544 C8_P_btm.t236 VSS 0.282615f
C6545 C8_P_btm.t42 VSS 0.282615f
C6546 C8_P_btm.t251 VSS 0.282615f
C6547 C8_P_btm.t64 VSS 0.282615f
C6548 C8_P_btm.t256 VSS 0.282615f
C6549 C8_P_btm.t203 VSS 0.313436f
C6550 C8_P_btm.t166 VSS 0.282615f
C6551 C8_P_btm.t133 VSS 0.313436f
C6552 C8_P_btm.t193 VSS 0.282615f
C6553 C8_P_btm.t45 VSS 0.282615f
C6554 C8_P_btm.t179 VSS 0.282615f
C6555 C8_P_btm.t239 VSS 0.313436f
C6556 C8_P_btm.t145 VSS 0.313436f
C6557 C8_P_btm.t92 VSS 0.282615f
C6558 C8_P_btm.t174 VSS 0.282615f
C6559 C8_P_btm.t103 VSS 0.282615f
C6560 C8_P_btm.t108 VSS 0.313436f
C6561 C8_P_btm.t125 VSS 0.282615f
C6562 C8_P_btm.t263 VSS 0.313436f
C6563 C8_P_btm.t148 VSS 0.282615f
C6564 C8_P_btm.t224 VSS 0.282615f
C6565 C8_P_btm.t135 VSS 0.282615f
C6566 C8_P_btm.t195 VSS 0.313436f
C6567 C8_P_btm.t106 VSS 0.313436f
C6568 C8_P_btm.t117 VSS 0.282615f
C6569 C8_P_btm.t270 VSS 0.282615f
C6570 C8_P_btm.t61 VSS 0.282615f
C6571 C8_P_btm.t132 VSS 0.313436f
C6572 C8_P_btm.t86 VSS 0.282615f
C6573 C8_P_btm.t205 VSS 0.313436f
C6574 C8_P_btm.t39 VSS 0.282615f
C6575 C8_P_btm.t67 VSS 0.282615f
C6576 C8_P_btm.t249 VSS 0.282615f
C6577 C8_P_btm.t44 VSS 0.313436f
C6578 C8_P_btm.t46 VSS 0.313436f
C6579 C8_P_btm.t188 VSS 0.282615f
C6580 C8_P_btm.t267 VSS 0.282615f
C6581 C8_P_btm.t88 VSS 0.313436f
C6582 C8_P_btm.t63 VSS 0.313436f
C6583 C8_P_btm.t19 VSS 0.282615f
C6584 C8_P_btm.t259 VSS 0.282615f
C6585 C8_P_btm.t131 VSS 0.282615f
C6586 C8_P_btm.t228 VSS 0.313436f
C6587 C8_P_btm.t101 VSS 0.282615f
C6588 C8_P_btm.t159 VSS 0.313436f
C6589 C8_P_btm.t220 VSS 0.282615f
C6590 C8_P_btm.t28 VSS 0.282615f
C6591 C8_P_btm.t207 VSS 0.282615f
C6592 C8_P_btm.t254 VSS 0.313436f
C6593 C8_P_btm.t231 VSS 0.282615f
C6594 C8_P_btm.t123 VSS 0.282615f
C6595 C8_P_btm.t245 VSS 0.282615f
C6596 C8_P_btm.t183 VSS 0.313436f
C6597 C8_P_btm.t9 VSS 0.325831f
C6598 C8_P_btm.n890 VSS 0.118587f
C6599 C8_P_btm.t264 VSS 0.313436f
C6600 C8_P_btm.t149 VSS 0.282615f
C6601 C8_P_btm.t225 VSS 0.282615f
C6602 C8_P_btm.t138 VSS 0.282615f
C6603 C8_P_btm.t196 VSS 0.313436f
C6604 C8_P_btm.t15 VSS 0.313963f
C6605 C8_P_btm.n903 VSS 0.165799f
C6606 a_9521_45982.n4 VSS 0.392617f
C6607 a_9521_45982.n9 VSS 0.317497f
C6608 a_9521_45982.n11 VSS 0.404961f
C6609 a_9521_45982.n12 VSS 0.26483f
C6610 a_9521_45982.n14 VSS 0.156779f
C6611 a_9521_45982.n15 VSS 0.134617f
C6612 a_9521_45982.n17 VSS 0.117587f
C6613 a_n2810_44894.n1 VSS 0.174752f
C6614 a_n2810_44894.t8 VSS 0.534733f
C6615 a_n2810_44894.t4 VSS 0.536087f
C6616 a_n2810_44894.t7 VSS 0.534733f
C6617 a_n2810_44894.t10 VSS 0.536087f
C6618 a_n2810_44894.t9 VSS 0.534733f
C6619 a_n2810_44894.t5 VSS 0.536087f
C6620 a_n2810_44894.n2 VSS 0.256967f
C6621 a_n2810_44894.t6 VSS 0.534733f
C6622 a_n2810_44894.n3 VSS 0.265637f
C6623 a_n2810_44894.n4 VSS 0.309901f
C6624 a_n2810_44894.n5 VSS 0.277546f
C6625 a_n2810_44894.n6 VSS 0.256967f
C6626 a_n2810_44894.n7 VSS 0.277546f
C6627 a_n2810_44894.n8 VSS 0.256967f
C6628 a_n2810_44894.t11 VSS 0.550065f
C6629 a_n2810_44894.n9 VSS 0.496742f
C6630 a_n2810_44894.n10 VSS 6.00762f
C6631 a_n2810_44894.n11 VSS 5.11317f
C6632 C10_N_btm.n0 VSS 0.147281f
C6633 C10_N_btm.n1 VSS 0.142447f
C6634 C10_N_btm.n2 VSS 0.448097f
C6635 C10_N_btm.n3 VSS 0.142447f
C6636 C10_N_btm.n4 VSS 0.230042f
C6637 C10_N_btm.n5 VSS 0.142447f
C6638 C10_N_btm.n6 VSS 0.230042f
C6639 C10_N_btm.n7 VSS 0.142447f
C6640 C10_N_btm.n8 VSS 0.230042f
C6641 C10_N_btm.n9 VSS 0.142447f
C6642 C10_N_btm.n10 VSS 0.230042f
C6643 C10_N_btm.n11 VSS 0.142447f
C6644 C10_N_btm.n12 VSS 0.229719f
C6645 C10_N_btm.n13 VSS 0.142447f
C6646 C10_N_btm.n14 VSS 0.39544f
C6647 C10_N_btm.n15 VSS 0.216437f
C6648 C10_N_btm.n16 VSS 0.21129f
C6649 C10_N_btm.n17 VSS 0.316949f
C6650 C10_N_btm.n18 VSS 0.21129f
C6651 C10_N_btm.n19 VSS 0.16285f
C6652 C10_N_btm.n20 VSS 0.21129f
C6653 C10_N_btm.n21 VSS 0.184948f
C6654 C10_N_btm.n22 VSS 0.258762f
C6655 C10_N_btm.n23 VSS 0.25913f
C6656 C10_N_btm.n24 VSS 0.220601f
C6657 C10_N_btm.n25 VSS 0.218927f
C6658 C10_N_btm.n26 VSS 0.213708f
C6659 C10_N_btm.n27 VSS 0.323008f
C6660 C10_N_btm.n28 VSS 0.213708f
C6661 C10_N_btm.n29 VSS 0.166325f
C6662 C10_N_btm.n30 VSS 0.213708f
C6663 C10_N_btm.n31 VSS 0.186482f
C6664 C10_N_btm.n32 VSS 0.94021f
C6665 C10_N_btm.t1061 VSS 0.216874f
C6666 C10_N_btm.t1074 VSS 0.216874f
C6667 C10_N_btm.t1069 VSS 0.216874f
C6668 C10_N_btm.t1067 VSS 0.216874f
C6669 C10_N_btm.t1079 VSS 0.216874f
C6670 C10_N_btm.t1065 VSS 0.216874f
C6671 C10_N_btm.t1071 VSS 0.216874f
C6672 C10_N_btm.t1062 VSS 0.216874f
C6673 C10_N_btm.t1070 VSS 0.216874f
C6674 C10_N_btm.t298 VSS 0.208624f
C6675 C10_N_btm.t1059 VSS 0.216874f
C6676 C10_N_btm.t632 VSS 0.208624f
C6677 C10_N_btm.t857 VSS 0.208624f
C6678 C10_N_btm.t634 VSS 0.208624f
C6679 C10_N_btm.t797 VSS 0.18811f
C6680 C10_N_btm.t449 VSS 0.18811f
C6681 C10_N_btm.t692 VSS 0.18811f
C6682 C10_N_btm.t926 VSS 0.18811f
C6683 C10_N_btm.t635 VSS 0.18811f
C6684 C10_N_btm.t870 VSS 0.18811f
C6685 C10_N_btm.t493 VSS 0.18811f
C6686 C10_N_btm.t813 VSS 0.18811f
C6687 C10_N_btm.t477 VSS 0.208624f
C6688 C10_N_btm.t207 VSS 0.208624f
C6689 C10_N_btm.t96 VSS 0.18811f
C6690 C10_N_btm.t678 VSS 0.18811f
C6691 C10_N_btm.t913 VSS 0.18811f
C6692 C10_N_btm.t101 VSS 0.18811f
C6693 C10_N_btm.t860 VSS 0.18811f
C6694 C10_N_btm.t52 VSS 0.18811f
C6695 C10_N_btm.t262 VSS 0.18811f
C6696 C10_N_btm.t979 VSS 0.18811f
C6697 C10_N_btm.t499 VSS 0.208624f
C6698 C10_N_btm.t410 VSS 0.208624f
C6699 C10_N_btm.t182 VSS 0.18811f
C6700 C10_N_btm.t897 VSS 0.18811f
C6701 C10_N_btm.t80 VSS 0.18811f
C6702 C10_N_btm.t292 VSS 0.18811f
C6703 C10_N_btm.t34 VSS 0.18811f
C6704 C10_N_btm.t249 VSS 0.18811f
C6705 C10_N_btm.t464 VSS 0.18811f
C6706 C10_N_btm.t194 VSS 0.18811f
C6707 C10_N_btm.t435 VSS 0.208624f
C6708 C10_N_btm.t628 VSS 0.208624f
C6709 C10_N_btm.t385 VSS 0.18811f
C6710 C10_N_btm.t67 VSS 0.18811f
C6711 C10_N_btm.t282 VSS 0.18811f
C6712 C10_N_btm.t506 VSS 0.18811f
C6713 C10_N_btm.t511 VSS 0.18811f
C6714 C10_N_btm.t446 VSS 0.18811f
C6715 C10_N_btm.t690 VSS 0.18811f
C6716 C10_N_btm.t396 VSS 0.18811f
C6717 C10_N_btm.t783 VSS 0.208624f
C6718 C10_N_btm.t972 VSS 0.208624f
C6719 C10_N_btm.t713 VSS 0.18811f
C6720 C10_N_btm.t1041 VSS 0.18811f
C6721 C10_N_btm.t614 VSS 0.18811f
C6722 C10_N_btm.t851 VSS 0.18811f
C6723 C10_N_btm.t552 VSS 0.18811f
C6724 C10_N_btm.t792 VSS 0.18811f
C6725 C10_N_btm.t478 VSS 0.18811f
C6726 C10_N_btm.t736 VSS 0.18811f
C6727 C10_N_btm.t531 VSS 0.208624f
C6728 C10_N_btm.t725 VSS 0.208624f
C6729 C10_N_btm.t498 VSS 0.18811f
C6730 C10_N_btm.t166 VSS 0.18811f
C6731 C10_N_btm.t377 VSS 0.18811f
C6732 C10_N_btm.t605 VSS 0.18811f
C6733 C10_N_btm.t326 VSS 0.18811f
C6734 C10_N_btm.t540 VSS 0.18811f
C6735 C10_N_btm.t388 VSS 0.18811f
C6736 C10_N_btm.t991 VSS 0.18811f
C6737 C10_N_btm.t758 VSS 0.208624f
C6738 C10_N_btm.t698 VSS 0.18811f
C6739 C10_N_btm.t360 VSS 0.18811f
C6740 C10_N_btm.t592 VSS 0.18811f
C6741 C10_N_btm.t827 VSS 0.18811f
C6742 C10_N_btm.t1057 VSS 0.18811f
C6743 C10_N_btm.t776 VSS 0.18811f
C6744 C10_N_btm.t1014 VSS 0.18811f
C6745 C10_N_btm.t710 VSS 0.18811f
C6746 C10_N_btm.t954 VSS 0.18811f
C6747 C10_N_btm.t608 VSS 0.18811f
C6748 C10_N_btm.t895 VSS 0.18811f
C6749 C10_N_btm.t78 VSS 0.18811f
C6750 C10_N_btm.t647 VSS 0.18811f
C6751 C10_N_btm.t878 VSS 0.18811f
C6752 C10_N_btm.t236 VSS 0.18811f
C6753 C10_N_btm.t821 VSS 0.18811f
C6754 C10_N_btm.t83 VSS 0.18811f
C6755 C10_N_btm.t274 VSS 0.18811f
C6756 C10_N_btm.t1008 VSS 0.18811f
C6757 C10_N_btm.t180 VSS 0.18811f
C6758 C10_N_btm.t951 VSS 0.18811f
C6759 C10_N_btm.t127 VSS 0.208624f
C6760 C10_N_btm.t395 VSS 0.208624f
C6761 C10_N_btm.t158 VSS 0.208624f
C6762 C10_N_btm.t333 VSS 0.208624f
C6763 C10_N_btm.t237 VSS 0.18811f
C6764 C10_N_btm.t317 VSS 0.18811f
C6765 C10_N_btm.t759 VSS 0.18811f
C6766 C10_N_btm.t232 VSS 0.18811f
C6767 C10_N_btm.t595 VSS 0.18811f
C6768 C10_N_btm.t173 VSS 0.18811f
C6769 C10_N_btm.t383 VSS 0.18811f
C6770 C10_N_btm.t670 VSS 0.18811f
C6771 C10_N_btm.t762 VSS 0.208624f
C6772 C10_N_btm.t959 VSS 0.208624f
C6773 C10_N_btm.t657 VSS 0.18811f
C6774 C10_N_btm.t944 VSS 0.18811f
C6775 C10_N_btm.t596 VSS 0.18811f
C6776 C10_N_btm.t835 VSS 0.18811f
C6777 C10_N_btm.t69 VSS 0.18811f
C6778 C10_N_btm.t782 VSS 0.18811f
C6779 C10_N_btm.t1020 VSS 0.18811f
C6780 C10_N_btm.t520 VSS 0.18811f
C6781 C10_N_btm.t937 VSS 0.208624f
C6782 C10_N_btm.t76 VSS 0.208624f
C6783 C10_N_btm.t824 VSS 0.18811f
C6784 C10_N_btm.t62 VSS 0.18811f
C6785 C10_N_btm.t771 VSS 0.18811f
C6786 C10_N_btm.t1021 VSS 0.18811f
C6787 C10_N_btm.t484 VSS 0.18811f
C6788 C10_N_btm.t952 VSS 0.18811f
C6789 C10_N_btm.t129 VSS 0.18811f
C6790 C10_N_btm.t391 VSS 0.18811f
C6791 C10_N_btm.t775 VSS 0.208624f
C6792 C10_N_btm.t514 VSS 0.208624f
C6793 C10_N_btm.t998 VSS 0.18811f
C6794 C10_N_btm.t240 VSS 0.18811f
C6795 C10_N_btm.t943 VSS 0.18811f
C6796 C10_N_btm.t120 VSS 0.18811f
C6797 C10_N_btm.t1045 VSS 0.18811f
C6798 C10_N_btm.t68 VSS 0.18811f
C6799 C10_N_btm.t283 VSS 0.18811f
C6800 C10_N_btm.t557 VSS 0.18811f
C6801 C10_N_btm.t227 VSS 0.208624f
C6802 C10_N_btm.t390 VSS 0.208624f
C6803 C10_N_btm.t468 VSS 0.18811f
C6804 C10_N_btm.t380 VSS 0.18811f
C6805 C10_N_btm.t60 VSS 0.18811f
C6806 C10_N_btm.t278 VSS 0.18811f
C6807 C10_N_btm.t544 VSS 0.18811f
C6808 C10_N_btm.t481 VSS 0.18811f
C6809 C10_N_btm.t442 VSS 0.18811f
C6810 C10_N_btm.t729 VSS 0.18811f
C6811 C10_N_btm.t372 VSS 0.208624f
C6812 C10_N_btm.t556 VSS 0.208624f
C6813 C10_N_btm.t269 VSS 0.18811f
C6814 C10_N_btm.t538 VSS 0.18811f
C6815 C10_N_btm.t235 VSS 0.18811f
C6816 C10_N_btm.t437 VSS 0.18811f
C6817 C10_N_btm.t716 VSS 0.18811f
C6818 C10_N_btm.t386 VSS 0.18811f
C6819 C10_N_btm.t615 VSS 0.18811f
C6820 C10_N_btm.t448 VSS 0.18811f
C6821 C10_N_btm.t1078 VSS 0.216874f
C6822 C10_N_btm.t1077 VSS 0.216874f
C6823 C10_N_btm.t1066 VSS 0.216874f
C6824 C10_N_btm.t1058 VSS 0.216874f
C6825 C10_N_btm.t1068 VSS 0.216874f
C6826 C10_N_btm.t1060 VSS 0.216874f
C6827 C10_N_btm.t1073 VSS 0.216874f
C6828 C10_N_btm.t1063 VSS 0.216874f
C6829 C10_N_btm.t1076 VSS 0.216874f
C6830 C10_N_btm.t1072 VSS 0.216874f
C6831 C10_N_btm.t139 VSS 0.208624f
C6832 C10_N_btm.t451 VSS 0.18811f
C6833 C10_N_btm.t189 VSS 0.18811f
C6834 C10_N_btm.t1025 VSS 0.18811f
C6835 C10_N_btm.t285 VSS 0.18811f
C6836 C10_N_btm.t118 VSS 0.18811f
C6837 C10_N_btm.t840 VSS 0.18811f
C6838 C10_N_btm.t123 VSS 0.18811f
C6839 C10_N_btm.t889 VSS 0.18811f
C6840 C10_N_btm.t1003 VSS 0.208624f
C6841 C10_N_btm.t1064 VSS 0.216874f
C6842 C10_N_btm.t178 VSS 0.18811f
C6843 C10_N_btm.t636 VSS 0.208624f
C6844 C10_N_btm.t871 VSS 0.18811f
C6845 C10_N_btm.t1054 VSS 0.18811f
C6846 C10_N_btm.t814 VSS 0.18811f
C6847 C10_N_btm.t480 VSS 0.18811f
C6848 C10_N_btm.t702 VSS 0.18811f
C6849 C10_N_btm.t995 VSS 0.18811f
C6850 C10_N_btm.t653 VSS 0.18811f
C6851 C10_N_btm.t883 VSS 0.18811f
C6852 C10_N_btm.t599 VSS 0.18811f
C6853 C10_N_btm.t831 VSS 0.208624f
C6854 C10_N_btm.t930 VSS 0.208624f
C6855 C10_N_btm.t208 VSS 0.18811f
C6856 C10_N_btm.t984 VSS 0.18811f
C6857 C10_N_btm.t746 VSS 0.18811f
C6858 C10_N_btm.t53 VSS 0.18811f
C6859 C10_N_btm.t802 VSS 0.18811f
C6860 C10_N_btm.t562 VSS 0.18811f
C6861 C10_N_btm.t915 VSS 0.18811f
C6862 C10_N_btm.t621 VSS 0.18811f
C6863 C10_N_btm.t966 VSS 0.18811f
C6864 C10_N_btm.t728 VSS 0.208624f
C6865 C10_N_btm.t600 VSS 0.18811f
C6866 C10_N_btm.t463 VSS 0.208624f
C6867 C10_N_btm.t695 VSS 0.18811f
C6868 C10_N_btm.t355 VSS 0.18811f
C6869 C10_N_btm.t646 VSS 0.18811f
C6870 C10_N_btm.t309 VSS 0.18811f
C6871 C10_N_btm.t527 VSS 0.18811f
C6872 C10_N_btm.t820 VSS 0.18811f
C6873 C10_N_btm.t490 VSS 0.18811f
C6874 C10_N_btm.t706 VSS 0.18811f
C6875 C10_N_btm.t1007 VSS 0.18811f
C6876 C10_N_btm.t662 VSS 0.208624f
C6877 C10_N_btm.t756 VSS 0.208624f
C6878 C10_N_btm.t213 VSS 0.18811f
C6879 C10_N_btm.t810 VSS 0.18811f
C6880 C10_N_btm.t569 VSS 0.18811f
C6881 C10_N_btm.t921 VSS 0.18811f
C6882 C10_N_btm.t630 VSS 0.18811f
C6883 C10_N_btm.t398 VSS 0.18811f
C6884 C10_N_btm.t740 VSS 0.18811f
C6885 C10_N_btm.t447 VSS 0.18811f
C6886 C10_N_btm.t794 VSS 0.18811f
C6887 C10_N_btm.t555 VSS 0.208624f
C6888 C10_N_btm.t429 VSS 0.18811f
C6889 C10_N_btm.t303 VSS 0.208624f
C6890 C10_N_btm.t1056 VSS 0.18811f
C6891 C10_N_btm.t202 VSS 0.18811f
C6892 C10_N_btm.t483 VSS 0.18811f
C6893 C10_N_btm.t159 VSS 0.18811f
C6894 C10_N_btm.t367 VSS 0.18811f
C6895 C10_N_btm.t654 VSS 0.18811f
C6896 C10_N_btm.t318 VSS 0.18811f
C6897 C10_N_btm.t534 VSS 0.18811f
C6898 C10_N_btm.t832 VSS 0.18811f
C6899 C10_N_btm.t597 VSS 0.208624f
C6900 C10_N_btm.t151 VSS 0.208624f
C6901 C10_N_btm.t466 VSS 0.18811f
C6902 C10_N_btm.t195 VSS 0.18811f
C6903 C10_N_btm.t47 VSS 0.18811f
C6904 C10_N_btm.t291 VSS 0.18811f
C6905 C10_N_btm.t35 VSS 0.18811f
C6906 C10_N_btm.t844 VSS 0.18811f
C6907 C10_N_btm.t131 VSS 0.18811f
C6908 C10_N_btm.t898 VSS 0.18811f
C6909 C10_N_btm.t91 VSS 0.18811f
C6910 C10_N_btm.t1016 VSS 0.208624f
C6911 C10_N_btm.t270 VSS 0.18811f
C6912 C10_N_btm.t150 VSS 0.208624f
C6913 C10_N_btm.t356 VSS 0.18811f
C6914 C10_N_btm.t85 VSS 0.18811f
C6915 C10_N_btm.t310 VSS 0.18811f
C6916 C10_N_btm.t941 VSS 0.18811f
C6917 C10_N_btm.t210 VSS 0.18811f
C6918 C10_N_btm.t494 VSS 0.18811f
C6919 C10_N_btm.t165 VSS 0.18811f
C6920 C10_N_btm.t376 VSS 0.18811f
C6921 C10_N_btm.t663 VSS 0.18811f
C6922 C10_N_btm.t324 VSS 0.208624f
C6923 C10_N_btm.t46 VSS 0.208624f
C6924 C10_N_btm.t304 VSS 0.18811f
C6925 C10_N_btm.t45 VSS 0.18811f
C6926 C10_N_btm.t854 VSS 0.18811f
C6927 C10_N_btm.t138 VSS 0.18811f
C6928 C10_N_btm.t909 VSS 0.18811f
C6929 C10_N_btm.t674 VSS 0.18811f
C6930 C10_N_btm.t1024 VSS 0.18811f
C6931 C10_N_btm.t720 VSS 0.18811f
C6932 C10_N_btm.t110 VSS 0.18811f
C6933 C10_N_btm.t838 VSS 0.208624f
C6934 C10_N_btm.t475 VSS 0.18811f
C6935 C10_N_btm.t561 VSS 0.208624f
C6936 C10_N_btm.t801 VSS 0.18811f
C6937 C10_N_btm.t455 VSS 0.18811f
C6938 C10_N_btm.t745 VSS 0.18811f
C6939 C10_N_btm.t402 VSS 0.18811f
C6940 C10_N_btm.t640 VSS 0.18811f
C6941 C10_N_btm.t929 VSS 0.18811f
C6942 C10_N_btm.t577 VSS 0.18811f
C6943 C10_N_btm.t816 VSS 0.18811f
C6944 C10_N_btm.t1033 VSS 0.18811f
C6945 C10_N_btm.t763 VSS 0.208624f
C6946 C10_N_btm.t863 VSS 0.208624f
C6947 C10_N_btm.t152 VSS 0.18811f
C6948 C10_N_btm.t917 VSS 0.18811f
C6949 C10_N_btm.t682 VSS 0.18811f
C6950 C10_N_btm.t55 VSS 0.18811f
C6951 C10_N_btm.t733 VSS 0.18811f
C6952 C10_N_btm.t1030 VSS 0.18811f
C6953 C10_N_btm.t845 VSS 0.18811f
C6954 C10_N_btm.t548 VSS 0.18811f
C6955 C10_N_btm.t899 VSS 0.18811f
C6956 C10_N_btm.t669 VSS 0.208624f
C6957 C10_N_btm.t999 VSS 0.18811f
C6958 C10_N_btm.t397 VSS 0.208624f
C6959 C10_N_btm.t629 VSS 0.18811f
C6960 C10_N_btm.t296 VSS 0.18811f
C6961 C10_N_btm.t568 VSS 0.18811f
C6962 C10_N_btm.t250 VSS 0.18811f
C6963 C10_N_btm.t470 VSS 0.18811f
C6964 C10_N_btm.t755 VSS 0.18811f
C6965 C10_N_btm.t413 VSS 0.18811f
C6966 C10_N_btm.t649 VSS 0.18811f
C6967 C10_N_btm.t938 VSS 0.18811f
C6968 C10_N_btm.t588 VSS 0.208624f
C6969 C10_N_btm.t691 VSS 0.208624f
C6970 C10_N_btm.t51 VSS 0.18811f
C6971 C10_N_btm.t743 VSS 0.18811f
C6972 C10_N_btm.t509 VSS 0.18811f
C6973 C10_N_btm.t855 VSS 0.18811f
C6974 C10_N_btm.t559 VSS 0.18811f
C6975 C10_N_btm.t338 VSS 0.18811f
C6976 C10_N_btm.t675 VSS 0.18811f
C6977 C10_N_btm.t1049 VSS 0.18811f
C6978 C10_N_btm.t721 VSS 0.18811f
C6979 C10_N_btm.t892 VSS 0.208624f
C6980 C10_N_btm.t366 VSS 0.18811f
C6981 C10_N_btm.t992 VSS 0.208624f
C6982 C10_N_btm.t456 VSS 0.18811f
C6983 C10_N_btm.t144 VSS 0.18811f
C6984 C10_N_btm.t403 VSS 0.18811f
C6985 C10_N_btm.t97 VSS 0.18811f
C6986 C10_N_btm.t307 VSS 0.18811f
C6987 C10_N_btm.t578 VSS 0.18811f
C6988 C10_N_btm.t260 VSS 0.18811f
C6989 C10_N_btm.t489 VSS 0.18811f
C6990 C10_N_btm.t764 VSS 0.18811f
C6991 C10_N_btm.t423 VSS 0.208624f
C6992 C10_N_btm.t689 VSS 0.208624f
C6993 C10_N_btm.t289 VSS 0.18811f
C6994 C10_N_btm.t567 VSS 0.18811f
C6995 C10_N_btm.t247 VSS 0.18811f
C6996 C10_N_btm.t462 VSS 0.18811f
C6997 C10_N_btm.t752 VSS 0.18811f
C6998 C10_N_btm.t407 VSS 0.18811f
C6999 C10_N_btm.t645 VSS 0.18811f
C7000 C10_N_btm.t934 VSS 0.18811f
C7001 C10_N_btm.t585 VSS 0.208624f
C7002 C10_N_btm.t1046 VSS 0.208624f
C7003 C10_N_btm.t864 VSS 0.18811f
C7004 C10_N_btm.t565 VSS 0.18811f
C7005 C10_N_btm.t343 VSS 0.18811f
C7006 C10_N_btm.t683 VSS 0.18811f
C7007 C10_N_btm.t393 VSS 0.18811f
C7008 C10_N_btm.t181 VSS 0.18811f
C7009 C10_N_btm.t502 VSS 0.18811f
C7010 C10_N_btm.t496 VSS 0.18811f
C7011 C10_N_btm.t549 VSS 0.18811f
C7012 C10_N_btm.t332 VSS 0.208624f
C7013 C10_N_btm.t624 VSS 0.18811f
C7014 C10_N_btm.t619 VSS 0.208624f
C7015 C10_N_btm.t714 VSS 0.18811f
C7016 C10_N_btm.t1043 VSS 0.18811f
C7017 C10_N_btm.t673 VSS 0.18811f
C7018 C10_N_btm.t337 VSS 0.18811f
C7019 C10_N_btm.t554 VSS 0.18811f
C7020 C10_N_btm.t850 VSS 0.18811f
C7021 C10_N_btm.t505 VSS 0.18811f
C7022 C10_N_btm.t739 VSS 0.18811f
C7023 C10_N_btm.t1035 VSS 0.18811f
C7024 C10_N_btm.t328 VSS 0.208624f
C7025 C10_N_btm.t667 VSS 0.18811f
C7026 C10_N_btm.t381 VSS 0.18811f
C7027 C10_N_btm.t169 VSS 0.18811f
C7028 C10_N_btm.t501 VSS 0.18811f
C7029 C10_N_btm.t225 VSS 0.18811f
C7030 C10_N_btm.t903 VSS 0.18811f
C7031 C10_N_btm.t315 VSS 0.18811f
C7032 C10_N_btm.t109 VSS 0.18811f
C7033 C10_N_btm.t359 VSS 0.18811f
C7034 C10_N_btm.t155 VSS 0.208624f
C7035 C10_N_btm.t886 VSS 0.208624f
C7036 C10_N_btm.t580 VSS 0.18811f
C7037 C10_N_btm.t873 VSS 0.18811f
C7038 C10_N_btm.t58 VSS 0.18811f
C7039 C10_N_btm.t765 VSS 0.18811f
C7040 C10_N_btm.t1000 VSS 0.18811f
C7041 C10_N_btm.t246 VSS 0.18811f
C7042 C10_N_btm.t945 VSS 0.18811f
C7043 C10_N_btm.t122 VSS 0.18811f
C7044 C10_N_btm.t887 VSS 0.18811f
C7045 C10_N_btm.t71 VSS 0.18811f
C7046 C10_N_btm.t284 VSS 0.18811f
C7047 C10_N_btm.t94 VSS 0.18811f
C7048 C10_N_btm.t598 VSS 0.18811f
C7049 C10_N_btm.t450 VSS 0.18811f
C7050 C10_N_btm.t136 VSS 0.18811f
C7051 C10_N_btm.t400 VSS 0.18811f
C7052 C10_N_btm.t90 VSS 0.18811f
C7053 C10_N_btm.t302 VSS 0.18811f
C7054 C10_N_btm.t574 VSS 0.18811f
C7055 C10_N_btm.t257 VSS 0.18811f
C7056 C10_N_btm.t482 VSS 0.18811f
C7057 C10_N_btm.t760 VSS 0.18811f
C7058 C10_N_btm.t421 VSS 0.208624f
C7059 C10_N_btm.t980 VSS 0.208624f
C7060 C10_N_btm.t264 VSS 0.208624f
C7061 C10_N_btm.t925 VSS 0.18811f
C7062 C10_N_btm.t575 VSS 0.18811f
C7063 C10_N_btm.t815 VSS 0.18811f
C7064 C10_N_btm.t573 VSS 0.18811f
C7065 C10_N_btm.t761 VSS 0.18811f
C7066 C10_N_btm.t996 VSS 0.18811f
C7067 C10_N_btm.t176 VSS 0.18811f
C7068 C10_N_btm.t942 VSS 0.18811f
C7069 C10_N_btm.t774 VSS 0.18811f
C7070 C10_N_btm.t833 VSS 0.18811f
C7071 C10_N_btm.t66 VSS 0.18811f
C7072 C10_N_btm.t281 VSS 0.18811f
C7073 C10_N_btm.t486 VSS 0.18811f
C7074 C10_N_btm.t703 VSS 0.18811f
C7075 C10_N_btm.t997 VSS 0.18811f
C7076 C10_N_btm.t655 VSS 0.18811f
C7077 C10_N_btm.t884 VSS 0.18811f
C7078 C10_N_btm.t1032 VSS 0.18811f
C7079 C10_N_btm.t412 VSS 0.18811f
C7080 C10_N_btm.t532 VSS 0.18811f
C7081 C10_N_btm.t781 VSS 0.18811f
C7082 C10_N_btm.t1018 VSS 0.18811f
C7083 C10_N_btm.t185 VSS 0.18811f
C7084 C10_N_btm.t900 VSS 0.18811f
C7085 C10_N_btm.t1051 VSS 0.18811f
C7086 C10_N_btm.t349 VSS 0.18811f
C7087 C10_N_btm.t37 VSS 0.18811f
C7088 C10_N_btm.t295 VSS 0.18811f
C7089 C10_N_btm.t95 VSS 0.18811f
C7090 C10_N_btm.t196 VSS 0.18811f
C7091 C10_N_btm.t469 VSS 0.18811f
C7092 C10_N_btm.t153 VSS 0.18811f
C7093 C10_N_btm.t357 VSS 0.18811f
C7094 C10_N_btm.t589 VSS 0.18811f
C7095 C10_N_btm.t313 VSS 0.18811f
C7096 C10_N_btm.t530 VSS 0.18811f
C7097 C10_N_btm.t214 VSS 0.18811f
C7098 C10_N_btm.t497 VSS 0.18811f
C7099 C10_N_btm.t709 VSS 0.18811f
C7100 C10_N_btm.t416 VSS 0.18811f
C7101 C10_N_btm.t699 VSS 0.18811f
C7102 C10_N_btm.t940 VSS 0.18811f
C7103 C10_N_btm.t591 VSS 0.18811f
C7104 C10_N_btm.t826 VSS 0.18811f
C7105 C10_N_btm.t64 VSS 0.18811f
C7106 C10_N_btm.t777 VSS 0.18811f
C7107 C10_N_btm.t1029 VSS 0.18811f
C7108 C10_N_btm.t711 VSS 0.18811f
C7109 C10_N_btm.t955 VSS 0.18811f
C7110 C10_N_btm.t130 VSS 0.18811f
C7111 C10_N_btm.t894 VSS 0.18811f
C7112 C10_N_btm.t79 VSS 0.18811f
C7113 C10_N_btm.t290 VSS 0.18811f
C7114 C10_N_btm.t40 VSS 0.18811f
C7115 C10_N_btm.t248 VSS 0.18811f
C7116 C10_N_btm.t967 VSS 0.18811f
C7117 C10_N_btm.t149 VSS 0.18811f
C7118 C10_N_btm.t408 VSS 0.18811f
C7119 C10_N_btm.t105 VSS 0.18811f
C7120 C10_N_btm.t311 VSS 0.18811f
C7121 C10_N_btm.t586 VSS 0.18811f
C7122 C10_N_btm.t146 VSS 0.208624f
C7123 C10_N_btm.t212 VSS 0.208624f
C7124 C10_N_btm.t100 VSS 0.18811f
C7125 C10_N_btm.t800 VSS 0.18811f
C7126 C10_N_btm.t975 VSS 0.18811f
C7127 C10_N_btm.t209 VSS 0.18811f
C7128 C10_N_btm.t983 VSS 0.18811f
C7129 C10_N_btm.t164 VSS 0.18811f
C7130 C10_N_btm.t183 VSS 0.18811f
C7131 C10_N_btm.t226 VSS 0.18811f
C7132 C10_N_btm.t323 VSS 0.18811f
C7133 C10_N_btm.t198 VSS 0.18811f
C7134 C10_N_btm.t271 VSS 0.18811f
C7135 C10_N_btm.t772 VSS 0.18811f
C7136 C10_N_btm.t312 VSS 0.18811f
C7137 C10_N_btm.t528 VSS 0.18811f
C7138 C10_N_btm.t822 VSS 0.18811f
C7139 C10_N_btm.t495 VSS 0.18811f
C7140 C10_N_btm.t707 VSS 0.18811f
C7141 C10_N_btm.t1009 VSS 0.18811f
C7142 C10_N_btm.t664 VSS 0.18811f
C7143 C10_N_btm.t890 VSS 0.18811f
C7144 C10_N_btm.t603 VSS 0.18811f
C7145 C10_N_btm.t841 VSS 0.18811f
C7146 C10_N_btm.t221 VSS 0.18811f
C7147 C10_N_btm.t722 VSS 0.18811f
C7148 C10_N_btm.t1028 VSS 0.18811f
C7149 C10_N_btm.t191 VSS 0.18811f
C7150 C10_N_btm.t910 VSS 0.18811f
C7151 C10_N_btm.t141 VSS 0.18811f
C7152 C10_N_btm.t856 VSS 0.18811f
C7153 C10_N_btm.t49 VSS 0.18811f
C7154 C10_N_btm.t306 VSS 0.18811f
C7155 C10_N_btm.t54 VSS 0.18811f
C7156 C10_N_btm.t203 VSS 0.18811f
C7157 C10_N_btm.t424 VSS 0.18811f
C7158 C10_N_btm.t161 VSS 0.18811f
C7159 C10_N_btm.t369 VSS 0.18811f
C7160 C10_N_btm.t245 VSS 0.18811f
C7161 C10_N_btm.t319 VSS 0.18811f
C7162 C10_N_btm.t536 VSS 0.18811f
C7163 C10_N_btm.t263 VSS 0.18811f
C7164 C10_N_btm.t523 VSS 0.18811f
C7165 C10_N_btm.t767 VSS 0.18811f
C7166 C10_N_btm.t426 VSS 0.18811f
C7167 C10_N_btm.t659 VSS 0.18811f
C7168 C10_N_btm.t946 VSS 0.18811f
C7169 C10_N_btm.t601 VSS 0.18811f
C7170 C10_N_btm.t837 VSS 0.18811f
C7171 C10_N_btm.t539 VSS 0.18811f
C7172 C10_N_btm.t786 VSS 0.18811f
C7173 C10_N_btm.t1022 VSS 0.18811f
C7174 C10_N_btm.t718 VSS 0.18811f
C7175 C10_N_btm.t963 VSS 0.18811f
C7176 C10_N_btm.t137 VSS 0.18811f
C7177 C10_N_btm.t853 VSS 0.18811f
C7178 C10_N_btm.t92 VSS 0.18811f
C7179 C10_N_btm.t795 VSS 0.18811f
C7180 C10_N_btm.t43 VSS 0.18811f
C7181 C10_N_btm.t258 VSS 0.18811f
C7182 C10_N_btm.t977 VSS 0.18811f
C7183 C10_N_btm.t160 VSS 0.18811f
C7184 C10_N_btm.t422 VSS 0.18811f
C7185 C10_N_btm.t791 VSS 0.208624f
C7186 C10_N_btm.t82 VSS 0.18811f
C7187 C10_N_btm.t846 VSS 0.18811f
C7188 C10_N_btm.t610 VSS 0.18811f
C7189 C10_N_btm.t958 VSS 0.18811f
C7190 C10_N_btm.t668 VSS 0.18811f
C7191 C10_N_btm.t430 VSS 0.18811f
C7192 C10_N_btm.t780 VSS 0.18811f
C7193 C10_N_btm.t519 VSS 0.18811f
C7194 C10_N_btm.t830 VSS 0.18811f
C7195 C10_N_btm.t594 VSS 0.18811f
C7196 C10_N_btm.t362 VSS 0.18811f
C7197 C10_N_btm.t652 VSS 0.18811f
C7198 C10_N_btm.t419 VSS 0.18811f
C7199 C10_N_btm.t199 VSS 0.18811f
C7200 C10_N_btm.t479 VSS 0.18811f
C7201 C10_N_btm.t254 VSS 0.18811f
C7202 C10_N_btm.t572 VSS 0.18811f
C7203 C10_N_btm.t300 VSS 0.18811f
C7204 C10_N_btm.t87 VSS 0.18811f
C7205 C10_N_btm.t399 VSS 0.18811f
C7206 C10_N_btm.t186 VSS 0.18811f
C7207 C10_N_btm.t960 VSS 0.18811f
C7208 C10_N_btm.t197 VSS 0.18811f
C7209 C10_N_btm.t111 VSS 0.18811f
C7210 C10_N_btm.t734 VSS 0.18811f
C7211 C10_N_btm.t38 VSS 0.18811f
C7212 C10_N_btm.t847 VSS 0.18811f
C7213 C10_N_btm.t84 VSS 0.18811f
C7214 C10_N_btm.t901 VSS 0.18811f
C7215 C10_N_btm.t671 VSS 0.18811f
C7216 C10_N_btm.t1019 VSS 0.18811f
C7217 C10_N_btm.t712 VSS 0.18811f
C7218 C10_N_btm.t612 VSS 0.18811f
C7219 C10_N_btm.t834 VSS 0.18811f
C7220 C10_N_btm.t535 VSS 0.18811f
C7221 C10_N_btm.t885 VSS 0.18811f
C7222 C10_N_btm.t656 VSS 0.18811f
C7223 C10_N_btm.t368 VSS 0.18811f
C7224 C10_N_btm.t704 VSS 0.18811f
C7225 C10_N_btm.t487 VSS 0.18811f
C7226 C10_N_btm.t259 VSS 0.18811f
C7227 C10_N_btm.t521 VSS 0.18811f
C7228 C10_N_btm.t305 VSS 0.18811f
C7229 C10_N_btm.t639 VSS 0.18811f
C7230 C10_N_btm.t351 VSS 0.18811f
C7231 C10_N_btm.t140 VSS 0.18811f
C7232 C10_N_btm.t453 VSS 0.18811f
C7233 C10_N_btm.t190 VSS 0.18811f
C7234 C10_N_btm.t508 VSS 0.18811f
C7235 C10_N_btm.t1015 VSS 0.18811f
C7236 C10_N_btm.t778 VSS 0.18811f
C7237 C10_N_btm.t518 VSS 0.18811f
C7238 C10_N_btm.t828 VSS 0.18811f
C7239 C10_N_btm.t593 VSS 0.18811f
C7240 C10_N_btm.t882 VSS 0.18811f
C7241 C10_N_btm.t651 VSS 0.18811f
C7242 C10_N_btm.t418 VSS 0.18811f
C7243 C10_N_btm.t701 VSS 0.18811f
C7244 C10_N_btm.t473 VSS 0.18811f
C7245 C10_N_btm.t253 VSS 0.18811f
C7246 C10_N_btm.t571 VSS 0.18811f
C7247 C10_N_btm.t299 VSS 0.18811f
C7248 C10_N_btm.t633 VSS 0.208624f
C7249 C10_N_btm.t862 VSS 0.18811f
C7250 C10_N_btm.t806 VSS 0.208624f
C7251 C10_N_btm.t461 VSS 0.18811f
C7252 C10_N_btm.t750 VSS 0.18811f
C7253 C10_N_btm.t406 VSS 0.18811f
C7254 C10_N_btm.t644 VSS 0.18811f
C7255 C10_N_btm.t877 VSS 0.18811f
C7256 C10_N_btm.t584 VSS 0.18811f
C7257 C10_N_btm.t819 VSS 0.18811f
C7258 C10_N_btm.t116 VSS 0.18811f
C7259 C10_N_btm.t770 VSS 0.18811f
C7260 C10_N_btm.t1005 VSS 0.18811f
C7261 C10_N_btm.t661 VSS 0.18811f
C7262 C10_N_btm.t949 VSS 0.18811f
C7263 C10_N_btm.t125 VSS 0.18811f
C7264 C10_N_btm.t242 VSS 0.18811f
C7265 C10_N_btm.t438 VSS 0.18811f
C7266 C10_N_btm.t719 VSS 0.18811f
C7267 C10_N_btm.t1047 VSS 0.18811f
C7268 C10_N_btm.t616 VSS 0.18811f
C7269 C10_N_btm.t908 VSS 0.18811f
C7270 C10_N_btm.t558 VSS 0.18811f
C7271 C10_N_btm.t796 VSS 0.18811f
C7272 C10_N_btm.t507 VSS 0.18811f
C7273 C10_N_btm.t742 VSS 0.18811f
C7274 C10_N_btm.t978 VSS 0.18811f
C7275 C10_N_btm.t631 VSS 0.18811f
C7276 C10_N_btm.t923 VSS 0.18811f
C7277 C10_N_btm.t216 VSS 0.18811f
C7278 C10_N_btm.t811 VSS 0.18811f
C7279 C10_N_btm.t230 VSS 0.18811f
C7280 C10_N_btm.t374 VSS 0.18811f
C7281 C10_N_btm.t990 VSS 0.18811f
C7282 C10_N_btm.t231 VSS 0.18811f
C7283 C10_N_btm.t939 VSS 0.18811f
C7284 C10_N_btm.t492 VSS 0.18811f
C7285 C10_N_btm.t334 VSS 0.18811f
C7286 C10_N_btm.t63 VSS 0.18811f
C7287 C10_N_btm.t280 VSS 0.18811f
C7288 C10_N_btm.t1026 VSS 0.18811f
C7289 C10_N_btm.t491 VSS 0.18811f
C7290 C10_N_btm.t444 VSS 0.18811f
C7291 C10_N_btm.t175 VSS 0.18811f
C7292 C10_N_btm.t432 VSS 0.18811f
C7293 C10_N_btm.t672 VSS 0.18811f
C7294 C10_N_btm.t336 VSS 0.18811f
C7295 C10_N_btm.t553 VSS 0.18811f
C7296 C10_N_btm.t849 VSS 0.18811f
C7297 C10_N_btm.t504 VSS 0.18811f
C7298 C10_N_btm.t737 VSS 0.18811f
C7299 C10_N_btm.t445 VSS 0.18811f
C7300 C10_N_btm.t688 VSS 0.18811f
C7301 C10_N_btm.t919 VSS 0.18811f
C7302 C10_N_btm.t626 VSS 0.18811f
C7303 C10_N_btm.t869 VSS 0.18811f
C7304 C10_N_btm.t114 VSS 0.18811f
C7305 C10_N_btm.t754 VSS 0.18811f
C7306 C10_N_btm.t812 VSS 0.18811f
C7307 C10_N_btm.t696 VSS 0.18811f
C7308 C10_N_btm.t936 VSS 0.18811f
C7309 C10_N_btm.t170 VSS 0.18811f
C7310 C10_N_btm.t879 VSS 0.18811f
C7311 C10_N_btm.t61 VSS 0.18811f
C7312 C10_N_btm.t329 VSS 0.18811f
C7313 C10_N_btm.t117 VSS 0.208624f
C7314 C10_N_btm.t964 VSS 0.208624f
C7315 C10_N_btm.t620 VSS 0.18811f
C7316 C10_N_btm.t1023 VSS 0.18811f
C7317 C10_N_btm.t787 VSS 0.18811f
C7318 C10_N_btm.t72 VSS 0.18811f
C7319 C10_N_btm.t839 VSS 0.18811f
C7320 C10_N_btm.t602 VSS 0.18811f
C7321 C10_N_btm.t947 VSS 0.18811f
C7322 C10_N_btm.t660 VSS 0.18811f
C7323 C10_N_btm.t1002 VSS 0.18811f
C7324 C10_N_btm.t768 VSS 0.18811f
C7325 C10_N_btm.t524 VSS 0.18811f
C7326 C10_N_btm.t818 VSS 0.18811f
C7327 C10_N_btm.t582 VSS 0.18811f
C7328 C10_N_btm.t353 VSS 0.18811f
C7329 C10_N_btm.t643 VSS 0.18811f
C7330 C10_N_btm.t405 VSS 0.18811f
C7331 C10_N_btm.t749 VSS 0.18811f
C7332 C10_N_btm.t460 VSS 0.18811f
C7333 C10_N_btm.t1031 VSS 0.18811f
C7334 C10_N_btm.t566 VSS 0.18811f
C7335 C10_N_btm.t344 VSS 0.18811f
C7336 C10_N_btm.t77 VSS 0.18811f
C7337 C10_N_btm.t352 VSS 0.18811f
C7338 C10_N_btm.t142 VSS 0.18811f
C7339 C10_N_btm.t911 VSS 0.18811f
C7340 C10_N_btm.t192 VSS 0.18811f
C7341 C10_N_btm.t1037 VSS 0.18811f
C7342 C10_N_btm.t1013 VSS 0.18811f
C7343 C10_N_btm.t238 VSS 0.18811f
C7344 C10_N_btm.t842 VSS 0.18811f
C7345 C10_N_btm.t128 VSS 0.18811f
C7346 C10_N_btm.t891 VSS 0.18811f
C7347 C10_N_btm.t665 VSS 0.18811f
C7348 C10_N_btm.t1010 VSS 0.18811f
C7349 C10_N_btm.t708 VSS 0.18811f
C7350 C10_N_btm.t41 VSS 0.18811f
C7351 C10_N_btm.t823 VSS 0.18811f
C7352 C10_N_btm.t529 VSS 0.18811f
C7353 C10_N_btm.t880 VSS 0.18811f
C7354 C10_N_btm.t648 VSS 0.18811f
C7355 C10_N_btm.t411 VSS 0.18811f
C7356 C10_N_btm.t697 VSS 0.18811f
C7357 C10_N_btm.t465 VSS 0.18811f
C7358 C10_N_btm.t809 VSS 0.18811f
C7359 C10_N_btm.t1050 VSS 0.18811f
C7360 C10_N_btm.t143 VSS 0.18811f
C7361 C10_N_btm.t627 VSS 0.18811f
C7362 C10_N_btm.t348 VSS 0.18811f
C7363 C10_N_btm.t133 VSS 0.18811f
C7364 C10_N_btm.t788 VSS 0.18811f
C7365 C10_N_btm.t541 VSS 0.18811f
C7366 C10_N_btm.t275 VSS 0.18811f
C7367 C10_N_btm.t606 VSS 0.18811f
C7368 C10_N_btm.t378 VSS 0.18811f
C7369 C10_N_btm.t666 VSS 0.18811f
C7370 C10_N_btm.t427 VSS 0.18811f
C7371 C10_N_btm.t217 VSS 0.18811f
C7372 C10_N_btm.t510 VSS 0.18811f
C7373 C10_N_btm.t266 VSS 0.18811f
C7374 C10_N_btm.t89 VSS 0.18811f
C7375 C10_N_btm.t358 VSS 0.18811f
C7376 C10_N_btm.t108 VSS 0.18811f
C7377 C10_N_btm.t414 VSS 0.208624f
C7378 C10_N_btm.t637 VSS 0.18811f
C7379 C10_N_btm.t579 VSS 0.208624f
C7380 C10_N_btm.t261 VSS 0.18811f
C7381 C10_N_btm.t522 VSS 0.18811f
C7382 C10_N_btm.t204 VSS 0.18811f
C7383 C10_N_btm.t425 VSS 0.18811f
C7384 C10_N_btm.t658 VSS 0.18811f
C7385 C10_N_btm.t371 VSS 0.18811f
C7386 C10_N_btm.t294 VSS 0.18811f
C7387 C10_N_btm.t836 VSS 0.18811f
C7388 C10_N_btm.t537 VSS 0.18811f
C7389 C10_N_btm.t784 VSS 0.18811f
C7390 C10_N_btm.t436 VSS 0.18811f
C7391 C10_N_btm.t715 VSS 0.18811f
C7392 C10_N_btm.t961 VSS 0.18811f
C7393 C10_N_btm.t382 VSS 0.18811f
C7394 C10_N_btm.t609 VSS 0.18811f
C7395 C10_N_btm.t896 VSS 0.18811f
C7396 C10_N_btm.t545 VSS 0.18811f
C7397 C10_N_btm.t790 VSS 0.18811f
C7398 C10_N_btm.t1034 VSS 0.18811f
C7399 C10_N_btm.t730 VSS 0.18811f
C7400 C10_N_btm.t968 VSS 0.18811f
C7401 C10_N_btm.t680 VSS 0.18811f
C7402 C10_N_btm.t916 VSS 0.18811f
C7403 C10_N_btm.t107 VSS 0.18811f
C7404 C10_N_btm.t803 VSS 0.18811f
C7405 C10_N_btm.t56 VSS 0.18811f
C7406 C10_N_btm.t265 VSS 0.18811f
C7407 C10_N_btm.t985 VSS 0.18811f
C7408 C10_N_btm.t211 VSS 0.18811f
C7409 C10_N_btm.t931 VSS 0.18811f
C7410 C10_N_btm.t229 VSS 0.18811f
C7411 C10_N_btm.t375 VSS 0.18811f
C7412 C10_N_btm.t57 VSS 0.18811f
C7413 C10_N_btm.t272 VSS 0.18811f
C7414 C10_N_btm.t905 VSS 0.18811f
C7415 C10_N_btm.t243 VSS 0.18811f
C7416 C10_N_btm.t439 VSS 0.18811f
C7417 C10_N_btm.t121 VSS 0.18811f
C7418 C10_N_btm.t387 VSS 0.18811f
C7419 C10_N_btm.t617 VSS 0.18811f
C7420 C10_N_btm.t325 VSS 0.18811f
C7421 C10_N_btm.t604 VSS 0.18811f
C7422 C10_N_btm.t843 VSS 0.18811f
C7423 C10_N_btm.t974 VSS 0.18811f
C7424 C10_N_btm.t724 VSS 0.18811f
C7425 C10_N_btm.t48 VSS 0.18811f
C7426 C10_N_btm.t677 VSS 0.18811f
C7427 C10_N_btm.t912 VSS 0.18811f
C7428 C10_N_btm.t618 VSS 0.18811f
C7429 C10_N_btm.t858 VSS 0.18811f
C7430 C10_N_btm.t50 VSS 0.18811f
C7431 C10_N_btm.t394 VSS 0.18811f
C7432 C10_N_btm.t1055 VSS 0.18811f
C7433 C10_N_btm.t205 VSS 0.18811f
C7434 C10_N_btm.t928 VSS 0.18811f
C7435 C10_N_btm.t162 VSS 0.18811f
C7436 C10_N_btm.t872 VSS 0.18811f
C7437 C10_N_btm.t516 VSS 0.18811f
C7438 C10_N_btm.t321 VSS 0.18811f
C7439 C10_N_btm.t361 VSS 0.18811f
C7440 C10_N_btm.t239 VSS 0.18811f
C7441 C10_N_btm.t757 VSS 0.18811f
C7442 C10_N_btm.t177 VSS 0.208624f
C7443 C10_N_btm.t1044 VSS 0.208624f
C7444 C10_N_btm.t861 VSS 0.18811f
C7445 C10_N_btm.t563 VSS 0.18811f
C7446 C10_N_btm.t342 VSS 0.18811f
C7447 C10_N_btm.t679 VSS 0.18811f
C7448 C10_N_btm.t389 VSS 0.18811f
C7449 C10_N_btm.t179 VSS 0.18811f
C7450 C10_N_btm.t1012 VSS 0.18811f
C7451 C10_N_btm.t474 VSS 0.18811f
C7452 C10_N_btm.t543 VSS 0.18811f
C7453 C10_N_btm.t327 VSS 0.18811f
C7454 C10_N_btm.t233 VSS 0.18811f
C7455 C10_N_btm.t379 VSS 0.18811f
C7456 C10_N_btm.t167 VSS 0.18811f
C7457 C10_N_btm.t987 VSS 0.18811f
C7458 C10_N_btm.t224 VSS 0.18811f
C7459 C10_N_btm.t924 VSS 0.18811f
C7460 C10_N_btm.t314 VSS 0.18811f
C7461 C10_N_btm.t102 VSS 0.18811f
C7462 C10_N_btm.t867 VSS 0.18811f
C7463 C10_N_btm.t154 VSS 0.18811f
C7464 C10_N_btm.t969 VSS 0.18811f
C7465 C10_N_btm.t686 VSS 0.18811f
C7466 C10_N_btm.t986 VSS 0.18811f
C7467 C10_N_btm.t747 VSS 0.18811f
C7468 C10_N_btm.t457 VSS 0.18811f
C7469 C10_N_btm.t804 VSS 0.18811f
C7470 C10_N_btm.t564 VSS 0.18811f
C7471 C10_N_btm.t865 VSS 0.18811f
C7472 C10_N_btm.t622 VSS 0.18811f
C7473 C10_N_btm.t392 VSS 0.18811f
C7474 C10_N_btm.t732 VSS 0.18811f
C7475 C10_N_btm.t443 VSS 0.18811f
C7476 C10_N_btm.t488 VSS 0.18811f
C7477 C10_N_btm.t547 VSS 0.18811f
C7478 C10_N_btm.t279 VSS 0.18811f
C7479 C10_N_btm.t611 VSS 0.18811f
C7480 C10_N_btm.t1039 VSS 0.18811f
C7481 C10_N_btm.t485 VSS 0.18811f
C7482 C10_N_btm.t431 VSS 0.18811f
C7483 C10_N_btm.t228 VSS 0.18811f
C7484 C10_N_btm.t793 VSS 0.18811f
C7485 C10_N_btm.t268 VSS 0.18811f
C7486 C10_N_btm.t220 VSS 0.18811f
C7487 C10_N_btm.t365 VSS 0.18811f
C7488 C10_N_btm.t119 VSS 0.18811f
C7489 C10_N_btm.t922 VSS 0.18811f
C7490 C10_N_btm.t201 VSS 0.18811f
C7491 C10_N_btm.t976 VSS 0.18811f
C7492 C10_N_btm.t741 VSS 0.18811f
C7493 C10_N_btm.t440 VSS 0.18811f
C7494 C10_N_btm.t471 VSS 0.18811f
C7495 C10_N_btm.t1011 VSS 0.18811f
C7496 C10_N_btm.t276 VSS 0.18811f
C7497 C10_N_btm.t59 VSS 0.18811f
C7498 C10_N_btm.t330 VSS 0.18811f
C7499 C10_N_btm.t241 VSS 0.18811f
C7500 C10_N_btm.t935 VSS 0.18811f
C7501 C10_N_btm.t171 VSS 0.18811f
C7502 C10_N_btm.t989 VSS 0.18811f
C7503 C10_N_btm.t753 VSS 0.18811f
C7504 C10_N_btm.t93 VSS 0.18811f
C7505 C10_N_btm.t808 VSS 0.18811f
C7506 C10_N_btm.t112 VSS 0.208624f
C7507 C10_N_btm.t417 VSS 0.18811f
C7508 C10_N_btm.t370 VSS 0.208624f
C7509 C10_N_btm.t476 VSS 0.18811f
C7510 C10_N_btm.t320 VSS 0.18811f
C7511 C10_N_btm.t738 VSS 0.18811f
C7512 C10_N_btm.t234 VSS 0.18811f
C7513 C10_N_btm.t433 VSS 0.18811f
C7514 C10_N_btm.t174 VSS 0.18811f
C7515 C10_N_btm.t384 VSS 0.18811f
C7516 C10_N_btm.t613 VSS 0.18811f
C7517 C10_N_btm.t335 VSS 0.18811f
C7518 C10_N_btm.t550 VSS 0.208624f
C7519 C10_N_btm.t73 VSS 0.208624f
C7520 C10_N_btm.t888 VSS 0.18811f
C7521 C10_N_btm.t124 VSS 0.18811f
C7522 C10_N_btm.t948 VSS 0.18811f
C7523 C10_N_btm.t705 VSS 0.18811f
C7524 C10_N_btm.t1004 VSS 0.18811f
C7525 C10_N_btm.t769 VSS 0.18811f
C7526 C10_N_btm.t525 VSS 0.18811f
C7527 C10_N_btm.t874 VSS 0.18811f
C7528 C10_N_btm.t583 VSS 0.18811f
C7529 C10_N_btm.t932 VSS 0.208624f
C7530 C10_N_btm.t215 VSS 0.18811f
C7531 C10_N_btm.t512 VSS 0.208624f
C7532 C10_N_btm.t172 VSS 0.18811f
C7533 C10_N_btm.t428 VSS 0.18811f
C7534 C10_N_btm.t244 VSS 0.18811f
C7535 C10_N_btm.t331 VSS 0.18811f
C7536 C10_N_btm.t546 VSS 0.18811f
C7537 C10_N_btm.t277 VSS 0.18811f
C7538 C10_N_btm.t1027 VSS 0.18811f
C7539 C10_N_btm.t731 VSS 0.18811f
C7540 C10_N_btm.t441 VSS 0.18811f
C7541 C10_N_btm.t681 VSS 0.208624f
C7542 C10_N_btm.t293 VSS 0.208624f
C7543 C10_N_btm.t81 VSS 0.18811f
C7544 C10_N_btm.t347 VSS 0.18811f
C7545 C10_N_btm.t132 VSS 0.18811f
C7546 C10_N_btm.t957 VSS 0.18811f
C7547 C10_N_btm.t184 VSS 0.18811f
C7548 C10_N_btm.t1017 VSS 0.18811f
C7549 C10_N_btm.t779 VSS 0.18811f
C7550 C10_N_btm.t65 VSS 0.18811f
C7551 C10_N_btm.t829 VSS 0.18811f
C7552 C10_N_btm.t500 VSS 0.208624f
C7553 C10_N_btm.t434 VSS 0.18811f
C7554 C10_N_btm.t273 VSS 0.208624f
C7555 C10_N_btm.t1006 VSS 0.18811f
C7556 C10_N_btm.t467 VSS 0.18811f
C7557 C10_N_btm.t950 VSS 0.18811f
C7558 C10_N_btm.t126 VSS 0.18811f
C7559 C10_N_btm.t341 VSS 0.18811f
C7560 C10_N_btm.t75 VSS 0.18811f
C7561 C10_N_btm.t286 VSS 0.18811f
C7562 C10_N_btm.t1042 VSS 0.18811f
C7563 C10_N_btm.t906 VSS 0.18811f
C7564 C10_N_btm.t454 VSS 0.208624f
C7565 C10_N_btm.t104 VSS 0.208624f
C7566 C10_N_btm.t914 VSS 0.18811f
C7567 C10_N_btm.t147 VSS 0.18811f
C7568 C10_N_btm.t965 VSS 0.18811f
C7569 C10_N_btm.t727 VSS 0.18811f
C7570 C10_N_btm.t223 VSS 0.18811f
C7571 C10_N_btm.t789 VSS 0.18811f
C7572 C10_N_btm.t542 VSS 0.18811f
C7573 C10_N_btm.t893 VSS 0.18811f
C7574 C10_N_btm.t607 VSS 0.18811f
C7575 C10_N_btm.t953 VSS 0.208624f
C7576 C10_N_btm.t993 VSS 0.18811f
C7577 C10_N_btm.t70 VSS 0.208624f
C7578 C10_N_btm.t785 VSS 0.18811f
C7579 C10_N_btm.t86 VSS 0.18811f
C7580 C10_N_btm.t717 VSS 0.18811f
C7581 C10_N_btm.t962 VSS 0.18811f
C7582 C10_N_btm.t135 VSS 0.18811f
C7583 C10_N_btm.t907 VSS 0.18811f
C7584 C10_N_btm.t88 VSS 0.18811f
C7585 C10_N_btm.t301 VSS 0.18811f
C7586 C10_N_btm.t44 VSS 0.18811f
C7587 C10_N_btm.t256 VSS 0.208624f
C7588 C10_N_btm.t927 VSS 0.208624f
C7589 C10_N_btm.t693 VSS 0.18811f
C7590 C10_N_btm.t981 VSS 0.18811f
C7591 C10_N_btm.t744 VSS 0.18811f
C7592 C10_N_btm.t1040 VSS 0.18811f
C7593 C10_N_btm.t798 VSS 0.18811f
C7594 C10_N_btm.t560 VSS 0.18811f
C7595 C10_N_btm.t339 VSS 0.18811f
C7596 C10_N_btm.t676 VSS 0.18811f
C7597 C10_N_btm.t1052 VSS 0.18811f
C7598 C10_N_btm.t723 VSS 0.208624f
C7599 C10_N_btm.t956 VSS 0.18811f
C7600 C10_N_btm.t902 VSS 0.208624f
C7601 C10_N_btm.t551 VSS 0.18811f
C7602 C10_N_btm.t848 VSS 0.18811f
C7603 C10_N_btm.t503 VSS 0.18811f
C7604 C10_N_btm.t735 VSS 0.18811f
C7605 C10_N_btm.t971 VSS 0.18811f
C7606 C10_N_btm.t687 VSS 0.18811f
C7607 C10_N_btm.t918 VSS 0.18811f
C7608 C10_N_btm.t113 VSS 0.18811f
C7609 C10_N_btm.t868 VSS 0.18811f
C7610 C10_N_btm.t106 VSS 0.208624f
C7611 C10_N_btm.t576 VSS 0.208624f
C7612 C10_N_btm.t350 VSS 0.18811f
C7613 C10_N_btm.t638 VSS 0.18811f
C7614 C10_N_btm.t401 VSS 0.18811f
C7615 C10_N_btm.t188 VSS 0.18811f
C7616 C10_N_btm.t452 VSS 0.18811f
C7617 C10_N_btm.t773 VSS 0.18811f
C7618 C10_N_btm.t103 VSS 0.18811f
C7619 C10_N_btm.t340 VSS 0.18811f
C7620 C10_N_btm.t74 VSS 0.18811f
C7621 C10_N_btm.t1053 VSS 0.208624f
C7622 C10_N_btm.t726 VSS 0.18811f
C7623 C10_N_btm.t684 VSS 0.208624f
C7624 C10_N_btm.t345 VSS 0.18811f
C7625 C10_N_btm.t623 VSS 0.18811f
C7626 C10_N_btm.t287 VSS 0.18811f
C7627 C10_N_btm.t1048 VSS 0.18811f
C7628 C10_N_btm.t751 VSS 0.18811f
C7629 C10_N_btm.t459 VSS 0.18811f
C7630 C10_N_btm.t694 VSS 0.18811f
C7631 C10_N_btm.t933 VSS 0.18811f
C7632 C10_N_btm.t642 VSS 0.18811f
C7633 C10_N_btm.t876 VSS 0.208624f
C7634 C10_N_btm.t364 VSS 0.208624f
C7635 C10_N_btm.t157 VSS 0.18811f
C7636 C10_N_btm.t420 VSS 0.18811f
C7637 C10_N_btm.t200 VSS 0.18811f
C7638 C10_N_btm.t39 VSS 0.18811f
C7639 C10_N_btm.t255 VSS 0.18811f
C7640 C10_N_btm.t42 VSS 0.18811f
C7641 C10_N_btm.t852 VSS 0.18811f
C7642 C10_N_btm.t134 VSS 0.18811f
C7643 C10_N_btm.t904 VSS 0.18811f
C7644 C10_N_btm.t187 VSS 0.208624f
C7645 C10_N_btm.t1038 VSS 0.18811f
C7646 C10_N_btm.t346 VSS 0.208624f
C7647 C10_N_btm.t517 VSS 0.18811f
C7648 C10_N_btm.t288 VSS 0.18811f
C7649 C10_N_btm.t1036 VSS 0.18811f
C7650 C10_N_btm.t193 VSS 0.18811f
C7651 C10_N_btm.t409 VSS 0.18811f
C7652 C10_N_btm.t148 VSS 0.18811f
C7653 C10_N_btm.t354 VSS 0.18811f
C7654 C10_N_btm.t587 VSS 0.18811f
C7655 C10_N_btm.t308 VSS 0.18811f
C7656 C10_N_btm.t526 VSS 0.208624f
C7657 C10_N_btm.t322 VSS 0.208624f
C7658 C10_N_btm.t570 VSS 0.18811f
C7659 C10_N_btm.t251 VSS 0.18811f
C7660 C10_N_btm.t472 VSS 0.18811f
C7661 C10_N_btm.t700 VSS 0.18811f
C7662 C10_N_btm.t415 VSS 0.18811f
C7663 C10_N_btm.t650 VSS 0.18811f
C7664 C10_N_btm.t881 VSS 0.18811f
C7665 C10_N_btm.t590 VSS 0.18811f
C7666 C10_N_btm.t825 VSS 0.208624f
C7667 C10_N_btm.t168 VSS 0.208624f
C7668 C10_N_btm.t988 VSS 0.18811f
C7669 C10_N_btm.t218 VSS 0.18811f
C7670 C10_N_btm.t920 VSS 0.18811f
C7671 C10_N_btm.t807 VSS 0.18811f
C7672 C10_N_btm.t99 VSS 0.18811f
C7673 C10_N_btm.t866 VSS 0.18811f
C7674 C10_N_btm.t625 VSS 0.18811f
C7675 C10_N_btm.t970 VSS 0.18811f
C7676 C10_N_btm.t685 VSS 0.18811f
C7677 C10_N_btm.t222 VSS 0.208624f
C7678 C10_N_btm.t297 VSS 0.18811f
C7679 C10_N_btm.t145 VSS 0.208624f
C7680 C10_N_btm.t859 VSS 0.18811f
C7681 C10_N_btm.t98 VSS 0.18811f
C7682 C10_N_btm.t799 VSS 0.18811f
C7683 C10_N_btm.t994 VSS 0.18811f
C7684 C10_N_btm.t206 VSS 0.18811f
C7685 C10_N_btm.t982 VSS 0.18811f
C7686 C10_N_btm.t163 VSS 0.18811f
C7687 C10_N_btm.t373 VSS 0.18811f
C7688 C10_N_btm.t219 VSS 0.18811f
C7689 C10_N_btm.t1001 VSS 0.208624f
C7690 C10_N_btm.t766 VSS 0.18811f
C7691 C10_N_btm.t515 VSS 0.18811f
C7692 C10_N_btm.t817 VSS 0.18811f
C7693 C10_N_btm.t581 VSS 0.18811f
C7694 C10_N_btm.t875 VSS 0.18811f
C7695 C10_N_btm.t641 VSS 0.18811f
C7696 C10_N_btm.t404 VSS 0.18811f
C7697 C10_N_btm.t748 VSS 0.18811f
C7698 C10_N_btm.t458 VSS 0.18811f
C7699 C10_N_btm.t805 VSS 0.208624f
C7700 C10_N_btm.t36 VSS 0.18811f
C7701 C10_N_btm.t252 VSS 0.18811f
C7702 C10_N_btm.t973 VSS 0.18811f
C7703 C10_N_btm.t156 VSS 0.18811f
C7704 C10_N_btm.t363 VSS 0.18811f
C7705 C10_N_btm.t115 VSS 0.18811f
C7706 C10_N_btm.t316 VSS 0.18811f
C7707 C10_N_btm.t533 VSS 0.18811f
C7708 C10_N_btm.t267 VSS 0.18811f
C7709 C10_N_btm.t513 VSS 0.208624f
C7710 C10_N_btm.t1075 VSS 0.208975f
C7711 C10_N_btm.n3897 VSS 0.100561f
C7712 a_n1522_42718.t4 VSS 1.6089f
C7713 a_n1522_42718.n1 VSS 11.891701f
C7714 C10_P_btm.n0 VSS 0.147281f
C7715 C10_P_btm.n1 VSS 0.142447f
C7716 C10_P_btm.n2 VSS 0.448098f
C7717 C10_P_btm.n3 VSS 0.142447f
C7718 C10_P_btm.n4 VSS 0.230043f
C7719 C10_P_btm.n5 VSS 0.142447f
C7720 C10_P_btm.n6 VSS 0.230043f
C7721 C10_P_btm.n7 VSS 0.142447f
C7722 C10_P_btm.n8 VSS 0.230043f
C7723 C10_P_btm.n9 VSS 0.142447f
C7724 C10_P_btm.n10 VSS 0.230043f
C7725 C10_P_btm.n11 VSS 0.142447f
C7726 C10_P_btm.n12 VSS 0.229719f
C7727 C10_P_btm.n13 VSS 0.142447f
C7728 C10_P_btm.n14 VSS 0.395441f
C7729 C10_P_btm.n15 VSS 0.216437f
C7730 C10_P_btm.n16 VSS 0.21129f
C7731 C10_P_btm.n17 VSS 0.31695f
C7732 C10_P_btm.n18 VSS 0.21129f
C7733 C10_P_btm.n19 VSS 0.16285f
C7734 C10_P_btm.n20 VSS 0.21129f
C7735 C10_P_btm.n21 VSS 0.184948f
C7736 C10_P_btm.n22 VSS 0.258762f
C7737 C10_P_btm.n23 VSS 0.25913f
C7738 C10_P_btm.n24 VSS 0.220601f
C7739 C10_P_btm.n25 VSS 0.213709f
C7740 C10_P_btm.n26 VSS 0.218928f
C7741 C10_P_btm.n27 VSS 0.213709f
C7742 C10_P_btm.n28 VSS 0.323009f
C7743 C10_P_btm.n29 VSS 0.213709f
C7744 C10_P_btm.n30 VSS 0.166325f
C7745 C10_P_btm.n31 VSS 0.186482f
C7746 C10_P_btm.n32 VSS 0.93945f
C7747 C10_P_btm.t19 VSS 0.216875f
C7748 C10_P_btm.t24 VSS 0.216875f
C7749 C10_P_btm.t21 VSS 0.216875f
C7750 C10_P_btm.t13 VSS 0.216875f
C7751 C10_P_btm.t14 VSS 0.216875f
C7752 C10_P_btm.t20 VSS 0.216875f
C7753 C10_P_btm.t25 VSS 0.216875f
C7754 C10_P_btm.t16 VSS 0.216875f
C7755 C10_P_btm.t23 VSS 0.216875f
C7756 C10_P_btm.t364 VSS 0.208624f
C7757 C10_P_btm.t72 VSS 0.208624f
C7758 C10_P_btm.t340 VSS 0.208624f
C7759 C10_P_btm.t111 VSS 0.18811f
C7760 C10_P_btm.t826 VSS 0.18811f
C7761 C10_P_btm.t894 VSS 0.18811f
C7762 C10_P_btm.t230 VSS 0.18811f
C7763 C10_P_btm.t1001 VSS 0.18811f
C7764 C10_P_btm.t169 VSS 0.18811f
C7765 C10_P_btm.t390 VSS 0.18811f
C7766 C10_P_btm.t483 VSS 0.18811f
C7767 C10_P_btm.t997 VSS 0.208624f
C7768 C10_P_btm.t122 VSS 0.208624f
C7769 C10_P_btm.t938 VSS 0.18811f
C7770 C10_P_btm.t606 VSS 0.18811f
C7771 C10_P_btm.t837 VSS 0.18811f
C7772 C10_P_btm.t266 VSS 0.18811f
C7773 C10_P_btm.t789 VSS 0.18811f
C7774 C10_P_btm.t1012 VSS 0.18811f
C7775 C10_P_btm.t179 VSS 0.18811f
C7776 C10_P_btm.t956 VSS 0.18811f
C7777 C10_P_btm.t786 VSS 0.208624f
C7778 C10_P_btm.t971 VSS 0.208624f
C7779 C10_P_btm.t727 VSS 0.18811f
C7780 C10_P_btm.t1039 VSS 0.18811f
C7781 C10_P_btm.t624 VSS 0.18811f
C7782 C10_P_btm.t848 VSS 0.18811f
C7783 C10_P_btm.t558 VSS 0.18811f
C7784 C10_P_btm.t800 VSS 0.18811f
C7785 C10_P_btm.t1020 VSS 0.18811f
C7786 C10_P_btm.t740 VSS 0.18811f
C7787 C10_P_btm.t556 VSS 0.208624f
C7788 C10_P_btm.t751 VSS 0.208624f
C7789 C10_P_btm.t503 VSS 0.18811f
C7790 C10_P_btm.t171 VSS 0.18811f
C7791 C10_P_btm.t393 VSS 0.18811f
C7792 C10_P_btm.t637 VSS 0.18811f
C7793 C10_P_btm.t345 VSS 0.18811f
C7794 C10_P_btm.t572 VSS 0.18811f
C7795 C10_P_btm.t812 VSS 0.18811f
C7796 C10_P_btm.t1052 VSS 0.18811f
C7797 C10_P_btm.t140 VSS 0.208624f
C7798 C10_P_btm.t328 VSS 0.208624f
C7799 C10_P_btm.t91 VSS 0.18811f
C7800 C10_P_btm.t817 VSS 0.18811f
C7801 C10_P_btm.t45 VSS 0.18811f
C7802 C10_P_btm.t210 VSS 0.18811f
C7803 C10_P_btm.t989 VSS 0.18811f
C7804 C10_P_btm.t158 VSS 0.18811f
C7805 C10_P_btm.t1041 VSS 0.18811f
C7806 C10_P_btm.t217 VSS 0.18811f
C7807 C10_P_btm.t404 VSS 0.208624f
C7808 C10_P_btm.t602 VSS 0.208624f
C7809 C10_P_btm.t354 VSS 0.18811f
C7810 C10_P_btm.t236 VSS 0.18811f
C7811 C10_P_btm.t250 VSS 0.18811f
C7812 C10_P_btm.t484 VSS 0.18811f
C7813 C10_P_btm.t194 VSS 0.18811f
C7814 C10_P_btm.t423 VSS 0.18811f
C7815 C10_P_btm.t655 VSS 0.18811f
C7816 C10_P_btm.t371 VSS 0.18811f
C7817 C10_P_btm.t526 VSS 0.208624f
C7818 C10_P_btm.t480 VSS 0.18811f
C7819 C10_P_btm.t138 VSS 0.18811f
C7820 C10_P_btm.t369 VSS 0.18811f
C7821 C10_P_btm.t600 VSS 0.18811f
C7822 C10_P_btm.t308 VSS 0.18811f
C7823 C10_P_btm.t541 VSS 0.18811f
C7824 C10_P_btm.t784 VSS 0.18811f
C7825 C10_P_btm.t629 VSS 0.18811f
C7826 C10_P_btm.t725 VSS 0.18811f
C7827 C10_P_btm.t1037 VSS 0.18811f
C7828 C10_P_btm.t674 VSS 0.18811f
C7829 C10_P_btm.t904 VSS 0.18811f
C7830 C10_P_btm.t350 VSS 0.18811f
C7831 C10_P_btm.t584 VSS 0.18811f
C7832 C10_P_btm.t869 VSS 0.18811f
C7833 C10_P_btm.t523 VSS 0.18811f
C7834 C10_P_btm.t760 VSS 0.18811f
C7835 C10_P_btm.t41 VSS 0.18811f
C7836 C10_P_btm.t707 VSS 0.18811f
C7837 C10_P_btm.t935 VSS 0.18811f
C7838 C10_P_btm.t653 VSS 0.18811f
C7839 C10_P_btm.t885 VSS 0.208624f
C7840 C10_P_btm.t749 VSS 0.208624f
C7841 C10_P_btm.t1023 VSS 0.208624f
C7842 C10_P_btm.t697 VSS 0.18811f
C7843 C10_P_btm.t355 VSS 0.18811f
C7844 C10_P_btm.t587 VSS 0.18811f
C7845 C10_P_btm.t821 VSS 0.18811f
C7846 C10_P_btm.t527 VSS 0.18811f
C7847 C10_P_btm.t764 VSS 0.18811f
C7848 C10_P_btm.t996 VSS 0.18811f
C7849 C10_P_btm.t711 VSS 0.18811f
C7850 C10_P_btm.t937 VSS 0.18811f
C7851 C10_P_btm.t604 VSS 0.18811f
C7852 C10_P_btm.t888 VSS 0.18811f
C7853 C10_P_btm.t513 VSS 0.18811f
C7854 C10_P_btm.t186 VSS 0.18811f
C7855 C10_P_btm.t410 VSS 0.18811f
C7856 C10_P_btm.t700 VSS 0.18811f
C7857 C10_P_btm.t358 VSS 0.18811f
C7858 C10_P_btm.t590 VSS 0.18811f
C7859 C10_P_btm.t879 VSS 0.18811f
C7860 C10_P_btm.t533 VSS 0.18811f
C7861 C10_P_btm.t772 VSS 0.18811f
C7862 C10_P_btm.t495 VSS 0.18811f
C7863 C10_P_btm.t716 VSS 0.18811f
C7864 C10_P_btm.t943 VSS 0.18811f
C7865 C10_P_btm.t611 VSS 0.18811f
C7866 C10_P_btm.t893 VSS 0.18811f
C7867 C10_P_btm.t62 VSS 0.18811f
C7868 C10_P_btm.t793 VSS 0.18811f
C7869 C10_P_btm.t490 VSS 0.18811f
C7870 C10_P_btm.t731 VSS 0.18811f
C7871 C10_P_btm.t959 VSS 0.18811f
C7872 C10_P_btm.t181 VSS 0.18811f
C7873 C10_P_btm.t909 VSS 0.18811f
C7874 C10_P_btm.t75 VSS 0.18811f
C7875 C10_P_btm.t294 VSS 0.18811f
C7876 C10_P_btm.t116 VSS 0.18811f
C7877 C10_P_btm.t248 VSS 0.18811f
C7878 C10_P_btm.t975 VSS 0.18811f
C7879 C10_P_btm.t192 VSS 0.18811f
C7880 C10_P_btm.t421 VSS 0.18811f
C7881 C10_P_btm.t126 VSS 0.18811f
C7882 C10_P_btm.t406 VSS 0.18811f
C7883 C10_P_btm.t644 VSS 0.18811f
C7884 C10_P_btm.t296 VSS 0.18811f
C7885 C10_P_btm.t529 VSS 0.18811f
C7886 C10_P_btm.t823 VSS 0.18811f
C7887 C10_P_btm.t488 VSS 0.18811f
C7888 C10_P_btm.t713 VSS 0.18811f
C7889 C10_P_btm.t425 VSS 0.18811f
C7890 C10_P_btm.t660 VSS 0.18811f
C7891 C10_P_btm.t890 VSS 0.18811f
C7892 C10_P_btm.t607 VSS 0.18811f
C7893 C10_P_btm.t838 VSS 0.18811f
C7894 C10_P_btm.t147 VSS 0.18811f
C7895 C10_P_btm.t730 VSS 0.18811f
C7896 C10_P_btm.t1018 VSS 0.18811f
C7897 C10_P_btm.t677 VSS 0.18811f
C7898 C10_P_btm.t908 VSS 0.18811f
C7899 C10_P_btm.t123 VSS 0.18811f
C7900 C10_P_btm.t851 VSS 0.18811f
C7901 C10_P_btm.t101 VSS 0.18811f
C7902 C10_P_btm.t291 VSS 0.18811f
C7903 C10_P_btm.t968 VSS 0.208624f
C7904 C10_P_btm.t857 VSS 0.208624f
C7905 C10_P_btm.t914 VSS 0.18811f
C7906 C10_P_btm.t571 VSS 0.18811f
C7907 C10_P_btm.t810 VSS 0.18811f
C7908 C10_P_btm.t46 VSS 0.18811f
C7909 C10_P_btm.t750 VSS 0.18811f
C7910 C10_P_btm.t981 VSS 0.18811f
C7911 C10_P_btm.t149 VSS 0.18811f
C7912 C10_P_btm.t926 VSS 0.18811f
C7913 C10_P_btm.t106 VSS 0.18811f
C7914 C10_P_btm.t825 VSS 0.18811f
C7915 C10_P_btm.t100 VSS 0.18811f
C7916 C10_P_btm.t269 VSS 0.18811f
C7917 C10_P_btm.t108 VSS 0.18811f
C7918 C10_P_btm.t1030 VSS 0.18811f
C7919 C10_P_btm.t524 VSS 0.18811f
C7920 C10_P_btm.t190 VSS 0.18811f
C7921 C10_P_btm.t418 VSS 0.18811f
C7922 C10_P_btm.t708 VSS 0.18811f
C7923 C10_P_btm.t367 VSS 0.18811f
C7924 C10_P_btm.t598 VSS 0.18811f
C7925 C10_P_btm.t306 VSS 0.18811f
C7926 C10_P_btm.t539 VSS 0.18811f
C7927 C10_P_btm.t782 VSS 0.18811f
C7928 C10_P_btm.t441 VSS 0.18811f
C7929 C10_P_btm.t723 VSS 0.18811f
C7930 C10_P_btm.t953 VSS 0.18811f
C7931 C10_P_btm.t621 VSS 0.18811f
C7932 C10_P_btm.t902 VSS 0.18811f
C7933 C10_P_btm.t555 VSS 0.18811f
C7934 C10_P_btm.t798 VSS 0.18811f
C7935 C10_P_btm.t531 VSS 0.18811f
C7936 C10_P_btm.t738 VSS 0.18811f
C7937 C10_P_btm.t969 VSS 0.18811f
C7938 C10_P_btm.t132 VSS 0.18811f
C7939 C10_P_btm.t915 VSS 0.18811f
C7940 C10_P_btm.t86 VSS 0.18811f
C7941 C10_P_btm.t811 VSS 0.18811f
C7942 C10_P_btm.t33 VSS 0.18811f
C7943 C10_P_btm.t254 VSS 0.18811f
C7944 C10_P_btm.t1022 VSS 0.18811f
C7945 C10_P_btm.t630 VSS 0.18811f
C7946 C10_P_btm.t471 VSS 0.18811f
C7947 C10_P_btm.t135 VSS 0.18811f
C7948 C10_P_btm.t365 VSS 0.18811f
C7949 C10_P_btm.t650 VSS 0.18811f
C7950 C10_P_btm.t304 VSS 0.18811f
C7951 C10_P_btm.t537 VSS 0.18811f
C7952 C10_P_btm.t256 VSS 0.18811f
C7953 C10_P_btm.t516 VSS 0.18811f
C7954 C10_P_btm.t720 VSS 0.18811f
C7955 C10_P_btm.t436 VSS 0.18811f
C7956 C10_P_btm.t671 VSS 0.18811f
C7957 C10_P_btm.t900 VSS 0.18811f
C7958 C10_P_btm.t553 VSS 0.18811f
C7959 C10_P_btm.t846 VSS 0.18811f
C7960 C10_P_btm.t1029 VSS 0.18811f
C7961 C10_P_btm.t737 VSS 0.18811f
C7962 C10_P_btm.t1016 VSS 0.18811f
C7963 C10_P_btm.t687 VSS 0.18811f
C7964 C10_P_btm.t913 VSS 0.18811f
C7965 C10_P_btm.t130 VSS 0.18811f
C7966 C10_P_btm.t859 VSS 0.208624f
C7967 C10_P_btm.t840 VSS 0.18811f
C7968 C10_P_btm.t545 VSS 0.18811f
C7969 C10_P_btm.t316 VSS 0.18811f
C7970 C10_P_btm.t662 VSS 0.18811f
C7971 C10_P_btm.t89 VSS 0.18811f
C7972 C10_P_btm.t144 VSS 0.18811f
C7973 C10_P_btm.t493 VSS 0.18811f
C7974 C10_P_btm.t199 VSS 0.18811f
C7975 C10_P_btm.t1055 VSS 0.18811f
C7976 C10_P_btm.t297 VSS 0.18811f
C7977 C10_P_btm.t80 VSS 0.18811f
C7978 C10_P_btm.t356 VSS 0.18811f
C7979 C10_P_btm.t128 VSS 0.18811f
C7980 C10_P_btm.t963 VSS 0.18811f
C7981 C10_P_btm.t90 VSS 0.18811f
C7982 C10_P_btm.t1013 VSS 0.18811f
C7983 C10_P_btm.t283 VSS 0.18811f
C7984 C10_P_btm.t95 VSS 0.18811f
C7985 C10_P_btm.t843 VSS 0.18811f
C7986 C10_P_btm.t498 VSS 0.18811f
C7987 C10_P_btm.t947 VSS 0.18811f
C7988 C10_P_btm.t667 VSS 0.18811f
C7989 C10_P_btm.t960 VSS 0.18811f
C7990 C10_P_btm.t732 VSS 0.18811f
C7991 C10_P_btm.t450 VSS 0.18811f
C7992 C10_P_btm.t794 VSS 0.18811f
C7993 C10_P_btm.t547 VSS 0.18811f
C7994 C10_P_btm.t842 VSS 0.18811f
C7995 C10_P_btm.t612 VSS 0.18811f
C7996 C10_P_btm.t376 VSS 0.18811f
C7997 C10_P_btm.t717 VSS 0.18811f
C7998 C10_P_btm.t430 VSS 0.18811f
C7999 C10_P_btm.t201 VSS 0.18811f
C8000 C10_P_btm.t534 VSS 0.18811f
C8001 C10_P_btm.t253 VSS 0.18811f
C8002 C10_P_btm.t591 VSS 0.18811f
C8003 C10_P_btm.t359 VSS 0.18811f
C8004 C10_P_btm.t84 VSS 0.18811f
C8005 C10_P_btm.t411 VSS 0.18811f
C8006 C10_P_btm.t187 VSS 0.18811f
C8007 C10_P_btm.t1017 VSS 0.18811f
C8008 C10_P_btm.t501 VSS 0.18811f
C8009 C10_P_btm.t44 VSS 0.18811f
C8010 C10_P_btm.t347 VSS 0.18811f
C8011 C10_P_btm.t68 VSS 0.18811f
C8012 C10_P_btm.t901 VSS 0.18811f
C8013 C10_P_btm.t175 VSS 0.18811f
C8014 C10_P_btm.t952 VSS 0.18811f
C8015 C10_P_btm.t722 VSS 0.18811f
C8016 C10_P_btm.t785 VSS 0.18811f
C8017 C10_P_btm.t542 VSS 0.18811f
C8018 C10_P_btm.t259 VSS 0.18811f
C8019 C10_P_btm.t601 VSS 0.18811f
C8020 C10_P_btm.t370 VSS 0.18811f
C8021 C10_P_btm.t654 VSS 0.18811f
C8022 C10_P_btm.t422 VSS 0.18811f
C8023 C10_P_btm.t193 VSS 0.18811f
C8024 C10_P_btm.t481 VSS 0.18811f
C8025 C10_P_btm.t249 VSS 0.18811f
C8026 C10_P_btm.t219 VSS 0.18811f
C8027 C10_P_btm.t352 VSS 0.18811f
C8028 C10_P_btm.t76 VSS 0.18811f
C8029 C10_P_btm.t402 VSS 0.208624f
C8030 C10_P_btm.t636 VSS 0.18811f
C8031 C10_P_btm.t576 VSS 0.208624f
C8032 C10_P_btm.t511 VSS 0.18811f
C8033 C10_P_btm.t519 VSS 0.18811f
C8034 C10_P_btm.t188 VSS 0.18811f
C8035 C10_P_btm.t414 VSS 0.18811f
C8036 C10_P_btm.t647 VSS 0.18811f
C8037 C10_P_btm.t361 VSS 0.18811f
C8038 C10_P_btm.t594 VSS 0.18811f
C8039 C10_P_btm.t827 VSS 0.18811f
C8040 C10_P_btm.t535 VSS 0.18811f
C8041 C10_P_btm.t774 VSS 0.18811f
C8042 C10_P_btm.t434 VSS 0.18811f
C8043 C10_P_btm.t718 VSS 0.18811f
C8044 C10_P_btm.t945 VSS 0.18811f
C8045 C10_P_btm.t983 VSS 0.18811f
C8046 C10_P_btm.t155 VSS 0.18811f
C8047 C10_P_btm.t437 VSS 0.18811f
C8048 C10_P_btm.t113 VSS 0.18811f
C8049 C10_P_btm.t324 VSS 0.18811f
C8050 C10_P_btm.t618 VSS 0.18811f
C8051 C10_P_btm.t275 VSS 0.18811f
C8052 C10_P_btm.t502 VSS 0.18811f
C8053 C10_P_btm.t232 VSS 0.18811f
C8054 C10_P_btm.t455 VSS 0.18811f
C8055 C10_P_btm.t688 VSS 0.18811f
C8056 C10_P_btm.t343 VSS 0.18811f
C8057 C10_P_btm.t635 VSS 0.18811f
C8058 C10_P_btm.t858 VSS 0.18811f
C8059 C10_P_btm.t1050 VSS 0.18811f
C8060 C10_P_btm.t809 VSS 0.18811f
C8061 C10_P_btm.t463 VSS 0.18811f
C8062 C10_P_btm.t698 VSS 0.18811f
C8063 C10_P_btm.t980 VSS 0.18811f
C8064 C10_P_btm.t643 VSS 0.18811f
C8065 C10_P_btm.t876 VSS 0.18811f
C8066 C10_P_btm.t97 VSS 0.18811f
C8067 C10_P_btm.t820 VSS 0.18811f
C8068 C10_P_btm.t898 VSS 0.18811f
C8069 C10_P_btm.t712 VSS 0.18811f
C8070 C10_P_btm.t995 VSS 0.18811f
C8071 C10_P_btm.t166 VSS 0.18811f
C8072 C10_P_btm.t927 VSS 0.18811f
C8073 C10_P_btm.t150 VSS 0.18811f
C8074 C10_P_btm.t379 VSS 0.18811f
C8075 C10_P_btm.t112 VSS 0.18811f
C8076 C10_P_btm.t274 VSS 0.18811f
C8077 C10_P_btm.t550 VSS 0.18811f
C8078 C10_P_btm.t229 VSS 0.18811f
C8079 C10_P_btm.t453 VSS 0.18811f
C8080 C10_P_btm.t168 VSS 0.18811f
C8081 C10_P_btm.t389 VSS 0.18811f
C8082 C10_P_btm.t633 VSS 0.18811f
C8083 C10_P_btm.t337 VSS 0.18811f
C8084 C10_P_btm.t569 VSS 0.18811f
C8085 C10_P_btm.t807 VSS 0.18811f
C8086 C10_P_btm.t462 VSS 0.18811f
C8087 C10_P_btm.t746 VSS 0.18811f
C8088 C10_P_btm.t400 VSS 0.18811f
C8089 C10_P_btm.t642 VSS 0.18811f
C8090 C10_P_btm.t923 VSS 0.18811f
C8091 C10_P_btm.t585 VSS 0.18811f
C8092 C10_P_btm.t818 VSS 0.18811f
C8093 C10_P_btm.t54 VSS 0.18811f
C8094 C10_P_btm.t761 VSS 0.208624f
C8095 C10_P_btm.t672 VSS 0.208624f
C8096 C10_P_btm.t1003 VSS 0.18811f
C8097 C10_P_btm.t721 VSS 0.18811f
C8098 C10_P_btm.t517 VSS 0.18811f
C8099 C10_P_btm.t830 VSS 0.18811f
C8100 C10_P_btm.t538 VSS 0.18811f
C8101 C10_P_btm.t305 VSS 0.18811f
C8102 C10_P_btm.t651 VSS 0.18811f
C8103 C10_P_btm.t366 VSS 0.18811f
C8104 C10_P_btm.t705 VSS 0.18811f
C8105 C10_P_btm.t477 VSS 0.18811f
C8106 C10_P_btm.t769 VSS 0.18811f
C8107 C10_P_btm.t521 VSS 0.18811f
C8108 C10_P_btm.t289 VSS 0.18811f
C8109 C10_P_btm.t71 VSS 0.18811f
C8110 C10_P_btm.t349 VSS 0.18811f
C8111 C10_P_btm.t120 VSS 0.18811f
C8112 C10_P_btm.t459 VSS 0.18811f
C8113 C10_P_btm.t178 VSS 0.18811f
C8114 C10_P_btm.t1009 VSS 0.18811f
C8115 C10_P_btm.t280 VSS 0.18811f
C8116 C10_P_btm.t771 VSS 0.18811f
C8117 C10_P_btm.t834 VSS 0.18811f
C8118 C10_P_btm.t69 VSS 0.18811f
C8119 C10_P_btm.t903 VSS 0.18811f
C8120 C10_P_btm.t622 VSS 0.18811f
C8121 C10_P_btm.t954 VSS 0.18811f
C8122 C10_P_btm.t724 VSS 0.18811f
C8123 C10_P_btm.t1007 VSS 0.18811f
C8124 C10_P_btm.t783 VSS 0.18811f
C8125 C10_P_btm.t540 VSS 0.18811f
C8126 C10_P_btm.t886 VSS 0.18811f
C8127 C10_P_btm.t599 VSS 0.18811f
C8128 C10_P_btm.t368 VSS 0.18811f
C8129 C10_P_btm.t709 VSS 0.18811f
C8130 C10_P_btm.t419 VSS 0.18811f
C8131 C10_P_btm.t762 VSS 0.18811f
C8132 C10_P_btm.t525 VSS 0.18811f
C8133 C10_P_btm.t247 VSS 0.18811f
C8134 C10_P_btm.t586 VSS 0.18811f
C8135 C10_P_btm.t351 VSS 0.18811f
C8136 C10_P_btm.t124 VSS 0.18811f
C8137 C10_P_btm.t401 VSS 0.18811f
C8138 C10_P_btm.t180 VSS 0.18811f
C8139 C10_P_btm.t515 VSS 0.18811f
C8140 C10_P_btm.t486 VSS 0.18811f
C8141 C10_P_btm.t1031 VSS 0.18811f
C8142 C10_P_btm.t338 VSS 0.18811f
C8143 C10_P_btm.t61 VSS 0.18811f
C8144 C10_P_btm.t892 VSS 0.18811f
C8145 C10_P_btm.t554 VSS 0.18811f
C8146 C10_P_btm.t326 VSS 0.18811f
C8147 C10_P_btm.t119 VSS 0.18811f
C8148 C10_P_btm.t382 VSS 0.18811f
C8149 C10_P_btm.t157 VSS 0.18811f
C8150 C10_P_btm.t440 VSS 0.18811f
C8151 C10_P_btm.t207 VSS 0.18811f
C8152 C10_P_btm.t1034 VSS 0.18811f
C8153 C10_P_btm.t258 VSS 0.18811f
C8154 C10_P_btm.t42 VSS 0.18811f
C8155 C10_P_btm.t864 VSS 0.18811f
C8156 C10_P_btm.t136 VSS 0.18811f
C8157 C10_P_btm.t918 VSS 0.18811f
C8158 C10_P_btm.t189 VSS 0.208624f
C8159 C10_P_btm.t405 VSS 0.18811f
C8160 C10_P_btm.t360 VSS 0.208624f
C8161 C10_P_btm.t32 VSS 0.18811f
C8162 C10_P_btm.t299 VSS 0.18811f
C8163 C10_P_btm.t38 VSS 0.18811f
C8164 C10_P_btm.t202 VSS 0.18811f
C8165 C10_P_btm.t431 VSS 0.18811f
C8166 C10_P_btm.t148 VSS 0.18811f
C8167 C10_P_btm.t377 VSS 0.18811f
C8168 C10_P_btm.t613 VSS 0.18811f
C8169 C10_P_btm.t320 VSS 0.18811f
C8170 C10_P_btm.t548 VSS 0.18811f
C8171 C10_P_btm.t216 VSS 0.18811f
C8172 C10_P_btm.t965 VSS 0.18811f
C8173 C10_P_btm.t733 VSS 0.18811f
C8174 C10_P_btm.t102 VSS 0.18811f
C8175 C10_P_btm.t315 VSS 0.18811f
C8176 C10_P_btm.t608 VSS 0.18811f
C8177 C10_P_btm.t265 VSS 0.18811f
C8178 C10_P_btm.t768 VSS 0.18811f
C8179 C10_P_btm.t790 VSS 0.18811f
C8180 C10_P_btm.t447 VSS 0.18811f
C8181 C10_P_btm.t678 VSS 0.18811f
C8182 C10_P_btm.t1043 VSS 0.18811f
C8183 C10_P_btm.t627 VSS 0.18811f
C8184 C10_P_btm.t852 VSS 0.18811f
C8185 C10_P_btm.t508 VSS 0.18811f
C8186 C10_P_btm.t801 VSS 0.18811f
C8187 C10_P_btm.t1024 VSS 0.18811f
C8188 C10_P_btm.t691 VSS 0.18811f
C8189 C10_P_btm.t972 VSS 0.18811f
C8190 C10_P_btm.t640 VSS 0.18811f
C8191 C10_P_btm.t863 VSS 0.18811f
C8192 C10_P_btm.t85 VSS 0.18811f
C8193 C10_P_btm.t814 VSS 0.18811f
C8194 C10_P_btm.t476 VSS 0.18811f
C8195 C10_P_btm.t206 VSS 0.18811f
C8196 C10_P_btm.t984 VSS 0.18811f
C8197 C10_P_btm.t156 VSS 0.18811f
C8198 C10_P_btm.t881 VSS 0.18811f
C8199 C10_P_btm.t114 VSS 0.18811f
C8200 C10_P_btm.t325 VSS 0.18811f
C8201 C10_P_btm.t47 VSS 0.18811f
C8202 C10_P_btm.t309 VSS 0.18811f
C8203 C10_P_btm.t543 VSS 0.18811f
C8204 C10_P_btm.t208 VSS 0.18811f
C8205 C10_P_btm.t442 VSS 0.18811f
C8206 C10_P_btm.t726 VSS 0.18811f
C8207 C10_P_btm.t383 VSS 0.18811f
C8208 C10_P_btm.t623 VSS 0.18811f
C8209 C10_P_btm.t327 VSS 0.18811f
C8210 C10_P_btm.t557 VSS 0.18811f
C8211 C10_P_btm.t799 VSS 0.18811f
C8212 C10_P_btm.t504 VSS 0.18811f
C8213 C10_P_btm.t739 VSS 0.18811f
C8214 C10_P_btm.t970 VSS 0.18811f
C8215 C10_P_btm.t639 VSS 0.18811f
C8216 C10_P_btm.t916 VSS 0.18811f
C8217 C10_P_btm.t574 VSS 0.18811f
C8218 C10_P_btm.t813 VSS 0.18811f
C8219 C10_P_btm.t35 VSS 0.18811f
C8220 C10_P_btm.t755 VSS 0.18811f
C8221 C10_P_btm.t982 VSS 0.18811f
C8222 C10_P_btm.t203 VSS 0.18811f
C8223 C10_P_btm.t930 VSS 0.208624f
C8224 C10_P_btm.t98 VSS 0.208624f
C8225 C10_P_btm.t413 VSS 0.208624f
C8226 C10_P_btm.t615 VSS 0.208624f
C8227 C10_P_btm.t300 VSS 0.18811f
C8228 C10_P_btm.t593 VSS 0.18811f
C8229 C10_P_btm.t255 VSS 0.18811f
C8230 C10_P_btm.t499 VSS 0.18811f
C8231 C10_P_btm.t773 VSS 0.18811f
C8232 C10_P_btm.t433 VSS 0.18811f
C8233 C10_P_btm.t666 VSS 0.18811f
C8234 C10_P_btm.t944 VSS 0.18811f
C8235 C10_P_btm.t107 VSS 0.208624f
C8236 C10_P_btm.t472 VSS 0.208624f
C8237 C10_P_btm.t998 VSS 0.18811f
C8238 C10_P_btm.t225 VSS 0.18811f
C8239 C10_P_btm.t940 VSS 0.18811f
C8240 C10_P_btm.t246 VSS 0.18811f
C8241 C10_P_btm.t1051 VSS 0.18811f
C8242 C10_P_btm.t58 VSS 0.18811f
C8243 C10_P_btm.t281 VSS 0.18811f
C8244 C10_P_btm.t567 VSS 0.18811f
C8245 C10_P_btm.t933 VSS 0.208624f
C8246 C10_P_btm.t66 VSS 0.208624f
C8247 C10_P_btm.t833 VSS 0.18811f
C8248 C10_P_btm.t235 VSS 0.18811f
C8249 C10_P_btm.t780 VSS 0.18811f
C8250 C10_P_btm.t1006 VSS 0.18811f
C8251 C10_P_btm.t238 VSS 0.18811f
C8252 C10_P_btm.t950 VSS 0.18811f
C8253 C10_P_btm.t770 VSS 0.18811f
C8254 C10_P_btm.t395 VSS 0.18811f
C8255 C10_P_btm.t766 VSS 0.208624f
C8256 C10_P_btm.t957 VSS 0.208624f
C8257 C10_P_btm.t663 VSS 0.18811f
C8258 C10_P_btm.t941 VSS 0.18811f
C8259 C10_P_btm.t609 VSS 0.18811f
C8260 C10_P_btm.t841 VSS 0.18811f
C8261 C10_P_btm.t59 VSS 0.18811f
C8262 C10_P_btm.t791 VSS 0.18811f
C8263 C10_P_btm.t1027 VSS 0.18811f
C8264 C10_P_btm.t482 VSS 0.18811f
C8265 C10_P_btm.t596 VSS 0.208624f
C8266 C10_P_btm.t797 VSS 0.208624f
C8267 C10_P_btm.t522 VSS 0.18811f
C8268 C10_P_btm.t781 VSS 0.18811f
C8269 C10_P_btm.t439 VSS 0.18811f
C8270 C10_P_btm.t673 VSS 0.18811f
C8271 C10_P_btm.t951 VSS 0.18811f
C8272 C10_P_btm.t620 VSS 0.18811f
C8273 C10_P_btm.t847 VSS 0.18811f
C8274 C10_P_btm.t67 VSS 0.18811f
C8275 C10_P_btm.t426 VSS 0.208624f
C8276 C10_P_btm.t628 VSS 0.208624f
C8277 C10_P_btm.t318 VSS 0.18811f
C8278 C10_P_btm.t610 VSS 0.18811f
C8279 C10_P_btm.t268 VSS 0.18811f
C8280 C10_P_btm.t867 VSS 0.18811f
C8281 C10_P_btm.t792 VSS 0.18811f
C8282 C10_P_btm.t449 VSS 0.18811f
C8283 C10_P_btm.t679 VSS 0.18811f
C8284 C10_P_btm.t958 VSS 0.18811f
C8285 C10_P_btm.t10 VSS 0.216875f
C8286 C10_P_btm.t27 VSS 0.216875f
C8287 C10_P_btm.t12 VSS 0.216875f
C8288 C10_P_btm.t28 VSS 0.216875f
C8289 C10_P_btm.t22 VSS 0.216875f
C8290 C10_P_btm.t26 VSS 0.216875f
C8291 C10_P_btm.t31 VSS 0.216875f
C8292 C10_P_btm.t18 VSS 0.216875f
C8293 C10_P_btm.t15 VSS 0.216875f
C8294 C10_P_btm.t11 VSS 0.216875f
C8295 C10_P_btm.t464 VSS 0.208624f
C8296 C10_P_btm.t332 VSS 0.18811f
C8297 C10_P_btm.t491 VSS 0.18811f
C8298 C10_P_btm.t887 VSS 0.18811f
C8299 C10_P_btm.t162 VSS 0.18811f
C8300 C10_P_btm.t936 VSS 0.18811f
C8301 C10_P_btm.t710 VSS 0.18811f
C8302 C10_P_btm.t1053 VSS 0.18811f
C8303 C10_P_btm.t763 VSS 0.18811f
C8304 C10_P_btm.t29 VSS 0.216875f
C8305 C10_P_btm.t872 VSS 0.208624f
C8306 C10_P_btm.t87 VSS 0.18811f
C8307 C10_P_btm.t170 VSS 0.208624f
C8308 C10_P_btm.t392 VSS 0.18811f
C8309 C10_P_btm.t63 VSS 0.18811f
C8310 C10_P_btm.t342 VSS 0.18811f
C8311 C10_P_btm.t242 VSS 0.18811f
C8312 C10_P_btm.t489 VSS 0.18811f
C8313 C10_P_btm.t1048 VSS 0.18811f
C8314 C10_P_btm.t182 VSS 0.18811f
C8315 C10_P_btm.t403 VSS 0.18811f
C8316 C10_P_btm.t696 VSS 0.18811f
C8317 C10_P_btm.t353 VSS 0.208624f
C8318 C10_P_btm.t257 VSS 0.208624f
C8319 C10_P_btm.t597 VSS 0.18811f
C8320 C10_P_btm.t307 VSS 0.18811f
C8321 C10_P_btm.t88 VSS 0.18811f
C8322 C10_P_btm.t416 VSS 0.18811f
C8323 C10_P_btm.t137 VSS 0.18811f
C8324 C10_P_btm.t973 VSS 0.18811f
C8325 C10_P_btm.t966 VSS 0.18811f
C8326 C10_P_btm.t1025 VSS 0.18811f
C8327 C10_P_btm.t292 VSS 0.18811f
C8328 C10_P_btm.t73 VSS 0.208624f
C8329 C10_P_btm.t665 VSS 0.18811f
C8330 C10_P_btm.t329 VSS 0.208624f
C8331 C10_P_btm.t561 VSS 0.18811f
C8332 C10_P_btm.t244 VSS 0.18811f
C8333 C10_P_btm.t506 VSS 0.18811f
C8334 C10_P_btm.t176 VSS 0.18811f
C8335 C10_P_btm.t396 VSS 0.18811f
C8336 C10_P_btm.t690 VSS 0.18811f
C8337 C10_P_btm.t348 VSS 0.18811f
C8338 C10_P_btm.t575 VSS 0.18811f
C8339 C10_P_btm.t862 VSS 0.18811f
C8340 C10_P_btm.t1054 VSS 0.208624f
C8341 C10_P_btm.t427 VSS 0.208624f
C8342 C10_P_btm.t767 VSS 0.18811f
C8343 C10_P_btm.t496 VSS 0.18811f
C8344 C10_P_btm.t251 VSS 0.18811f
C8345 C10_P_btm.t588 VSS 0.18811f
C8346 C10_P_btm.t298 VSS 0.18811f
C8347 C10_P_btm.t82 VSS 0.18811f
C8348 C10_P_btm.t407 VSS 0.18811f
C8349 C10_P_btm.t131 VSS 0.18811f
C8350 C10_P_btm.t466 VSS 0.18811f
C8351 C10_P_btm.t494 VSS 0.208624f
C8352 C10_P_btm.t412 VSS 0.18811f
C8353 C10_P_btm.t1019 VSS 0.208624f
C8354 C10_P_btm.t736 VSS 0.18811f
C8355 C10_P_btm.t391 VSS 0.18811f
C8356 C10_P_btm.t685 VSS 0.18811f
C8357 C10_P_btm.t341 VSS 0.18811f
C8358 C10_P_btm.t570 VSS 0.18811f
C8359 C10_P_btm.t855 VSS 0.18811f
C8360 C10_P_btm.t1046 VSS 0.18811f
C8361 C10_P_btm.t748 VSS 0.18811f
C8362 C10_P_btm.t221 VSS 0.18811f
C8363 C10_P_btm.t695 VSS 0.208624f
C8364 C10_P_btm.t664 VSS 0.208624f
C8365 C10_P_btm.t323 VSS 0.18811f
C8366 C10_P_btm.t115 VSS 0.18811f
C8367 C10_P_btm.t880 VSS 0.18811f
C8368 C10_P_btm.t154 VSS 0.18811f
C8369 C10_P_btm.t931 VSS 0.18811f
C8370 C10_P_btm.t701 VSS 0.18811f
C8371 C10_P_btm.t109 VSS 0.18811f
C8372 C10_P_btm.t756 VSS 0.18811f
C8373 C10_P_btm.t39 VSS 0.18811f
C8374 C10_P_btm.t860 VSS 0.208624f
C8375 C10_P_btm.t1000 VSS 0.18811f
C8376 C10_P_btm.t676 VSS 0.208624f
C8377 C10_P_btm.t906 VSS 0.18811f
C8378 C10_P_btm.t560 VSS 0.18811f
C8379 C10_P_btm.t850 VSS 0.18811f
C8380 C10_P_btm.t505 VSS 0.18811f
C8381 C10_P_btm.t741 VSS 0.18811f
C8382 C10_P_btm.t1021 VSS 0.18811f
C8383 C10_P_btm.t689 VSS 0.18811f
C8384 C10_P_btm.t917 VSS 0.18811f
C8385 C10_P_btm.t134 VSS 0.18811f
C8386 C10_P_btm.t861 VSS 0.208624f
C8387 C10_P_btm.t163 VSS 0.208624f
C8388 C10_P_btm.t757 VSS 0.18811f
C8389 C10_P_btm.t213 VSS 0.18811f
C8390 C10_P_btm.t220 VSS 0.18811f
C8391 C10_P_btm.t314 VSS 0.18811f
C8392 C10_P_btm.t92 VSS 0.18811f
C8393 C10_P_btm.t873 VSS 0.18811f
C8394 C10_P_btm.t143 VSS 0.18811f
C8395 C10_P_btm.t925 VSS 0.18811f
C8396 C10_P_btm.t198 VSS 0.18811f
C8397 C10_P_btm.t1026 VSS 0.208624f
C8398 C10_P_btm.t214 VSS 0.18811f
C8399 C10_P_btm.t469 VSS 0.208624f
C8400 C10_P_btm.t460 VSS 0.18811f
C8401 C10_P_btm.t125 VSS 0.18811f
C8402 C10_P_btm.t399 VSS 0.18811f
C8403 C10_P_btm.t74 VSS 0.18811f
C8404 C10_P_btm.t293 VSS 0.18811f
C8405 C10_P_btm.t583 VSS 0.18811f
C8406 C10_P_btm.t1011 VSS 0.18811f
C8407 C10_P_btm.t478 VSS 0.18811f
C8408 C10_P_btm.t759 VSS 0.18811f
C8409 C10_P_btm.t417 VSS 0.208624f
C8410 C10_P_btm.t321 VSS 0.208624f
C8411 C10_P_btm.t670 VSS 0.18811f
C8412 C10_P_btm.t380 VSS 0.18811f
C8413 C10_P_btm.t152 VSS 0.18811f
C8414 C10_P_btm.t510 VSS 0.18811f
C8415 C10_P_btm.t204 VSS 0.18811f
C8416 C10_P_btm.t53 VSS 0.18811f
C8417 C10_P_btm.t302 VSS 0.18811f
C8418 C10_P_btm.t36 VSS 0.18811f
C8419 C10_P_btm.t363 VSS 0.18811f
C8420 C10_P_btm.t133 VSS 0.208624f
C8421 C10_P_btm.t272 VSS 0.18811f
C8422 C10_P_btm.t394 VSS 0.208624f
C8423 C10_P_btm.t638 VSS 0.18811f
C8424 C10_P_btm.t285 VSS 0.18811f
C8425 C10_P_btm.t573 VSS 0.18811f
C8426 C10_P_btm.t497 VSS 0.18811f
C8427 C10_P_btm.t468 VSS 0.18811f
C8428 C10_P_btm.t752 VSS 0.18811f
C8429 C10_P_btm.t408 VSS 0.18811f
C8430 C10_P_btm.t645 VSS 0.18811f
C8431 C10_P_btm.t928 VSS 0.18811f
C8432 C10_P_btm.t589 VSS 0.208624f
C8433 C10_P_btm.t754 VSS 0.208624f
C8434 C10_P_btm.t835 VSS 0.18811f
C8435 C10_P_btm.t544 VSS 0.18811f
C8436 C10_P_btm.t312 VSS 0.18811f
C8437 C10_P_btm.t657 VSS 0.18811f
C8438 C10_P_btm.t373 VSS 0.18811f
C8439 C10_P_btm.t142 VSS 0.18811f
C8440 C10_P_btm.t485 VSS 0.18811f
C8441 C10_P_btm.t197 VSS 0.18811f
C8442 C10_P_btm.t528 VSS 0.18811f
C8443 C10_P_btm.t295 VSS 0.208624f
C8444 C10_P_btm.t646 VSS 0.18811f
C8445 C10_P_btm.t319 VSS 0.208624f
C8446 C10_P_btm.t546 VSS 0.18811f
C8447 C10_P_btm.t215 VSS 0.18811f
C8448 C10_P_btm.t929 VSS 0.18811f
C8449 C10_P_btm.t167 VSS 0.18811f
C8450 C10_P_btm.t1045 VSS 0.18811f
C8451 C10_P_btm.t680 VSS 0.18811f
C8452 C10_P_btm.t335 VSS 0.18811f
C8453 C10_P_btm.t564 VSS 0.18811f
C8454 C10_P_btm.t853 VSS 0.18811f
C8455 C10_P_btm.t1038 VSS 0.208624f
C8456 C10_P_btm.t375 VSS 0.208624f
C8457 C10_P_btm.t56 VSS 0.18811f
C8458 C10_P_btm.t263 VSS 0.18811f
C8459 C10_P_btm.t992 VSS 0.18811f
C8460 C10_P_btm.t161 VSS 0.18811f
C8461 C10_P_btm.t445 VSS 0.18811f
C8462 C10_P_btm.t231 VSS 0.18811f
C8463 C10_P_btm.t331 VSS 0.18811f
C8464 C10_P_btm.t626 VSS 0.18811f
C8465 C10_P_btm.t277 VSS 0.208624f
C8466 C10_P_btm.t415 VSS 0.208624f
C8467 C10_P_btm.t374 VSS 0.18811f
C8468 C10_P_btm.t467 VSS 0.18811f
C8469 C10_P_btm.t518 VSS 0.18811f
C8470 C10_P_btm.t577 VSS 0.18811f
C8471 C10_P_btm.t287 VSS 0.18811f
C8472 C10_P_btm.t70 VSS 0.18811f
C8473 C10_P_btm.t397 VSS 0.18811f
C8474 C10_P_btm.t967 VSS 0.18811f
C8475 C10_P_btm.t456 VSS 0.18811f
C8476 C10_P_btm.t245 VSS 0.208624f
C8477 C10_P_btm.t313 VSS 0.18811f
C8478 C10_P_btm.t184 VSS 0.208624f
C8479 C10_P_btm.t409 VSS 0.18811f
C8480 C10_P_btm.t83 VSS 0.18811f
C8481 C10_P_btm.t357 VSS 0.18811f
C8482 C10_P_btm.t1033 VSS 0.18811f
C8483 C10_P_btm.t252 VSS 0.18811f
C8484 C10_P_btm.t532 VSS 0.18811f
C8485 C10_P_btm.t200 VSS 0.18811f
C8486 C10_P_btm.t428 VSS 0.18811f
C8487 C10_P_btm.t715 VSS 0.18811f
C8488 C10_P_btm.t51 VSS 0.208624f
C8489 C10_P_btm.t372 VSS 0.18811f
C8490 C10_P_btm.t99 VSS 0.18811f
C8491 C10_P_btm.t922 VSS 0.18811f
C8492 C10_P_btm.t195 VSS 0.18811f
C8493 C10_P_btm.t978 VSS 0.18811f
C8494 C10_P_btm.t745 VSS 0.18811f
C8495 C10_P_btm.t514 VSS 0.18811f
C8496 C10_P_btm.t806 VSS 0.18811f
C8497 C10_P_btm.t78 VSS 0.18811f
C8498 C10_P_btm.t911 VSS 0.208624f
C8499 C10_P_btm.t592 VSS 0.208624f
C8500 C10_P_btm.t288 VSS 0.18811f
C8501 C10_P_btm.t581 VSS 0.18811f
C8502 C10_P_btm.t815 VSS 0.18811f
C8503 C10_P_btm.t470 VSS 0.18811f
C8504 C10_P_btm.t704 VSS 0.18811f
C8505 C10_P_btm.t986 VSS 0.18811f
C8506 C10_P_btm.t649 VSS 0.18811f
C8507 C10_P_btm.t883 VSS 0.18811f
C8508 C10_P_btm.t595 VSS 0.18811f
C8509 C10_P_btm.t829 VSS 0.18811f
C8510 C10_P_btm.t578 VSS 0.18811f
C8511 C10_P_btm.t777 VSS 0.18811f
C8512 C10_P_btm.t1002 VSS 0.18811f
C8513 C10_P_btm.t172 VSS 0.18811f
C8514 C10_P_btm.t899 VSS 0.18811f
C8515 C10_P_btm.t512 VSS 0.18811f
C8516 C10_P_btm.t845 VSS 0.18811f
C8517 C10_P_btm.t48 VSS 0.18811f
C8518 C10_P_btm.t284 VSS 0.18811f
C8519 C10_P_btm.t1015 VSS 0.18811f
C8520 C10_P_btm.t185 VSS 0.18811f
C8521 C10_P_btm.t465 VSS 0.18811f
C8522 C10_P_btm.t129 VSS 0.208624f
C8523 C10_P_btm.t241 VSS 0.208624f
C8524 C10_P_btm.t559 VSS 0.18811f
C8525 C10_P_btm.t278 VSS 0.18811f
C8526 C10_P_btm.t474 VSS 0.18811f
C8527 C10_P_btm.t384 VSS 0.18811f
C8528 C10_P_btm.t227 VSS 0.18811f
C8529 C10_P_btm.t934 VSS 0.18811f
C8530 C10_P_btm.t209 VSS 0.18811f
C8531 C10_P_btm.t991 VSS 0.18811f
C8532 C10_P_btm.t262 VSS 0.18811f
C8533 C10_P_btm.t50 VSS 0.18811f
C8534 C10_P_btm.t429 VSS 0.18811f
C8535 C10_P_btm.t96 VSS 0.18811f
C8536 C10_P_btm.t921 VSS 0.18811f
C8537 C10_P_btm.t694 VSS 0.18811f
C8538 C10_P_btm.t977 VSS 0.18811f
C8539 C10_P_btm.t744 VSS 0.18811f
C8540 C10_P_btm.t475 VSS 0.18811f
C8541 C10_P_btm.t805 VSS 0.18811f
C8542 C10_P_btm.t568 VSS 0.18811f
C8543 C10_P_btm.t910 VSS 0.18811f
C8544 C10_P_btm.t682 VSS 0.18811f
C8545 C10_P_btm.t388 VSS 0.18811f
C8546 C10_P_btm.t692 VSS 0.18811f
C8547 C10_P_btm.t457 VSS 0.18811f
C8548 C10_P_btm.t177 VSS 0.18811f
C8549 C10_P_btm.t1036 VSS 0.18811f
C8550 C10_P_btm.t279 VSS 0.18811f
C8551 C10_P_btm.t563 VSS 0.18811f
C8552 C10_P_btm.t334 VSS 0.18811f
C8553 C10_P_btm.t239 VSS 0.18811f
C8554 C10_P_btm.t448 VSS 0.18811f
C8555 C10_P_btm.t165 VSS 0.18811f
C8556 C10_P_btm.t994 VSS 0.18811f
C8557 C10_P_btm.t267 VSS 0.18811f
C8558 C10_P_btm.t961 VSS 0.18811f
C8559 C10_P_btm.t317 VSS 0.18811f
C8560 C10_P_btm.t105 VSS 0.18811f
C8561 C10_P_btm.t875 VSS 0.18811f
C8562 C10_P_btm.t146 VSS 0.18811f
C8563 C10_P_btm.t979 VSS 0.18811f
C8564 C10_P_btm.t747 VSS 0.18811f
C8565 C10_P_btm.t1035 VSS 0.18811f
C8566 C10_P_btm.t808 VSS 0.18811f
C8567 C10_P_btm.t81 VSS 0.18811f
C8568 C10_P_btm.t856 VSS 0.18811f
C8569 C10_P_btm.t634 VSS 0.18811f
C8570 C10_P_btm.t964 VSS 0.18811f
C8571 C10_P_btm.t686 VSS 0.18811f
C8572 C10_P_btm.t454 VSS 0.18811f
C8573 C10_P_btm.t233 VSS 0.18811f
C8574 C10_P_btm.t579 VSS 0.18811f
C8575 C10_P_btm.t776 VSS 0.18811f
C8576 C10_P_btm.t218 VSS 0.18811f
C8577 C10_P_btm.t882 VSS 0.18811f
C8578 C10_P_btm.t117 VSS 0.18811f
C8579 C10_P_btm.t932 VSS 0.18811f
C8580 C10_P_btm.t702 VSS 0.18811f
C8581 C10_P_btm.t985 VSS 0.18811f
C8582 C10_P_btm.t183 VSS 0.18811f
C8583 C10_P_btm.t520 VSS 0.18811f
C8584 C10_P_btm.t865 VSS 0.18811f
C8585 C10_P_btm.t580 VSS 0.18811f
C8586 C10_P_btm.t919 VSS 0.208624f
C8587 C10_P_btm.t191 VSS 0.18811f
C8588 C10_P_btm.t145 VSS 0.208624f
C8589 C10_P_btm.t874 VSS 0.18811f
C8590 C10_P_btm.t103 VSS 0.18811f
C8591 C10_P_btm.t819 VSS 0.18811f
C8592 C10_P_btm.t974 VSS 0.18811f
C8593 C10_P_btm.t212 VSS 0.18811f
C8594 C10_P_btm.t753 VSS 0.18811f
C8595 C10_P_btm.t164 VSS 0.18811f
C8596 C10_P_btm.t386 VSS 0.18811f
C8597 C10_P_btm.t234 VSS 0.18811f
C8598 C10_P_btm.t333 VSS 0.208624f
C8599 C10_P_btm.t987 VSS 0.208624f
C8600 C10_P_btm.t758 VSS 0.18811f
C8601 C10_P_btm.t34 VSS 0.18811f
C8602 C10_P_btm.t816 VSS 0.18811f
C8603 C10_P_btm.t582 VSS 0.18811f
C8604 C10_P_btm.t866 VSS 0.18811f
C8605 C10_P_btm.t641 VSS 0.18811f
C8606 C10_P_btm.t398 VSS 0.18811f
C8607 C10_P_btm.t742 VSS 0.18811f
C8608 C10_P_btm.t458 VSS 0.18811f
C8609 C10_P_btm.t802 VSS 0.208624f
C8610 C10_P_btm.t77 VSS 0.18811f
C8611 C10_P_btm.t432 VSS 0.208624f
C8612 C10_P_btm.t110 VSS 0.18811f
C8613 C10_P_btm.t378 VSS 0.18811f
C8614 C10_P_btm.t104 VSS 0.18811f
C8615 C10_P_btm.t270 VSS 0.18811f
C8616 C10_P_btm.t993 VSS 0.18811f
C8617 C10_P_btm.t222 VSS 0.18811f
C8618 C10_P_btm.t451 VSS 0.18811f
C8619 C10_P_btm.t683 VSS 0.18811f
C8620 C10_P_btm.t387 VSS 0.18811f
C8621 C10_P_btm.t310 VSS 0.208624f
C8622 C10_P_btm.t1008 VSS 0.208624f
C8623 C10_P_btm.t788 VSS 0.18811f
C8624 C10_P_btm.t344 VSS 0.18811f
C8625 C10_P_btm.t836 VSS 0.18811f
C8626 C10_P_btm.t605 VSS 0.18811f
C8627 C10_P_btm.t889 VSS 0.18811f
C8628 C10_P_btm.t658 VSS 0.18811f
C8629 C10_P_btm.t424 VSS 0.18811f
C8630 C10_P_btm.t765 VSS 0.18811f
C8631 C10_P_btm.t487 VSS 0.18811f
C8632 C10_P_btm.t822 VSS 0.208624f
C8633 C10_P_btm.t870 VSS 0.18811f
C8634 C10_P_btm.t734 VSS 0.208624f
C8635 C10_P_btm.t1047 VSS 0.18811f
C8636 C10_P_btm.t681 VSS 0.18811f
C8637 C10_P_btm.t336 VSS 0.18811f
C8638 C10_P_btm.t565 VSS 0.18811f
C8639 C10_P_btm.t803 VSS 0.18811f
C8640 C10_P_btm.t1040 VSS 0.18811f
C8641 C10_P_btm.t743 VSS 0.18811f
C8642 C10_P_btm.t976 VSS 0.18811f
C8643 C10_P_btm.t693 VSS 0.18811f
C8644 C10_P_btm.t920 VSS 0.208624f
C8645 C10_P_btm.t868 VSS 0.208624f
C8646 C10_P_btm.t93 VSS 0.18811f
C8647 C10_P_btm.t290 VSS 0.18811f
C8648 C10_P_btm.t43 VSS 0.18811f
C8649 C10_P_btm.t907 VSS 0.18811f
C8650 C10_P_btm.t121 VSS 0.18811f
C8651 C10_P_btm.t955 VSS 0.18811f
C8652 C10_P_btm.t729 VSS 0.18811f
C8653 C10_P_btm.t420 VSS 0.18811f
C8654 C10_P_btm.t787 VSS 0.18811f
C8655 C10_P_btm.t1032 VSS 0.208624f
C8656 C10_P_btm.t237 VSS 0.18811f
C8657 C10_P_btm.t946 VSS 0.208624f
C8658 C10_P_btm.t616 VSS 0.18811f
C8659 C10_P_btm.t895 VSS 0.18811f
C8660 C10_P_btm.t551 VSS 0.18811f
C8661 C10_P_btm.t795 VSS 0.18811f
C8662 C10_P_btm.t1028 VSS 0.18811f
C8663 C10_P_btm.t735 VSS 0.18811f
C8664 C10_P_btm.t962 VSS 0.18811f
C8665 C10_P_btm.t127 VSS 0.18811f
C8666 C10_P_btm.t912 VSS 0.18811f
C8667 C10_P_btm.t79 VSS 0.208624f
C8668 C10_P_btm.t461 VSS 0.208624f
C8669 C10_P_btm.t479 VSS 0.18811f
C8670 C10_P_btm.t1044 VSS 0.18811f
C8671 C10_P_btm.t282 VSS 0.18811f
C8672 C10_P_btm.t60 VSS 0.18811f
C8673 C10_P_btm.t339 VSS 0.18811f
C8674 C10_P_btm.t473 VSS 0.18811f
C8675 C10_P_btm.t942 VSS 0.18811f
C8676 C10_P_btm.t226 VSS 0.18811f
C8677 C10_P_btm.t999 VSS 0.18811f
C8678 C10_P_btm.t273 VSS 0.208624f
C8679 C10_P_btm.t443 VSS 0.18811f
C8680 C10_P_btm.t118 VSS 0.208624f
C8681 C10_P_btm.t831 VSS 0.18811f
C8682 C10_P_btm.t228 VSS 0.18811f
C8683 C10_P_btm.t779 VSS 0.18811f
C8684 C10_P_btm.t1004 VSS 0.18811f
C8685 C10_P_btm.t173 VSS 0.18811f
C8686 C10_P_btm.t949 VSS 0.18811f
C8687 C10_P_btm.t631 VSS 0.18811f
C8688 C10_P_btm.t346 VSS 0.18811f
C8689 C10_P_btm.t65 VSS 0.18811f
C8690 C10_P_btm.t286 VSS 0.208624f
C8691 C10_P_btm.t804 VSS 0.208624f
C8692 C10_P_btm.t566 VSS 0.18811f
C8693 C10_P_btm.t854 VSS 0.18811f
C8694 C10_P_btm.t632 VSS 0.18811f
C8695 C10_P_btm.t1049 VSS 0.18811f
C8696 C10_P_btm.t684 VSS 0.18811f
C8697 C10_P_btm.t452 VSS 0.18811f
C8698 C10_P_btm.t223 VSS 0.18811f
C8699 C10_P_btm.t549 VSS 0.18811f
C8700 C10_P_btm.t271 VSS 0.18811f
C8701 C10_P_btm.t614 VSS 0.208624f
C8702 C10_P_btm.t659 VSS 0.18811f
C8703 C10_P_btm.t311 VSS 0.208624f
C8704 C10_P_btm.t49 VSS 0.18811f
C8705 C10_P_btm.t261 VSS 0.18811f
C8706 C10_P_btm.t990 VSS 0.18811f
C8707 C10_P_btm.t159 VSS 0.18811f
C8708 C10_P_btm.t1042 VSS 0.18811f
C8709 C10_P_btm.t224 VSS 0.18811f
C8710 C10_P_btm.t330 VSS 0.18811f
C8711 C10_P_btm.t562 VSS 0.18811f
C8712 C10_P_btm.t276 VSS 0.18811f
C8713 C10_P_btm.t507 VSS 0.208624f
C8714 C10_P_btm.t1014 VSS 0.208624f
C8715 C10_P_btm.t796 VSS 0.18811f
C8716 C10_P_btm.t64 VSS 0.18811f
C8717 C10_P_btm.t844 VSS 0.18811f
C8718 C10_P_btm.t617 VSS 0.18811f
C8719 C10_P_btm.t896 VSS 0.18811f
C8720 C10_P_btm.t668 VSS 0.18811f
C8721 C10_P_btm.t435 VSS 0.18811f
C8722 C10_P_btm.t775 VSS 0.18811f
C8723 C10_P_btm.t500 VSS 0.18811f
C8724 C10_P_btm.t828 VSS 0.208624f
C8725 C10_P_btm.t878 VSS 0.18811f
C8726 C10_P_btm.t656 VSS 0.208624f
C8727 C10_P_btm.t151 VSS 0.18811f
C8728 C10_P_btm.t603 VSS 0.18811f
C8729 C10_P_btm.t260 VSS 0.18811f
C8730 C10_P_btm.t699 VSS 0.18811f
C8731 C10_P_btm.t728 VSS 0.18811f
C8732 C10_P_btm.t444 VSS 0.18811f
C8733 C10_P_btm.t675 VSS 0.18811f
C8734 C10_P_btm.t905 VSS 0.18811f
C8735 C10_P_btm.t625 VSS 0.18811f
C8736 C10_P_btm.t849 VSS 0.208624f
C8737 C10_P_btm.t139 VSS 0.208624f
C8738 C10_P_btm.t303 VSS 0.18811f
C8739 C10_P_btm.t94 VSS 0.18811f
C8740 C10_P_btm.t205 VSS 0.18811f
C8741 C10_P_btm.t438 VSS 0.18811f
C8742 C10_P_btm.t153 VSS 0.18811f
C8743 C10_P_btm.t381 VSS 0.18811f
C8744 C10_P_btm.t619 VSS 0.18811f
C8745 C10_P_btm.t322 VSS 0.18811f
C8746 C10_P_btm.t552 VSS 0.208624f
C8747 C10_P_btm.t174 VSS 0.208624f
C8748 C10_P_btm.t1005 VSS 0.18811f
C8749 C10_P_btm.t240 VSS 0.18811f
C8750 C10_P_btm.t1010 VSS 0.18811f
C8751 C10_P_btm.t832 VSS 0.18811f
C8752 C10_P_btm.t243 VSS 0.18811f
C8753 C10_P_btm.t884 VSS 0.18811f
C8754 C10_P_btm.t652 VSS 0.18811f
C8755 C10_P_btm.t988 VSS 0.18811f
C8756 C10_P_btm.t706 VSS 0.18811f
C8757 C10_P_btm.t37 VSS 0.208624f
C8758 C10_P_btm.t40 VSS 0.18811f
C8759 C10_P_btm.t877 VSS 0.208624f
C8760 C10_P_btm.t530 VSS 0.18811f
C8761 C10_P_btm.t824 VSS 0.18811f
C8762 C10_P_btm.t492 VSS 0.18811f
C8763 C10_P_btm.t714 VSS 0.18811f
C8764 C10_P_btm.t939 VSS 0.18811f
C8765 C10_P_btm.t661 VSS 0.18811f
C8766 C10_P_btm.t891 VSS 0.18811f
C8767 C10_P_btm.t57 VSS 0.18811f
C8768 C10_P_btm.t839 VSS 0.18811f
C8769 C10_P_btm.t385 VSS 0.208624f
C8770 C10_P_btm.t160 VSS 0.18811f
C8771 C10_P_btm.t446 VSS 0.18811f
C8772 C10_P_btm.t211 VSS 0.18811f
C8773 C10_P_btm.t52 VSS 0.18811f
C8774 C10_P_btm.t264 VSS 0.18811f
C8775 C10_P_btm.t55 VSS 0.18811f
C8776 C10_P_btm.t871 VSS 0.18811f
C8777 C10_P_btm.t141 VSS 0.18811f
C8778 C10_P_btm.t924 VSS 0.18811f
C8779 C10_P_btm.t196 VSS 0.208624f
C8780 C10_P_btm.t30 VSS 0.216875f
C8781 C10_P_btm.t703 VSS 0.208624f
C8782 C10_P_btm.t362 VSS 0.18811f
C8783 C10_P_btm.t648 VSS 0.18811f
C8784 C10_P_btm.t301 VSS 0.18811f
C8785 C10_P_btm.t536 VSS 0.18811f
C8786 C10_P_btm.t778 VSS 0.18811f
C8787 C10_P_btm.t509 VSS 0.18811f
C8788 C10_P_btm.t719 VSS 0.18811f
C8789 C10_P_btm.t948 VSS 0.18811f
C8790 C10_P_btm.t669 VSS 0.18811f
C8791 C10_P_btm.t897 VSS 0.208624f
C8792 C10_P_btm.t17 VSS 0.208975f
C8793 C10_P_btm.n3897 VSS 0.100784f
C8794 VDD.n5 VSS 0.399626f
C8795 VDD.t3216 VSS 0.197243f
C8796 VDD.t3120 VSS 0.197241f
C8797 VDD.t3185 VSS 0.198209f
C8798 VDD.n9 VSS 0.204946f
C8799 VDD.t1318 VSS 0.105641f
C8800 VDD.t2720 VSS 0.174244f
C8801 VDD.n27 VSS 0.219516f
C8802 VDD.n28 VSS 0.508669f
C8803 VDD.n29 VSS 0.197477f
C8804 VDD.n30 VSS 0.181171f
C8805 VDD.n31 VSS 0.172458f
C8806 VDD.n32 VSS 0.172458f
C8807 VDD.n33 VSS 0.203068f
C8808 VDD.n34 VSS 0.226793f
C8809 VDD.n35 VSS 0.528149f
C8810 VDD.t157 VSS 0.595346f
C8811 VDD.t3087 VSS 0.644138f
C8812 VDD.t3058 VSS 0.644138f
C8813 VDD.t2040 VSS 0.644138f
C8814 VDD.t3078 VSS 0.644138f
C8815 VDD.t144 VSS 0.64813f
C8816 VDD.t3039 VSS 0.496412f
C8817 VDD.t2039 VSS 0.340701f
C8818 VDD.t2038 VSS 0.340701f
C8819 VDD.t88 VSS 0.340701f
C8820 VDD.t86 VSS 0.340701f
C8821 VDD.t89 VSS 0.340701f
C8822 VDD.t87 VSS 0.340701f
C8823 VDD.t579 VSS 0.340701f
C8824 VDD.t578 VSS 0.340701f
C8825 VDD.t583 VSS 0.20096f
C8826 VDD.n37 VSS 0.139741f
C8827 VDD.t584 VSS 0.270165f
C8828 VDD.t581 VSS 0.340701f
C8829 VDD.t582 VSS 0.340701f
C8830 VDD.t577 VSS 0.340701f
C8831 VDD.t580 VSS 0.340701f
C8832 VDD.t3003 VSS 0.340701f
C8833 VDD.t3005 VSS 0.340701f
C8834 VDD.t2991 VSS 0.340701f
C8835 VDD.t2998 VSS 0.340701f
C8836 VDD.t3000 VSS 0.340701f
C8837 VDD.t3004 VSS 0.340701f
C8838 VDD.t2992 VSS 0.340701f
C8839 VDD.t2997 VSS 0.340701f
C8840 VDD.t2990 VSS 0.340701f
C8841 VDD.t2993 VSS 0.340701f
C8842 VDD.t2999 VSS 0.340701f
C8843 VDD.t3001 VSS 0.340701f
C8844 VDD.t2995 VSS 0.340701f
C8845 VDD.t2996 VSS 0.340701f
C8846 VDD.t2994 VSS 0.340701f
C8847 VDD.t3002 VSS 0.437214f
C8848 VDD.n38 VSS 0.521253f
C8849 VDD.n39 VSS 0.197665f
C8850 VDD.n40 VSS 0.19461f
C8851 VDD.n41 VSS 0.176023f
C8852 VDD.n42 VSS 0.489f
C8853 VDD.n43 VSS 0.372762f
C8854 VDD.n44 VSS 1.05127f
C8855 VDD.n45 VSS 1.4343f
C8856 VDD.t2762 VSS 0.174244f
C8857 VDD.t824 VSS 0.105641f
C8858 VDD.n63 VSS 0.48901f
C8859 VDD.n64 VSS 0.508669f
C8860 VDD.n65 VSS 0.176023f
C8861 VDD.n66 VSS 0.181171f
C8862 VDD.n67 VSS 0.172458f
C8863 VDD.n68 VSS 0.172458f
C8864 VDD.n69 VSS 0.197484f
C8865 VDD.n70 VSS 0.203082f
C8866 VDD.n71 VSS 0.226772f
C8867 VDD.n72 VSS 0.528149f
C8868 VDD.t143 VSS 0.595346f
C8869 VDD.t2975 VSS 0.644138f
C8870 VDD.t3070 VSS 0.644138f
C8871 VDD.t412 VSS 0.644138f
C8872 VDD.t172 VSS 0.644138f
C8873 VDD.t2976 VSS 0.64813f
C8874 VDD.t602 VSS 0.496412f
C8875 VDD.t254 VSS 0.340701f
C8876 VDD.t255 VSS 0.340701f
C8877 VDD.t2933 VSS 0.340701f
C8878 VDD.t2932 VSS 0.340701f
C8879 VDD.t2930 VSS 0.340701f
C8880 VDD.t2931 VSS 0.340701f
C8881 VDD.t2053 VSS 0.340701f
C8882 VDD.t2057 VSS 0.340701f
C8883 VDD.t2055 VSS 0.20096f
C8884 VDD.n74 VSS 0.139741f
C8885 VDD.t2056 VSS 0.270165f
C8886 VDD.t2051 VSS 0.340701f
C8887 VDD.t2058 VSS 0.340701f
C8888 VDD.t2054 VSS 0.340701f
C8889 VDD.t2052 VSS 0.340701f
C8890 VDD.t521 VSS 0.340701f
C8891 VDD.t529 VSS 0.340701f
C8892 VDD.t522 VSS 0.340701f
C8893 VDD.t528 VSS 0.340701f
C8894 VDD.t518 VSS 0.340701f
C8895 VDD.t520 VSS 0.340701f
C8896 VDD.t516 VSS 0.340701f
C8897 VDD.t524 VSS 0.340701f
C8898 VDD.t530 VSS 0.340701f
C8899 VDD.t526 VSS 0.340701f
C8900 VDD.t531 VSS 0.340701f
C8901 VDD.t527 VSS 0.340701f
C8902 VDD.t523 VSS 0.340701f
C8903 VDD.t519 VSS 0.340701f
C8904 VDD.t525 VSS 0.340701f
C8905 VDD.t517 VSS 0.437214f
C8906 VDD.n75 VSS 0.521253f
C8907 VDD.n76 VSS 0.197665f
C8908 VDD.n77 VSS 0.19461f
C8909 VDD.n78 VSS 0.219513f
C8910 VDD.n79 VSS 0.372803f
C8911 VDD.n80 VSS 1.0866f
C8912 VDD.t3189 VSS 0.198208f
C8913 VDD.n81 VSS 0.390552f
C8914 VDD.n82 VSS 0.399389f
C8915 VDD.t3188 VSS 0.197241f
C8916 VDD.t3174 VSS 0.197243f
C8917 VDD.n86 VSS 2.41015f
C8918 VDD.n87 VSS 0.359186f
C8919 VDD.n88 VSS 0.142013f
C8920 VDD.n89 VSS 0.933884f
C8921 VDD.n104 VSS 0.933884f
C8922 VDD.n105 VSS 0.141077f
C8923 VDD.n106 VSS 0.344308f
C8924 VDD.n107 VSS 0.103881f
C8925 VDD.n108 VSS 0.127011f
C8926 VDD.t146 VSS 10.3255f
C8927 VDD.t148 VSS 10.3255f
C8928 VDD.n109 VSS 0.147198f
C8929 VDD.n110 VSS 0.104018f
C8930 VDD.t2794 VSS 0.103345f
C8931 VDD.t1802 VSS 0.136262f
C8932 VDD.t64 VSS 0.119803f
C8933 VDD.t726 VSS 0.143917f
C8934 VDD.t642 VSS 0.163656f
C8935 VDD.n123 VSS 0.169999f
C8936 VDD.t2792 VSS 0.130036f
C8937 VDD.n132 VSS 0.350339f
C8938 VDD.n133 VSS 3.85796f
C8939 VDD.n134 VSS 0.156352f
C8940 VDD.n135 VSS 0.127218f
C8941 VDD.n136 VSS 4.02892f
C8942 VDD.n137 VSS 0.127011f
C8943 VDD.n138 VSS 0.134395f
C8944 VDD.n139 VSS 0.338605f
C8945 VDD.n141 VSS 0.145543f
C8946 VDD.n142 VSS 0.152384f
C8947 VDD.n144 VSS 0.377186f
C8948 VDD.n145 VSS 0.296901f
C8949 VDD.n146 VSS 0.200448f
C8950 VDD.t151 VSS 13.2771f
C8951 VDD.n147 VSS 0.200448f
C8952 VDD.n148 VSS 0.198303f
C8953 VDD.n149 VSS 0.682538f
C8954 VDD.n150 VSS 0.374374f
C8955 VDD.t2940 VSS 0.143871f
C8956 VDD.n151 VSS 0.502169f
C8957 VDD.n152 VSS 0.933884f
C8958 VDD.t2938 VSS 0.183093f
C8959 VDD.n155 VSS 0.545063f
C8960 VDD.n169 VSS 0.214529f
C8961 VDD.n171 VSS 0.500329f
C8962 VDD.t147 VSS 0.183093f
C8963 VDD.n174 VSS 0.933884f
C8964 VDD.t150 VSS 0.143871f
C8965 VDD.n175 VSS 0.502169f
C8966 VDD.n176 VSS 0.275367f
C8967 VDD.n177 VSS 0.432717f
C8968 VDD.n178 VSS 5.83461f
C8969 VDD.t452 VSS 0.122079f
C8970 VDD.t451 VSS 0.124007f
C8971 VDD.n179 VSS 0.316573f
C8972 VDD.t454 VSS 0.122361f
C8973 VDD.t455 VSS 0.124313f
C8974 VDD.n180 VSS 0.309585f
C8975 VDD.n181 VSS 0.365643f
C8976 VDD.n182 VSS 0.483305f
C8977 VDD.n183 VSS 0.118962f
C8978 VDD.n189 VSS 0.345f
C8979 VDD.n193 VSS 0.163438f
C8980 VDD.n198 VSS 0.103813f
C8981 VDD.t2919 VSS 0.134816f
C8982 VDD.n205 VSS 0.105075f
C8983 VDD.n206 VSS 0.11908f
C8984 VDD.n207 VSS 0.15281f
C8985 VDD.n215 VSS 0.346552f
C8986 VDD.t2241 VSS 0.783951f
C8987 VDD.t2243 VSS 0.407444f
C8988 VDD.t2254 VSS 0.407444f
C8989 VDD.t2255 VSS 0.35436f
C8990 VDD.t2249 VSS 0.35436f
C8991 VDD.t2246 VSS 0.407444f
C8992 VDD.t2252 VSS 0.407444f
C8993 VDD.t2247 VSS 0.720035f
C8994 VDD.t2244 VSS 0.720034f
C8995 VDD.t2240 VSS 0.407444f
C8996 VDD.t2250 VSS 0.407444f
C8997 VDD.t2251 VSS 0.35436f
C8998 VDD.t2242 VSS 0.35436f
C8999 VDD.t2245 VSS 0.407444f
C9000 VDD.t2248 VSS 0.407444f
C9001 VDD.t2253 VSS 0.806546f
C9002 VDD.t2917 VSS 0.159305f
C9003 VDD.t448 VSS 0.746798f
C9004 VDD.n222 VSS 0.107107f
C9005 VDD.t2941 VSS 0.125461f
C9006 VDD.n227 VSS 0.11869f
C9007 VDD.t145 VSS 0.125461f
C9008 VDD.n229 VSS 0.11869f
C9009 VDD.n235 VSS 0.295819f
C9010 VDD.n236 VSS 0.127858f
C9011 VDD.t447 VSS 0.115153f
C9012 VDD.n248 VSS 0.110367f
C9013 VDD.n253 VSS 0.165741f
C9014 VDD.n256 VSS 0.165741f
C9015 VDD.t2494 VSS 0.163193f
C9016 VDD.t2286 VSS 0.146208f
C9017 VDD.n258 VSS 0.18361f
C9018 VDD.t2580 VSS 0.146208f
C9019 VDD.t2646 VSS 0.163193f
C9020 VDD.n270 VSS 0.357352f
C9021 VDD.n272 VSS 0.626421f
C9022 VDD.n273 VSS 0.280223f
C9023 VDD.t457 VSS 0.115153f
C9024 VDD.n277 VSS 0.10889f
C9025 VDD.t437 VSS 0.115153f
C9026 VDD.n280 VSS 0.10889f
C9027 VDD.t459 VSS 0.115153f
C9028 VDD.n284 VSS 0.10889f
C9029 VDD.t445 VSS 0.115153f
C9030 VDD.n289 VSS 0.10889f
C9031 VDD.t435 VSS 0.115153f
C9032 VDD.n292 VSS 0.10889f
C9033 VDD.t449 VSS 0.115153f
C9034 VDD.n296 VSS 0.10889f
C9035 VDD.t461 VSS 0.115153f
C9036 VDD.n301 VSS 0.10889f
C9037 VDD.t439 VSS 0.115153f
C9038 VDD.n304 VSS 0.10889f
C9039 VDD.t443 VSS 0.115153f
C9040 VDD.n308 VSS 0.10889f
C9041 VDD.t441 VSS 0.115153f
C9042 VDD.n313 VSS 0.10889f
C9043 VDD.n318 VSS 0.298427f
C9044 VDD.t460 VSS 0.746798f
C9045 VDD.t438 VSS 0.746798f
C9046 VDD.t442 VSS 0.746798f
C9047 VDD.t440 VSS 0.746798f
C9048 VDD.t453 VSS 0.768707f
C9049 VDD.n319 VSS 0.397119f
C9050 VDD.n320 VSS 0.105573f
C9051 VDD.t434 VSS 0.746798f
C9052 VDD.t444 VSS 0.746798f
C9053 VDD.t458 VSS 0.746798f
C9054 VDD.t436 VSS 0.641093f
C9055 VDD.n321 VSS 0.384841f
C9056 VDD.t456 VSS 0.479104f
C9057 VDD.t446 VSS 0.746798f
C9058 VDD.t450 VSS 0.699972f
C9059 VDD.n322 VSS 0.108437f
C9060 VDD.n323 VSS 0.289069f
C9061 VDD.n325 VSS 0.160304f
C9062 VDD.n326 VSS 0.214626f
C9063 VDD.n327 VSS 0.449714f
C9064 VDD.n328 VSS 0.226567f
C9065 VDD.n329 VSS 0.634214f
C9066 VDD.n330 VSS 3.66081f
C9067 VDD.n339 VSS 0.248022f
C9068 VDD.t58 VSS 0.431687f
C9069 VDD.n347 VSS 0.132334f
C9070 VDD.t61 VSS 0.44032f
C9071 VDD.t3035 VSS 0.338494f
C9072 VDD.t2927 VSS 0.113833f
C9073 VDD.t2768 VSS 0.113022f
C9074 VDD.n389 VSS 0.132548f
C9075 VDD.t464 VSS 0.338494f
C9076 VDD.n393 VSS 0.211863f
C9077 VDD.n396 VSS 0.155125f
C9078 VDD.n397 VSS 0.124392f
C9079 VDD.n398 VSS 0.10056f
C9080 VDD.n402 VSS 0.147431f
C9081 VDD.n405 VSS 0.12216f
C9082 VDD.n430 VSS 0.232929f
C9083 VDD.n431 VSS 0.188399f
C9084 VDD.n437 VSS 2.51755f
C9085 VDD.n438 VSS 2.61527f
C9086 VDD.t2348 VSS 0.142769f
C9087 VDD.t94 VSS 0.120952f
C9088 VDD.t335 VSS 0.10411f
C9089 VDD.t358 VSS 0.10411f
C9090 VDD.n628 VSS 0.11419f
C9091 VDD.t1783 VSS 0.104876f
C9092 VDD.t1541 VSS 0.108321f
C9093 VDD.t2473 VSS 0.142003f
C9094 VDD.t2382 VSS 0.212048f
C9095 VDD.t1971 VSS 0.141621f
C9096 VDD.n645 VSS 0.137209f
C9097 VDD.t3019 VSS 0.110234f
C9098 VDD.t1442 VSS 0.105641f
C9099 VDD.t2607 VSS 0.141621f
C9100 VDD.t2529 VSS 0.141621f
C9101 VDD.t1150 VSS 0.175303f
C9102 VDD.t2369 VSS 0.14851f
C9103 VDD.t901 VSS 0.113679f
C9104 VDD.t651 VSS 0.124014f
C9105 VDD.t227 VSS 0.121717f
C9106 VDD.t1107 VSS 0.102579f
C9107 VDD.n701 VSS 0.137209f
C9108 VDD.t3067 VSS 0.102197f
C9109 VDD.t1485 VSS 0.113297f
C9110 VDD.t2271 VSS 0.140855f
C9111 VDD.t1305 VSS 0.129372f
C9112 VDD.t2258 VSS 0.223914f
C9113 VDD.n817 VSS 0.100894f
C9114 VDD.n874 VSS 0.121516f
C9115 VDD.t681 VSS 0.108321f
C9116 VDD.t972 VSS 0.108321f
C9117 VDD.t603 VSS 0.122483f
C9118 VDD.t2634 VSS 0.106407f
C9119 VDD.t2222 VSS 0.103728f
C9120 VDD.t1366 VSS 0.10411f
C9121 VDD.t2563 VSS 0.102197f
C9122 VDD.t710 VSS 0.135114f
C9123 VDD.n875 VSS 0.172423f
C9124 VDD.t1985 VSS 0.122483f
C9125 VDD.t2261 VSS 0.106407f
C9126 VDD.t2414 VSS 0.145831f
C9127 VDD.t1918 VSS 0.117998f
C9128 VDD.n1230 VSS 0.123812f
C9129 VDD.t344 VSS 0.105641f
C9130 VDD.t2517 VSS 0.223914f
C9131 VDD.t66 VSS 0.105641f
C9132 VDD.t2470 VSS 0.106407f
C9133 VDD.t2509 VSS 0.141621f
C9134 VDD.n1257 VSS 0.844243f
C9135 VDD.t3225 VSS 0.147331f
C9136 VDD.t1163 VSS 0.10679f
C9137 VDD.t2663 VSS 0.110617f
C9138 VDD.t12 VSS 0.10411f
C9139 VDD.t1307 VSS 0.109469f
C9140 VDD.t592 VSS 0.102197f
C9141 VDD.t2296 VSS 0.223914f
C9142 VDD.t1062 VSS 0.121334f
C9143 VDD.t873 VSS 0.108703f
C9144 VDD.t3236 VSS 0.147331f
C9145 VDD.t3182 VSS 0.147331f
C9146 VDD.n1624 VSS 0.106306f
C9147 VDD.t2650 VSS 0.209752f
C9148 VDD.t2556 VSS 0.212814f
C9149 VDD.t2506 VSS 0.285921f
C9150 VDD.t137 VSS 0.283624f
C9151 VDD.t1364 VSS 0.104876f
C9152 VDD.t1216 VSS 0.102197f
C9153 VDD.t1823 VSS 0.102579f
C9154 VDD.t2523 VSS 0.140855f
C9155 VDD.n1676 VSS 0.130629f
C9156 VDD.n1923 VSS 0.100894f
C9157 VDD.t2417 VSS 0.223914f
C9158 VDD.t879 VSS 0.121334f
C9159 VDD.t2122 VSS 0.108703f
C9160 VDD.t735 VSS 0.104493f
C9161 VDD.t1140 VSS 0.109086f
C9162 VDD.t3029 VSS 0.104876f
C9163 VDD.t3027 VSS 0.105641f
C9164 VDD.t260 VSS 0.105641f
C9165 VDD.t262 VSS 0.105641f
C9166 VDD.t129 VSS 0.105641f
C9167 VDD.t2428 VSS 0.1776f
C9168 VDD.t2572 VSS 0.299317f
C9169 VDD.n2059 VSS 0.200144f
C9170 VDD.n2087 VSS 0.470888f
C9171 VDD.n2113 VSS 0.137486f
C9172 VDD.t3149 VSS 0.147331f
C9173 VDD.n2226 VSS 0.11419f
C9174 VDD.t3195 VSS 0.147331f
C9175 VDD.t99 VSS 0.107172f
C9176 VDD.t423 VSS 0.103345f
C9177 VDD.t2601 VSS 0.229655f
C9178 VDD.t2643 VSS 0.211283f
C9179 VDD.t350 VSS 0.103345f
C9180 VDD.t2114 VSS 0.134348f
C9181 VDD.t1192 VSS 0.13741f
C9182 VDD.t1274 VSS 0.106407f
C9183 VDD.t1786 VSS 0.104876f
C9184 VDD.t2016 VSS 0.107938f
C9185 VDD.t2694 VSS 0.106407f
C9186 VDD.t3023 VSS 0.112531f
C9187 VDD.n2287 VSS 0.111874f
C9188 VDD.t3235 VSS 0.147331f
C9189 VDD.t957 VSS 0.109852f
C9190 VDD.t1118 VSS 0.113679f
C9191 VDD.t557 VSS 0.121334f
C9192 VDD.t692 VSS 0.127459f
C9193 VDD.t2673 VSS 0.128224f
C9194 VDD.t2613 VSS 0.158462f
C9195 VDD.t3219 VSS 0.147331f
C9196 VDD.t44 VSS 0.112914f
C9197 VDD.t2476 VSS 0.176834f
C9198 VDD.t2388 VSS 0.282476f
C9199 VDD.t2877 VSS 0.193676f
C9200 VDD.n2369 VSS 0.127013f
C9201 VDD.t1196 VSS 0.107172f
C9202 VDD.t2409 VSS 0.109852f
C9203 VDD.t2590 VSS 0.193676f
C9204 VDD.n2376 VSS 0.148218f
C9205 VDD.t3139 VSS 0.147331f
C9206 VDD.t2290 VSS 0.223914f
C9207 VDD.t1284 VSS 0.121334f
C9208 VDD.t538 VSS 0.108703f
C9209 VDD.t3209 VSS 0.147331f
C9210 VDD.t3138 VSS 0.147331f
C9211 VDD.t3133 VSS 0.150109f
C9212 VDD.t3063 VSS 0.209752f
C9213 VDD.t2550 VSS 0.248027f
C9214 VDD.t2363 VSS 0.352138f
C9215 VDD.t2566 VSS 0.422565f
C9216 VDD.t2268 VSS 0.22889f
C9217 VDD.t1047 VSS 0.108321f
C9218 VDD.t1811 VSS 0.107555f
C9219 VDD.t1977 VSS 0.107555f
C9220 VDD.t1975 VSS 0.10411f
C9221 VDD.t2704 VSS 0.10411f
C9222 VDD.t981 VSS 0.200948f
C9223 VDD.n2494 VSS 0.253494f
C9224 VDD.t1935 VSS 0.130521f
C9225 VDD.t1926 VSS 0.130138f
C9226 VDD.t2596 VSS 0.102579f
C9227 VDD.t267 VSS 0.134731f
C9228 VDD.t2366 VSS 0.223914f
C9229 VDD.t1303 VSS 0.121334f
C9230 VDD.t306 VSS 0.108703f
C9231 VDD.t671 VSS 0.104493f
C9232 VDD.t1422 VSS 0.109086f
C9233 VDD.t2873 VSS 0.104876f
C9234 VDD.t2870 VSS 0.105641f
C9235 VDD.t280 VSS 0.105641f
C9236 VDD.t278 VSS 0.105641f
C9237 VDD.t70 VSS 0.105641f
C9238 VDD.t72 VSS 0.10411f
C9239 VDD.t2422 VSS 0.1776f
C9240 VDD.t2357 VSS 0.193676f
C9241 VDD.t2336 VSS 0.158462f
C9242 VDD.n2867 VSS 0.179604f
C9243 VDD.n2892 VSS 0.470888f
C9244 VDD.t2320 VSS 0.223914f
C9245 VDD.t1857 VSS 0.121334f
C9246 VDD.t125 VSS 0.108703f
C9247 VDD.t3220 VSS 0.147331f
C9248 VDD.t3143 VSS 0.147331f
C9249 VDD.t3238 VSS 0.147331f
C9250 VDD.t3199 VSS 0.147331f
C9251 VDD.t264 VSS 0.24841f
C9252 VDD.t2628 VSS 0.247262f
C9253 VDD.t2526 VSS 0.422565f
C9254 VDD.t2274 VSS 0.422565f
C9255 VDD.t2622 VSS 0.22889f
C9256 VDD.t2030 VSS 0.109086f
C9257 VDD.t406 VSS 0.131669f
C9258 VDD.t402 VSS 0.111383f
C9259 VDD.t731 VSS 0.123248f
C9260 VDD.t548 VSS 0.104876f
C9261 VDD.n3134 VSS 0.257175f
C9262 VDD.n3295 VSS 0.112239f
C9263 VDD.t411 VSS 0.105641f
C9264 VDD.t3025 VSS 0.10411f
C9265 VDD.t2967 VSS 0.108703f
C9266 VDD.t22 VSS 0.100665f
C9267 VDD.t2675 VSS 0.10679f
C9268 VDD.t2520 VSS 0.159993f
C9269 VDD.t1330 VSS 0.106407f
C9270 VDD.t1134 VSS 0.100665f
C9271 VDD.t364 VSS 0.10411f
C9272 VDD.t1601 VSS 0.114445f
C9273 VDD.n3423 VSS 0.107263f
C9274 VDD.t356 VSS 0.102197f
C9275 VDD.t2299 VSS 0.223914f
C9276 VDD.t1595 VSS 0.121334f
C9277 VDD.t368 VSS 0.108703f
C9278 VDD.t1453 VSS 0.104493f
C9279 VDD.t113 VSS 0.283624f
C9280 VDD.t2283 VSS 0.528972f
C9281 VDD.t2333 VSS 0.388117f
C9282 VDD.t366 VSS 0.123248f
C9283 VDD.t3128 VSS 0.147331f
C9284 VDD.t3217 VSS 0.147331f
C9285 VDD.n3585 VSS 0.13552f
C9286 VDD.n3658 VSS 0.470888f
C9287 VDD.t3126 VSS 0.147331f
C9288 VDD.t3212 VSS 0.148035f
C9289 VDD.t3221 VSS 0.147331f
C9290 VDD.t3114 VSS 0.147331f
C9291 VDD.n3791 VSS 0.11419f
C9292 VDD.t3150 VSS 0.147798f
C9293 VDD.t2287 VSS 0.223914f
C9294 VDD.t1136 VSS 0.121334f
C9295 VDD.t314 VSS 0.108321f
C9296 VDD.t162 VSS 0.149276f
C9297 VDD.t1148 VSS 0.157314f
C9298 VDD.t84 VSS 0.140855f
C9299 VDD.t2479 VSS 0.247645f
C9300 VDD.t2323 VSS 0.141621f
C9301 VDD.n3837 VSS 0.124195f
C9302 VDD.t298 VSS 0.102579f
C9303 VDD.t1372 VSS 0.100665f
C9304 VDD.t26 VSS 0.107555f
C9305 VDD.t2748 VSS 0.108321f
C9306 VDD.n3838 VSS 0.113258f
C9307 VDD.t2302 VSS 0.141621f
C9308 VDD.t2811 VSS 0.141621f
C9309 VDD.t717 VSS 0.177217f
C9310 VDD.t2455 VSS 0.180279f
C9311 VDD.t2277 VSS 0.247262f
C9312 VDD.t587 VSS 0.2442f
C9313 VDD.n3839 VSS 0.133381f
C9314 VDD.t117 VSS 0.110234f
C9315 VDD.t1340 VSS 0.107172f
C9316 VDD.t2425 VSS 0.188317f
C9317 VDD.t2503 VSS 0.193676f
C9318 VDD.n3840 VSS 0.182423f
C9319 VDD.t2400 VSS 0.264869f
C9320 VDD.t683 VSS 0.173772f
C9321 VDD.t1895 VSS 0.104493f
C9322 VDD.t1896 VSS 0.143917f
C9323 VDD.t1809 VSS 0.210517f
C9324 VDD.t2360 VSS 0.253386f
C9325 VDD.t2500 VSS 0.193676f
C9326 VDD.n3841 VSS 0.19003f
C9327 VDD.t155 VSS 0.143152f
C9328 VDD.t2461 VSS 0.247645f
C9329 VDD.t2443 VSS 0.352138f
C9330 VDD.t2487 VSS 0.247262f
C9331 VDD.t2828 VSS 0.140855f
C9332 VDD.t1019 VSS 0.124014f
C9333 VDD.t276 VSS 0.108321f
C9334 VDD.n3877 VSS 0.127013f
C9335 VDD.t3121 VSS 0.150126f
C9336 VDD.t3119 VSS 0.147331f
C9337 VDD.n3918 VSS 0.127013f
C9338 VDD.n4030 VSS 0.106306f
C9339 VDD.n4181 VSS 0.127013f
C9340 VDD.t923 VSS 0.114062f
C9341 VDD.t195 VSS 0.106407f
C9342 VDD.t2110 VSS 0.173772f
C9343 VDD.t2631 VSS 0.145831f
C9344 VDD.t2020 VSS 0.174538f
C9345 VDD.t2593 VSS 0.149276f
C9346 VDD.t323 VSS 0.12631f
C9347 VDD.t1603 VSS 0.110617f
C9348 VDD.t2001 VSS 0.142769f
C9349 VDD.t2434 VSS 0.250707f
C9350 VDD.t2514 VSS 0.28171f
C9351 VDD.t2351 VSS 0.248027f
C9352 VDD.t1517 VSS 0.139324f
C9353 VDD.t2581 VSS 0.123248f
C9354 VDD.n4251 VSS 0.137592f
C9355 VDD.t3159 VSS 0.147331f
C9356 VDD.t321 VSS 0.104493f
C9357 VDD.t562 VSS 0.102579f
C9358 VDD.t1232 VSS 0.130521f
C9359 VDD.t675 VSS 0.106407f
C9360 VDD.t975 VSS 0.118655f
C9361 VDD.t893 VSS 0.118655f
C9362 VDD.t2342 VSS 0.223914f
C9363 VDD.t270 VSS 0.108321f
C9364 VDD.t20 VSS 0.105641f
C9365 VDD.t617 VSS 0.104876f
C9366 VDD.t2440 VSS 0.145831f
C9367 VDD.t1947 VSS 0.107555f
C9368 VDD.n4364 VSS 0.121516f
C9369 VDD.t3191 VSS 0.147331f
C9370 VDD.n4467 VSS 0.49361f
C9371 a_8912_37509.t25 VSS 0.784296f
C9372 a_8912_37509.t30 VSS 0.177274f
C9373 a_8912_37509.t35 VSS 0.177274f
C9374 a_8912_37509.n0 VSS 0.494639f
C9375 a_8912_37509.n1 VSS 2.08091f
C9376 a_8912_37509.t22 VSS 0.177274f
C9377 a_8912_37509.t36 VSS 0.177274f
C9378 a_8912_37509.n2 VSS 0.494639f
C9379 a_8912_37509.n3 VSS 1.04163f
C9380 a_8912_37509.t28 VSS 0.177274f
C9381 a_8912_37509.t26 VSS 0.177274f
C9382 a_8912_37509.n4 VSS 0.494639f
C9383 a_8912_37509.n5 VSS 1.04724f
C9384 a_8912_37509.t34 VSS 0.779123f
C9385 a_8912_37509.n6 VSS 1.13411f
C9386 a_8912_37509.t7 VSS 0.779123f
C9387 a_8912_37509.n7 VSS 1.12851f
C9388 a_8912_37509.t19 VSS 0.177274f
C9389 a_8912_37509.t15 VSS 0.177274f
C9390 a_8912_37509.n8 VSS 0.494639f
C9391 a_8912_37509.n9 VSS 1.04163f
C9392 a_8912_37509.t18 VSS 0.177274f
C9393 a_8912_37509.t10 VSS 0.177274f
C9394 a_8912_37509.n10 VSS 0.494639f
C9395 a_8912_37509.n11 VSS 1.04163f
C9396 a_8912_37509.t17 VSS 0.177274f
C9397 a_8912_37509.t9 VSS 0.177274f
C9398 a_8912_37509.n12 VSS 0.494639f
C9399 a_8912_37509.n13 VSS 1.04163f
C9400 a_8912_37509.t11 VSS 0.779123f
C9401 a_8912_37509.n14 VSS 1.59247f
C9402 a_8912_37509.n15 VSS 0.760578f
C9403 a_8912_37509.n16 VSS 0.459486f
C9404 a_8912_37509.t4 VSS 0.890777f
C9405 a_8912_37509.n17 VSS 0.548555f
C9406 a_8912_37509.t3 VSS 0.890777f
C9407 a_8912_37509.t1 VSS 0.890777f
C9408 a_8912_37509.n18 VSS 1.34409f
C9409 a_8912_37509.t5 VSS 0.890777f
C9410 a_8912_37509.n19 VSS 1.31827f
C9411 a_8912_37509.n20 VSS 0.502978f
C9412 a_8912_37509.n21 VSS 0.453882f
C9413 a_8912_37509.n22 VSS 1.31827f
C9414 a_8912_37509.n23 VSS 0.475921f
C9415 a_8912_37509.t2 VSS 0.890777f
C9416 a_8912_37509.n24 VSS 1.31827f
C9417 a_8912_37509.n25 VSS 0.481525f
C9418 a_8912_37509.n26 VSS 0.330231f
C9419 a_8912_37509.n27 VSS 1.31827f
C9420 a_8912_37509.n28 VSS 0.308192f
C9421 a_8912_37509.t16 VSS 0.772205f
C9422 a_8912_37509.t6 VSS 0.177274f
C9423 a_8912_37509.t14 VSS 0.177274f
C9424 a_8912_37509.n29 VSS 0.48185f
C9425 a_8912_37509.n30 VSS 1.95207f
C9426 a_8912_37509.t13 VSS 0.177274f
C9427 a_8912_37509.t20 VSS 0.177274f
C9428 a_8912_37509.n31 VSS 0.48185f
C9429 a_8912_37509.n32 VSS 0.977562f
C9430 a_8912_37509.t21 VSS 0.177274f
C9431 a_8912_37509.t12 VSS 0.177274f
C9432 a_8912_37509.n33 VSS 0.48185f
C9433 a_8912_37509.n34 VSS 0.983166f
C9434 a_8912_37509.t8 VSS 0.76733f
C9435 a_8912_37509.n35 VSS 1.06904f
C9436 a_8912_37509.t24 VSS 0.76733f
C9437 a_8912_37509.n36 VSS 1.06344f
C9438 a_8912_37509.t23 VSS 0.177274f
C9439 a_8912_37509.t32 VSS 0.177274f
C9440 a_8912_37509.n37 VSS 0.48185f
C9441 a_8912_37509.n38 VSS 0.977562f
C9442 a_8912_37509.t33 VSS 0.177274f
C9443 a_8912_37509.t31 VSS 0.177274f
C9444 a_8912_37509.n39 VSS 0.48185f
C9445 a_8912_37509.n40 VSS 0.983166f
C9446 a_8912_37509.t37 VSS 0.177274f
C9447 a_8912_37509.t27 VSS 0.177274f
C9448 a_8912_37509.n41 VSS 0.48185f
C9449 a_8912_37509.n42 VSS 0.977562f
C9450 a_8912_37509.t29 VSS 0.76733f
C9451 a_8912_37509.n43 VSS 1.51956f
C9452 a_8912_37509.n44 VSS 0.736298f
C9453 a_8912_37509.n45 VSS 1.31827f
C9454 a_8912_37509.t0 VSS 0.890777f
C9455 a_5088_37509.t16 VSS 0.140614f
C9456 a_5088_37509.t10 VSS 0.140614f
C9457 a_5088_37509.n0 VSS 0.381085f
C9458 a_5088_37509.t8 VSS 0.140614f
C9459 a_5088_37509.t4 VSS 0.140614f
C9460 a_5088_37509.n1 VSS 0.376291f
C9461 a_5088_37509.n2 VSS 1.35312f
C9462 a_5088_37509.t18 VSS 0.140614f
C9463 a_5088_37509.t12 VSS 0.140614f
C9464 a_5088_37509.n3 VSS 0.376291f
C9465 a_5088_37509.n4 VSS 0.701585f
C9466 a_5088_37509.t17 VSS 0.140614f
C9467 a_5088_37509.t7 VSS 0.140614f
C9468 a_5088_37509.n5 VSS 0.376291f
C9469 a_5088_37509.n6 VSS 0.698353f
C9470 a_5088_37509.t11 VSS 0.140614f
C9471 a_5088_37509.t19 VSS 0.140614f
C9472 a_5088_37509.n7 VSS 0.364369f
C9473 a_5088_37509.t9 VSS 0.140614f
C9474 a_5088_37509.t15 VSS 0.140614f
C9475 a_5088_37509.n8 VSS 0.360133f
C9476 a_5088_37509.n9 VSS 1.18972f
C9477 a_5088_37509.t13 VSS 0.140614f
C9478 a_5088_37509.t5 VSS 0.140614f
C9479 a_5088_37509.n10 VSS 0.360133f
C9480 a_5088_37509.n11 VSS 0.619605f
C9481 a_5088_37509.t14 VSS 0.140614f
C9482 a_5088_37509.t6 VSS 0.140614f
C9483 a_5088_37509.n12 VSS 0.360133f
C9484 a_5088_37509.n13 VSS 1.42395f
C9485 a_5088_37509.n14 VSS 1.64996f
C9486 a_5088_37509.t3 VSS 0.193609f
C9487 a_5088_37509.n15 VSS 1.98688f
C9488 a_5088_37509.t1 VSS 0.194513f
C9489 a_5088_37509.n16 VSS 0.755758f
C9490 a_5088_37509.n17 VSS 0.121722f
C9491 VDAC_P.t1085 VSS 0.102851f
C9492 VDAC_P.t1050 VSS 0.102808f
C9493 VDAC_P.n0 VSS 0.114955f
C9494 VDAC_P.t90 VSS 0.102808f
C9495 VDAC_P.t456 VSS 0.102808f
C9496 VDAC_P.n2 VSS 0.113566f
C9497 VDAC_P.t320 VSS 0.102851f
C9498 VDAC_P.t2131 VSS 0.102808f
C9499 VDAC_P.n3 VSS 0.114955f
C9500 VDAC_P.t2091 VSS 0.102808f
C9501 VDAC_P.t1537 VSS 0.102808f
C9502 VDAC_P.t602 VSS 0.102843f
C9503 VDAC_P.t668 VSS 0.102808f
C9504 VDAC_P.n7 VSS 0.119912f
C9505 VDAC_P.t1081 VSS 0.102808f
C9506 VDAC_P.t221 VSS 0.102808f
C9507 VDAC_P.n9 VSS -0.13856f
C9508 VDAC_P.t2078 VSS 0.102808f
C9509 VDAC_P.t1087 VSS 0.102808f
C9510 VDAC_P.t165 VSS 0.102808f
C9511 VDAC_P.t941 VSS 0.102809f
C9512 VDAC_P.n14 VSS 0.422942f
C9513 VDAC_P.n15 VSS 0.267586f
C9514 VDAC_P.n16 VSS 0.261329f
C9515 VDAC_P.n17 VSS 0.368082f
C9516 VDAC_P.n18 VSS 0.267586f
C9517 VDAC_P.n19 VSS 0.261329f
C9518 VDAC_P.n20 VSS 0.368612f
C9519 VDAC_P.n21 VSS 0.372189f
C9520 VDAC_P.n22 VSS 2.31056f
C9521 VDAC_P.t599 VSS 0.10586f
C9522 VDAC_P.n23 VSS 0.137296f
C9523 VDAC_P.t694 VSS 0.10586f
C9524 VDAC_P.n24 VSS 0.12686f
C9525 VDAC_P.t1377 VSS 0.10586f
C9526 VDAC_P.n25 VSS 0.132855f
C9527 VDAC_P.t1586 VSS 0.10586f
C9528 VDAC_P.n26 VSS 0.132855f
C9529 VDAC_P.t1272 VSS 0.10586f
C9530 VDAC_P.n27 VSS 0.132855f
C9531 VDAC_P.t1026 VSS 0.10586f
C9532 VDAC_P.n28 VSS 0.132855f
C9533 VDAC_P.t1744 VSS 0.10586f
C9534 VDAC_P.n29 VSS 0.132855f
C9535 VDAC_P.t2117 VSS 0.10586f
C9536 VDAC_P.n30 VSS 0.132855f
C9537 VDAC_P.t670 VSS 0.10586f
C9538 VDAC_P.n31 VSS 0.132855f
C9539 VDAC_P.t1100 VSS 0.10586f
C9540 VDAC_P.n32 VSS 0.132855f
C9541 VDAC_P.t786 VSS 0.10586f
C9542 VDAC_P.n33 VSS 0.132855f
C9543 VDAC_P.t1152 VSS 0.10586f
C9544 VDAC_P.n34 VSS 0.132855f
C9545 VDAC_P.t517 VSS 0.10586f
C9546 VDAC_P.n35 VSS 0.132855f
C9547 VDAC_P.t824 VSS 0.10586f
C9548 VDAC_P.n36 VSS 0.132855f
C9549 VDAC_P.t285 VSS 0.10586f
C9550 VDAC_P.n37 VSS 0.132855f
C9551 VDAC_P.t1635 VSS 0.10586f
C9552 VDAC_P.n38 VSS 0.132855f
C9553 VDAC_P.t1212 VSS 0.10586f
C9554 VDAC_P.n39 VSS 0.132855f
C9555 VDAC_P.t455 VSS 0.10586f
C9556 VDAC_P.n40 VSS 0.132855f
C9557 VDAC_P.t2052 VSS 0.10586f
C9558 VDAC_P.n41 VSS 0.132855f
C9559 VDAC_P.t255 VSS 0.10586f
C9560 VDAC_P.n42 VSS 0.132855f
C9561 VDAC_P.t1385 VSS 0.10586f
C9562 VDAC_P.n43 VSS 0.132855f
C9563 VDAC_P.t535 VSS 0.10586f
C9564 VDAC_P.n44 VSS 0.132855f
C9565 VDAC_P.t225 VSS 0.10586f
C9566 VDAC_P.n45 VSS 0.132855f
C9567 VDAC_P.t2038 VSS 0.10586f
C9568 VDAC_P.n46 VSS 0.132855f
C9569 VDAC_P.t1627 VSS 0.10586f
C9570 VDAC_P.n47 VSS 0.132855f
C9571 VDAC_P.t171 VSS 0.10586f
C9572 VDAC_P.n48 VSS 0.132855f
C9573 VDAC_P.t1162 VSS 0.10586f
C9574 VDAC_P.n49 VSS 0.132855f
C9575 VDAC_P.t67 VSS 0.10586f
C9576 VDAC_P.n50 VSS 0.132855f
C9577 VDAC_P.t810 VSS 0.10586f
C9578 VDAC_P.n51 VSS 0.132855f
C9579 VDAC_P.t1381 VSS 0.10586f
C9580 VDAC_P.n52 VSS 0.132855f
C9581 VDAC_P.t474 VSS 0.10586f
C9582 VDAC_P.n53 VSS 0.132855f
C9583 VDAC_P.t1752 VSS 0.10586f
C9584 VDAC_P.n54 VSS 0.132855f
C9585 VDAC_P.t1145 VSS 0.10586f
C9586 VDAC_P.n55 VSS 0.132855f
C9587 VDAC_P.t162 VSS 0.10586f
C9588 VDAC_P.n56 VSS 0.132855f
C9589 VDAC_P.t300 VSS 0.10586f
C9590 VDAC_P.n57 VSS 0.132855f
C9591 VDAC_P.t1550 VSS 0.10586f
C9592 VDAC_P.n58 VSS 0.132855f
C9593 VDAC_P.t740 VSS 0.10586f
C9594 VDAC_P.n59 VSS 0.132855f
C9595 VDAC_P.t82 VSS 0.10586f
C9596 VDAC_P.n60 VSS 0.132855f
C9597 VDAC_P.t1640 VSS 0.10586f
C9598 VDAC_P.n61 VSS 0.132855f
C9599 VDAC_P.t1989 VSS 0.10586f
C9600 VDAC_P.n62 VSS 0.132855f
C9601 VDAC_P.t536 VSS 0.10586f
C9602 VDAC_P.n63 VSS 0.132855f
C9603 VDAC_P.t1276 VSS 0.10586f
C9604 VDAC_P.n64 VSS 0.132855f
C9605 VDAC_P.t885 VSS 0.10586f
C9606 VDAC_P.n65 VSS 0.132855f
C9607 VDAC_P.t1204 VSS 0.10586f
C9608 VDAC_P.n66 VSS 0.132855f
C9609 VDAC_P.t1847 VSS 0.10586f
C9610 VDAC_P.n67 VSS 0.132855f
C9611 VDAC_P.t120 VSS 0.10586f
C9612 VDAC_P.n68 VSS 0.132855f
C9613 VDAC_P.t1955 VSS 0.10586f
C9614 VDAC_P.n69 VSS 0.132855f
C9615 VDAC_P.t397 VSS 0.10586f
C9616 VDAC_P.n70 VSS 0.132855f
C9617 VDAC_P.t12 VSS 0.10586f
C9618 VDAC_P.n71 VSS 0.132855f
C9619 VDAC_P.t819 VSS 0.10586f
C9620 VDAC_P.n72 VSS 0.132855f
C9621 VDAC_P.t169 VSS 0.10586f
C9622 VDAC_P.n73 VSS 0.132855f
C9623 VDAC_P.t1123 VSS 0.10586f
C9624 VDAC_P.n74 VSS 0.132855f
C9625 VDAC_P.t1278 VSS 0.10586f
C9626 VDAC_P.n75 VSS 0.132855f
C9627 VDAC_P.t444 VSS 0.10586f
C9628 VDAC_P.n76 VSS 0.132855f
C9629 VDAC_P.t1510 VSS 0.10586f
C9630 VDAC_P.n77 VSS 0.132855f
C9631 VDAC_P.t560 VSS 0.10586f
C9632 VDAC_P.n78 VSS 0.132855f
C9633 VDAC_P.t870 VSS 0.10586f
C9634 VDAC_P.n79 VSS 0.132855f
C9635 VDAC_P.t1544 VSS 0.10586f
C9636 VDAC_P.n80 VSS 0.132855f
C9637 VDAC_P.t1049 VSS 0.10586f
C9638 VDAC_P.n81 VSS 0.132855f
C9639 VDAC_P.t272 VSS 0.10586f
C9640 VDAC_P.n82 VSS 0.132855f
C9641 VDAC_P.t26 VSS 0.10586f
C9642 VDAC_P.n83 VSS 0.132855f
C9643 VDAC_P.t875 VSS 0.10586f
C9644 VDAC_P.n84 VSS 0.132855f
C9645 VDAC_P.t980 VSS 0.10586f
C9646 VDAC_P.n85 VSS 0.132855f
C9647 VDAC_P.t1829 VSS 0.10586f
C9648 VDAC_P.n86 VSS 0.132855f
C9649 VDAC_P.t1408 VSS 0.10586f
C9650 VDAC_P.n87 VSS 0.12686f
C9651 VDAC_P.t241 VSS 0.10586f
C9652 VDAC_P.n88 VSS 0.12686f
C9653 VDAC_P.t718 VSS 0.10586f
C9654 VDAC_P.n89 VSS 0.12686f
C9655 VDAC_P.t2065 VSS 0.10586f
C9656 VDAC_P.n90 VSS 0.12686f
C9657 VDAC_P.t347 VSS 0.10586f
C9658 VDAC_P.n91 VSS 0.12686f
C9659 VDAC_P.t2036 VSS 0.10586f
C9660 VDAC_P.n92 VSS 0.12686f
C9661 VDAC_P.t431 VSS 0.10586f
C9662 VDAC_P.n93 VSS 0.12686f
C9663 VDAC_P.t1214 VSS 0.10586f
C9664 VDAC_P.n94 VSS 0.12686f
C9665 VDAC_P.t1003 VSS 0.10586f
C9666 VDAC_P.n95 VSS 0.12686f
C9667 VDAC_P.t621 VSS 0.10586f
C9668 VDAC_P.n96 VSS 0.12686f
C9669 VDAC_P.t1236 VSS 0.10586f
C9670 VDAC_P.n97 VSS 0.12686f
C9671 VDAC_P.t1549 VSS 0.10586f
C9672 VDAC_P.n98 VSS 0.12686f
C9673 VDAC_P.t2032 VSS 0.10586f
C9674 VDAC_P.n99 VSS 0.12686f
C9675 VDAC_P.t951 VSS 0.10586f
C9676 VDAC_P.n100 VSS 0.12686f
C9677 VDAC_P.t1115 VSS 0.10586f
C9678 VDAC_P.n101 VSS 0.12686f
C9679 VDAC_P.t956 VSS 0.10586f
C9680 VDAC_P.n102 VSS 0.12686f
C9681 VDAC_P.t117 VSS 0.10586f
C9682 VDAC_P.n103 VSS 0.12686f
C9683 VDAC_P.t500 VSS 0.10586f
C9684 VDAC_P.n104 VSS 0.12686f
C9685 VDAC_P.t53 VSS 0.10586f
C9686 VDAC_P.n105 VSS 0.12686f
C9687 VDAC_P.t1670 VSS 0.10586f
C9688 VDAC_P.n106 VSS 0.12686f
C9689 VDAC_P.t418 VSS 0.10586f
C9690 VDAC_P.n107 VSS 0.12686f
C9691 VDAC_P.t1581 VSS 0.10586f
C9692 VDAC_P.n108 VSS 0.12686f
C9693 VDAC_P.t1972 VSS 0.10586f
C9694 VDAC_P.n109 VSS 0.12686f
C9695 VDAC_P.t538 VSS 0.10586f
C9696 VDAC_P.n110 VSS 0.12686f
C9697 VDAC_P.t925 VSS 0.10586f
C9698 VDAC_P.n111 VSS 0.12686f
C9699 VDAC_P.t198 VSS 0.10586f
C9700 VDAC_P.n112 VSS 0.12686f
C9701 VDAC_P.t211 VSS 0.10586f
C9702 VDAC_P.n113 VSS 0.12686f
C9703 VDAC_P.t1376 VSS 0.10586f
C9704 VDAC_P.n114 VSS 0.12686f
C9705 VDAC_P.t591 VSS 0.10586f
C9706 VDAC_P.n115 VSS 0.12686f
C9707 VDAC_P.t87 VSS 0.10586f
C9708 VDAC_P.n116 VSS 0.12686f
C9709 VDAC_P.t1251 VSS 0.10586f
C9710 VDAC_P.n117 VSS 0.132855f
C9711 VDAC_P.t919 VSS 0.10586f
C9712 VDAC_P.n118 VSS 0.132855f
C9713 VDAC_P.t1147 VSS 0.10586f
C9714 VDAC_P.n119 VSS 0.132855f
C9715 VDAC_P.t421 VSS 0.10586f
C9716 VDAC_P.n120 VSS 0.132855f
C9717 VDAC_P.t1041 VSS 0.10586f
C9718 VDAC_P.n121 VSS 0.132855f
C9719 VDAC_P.t761 VSS 0.10586f
C9720 VDAC_P.n122 VSS 0.132855f
C9721 VDAC_P.t43 VSS 0.10586f
C9722 VDAC_P.n123 VSS 0.132855f
C9723 VDAC_P.t2020 VSS 0.10586f
C9724 VDAC_P.n124 VSS 0.132855f
C9725 VDAC_P.t933 VSS 0.10586f
C9726 VDAC_P.n125 VSS 0.132855f
C9727 VDAC_P.t164 VSS 0.10586f
C9728 VDAC_P.n126 VSS 0.132855f
C9729 VDAC_P.t1631 VSS 0.10586f
C9730 VDAC_P.n127 VSS 0.132855f
C9731 VDAC_P.t2134 VSS 0.10586f
C9732 VDAC_P.n128 VSS 0.132855f
C9733 VDAC_P.t152 VSS 0.10586f
C9734 VDAC_P.n129 VSS 0.132855f
C9735 VDAC_P.t1074 VSS 0.10586f
C9736 VDAC_P.n130 VSS 0.132855f
C9737 VDAC_P.t480 VSS 0.10586f
C9738 VDAC_P.n131 VSS 0.132855f
C9739 VDAC_P.t1046 VSS 0.10586f
C9740 VDAC_P.n132 VSS 0.132855f
C9741 VDAC_P.t704 VSS 0.10586f
C9742 VDAC_P.n133 VSS 0.132855f
C9743 VDAC_P.t430 VSS 0.10586f
C9744 VDAC_P.n134 VSS 0.132855f
C9745 VDAC_P.t713 VSS 0.10586f
C9746 VDAC_P.n135 VSS 0.132855f
C9747 VDAC_P.t202 VSS 0.10586f
C9748 VDAC_P.n136 VSS 0.132855f
C9749 VDAC_P.t1191 VSS 0.10586f
C9750 VDAC_P.n137 VSS 0.132855f
C9751 VDAC_P.t614 VSS 0.10586f
C9752 VDAC_P.n138 VSS 0.132855f
C9753 VDAC_P.t19 VSS 0.10586f
C9754 VDAC_P.n139 VSS 0.132855f
C9755 VDAC_P.t785 VSS 0.10586f
C9756 VDAC_P.n140 VSS 0.132855f
C9757 VDAC_P.t862 VSS 0.10586f
C9758 VDAC_P.n141 VSS 0.132855f
C9759 VDAC_P.t1429 VSS 0.10586f
C9760 VDAC_P.n142 VSS 0.132855f
C9761 VDAC_P.t1889 VSS 0.10586f
C9762 VDAC_P.n143 VSS 0.132855f
C9763 VDAC_P.t103 VSS 0.10586f
C9764 VDAC_P.n144 VSS 0.132855f
C9765 VDAC_P.t467 VSS 0.10586f
C9766 VDAC_P.n145 VSS 0.132855f
C9767 VDAC_P.t571 VSS 0.10586f
C9768 VDAC_P.n146 VSS 0.132855f
C9769 VDAC_P.t1573 VSS 0.10586f
C9770 VDAC_P.n147 VSS 0.132855f
C9771 VDAC_P.t2115 VSS 0.10586f
C9772 VDAC_P.n148 VSS 0.132855f
C9773 VDAC_P.t747 VSS 0.10586f
C9774 VDAC_P.n149 VSS 0.132855f
C9775 VDAC_P.t1917 VSS 0.10586f
C9776 VDAC_P.n150 VSS 0.132855f
C9777 VDAC_P.t1828 VSS 0.10586f
C9778 VDAC_P.n151 VSS 0.132855f
C9779 VDAC_P.t1811 VSS 0.10586f
C9780 VDAC_P.n152 VSS 0.132855f
C9781 VDAC_P.t908 VSS 0.10586f
C9782 VDAC_P.n153 VSS 0.132855f
C9783 VDAC_P.t1601 VSS 0.10586f
C9784 VDAC_P.n154 VSS 0.132855f
C9785 VDAC_P.t1436 VSS 0.10586f
C9786 VDAC_P.n155 VSS 0.132855f
C9787 VDAC_P.t1904 VSS 0.10586f
C9788 VDAC_P.n156 VSS 0.132855f
C9789 VDAC_P.t279 VSS 0.10586f
C9790 VDAC_P.n157 VSS 0.132855f
C9791 VDAC_P.t1808 VSS 0.10586f
C9792 VDAC_P.n158 VSS 0.132855f
C9793 VDAC_P.t1850 VSS 0.10586f
C9794 VDAC_P.n159 VSS 0.132855f
C9795 VDAC_P.t1860 VSS 0.10586f
C9796 VDAC_P.n160 VSS 0.132855f
C9797 VDAC_P.t1410 VSS 0.10586f
C9798 VDAC_P.n161 VSS 0.132855f
C9799 VDAC_P.t107 VSS 0.10586f
C9800 VDAC_P.n162 VSS 0.132855f
C9801 VDAC_P.t174 VSS 0.10586f
C9802 VDAC_P.n163 VSS 0.132855f
C9803 VDAC_P.t11 VSS 0.10586f
C9804 VDAC_P.n164 VSS 0.132855f
C9805 VDAC_P.t1920 VSS 0.10586f
C9806 VDAC_P.n165 VSS 0.132855f
C9807 VDAC_P.t970 VSS 0.10586f
C9808 VDAC_P.n166 VSS 0.132855f
C9809 VDAC_P.t727 VSS 0.10586f
C9810 VDAC_P.n167 VSS 0.132855f
C9811 VDAC_P.t1682 VSS 0.10586f
C9812 VDAC_P.n168 VSS 0.132855f
C9813 VDAC_P.t353 VSS 0.10586f
C9814 VDAC_P.n169 VSS 0.132855f
C9815 VDAC_P.t903 VSS 0.10586f
C9816 VDAC_P.n170 VSS 0.132855f
C9817 VDAC_P.t569 VSS 0.10586f
C9818 VDAC_P.n171 VSS 0.132855f
C9819 VDAC_P.t1679 VSS 0.10586f
C9820 VDAC_P.n172 VSS 0.132855f
C9821 VDAC_P.t998 VSS 0.10586f
C9822 VDAC_P.n173 VSS 0.132855f
C9823 VDAC_P.t1463 VSS 0.10586f
C9824 VDAC_P.n174 VSS 0.132855f
C9825 VDAC_P.t2025 VSS 0.10586f
C9826 VDAC_P.n175 VSS 0.132855f
C9827 VDAC_P.t1357 VSS 0.10586f
C9828 VDAC_P.n176 VSS 0.132855f
C9829 VDAC_P.t473 VSS 0.10586f
C9830 VDAC_P.n177 VSS 0.132855f
C9831 VDAC_P.t1764 VSS 0.10586f
C9832 VDAC_P.n178 VSS 0.132855f
C9833 VDAC_P.t447 VSS 0.10586f
C9834 VDAC_P.n179 VSS 0.12686f
C9835 VDAC_P.t1800 VSS 0.10586f
C9836 VDAC_P.n180 VSS 0.132855f
C9837 VDAC_P.t1038 VSS 0.10586f
C9838 VDAC_P.n181 VSS 0.132855f
C9839 VDAC_P.t1344 VSS 0.10586f
C9840 VDAC_P.n182 VSS 0.132855f
C9841 VDAC_P.t1622 VSS 0.10586f
C9842 VDAC_P.n183 VSS 0.132855f
C9843 VDAC_P.t657 VSS 0.10586f
C9844 VDAC_P.n184 VSS 0.132855f
C9845 VDAC_P.t1398 VSS 0.10586f
C9846 VDAC_P.n185 VSS 0.132855f
C9847 VDAC_P.t317 VSS 0.10586f
C9848 VDAC_P.n186 VSS 0.132855f
C9849 VDAC_P.t1639 VSS 0.10586f
C9850 VDAC_P.n187 VSS 0.132855f
C9851 VDAC_P.t158 VSS 0.10586f
C9852 VDAC_P.n188 VSS 0.132855f
C9853 VDAC_P.t1529 VSS 0.10586f
C9854 VDAC_P.n189 VSS 0.132855f
C9855 VDAC_P.t234 VSS 0.10586f
C9856 VDAC_P.n190 VSS 0.132855f
C9857 VDAC_P.t1419 VSS 0.10586f
C9858 VDAC_P.n191 VSS 0.132855f
C9859 VDAC_P.t1873 VSS 0.10586f
C9860 VDAC_P.n192 VSS 0.132855f
C9861 VDAC_P.t1953 VSS 0.10586f
C9862 VDAC_P.n193 VSS 0.132855f
C9863 VDAC_P.t1060 VSS 0.10586f
C9864 VDAC_P.n194 VSS 0.132855f
C9865 VDAC_P.t442 VSS 0.10586f
C9866 VDAC_P.n195 VSS 0.132855f
C9867 VDAC_P.t1188 VSS 0.10586f
C9868 VDAC_P.n196 VSS 0.132855f
C9869 VDAC_P.t1258 VSS 0.10586f
C9870 VDAC_P.n197 VSS 0.132855f
C9871 VDAC_P.t625 VSS 0.10586f
C9872 VDAC_P.n198 VSS 0.132855f
C9873 VDAC_P.t1040 VSS 0.10586f
C9874 VDAC_P.n199 VSS 0.132855f
C9875 VDAC_P.t1970 VSS 0.10586f
C9876 VDAC_P.n200 VSS 0.132855f
C9877 VDAC_P.t1624 VSS 0.10586f
C9878 VDAC_P.n201 VSS 0.132855f
C9879 VDAC_P.t1750 VSS 0.10586f
C9880 VDAC_P.n202 VSS 0.132855f
C9881 VDAC_P.t693 VSS 0.10586f
C9882 VDAC_P.n203 VSS 0.132855f
C9883 VDAC_P.t1318 VSS 0.10586f
C9884 VDAC_P.n204 VSS 0.132855f
C9885 VDAC_P.t333 VSS 0.10586f
C9886 VDAC_P.n205 VSS 0.132855f
C9887 VDAC_P.t1705 VSS 0.10586f
C9888 VDAC_P.n206 VSS 0.132855f
C9889 VDAC_P.t2034 VSS 0.10586f
C9890 VDAC_P.n207 VSS 0.132855f
C9891 VDAC_P.t77 VSS 0.10586f
C9892 VDAC_P.n208 VSS 0.132855f
C9893 VDAC_P.t1810 VSS 0.10586f
C9894 VDAC_P.n209 VSS 0.132855f
C9895 VDAC_P.t197 VSS 0.10586f
C9896 VDAC_P.n210 VSS 0.132855f
C9897 VDAC_P.t985 VSS 0.10586f
C9898 VDAC_P.n211 VSS 0.132855f
C9899 VDAC_P.t339 VSS 0.10586f
C9900 VDAC_P.n212 VSS 0.132855f
C9901 VDAC_P.t1729 VSS 0.10586f
C9902 VDAC_P.n213 VSS 0.132855f
C9903 VDAC_P.t92 VSS 0.10586f
C9904 VDAC_P.n214 VSS 0.132855f
C9905 VDAC_P.t1623 VSS 0.10586f
C9906 VDAC_P.n215 VSS 0.132855f
C9907 VDAC_P.t2081 VSS 0.10586f
C9908 VDAC_P.n216 VSS 0.132855f
C9909 VDAC_P.t1405 VSS 0.10586f
C9910 VDAC_P.n217 VSS 0.132855f
C9911 VDAC_P.t1001 VSS 0.10586f
C9912 VDAC_P.n218 VSS 0.132855f
C9913 VDAC_P.t1128 VSS 0.10586f
C9914 VDAC_P.n219 VSS 0.132855f
C9915 VDAC_P.t1841 VSS 0.10586f
C9916 VDAC_P.n220 VSS 0.132855f
C9917 VDAC_P.t1028 VSS 0.10586f
C9918 VDAC_P.n221 VSS 0.132855f
C9919 VDAC_P.t390 VSS 0.10586f
C9920 VDAC_P.n222 VSS 0.132855f
C9921 VDAC_P.t316 VSS 0.10586f
C9922 VDAC_P.n223 VSS 0.132855f
C9923 VDAC_P.t1032 VSS 0.10586f
C9924 VDAC_P.n224 VSS 0.132855f
C9925 VDAC_P.t1101 VSS 0.10586f
C9926 VDAC_P.n225 VSS 0.132855f
C9927 VDAC_P.t424 VSS 0.10586f
C9928 VDAC_P.n226 VSS 0.132855f
C9929 VDAC_P.t886 VSS 0.10586f
C9930 VDAC_P.n227 VSS 0.132855f
C9931 VDAC_P.t584 VSS 0.10586f
C9932 VDAC_P.n228 VSS 0.132855f
C9933 VDAC_P.t1538 VSS 0.10586f
C9934 VDAC_P.n229 VSS 0.132855f
C9935 VDAC_P.t637 VSS 0.10586f
C9936 VDAC_P.n230 VSS 0.132855f
C9937 VDAC_P.t346 VSS 0.10586f
C9938 VDAC_P.n231 VSS 0.132855f
C9939 VDAC_P.t1139 VSS 0.10586f
C9940 VDAC_P.n232 VSS 0.132855f
C9941 VDAC_P.t1591 VSS 0.10586f
C9942 VDAC_P.n233 VSS 0.132855f
C9943 VDAC_P.t1802 VSS 0.10586f
C9944 VDAC_P.n234 VSS 0.132855f
C9945 VDAC_P.t757 VSS 0.10586f
C9946 VDAC_P.n235 VSS 0.132855f
C9947 VDAC_P.t222 VSS 0.10586f
C9948 VDAC_P.n236 VSS 0.132855f
C9949 VDAC_P.t1269 VSS 0.10586f
C9950 VDAC_P.n237 VSS 0.132855f
C9951 VDAC_P.t253 VSS 0.10586f
C9952 VDAC_P.n238 VSS 0.132855f
C9953 VDAC_P.t1167 VSS 0.10586f
C9954 VDAC_P.n239 VSS 0.132855f
C9955 VDAC_P.t1621 VSS 0.10586f
C9956 VDAC_P.n240 VSS 0.132855f
C9957 VDAC_P.t540 VSS 0.10586f
C9958 VDAC_P.n241 VSS 0.132855f
C9959 VDAC_P.t771 VSS 0.10586f
C9960 VDAC_P.n242 VSS 0.12686f
C9961 VDAC_P.t35 VSS 0.10586f
C9962 VDAC_P.n243 VSS 0.132855f
C9963 VDAC_P.t948 VSS 0.10586f
C9964 VDAC_P.n244 VSS 0.132855f
C9965 VDAC_P.t1713 VSS 0.10586f
C9966 VDAC_P.n245 VSS 0.132855f
C9967 VDAC_P.t22 VSS 0.10586f
C9968 VDAC_P.n246 VSS 0.132855f
C9969 VDAC_P.t1936 VSS 0.10586f
C9970 VDAC_P.n247 VSS 0.132855f
C9971 VDAC_P.t1045 VSS 0.10586f
C9972 VDAC_P.n248 VSS 0.132855f
C9973 VDAC_P.t400 VSS 0.10586f
C9974 VDAC_P.n249 VSS 0.132855f
C9975 VDAC_P.t1694 VSS 0.10586f
C9976 VDAC_P.n250 VSS 0.132855f
C9977 VDAC_P.t2116 VSS 0.10586f
C9978 VDAC_P.n251 VSS 0.132855f
C9979 VDAC_P.t1490 VSS 0.10586f
C9980 VDAC_P.n252 VSS 0.132855f
C9981 VDAC_P.t1340 VSS 0.10586f
C9982 VDAC_P.n253 VSS 0.132855f
C9983 VDAC_P.t1262 VSS 0.10586f
C9984 VDAC_P.n254 VSS 0.132855f
C9985 VDAC_P.t1113 VSS 0.10586f
C9986 VDAC_P.n255 VSS 0.132855f
C9987 VDAC_P.t1763 VSS 0.10586f
C9988 VDAC_P.n256 VSS 0.132855f
C9989 VDAC_P.t2108 VSS 0.10586f
C9990 VDAC_P.n257 VSS 0.132855f
C9991 VDAC_P.t1302 VSS 0.10586f
C9992 VDAC_P.n258 VSS 0.132855f
C9993 VDAC_P.t2113 VSS 0.10586f
C9994 VDAC_P.n259 VSS 0.132855f
C9995 VDAC_P.t1736 VSS 0.10586f
C9996 VDAC_P.n260 VSS 0.132855f
C9997 VDAC_P.t2010 VSS 0.10586f
C9998 VDAC_P.n261 VSS 0.132855f
C9999 VDAC_P.t1256 VSS 0.10586f
C10000 VDAC_P.n262 VSS 0.132855f
C10001 VDAC_P.t1582 VSS 0.10586f
C10002 VDAC_P.n263 VSS 0.132855f
C10003 VDAC_P.t1636 VSS 0.10586f
C10004 VDAC_P.n264 VSS 0.132855f
C10005 VDAC_P.t1354 VSS 0.10586f
C10006 VDAC_P.n265 VSS 0.132855f
C10007 VDAC_P.t313 VSS 0.10586f
C10008 VDAC_P.n266 VSS 0.132855f
C10009 VDAC_P.t1840 VSS 0.10586f
C10010 VDAC_P.n267 VSS 0.132855f
C10011 VDAC_P.t2066 VSS 0.10586f
C10012 VDAC_P.n268 VSS 0.132855f
C10013 VDAC_P.t1515 VSS 0.10586f
C10014 VDAC_P.n269 VSS 0.132855f
C10015 VDAC_P.t1638 VSS 0.10586f
C10016 VDAC_P.n270 VSS 0.132855f
C10017 VDAC_P.t1399 VSS 0.10586f
C10018 VDAC_P.n271 VSS 0.132855f
C10019 VDAC_P.t1422 VSS 0.10586f
C10020 VDAC_P.n272 VSS 0.132855f
C10021 VDAC_P.t319 VSS 0.10586f
C10022 VDAC_P.n273 VSS 0.132855f
C10023 VDAC_P.t889 VSS 0.10586f
C10024 VDAC_P.n274 VSS 0.132855f
C10025 VDAC_P.t21 VSS 0.10586f
C10026 VDAC_P.n275 VSS 0.132855f
C10027 VDAC_P.t1543 VSS 0.10586f
C10028 VDAC_P.n276 VSS 0.132855f
C10029 VDAC_P.t521 VSS 0.10586f
C10030 VDAC_P.n277 VSS 0.132855f
C10031 VDAC_P.t729 VSS 0.10586f
C10032 VDAC_P.n278 VSS 0.132855f
C10033 VDAC_P.t959 VSS 0.10586f
C10034 VDAC_P.n279 VSS 0.132855f
C10035 VDAC_P.t1229 VSS 0.10586f
C10036 VDAC_P.n280 VSS 0.132855f
C10037 VDAC_P.t1785 VSS 0.10586f
C10038 VDAC_P.n281 VSS 0.132855f
C10039 VDAC_P.t1292 VSS 0.10586f
C10040 VDAC_P.n282 VSS 0.132855f
C10041 VDAC_P.t841 VSS 0.10586f
C10042 VDAC_P.n283 VSS 0.132855f
C10043 VDAC_P.t1852 VSS 0.10586f
C10044 VDAC_P.n284 VSS 0.132855f
C10045 VDAC_P.t1080 VSS 0.10586f
C10046 VDAC_P.n285 VSS 0.132855f
C10047 VDAC_P.t2005 VSS 0.10586f
C10048 VDAC_P.n286 VSS 0.132855f
C10049 VDAC_P.t632 VSS 0.10586f
C10050 VDAC_P.n287 VSS 0.132855f
C10051 VDAC_P.t1786 VSS 0.10586f
C10052 VDAC_P.n288 VSS 0.132855f
C10053 VDAC_P.t1588 VSS 0.10586f
C10054 VDAC_P.n289 VSS 0.132855f
C10055 VDAC_P.t1350 VSS 0.10586f
C10056 VDAC_P.n290 VSS 0.132855f
C10057 VDAC_P.t364 VSS 0.10586f
C10058 VDAC_P.n291 VSS 0.132855f
C10059 VDAC_P.t582 VSS 0.10586f
C10060 VDAC_P.n292 VSS 0.132855f
C10061 VDAC_P.t282 VSS 0.10586f
C10062 VDAC_P.n293 VSS 0.132855f
C10063 VDAC_P.t920 VSS 0.10586f
C10064 VDAC_P.n294 VSS 0.132855f
C10065 VDAC_P.t142 VSS 0.10586f
C10066 VDAC_P.n295 VSS 0.132855f
C10067 VDAC_P.t1395 VSS 0.10586f
C10068 VDAC_P.n296 VSS 0.132855f
C10069 VDAC_P.t374 VSS 0.10586f
C10070 VDAC_P.n297 VSS 0.132855f
C10071 VDAC_P.t661 VSS 0.10586f
C10072 VDAC_P.n298 VSS 0.132855f
C10073 VDAC_P.t1198 VSS 0.10586f
C10074 VDAC_P.n299 VSS 0.132855f
C10075 VDAC_P.t13 VSS 0.10586f
C10076 VDAC_P.n300 VSS 0.132855f
C10077 VDAC_P.t129 VSS 0.10586f
C10078 VDAC_P.n301 VSS 0.132855f
C10079 VDAC_P.t1914 VSS 0.10586f
C10080 VDAC_P.n302 VSS 0.132855f
C10081 VDAC_P.t1427 VSS 0.10586f
C10082 VDAC_P.n303 VSS 0.132855f
C10083 VDAC_P.t519 VSS 0.10586f
C10084 VDAC_P.n304 VSS 0.132855f
C10085 VDAC_P.t1329 VSS 0.10586f
C10086 VDAC_P.n305 VSS 0.12686f
C10087 VDAC_P.t1590 VSS 0.10586f
C10088 VDAC_P.n306 VSS 0.132855f
C10089 VDAC_P.t1379 VSS 0.10586f
C10090 VDAC_P.n307 VSS 0.132855f
C10091 VDAC_P.t1370 VSS 0.10586f
C10092 VDAC_P.n308 VSS 0.132855f
C10093 VDAC_P.t1171 VSS 0.10586f
C10094 VDAC_P.n309 VSS 0.132855f
C10095 VDAC_P.t827 VSS 0.10586f
C10096 VDAC_P.n310 VSS 0.132855f
C10097 VDAC_P.t30 VSS 0.10586f
C10098 VDAC_P.n311 VSS 0.132855f
C10099 VDAC_P.t401 VSS 0.10586f
C10100 VDAC_P.n312 VSS 0.132855f
C10101 VDAC_P.t1977 VSS 0.10586f
C10102 VDAC_P.n313 VSS 0.132855f
C10103 VDAC_P.t71 VSS 0.10586f
C10104 VDAC_P.n314 VSS 0.132855f
C10105 VDAC_P.t1861 VSS 0.10586f
C10106 VDAC_P.n315 VSS 0.132855f
C10107 VDAC_P.t613 VSS 0.10586f
C10108 VDAC_P.n316 VSS 0.132855f
C10109 VDAC_P.t1757 VSS 0.10586f
C10110 VDAC_P.n317 VSS 0.132855f
C10111 VDAC_P.t252 VSS 0.10586f
C10112 VDAC_P.n318 VSS 0.132855f
C10113 VDAC_P.t672 VSS 0.10586f
C10114 VDAC_P.n319 VSS 0.132855f
C10115 VDAC_P.t1610 VSS 0.10586f
C10116 VDAC_P.n320 VSS 0.132855f
C10117 VDAC_P.t367 VSS 0.10586f
C10118 VDAC_P.n321 VSS 0.132855f
C10119 VDAC_P.t706 VSS 0.10586f
C10120 VDAC_P.n322 VSS 0.132855f
C10121 VDAC_P.t1179 VSS 0.10586f
C10122 VDAC_P.n323 VSS 0.132855f
C10123 VDAC_P.t1735 VSS 0.10586f
C10124 VDAC_P.n324 VSS 0.132855f
C10125 VDAC_P.t1062 VSS 0.10586f
C10126 VDAC_P.n325 VSS 0.132855f
C10127 VDAC_P.t777 VSS 0.10586f
C10128 VDAC_P.n326 VSS 0.132855f
C10129 VDAC_P.t86 VSS 0.10586f
C10130 VDAC_P.n327 VSS 0.132855f
C10131 VDAC_P.t201 VSS 0.10586f
C10132 VDAC_P.n328 VSS 0.132855f
C10133 VDAC_P.t949 VSS 0.10586f
C10134 VDAC_P.n329 VSS 0.132855f
C10135 VDAC_P.t1209 VSS 0.10586f
C10136 VDAC_P.n330 VSS 0.132855f
C10137 VDAC_P.t245 VSS 0.10586f
C10138 VDAC_P.n331 VSS 0.132855f
C10139 VDAC_P.t556 VSS 0.10586f
C10140 VDAC_P.n332 VSS 0.132855f
C10141 VDAC_P.t1561 VSS 0.10586f
C10142 VDAC_P.n333 VSS 0.132855f
C10143 VDAC_P.t289 VSS 0.10586f
C10144 VDAC_P.n334 VSS 0.132855f
C10145 VDAC_P.t383 VSS 0.10586f
C10146 VDAC_P.n335 VSS 0.132855f
C10147 VDAC_P.t965 VSS 0.10586f
C10148 VDAC_P.n336 VSS 0.132855f
C10149 VDAC_P.t336 VSS 0.10586f
C10150 VDAC_P.n337 VSS 0.132855f
C10151 VDAC_P.t1797 VSS 0.10586f
C10152 VDAC_P.n338 VSS 0.132855f
C10153 VDAC_P.t1484 VSS 0.10586f
C10154 VDAC_P.n339 VSS 0.132855f
C10155 VDAC_P.t1158 VSS 0.10586f
C10156 VDAC_P.n340 VSS 0.132855f
C10157 VDAC_P.t2122 VSS 0.10586f
C10158 VDAC_P.n341 VSS 0.132855f
C10159 VDAC_P.t1848 VSS 0.10586f
C10160 VDAC_P.n342 VSS 0.132855f
C10161 VDAC_P.t1929 VSS 0.10586f
C10162 VDAC_P.n343 VSS 0.132855f
C10163 VDAC_P.t368 VSS 0.10586f
C10164 VDAC_P.n344 VSS 0.132855f
C10165 VDAC_P.t834 VSS 0.10586f
C10166 VDAC_P.n345 VSS 0.132855f
C10167 VDAC_P.t868 VSS 0.10586f
C10168 VDAC_P.n346 VSS 0.132855f
C10169 VDAC_P.t1594 VSS 0.10586f
C10170 VDAC_P.n347 VSS 0.132855f
C10171 VDAC_P.t1277 VSS 0.10586f
C10172 VDAC_P.n348 VSS 0.132855f
C10173 VDAC_P.t170 VSS 0.10586f
C10174 VDAC_P.n349 VSS 0.132855f
C10175 VDAC_P.t2082 VSS 0.10586f
C10176 VDAC_P.n350 VSS 0.132855f
C10177 VDAC_P.t1629 VSS 0.10586f
C10178 VDAC_P.n351 VSS 0.132855f
C10179 VDAC_P.t490 VSS 0.10586f
C10180 VDAC_P.n352 VSS 0.132855f
C10181 VDAC_P.t1407 VSS 0.10586f
C10182 VDAC_P.n353 VSS 0.132855f
C10183 VDAC_P.t1650 VSS 0.10586f
C10184 VDAC_P.n354 VSS 0.132855f
C10185 VDAC_P.t1309 VSS 0.10586f
C10186 VDAC_P.n355 VSS 0.132855f
C10187 VDAC_P.t1761 VSS 0.10586f
C10188 VDAC_P.n356 VSS 0.132855f
C10189 VDAC_P.t1201 VSS 0.10586f
C10190 VDAC_P.n357 VSS 0.132855f
C10191 VDAC_P.t843 VSS 0.10586f
C10192 VDAC_P.n358 VSS 0.132855f
C10193 VDAC_P.t2111 VSS 0.10586f
C10194 VDAC_P.n359 VSS 0.132855f
C10195 VDAC_P.t735 VSS 0.10586f
C10196 VDAC_P.n360 VSS 0.132855f
C10197 VDAC_P.t523 VSS 0.10586f
C10198 VDAC_P.n361 VSS 0.132855f
C10199 VDAC_P.t1339 VSS 0.10586f
C10200 VDAC_P.n362 VSS 0.132855f
C10201 VDAC_P.t911 VSS 0.10586f
C10202 VDAC_P.n363 VSS 0.132855f
C10203 VDAC_P.t1620 VSS 0.10586f
C10204 VDAC_P.n364 VSS 0.132855f
C10205 VDAC_P.t859 VSS 0.10586f
C10206 VDAC_P.n365 VSS 0.132855f
C10207 VDAC_P.t550 VSS 0.10586f
C10208 VDAC_P.n366 VSS 0.132855f
C10209 VDAC_P.t1142 VSS 0.10586f
C10210 VDAC_P.n367 VSS 0.132855f
C10211 VDAC_P.t2037 VSS 0.10586f
C10212 VDAC_P.n368 VSS 0.12686f
C10213 VDAC_P.t412 VSS 0.10586f
C10214 VDAC_P.n369 VSS 0.132855f
C10215 VDAC_P.t1174 VSS 0.10586f
C10216 VDAC_P.n370 VSS 0.132855f
C10217 VDAC_P.t2051 VSS 0.10586f
C10218 VDAC_P.n371 VSS 0.132855f
C10219 VDAC_P.t744 VSS 0.10586f
C10220 VDAC_P.n372 VSS 0.132855f
C10221 VDAC_P.t1666 VSS 0.10586f
C10222 VDAC_P.n373 VSS 0.132855f
C10223 VDAC_P.t276 VSS 0.10586f
C10224 VDAC_P.n374 VSS 0.132855f
C10225 VDAC_P.t1462 VSS 0.10586f
C10226 VDAC_P.n375 VSS 0.132855f
C10227 VDAC_P.t1211 VSS 0.10586f
C10228 VDAC_P.n376 VSS 0.132855f
C10229 VDAC_P.t634 VSS 0.10586f
C10230 VDAC_P.n377 VSS 0.132855f
C10231 VDAC_P.t1095 VSS 0.10586f
C10232 VDAC_P.n378 VSS 0.132855f
C10233 VDAC_P.t1584 VSS 0.10586f
C10234 VDAC_P.n379 VSS 0.132855f
C10235 VDAC_P.t58 VSS 0.10586f
C10236 VDAC_P.n380 VSS 0.132855f
C10237 VDAC_P.t739 VSS 0.10586f
C10238 VDAC_P.n381 VSS 0.132855f
C10239 VDAC_P.t1036 VSS 0.10586f
C10240 VDAC_P.n382 VSS 0.132855f
C10241 VDAC_P.t626 VSS 0.10586f
C10242 VDAC_P.n383 VSS 0.132855f
C10243 VDAC_P.t615 VSS 0.10586f
C10244 VDAC_P.n384 VSS 0.132855f
C10245 VDAC_P.t1984 VSS 0.10586f
C10246 VDAC_P.n385 VSS 0.132855f
C10247 VDAC_P.t982 VSS 0.10586f
C10248 VDAC_P.n386 VSS 0.132855f
C10249 VDAC_P.t1553 VSS 0.10586f
C10250 VDAC_P.n387 VSS 0.132855f
C10251 VDAC_P.t1714 VSS 0.10586f
C10252 VDAC_P.n388 VSS 0.132855f
C10253 VDAC_P.t69 VSS 0.10586f
C10254 VDAC_P.n389 VSS 0.132855f
C10255 VDAC_P.t398 VSS 0.10586f
C10256 VDAC_P.n390 VSS 0.132855f
C10257 VDAC_P.t631 VSS 0.10586f
C10258 VDAC_P.n391 VSS 0.132855f
C10259 VDAC_P.t1691 VSS 0.10586f
C10260 VDAC_P.n392 VSS 0.132855f
C10261 VDAC_P.t1010 VSS 0.10586f
C10262 VDAC_P.n393 VSS 0.132855f
C10263 VDAC_P.t803 VSS 0.10586f
C10264 VDAC_P.n394 VSS 0.132855f
C10265 VDAC_P.t1033 VSS 0.10586f
C10266 VDAC_P.n395 VSS 0.132855f
C10267 VDAC_P.t363 VSS 0.10586f
C10268 VDAC_P.n396 VSS 0.132855f
C10269 VDAC_P.t265 VSS 0.10586f
C10270 VDAC_P.n397 VSS 0.132855f
C10271 VDAC_P.t105 VSS 0.10586f
C10272 VDAC_P.n398 VSS 0.132855f
C10273 VDAC_P.t449 VSS 0.10586f
C10274 VDAC_P.n399 VSS 0.132855f
C10275 VDAC_P.t1868 VSS 0.10586f
C10276 VDAC_P.n400 VSS 0.132855f
C10277 VDAC_P.t1609 VSS 0.10586f
C10278 VDAC_P.n401 VSS 0.132855f
C10279 VDAC_P.t2061 VSS 0.10586f
C10280 VDAC_P.n402 VSS 0.132855f
C10281 VDAC_P.t768 VSS 0.10586f
C10282 VDAC_P.n403 VSS 0.132855f
C10283 VDAC_P.t991 VSS 0.10586f
C10284 VDAC_P.n404 VSS 0.132855f
C10285 VDAC_P.t548 VSS 0.10586f
C10286 VDAC_P.n405 VSS 0.132855f
C10287 VDAC_P.t1743 VSS 0.10586f
C10288 VDAC_P.n406 VSS 0.132855f
C10289 VDAC_P.t612 VSS 0.10586f
C10290 VDAC_P.n407 VSS 0.132855f
C10291 VDAC_P.t182 VSS 0.10586f
C10292 VDAC_P.n408 VSS 0.132855f
C10293 VDAC_P.t1308 VSS 0.10586f
C10294 VDAC_P.n409 VSS 0.132855f
C10295 VDAC_P.t618 VSS 0.10586f
C10296 VDAC_P.n410 VSS 0.132855f
C10297 VDAC_P.t1083 VSS 0.10586f
C10298 VDAC_P.n411 VSS 0.132855f
C10299 VDAC_P.t1528 VSS 0.10586f
C10300 VDAC_P.n412 VSS 0.132855f
C10301 VDAC_P.t1698 VSS 0.10586f
C10302 VDAC_P.n413 VSS 0.132855f
C10303 VDAC_P.t731 VSS 0.10586f
C10304 VDAC_P.n414 VSS 0.132855f
C10305 VDAC_P.t762 VSS 0.10586f
C10306 VDAC_P.n415 VSS 0.132855f
C10307 VDAC_P.t629 VSS 0.10586f
C10308 VDAC_P.n416 VSS 0.132855f
C10309 VDAC_P.t338 VSS 0.10586f
C10310 VDAC_P.n417 VSS 0.132855f
C10311 VDAC_P.t45 VSS 0.10586f
C10312 VDAC_P.n418 VSS 0.132855f
C10313 VDAC_P.t1575 VSS 0.10586f
C10314 VDAC_P.n419 VSS 0.132855f
C10315 VDAC_P.t1974 VSS 0.10586f
C10316 VDAC_P.n420 VSS 0.132855f
C10317 VDAC_P.t1469 VSS 0.10586f
C10318 VDAC_P.n421 VSS 0.132855f
C10319 VDAC_P.t1921 VSS 0.10586f
C10320 VDAC_P.n422 VSS 0.132855f
C10321 VDAC_P.t1255 VSS 0.10586f
C10322 VDAC_P.n423 VSS 0.132855f
C10323 VDAC_P.t921 VSS 0.10586f
C10324 VDAC_P.n424 VSS 0.132855f
C10325 VDAC_P.t309 VSS 0.10586f
C10326 VDAC_P.n425 VSS 0.132855f
C10327 VDAC_P.t817 VSS 0.10586f
C10328 VDAC_P.n426 VSS 0.132855f
C10329 VDAC_P.t1820 VSS 0.10586f
C10330 VDAC_P.n427 VSS 0.132855f
C10331 VDAC_P.t51 VSS 0.10586f
C10332 VDAC_P.n428 VSS 0.132855f
C10333 VDAC_P.t509 VSS 0.10586f
C10334 VDAC_P.n429 VSS 0.132855f
C10335 VDAC_P.t1480 VSS 0.10586f
C10336 VDAC_P.n430 VSS 0.132855f
C10337 VDAC_P.t1843 VSS 0.10586f
C10338 VDAC_P.n431 VSS 0.12686f
C10339 VDAC_P.t1157 VSS 0.10586f
C10340 VDAC_P.n432 VSS 0.132855f
C10341 VDAC_P.t871 VSS 0.10586f
C10342 VDAC_P.n433 VSS 0.132855f
C10343 VDAC_P.t534 VSS 0.10586f
C10344 VDAC_P.n434 VSS 0.132855f
C10345 VDAC_P.t1507 VSS 0.10586f
C10346 VDAC_P.n435 VSS 0.132855f
C10347 VDAC_P.t993 VSS 0.10586f
C10348 VDAC_P.n436 VSS 0.132855f
C10349 VDAC_P.t1389 VSS 0.10586f
C10350 VDAC_P.n437 VSS 0.132855f
C10351 VDAC_P.t1849 VSS 0.10586f
C10352 VDAC_P.n438 VSS 0.132855f
C10353 VDAC_P.t1220 VSS 0.10586f
C10354 VDAC_P.n439 VSS 0.132855f
C10355 VDAC_P.t457 VSS 0.10586f
C10356 VDAC_P.n440 VSS 0.132855f
C10357 VDAC_P.t700 VSS 0.10586f
C10358 VDAC_P.n441 VSS 0.132855f
C10359 VDAC_P.t1531 VSS 0.10586f
C10360 VDAC_P.n442 VSS 0.132855f
C10361 VDAC_P.t1059 VSS 0.10586f
C10362 VDAC_P.n443 VSS 0.132855f
C10363 VDAC_P.t1648 VSS 0.10586f
C10364 VDAC_P.n444 VSS 0.132855f
C10365 VDAC_P.t458 VSS 0.10586f
C10366 VDAC_P.n445 VSS 0.132855f
C10367 VDAC_P.t1353 VSS 0.10586f
C10368 VDAC_P.n446 VSS 0.132855f
C10369 VDAC_P.t1911 VSS 0.10586f
C10370 VDAC_P.n447 VSS 0.132855f
C10371 VDAC_P.t1247 VSS 0.10586f
C10372 VDAC_P.n448 VSS 0.132855f
C10373 VDAC_P.t1701 VSS 0.10586f
C10374 VDAC_P.n449 VSS 0.132855f
C10375 VDAC_P.t1612 VSS 0.10586f
C10376 VDAC_P.n450 VSS 0.132855f
C10377 VDAC_P.t1593 VSS 0.10586f
C10378 VDAC_P.n451 VSS 0.132855f
C10379 VDAC_P.t2047 VSS 0.10586f
C10380 VDAC_P.n452 VSS 0.132855f
C10381 VDAC_P.t393 VSS 0.10586f
C10382 VDAC_P.n453 VSS 0.132855f
C10383 VDAC_P.t267 VSS 0.10586f
C10384 VDAC_P.n454 VSS 0.132855f
C10385 VDAC_P.t516 VSS 0.10586f
C10386 VDAC_P.n455 VSS 0.132855f
C10387 VDAC_P.t453 VSS 0.10586f
C10388 VDAC_P.n456 VSS 0.132855f
C10389 VDAC_P.t44 VSS 0.10586f
C10390 VDAC_P.n457 VSS 0.132855f
C10391 VDAC_P.t1230 VSS 0.10586f
C10392 VDAC_P.n458 VSS 0.132855f
C10393 VDAC_P.t1053 VSS 0.10586f
C10394 VDAC_P.n459 VSS 0.132855f
C10395 VDAC_P.t1008 VSS 0.10586f
C10396 VDAC_P.n460 VSS 0.132855f
C10397 VDAC_P.t1973 VSS 0.10586f
C10398 VDAC_P.n461 VSS 0.132855f
C10399 VDAC_P.t576 VSS 0.10586f
C10400 VDAC_P.n462 VSS 0.132855f
C10401 VDAC_P.t1718 VSS 0.10586f
C10402 VDAC_P.n463 VSS 0.132855f
C10403 VDAC_P.t356 VSS 0.10586f
C10404 VDAC_P.n464 VSS 0.132855f
C10405 VDAC_P.t1290 VSS 0.10586f
C10406 VDAC_P.n465 VSS 0.132855f
C10407 VDAC_P.t1129 VSS 0.10586f
C10408 VDAC_P.n466 VSS 0.132855f
C10409 VDAC_P.t2112 VSS 0.10586f
C10410 VDAC_P.n467 VSS 0.132855f
C10411 VDAC_P.t1014 VSS 0.10586f
C10412 VDAC_P.n468 VSS 0.132855f
C10413 VDAC_P.t1224 VSS 0.10586f
C10414 VDAC_P.n469 VSS 0.132855f
C10415 VDAC_P.t1774 VSS 0.10586f
C10416 VDAC_P.n470 VSS 0.132855f
C10417 VDAC_P.t699 VSS 0.10586f
C10418 VDAC_P.n471 VSS 0.132855f
C10419 VDAC_P.t782 VSS 0.10586f
C10420 VDAC_P.n472 VSS 0.132855f
C10421 VDAC_P.t1345 VSS 0.10586f
C10422 VDAC_P.n473 VSS 0.132855f
C10423 VDAC_P.t1801 VSS 0.10586f
C10424 VDAC_P.n474 VSS 0.132855f
C10425 VDAC_P.t583 VSS 0.10586f
C10426 VDAC_P.n475 VSS 0.132855f
C10427 VDAC_P.t1587 VSS 0.10586f
C10428 VDAC_P.n476 VSS 0.132855f
C10429 VDAC_P.t1500 VSS 0.10586f
C10430 VDAC_P.n477 VSS 0.132855f
C10431 VDAC_P.t755 VSS 0.10586f
C10432 VDAC_P.n478 VSS 0.132855f
C10433 VDAC_P.t505 VSS 0.10586f
C10434 VDAC_P.n479 VSS 0.132855f
C10435 VDAC_P.t49 VSS 0.10586f
C10436 VDAC_P.n480 VSS 0.132855f
C10437 VDAC_P.t1825 VSS 0.10586f
C10438 VDAC_P.n481 VSS 0.132855f
C10439 VDAC_P.t1996 VSS 0.10586f
C10440 VDAC_P.n482 VSS 0.132855f
C10441 VDAC_P.t873 VSS 0.10586f
C10442 VDAC_P.n483 VSS 0.132855f
C10443 VDAC_P.t24 VSS 0.10586f
C10444 VDAC_P.n484 VSS 0.132855f
C10445 VDAC_P.t1968 VSS 0.10586f
C10446 VDAC_P.n485 VSS 0.132855f
C10447 VDAC_P.t1967 VSS 0.10586f
C10448 VDAC_P.n486 VSS 0.132855f
C10449 VDAC_P.t216 VSS 0.10586f
C10450 VDAC_P.n487 VSS 0.132855f
C10451 VDAC_P.t1855 VSS 0.10586f
C10452 VDAC_P.n488 VSS 0.132855f
C10453 VDAC_P.t1300 VSS 0.10586f
C10454 VDAC_P.n489 VSS 0.132855f
C10455 VDAC_P.t74 VSS 0.10586f
C10456 VDAC_P.n490 VSS 0.132855f
C10457 VDAC_P.t828 VSS 0.10586f
C10458 VDAC_P.n491 VSS 0.132855f
C10459 VDAC_P.t2096 VSS 0.10586f
C10460 VDAC_P.n492 VSS 0.132855f
C10461 VDAC_P.t573 VSS 0.10586f
C10462 VDAC_P.n493 VSS 0.132855f
C10463 VDAC_P.t440 VSS 0.10586f
C10464 VDAC_P.n494 VSS 0.12686f
C10465 VDAC_P.t1384 VSS 0.10586f
C10466 VDAC_P.n495 VSS 0.132855f
C10467 VDAC_P.t1858 VSS 0.10586f
C10468 VDAC_P.n496 VSS 0.132855f
C10469 VDAC_P.t1892 VSS 0.10586f
C10470 VDAC_P.n497 VSS 0.132855f
C10471 VDAC_P.t726 VSS 0.10586f
C10472 VDAC_P.n498 VSS 0.132855f
C10473 VDAC_P.t1193 VSS 0.10586f
C10474 VDAC_P.n499 VSS 0.132855f
C10475 VDAC_P.t322 VSS 0.10586f
C10476 VDAC_P.n500 VSS 0.132855f
C10477 VDAC_P.t23 VSS 0.10586f
C10478 VDAC_P.n501 VSS 0.132855f
C10479 VDAC_P.t1545 VSS 0.10586f
C10480 VDAC_P.n502 VSS 0.132855f
C10481 VDAC_P.t974 VSS 0.10586f
C10482 VDAC_P.n503 VSS 0.132855f
C10483 VDAC_P.t1431 VSS 0.10586f
C10484 VDAC_P.n504 VSS 0.132855f
C10485 VDAC_P.t394 VSS 0.10586f
C10486 VDAC_P.n505 VSS 0.132855f
C10487 VDAC_P.t191 VSS 0.10586f
C10488 VDAC_P.n506 VSS 0.132855f
C10489 VDAC_P.t907 VSS 0.10586f
C10490 VDAC_P.n507 VSS 0.132855f
C10491 VDAC_P.t690 VSS 0.10586f
C10492 VDAC_P.n508 VSS 0.132855f
C10493 VDAC_P.t1165 VSS 0.10586f
C10494 VDAC_P.n509 VSS 0.132855f
C10495 VDAC_P.t1719 VSS 0.10586f
C10496 VDAC_P.n510 VSS 0.132855f
C10497 VDAC_P.t2062 VSS 0.10586f
C10498 VDAC_P.n511 VSS 0.132855f
C10499 VDAC_P.t1513 VSS 0.10586f
C10500 VDAC_P.n512 VSS 0.132855f
C10501 VDAC_P.t1047 VSS 0.10586f
C10502 VDAC_P.n513 VSS 0.132855f
C10503 VDAC_P.t1397 VSS 0.10586f
C10504 VDAC_P.n514 VSS 0.132855f
C10505 VDAC_P.t485 VSS 0.10586f
C10506 VDAC_P.n515 VSS 0.132855f
C10507 VDAC_P.t1297 VSS 0.10586f
C10508 VDAC_P.n516 VSS 0.132855f
C10509 VDAC_P.t1749 VSS 0.10586f
C10510 VDAC_P.n517 VSS 0.132855f
C10511 VDAC_P.t1660 VSS 0.10586f
C10512 VDAC_P.n518 VSS 0.132855f
C10513 VDAC_P.t1541 VSS 0.10586f
C10514 VDAC_P.n519 VSS 0.132855f
C10515 VDAC_P.t545 VSS 0.10586f
C10516 VDAC_P.n520 VSS 0.132855f
C10517 VDAC_P.t1680 VSS 0.10586f
C10518 VDAC_P.n521 VSS 0.132855f
C10519 VDAC_P.t493 VSS 0.10586f
C10520 VDAC_P.n522 VSS 0.132855f
C10521 VDAC_P.t1200 VSS 0.10586f
C10522 VDAC_P.n523 VSS 0.132855f
C10523 VDAC_P.t1783 VSS 0.10586f
C10524 VDAC_P.n524 VSS 0.132855f
C10525 VDAC_P.t652 VSS 0.10586f
C10526 VDAC_P.n525 VSS 0.132855f
C10527 VDAC_P.t354 VSS 0.10586f
C10528 VDAC_P.n526 VSS 0.132855f
C10529 VDAC_P.t2106 VSS 0.10586f
C10530 VDAC_P.n527 VSS 0.132855f
C10531 VDAC_P.t1792 VSS 0.10586f
C10532 VDAC_P.n528 VSS 0.132855f
C10533 VDAC_P.t1834 VSS 0.10586f
C10534 VDAC_P.n529 VSS 0.132855f
C10535 VDAC_P.t352 VSS 0.10586f
C10536 VDAC_P.n530 VSS 0.132855f
C10537 VDAC_P.t1618 VSS 0.10586f
C10538 VDAC_P.n531 VSS 0.132855f
C10539 VDAC_P.t1772 VSS 0.10586f
C10540 VDAC_P.n532 VSS 0.132855f
C10541 VDAC_P.t1390 VSS 0.10586f
C10542 VDAC_P.n533 VSS 0.132855f
C10543 VDAC_P.t605 VSS 0.10586f
C10544 VDAC_P.n534 VSS 0.132855f
C10545 VDAC_P.t166 VSS 0.10586f
C10546 VDAC_P.n535 VSS 0.132855f
C10547 VDAC_P.t1159 VSS 0.10586f
C10548 VDAC_P.n536 VSS 0.132855f
C10549 VDAC_P.t821 VSS 0.10586f
C10550 VDAC_P.n537 VSS 0.132855f
C10551 VDAC_P.t938 VSS 0.10586f
C10552 VDAC_P.n538 VSS 0.132855f
C10553 VDAC_P.t369 VSS 0.10586f
C10554 VDAC_P.n539 VSS 0.132855f
C10555 VDAC_P.t1959 VSS 0.10586f
C10556 VDAC_P.n540 VSS 0.132855f
C10557 VDAC_P.t1291 VSS 0.10586f
C10558 VDAC_P.n541 VSS 0.132855f
C10559 VDAC_P.t1747 VSS 0.10586f
C10560 VDAC_P.n542 VSS 0.132855f
C10561 VDAC_P.t607 VSS 0.10586f
C10562 VDAC_P.n543 VSS 0.132855f
C10563 VDAC_P.t1643 VSS 0.10586f
C10564 VDAC_P.n544 VSS 0.132855f
C10565 VDAC_P.t1061 VSS 0.10586f
C10566 VDAC_P.n545 VSS 0.132855f
C10567 VDAC_P.t75 VSS 0.10586f
C10568 VDAC_P.n546 VSS 0.132855f
C10569 VDAC_P.t1991 VSS 0.10586f
C10570 VDAC_P.n547 VSS 0.132855f
C10571 VDAC_P.t64 VSS 0.10586f
C10572 VDAC_P.n548 VSS 0.132855f
C10573 VDAC_P.t465 VSS 0.10586f
C10574 VDAC_P.n549 VSS 0.132855f
C10575 VDAC_P.t1476 VSS 0.10586f
C10576 VDAC_P.n550 VSS 0.132855f
C10577 VDAC_P.t1677 VSS 0.10586f
C10578 VDAC_P.n551 VSS 0.132855f
C10579 VDAC_P.t1079 VSS 0.10586f
C10580 VDAC_P.n552 VSS 0.132855f
C10581 VDAC_P.t566 VSS 0.10586f
C10582 VDAC_P.n553 VSS 0.132855f
C10583 VDAC_P.t2023 VSS 0.10586f
C10584 VDAC_P.n554 VSS 0.132855f
C10585 VDAC_P.t1312 VSS 0.10586f
C10586 VDAC_P.n555 VSS 0.132855f
C10587 VDAC_P.t1814 VSS 0.10586f
C10588 VDAC_P.n556 VSS 0.132855f
C10589 VDAC_P.t1748 VSS 0.10586f
C10590 VDAC_P.n557 VSS 0.12686f
C10591 VDAC_P.t1727 VSS 0.10586f
C10592 VDAC_P.n558 VSS 0.132855f
C10593 VDAC_P.t2060 VSS 0.10586f
C10594 VDAC_P.n559 VSS 0.132855f
C10595 VDAC_P.t825 VSS 0.10586f
C10596 VDAC_P.n560 VSS 0.132855f
C10597 VDAC_P.t2077 VSS 0.10586f
C10598 VDAC_P.n561 VSS 0.132855f
C10599 VDAC_P.t40 VSS 0.10586f
C10600 VDAC_P.n562 VSS 0.132855f
C10601 VDAC_P.t271 VSS 0.10586f
C10602 VDAC_P.n563 VSS 0.132855f
C10603 VDAC_P.t96 VSS 0.10586f
C10604 VDAC_P.n564 VSS 0.132855f
C10605 VDAC_P.t1518 VSS 0.10586f
C10606 VDAC_P.n565 VSS 0.132855f
C10607 VDAC_P.t1332 VSS 0.10586f
C10608 VDAC_P.n566 VSS 0.132855f
C10609 VDAC_P.t1286 VSS 0.10586f
C10610 VDAC_P.n567 VSS 0.132855f
C10611 VDAC_P.t2103 VSS 0.10586f
C10612 VDAC_P.n568 VSS 0.132855f
C10613 VDAC_P.t288 VSS 0.10586f
C10614 VDAC_P.n569 VSS 0.132855f
C10615 VDAC_P.t274 VSS 0.10586f
C10616 VDAC_P.n570 VSS 0.132855f
C10617 VDAC_P.t264 VSS 0.10586f
C10618 VDAC_P.n571 VSS 0.132855f
C10619 VDAC_P.t1910 VSS 0.10586f
C10620 VDAC_P.n572 VSS 0.132855f
C10621 VDAC_P.t1533 VSS 0.10586f
C10622 VDAC_P.n573 VSS 0.132855f
C10623 VDAC_P.t854 VSS 0.10586f
C10624 VDAC_P.n574 VSS 0.132855f
C10625 VDAC_P.t1327 VSS 0.10586f
C10626 VDAC_P.n575 VSS 0.132855f
C10627 VDAC_P.t259 VSS 0.10586f
C10628 VDAC_P.n576 VSS 0.132855f
C10629 VDAC_P.t1221 VSS 0.10586f
C10630 VDAC_P.n577 VSS 0.132855f
C10631 VDAC_P.t853 VSS 0.10586f
C10632 VDAC_P.n578 VSS 0.132855f
C10633 VDAC_P.t297 VSS 0.10586f
C10634 VDAC_P.n579 VSS 0.132855f
C10635 VDAC_P.t797 VSS 0.10586f
C10636 VDAC_P.n580 VSS 0.132855f
C10637 VDAC_P.t527 VSS 0.10586f
C10638 VDAC_P.n581 VSS 0.132855f
C10639 VDAC_P.t1355 VSS 0.10586f
C10640 VDAC_P.n582 VSS 0.132855f
C10641 VDAC_P.t499 VSS 0.10586f
C10642 VDAC_P.n583 VSS 0.132855f
C10643 VDAC_P.t244 VSS 0.10586f
C10644 VDAC_P.n584 VSS 0.132855f
C10645 VDAC_P.t1703 VSS 0.10586f
C10646 VDAC_P.n585 VSS 0.132855f
C10647 VDAC_P.t428 VSS 0.10586f
C10648 VDAC_P.n586 VSS 0.132855f
C10649 VDAC_P.t1595 VSS 0.10586f
C10650 VDAC_P.n587 VSS 0.132855f
C10651 VDAC_P.t2049 VSS 0.10586f
C10652 VDAC_P.n588 VSS 0.132855f
C10653 VDAC_P.t488 VSS 0.10586f
C10654 VDAC_P.n589 VSS 0.132855f
C10655 VDAC_P.t1941 VSS 0.10586f
C10656 VDAC_P.n590 VSS 0.132855f
C10657 VDAC_P.t1012 VSS 0.10586f
C10658 VDAC_P.n591 VSS 0.132855f
C10659 VDAC_P.t1454 VSS 0.10586f
C10660 VDAC_P.n592 VSS 0.132855f
C10661 VDAC_P.t2092 VSS 0.10586f
C10662 VDAC_P.n593 VSS 0.132855f
C10663 VDAC_P.t1234 VSS 0.10586f
C10664 VDAC_P.n594 VSS 0.132855f
C10665 VDAC_P.t541 VSS 0.10586f
C10666 VDAC_P.n595 VSS 0.132855f
C10667 VDAC_P.t1992 VSS 0.10586f
C10668 VDAC_P.n596 VSS 0.132855f
C10669 VDAC_P.t1942 VSS 0.10586f
C10670 VDAC_P.n597 VSS 0.132855f
C10671 VDAC_P.t752 VSS 0.10586f
C10672 VDAC_P.n598 VSS 0.132855f
C10673 VDAC_P.t962 VSS 0.10586f
C10674 VDAC_P.n599 VSS 0.132855f
C10675 VDAC_P.t115 VSS 0.10586f
C10676 VDAC_P.n600 VSS 0.132855f
C10677 VDAC_P.t1474 VSS 0.10586f
C10678 VDAC_P.n601 VSS 0.132855f
C10679 VDAC_P.t1217 VSS 0.10586f
C10680 VDAC_P.n602 VSS 0.132855f
C10681 VDAC_P.t463 VSS 0.10586f
C10682 VDAC_P.n603 VSS 0.132855f
C10683 VDAC_P.t1099 VSS 0.10586f
C10684 VDAC_P.n604 VSS 0.132855f
C10685 VDAC_P.t1563 VSS 0.10586f
C10686 VDAC_P.n605 VSS 0.132855f
C10687 VDAC_P.t510 VSS 0.10586f
C10688 VDAC_P.n606 VSS 0.132855f
C10689 VDAC_P.t1455 VSS 0.10586f
C10690 VDAC_P.n607 VSS 0.132855f
C10691 VDAC_P.t1907 VSS 0.10586f
C10692 VDAC_P.n608 VSS 0.132855f
C10693 VDAC_P.t687 VSS 0.10586f
C10694 VDAC_P.n609 VSS 0.132855f
C10695 VDAC_P.t915 VSS 0.10586f
C10696 VDAC_P.n610 VSS 0.132855f
C10697 VDAC_P.t76 VSS 0.10586f
C10698 VDAC_P.n611 VSS 0.132855f
C10699 VDAC_P.t223 VSS 0.10586f
C10700 VDAC_P.n612 VSS 0.132855f
C10701 VDAC_P.t732 VSS 0.10586f
C10702 VDAC_P.n613 VSS 0.132855f
C10703 VDAC_P.t1485 VSS 0.10586f
C10704 VDAC_P.n614 VSS 0.132855f
C10705 VDAC_P.t1937 VSS 0.10586f
C10706 VDAC_P.n615 VSS 0.132855f
C10707 VDAC_P.t200 VSS 0.10586f
C10708 VDAC_P.n616 VSS 0.132855f
C10709 VDAC_P.t1827 VSS 0.10586f
C10710 VDAC_P.n617 VSS 0.132855f
C10711 VDAC_P.t2028 VSS 0.10586f
C10712 VDAC_P.n618 VSS 0.132855f
C10713 VDAC_P.t50 VSS 0.10586f
C10714 VDAC_P.n619 VSS 0.132855f
C10715 VDAC_P.t1884 VSS 0.10586f
C10716 VDAC_P.n620 VSS 0.12686f
C10717 VDAC_P.t906 VSS 0.10586f
C10718 VDAC_P.n621 VSS 0.132855f
C10719 VDAC_P.t1477 VSS 0.10586f
C10720 VDAC_P.n622 VSS 0.132855f
C10721 VDAC_P.t1570 VSS 0.10586f
C10722 VDAC_P.n623 VSS 0.132855f
C10723 VDAC_P.t337 VSS 0.10586f
C10724 VDAC_P.n624 VSS 0.132855f
C10725 VDAC_P.t239 VSS 0.10586f
C10726 VDAC_P.n625 VSS 0.132855f
C10727 VDAC_P.t311 VSS 0.10586f
C10728 VDAC_P.n626 VSS 0.132855f
C10729 VDAC_P.t1615 VSS 0.10586f
C10730 VDAC_P.n627 VSS 0.132855f
C10731 VDAC_P.t537 VSS 0.10586f
C10732 VDAC_P.n628 VSS 0.132855f
C10733 VDAC_P.t213 VSS 0.10586f
C10734 VDAC_P.n629 VSS 0.132855f
C10735 VDAC_P.t511 VSS 0.10586f
C10736 VDAC_P.n630 VSS 0.132855f
C10737 VDAC_P.t1293 VSS 0.10586f
C10738 VDAC_P.n631 VSS 0.132855f
C10739 VDAC_P.t939 VSS 0.10586f
C10740 VDAC_P.n632 VSS 0.132855f
C10741 VDAC_P.t628 VSS 0.10586f
C10742 VDAC_P.n633 VSS 0.132855f
C10743 VDAC_P.t609 VSS 0.10586f
C10744 VDAC_P.n634 VSS 0.132855f
C10745 VDAC_P.t839 VSS 0.10586f
C10746 VDAC_P.n635 VSS 0.132855f
C10747 VDAC_P.t1596 VSS 0.10586f
C10748 VDAC_P.n636 VSS 0.132855f
C10749 VDAC_P.t217 VSS 0.10586f
C10750 VDAC_P.n637 VSS 0.132855f
C10751 VDAC_P.t1013 VSS 0.10586f
C10752 VDAC_P.n638 VSS 0.132855f
C10753 VDAC_P.t1672 VSS 0.10586f
C10754 VDAC_P.n639 VSS 0.132855f
C10755 VDAC_P.t1887 VSS 0.10586f
C10756 VDAC_P.n640 VSS 0.132855f
C10757 VDAC_P.t404 VSS 0.10586f
C10758 VDAC_P.n641 VSS 0.132855f
C10759 VDAC_P.t905 VSS 0.10586f
C10760 VDAC_P.n642 VSS 0.132855f
C10761 VDAC_P.t1260 VSS 0.10586f
C10762 VDAC_P.n643 VSS 0.132855f
C10763 VDAC_P.t1122 VSS 0.10586f
C10764 VDAC_P.n644 VSS 0.132855f
C10765 VDAC_P.t1029 VSS 0.10586f
C10766 VDAC_P.n645 VSS 0.132855f
C10767 VDAC_P.t248 VSS 0.10586f
C10768 VDAC_P.n646 VSS 0.132855f
C10769 VDAC_P.t930 VSS 0.10586f
C10770 VDAC_P.n647 VSS 0.132855f
C10771 VDAC_P.t84 VSS 0.10586f
C10772 VDAC_P.n648 VSS 0.132855f
C10773 VDAC_P.t822 VSS 0.10586f
C10774 VDAC_P.n649 VSS 0.132855f
C10775 VDAC_P.t460 VSS 0.10586f
C10776 VDAC_P.n650 VSS 0.132855f
C10777 VDAC_P.t1182 VSS 0.10586f
C10778 VDAC_P.n651 VSS 0.132855f
C10779 VDAC_P.t1181 VSS 0.10586f
C10780 VDAC_P.n652 VSS 0.132855f
C10781 VDAC_P.t496 VSS 0.10586f
C10782 VDAC_P.n653 VSS 0.132855f
C10783 VDAC_P.t1894 VSS 0.10586f
C10784 VDAC_P.n654 VSS 0.132855f
C10785 VDAC_P.t723 VSS 0.10586f
C10786 VDAC_P.n655 VSS 0.132855f
C10787 VDAC_P.t438 VSS 0.10586f
C10788 VDAC_P.n656 VSS 0.132855f
C10789 VDAC_P.t1319 VSS 0.10586f
C10790 VDAC_P.n657 VSS 0.132855f
C10791 VDAC_P.t66 VSS 0.10586f
C10792 VDAC_P.n658 VSS 0.132855f
C10793 VDAC_P.t1213 VSS 0.10586f
C10794 VDAC_P.n659 VSS 0.132855f
C10795 VDAC_P.t233 VSS 0.10586f
C10796 VDAC_P.n660 VSS 0.132855f
C10797 VDAC_P.t10 VSS 0.10586f
C10798 VDAC_P.n661 VSS 0.132855f
C10799 VDAC_P.t835 VSS 0.10586f
C10800 VDAC_P.n662 VSS 0.132855f
C10801 VDAC_P.t2093 VSS 0.10586f
C10802 VDAC_P.n663 VSS 0.132855f
C10803 VDAC_P.t377 VSS 0.10586f
C10804 VDAC_P.n664 VSS 0.132855f
C10805 VDAC_P.t491 VSS 0.10586f
C10806 VDAC_P.n665 VSS 0.132855f
C10807 VDAC_P.t600 VSS 0.10586f
C10808 VDAC_P.n666 VSS 0.132855f
C10809 VDAC_P.t901 VSS 0.10586f
C10810 VDAC_P.n667 VSS 0.132855f
C10811 VDAC_P.t1164 VSS 0.10586f
C10812 VDAC_P.n668 VSS 0.132855f
C10813 VDAC_P.t131 VSS 0.10586f
C10814 VDAC_P.n669 VSS 0.132855f
C10815 VDAC_P.t553 VSS 0.10586f
C10816 VDAC_P.n670 VSS 0.132855f
C10817 VDAC_P.t464 VSS 0.10586f
C10818 VDAC_P.n671 VSS 0.132855f
C10819 VDAC_P.t277 VSS 0.10586f
C10820 VDAC_P.n672 VSS 0.132855f
C10821 VDAC_P.t1304 VSS 0.10586f
C10822 VDAC_P.n673 VSS 0.132855f
C10823 VDAC_P.t1606 VSS 0.10586f
C10824 VDAC_P.n674 VSS 0.132855f
C10825 VDAC_P.t1676 VSS 0.10586f
C10826 VDAC_P.n675 VSS 0.132855f
C10827 VDAC_P.t1378 VSS 0.10586f
C10828 VDAC_P.n676 VSS 0.132855f
C10829 VDAC_P.t1116 VSS 0.10586f
C10830 VDAC_P.n677 VSS 0.132855f
C10831 VDAC_P.t144 VSS 0.10586f
C10832 VDAC_P.n678 VSS 0.132855f
C10833 VDAC_P.t286 VSS 0.10586f
C10834 VDAC_P.n679 VSS 0.132855f
C10835 VDAC_P.t72 VSS 0.10586f
C10836 VDAC_P.n680 VSS 0.132855f
C10837 VDAC_P.t130 VSS 0.10586f
C10838 VDAC_P.n681 VSS 0.132855f
C10839 VDAC_P.t719 VSS 0.10586f
C10840 VDAC_P.n682 VSS 0.132855f
C10841 VDAC_P.t738 VSS 0.10586f
C10842 VDAC_P.n683 VSS 0.12686f
C10843 VDAC_P.t1516 VSS 0.10586f
C10844 VDAC_P.n684 VSS 0.132855f
C10845 VDAC_P.t1366 VSS 0.10586f
C10846 VDAC_P.n685 VSS 0.132855f
C10847 VDAC_P.t1628 VSS 0.10586f
C10848 VDAC_P.n686 VSS 0.132855f
C10849 VDAC_P.t1856 VSS 0.10586f
C10850 VDAC_P.n687 VSS 0.132855f
C10851 VDAC_P.t258 VSS 0.10586f
C10852 VDAC_P.n688 VSS 0.132855f
C10853 VDAC_P.t1400 VSS 0.10586f
C10854 VDAC_P.n689 VSS 0.132855f
C10855 VDAC_P.t230 VSS 0.10586f
C10856 VDAC_P.n690 VSS 0.132855f
C10857 VDAC_P.t1303 VSS 0.10586f
C10858 VDAC_P.n691 VSS 0.132855f
C10859 VDAC_P.t1434 VSS 0.10586f
C10860 VDAC_P.n692 VSS 0.132855f
C10861 VDAC_P.t101 VSS 0.10586f
C10862 VDAC_P.n693 VSS 0.132855f
C10863 VDAC_P.t88 VSS 0.10586f
C10864 VDAC_P.n694 VSS 0.132855f
C10865 VDAC_P.t555 VSS 0.10586f
C10866 VDAC_P.n695 VSS 0.132855f
C10867 VDAC_P.t1547 VSS 0.10586f
C10868 VDAC_P.n696 VSS 0.132855f
C10869 VDAC_P.t270 VSS 0.10586f
C10870 VDAC_P.n697 VSS 0.132855f
C10871 VDAC_P.t207 VSS 0.10586f
C10872 VDAC_P.n698 VSS 0.132855f
C10873 VDAC_P.t1025 VSS 0.10586f
C10874 VDAC_P.n699 VSS 0.132855f
C10875 VDAC_P.t691 VSS 0.10586f
C10876 VDAC_P.n700 VSS 0.132855f
C10877 VDAC_P.t1805 VSS 0.10586f
C10878 VDAC_P.n701 VSS 0.132855f
C10879 VDAC_P.t884 VSS 0.10586f
C10880 VDAC_P.n702 VSS 0.132855f
C10881 VDAC_P.t865 VSS 0.10586f
C10882 VDAC_P.n703 VSS 0.132855f
C10883 VDAC_P.t156 VSS 0.10586f
C10884 VDAC_P.n704 VSS 0.132855f
C10885 VDAC_P.t811 VSS 0.10586f
C10886 VDAC_P.n705 VSS 0.132855f
C10887 VDAC_P.t533 VSS 0.10586f
C10888 VDAC_P.n706 VSS 0.132855f
C10889 VDAC_P.t736 VSS 0.10586f
C10890 VDAC_P.n707 VSS 0.132855f
C10891 VDAC_P.t931 VSS 0.10586f
C10892 VDAC_P.n708 VSS 0.132855f
C10893 VDAC_P.t1988 VSS 0.10586f
C10894 VDAC_P.n709 VSS 0.132855f
C10895 VDAC_P.t206 VSS 0.10586f
C10896 VDAC_P.n710 VSS 0.132855f
C10897 VDAC_P.t2012 VSS 0.10586f
C10898 VDAC_P.n711 VSS 0.132855f
C10899 VDAC_P.t630 VSS 0.10586f
C10900 VDAC_P.n712 VSS 0.132855f
C10901 VDAC_P.t2079 VSS 0.10586f
C10902 VDAC_P.n713 VSS 0.132855f
C10903 VDAC_P.t1568 VSS 0.10586f
C10904 VDAC_P.n714 VSS 0.132855f
C10905 VDAC_P.t506 VSS 0.10586f
C10906 VDAC_P.n715 VSS 0.132855f
C10907 VDAC_P.t1120 VSS 0.10586f
C10908 VDAC_P.n716 VSS 0.132855f
C10909 VDAC_P.t774 VSS 0.10586f
C10910 VDAC_P.n717 VSS 0.132855f
C10911 VDAC_P.t1239 VSS 0.10586f
C10912 VDAC_P.n718 VSS 0.132855f
C10913 VDAC_P.t658 VSS 0.10586f
C10914 VDAC_P.n719 VSS 0.132855f
C10915 VDAC_P.t303 VSS 0.10586f
C10916 VDAC_P.n720 VSS 0.132855f
C10917 VDAC_P.t448 VSS 0.10586f
C10918 VDAC_P.n721 VSS 0.132855f
C10919 VDAC_P.t1998 VSS 0.10586f
C10920 VDAC_P.n722 VSS 0.132855f
C10921 VDAC_P.t209 VSS 0.10586f
C10922 VDAC_P.n723 VSS 0.132855f
C10923 VDAC_P.t242 VSS 0.10586f
C10924 VDAC_P.n724 VSS 0.132855f
C10925 VDAC_P.t741 VSS 0.10586f
C10926 VDAC_P.n725 VSS 0.132855f
C10927 VDAC_P.t967 VSS 0.10586f
C10928 VDAC_P.n726 VSS 0.132855f
C10929 VDAC_P.t47 VSS 0.10586f
C10930 VDAC_P.n727 VSS 0.132855f
C10931 VDAC_P.t1697 VSS 0.10586f
C10932 VDAC_P.n728 VSS 0.132855f
C10933 VDAC_P.t1548 VSS 0.10586f
C10934 VDAC_P.n729 VSS 0.132855f
C10935 VDAC_P.t807 VSS 0.10586f
C10936 VDAC_P.n730 VSS 0.132855f
C10937 VDAC_P.t91 VSS 0.10586f
C10938 VDAC_P.n731 VSS 0.132855f
C10939 VDAC_P.t119 VSS 0.10586f
C10940 VDAC_P.n732 VSS 0.132855f
C10941 VDAC_P.t1935 VSS 0.10586f
C10942 VDAC_P.n733 VSS 0.132855f
C10943 VDAC_P.t148 VSS 0.10586f
C10944 VDAC_P.n734 VSS 0.132855f
C10945 VDAC_P.t927 VSS 0.10586f
C10946 VDAC_P.n735 VSS 0.132855f
C10947 VDAC_P.t524 VSS 0.10586f
C10948 VDAC_P.n736 VSS 0.132855f
C10949 VDAC_P.t326 VSS 0.10586f
C10950 VDAC_P.n737 VSS 0.132855f
C10951 VDAC_P.t539 VSS 0.10586f
C10952 VDAC_P.n738 VSS 0.132855f
C10953 VDAC_P.t1000 VSS 0.10586f
C10954 VDAC_P.n739 VSS 0.132855f
C10955 VDAC_P.t513 VSS 0.10586f
C10956 VDAC_P.n740 VSS 0.132855f
C10957 VDAC_P.t296 VSS 0.10586f
C10958 VDAC_P.n741 VSS 0.132855f
C10959 VDAC_P.t1710 VSS 0.10586f
C10960 VDAC_P.n742 VSS 0.132855f
C10961 VDAC_P.t68 VSS 0.10586f
C10962 VDAC_P.n743 VSS 0.132855f
C10963 VDAC_P.t1282 VSS 0.10586f
C10964 VDAC_P.n744 VSS 0.132855f
C10965 VDAC_P.t1233 VSS 0.10586f
C10966 VDAC_P.n745 VSS 0.132855f
C10967 VDAC_P.t544 VSS 0.10586f
C10968 VDAC_P.n746 VSS 0.12686f
C10969 VDAC_P.t1124 VSS 0.10586f
C10970 VDAC_P.n747 VSS 0.132855f
C10971 VDAC_P.t1466 VSS 0.10586f
C10972 VDAC_P.n748 VSS 0.132855f
C10973 VDAC_P.t2076 VSS 0.10586f
C10974 VDAC_P.n749 VSS 0.132855f
C10975 VDAC_P.t2016 VSS 0.10586f
C10976 VDAC_P.n750 VSS 0.132855f
C10977 VDAC_P.t1958 VSS 0.10586f
C10978 VDAC_P.n751 VSS 0.132855f
C10979 VDAC_P.t808 VSS 0.10586f
C10980 VDAC_P.n752 VSS 0.132855f
C10981 VDAC_P.t1734 VSS 0.10586f
C10982 VDAC_P.n753 VSS 0.132855f
C10983 VDAC_P.t1347 VSS 0.10586f
C10984 VDAC_P.n754 VSS 0.132855f
C10985 VDAC_P.t778 VSS 0.10586f
C10986 VDAC_P.n755 VSS 0.132855f
C10987 VDAC_P.t1241 VSS 0.10586f
C10988 VDAC_P.n756 VSS 0.132855f
C10989 VDAC_P.t1082 VSS 0.10586f
C10990 VDAC_P.n757 VSS 0.132855f
C10991 VDAC_P.t581 VSS 0.10586f
C10992 VDAC_P.n758 VSS 0.132855f
C10993 VDAC_P.t1583 VSS 0.10586f
C10994 VDAC_P.n759 VSS 0.132855f
C10995 VDAC_P.t1273 VSS 0.10586f
C10996 VDAC_P.n760 VSS 0.132855f
C10997 VDAC_P.t879 VSS 0.10586f
C10998 VDAC_P.n761 VSS 0.132855f
C10999 VDAC_P.t292 VSS 0.10586f
C11000 VDAC_P.n762 VSS 0.132855f
C11001 VDAC_P.t427 VSS 0.10586f
C11002 VDAC_P.n763 VSS 0.132855f
C11003 VDAC_P.t1055 VSS 0.10586f
C11004 VDAC_P.n764 VSS 0.132855f
C11005 VDAC_P.t1016 VSS 0.10586f
C11006 VDAC_P.n765 VSS 0.132855f
C11007 VDAC_P.t1975 VSS 0.10586f
C11008 VDAC_P.n766 VSS 0.132855f
C11009 VDAC_P.t1136 VSS 0.10586f
C11010 VDAC_P.n767 VSS 0.132855f
C11011 VDAC_P.t1859 VSS 0.10586f
C11012 VDAC_P.n768 VSS 0.132855f
C11013 VDAC_P.t692 VSS 0.10586f
C11014 VDAC_P.n769 VSS 0.132855f
C11015 VDAC_P.t1294 VSS 0.10586f
C11016 VDAC_P.n770 VSS 0.132855f
C11017 VDAC_P.t2105 VSS 0.10586f
C11018 VDAC_P.n771 VSS 0.132855f
C11019 VDAC_P.t552 VSS 0.10586f
C11020 VDAC_P.n772 VSS 0.132855f
C11021 VDAC_P.t522 VSS 0.10586f
C11022 VDAC_P.n773 VSS 0.132855f
C11023 VDAC_P.t1232 VSS 0.10586f
C11024 VDAC_P.n774 VSS 0.132855f
C11025 VDAC_P.t466 VSS 0.10586f
C11026 VDAC_P.n775 VSS 0.132855f
C11027 VDAC_P.t804 VSS 0.10586f
C11028 VDAC_P.n776 VSS 0.132855f
C11029 VDAC_P.t358 VSS 0.10586f
C11030 VDAC_P.n777 VSS 0.132855f
C11031 VDAC_P.t1263 VSS 0.10586f
C11032 VDAC_P.n778 VSS 0.132855f
C11033 VDAC_P.t1134 VSS 0.10586f
C11034 VDAC_P.n779 VSS 0.132855f
C11035 VDAC_P.t1042 VSS 0.10586f
C11036 VDAC_P.n780 VSS 0.132855f
C11037 VDAC_P.t769 VSS 0.10586f
C11038 VDAC_P.n781 VSS 0.132855f
C11039 VDAC_P.t1846 VSS 0.10586f
C11040 VDAC_P.n782 VSS 0.132855f
C11041 VDAC_P.t1393 VSS 0.10586f
C11042 VDAC_P.n783 VSS 0.132855f
C11043 VDAC_P.t1406 VSS 0.10586f
C11044 VDAC_P.n784 VSS 0.132855f
C11045 VDAC_P.t659 VSS 0.10586f
C11046 VDAC_P.n785 VSS 0.132855f
C11047 VDAC_P.t887 VSS 0.10586f
C11048 VDAC_P.n786 VSS 0.132855f
C11049 VDAC_P.t1169 VSS 0.10586f
C11050 VDAC_P.n787 VSS 0.132855f
C11051 VDAC_P.t1723 VSS 0.10586f
C11052 VDAC_P.n788 VSS 0.132855f
C11053 VDAC_P.t988 VSS 0.10586f
C11054 VDAC_P.n789 VSS 0.132855f
C11055 VDAC_P.t121 VSS 0.10586f
C11056 VDAC_P.n790 VSS 0.132855f
C11057 VDAC_P.t1971 VSS 0.10586f
C11058 VDAC_P.n791 VSS 0.132855f
C11059 VDAC_P.t408 VSS 0.10586f
C11060 VDAC_P.n792 VSS 0.132855f
C11061 VDAC_P.t1857 VSS 0.10586f
C11062 VDAC_P.n793 VSS 0.132855f
C11063 VDAC_P.t676 VSS 0.10586f
C11064 VDAC_P.n794 VSS 0.132855f
C11065 VDAC_P.t459 VSS 0.10586f
C11066 VDAC_P.n795 VSS 0.132855f
C11067 VDAC_P.t1724 VSS 0.10586f
C11068 VDAC_P.n796 VSS 0.132855f
C11069 VDAC_P.t2104 VSS 0.10586f
C11070 VDAC_P.n797 VSS 0.132855f
C11071 VDAC_P.t287 VSS 0.10586f
C11072 VDAC_P.n798 VSS 0.132855f
C11073 VDAC_P.t80 VSS 0.10586f
C11074 VDAC_P.n799 VSS 0.132855f
C11075 VDAC_P.t246 VSS 0.10586f
C11076 VDAC_P.n800 VSS 0.132855f
C11077 VDAC_P.t1556 VSS 0.10586f
C11078 VDAC_P.n801 VSS 0.132855f
C11079 VDAC_P.t34 VSS 0.10586f
C11080 VDAC_P.n802 VSS 0.132855f
C11081 VDAC_P.t1324 VSS 0.10586f
C11082 VDAC_P.n803 VSS 0.132855f
C11083 VDAC_P.t578 VSS 0.10586f
C11084 VDAC_P.n804 VSS 0.132855f
C11085 VDAC_P.t1155 VSS 0.10586f
C11086 VDAC_P.n805 VSS 0.132855f
C11087 VDAC_P.t472 VSS 0.10586f
C11088 VDAC_P.n806 VSS 0.132855f
C11089 VDAC_P.t1838 VSS 0.10586f
C11090 VDAC_P.n807 VSS 0.132855f
C11091 VDAC_P.t1503 VSS 0.10586f
C11092 VDAC_P.n808 VSS 0.132855f
C11093 VDAC_P.t826 VSS 0.10586f
C11094 VDAC_P.n809 VSS 0.12686f
C11095 VDAC_P.t1874 VSS 0.10586f
C11096 VDAC_P.n810 VSS 0.132855f
C11097 VDAC_P.t1521 VSS 0.10586f
C11098 VDAC_P.n811 VSS 0.132855f
C11099 VDAC_P.t838 VSS 0.10586f
C11100 VDAC_P.n812 VSS 0.132855f
C11101 VDAC_P.t1307 VSS 0.10586f
C11102 VDAC_P.n813 VSS 0.132855f
C11103 VDAC_P.t461 VSS 0.10586f
C11104 VDAC_P.n814 VSS 0.132855f
C11105 VDAC_P.t1199 VSS 0.10586f
C11106 VDAC_P.n815 VSS 0.132855f
C11107 VDAC_P.t435 VSS 0.10586f
C11108 VDAC_P.n816 VSS 0.132855f
C11109 VDAC_P.t93 VSS 0.10586f
C11110 VDAC_P.n817 VSS 0.132855f
C11111 VDAC_P.t1551 VSS 0.10586f
C11112 VDAC_P.n818 VSS 0.132855f
C11113 VDAC_P.t1017 VSS 0.10586f
C11114 VDAC_P.n819 VSS 0.132855f
C11115 VDAC_P.t683 VSS 0.10586f
C11116 VDAC_P.n820 VSS 0.132855f
C11117 VDAC_P.t1893 VSS 0.10586f
C11118 VDAC_P.n821 VSS 0.132855f
C11119 VDAC_P.t1604 VSS 0.10586f
C11120 VDAC_P.n822 VSS 0.132855f
C11121 VDAC_P.t1467 VSS 0.10586f
C11122 VDAC_P.n823 VSS 0.132855f
C11123 VDAC_P.t973 VSS 0.10586f
C11124 VDAC_P.n824 VSS 0.132855f
C11125 VDAC_P.t192 VSS 0.10586f
C11126 VDAC_P.n825 VSS 0.132855f
C11127 VDAC_P.t1813 VSS 0.10586f
C11128 VDAC_P.n826 VSS 0.132855f
C11129 VDAC_P.t1804 VSS 0.10586f
C11130 VDAC_P.n827 VSS 0.132855f
C11131 VDAC_P.t370 VSS 0.10586f
C11132 VDAC_P.n828 VSS 0.132855f
C11133 VDAC_P.t284 VSS 0.10586f
C11134 VDAC_P.n829 VSS 0.132855f
C11135 VDAC_P.t1912 VSS 0.10586f
C11136 VDAC_P.n830 VSS 0.132855f
C11137 VDAC_P.t2053 VSS 0.10586f
C11138 VDAC_P.n831 VSS 0.132855f
C11139 VDAC_P.t1472 VSS 0.10586f
C11140 VDAC_P.n832 VSS 0.132855f
C11141 VDAC_P.t1674 VSS 0.10586f
C11142 VDAC_P.n833 VSS 0.132855f
C11143 VDAC_P.t1140 VSS 0.10586f
C11144 VDAC_P.n834 VSS 0.132855f
C11145 VDAC_P.t750 VSS 0.10586f
C11146 VDAC_P.n835 VSS 0.132855f
C11147 VDAC_P.t325 VSS 0.10586f
C11148 VDAC_P.n836 VSS 0.132855f
C11149 VDAC_P.t528 VSS 0.10586f
C11150 VDAC_P.n837 VSS 0.132855f
C11151 VDAC_P.t563 VSS 0.10586f
C11152 VDAC_P.n838 VSS 0.132855f
C11153 VDAC_P.t1600 VSS 0.10586f
C11154 VDAC_P.n839 VSS 0.132855f
C11155 VDAC_P.t1738 VSS 0.10586f
C11156 VDAC_P.n840 VSS 0.132855f
C11157 VDAC_P.t1453 VSS 0.10586f
C11158 VDAC_P.n841 VSS 0.132855f
C11159 VDAC_P.t122 VSS 0.10586f
C11160 VDAC_P.n842 VSS 0.132855f
C11161 VDAC_P.t1243 VSS 0.10586f
C11162 VDAC_P.n843 VSS 0.132855f
C11163 VDAC_P.t445 VSS 0.10586f
C11164 VDAC_P.n844 VSS 0.132855f
C11165 VDAC_P.t1137 VSS 0.10586f
C11166 VDAC_P.n845 VSS 0.132855f
C11167 VDAC_P.t1585 VSS 0.10586f
C11168 VDAC_P.n846 VSS 0.132855f
C11169 VDAC_P.t910 VSS 0.10586f
C11170 VDAC_P.n847 VSS 0.132855f
C11171 VDAC_P.t1483 VSS 0.10586f
C11172 VDAC_P.n848 VSS 0.132855f
C11173 VDAC_P.t981 VSS 0.10586f
C11174 VDAC_P.n849 VSS 0.132855f
C11175 VDAC_P.t1359 VSS 0.10586f
C11176 VDAC_P.n850 VSS 0.132855f
C11177 VDAC_P.t971 VSS 0.10586f
C11178 VDAC_P.n851 VSS 0.132855f
C11179 VDAC_P.t468 VSS 0.10586f
C11180 VDAC_P.n852 VSS 0.132855f
C11181 VDAC_P.t867 VSS 0.10586f
C11182 VDAC_P.n853 VSS 0.132855f
C11183 VDAC_P.t1692 VSS 0.10586f
C11184 VDAC_P.n854 VSS 0.132855f
C11185 VDAC_P.t314 VSS 0.10586f
C11186 VDAC_P.n855 VSS 0.132855f
C11187 VDAC_P.t1039 VSS 0.10586f
C11188 VDAC_P.n856 VSS 0.132855f
C11189 VDAC_P.t384 VSS 0.10586f
C11190 VDAC_P.n857 VSS 0.132855f
C11191 VDAC_P.t507 VSS 0.10586f
C11192 VDAC_P.n858 VSS 0.132855f
C11193 VDAC_P.t2004 VSS 0.10586f
C11194 VDAC_P.n859 VSS 0.132855f
C11195 VDAC_P.t1458 VSS 0.10586f
C11196 VDAC_P.n860 VSS 0.132855f
C11197 VDAC_P.t2124 VSS 0.10586f
C11198 VDAC_P.n861 VSS 0.132855f
C11199 VDAC_P.t1238 VSS 0.10586f
C11200 VDAC_P.n862 VSS 0.132855f
C11201 VDAC_P.t1093 VSS 0.10586f
C11202 VDAC_P.n863 VSS 0.132855f
C11203 VDAC_P.t416 VSS 0.10586f
C11204 VDAC_P.n864 VSS 0.132855f
C11205 VDAC_P.t1946 VSS 0.10586f
C11206 VDAC_P.n865 VSS 0.132855f
C11207 VDAC_P.t304 VSS 0.10586f
C11208 VDAC_P.n866 VSS 0.132855f
C11209 VDAC_P.t402 VSS 0.10586f
C11210 VDAC_P.n867 VSS 0.132855f
C11211 VDAC_P.t685 VSS 0.10586f
C11212 VDAC_P.n868 VSS 0.132855f
C11213 VDAC_P.t186 VSS 0.10586f
C11214 VDAC_P.n869 VSS 0.132855f
C11215 VDAC_P.t1131 VSS 0.10586f
C11216 VDAC_P.n870 VSS 0.132855f
C11217 VDAC_P.t1693 VSS 0.10586f
C11218 VDAC_P.n871 VSS 0.132855f
C11219 VDAC_P.t2002 VSS 0.10586f
C11220 VDAC_P.n872 VSS 0.12686f
C11221 VDAC_P.t451 VSS 0.10586f
C11222 VDAC_P.n873 VSS 0.132855f
C11223 VDAC_P.t1964 VSS 0.10586f
C11224 VDAC_P.n874 VSS 0.132855f
C11225 VDAC_P.t823 VSS 0.10586f
C11226 VDAC_P.n875 VSS 0.132855f
C11227 VDAC_P.t2067 VSS 0.10586f
C11228 VDAC_P.n876 VSS 0.132855f
C11229 VDAC_P.t1536 VSS 0.10586f
C11230 VDAC_P.n877 VSS 0.132855f
C11231 VDAC_P.t1963 VSS 0.10586f
C11232 VDAC_P.n878 VSS 0.132855f
C11233 VDAC_P.t2132 VSS 0.10586f
C11234 VDAC_P.n879 VSS 0.132855f
C11235 VDAC_P.t1502 VSS 0.10586f
C11236 VDAC_P.n880 VSS 0.132855f
C11237 VDAC_P.t644 VSS 0.10586f
C11238 VDAC_P.n881 VSS 0.132855f
C11239 VDAC_P.t650 VSS 0.10586f
C11240 VDAC_P.n882 VSS 0.132855f
C11241 VDAC_P.t2097 VSS 0.10586f
C11242 VDAC_P.n883 VSS 0.132855f
C11243 VDAC_P.t32 VSS 0.10586f
C11244 VDAC_P.n884 VSS 0.132855f
C11245 VDAC_P.t1982 VSS 0.10586f
C11246 VDAC_P.n885 VSS 0.132855f
C11247 VDAC_P.t1653 VSS 0.10586f
C11248 VDAC_P.n886 VSS 0.132855f
C11249 VDAC_P.t547 VSS 0.10586f
C11250 VDAC_P.n887 VSS 0.132855f
C11251 VDAC_P.t2120 VSS 0.10586f
C11252 VDAC_P.n888 VSS 0.132855f
C11253 VDAC_P.t2003 VSS 0.10586f
C11254 VDAC_P.n889 VSS 0.132855f
C11255 VDAC_P.t328 VSS 0.10586f
C11256 VDAC_P.n890 VSS 0.132855f
C11257 VDAC_P.t1778 VSS 0.10586f
C11258 VDAC_P.n891 VSS 0.132855f
C11259 VDAC_P.t1572 VSS 0.10586f
C11260 VDAC_P.n892 VSS 0.132855f
C11261 VDAC_P.t1346 VSS 0.10586f
C11262 VDAC_P.n893 VSS 0.132855f
C11263 VDAC_P.t1356 VSS 0.10586f
C11264 VDAC_P.n894 VSS 0.132855f
C11265 VDAC_P.t1130 VSS 0.10586f
C11266 VDAC_P.n895 VSS 0.132855f
C11267 VDAC_P.t2054 VSS 0.10586f
C11268 VDAC_P.n896 VSS 0.132855f
C11269 VDAC_P.t360 VSS 0.10586f
C11270 VDAC_P.n897 VSS 0.132855f
C11271 VDAC_P.t482 VSS 0.10586f
C11272 VDAC_P.n898 VSS 0.132855f
C11273 VDAC_P.t1391 VSS 0.10586f
C11274 VDAC_P.n899 VSS 0.132855f
C11275 VDAC_P.t1402 VSS 0.10586f
C11276 VDAC_P.n900 VSS 0.132855f
C11277 VDAC_P.t1289 VSS 0.10586f
C11278 VDAC_P.n901 VSS 0.132855f
C11279 VDAC_P.t610 VSS 0.10586f
C11280 VDAC_P.n902 VSS 0.132855f
C11281 VDAC_P.t1070 VSS 0.10586f
C11282 VDAC_P.n903 VSS 0.132855f
C11283 VDAC_P.t1641 VSS 0.10586f
C11284 VDAC_P.n904 VSS 0.132855f
C11285 VDAC_P.t498 VSS 0.10586f
C11286 VDAC_P.n905 VSS 0.132855f
C11287 VDAC_P.t1423 VSS 0.10586f
C11288 VDAC_P.n906 VSS 0.132855f
C11289 VDAC_P.t1879 VSS 0.10586f
C11290 VDAC_P.n907 VSS 0.132855f
C11291 VDAC_P.t677 VSS 0.10586f
C11292 VDAC_P.n908 VSS 0.132855f
C11293 VDAC_P.t1773 VSS 0.10586f
C11294 VDAC_P.n909 VSS 0.132855f
C11295 VDAC_P.t1107 VSS 0.10586f
C11296 VDAC_P.n910 VSS 0.132855f
C11297 VDAC_P.t1675 VSS 0.10586f
C11298 VDAC_P.n911 VSS 0.132855f
C11299 VDAC_P.t2127 VSS 0.10586f
C11300 VDAC_P.n912 VSS 0.132855f
C11301 VDAC_P.t407 VSS 0.10586f
C11302 VDAC_P.n913 VSS 0.132855f
C11303 VDAC_P.t2099 VSS 0.10586f
C11304 VDAC_P.n914 VSS 0.132855f
C11305 VDAC_P.t1688 VSS 0.10586f
C11306 VDAC_P.n915 VSS 0.132855f
C11307 VDAC_P.t1891 VSS 0.10586f
C11308 VDAC_P.n916 VSS 0.132855f
C11309 VDAC_P.t788 VSS 0.10586f
C11310 VDAC_P.n917 VSS 0.132855f
C11311 VDAC_P.t1562 VSS 0.10586f
C11312 VDAC_P.n918 VSS 0.132855f
C11313 VDAC_P.t108 VSS 0.10586f
C11314 VDAC_P.n919 VSS 0.132855f
C11315 VDAC_P.t1126 VSS 0.10586f
C11316 VDAC_P.n920 VSS 0.132855f
C11317 VDAC_P.t65 VSS 0.10586f
C11318 VDAC_P.n921 VSS 0.132855f
C11319 VDAC_P.t912 VSS 0.10586f
C11320 VDAC_P.n922 VSS 0.132855f
C11321 VDAC_P.t254 VSS 0.10586f
C11322 VDAC_P.n923 VSS 0.132855f
C11323 VDAC_P.t680 VSS 0.10586f
C11324 VDAC_P.n924 VSS 0.132855f
C11325 VDAC_P.t426 VSS 0.10586f
C11326 VDAC_P.n925 VSS 0.132855f
C11327 VDAC_P.t1285 VSS 0.10586f
C11328 VDAC_P.n926 VSS 0.132855f
C11329 VDAC_P.t606 VSS 0.10586f
C11330 VDAC_P.n927 VSS 0.132855f
C11331 VDAC_P.t1183 VSS 0.10586f
C11332 VDAC_P.n928 VSS 0.132855f
C11333 VDAC_P.t968 VSS 0.10586f
C11334 VDAC_P.n929 VSS 0.132855f
C11335 VDAC_P.t1898 VSS 0.10586f
C11336 VDAC_P.n930 VSS 0.132855f
C11337 VDAC_P.t403 VSS 0.10586f
C11338 VDAC_P.n931 VSS 0.132855f
C11339 VDAC_P.t850 VSS 0.10586f
C11340 VDAC_P.n932 VSS 0.132855f
C11341 VDAC_P.t351 VSS 0.10586f
C11342 VDAC_P.n933 VSS 0.132855f
C11343 VDAC_P.t1871 VSS 0.10586f
C11344 VDAC_P.n934 VSS 0.132855f
C11345 VDAC_P.t1215 VSS 0.10586f
C11346 VDAC_P.n935 VSS 0.12686f
C11347 VDAC_P.t1526 VSS 0.10586f
C11348 VDAC_P.n936 VSS 0.132855f
C11349 VDAC_P.t357 VSS 0.10586f
C11350 VDAC_P.n937 VSS 0.132855f
C11351 VDAC_P.t1298 VSS 0.10586f
C11352 VDAC_P.n938 VSS 0.132855f
C11353 VDAC_P.t1133 VSS 0.10586f
C11354 VDAC_P.n939 VSS 0.132855f
C11355 VDAC_P.t805 VSS 0.10586f
C11356 VDAC_P.n940 VSS 0.132855f
C11357 VDAC_P.t1018 VSS 0.10586f
C11358 VDAC_P.n941 VSS 0.132855f
C11359 VDAC_P.t391 VSS 0.10586f
C11360 VDAC_P.n942 VSS 0.132855f
C11361 VDAC_P.t1931 VSS 0.10586f
C11362 VDAC_P.n943 VSS 0.132855f
C11363 VDAC_P.t1371 VSS 0.10586f
C11364 VDAC_P.n944 VSS 0.132855f
C11365 VDAC_P.t477 VSS 0.10586f
C11366 VDAC_P.n945 VSS 0.132855f
C11367 VDAC_P.t1163 VSS 0.10586f
C11368 VDAC_P.n946 VSS 0.132855f
C11369 VDAC_P.t1717 VSS 0.10586f
C11370 VDAC_P.n947 VSS 0.132855f
C11371 VDAC_P.t2126 VSS 0.10586f
C11372 VDAC_P.n948 VSS 0.132855f
C11373 VDAC_P.t1425 VSS 0.10586f
C11374 VDAC_P.n949 VSS 0.132855f
C11375 VDAC_P.t955 VSS 0.10586f
C11376 VDAC_P.n950 VSS 0.132855f
C11377 VDAC_P.t1176 VSS 0.10586f
C11378 VDAC_P.n951 VSS 0.132855f
C11379 VDAC_P.t1775 VSS 0.10586f
C11380 VDAC_P.n952 VSS 0.132855f
C11381 VDAC_P.t1196 VSS 0.10586f
C11382 VDAC_P.n953 VSS 0.132855f
C11383 VDAC_P.t190 VSS 0.10586f
C11384 VDAC_P.n954 VSS 0.132855f
C11385 VDAC_P.t2129 VSS 0.10586f
C11386 VDAC_P.n955 VSS 0.132855f
C11387 VDAC_P.t904 VSS 0.10586f
C11388 VDAC_P.n956 VSS 0.132855f
C11389 VDAC_P.t2021 VSS 0.10586f
C11390 VDAC_P.n957 VSS 0.132855f
C11391 VDAC_P.t48 VSS 0.10586f
C11392 VDAC_P.n958 VSS 0.132855f
C11393 VDAC_P.t818 VSS 0.10586f
C11394 VDAC_P.n959 VSS 0.132855f
C11395 VDAC_P.t236 VSS 0.10586f
C11396 VDAC_P.n960 VSS 0.132855f
C11397 VDAC_P.t366 VSS 0.10586f
C11398 VDAC_P.n961 VSS 0.132855f
C11399 VDAC_P.t603 VSS 0.10586f
C11400 VDAC_P.n962 VSS 0.132855f
C11401 VDAC_P.t1888 VSS 0.10586f
C11402 VDAC_P.n963 VSS 0.132855f
C11403 VDAC_P.t2094 VSS 0.10586f
C11404 VDAC_P.n964 VSS 0.132855f
C11405 VDAC_P.t1440 VSS 0.10586f
C11406 VDAC_P.n965 VSS 0.132855f
C11407 VDAC_P.t1662 VSS 0.10586f
C11408 VDAC_P.n966 VSS 0.132855f
C11409 VDAC_P.t1411 VSS 0.10586f
C11410 VDAC_P.n967 VSS 0.132855f
C11411 VDAC_P.t1450 VSS 0.10586f
C11412 VDAC_P.n968 VSS 0.132855f
C11413 VDAC_P.t323 VSS 0.10586f
C11414 VDAC_P.n969 VSS 0.132855f
C11415 VDAC_P.t1663 VSS 0.10586f
C11416 VDAC_P.n970 VSS 0.132855f
C11417 VDAC_P.t161 VSS 0.10586f
C11418 VDAC_P.n971 VSS 0.132855f
C11419 VDAC_P.t1559 VSS 0.10586f
C11420 VDAC_P.n972 VSS 0.132855f
C11421 VDAC_P.t878 VSS 0.10586f
C11422 VDAC_P.n973 VSS 0.132855f
C11423 VDAC_P.t1447 VSS 0.10586f
C11424 VDAC_P.n974 VSS 0.132855f
C11425 VDAC_P.t1901 VSS 0.10586f
C11426 VDAC_P.n975 VSS 0.132855f
C11427 VDAC_P.t1321 VSS 0.10586f
C11428 VDAC_P.n976 VSS 0.132855f
C11429 VDAC_P.t489 VSS 0.10586f
C11430 VDAC_P.n977 VSS 0.132855f
C11431 VDAC_P.t1444 VSS 0.10586f
C11432 VDAC_P.n978 VSS 0.132855f
C11433 VDAC_P.t849 VSS 0.10586f
C11434 VDAC_P.n979 VSS 0.132855f
C11435 VDAC_P.t2121 VSS 0.10586f
C11436 VDAC_P.n980 VSS 0.132855f
C11437 VDAC_P.t1098 VSS 0.10586f
C11438 VDAC_P.n981 VSS 0.132855f
C11439 VDAC_P.t2015 VSS 0.10586f
C11440 VDAC_P.n982 VSS 0.132855f
C11441 VDAC_P.t1296 VSS 0.10586f
C11442 VDAC_P.n983 VSS 0.132855f
C11443 VDAC_P.t1905 VSS 0.10586f
C11444 VDAC_P.n984 VSS 0.132855f
C11445 VDAC_P.t1700 VSS 0.10586f
C11446 VDAC_P.n985 VSS 0.132855f
C11447 VDAC_P.t70 VSS 0.10586f
C11448 VDAC_P.n986 VSS 0.132855f
C11449 VDAC_P.t780 VSS 0.10586f
C11450 VDAC_P.n987 VSS 0.132855f
C11451 VDAC_P.t594 VSS 0.10586f
C11452 VDAC_P.n988 VSS 0.132855f
C11453 VDAC_P.t1054 VSS 0.10586f
C11454 VDAC_P.n989 VSS 0.132855f
C11455 VDAC_P.t720 VSS 0.10586f
C11456 VDAC_P.n990 VSS 0.132855f
C11457 VDAC_P.t950 VSS 0.10586f
C11458 VDAC_P.n991 VSS 0.132855f
C11459 VDAC_P.t1940 VSS 0.10586f
C11460 VDAC_P.n992 VSS 0.132855f
C11461 VDAC_P.t734 VSS 0.10586f
C11462 VDAC_P.n993 VSS 0.132855f
C11463 VDAC_P.t667 VSS 0.10586f
C11464 VDAC_P.n994 VSS 0.132855f
C11465 VDAC_P.t1218 VSS 0.10586f
C11466 VDAC_P.n995 VSS 0.132855f
C11467 VDAC_P.t293 VSS 0.10586f
C11468 VDAC_P.n996 VSS 0.132855f
C11469 VDAC_P.t1655 VSS 0.10586f
C11470 VDAC_P.n997 VSS 0.132855f
C11471 VDAC_P.t266 VSS 0.10586f
C11472 VDAC_P.n998 VSS 0.12686f
C11473 VDAC_P.t789 VSS 0.10586f
C11474 VDAC_P.n999 VSS 0.132855f
C11475 VDAC_P.t1067 VSS 0.10586f
C11476 VDAC_P.n1000 VSS 0.132855f
C11477 VDAC_P.t733 VSS 0.10586f
C11478 VDAC_P.n1001 VSS 0.132855f
C11479 VDAC_P.t261 VSS 0.10586f
C11480 VDAC_P.n1002 VSS 0.132855f
C11481 VDAC_P.t420 VSS 0.10586f
C11482 VDAC_P.n1003 VSS 0.132855f
C11483 VDAC_P.t1791 VSS 0.10586f
C11484 VDAC_P.n1004 VSS 0.132855f
C11485 VDAC_P.t1388 VSS 0.10586f
C11486 VDAC_P.n1005 VSS 0.132855f
C11487 VDAC_P.t1138 VSS 0.10586f
C11488 VDAC_P.n1006 VSS 0.132855f
C11489 VDAC_P.t388 VSS 0.10586f
C11490 VDAC_P.n1007 VSS 0.132855f
C11491 VDAC_P.t1816 VSS 0.10586f
C11492 VDAC_P.n1008 VSS 0.132855f
C11493 VDAC_P.t1923 VSS 0.10586f
C11494 VDAC_P.n1009 VSS 0.132855f
C11495 VDAC_P.t1360 VSS 0.10586f
C11496 VDAC_P.n1010 VSS 0.132855f
C11497 VDAC_P.t1626 VSS 0.10586f
C11498 VDAC_P.n1011 VSS 0.132855f
C11499 VDAC_P.t1619 VSS 0.10586f
C11500 VDAC_P.n1012 VSS 0.132855f
C11501 VDAC_P.t2071 VSS 0.10586f
C11502 VDAC_P.n1013 VSS 0.132855f
C11503 VDAC_P.t512 VSS 0.10586f
C11504 VDAC_P.n1014 VSS 0.132855f
C11505 VDAC_P.t997 VSS 0.10586f
C11506 VDAC_P.n1015 VSS 0.132855f
C11507 VDAC_P.t1096 VSS 0.10586f
C11508 VDAC_P.n1016 VSS 0.132855f
C11509 VDAC_P.t238 VSS 0.10586f
C11510 VDAC_P.n1017 VSS 0.132855f
C11511 VDAC_P.t660 VSS 0.10586f
C11512 VDAC_P.n1018 VSS 0.132855f
C11513 VDAC_P.t654 VSS 0.10586f
C11514 VDAC_P.n1019 VSS 0.132855f
C11515 VDAC_P.t124 VSS 0.10586f
C11516 VDAC_P.n1020 VSS 0.132855f
C11517 VDAC_P.t2088 VSS 0.10586f
C11518 VDAC_P.n1021 VSS 0.132855f
C11519 VDAC_P.t518 VSS 0.10586f
C11520 VDAC_P.n1022 VSS 0.132855f
C11521 VDAC_P.t1216 VSS 0.10586f
C11522 VDAC_P.n1023 VSS 0.132855f
C11523 VDAC_P.t898 VSS 0.10586f
C11524 VDAC_P.n1024 VSS 0.132855f
C11525 VDAC_P.t697 VSS 0.10586f
C11526 VDAC_P.n1025 VSS 0.132855f
C11527 VDAC_P.t110 VSS 0.10586f
C11528 VDAC_P.n1026 VSS 0.132855f
C11529 VDAC_P.t1259 VSS 0.10586f
C11530 VDAC_P.n1027 VSS 0.132855f
C11531 VDAC_P.t574 VSS 0.10586f
C11532 VDAC_P.n1028 VSS 0.132855f
C11533 VDAC_P.t2046 VSS 0.10586f
C11534 VDAC_P.n1029 VSS 0.132855f
C11535 VDAC_P.t423 VSS 0.10586f
C11536 VDAC_P.n1030 VSS 0.132855f
C11537 VDAC_P.t1830 VSS 0.10586f
C11538 VDAC_P.n1031 VSS 0.132855f
C11539 VDAC_P.t113 VSS 0.10586f
C11540 VDAC_P.n1032 VSS 0.132855f
C11541 VDAC_P.t937 VSS 0.10586f
C11542 VDAC_P.n1033 VSS 0.132855f
C11543 VDAC_P.t185 VSS 0.10586f
C11544 VDAC_P.n1034 VSS 0.132855f
C11545 VDAC_P.t1741 VSS 0.10586f
C11546 VDAC_P.n1035 VSS 0.132855f
C11547 VDAC_P.t8 VSS 0.10586f
C11548 VDAC_P.n1036 VSS 0.132855f
C11549 VDAC_P.t833 VSS 0.10586f
C11550 VDAC_P.n1037 VSS 0.132855f
C11551 VDAC_P.t2089 VSS 0.10586f
C11552 VDAC_P.n1038 VSS 0.132855f
C11553 VDAC_P.t1509 VSS 0.10586f
C11554 VDAC_P.n1039 VSS 0.132855f
C11555 VDAC_P.t2063 VSS 0.10586f
C11556 VDAC_P.n1040 VSS 0.132855f
C11557 VDAC_P.t1520 VSS 0.10586f
C11558 VDAC_P.n1041 VSS 0.132855f
C11559 VDAC_P.t85 VSS 0.10586f
C11560 VDAC_P.n1042 VSS 0.132855f
C11561 VDAC_P.t180 VSS 0.10586f
C11562 VDAC_P.n1043 VSS 0.132855f
C11563 VDAC_P.t1494 VSS 0.10586f
C11564 VDAC_P.n1044 VSS 0.132855f
C11565 VDAC_P.t380 VSS 0.10586f
C11566 VDAC_P.n1045 VSS 0.132855f
C11567 VDAC_P.t2072 VSS 0.10586f
C11568 VDAC_P.n1046 VSS 0.132855f
C11569 VDAC_P.t157 VSS 0.10586f
C11570 VDAC_P.n1047 VSS 0.132855f
C11571 VDAC_P.t232 VSS 0.10586f
C11572 VDAC_P.n1048 VSS 0.132855f
C11573 VDAC_P.t894 VSS 0.10586f
C11574 VDAC_P.n1049 VSS 0.132855f
C11575 VDAC_P.t1168 VSS 0.10586f
C11576 VDAC_P.n1050 VSS 0.132855f
C11577 VDAC_P.t410 VSS 0.10586f
C11578 VDAC_P.n1051 VSS 0.132855f
C11579 VDAC_P.t1253 VSS 0.10586f
C11580 VDAC_P.n1052 VSS 0.132855f
C11581 VDAC_P.t298 VSS 0.10586f
C11582 VDAC_P.n1053 VSS 0.132855f
C11583 VDAC_P.t1151 VSS 0.10586f
C11584 VDAC_P.n1054 VSS 0.132855f
C11585 VDAC_P.t1768 VSS 0.10586f
C11586 VDAC_P.n1055 VSS 0.132855f
C11587 VDAC_P.t42 VSS 0.10586f
C11588 VDAC_P.n1056 VSS 0.132855f
C11589 VDAC_P.t763 VSS 0.10586f
C11590 VDAC_P.n1057 VSS 0.132855f
C11591 VDAC_P.t422 VSS 0.10586f
C11592 VDAC_P.n1058 VSS 0.132855f
C11593 VDAC_P.t341 VSS 0.10586f
C11594 VDAC_P.n1059 VSS 0.132855f
C11595 VDAC_P.t935 VSS 0.10586f
C11596 VDAC_P.n1060 VSS 0.132855f
C11597 VDAC_P.t1177 VSS 0.10586f
C11598 VDAC_P.n1061 VSS 0.12686f
C11599 VDAC_P.t840 VSS 0.10586f
C11600 VDAC_P.n1062 VSS 0.132855f
C11601 VDAC_P.t514 VSS 0.10586f
C11602 VDAC_P.n1063 VSS 0.132855f
C11603 VDAC_P.t312 VSS 0.10586f
C11604 VDAC_P.n1064 VSS 0.132855f
C11605 VDAC_P.t1554 VSS 0.10586f
C11606 VDAC_P.n1065 VSS 0.132855f
C11607 VDAC_P.t181 VSS 0.10586f
C11608 VDAC_P.n1066 VSS 0.132855f
C11609 VDAC_P.t1322 VSS 0.10586f
C11610 VDAC_P.n1067 VSS 0.132855f
C11611 VDAC_P.t589 VSS 0.10586f
C11612 VDAC_P.n1068 VSS 0.132855f
C11613 VDAC_P.t1603 VSS 0.10586f
C11614 VDAC_P.n1069 VSS 0.132855f
C11615 VDAC_P.t530 VSS 0.10586f
C11616 VDAC_P.n1070 VSS 0.132855f
C11617 VDAC_P.t1497 VSS 0.10586f
C11618 VDAC_P.n1071 VSS 0.132855f
C11619 VDAC_P.t1598 VSS 0.10586f
C11620 VDAC_P.n1072 VSS 0.132855f
C11621 VDAC_P.t1383 VSS 0.10586f
C11622 VDAC_P.n1073 VSS 0.132855f
C11623 VDAC_P.t481 VSS 0.10586f
C11624 VDAC_P.n1074 VSS 0.132855f
C11625 VDAC_P.t1762 VSS 0.10586f
C11626 VDAC_P.n1075 VSS 0.132855f
C11627 VDAC_P.t1361 VSS 0.10586f
C11628 VDAC_P.n1076 VSS 0.132855f
C11629 VDAC_P.t501 VSS 0.10586f
C11630 VDAC_P.n1077 VSS 0.132855f
C11631 VDAC_P.t641 VSS 0.10586f
C11632 VDAC_P.n1078 VSS 0.132855f
C11633 VDAC_P.t133 VSS 0.10586f
C11634 VDAC_P.n1079 VSS 0.132855f
C11635 VDAC_P.t1836 VSS 0.10586f
C11636 VDAC_P.n1080 VSS 0.132855f
C11637 VDAC_P.t1605 VSS 0.10586f
C11638 VDAC_P.n1081 VSS 0.132855f
C11639 VDAC_P.t1043 VSS 0.10586f
C11640 VDAC_P.n1082 VSS 0.132855f
C11641 VDAC_P.t1499 VSS 0.10586f
C11642 VDAC_P.n1083 VSS 0.132855f
C11643 VDAC_P.t1951 VSS 0.10586f
C11644 VDAC_P.n1084 VSS 0.132855f
C11645 VDAC_P.t2068 VSS 0.10586f
C11646 VDAC_P.n1085 VSS 0.132855f
C11647 VDAC_P.t883 VSS 0.10586f
C11648 VDAC_P.n1086 VSS 0.132855f
C11649 VDAC_P.t1172 VSS 0.10586f
C11650 VDAC_P.n1087 VSS 0.132855f
C11651 VDAC_P.t334 VSS 0.10586f
C11652 VDAC_P.n1088 VSS 0.132855f
C11653 VDAC_P.t1057 VSS 0.10586f
C11654 VDAC_P.n1089 VSS 0.132855f
C11655 VDAC_P.t2048 VSS 0.10586f
C11656 VDAC_P.n1090 VSS 0.132855f
C11657 VDAC_P.t1987 VSS 0.10586f
C11658 VDAC_P.n1091 VSS 0.132855f
C11659 VDAC_P.t1160 VSS 0.10586f
C11660 VDAC_P.n1092 VSS 0.132855f
C11661 VDAC_P.t1746 VSS 0.10586f
C11662 VDAC_P.n1093 VSS 0.132855f
C11663 VDAC_P.t1428 VSS 0.10586f
C11664 VDAC_P.n1094 VSS 0.132855f
C11665 VDAC_P.t350 VSS 0.10586f
C11666 VDAC_P.n1095 VSS 0.132855f
C11667 VDAC_P.t585 VSS 0.10586f
C11668 VDAC_P.n1096 VSS 0.132855f
C11669 VDAC_P.t562 VSS 0.10586f
C11670 VDAC_P.n1097 VSS 0.132855f
C11671 VDAC_P.t278 VSS 0.10586f
C11672 VDAC_P.n1098 VSS 0.132855f
C11673 VDAC_P.t1288 VSS 0.10586f
C11674 VDAC_P.n1099 VSS 0.132855f
C11675 VDAC_P.t918 VSS 0.10586f
C11676 VDAC_P.n1100 VSS 0.132855f
C11677 VDAC_P.t703 VSS 0.10586f
C11678 VDAC_P.n1101 VSS 0.132855f
C11679 VDAC_P.t790 VSS 0.10586f
C11680 VDAC_P.n1102 VSS 0.132855f
C11681 VDAC_P.t361 VSS 0.10586f
C11682 VDAC_P.n1103 VSS 0.132855f
C11683 VDAC_P.t251 VSS 0.10586f
C11684 VDAC_P.n1104 VSS 0.132855f
C11685 VDAC_P.t63 VSS 0.10586f
C11686 VDAC_P.n1105 VSS 0.132855f
C11687 VDAC_P.t815 VSS 0.10586f
C11688 VDAC_P.n1106 VSS 0.132855f
C11689 VDAC_P.t1180 VSS 0.10586f
C11690 VDAC_P.n1107 VSS 0.132855f
C11691 VDAC_P.t1495 VSS 0.10586f
C11692 VDAC_P.n1108 VSS 0.132855f
C11693 VDAC_P.t1949 VSS 0.10586f
C11694 VDAC_P.n1109 VSS 0.132855f
C11695 VDAC_P.t705 VSS 0.10586f
C11696 VDAC_P.n1110 VSS 0.132855f
C11697 VDAC_P.t1839 VSS 0.10586f
C11698 VDAC_P.n1111 VSS 0.132855f
C11699 VDAC_P.t580 VSS 0.10586f
C11700 VDAC_P.n1112 VSS 0.132855f
C11701 VDAC_P.t1733 VSS 0.10586f
C11702 VDAC_P.n1113 VSS 0.132855f
C11703 VDAC_P.t572 VSS 0.10586f
C11704 VDAC_P.n1114 VSS 0.132855f
C11705 VDAC_P.t2024 VSS 0.10586f
C11706 VDAC_P.n1115 VSS 0.132855f
C11707 VDAC_P.t89 VSS 0.10586f
C11708 VDAC_P.n1116 VSS 0.132855f
C11709 VDAC_P.t816 VSS 0.10586f
C11710 VDAC_P.n1117 VSS 0.132855f
C11711 VDAC_P.t947 VSS 0.10586f
C11712 VDAC_P.n1118 VSS 0.132855f
C11713 VDAC_P.t708 VSS 0.10586f
C11714 VDAC_P.n1119 VSS 0.132855f
C11715 VDAC_P.t1534 VSS 0.10586f
C11716 VDAC_P.n1120 VSS 0.132855f
C11717 VDAC_P.t1020 VSS 0.10586f
C11718 VDAC_P.n1121 VSS 0.132855f
C11719 VDAC_P.t1086 VSS 0.10586f
C11720 VDAC_P.n1122 VSS 0.132855f
C11721 VDAC_P.t305 VSS 0.10586f
C11722 VDAC_P.n1123 VSS 0.132855f
C11723 VDAC_P.t240 VSS 0.10586f
C11724 VDAC_P.n1124 VSS 0.12686f
C11725 VDAC_P.t1219 VSS 0.10586f
C11726 VDAC_P.n1125 VSS 0.132855f
C11727 VDAC_P.t1769 VSS 0.10586f
C11728 VDAC_P.n1126 VSS 0.132855f
C11729 VDAC_P.t565 VSS 0.10586f
C11730 VDAC_P.n1127 VSS 0.132855f
C11731 VDAC_P.t31 VSS 0.10586f
C11732 VDAC_P.n1128 VSS 0.132855f
C11733 VDAC_P.t2017 VSS 0.10586f
C11734 VDAC_P.n1129 VSS 0.132855f
C11735 VDAC_P.t385 VSS 0.10586f
C11736 VDAC_P.n1130 VSS 0.132855f
C11737 VDAC_P.t263 VSS 0.10586f
C11738 VDAC_P.n1131 VSS 0.132855f
C11739 VDAC_P.t1716 VSS 0.10586f
C11740 VDAC_P.n1132 VSS 0.132855f
C11741 VDAC_P.t1803 VSS 0.10586f
C11742 VDAC_P.n1133 VSS 0.132855f
C11743 VDAC_P.t1580 VSS 0.10586f
C11744 VDAC_P.n1134 VSS 0.132855f
C11745 VDAC_P.t419 VSS 0.10586f
C11746 VDAC_P.n1135 VSS 0.132855f
C11747 VDAC_P.t1372 VSS 0.10586f
C11748 VDAC_P.n1136 VSS 0.132855f
C11749 VDAC_P.t1864 VSS 0.10586f
C11750 VDAC_P.n1137 VSS 0.132855f
C11751 VDAC_P.t1089 VSS 0.10586f
C11752 VDAC_P.n1138 VSS 0.132855f
C11753 VDAC_P.t1555 VSS 0.10586f
C11754 VDAC_P.n1139 VSS 0.132855f
C11755 VDAC_P.t1069 VSS 0.10586f
C11756 VDAC_P.n1140 VSS 0.132855f
C11757 VDAC_P.t1441 VSS 0.10586f
C11758 VDAC_P.n1141 VSS 0.132855f
C11759 VDAC_P.t1897 VSS 0.10586f
C11760 VDAC_P.n1142 VSS 0.132855f
C11761 VDAC_P.t1248 VSS 0.10586f
C11762 VDAC_P.n1143 VSS 0.132855f
C11763 VDAC_P.t1793 VSS 0.10586f
C11764 VDAC_P.n1144 VSS 0.132855f
C11765 VDAC_P.t748 VSS 0.10586f
C11766 VDAC_P.n1145 VSS 0.132855f
C11767 VDAC_P.t443 VSS 0.10586f
C11768 VDAC_P.n1146 VSS 0.132855f
C11769 VDAC_P.t2114 VSS 0.10586f
C11770 VDAC_P.n1147 VSS 0.132855f
C11771 VDAC_P.t1832 VSS 0.10586f
C11772 VDAC_P.n1148 VSS 0.132855f
C11773 VDAC_P.t977 VSS 0.10586f
C11774 VDAC_P.n1149 VSS 0.132855f
C11775 VDAC_P.t1368 VSS 0.10586f
C11776 VDAC_P.n1150 VSS 0.132855f
C11777 VDAC_P.t1634 VSS 0.10586f
C11778 VDAC_P.n1151 VSS 0.132855f
C11779 VDAC_P.t972 VSS 0.10586f
C11780 VDAC_P.n1152 VSS 0.132855f
C11781 VDAC_P.t1418 VSS 0.10586f
C11782 VDAC_P.n1153 VSS 0.132855f
C11783 VDAC_P.t9 VSS 0.10586f
C11784 VDAC_P.n1154 VSS 0.132855f
C11785 VDAC_P.t504 VSS 0.10586f
C11786 VDAC_P.n1155 VSS 0.132855f
C11787 VDAC_P.t17 VSS 0.10586f
C11788 VDAC_P.n1156 VSS 0.132855f
C11789 VDAC_P.t1504 VSS 0.10586f
C11790 VDAC_P.n1157 VSS 0.132855f
C11791 VDAC_P.t54 VSS 0.10586f
C11792 VDAC_P.n1158 VSS 0.132855f
C11793 VDAC_P.t1331 VSS 0.10586f
C11794 VDAC_P.n1159 VSS 0.132855f
C11795 VDAC_P.t758 VSS 0.10586f
C11796 VDAC_P.n1160 VSS 0.132855f
C11797 VDAC_P.t1227 VSS 0.10586f
C11798 VDAC_P.n1161 VSS 0.132855f
C11799 VDAC_P.t2064 VSS 0.10586f
C11800 VDAC_P.n1162 VSS 0.132855f
C11801 VDAC_P.t299 VSS 0.10586f
C11802 VDAC_P.n1163 VSS 0.132855f
C11803 VDAC_P.t1571 VSS 0.10586f
C11804 VDAC_P.n1164 VSS 0.132855f
C11805 VDAC_P.t1926 VSS 0.10586f
C11806 VDAC_P.n1165 VSS 0.132855f
C11807 VDAC_P.t123 VSS 0.10586f
C11808 VDAC_P.n1166 VSS 0.132855f
C11809 VDAC_P.t1015 VSS 0.10586f
C11810 VDAC_P.n1167 VSS 0.132855f
C11811 VDAC_P.t681 VSS 0.10586f
C11812 VDAC_P.n1168 VSS 0.132855f
C11813 VDAC_P.t83 VSS 0.10586f
C11814 VDAC_P.n1169 VSS 0.132855f
C11815 VDAC_P.t52 VSS 0.10586f
C11816 VDAC_P.n1170 VSS 0.132855f
C11817 VDAC_P.t1683 VSS 0.10586f
C11818 VDAC_P.n1171 VSS 0.132855f
C11819 VDAC_P.t864 VSS 0.10586f
C11820 VDAC_P.n1172 VSS 0.132855f
C11821 VDAC_P.t801 VSS 0.10586f
C11822 VDAC_P.n1173 VSS 0.132855f
C11823 VDAC_P.t529 VSS 0.10586f
C11824 VDAC_P.n1174 VSS 0.132855f
C11825 VDAC_P.t1352 VSS 0.10586f
C11826 VDAC_P.n1175 VSS 0.132855f
C11827 VDAC_P.t1919 VSS 0.10586f
C11828 VDAC_P.n1176 VSS 0.132855f
C11829 VDAC_P.t932 VSS 0.10586f
C11830 VDAC_P.n1177 VSS 0.132855f
C11831 VDAC_P.t114 VSS 0.10586f
C11832 VDAC_P.n1178 VSS 0.132855f
C11833 VDAC_P.t796 VSS 0.10586f
C11834 VDAC_P.n1179 VSS 0.132855f
C11835 VDAC_P.t1190 VSS 0.10586f
C11836 VDAC_P.n1180 VSS 0.132855f
C11837 VDAC_P.t2057 VSS 0.10586f
C11838 VDAC_P.n1181 VSS 0.132855f
C11839 VDAC_P.t1488 VSS 0.10586f
C11840 VDAC_P.n1182 VSS 0.132855f
C11841 VDAC_P.t1906 VSS 0.10586f
C11842 VDAC_P.n1183 VSS 0.132855f
C11843 VDAC_P.t1044 VSS 0.10586f
C11844 VDAC_P.n1184 VSS 0.132855f
C11845 VDAC_P.t754 VSS 0.10586f
C11846 VDAC_P.n1185 VSS 0.132855f
C11847 VDAC_P.t1325 VSS 0.10586f
C11848 VDAC_P.n1186 VSS 0.132855f
C11849 VDAC_P.t1250 VSS 0.10586f
C11850 VDAC_P.n1187 VSS 0.12686f
C11851 VDAC_P.t1981 VSS 0.10586f
C11852 VDAC_P.n1188 VSS 0.132855f
C11853 VDAC_P.t1608 VSS 0.10586f
C11854 VDAC_P.n1189 VSS 0.132855f
C11855 VDAC_P.t143 VSS 0.10586f
C11856 VDAC_P.n1190 VSS 0.132855f
C11857 VDAC_P.t1396 VSS 0.10586f
C11858 VDAC_P.n1191 VSS 0.132855f
C11859 VDAC_P.t1306 VSS 0.10586f
C11860 VDAC_P.n1192 VSS 0.132855f
C11861 VDAC_P.t60 VSS 0.10586f
C11862 VDAC_P.n1193 VSS 0.132855f
C11863 VDAC_P.t558 VSS 0.10586f
C11864 VDAC_P.n1194 VSS 0.132855f
C11865 VDAC_P.t1022 VSS 0.10586f
C11866 VDAC_P.n1195 VSS 0.132855f
C11867 VDAC_P.t1728 VSS 0.10586f
C11868 VDAC_P.n1196 VSS 0.132855f
C11869 VDAC_P.t1798 VSS 0.10586f
C11870 VDAC_P.n1197 VSS 0.132855f
C11871 VDAC_P.t436 VSS 0.10586f
C11872 VDAC_P.n1198 VSS 0.132855f
C11873 VDAC_P.t1578 VSS 0.10586f
C11874 VDAC_P.n1199 VSS 0.132855f
C11875 VDAC_P.t1267 VSS 0.10586f
C11876 VDAC_P.n1200 VSS 0.132855f
C11877 VDAC_P.t1281 VSS 0.10586f
C11878 VDAC_P.n1201 VSS 0.132855f
C11879 VDAC_P.t1737 VSS 0.10586f
C11880 VDAC_P.n1202 VSS 0.132855f
C11881 VDAC_P.t596 VSS 0.10586f
C11882 VDAC_P.n1203 VSS 0.132855f
C11883 VDAC_P.t229 VSS 0.10586f
C11884 VDAC_P.n1204 VSS 0.132855f
C11885 VDAC_P.t2085 VSS 0.10586f
C11886 VDAC_P.n1205 VSS 0.132855f
C11887 VDAC_P.t280 VSS 0.10586f
C11888 VDAC_P.n1206 VSS 0.132855f
C11889 VDAC_P.t1007 VSS 0.10586f
C11890 VDAC_P.n1207 VSS 0.132855f
C11891 VDAC_P.t592 VSS 0.10586f
C11892 VDAC_P.n1208 VSS 0.132855f
C11893 VDAC_P.t1869 VSS 0.10586f
C11894 VDAC_P.n1209 VSS 0.132855f
C11895 VDAC_P.t724 VSS 0.10586f
C11896 VDAC_P.n1210 VSS 0.132855f
C11897 VDAC_P.t1314 VSS 0.10586f
C11898 VDAC_P.n1211 VSS 0.132855f
C11899 VDAC_P.t2119 VSS 0.10586f
C11900 VDAC_P.n1212 VSS 0.132855f
C11901 VDAC_P.t1094 VSS 0.10586f
C11902 VDAC_P.n1213 VSS 0.132855f
C11903 VDAC_P.t2026 VSS 0.10586f
C11904 VDAC_P.n1214 VSS 0.132855f
C11905 VDAC_P.t1280 VSS 0.10586f
C11906 VDAC_P.n1215 VSS 0.132855f
C11907 VDAC_P.t1806 VSS 0.10586f
C11908 VDAC_P.n1216 VSS 0.132855f
C11909 VDAC_P.t1684 VSS 0.10586f
C11910 VDAC_P.n1217 VSS 0.132855f
C11911 VDAC_P.t362 VSS 0.10586f
C11912 VDAC_P.n1218 VSS 0.132855f
C11913 VDAC_P.t1271 VSS 0.10586f
C11914 VDAC_P.n1219 VSS 0.132855f
C11915 VDAC_P.t310 VSS 0.10586f
C11916 VDAC_P.n1220 VSS 0.132855f
C11917 VDAC_P.t2074 VSS 0.10586f
C11918 VDAC_P.n1221 VSS 0.132855f
C11919 VDAC_P.t773 VSS 0.10586f
C11920 VDAC_P.n1222 VSS 0.132855f
C11921 VDAC_P.t946 VSS 0.10586f
C11922 VDAC_P.n1223 VSS 0.132855f
C11923 VDAC_P.t1403 VSS 0.10586f
C11924 VDAC_P.n1224 VSS 0.132855f
C11925 VDAC_P.t730 VSS 0.10586f
C11926 VDAC_P.n1225 VSS 0.132855f
C11927 VDAC_P.t1301 VSS 0.10586f
C11928 VDAC_P.n1226 VSS 0.132855f
C11929 VDAC_P.t55 VSS 0.10586f
C11930 VDAC_P.n1227 VSS 0.132855f
C11931 VDAC_P.t601 VSS 0.10586f
C11932 VDAC_P.n1228 VSS 0.132855f
C11933 VDAC_P.t1731 VSS 0.10586f
C11934 VDAC_P.n1229 VSS 0.132855f
C11935 VDAC_P.t1084 VSS 0.10586f
C11936 VDAC_P.n1230 VSS 0.132855f
C11937 VDAC_P.t1523 VSS 0.10586f
C11938 VDAC_P.n1231 VSS 0.132855f
C11939 VDAC_P.t1979 VSS 0.10586f
C11940 VDAC_P.n1232 VSS 0.132855f
C11941 VDAC_P.t1592 VSS 0.10586f
C11942 VDAC_P.n1233 VSS 0.132855f
C11943 VDAC_P.t487 VSS 0.10586f
C11944 VDAC_P.n1234 VSS 0.132855f
C11945 VDAC_P.t1380 VSS 0.10586f
C11946 VDAC_P.n1235 VSS 0.132855f
C11947 VDAC_P.t1759 VSS 0.10586f
C11948 VDAC_P.n1236 VSS 0.132855f
C11949 VDAC_P.t508 VSS 0.10586f
C11950 VDAC_P.n1237 VSS 0.132855f
C11951 VDAC_P.t94 VSS 0.10586f
C11952 VDAC_P.n1238 VSS 0.132855f
C11953 VDAC_P.t2107 VSS 0.10586f
C11954 VDAC_P.n1239 VSS 0.132855f
C11955 VDAC_P.t1720 VSS 0.10586f
C11956 VDAC_P.n1240 VSS 0.132855f
C11957 VDAC_P.t138 VSS 0.10586f
C11958 VDAC_P.n1241 VSS 0.132855f
C11959 VDAC_P.t836 VSS 0.10586f
C11960 VDAC_P.n1242 VSS 0.132855f
C11961 VDAC_P.t802 VSS 0.10586f
C11962 VDAC_P.n1243 VSS 0.132855f
C11963 VDAC_P.t1452 VSS 0.10586f
C11964 VDAC_P.n1244 VSS 0.132855f
C11965 VDAC_P.t98 VSS 0.10586f
C11966 VDAC_P.n1245 VSS 0.132855f
C11967 VDAC_P.t99 VSS 0.10586f
C11968 VDAC_P.n1246 VSS 0.132855f
C11969 VDAC_P.t928 VSS 0.10586f
C11970 VDAC_P.n1247 VSS 0.132855f
C11971 VDAC_P.t942 VSS 0.10586f
C11972 VDAC_P.n1248 VSS 0.132855f
C11973 VDAC_P.t399 VSS 0.10586f
C11974 VDAC_P.n1249 VSS 0.132855f
C11975 VDAC_P.t830 VSS 0.10586f
C11976 VDAC_P.n1250 VSS 0.12686f
C11977 VDAC_P.t1702 VSS 0.10586f
C11978 VDAC_P.n1251 VSS 0.132855f
C11979 VDAC_P.t1435 VSS 0.10586f
C11980 VDAC_P.n1252 VSS 0.132855f
C11981 VDAC_P.t1498 VSS 0.10586f
C11982 VDAC_P.n1253 VSS 0.132855f
C11983 VDAC_P.t1231 VSS 0.10586f
C11984 VDAC_P.n1254 VSS 0.132855f
C11985 VDAC_P.t1685 VSS 0.10586f
C11986 VDAC_P.n1255 VSS 0.132855f
C11987 VDAC_P.t1117 VSS 0.10586f
C11988 VDAC_P.n1256 VSS 0.132855f
C11989 VDAC_P.t415 VSS 0.10586f
C11990 VDAC_P.n1257 VSS 0.132855f
C11991 VDAC_P.t2033 VSS 0.10586f
C11992 VDAC_P.n1258 VSS 0.132855f
C11993 VDAC_P.t749 VSS 0.10586f
C11994 VDAC_P.n1259 VSS 0.132855f
C11995 VDAC_P.t975 VSS 0.10586f
C11996 VDAC_P.n1260 VSS 0.132855f
C11997 VDAC_P.t335 VSS 0.10586f
C11998 VDAC_P.n1261 VSS 0.132855f
C11999 VDAC_P.t1815 VSS 0.10586f
C12000 VDAC_P.n1262 VSS 0.132855f
C12001 VDAC_P.t940 VSS 0.10586f
C12002 VDAC_P.n1263 VSS 0.132855f
C12003 VDAC_P.t294 VSS 0.10586f
C12004 VDAC_P.n1264 VSS 0.132855f
C12005 VDAC_P.t526 VSS 0.10586f
C12006 VDAC_P.n1265 VSS 0.132855f
C12007 VDAC_P.t809 VSS 0.10586f
C12008 VDAC_P.n1266 VSS 0.132855f
C12009 VDAC_P.t914 VSS 0.10586f
C12010 VDAC_P.n1267 VSS 0.132855f
C12011 VDAC_P.t1375 VSS 0.10586f
C12012 VDAC_P.n1268 VSS 0.132855f
C12013 VDAC_P.t983 VSS 0.10586f
C12014 VDAC_P.n1269 VSS 0.132855f
C12015 VDAC_P.t183 VSS 0.10586f
C12016 VDAC_P.n1270 VSS 0.132855f
C12017 VDAC_P.t877 VSS 0.10586f
C12018 VDAC_P.n1271 VSS 0.132855f
C12019 VDAC_P.t597 VSS 0.10586f
C12020 VDAC_P.n1272 VSS 0.132855f
C12021 VDAC_P.t227 VSS 0.10586f
C12022 VDAC_P.n1273 VSS 0.132855f
C12023 VDAC_P.t2075 VSS 0.10586f
C12024 VDAC_P.n1274 VSS 0.132855f
C12025 VDAC_P.t1401 VSS 0.10586f
C12026 VDAC_P.n1275 VSS 0.132855f
C12027 VDAC_P.t1969 VSS 0.10586f
C12028 VDAC_P.n1276 VSS 0.132855f
C12029 VDAC_P.t1112 VSS 0.10586f
C12030 VDAC_P.n1277 VSS 0.132855f
C12031 VDAC_P.t891 VSS 0.10586f
C12032 VDAC_P.n1278 VSS 0.132855f
C12033 VDAC_P.t1316 VSS 0.10586f
C12034 VDAC_P.n1279 VSS 0.132855f
C12035 VDAC_P.t1651 VSS 0.10586f
C12036 VDAC_P.n1280 VSS 0.132855f
C12037 VDAC_P.t1065 VSS 0.10586f
C12038 VDAC_P.n1281 VSS 0.132855f
C12039 VDAC_P.t1064 VSS 0.10586f
C12040 VDAC_P.n1282 VSS 0.132855f
C12041 VDAC_P.t1999 VSS 0.10586f
C12042 VDAC_P.n1283 VSS 0.132855f
C12043 VDAC_P.t624 VSS 0.10586f
C12044 VDAC_P.n1284 VSS 0.132855f
C12045 VDAC_P.t1566 VSS 0.10586f
C12046 VDAC_P.n1285 VSS 0.132855f
C12047 VDAC_P.t1540 VSS 0.10586f
C12048 VDAC_P.n1286 VSS 0.132855f
C12049 VDAC_P.t686 VSS 0.10586f
C12050 VDAC_P.n1287 VSS 0.132855f
C12051 VDAC_P.t95 VSS 0.10586f
C12052 VDAC_P.n1288 VSS 0.132855f
C12053 VDAC_P.t302 VSS 0.10586f
C12054 VDAC_P.n1289 VSS 0.132855f
C12055 VDAC_P.t2050 VSS 0.10586f
C12056 VDAC_P.n1290 VSS 0.132855f
C12057 VDAC_P.t872 VSS 0.10586f
C12058 VDAC_P.n1291 VSS 0.132855f
C12059 VDAC_P.t2006 VSS 0.10586f
C12060 VDAC_P.n1292 VSS 0.132855f
C12061 VDAC_P.t1479 VSS 0.10586f
C12062 VDAC_P.n1293 VSS 0.132855f
C12063 VDAC_P.t414 VSS 0.10586f
C12064 VDAC_P.n1294 VSS 0.132855f
C12065 VDAC_P.t1265 VSS 0.10586f
C12066 VDAC_P.n1295 VSS 0.132855f
C12067 VDAC_P.t1823 VSS 0.10586f
C12068 VDAC_P.n1296 VSS 0.132855f
C12069 VDAC_P.t1161 VSS 0.10586f
C12070 VDAC_P.n1297 VSS 0.132855f
C12071 VDAC_P.t1617 VSS 0.10586f
C12072 VDAC_P.n1298 VSS 0.132855f
C12073 VDAC_P.t2058 VSS 0.10586f
C12074 VDAC_P.n1299 VSS 0.132855f
C12075 VDAC_P.t1511 VSS 0.10586f
C12076 VDAC_P.n1300 VSS 0.132855f
C12077 VDAC_P.t995 VSS 0.10586f
C12078 VDAC_P.n1301 VSS 0.132855f
C12079 VDAC_P.t711 VSS 0.10586f
C12080 VDAC_P.n1302 VSS 0.132855f
C12081 VDAC_P.t1853 VSS 0.10586f
C12082 VDAC_P.n1303 VSS 0.132855f
C12083 VDAC_P.t1252 VSS 0.10586f
C12084 VDAC_P.n1304 VSS 0.132855f
C12085 VDAC_P.t1647 VSS 0.10586f
C12086 VDAC_P.n1305 VSS 0.132855f
C12087 VDAC_P.t764 VSS 0.10586f
C12088 VDAC_P.n1306 VSS 0.132855f
C12089 VDAC_P.t783 VSS 0.10586f
C12090 VDAC_P.n1307 VSS 0.132855f
C12091 VDAC_P.t151 VSS 0.10586f
C12092 VDAC_P.n1308 VSS 0.132855f
C12093 VDAC_P.t1664 VSS 0.10586f
C12094 VDAC_P.n1309 VSS 0.132855f
C12095 VDAC_P.t1883 VSS 0.10586f
C12096 VDAC_P.n1310 VSS 0.132855f
C12097 VDAC_P.t1508 VSS 0.10586f
C12098 VDAC_P.n1311 VSS 0.132855f
C12099 VDAC_P.t1558 VSS 0.10586f
C12100 VDAC_P.n1312 VSS 0.132855f
C12101 VDAC_P.t620 VSS 0.10586f
C12102 VDAC_P.n1313 VSS 0.12686f
C12103 VDAC_P.t1645 VSS 0.10586f
C12104 VDAC_P.n1314 VSS 0.132855f
C12105 VDAC_P.t1468 VSS 0.10586f
C12106 VDAC_P.n1315 VSS 0.132855f
C12107 VDAC_P.t405 VSS 0.10586f
C12108 VDAC_P.n1316 VSS 0.132855f
C12109 VDAC_P.t1011 VSS 0.10586f
C12110 VDAC_P.n1317 VSS 0.132855f
C12111 VDAC_P.t1184 VSS 0.10586f
C12112 VDAC_P.n1318 VSS 0.132855f
C12113 VDAC_P.t1881 VSS 0.10586f
C12114 VDAC_P.n1319 VSS 0.132855f
C12115 VDAC_P.t1492 VSS 0.10586f
C12116 VDAC_P.n1320 VSS 0.132855f
C12117 VDAC_P.t1326 VSS 0.10586f
C12118 VDAC_P.n1321 VSS 0.132855f
C12119 VDAC_P.t172 VSS 0.10586f
C12120 VDAC_P.n1322 VSS 0.132855f
C12121 VDAC_P.t1110 VSS 0.10586f
C12122 VDAC_P.n1323 VSS 0.132855f
C12123 VDAC_P.t1027 VSS 0.10586f
C12124 VDAC_P.n1324 VSS 0.132855f
C12125 VDAC_P.t1776 VSS 0.10586f
C12126 VDAC_P.n1325 VSS 0.132855f
C12127 VDAC_P.t1822 VSS 0.10586f
C12128 VDAC_P.n1326 VSS 0.132855f
C12129 VDAC_P.t210 VSS 0.10586f
C12130 VDAC_P.n1327 VSS 0.132855f
C12131 VDAC_P.t327 VSS 0.10586f
C12132 VDAC_P.n1328 VSS 0.132855f
C12133 VDAC_P.t1777 VSS 0.10586f
C12134 VDAC_P.n1329 VSS 0.132855f
C12135 VDAC_P.t1109 VSS 0.10586f
C12136 VDAC_P.n1330 VSS 0.132855f
C12137 VDAC_P.t413 VSS 0.10586f
C12138 VDAC_P.n1331 VSS 0.132855f
C12139 VDAC_P.t291 VSS 0.10586f
C12140 VDAC_P.n1332 VSS 0.132855f
C12141 VDAC_P.t745 VSS 0.10586f
C12142 VDAC_P.n1333 VSS 0.132855f
C12143 VDAC_P.t1915 VSS 0.10586f
C12144 VDAC_P.n1334 VSS 0.132855f
C12145 VDAC_P.t111 VSS 0.10586f
C12146 VDAC_P.n1335 VSS 0.132855f
C12147 VDAC_P.t1807 VSS 0.10586f
C12148 VDAC_P.n1336 VSS 0.132855f
C12149 VDAC_P.t1708 VSS 0.10586f
C12150 VDAC_P.n1337 VSS 0.132855f
C12151 VDAC_P.t813 VSS 0.10586f
C12152 VDAC_P.n1338 VSS 0.132855f
C12153 VDAC_P.t1948 VSS 0.10586f
C12154 VDAC_P.n1339 VSS 0.132855f
C12155 VDAC_P.t960 VSS 0.10586f
C12156 VDAC_P.n1340 VSS 0.132855f
C12157 VDAC_P.t987 VSS 0.10586f
C12158 VDAC_P.n1341 VSS 0.132855f
C12159 VDAC_P.t1448 VSS 0.10586f
C12160 VDAC_P.n1342 VSS 0.132855f
C12161 VDAC_P.t141 VSS 0.10586f
C12162 VDAC_P.n1343 VSS 0.132855f
C12163 VDAC_P.t564 VSS 0.10586f
C12164 VDAC_P.n1344 VSS 0.132855f
C12165 VDAC_P.t742 VSS 0.10586f
C12166 VDAC_P.n1345 VSS 0.132855f
C12167 VDAC_P.t554 VSS 0.10586f
C12168 VDAC_P.n1346 VSS 0.132855f
C12169 VDAC_P.t2008 VSS 0.10586f
C12170 VDAC_P.n1347 VSS 0.132855f
C12171 VDAC_P.t1950 VSS 0.10586f
C12172 VDAC_P.n1348 VSS 0.132855f
C12173 VDAC_P.t1576 VSS 0.10586f
C12174 VDAC_P.n1349 VSS 0.132855f
C12175 VDAC_P.t1730 VSS 0.10586f
C12176 VDAC_P.n1350 VSS 0.132855f
C12177 VDAC_P.t196 VSS 0.10586f
C12178 VDAC_P.n1351 VSS 0.132855f
C12179 VDAC_P.t1522 VSS 0.10586f
C12180 VDAC_P.n1352 VSS 0.132855f
C12181 VDAC_P.t331 VSS 0.10586f
C12182 VDAC_P.n1353 VSS 0.132855f
C12183 VDAC_P.t1246 VSS 0.10586f
C12184 VDAC_P.n1354 VSS 0.132855f
C12185 VDAC_P.t623 VSS 0.10586f
C12186 VDAC_P.n1355 VSS 0.132855f
C12187 VDAC_P.t1671 VSS 0.10586f
C12188 VDAC_P.n1356 VSS 0.132855f
C12189 VDAC_P.t994 VSS 0.10586f
C12190 VDAC_P.n1357 VSS 0.132855f
C12191 VDAC_P.t1457 VSS 0.10586f
C12192 VDAC_P.n1358 VSS 0.132855f
C12193 VDAC_P.t525 VSS 0.10586f
C12194 VDAC_P.n1359 VSS 0.132855f
C12195 VDAC_P.t689 VSS 0.10586f
C12196 VDAC_P.n1360 VSS 0.132855f
C12197 VDAC_P.t139 VSS 0.10586f
C12198 VDAC_P.n1361 VSS 0.132855f
C12199 VDAC_P.t1245 VSS 0.10586f
C12200 VDAC_P.n1362 VSS 0.132855f
C12201 VDAC_P.t1699 VSS 0.10586f
C12202 VDAC_P.n1363 VSS 0.132855f
C12203 VDAC_P.t348 VSS 0.10586f
C12204 VDAC_P.n1364 VSS 0.132855f
C12205 VDAC_P.t1589 VSS 0.10586f
C12206 VDAC_P.n1365 VSS 0.132855f
C12207 VDAC_P.t2045 VSS 0.10586f
C12208 VDAC_P.n1366 VSS 0.132855f
C12209 VDAC_P.t1416 VSS 0.10586f
C12210 VDAC_P.n1367 VSS 0.132855f
C12211 VDAC_P.t1831 VSS 0.10586f
C12212 VDAC_P.n1368 VSS 0.132855f
C12213 VDAC_P.t1956 VSS 0.10586f
C12214 VDAC_P.n1369 VSS 0.132855f
C12215 VDAC_P.t1725 VSS 0.10586f
C12216 VDAC_P.n1370 VSS 0.132855f
C12217 VDAC_P.t2130 VSS 0.10586f
C12218 VDAC_P.n1371 VSS 0.132855f
C12219 VDAC_P.t1222 VSS 0.10586f
C12220 VDAC_P.n1372 VSS 0.132855f
C12221 VDAC_P.t1051 VSS 0.10586f
C12222 VDAC_P.n1373 VSS 0.132855f
C12223 VDAC_P.t1552 VSS 0.10586f
C12224 VDAC_P.n1374 VSS 0.132855f
C12225 VDAC_P.t1934 VSS 0.10586f
C12226 VDAC_P.n1375 VSS 0.132855f
C12227 VDAC_P.t568 VSS 0.10586f
C12228 VDAC_P.n1376 VSS 0.12686f
C12229 VDAC_P.t1024 VSS 0.10586f
C12230 VDAC_P.n1377 VSS 0.132855f
C12231 VDAC_P.t1097 VSS 0.10586f
C12232 VDAC_P.n1378 VSS 0.132855f
C12233 VDAC_P.t224 VSS 0.10586f
C12234 VDAC_P.n1379 VSS 0.132855f
C12235 VDAC_P.t882 VSS 0.10586f
C12236 VDAC_P.n1380 VSS 0.132855f
C12237 VDAC_P.t193 VSS 0.10586f
C12238 VDAC_P.n1381 VSS 0.132855f
C12239 VDAC_P.t1530 VSS 0.10586f
C12240 VDAC_P.n1382 VSS 0.132855f
C12241 VDAC_P.t635 VSS 0.10586f
C12242 VDAC_P.n1383 VSS 0.132855f
C12243 VDAC_P.t1695 VSS 0.10586f
C12244 VDAC_P.n1384 VSS 0.132855f
C12245 VDAC_P.t1135 VSS 0.10586f
C12246 VDAC_P.n1385 VSS 0.132855f
C12247 VDAC_P.t417 VSS 0.10586f
C12248 VDAC_P.n1386 VSS 0.132855f
C12249 VDAC_P.t1790 VSS 0.10586f
C12250 VDAC_P.n1387 VSS 0.132855f
C12251 VDAC_P.t1481 VSS 0.10586f
C12252 VDAC_P.n1388 VSS 0.132855f
C12253 VDAC_P.t1933 VSS 0.10586f
C12254 VDAC_P.n1389 VSS 0.132855f
C12255 VDAC_P.t1244 VSS 0.10586f
C12256 VDAC_P.n1390 VSS 0.132855f
C12257 VDAC_P.t1872 VSS 0.10586f
C12258 VDAC_P.n1391 VSS 0.132855f
C12259 VDAC_P.t1058 VSS 0.10586f
C12260 VDAC_P.n1392 VSS 0.132855f
C12261 VDAC_P.t376 VSS 0.10586f
C12262 VDAC_P.n1393 VSS 0.132855f
C12263 VDAC_P.t1654 VSS 0.10586f
C12264 VDAC_P.n1394 VSS 0.132855f
C12265 VDAC_P.t1409 VSS 0.10586f
C12266 VDAC_P.n1395 VSS 0.132855f
C12267 VDAC_P.t1442 VSS 0.10586f
C12268 VDAC_P.n1396 VSS 0.132855f
C12269 VDAC_P.t1205 VSS 0.10586f
C12270 VDAC_P.n1397 VSS 0.132855f
C12271 VDAC_P.t178 VSS 0.10586f
C12272 VDAC_P.n1398 VSS 0.132855f
C12273 VDAC_P.t559 VSS 0.10586f
C12274 VDAC_P.n1399 VSS 0.132855f
C12275 VDAC_P.t1557 VSS 0.10586f
C12276 VDAC_P.n1400 VSS 0.132855f
C12277 VDAC_P.t1722 VSS 0.10586f
C12278 VDAC_P.n1401 VSS 0.132855f
C12279 VDAC_P.t1445 VSS 0.10586f
C12280 VDAC_P.n1402 VSS 0.132855f
C12281 VDAC_P.t1899 VSS 0.10586f
C12282 VDAC_P.n1403 VSS 0.132855f
C12283 VDAC_P.t179 VSS 0.10586f
C12284 VDAC_P.n1404 VSS 0.132855f
C12285 VDAC_P.t249 VSS 0.10586f
C12286 VDAC_P.n1405 VSS 0.132855f
C12287 VDAC_P.t577 VSS 0.10586f
C12288 VDAC_P.n1406 VSS 0.132855f
C12289 VDAC_P.t125 VSS 0.10586f
C12290 VDAC_P.n1407 VSS 0.132855f
C12291 VDAC_P.t2118 VSS 0.10586f
C12292 VDAC_P.n1408 VSS 0.132855f
C12293 VDAC_P.t751 VSS 0.10586f
C12294 VDAC_P.n1409 VSS 0.132855f
C12295 VDAC_P.t503 VSS 0.10586f
C12296 VDAC_P.n1410 VSS 0.132855f
C12297 VDAC_P.t260 VSS 0.10586f
C12298 VDAC_P.n1411 VSS 0.132855f
C12299 VDAC_P.t1821 VSS 0.10586f
C12300 VDAC_P.n1412 VSS 0.132855f
C12301 VDAC_P.t268 VSS 0.10586f
C12302 VDAC_P.n1413 VSS 0.132855f
C12303 VDAC_P.t127 VSS 0.10586f
C12304 VDAC_P.n1414 VSS 0.132855f
C12305 VDAC_P.t476 VSS 0.10586f
C12306 VDAC_P.n1415 VSS 0.132855f
C12307 VDAC_P.t984 VSS 0.10586f
C12308 VDAC_P.n1416 VSS 0.132855f
C12309 VDAC_P.t1035 VSS 0.10586f
C12310 VDAC_P.n1417 VSS 0.132855f
C12311 VDAC_P.t944 VSS 0.10586f
C12312 VDAC_P.n1418 VSS 0.132855f
C12313 VDAC_P.t1870 VSS 0.10586f
C12314 VDAC_P.n1419 VSS 0.132855f
C12315 VDAC_P.t1908 VSS 0.10586f
C12316 VDAC_P.n1420 VSS 0.132855f
C12317 VDAC_P.t1438 VSS 0.10586f
C12318 VDAC_P.n1421 VSS 0.132855f
C12319 VDAC_P.t1305 VSS 0.10586f
C12320 VDAC_P.n1422 VSS 0.132855f
C12321 VDAC_P.t102 VSS 0.10586f
C12322 VDAC_P.n1423 VSS 0.132855f
C12323 VDAC_P.t557 VSS 0.10586f
C12324 VDAC_P.n1424 VSS 0.132855f
C12325 VDAC_P.t992 VSS 0.10586f
C12326 VDAC_P.n1425 VSS 0.132855f
C12327 VDAC_P.t1930 VSS 0.10586f
C12328 VDAC_P.n1426 VSS 0.132855f
C12329 VDAC_P.t1437 VSS 0.10586f
C12330 VDAC_P.n1427 VSS 0.132855f
C12331 VDAC_P.t1706 VSS 0.10586f
C12332 VDAC_P.n1428 VSS 0.132855f
C12333 VDAC_P.t1337 VSS 0.10586f
C12334 VDAC_P.n1429 VSS 0.132855f
C12335 VDAC_P.t909 VSS 0.10586f
C12336 VDAC_P.n1430 VSS 0.132855f
C12337 VDAC_P.t301 VSS 0.10586f
C12338 VDAC_P.n1431 VSS 0.132855f
C12339 VDAC_P.t1687 VSS 0.10586f
C12340 VDAC_P.n1432 VSS 0.132855f
C12341 VDAC_P.t150 VSS 0.10586f
C12342 VDAC_P.n1433 VSS 0.132855f
C12343 VDAC_P.t389 VSS 0.10586f
C12344 VDAC_P.n1434 VSS 0.132855f
C12345 VDAC_P.t2035 VSS 0.10586f
C12346 VDAC_P.n1435 VSS 0.132855f
C12347 VDAC_P.t1363 VSS 0.10586f
C12348 VDAC_P.n1436 VSS 0.132855f
C12349 VDAC_P.t1817 VSS 0.10586f
C12350 VDAC_P.n1437 VSS 0.132855f
C12351 VDAC_P.t484 VSS 0.10586f
C12352 VDAC_P.n1438 VSS 0.132855f
C12353 VDAC_P.t869 VSS 0.10586f
C12354 VDAC_P.n1439 VSS 0.12686f
C12355 VDAC_P.t33 VSS 0.10586f
C12356 VDAC_P.n1440 VSS 0.132855f
C12357 VDAC_P.t945 VSS 0.10586f
C12358 VDAC_P.n1441 VSS 0.132855f
C12359 VDAC_P.t321 VSS 0.10586f
C12360 VDAC_P.n1442 VSS 0.132855f
C12361 VDAC_P.t1657 VSS 0.10586f
C12362 VDAC_P.n1443 VSS 0.132855f
C12363 VDAC_P.t2109 VSS 0.10586f
C12364 VDAC_P.n1444 VSS 0.132855f
C12365 VDAC_P.t409 VSS 0.10586f
C12366 VDAC_P.n1445 VSS 0.132855f
C12367 VDAC_P.t2007 VSS 0.10586f
C12368 VDAC_P.n1446 VSS 0.132855f
C12369 VDAC_P.t104 VSS 0.10586f
C12370 VDAC_P.n1447 VSS 0.132855f
C12371 VDAC_P.t961 VSS 0.10586f
C12372 VDAC_P.n1448 VSS 0.132855f
C12373 VDAC_P.t820 VSS 0.10586f
C12374 VDAC_P.n1449 VSS 0.132855f
C12375 VDAC_P.t1689 VSS 0.10586f
C12376 VDAC_P.n1450 VSS 0.132855f
C12377 VDAC_P.t716 VSS 0.10586f
C12378 VDAC_P.n1451 VSS 0.132855f
C12379 VDAC_P.t306 VSS 0.10586f
C12380 VDAC_P.n1452 VSS 0.132855f
C12381 VDAC_P.t772 VSS 0.10586f
C12382 VDAC_P.n1453 VSS 0.132855f
C12383 VDAC_P.t1334 VSS 0.10586f
C12384 VDAC_P.n1454 VSS 0.132855f
C12385 VDAC_P.t643 VSS 0.10586f
C12386 VDAC_P.n1455 VSS 0.132855f
C12387 VDAC_P.t1114 VSS 0.10586f
C12388 VDAC_P.n1456 VSS 0.132855f
C12389 VDAC_P.t1034 VSS 0.10586f
C12390 VDAC_P.n1457 VSS 0.132855f
C12391 VDAC_P.t1607 VSS 0.10586f
C12392 VDAC_P.n1458 VSS 0.132855f
C12393 VDAC_P.t926 VSS 0.10586f
C12394 VDAC_P.n1459 VSS 0.132855f
C12395 VDAC_P.t1387 VSS 0.10586f
C12396 VDAC_P.n1460 VSS 0.132855f
C12397 VDAC_P.t226 VSS 0.10586f
C12398 VDAC_P.n1461 VSS 0.132855f
C12399 VDAC_P.t655 VSS 0.10586f
C12400 VDAC_P.n1462 VSS 0.132855f
C12401 VDAC_P.t135 VSS 0.10586f
C12402 VDAC_P.n1463 VSS 0.132855f
C12403 VDAC_P.t546 VSS 0.10586f
C12404 VDAC_P.n1464 VSS 0.132855f
C12405 VDAC_P.t1637 VSS 0.10586f
C12406 VDAC_P.n1465 VSS 0.132855f
C12407 VDAC_P.t543 VSS 0.10586f
C12408 VDAC_P.n1466 VSS 0.132855f
C12409 VDAC_P.t1415 VSS 0.10586f
C12410 VDAC_P.n1467 VSS 0.132855f
C12411 VDAC_P.t273 VSS 0.10586f
C12412 VDAC_P.n1468 VSS 0.132855f
C12413 VDAC_P.t189 VSS 0.10586f
C12414 VDAC_P.n1469 VSS 0.132855f
C12415 VDAC_P.t897 VSS 0.10586f
C12416 VDAC_P.n1470 VSS 0.132855f
C12417 VDAC_P.t116 VSS 0.10586f
C12418 VDAC_P.n1471 VSS 0.132855f
C12419 VDAC_P.t1665 VSS 0.10586f
C12420 VDAC_P.n1472 VSS 0.132855f
C12421 VDAC_P.t551 VSS 0.10586f
C12422 VDAC_P.n1473 VSS 0.132855f
C12423 VDAC_P.t888 VSS 0.10586f
C12424 VDAC_P.n1474 VSS 0.132855f
C12425 VDAC_P.t1021 VSS 0.10586f
C12426 VDAC_P.n1475 VSS 0.132855f
C12427 VDAC_P.t344 VSS 0.10586f
C12428 VDAC_P.n1476 VSS 0.132855f
C12429 VDAC_P.t1799 VSS 0.10586f
C12430 VDAC_P.n1477 VSS 0.132855f
C12431 VDAC_P.t132 VSS 0.10586f
C12432 VDAC_P.n1478 VSS 0.132855f
C12433 VDAC_P.t698 VSS 0.10586f
C12434 VDAC_P.n1479 VSS 0.132855f
C12435 VDAC_P.t1132 VSS 0.10586f
C12436 VDAC_P.n1480 VSS 0.132855f
C12437 VDAC_P.t674 VSS 0.10586f
C12438 VDAC_P.n1481 VSS 0.132855f
C12439 VDAC_P.t1149 VSS 0.10586f
C12440 VDAC_P.n1482 VSS 0.132855f
C12441 VDAC_P.t136 VSS 0.10586f
C12442 VDAC_P.n1483 VSS 0.132855f
C12443 VDAC_P.t922 VSS 0.10586f
C12444 VDAC_P.n1484 VSS 0.132855f
C12445 VDAC_P.t395 VSS 0.10586f
C12446 VDAC_P.n1485 VSS 0.132855f
C12447 VDAC_P.t126 VSS 0.10586f
C12448 VDAC_P.n1486 VSS 0.132855f
C12449 VDAC_P.t1279 VSS 0.10586f
C12450 VDAC_P.n1487 VSS 0.132855f
C12451 VDAC_P.t1374 VSS 0.10586f
C12452 VDAC_P.n1488 VSS 0.132855f
C12453 VDAC_P.t1175 VSS 0.10586f
C12454 VDAC_P.n1489 VSS 0.132855f
C12455 VDAC_P.t429 VSS 0.10586f
C12456 VDAC_P.n1490 VSS 0.132855f
C12457 VDAC_P.t2086 VSS 0.10586f
C12458 VDAC_P.n1491 VSS 0.132855f
C12459 VDAC_P.t215 VSS 0.10586f
C12460 VDAC_P.n1492 VSS 0.132855f
C12461 VDAC_P.t1005 VSS 0.10586f
C12462 VDAC_P.n1493 VSS 0.132855f
C12463 VDAC_P.t349 VSS 0.10586f
C12464 VDAC_P.n1494 VSS 0.132855f
C12465 VDAC_P.t1867 VSS 0.10586f
C12466 VDAC_P.n1495 VSS 0.132855f
C12467 VDAC_P.t175 VSS 0.10586f
C12468 VDAC_P.n1496 VSS 0.132855f
C12469 VDAC_P.t845 VSS 0.10586f
C12470 VDAC_P.n1497 VSS 0.132855f
C12471 VDAC_P.t2044 VSS 0.10586f
C12472 VDAC_P.n1498 VSS 0.132855f
C12473 VDAC_P.t219 VSS 0.10586f
C12474 VDAC_P.n1499 VSS 0.132855f
C12475 VDAC_P.t2011 VSS 0.10586f
C12476 VDAC_P.n1500 VSS 0.132855f
C12477 VDAC_P.t880 VSS 0.10586f
C12478 VDAC_P.n1501 VSS 0.132855f
C12479 VDAC_P.t963 VSS 0.10586f
C12480 VDAC_P.n1502 VSS 0.12686f
C12481 VDAC_P.t283 VSS 0.10586f
C12482 VDAC_P.n1503 VSS 0.132855f
C12483 VDAC_P.t1960 VSS 0.10586f
C12484 VDAC_P.n1504 VSS 0.132855f
C12485 VDAC_P.t1965 VSS 0.10586f
C12486 VDAC_P.n1505 VSS 0.132855f
C12487 VDAC_P.t1088 VSS 0.10586f
C12488 VDAC_P.n1506 VSS 0.132855f
C12489 VDAC_P.t766 VSS 0.10586f
C12490 VDAC_P.n1507 VSS 0.132855f
C12491 VDAC_P.t340 VSS 0.10586f
C12492 VDAC_P.n1508 VSS 0.132855f
C12493 VDAC_P.t106 VSS 0.10586f
C12494 VDAC_P.n1509 VSS 0.132855f
C12495 VDAC_P.t575 VSS 0.10586f
C12496 VDAC_P.n1510 VSS 0.132855f
C12497 VDAC_P.t2080 VSS 0.10586f
C12498 VDAC_P.n1511 VSS 0.132855f
C12499 VDAC_P.t1986 VSS 0.10586f
C12500 VDAC_P.n1512 VSS 0.132855f
C12501 VDAC_P.t1208 VSS 0.10586f
C12502 VDAC_P.n1513 VSS 0.132855f
C12503 VDAC_P.t1766 VSS 0.10586f
C12504 VDAC_P.n1514 VSS 0.132855f
C12505 VDAC_P.t1365 VSS 0.10586f
C12506 VDAC_P.n1515 VSS 0.132855f
C12507 VDAC_P.t792 VSS 0.10586f
C12508 VDAC_P.n1516 VSS 0.132855f
C12509 VDAC_P.t874 VSS 0.10586f
C12510 VDAC_P.n1517 VSS 0.132855f
C12511 VDAC_P.t205 VSS 0.10586f
C12512 VDAC_P.n1518 VSS 0.132855f
C12513 VDAC_P.t1514 VSS 0.10586f
C12514 VDAC_P.n1519 VSS 0.132855f
C12515 VDAC_P.t1235 VSS 0.10586f
C12516 VDAC_P.n1520 VSS 0.132855f
C12517 VDAC_P.t1795 VSS 0.10586f
C12518 VDAC_P.n1521 VSS 0.132855f
C12519 VDAC_P.t1125 VSS 0.10586f
C12520 VDAC_P.n1522 VSS 0.132855f
C12521 VDAC_P.t1579 VSS 0.10586f
C12522 VDAC_P.n1523 VSS 0.132855f
C12523 VDAC_P.t1994 VSS 0.10586f
C12524 VDAC_P.n1524 VSS 0.132855f
C12525 VDAC_P.t1473 VSS 0.10586f
C12526 VDAC_P.n1525 VSS 0.132855f
C12527 VDAC_P.t1927 VSS 0.10586f
C12528 VDAC_P.n1526 VSS 0.132855f
C12529 VDAC_P.t1261 VSS 0.10586f
C12530 VDAC_P.n1527 VSS 0.132855f
C12531 VDAC_P.t1819 VSS 0.10586f
C12532 VDAC_P.n1528 VSS 0.132855f
C12533 VDAC_P.t1932 VSS 0.10586f
C12534 VDAC_P.n1529 VSS 0.132855f
C12535 VDAC_P.t1611 VSS 0.10586f
C12536 VDAC_P.n1530 VSS 0.132855f
C12537 VDAC_P.t290 VSS 0.10586f
C12538 VDAC_P.n1531 VSS 0.132855f
C12539 VDAC_P.t1505 VSS 0.10586f
C12540 VDAC_P.n1532 VSS 0.132855f
C12541 VDAC_P.t269 VSS 0.10586f
C12542 VDAC_P.n1533 VSS 0.132855f
C12543 VDAC_P.t1512 VSS 0.10586f
C12544 VDAC_P.n1534 VSS 0.132855f
C12545 VDAC_P.t483 VSS 0.10586f
C12546 VDAC_P.n1535 VSS 0.132855f
C12547 VDAC_P.t324 VSS 0.10586f
C12548 VDAC_P.n1536 VSS 0.132855f
C12549 VDAC_P.t646 VSS 0.10586f
C12550 VDAC_P.n1537 VSS 0.132855f
C12551 VDAC_P.t188 VSS 0.10586f
C12552 VDAC_P.n1538 VSS 0.132855f
C12553 VDAC_P.t1048 VSS 0.10586f
C12554 VDAC_P.n1539 VSS 0.132855f
C12555 VDAC_P.t1009 VSS 0.10586f
C12556 VDAC_P.n1540 VSS 0.132855f
C12557 VDAC_P.t432 VSS 0.10586f
C12558 VDAC_P.n1541 VSS 0.132855f
C12559 VDAC_P.t1758 VSS 0.10586f
C12560 VDAC_P.n1542 VSS 0.132855f
C12561 VDAC_P.t1076 VSS 0.10586f
C12562 VDAC_P.n1543 VSS 0.132855f
C12563 VDAC_P.t446 VSS 0.10586f
C12564 VDAC_P.n1544 VSS 0.132855f
C12565 VDAC_P.t1335 VSS 0.10586f
C12566 VDAC_P.n1545 VSS 0.132855f
C12567 VDAC_P.t1270 VSS 0.10586f
C12568 VDAC_P.n1546 VSS 0.132855f
C12569 VDAC_P.t1119 VSS 0.10586f
C12570 VDAC_P.n1547 VSS 0.132855f
C12571 VDAC_P.t235 VSS 0.10586f
C12572 VDAC_P.n1548 VSS 0.132855f
C12573 VDAC_P.t1002 VSS 0.10586f
C12574 VDAC_P.n1549 VSS 0.132855f
C12575 VDAC_P.t1471 VSS 0.10586f
C12576 VDAC_P.n1550 VSS 0.132855f
C12577 VDAC_P.t462 VSS 0.10586f
C12578 VDAC_P.n1551 VSS 0.132855f
C12579 VDAC_P.t695 VSS 0.10586f
C12580 VDAC_P.n1552 VSS 0.132855f
C12581 VDAC_P.t475 VSS 0.10586f
C12582 VDAC_P.n1553 VSS 0.132855f
C12583 VDAC_P.t1257 VSS 0.10586f
C12584 VDAC_P.n1554 VSS 0.132855f
C12585 VDAC_P.t1709 VSS 0.10586f
C12586 VDAC_P.n1555 VSS 0.132855f
C12587 VDAC_P.t20 VSS 0.10586f
C12588 VDAC_P.n1556 VSS 0.132855f
C12589 VDAC_P.t1501 VSS 0.10586f
C12590 VDAC_P.n1557 VSS 0.132855f
C12591 VDAC_P.t155 VSS 0.10586f
C12592 VDAC_P.n1558 VSS 0.132855f
C12593 VDAC_P.t707 VSS 0.10586f
C12594 VDAC_P.n1559 VSS 0.132855f
C12595 VDAC_P.t1845 VSS 0.10586f
C12596 VDAC_P.n1560 VSS 0.132855f
C12597 VDAC_P.t2084 VSS 0.10586f
C12598 VDAC_P.n1561 VSS 0.132855f
C12599 VDAC_P.t1739 VSS 0.10586f
C12600 VDAC_P.n1562 VSS 0.132855f
C12601 VDAC_P.t636 VSS 0.10586f
C12602 VDAC_P.n1563 VSS 0.132855f
C12603 VDAC_P.t642 VSS 0.10586f
C12604 VDAC_P.n1564 VSS 0.132855f
C12605 VDAC_P.t2087 VSS 0.10586f
C12606 VDAC_P.n1565 VSS 0.12686f
C12607 VDAC_P.t1902 VSS 0.10586f
C12608 VDAC_P.n1566 VSS 0.132855f
C12609 VDAC_P.t779 VSS 0.10586f
C12610 VDAC_P.n1567 VSS 0.132855f
C12611 VDAC_P.t1678 VSS 0.10586f
C12612 VDAC_P.n1568 VSS 0.132855f
C12613 VDAC_P.t1323 VSS 0.10586f
C12614 VDAC_P.n1569 VSS 0.132855f
C12615 VDAC_P.t899 VSS 0.10586f
C12616 VDAC_P.n1570 VSS 0.132855f
C12617 VDAC_P.t177 VSS 0.10586f
C12618 VDAC_P.n1571 VSS 0.132855f
C12619 VDAC_P.t1673 VSS 0.10586f
C12620 VDAC_P.n1572 VSS 0.132855f
C12621 VDAC_P.t159 VSS 0.10586f
C12622 VDAC_P.n1573 VSS 0.132855f
C12623 VDAC_P.t1565 VSS 0.10586f
C12624 VDAC_P.n1574 VSS 0.132855f
C12625 VDAC_P.t2019 VSS 0.10586f
C12626 VDAC_P.n1575 VSS 0.132855f
C12627 VDAC_P.t359 VSS 0.10586f
C12628 VDAC_P.n1576 VSS 0.132855f
C12629 VDAC_P.t969 VSS 0.10586f
C12630 VDAC_P.n1577 VSS 0.132855f
C12631 VDAC_P.t1732 VSS 0.10586f
C12632 VDAC_P.n1578 VSS 0.132855f
C12633 VDAC_P.t923 VSS 0.10586f
C12634 VDAC_P.n1579 VSS 0.132855f
C12635 VDAC_P.t492 VSS 0.10586f
C12636 VDAC_P.n1580 VSS 0.132855f
C12637 VDAC_P.t722 VSS 0.10586f
C12638 VDAC_P.n1581 VSS 0.132855f
C12639 VDAC_P.t14 VSS 0.10586f
C12640 VDAC_P.n1582 VSS 0.132855f
C12641 VDAC_P.t976 VSS 0.10586f
C12642 VDAC_P.n1583 VSS 0.132855f
C12643 VDAC_P.t15 VSS 0.10586f
C12644 VDAC_P.n1584 VSS 0.132855f
C12645 VDAC_P.t1496 VSS 0.10586f
C12646 VDAC_P.n1585 VSS 0.132855f
C12647 VDAC_P.t1690 VSS 0.10586f
C12648 VDAC_P.n1586 VSS 0.132855f
C12649 VDAC_P.t2100 VSS 0.10586f
C12650 VDAC_P.n1587 VSS 0.132855f
C12651 VDAC_P.t1486 VSS 0.10586f
C12652 VDAC_P.n1588 VSS 0.132855f
C12653 VDAC_P.t627 VSS 0.10586f
C12654 VDAC_P.n1589 VSS 0.132855f
C12655 VDAC_P.t2056 VSS 0.10586f
C12656 VDAC_P.n1590 VSS 0.132855f
C12657 VDAC_P.t1111 VSS 0.10586f
C12658 VDAC_P.n1591 VSS 0.132855f
C12659 VDAC_P.t799 VSS 0.10586f
C12660 VDAC_P.n1592 VSS 0.132855f
C12661 VDAC_P.t1754 VSS 0.10586f
C12662 VDAC_P.n1593 VSS 0.132855f
C12663 VDAC_P.t387 VSS 0.10586f
C12664 VDAC_P.n1594 VSS 0.132855f
C12665 VDAC_P.t218 VSS 0.10586f
C12666 VDAC_P.n1595 VSS 0.132855f
C12667 VDAC_P.t639 VSS 0.10586f
C12668 VDAC_P.n1596 VSS 0.132855f
C12669 VDAC_P.t1809 VSS 0.10586f
C12670 VDAC_P.n1597 VSS 0.132855f
C12671 VDAC_P.t307 VSS 0.10586f
C12672 VDAC_P.n1598 VSS 0.132855f
C12673 VDAC_P.t1599 VSS 0.10586f
C12674 VDAC_P.n1599 VSS 0.132855f
C12675 VDAC_P.t281 VSS 0.10586f
C12676 VDAC_P.n1600 VSS 0.132855f
C12677 VDAC_P.t1493 VSS 0.10586f
C12678 VDAC_P.n1601 VSS 0.132855f
C12679 VDAC_P.t1947 VSS 0.10586f
C12680 VDAC_P.n1602 VSS 0.132855f
C12681 VDAC_P.t1275 VSS 0.10586f
C12682 VDAC_P.n1603 VSS 0.132855f
C12683 VDAC_P.t1837 VSS 0.10586f
C12684 VDAC_P.n1604 VSS 0.132855f
C12685 VDAC_P.t1108 VSS 0.10586f
C12686 VDAC_P.n1605 VSS 0.132855f
C12687 VDAC_P.t1707 VSS 0.10586f
C12688 VDAC_P.n1606 VSS 0.132855f
C12689 VDAC_P.t140 VSS 0.10586f
C12690 VDAC_P.n1607 VSS 0.132855f
C12691 VDAC_P.t1186 VSS 0.10586f
C12692 VDAC_P.n1608 VSS 0.132855f
C12693 VDAC_P.t2055 VSS 0.10586f
C12694 VDAC_P.n1609 VSS 0.132855f
C12695 VDAC_P.t392 VSS 0.10586f
C12696 VDAC_P.n1610 VSS 0.132855f
C12697 VDAC_P.t262 VSS 0.10586f
C12698 VDAC_P.n1611 VSS 0.132855f
C12699 VDAC_P.t532 VSS 0.10586f
C12700 VDAC_P.n1612 VSS 0.132855f
C12701 VDAC_P.t1478 VSS 0.10586f
C12702 VDAC_P.n1613 VSS 0.132855f
C12703 VDAC_P.t1156 VSS 0.10586f
C12704 VDAC_P.n1614 VSS 0.132855f
C12705 VDAC_P.t638 VSS 0.10586f
C12706 VDAC_P.n1615 VSS 0.132855f
C12707 VDAC_P.t1103 VSS 0.10586f
C12708 VDAC_P.n1616 VSS 0.132855f
C12709 VDAC_P.t2040 VSS 0.10586f
C12710 VDAC_P.n1617 VSS 0.132855f
C12711 VDAC_P.t1962 VSS 0.10586f
C12712 VDAC_P.n1618 VSS 0.132855f
C12713 VDAC_P.t743 VSS 0.10586f
C12714 VDAC_P.n1619 VSS 0.132855f
C12715 VDAC_P.t1542 VSS 0.10586f
C12716 VDAC_P.n1620 VSS 0.132855f
C12717 VDAC_P.t1351 VSS 0.10586f
C12718 VDAC_P.n1621 VSS 0.132855f
C12719 VDAC_P.t1310 VSS 0.10586f
C12720 VDAC_P.n1622 VSS 0.132855f
C12721 VDAC_P.t1141 VSS 0.10586f
C12722 VDAC_P.n1623 VSS 0.132855f
C12723 VDAC_P.t237 VSS 0.10586f
C12724 VDAC_P.n1624 VSS 0.132855f
C12725 VDAC_P.t2022 VSS 0.10586f
C12726 VDAC_P.n1625 VSS 0.132855f
C12727 VDAC_P.t1489 VSS 0.10586f
C12728 VDAC_P.n1626 VSS 0.132855f
C12729 VDAC_P.t1037 VSS 0.10586f
C12730 VDAC_P.n1627 VSS 0.132855f
C12731 VDAC_P.t365 VSS 0.10586f
C12732 VDAC_P.n1628 VSS 0.12686f
C12733 VDAC_P.t881 VSS 0.10586f
C12734 VDAC_P.n1629 VSS 0.132855f
C12735 VDAC_P.t308 VSS 0.10586f
C12736 VDAC_P.n1630 VSS 0.132855f
C12737 VDAC_P.t1633 VSS 0.10586f
C12738 VDAC_P.n1631 VSS 0.132855f
C12739 VDAC_P.t2083 VSS 0.10586f
C12740 VDAC_P.n1632 VSS 0.132855f
C12741 VDAC_P.t1616 VSS 0.10586f
C12742 VDAC_P.n1633 VSS 0.132855f
C12743 VDAC_P.t1983 VSS 0.10586f
C12744 VDAC_P.n1634 VSS 0.132855f
C12745 VDAC_P.t168 VSS 0.10586f
C12746 VDAC_P.n1635 VSS 0.132855f
C12747 VDAC_P.t406 VSS 0.10586f
C12748 VDAC_P.n1636 VSS 0.132855f
C12749 VDAC_P.t372 VSS 0.10586f
C12750 VDAC_P.n1637 VSS 0.132855f
C12751 VDAC_P.t38 VSS 0.10586f
C12752 VDAC_P.n1638 VSS 0.132855f
C12753 VDAC_P.t1071 VSS 0.10586f
C12754 VDAC_P.n1639 VSS 0.132855f
C12755 VDAC_P.t1090 VSS 0.10586f
C12756 VDAC_P.n1640 VSS 0.132855f
C12757 VDAC_P.t2018 VSS 0.10586f
C12758 VDAC_P.n1641 VSS 0.132855f
C12759 VDAC_P.t59 VSS 0.10586f
C12760 VDAC_P.n1642 VSS 0.132855f
C12761 VDAC_P.t648 VSS 0.10586f
C12762 VDAC_P.n1643 VSS 0.132855f
C12763 VDAC_P.t250 VSS 0.10586f
C12764 VDAC_P.n1644 VSS 0.132855f
C12765 VDAC_P.t1668 VSS 0.10586f
C12766 VDAC_P.n1645 VSS 0.132855f
C12767 VDAC_P.t1358 VSS 0.10586f
C12768 VDAC_P.n1646 VSS 0.132855f
C12769 VDAC_P.t649 VSS 0.10586f
C12770 VDAC_P.n1647 VSS 0.132855f
C12771 VDAC_P.t590 VSS 0.10586f
C12772 VDAC_P.n1648 VSS 0.132855f
C12773 VDAC_P.t2070 VSS 0.10586f
C12774 VDAC_P.n1649 VSS 0.132855f
C12775 VDAC_P.t936 VSS 0.10586f
C12776 VDAC_P.n1650 VSS 0.132855f
C12777 VDAC_P.t486 VSS 0.10586f
C12778 VDAC_P.n1651 VSS 0.132855f
C12779 VDAC_P.t715 VSS 0.10586f
C12780 VDAC_P.n1652 VSS 0.132855f
C12781 VDAC_P.t1426 VSS 0.10586f
C12782 VDAC_P.n1653 VSS 0.132855f
C12783 VDAC_P.t187 VSS 0.10586f
C12784 VDAC_P.n1654 VSS 0.132855f
C12785 VDAC_P.t1755 VSS 0.10586f
C12786 VDAC_P.n1655 VSS 0.132855f
C12787 VDAC_P.t25 VSS 0.10586f
C12788 VDAC_P.n1656 VSS 0.132855f
C12789 VDAC_P.t231 VSS 0.10586f
C12790 VDAC_P.n1657 VSS 0.132855f
C12791 VDAC_P.t1922 VSS 0.10586f
C12792 VDAC_P.n1658 VSS 0.132855f
C12793 VDAC_P.t379 VSS 0.10586f
C12794 VDAC_P.n1659 VSS 0.132855f
C12795 VDAC_P.t2001 VSS 0.10586f
C12796 VDAC_P.n1660 VSS 0.132855f
C12797 VDAC_P.t1333 VSS 0.10586f
C12798 VDAC_P.n1661 VSS 0.132855f
C12799 VDAC_P.t1787 VSS 0.10586f
C12800 VDAC_P.n1662 VSS 0.132855f
C12801 VDAC_P.t684 VSS 0.10586f
C12802 VDAC_P.n1663 VSS 0.132855f
C12803 VDAC_P.t855 VSS 0.10586f
C12804 VDAC_P.n1664 VSS 0.132855f
C12805 VDAC_P.t450 VSS 0.10586f
C12806 VDAC_P.n1665 VSS 0.132855f
C12807 VDAC_P.t73 VSS 0.10586f
C12808 VDAC_P.n1666 VSS 0.132855f
C12809 VDAC_P.t2031 VSS 0.10586f
C12810 VDAC_P.n1667 VSS 0.132855f
C12811 VDAC_P.t688 VSS 0.10586f
C12812 VDAC_P.n1668 VSS 0.132855f
C12813 VDAC_P.t1895 VSS 0.10586f
C12814 VDAC_P.n1669 VSS 0.132855f
C12815 VDAC_P.t1240 VSS 0.10586f
C12816 VDAC_P.n1670 VSS 0.132855f
C12817 VDAC_P.t1574 VSS 0.10586f
C12818 VDAC_P.n1671 VSS 0.132855f
C12819 VDAC_P.t1420 VSS 0.10586f
C12820 VDAC_P.n1672 VSS 0.132855f
C12821 VDAC_P.t586 VSS 0.10586f
C12822 VDAC_P.n1673 VSS 0.132855f
C12823 VDAC_P.t595 VSS 0.10586f
C12824 VDAC_P.n1674 VSS 0.132855f
C12825 VDAC_P.t56 VSS 0.10586f
C12826 VDAC_P.n1675 VSS 0.132855f
C12827 VDAC_P.t1854 VSS 0.10586f
C12828 VDAC_P.n1676 VSS 0.132855f
C12829 VDAC_P.t696 VSS 0.10586f
C12830 VDAC_P.n1677 VSS 0.132855f
C12831 VDAC_P.t78 VSS 0.10586f
C12832 VDAC_P.n1678 VSS 0.132855f
C12833 VDAC_P.t345 VSS 0.10586f
C12834 VDAC_P.n1679 VSS 0.132855f
C12835 VDAC_P.t1414 VSS 0.10586f
C12836 VDAC_P.n1680 VSS 0.132855f
C12837 VDAC_P.t173 VSS 0.10586f
C12838 VDAC_P.n1681 VSS 0.132855f
C12839 VDAC_P.t433 VSS 0.10586f
C12840 VDAC_P.n1682 VSS 0.132855f
C12841 VDAC_P.t146 VSS 0.10586f
C12842 VDAC_P.n1683 VSS 0.132855f
C12843 VDAC_P.t1539 VSS 0.10586f
C12844 VDAC_P.n1684 VSS 0.132855f
C12845 VDAC_P.t858 VSS 0.10586f
C12846 VDAC_P.n1685 VSS 0.132855f
C12847 VDAC_P.t679 VSS 0.10586f
C12848 VDAC_P.n1686 VSS 0.132855f
C12849 VDAC_P.t57 VSS 0.10586f
C12850 VDAC_P.n1687 VSS 0.132855f
C12851 VDAC_P.t1225 VSS 0.10586f
C12852 VDAC_P.n1688 VSS 0.132855f
C12853 VDAC_P.t441 VSS 0.10586f
C12854 VDAC_P.n1689 VSS 0.132855f
C12855 VDAC_P.t1228 VSS 0.10586f
C12856 VDAC_P.n1690 VSS 0.132855f
C12857 VDAC_P.t1569 VSS 0.10586f
C12858 VDAC_P.n1691 VSS 0.12686f
C12859 VDAC_P.t1210 VSS 0.10586f
C12860 VDAC_P.n1692 VSS 0.132855f
C12861 VDAC_P.t1197 VSS 0.10586f
C12862 VDAC_P.n1693 VSS 0.132855f
C12863 VDAC_P.t1952 VSS 0.10586f
C12864 VDAC_P.n1694 VSS 0.132855f
C12865 VDAC_P.t978 VSS 0.10586f
C12866 VDAC_P.n1695 VSS 0.132855f
C12867 VDAC_P.t39 VSS 0.10586f
C12868 VDAC_P.n1696 VSS 0.132855f
C12869 VDAC_P.t866 VSS 0.10586f
C12870 VDAC_P.n1697 VSS 0.132855f
C12871 VDAC_P.t355 VSS 0.10586f
C12872 VDAC_P.n1698 VSS 0.132855f
C12873 VDAC_P.t1789 VSS 0.10586f
C12874 VDAC_P.n1699 VSS 0.132855f
C12875 VDAC_P.t329 VSS 0.10586f
C12876 VDAC_P.n1700 VSS 0.132855f
C12877 VDAC_P.t857 VSS 0.10586f
C12878 VDAC_P.n1701 VSS 0.132855f
C12879 VDAC_P.t1978 VSS 0.10586f
C12880 VDAC_P.n1702 VSS 0.132855f
C12881 VDAC_P.t1577 VSS 0.10586f
C12882 VDAC_P.n1703 VSS 0.132855f
C12883 VDAC_P.t1031 VSS 0.10586f
C12884 VDAC_P.n1704 VSS 0.132855f
C12885 VDAC_P.t1299 VSS 0.10586f
C12886 VDAC_P.n1705 VSS 0.132855f
C12887 VDAC_P.t1751 VSS 0.10586f
C12888 VDAC_P.n1706 VSS 0.132855f
C12889 VDAC_P.t1284 VSS 0.10586f
C12890 VDAC_P.n1707 VSS 0.132855f
C12891 VDAC_P.t1649 VSS 0.10586f
C12892 VDAC_P.n1708 VSS 0.132855f
C12893 VDAC_P.t1063 VSS 0.10586f
C12894 VDAC_P.n1709 VSS 0.132855f
C12895 VDAC_P.t1056 VSS 0.10586f
C12896 VDAC_P.n1710 VSS 0.132855f
C12897 VDAC_P.t1997 VSS 0.10586f
C12898 VDAC_P.n1711 VSS 0.132855f
C12899 VDAC_P.t176 VSS 0.10586f
C12900 VDAC_P.n1712 VSS 0.132855f
C12901 VDAC_P.t957 VSS 0.10586f
C12902 VDAC_P.n1713 VSS 0.132855f
C12903 VDAC_P.t1524 VSS 0.10586f
C12904 VDAC_P.n1714 VSS 0.132855f
C12905 VDAC_P.t1338 VSS 0.10586f
C12906 VDAC_P.n1715 VSS 0.132855f
C12907 VDAC_P.t587 VSS 0.10586f
C12908 VDAC_P.n1716 VSS 0.132855f
C12909 VDAC_P.t1118 VSS 0.10586f
C12910 VDAC_P.n1717 VSS 0.132855f
C12911 VDAC_P.t154 VSS 0.10586f
C12912 VDAC_P.n1718 VSS 0.132855f
C12913 VDAC_P.t1336 VSS 0.10586f
C12914 VDAC_P.n1719 VSS 0.132855f
C12915 VDAC_P.t478 VSS 0.10586f
C12916 VDAC_P.n1720 VSS 0.132855f
C12917 VDAC_P.t1812 VSS 0.10586f
C12918 VDAC_P.n1721 VSS 0.132855f
C12919 VDAC_P.t1394 VSS 0.10586f
C12920 VDAC_P.n1722 VSS 0.132855f
C12921 VDAC_P.t1283 VSS 0.10586f
C12922 VDAC_P.n1723 VSS 0.132855f
C12923 VDAC_P.t46 VSS 0.10586f
C12924 VDAC_P.n1724 VSS 0.132855f
C12925 VDAC_P.t1066 VSS 0.10586f
C12926 VDAC_P.n1725 VSS 0.132855f
C12927 VDAC_P.t1527 VSS 0.10586f
C12928 VDAC_P.n1726 VSS 0.132855f
C12929 VDAC_P.t494 VSS 0.10586f
C12930 VDAC_P.n1727 VSS 0.132855f
C12931 VDAC_P.t1417 VSS 0.10586f
C12932 VDAC_P.n1728 VSS 0.132855f
C12933 VDAC_P.t118 VSS 0.10586f
C12934 VDAC_P.n1729 VSS 0.132855f
C12935 VDAC_P.t673 VSS 0.10586f
C12936 VDAC_P.n1730 VSS 0.132855f
C12937 VDAC_P.t1767 VSS 0.10586f
C12938 VDAC_P.n1731 VSS 0.132855f
C12939 VDAC_P.t1187 VSS 0.10586f
C12940 VDAC_P.n1732 VSS 0.132855f
C12941 VDAC_P.t1745 VSS 0.10586f
C12942 VDAC_P.n1733 VSS 0.132855f
C12943 VDAC_P.t1404 VSS 0.10586f
C12944 VDAC_P.n1734 VSS 0.132855f
C12945 VDAC_P.t1535 VSS 0.10586f
C12946 VDAC_P.n1735 VSS 0.132855f
C12947 VDAC_P.t1993 VSS 0.10586f
C12948 VDAC_P.n1736 VSS 0.132855f
C12949 VDAC_P.t1656 VSS 0.10586f
C12950 VDAC_P.n1737 VSS 0.132855f
C12951 VDAC_P.t953 VSS 0.10586f
C12952 VDAC_P.n1738 VSS 0.132855f
C12953 VDAC_P.t756 VSS 0.10586f
C12954 VDAC_P.n1739 VSS 0.132855f
C12955 VDAC_P.t137 VSS 0.10586f
C12956 VDAC_P.n1740 VSS 0.132855f
C12957 VDAC_P.t588 VSS 0.10586f
C12958 VDAC_P.n1741 VSS 0.132855f
C12959 VDAC_P.t1106 VSS 0.10586f
C12960 VDAC_P.n1742 VSS 0.132855f
C12961 VDAC_P.t1077 VSS 0.10586f
C12962 VDAC_P.n1743 VSS 0.132855f
C12963 VDAC_P.t896 VSS 0.10586f
C12964 VDAC_P.n1744 VSS 0.132855f
C12965 VDAC_P.t1818 VSS 0.10586f
C12966 VDAC_P.n1745 VSS 0.132855f
C12967 VDAC_P.t1780 VSS 0.10586f
C12968 VDAC_P.n1746 VSS 0.132855f
C12969 VDAC_P.t1602 VSS 0.10586f
C12970 VDAC_P.n1747 VSS 0.132855f
C12971 VDAC_P.t844 VSS 0.10586f
C12972 VDAC_P.n1748 VSS 0.132855f
C12973 VDAC_P.t1170 VSS 0.10586f
C12974 VDAC_P.n1749 VSS 0.132855f
C12975 VDAC_P.t315 VSS 0.10586f
C12976 VDAC_P.n1750 VSS 0.132855f
C12977 VDAC_P.t1880 VSS 0.10586f
C12978 VDAC_P.n1751 VSS 0.132855f
C12979 VDAC_P.t1886 VSS 0.10586f
C12980 VDAC_P.n1752 VSS 0.132855f
C12981 VDAC_P.t1525 VSS 0.10586f
C12982 VDAC_P.n1753 VSS 0.132855f
C12983 VDAC_P.t1658 VSS 0.10586f
C12984 VDAC_P.n1754 VSS 0.12686f
C12985 VDAC_P.t199 VSS 0.10586f
C12986 VDAC_P.n1755 VSS 0.132855f
C12987 VDAC_P.t1961 VSS 0.10586f
C12988 VDAC_P.n1756 VSS 0.132855f
C12989 VDAC_P.t1295 VSS 0.10586f
C12990 VDAC_P.n1757 VSS 0.132855f
C12991 VDAC_P.t243 VSS 0.10586f
C12992 VDAC_P.n1758 VSS 0.132855f
C12993 VDAC_P.t1532 VSS 0.10586f
C12994 VDAC_P.n1759 VSS 0.132855f
C12995 VDAC_P.t837 VSS 0.10586f
C12996 VDAC_P.n1760 VSS 0.132855f
C12997 VDAC_P.t2095 VSS 0.10586f
C12998 VDAC_P.n1761 VSS 0.132855f
C12999 VDAC_P.t848 VSS 0.10586f
C13000 VDAC_P.n1762 VSS 0.132855f
C13001 VDAC_P.t1995 VSS 0.10586f
C13002 VDAC_P.n1763 VSS 0.132855f
C13003 VDAC_P.t608 VSS 0.10586f
C13004 VDAC_P.n1764 VSS 0.132855f
C13005 VDAC_P.t247 VSS 0.10586f
C13006 VDAC_P.n1765 VSS 0.132855f
C13007 VDAC_P.t212 VSS 0.10586f
C13008 VDAC_P.n1766 VSS 0.132855f
C13009 VDAC_P.t678 VSS 0.10586f
C13010 VDAC_P.n1767 VSS 0.132855f
C13011 VDAC_P.t759 VSS 0.10586f
C13012 VDAC_P.n1768 VSS 0.132855f
C13013 VDAC_P.t1943 VSS 0.10586f
C13014 VDAC_P.n1769 VSS 0.132855f
C13015 VDAC_P.t1432 VSS 0.10586f
C13016 VDAC_P.n1770 VSS 0.132855f
C13017 VDAC_P.t1833 VSS 0.10586f
C13018 VDAC_P.n1771 VSS 0.132855f
C13019 VDAC_P.t1068 VSS 0.10586f
C13020 VDAC_P.n1772 VSS 0.132855f
C13021 VDAC_P.t1446 VSS 0.10586f
C13022 VDAC_P.n1773 VSS 0.132855f
C13023 VDAC_P.t28 VSS 0.10586f
C13024 VDAC_P.n1774 VSS 0.132855f
C13025 VDAC_P.t2000 VSS 0.10586f
C13026 VDAC_P.n1775 VSS 0.132855f
C13027 VDAC_P.t2135 VSS 0.10586f
C13028 VDAC_P.n1776 VSS 0.132855f
C13029 VDAC_P.t1560 VSS 0.10586f
C13030 VDAC_P.n1777 VSS 0.132855f
C13031 VDAC_P.t1726 VSS 0.10586f
C13032 VDAC_P.n1778 VSS 0.132855f
C13033 VDAC_P.t1348 VSS 0.10586f
C13034 VDAC_P.n1779 VSS 0.132855f
C13035 VDAC_P.t214 VSS 0.10586f
C13036 VDAC_P.n1780 VSS 0.132855f
C13037 VDAC_P.t633 VSS 0.10586f
C13038 VDAC_P.n1781 VSS 0.132855f
C13039 VDAC_P.t1072 VSS 0.10586f
C13040 VDAC_P.n1782 VSS 0.132855f
C13041 VDAC_P.t1127 VSS 0.10586f
C13042 VDAC_P.n1783 VSS 0.132855f
C13043 VDAC_P.t1704 VSS 0.10586f
C13044 VDAC_P.n1784 VSS 0.132855f
C13045 VDAC_P.t902 VSS 0.10586f
C13046 VDAC_P.n1785 VSS 0.132855f
C13047 VDAC_P.t1475 VSS 0.10586f
C13048 VDAC_P.n1786 VSS 0.132855f
C13049 VDAC_P.t798 VSS 0.10586f
C13050 VDAC_P.n1787 VSS 0.132855f
C13051 VDAC_P.t645 VSS 0.10586f
C13052 VDAC_P.n1788 VSS 0.132855f
C13053 VDAC_P.t1715 VSS 0.10586f
C13054 VDAC_P.n1789 VSS 0.132855f
C13055 VDAC_P.t593 VSS 0.10586f
C13056 VDAC_P.n1790 VSS 0.132855f
C13057 VDAC_P.t1613 VSS 0.10586f
C13058 VDAC_P.n1791 VSS 0.132855f
C13059 VDAC_P.t934 VSS 0.10586f
C13060 VDAC_P.n1792 VSS 0.132855f
C13061 VDAC_P.t767 VSS 0.10586f
C13062 VDAC_P.n1793 VSS 0.132855f
C13063 VDAC_P.t1957 VSS 0.10586f
C13064 VDAC_P.n1794 VSS 0.132855f
C13065 VDAC_P.t1373 VSS 0.10586f
C13066 VDAC_P.n1795 VSS 0.132855f
C13067 VDAC_P.t147 VSS 0.10586f
C13068 VDAC_P.n1796 VSS 0.132855f
C13069 VDAC_P.t1924 VSS 0.10586f
C13070 VDAC_P.n1797 VSS 0.132855f
C13071 VDAC_P.t1721 VSS 0.10586f
C13072 VDAC_P.n1798 VSS 0.132855f
C13073 VDAC_P.t1078 VSS 0.10586f
C13074 VDAC_P.n1799 VSS 0.132855f
C13075 VDAC_P.t622 VSS 0.10586f
C13076 VDAC_P.n1800 VSS 0.132855f
C13077 VDAC_P.t2069 VSS 0.10586f
C13078 VDAC_P.n1801 VSS 0.132855f
C13079 VDAC_P.t784 VSS 0.10586f
C13080 VDAC_P.n1802 VSS 0.132855f
C13081 VDAC_P.t149 VSS 0.10586f
C13082 VDAC_P.n1803 VSS 0.132855f
C13083 VDAC_P.t160 VSS 0.10586f
C13084 VDAC_P.n1804 VSS 0.132855f
C13085 VDAC_P.t1506 VSS 0.10586f
C13086 VDAC_P.n1805 VSS 0.132855f
C13087 VDAC_P.t1268 VSS 0.10586f
C13088 VDAC_P.n1806 VSS 0.132855f
C13089 VDAC_P.t1274 VSS 0.10586f
C13090 VDAC_P.n1807 VSS 0.132855f
C13091 VDAC_P.t1121 VSS 0.10586f
C13092 VDAC_P.n1808 VSS 0.132855f
C13093 VDAC_P.t856 VSS 0.10586f
C13094 VDAC_P.n1809 VSS 0.132855f
C13095 VDAC_P.t1006 VSS 0.10586f
C13096 VDAC_P.n1810 VSS 0.132855f
C13097 VDAC_P.t616 VSS 0.10586f
C13098 VDAC_P.n1811 VSS 0.132855f
C13099 VDAC_P.t794 VSS 0.10586f
C13100 VDAC_P.n1812 VSS 0.132855f
C13101 VDAC_P.t195 VSS 0.10586f
C13102 VDAC_P.n1813 VSS 0.132855f
C13103 VDAC_P.t682 VSS 0.10586f
C13104 VDAC_P.n1814 VSS 0.132855f
C13105 VDAC_P.t1153 VSS 0.10586f
C13106 VDAC_P.n1815 VSS 0.132855f
C13107 VDAC_P.t1711 VSS 0.10586f
C13108 VDAC_P.n1816 VSS 0.132855f
C13109 VDAC_P.t2042 VSS 0.10586f
C13110 VDAC_P.n1817 VSS 0.12686f
C13111 VDAC_P.t18 VSS 0.10586f
C13112 VDAC_P.n1818 VSS 0.132855f
C13113 VDAC_P.t1194 VSS 0.10586f
C13114 VDAC_P.n1819 VSS 0.132855f
C13115 VDAC_P.t2059 VSS 0.10586f
C13116 VDAC_P.n1820 VSS 0.132855f
C13117 VDAC_P.t760 VSS 0.10586f
C13118 VDAC_P.n1821 VSS 0.132855f
C13119 VDAC_P.t1686 VSS 0.10586f
C13120 VDAC_P.n1822 VSS 0.132855f
C13121 VDAC_P.t36 VSS 0.10586f
C13122 VDAC_P.n1823 VSS 0.132855f
C13123 VDAC_P.t1482 VSS 0.10586f
C13124 VDAC_P.n1824 VSS 0.132855f
C13125 VDAC_P.t1223 VSS 0.10586f
C13126 VDAC_P.n1825 VSS 0.132855f
C13127 VDAC_P.t1254 VSS 0.10586f
C13128 VDAC_P.n1826 VSS 0.132855f
C13129 VDAC_P.t163 VSS 0.10586f
C13130 VDAC_P.n1827 VSS 0.132855f
C13131 VDAC_P.t128 VSS 0.10586f
C13132 VDAC_P.n1828 VSS 0.132855f
C13133 VDAC_P.t1966 VSS 0.10586f
C13134 VDAC_P.n1829 VSS 0.132855f
C13135 VDAC_P.t1459 VSS 0.10586f
C13136 VDAC_P.n1830 VSS 0.132855f
C13137 VDAC_P.t1681 VSS 0.10586f
C13138 VDAC_P.n1831 VSS 0.132855f
C13139 VDAC_P.t1367 VSS 0.10586f
C13140 VDAC_P.n1832 VSS 0.132855f
C13141 VDAC_P.t62 VSS 0.10586f
C13142 VDAC_P.n1833 VSS 0.132855f
C13143 VDAC_P.t2029 VSS 0.10586f
C13144 VDAC_P.n1834 VSS 0.132855f
C13145 VDAC_P.t1328 VSS 0.10586f
C13146 VDAC_P.n1835 VSS 0.132855f
C13147 VDAC_P.t1826 VSS 0.10586f
C13148 VDAC_P.n1836 VSS 0.132855f
C13149 VDAC_P.t916 VSS 0.10586f
C13150 VDAC_P.n1837 VSS 0.132855f
C13151 VDAC_P.t710 VSS 0.10586f
C13152 VDAC_P.n1838 VSS 0.132855f
C13153 VDAC_P.t1740 VSS 0.10586f
C13154 VDAC_P.n1839 VSS 0.132855f
C13155 VDAC_P.t1178 VSS 0.10586f
C13156 VDAC_P.n1840 VSS 0.132855f
C13157 VDAC_P.t2102 VSS 0.10586f
C13158 VDAC_P.n1841 VSS 0.132855f
C13159 VDAC_P.t1464 VSS 0.10586f
C13160 VDAC_P.n1842 VSS 0.132855f
C13161 VDAC_P.t1890 VSS 0.10586f
C13162 VDAC_P.n1843 VSS 0.132855f
C13163 VDAC_P.t375 VSS 0.10586f
C13164 VDAC_P.n1844 VSS 0.132855f
C13165 VDAC_P.t746 VSS 0.10586f
C13166 VDAC_P.n1845 VSS 0.132855f
C13167 VDAC_P.t1317 VSS 0.10586f
C13168 VDAC_P.n1846 VSS 0.132855f
C13169 VDAC_P.t1242 VSS 0.10586f
C13170 VDAC_P.n1847 VSS 0.132855f
C13171 VDAC_P.t295 VSS 0.10586f
C13172 VDAC_P.n1848 VSS 0.132855f
C13173 VDAC_P.t1667 VSS 0.10586f
C13174 VDAC_P.n1849 VSS 0.132855f
C13175 VDAC_P.t990 VSS 0.10586f
C13176 VDAC_P.n1850 VSS 0.132855f
C13177 VDAC_P.t1451 VSS 0.10586f
C13178 VDAC_P.n1851 VSS 0.132855f
C13179 VDAC_P.t497 VSS 0.10586f
C13180 VDAC_P.n1852 VSS 0.132855f
C13181 VDAC_P.t1343 VSS 0.10586f
C13182 VDAC_P.n1853 VSS 0.132855f
C13183 VDAC_P.t471 VSS 0.10586f
C13184 VDAC_P.n1854 VSS 0.132855f
C13185 VDAC_P.t97 VSS 0.10586f
C13186 VDAC_P.n1855 VSS 0.132855f
C13187 VDAC_P.t861 VSS 0.10586f
C13188 VDAC_P.n1856 VSS 0.132855f
C13189 VDAC_P.t220 VSS 0.10586f
C13190 VDAC_P.n1857 VSS 0.132855f
C13191 VDAC_P.t1567 VSS 0.10586f
C13192 VDAC_P.n1858 VSS 0.132855f
C13193 VDAC_P.t2123 VSS 0.10586f
C13194 VDAC_P.n1859 VSS 0.132855f
C13195 VDAC_P.t1760 VSS 0.10586f
C13196 VDAC_P.n1860 VSS 0.132855f
C13197 VDAC_P.t1913 VSS 0.10586f
C13198 VDAC_P.n1861 VSS 0.132855f
C13199 VDAC_P.t900 VSS 0.10586f
C13200 VDAC_P.n1862 VSS 0.132855f
C13201 VDAC_P.t814 VSS 0.10586f
C13202 VDAC_P.n1863 VSS 0.132855f
C13203 VDAC_P.t1644 VSS 0.10586f
C13204 VDAC_P.n1864 VSS 0.132855f
C13205 VDAC_P.t598 VSS 0.10586f
C13206 VDAC_P.n1865 VSS 0.132855f
C13207 VDAC_P.t604 VSS 0.10586f
C13208 VDAC_P.n1866 VSS 0.132855f
C13209 VDAC_P.t952 VSS 0.10586f
C13210 VDAC_P.n1867 VSS 0.132855f
C13211 VDAC_P.t1882 VSS 0.10586f
C13212 VDAC_P.n1868 VSS 0.132855f
C13213 VDAC_P.t728 VSS 0.10586f
C13214 VDAC_P.n1869 VSS 0.132855f
C13215 VDAC_P.t842 VSS 0.10586f
C13216 VDAC_P.n1870 VSS 0.132855f
C13217 VDAC_P.t1313 VSS 0.10586f
C13218 VDAC_P.n1871 VSS 0.132855f
C13219 VDAC_P.t330 VSS 0.10586f
C13220 VDAC_P.n1872 VSS 0.132855f
C13221 VDAC_P.t617 VSS 0.10586f
C13222 VDAC_P.n1873 VSS 0.132855f
C13223 VDAC_P.t520 VSS 0.10586f
C13224 VDAC_P.n1874 VSS 0.132855f
C13225 VDAC_P.t986 VSS 0.10586f
C13226 VDAC_P.n1875 VSS 0.132855f
C13227 VDAC_P.t793 VSS 0.10586f
C13228 VDAC_P.n1876 VSS 0.132855f
C13229 VDAC_P.t134 VSS 0.10586f
C13230 VDAC_P.n1877 VSS 0.132855f
C13231 VDAC_P.t1341 VSS 0.10586f
C13232 VDAC_P.n1878 VSS 0.132855f
C13233 VDAC_P.t145 VSS 0.10586f
C13234 VDAC_P.n1879 VSS 0.132855f
C13235 VDAC_P.t1237 VSS 0.10586f
C13236 VDAC_P.n1880 VSS 0.12686f
C13237 VDAC_P.t542 VSS 0.10586f
C13238 VDAC_P.n1881 VSS 0.132855f
C13239 VDAC_P.t829 VSS 0.10586f
C13240 VDAC_P.n1882 VSS 0.132855f
C13241 VDAC_P.t1878 VSS 0.10586f
C13242 VDAC_P.n1883 VSS 0.132855f
C13243 VDAC_P.t373 VSS 0.10586f
C13244 VDAC_P.n1884 VSS 0.132855f
C13245 VDAC_P.t1865 VSS 0.10586f
C13246 VDAC_P.n1885 VSS 0.132855f
C13247 VDAC_P.t669 VSS 0.10586f
C13248 VDAC_P.n1886 VSS 0.132855f
C13249 VDAC_P.t895 VSS 0.10586f
C13250 VDAC_P.n1887 VSS 0.132855f
C13251 VDAC_P.t1980 VSS 0.10586f
C13252 VDAC_P.n1888 VSS 0.132855f
C13253 VDAC_P.t1659 VSS 0.10586f
C13254 VDAC_P.n1889 VSS 0.132855f
C13255 VDAC_P.t549 VSS 0.10586f
C13256 VDAC_P.n1890 VSS 0.132855f
C13257 VDAC_P.t1443 VSS 0.10586f
C13258 VDAC_P.n1891 VSS 0.132855f
C13259 VDAC_P.t2009 VSS 0.10586f
C13260 VDAC_P.n1892 VSS 0.132855f
C13261 VDAC_P.t640 VSS 0.10586f
C13262 VDAC_P.n1893 VSS 0.132855f
C13263 VDAC_P.t958 VSS 0.10586f
C13264 VDAC_P.n1894 VSS 0.132855f
C13265 VDAC_P.t721 VSS 0.10586f
C13266 VDAC_P.n1895 VSS 0.132855f
C13267 VDAC_P.t1985 VSS 0.10586f
C13268 VDAC_P.n1896 VSS 0.132855f
C13269 VDAC_P.t1315 VSS 0.10586f
C13270 VDAC_P.n1897 VSS 0.132855f
C13271 VDAC_P.t1765 VSS 0.10586f
C13272 VDAC_P.n1898 VSS 0.132855f
C13273 VDAC_P.t1412 VSS 0.10586f
C13274 VDAC_P.n1899 VSS 0.132855f
C13275 VDAC_P.t437 VSS 0.10586f
C13276 VDAC_P.n1900 VSS 0.132855f
C13277 VDAC_P.t1073 VSS 0.10586f
C13278 VDAC_P.n1901 VSS 0.132855f
C13279 VDAC_P.t411 VSS 0.10586f
C13280 VDAC_P.n1902 VSS 0.132855f
C13281 VDAC_P.t2013 VSS 0.10586f
C13282 VDAC_P.n1903 VSS 0.132855f
C13283 VDAC_P.t184 VSS 0.10586f
C13284 VDAC_P.n1904 VSS 0.132855f
C13285 VDAC_P.t913 VSS 0.10586f
C13286 VDAC_P.n1905 VSS 0.132855f
C13287 VDAC_P.t852 VSS 0.10586f
C13288 VDAC_P.n1906 VSS 0.132855f
C13289 VDAC_P.t1362 VSS 0.10586f
C13290 VDAC_P.n1907 VSS 0.132855f
C13291 VDAC_P.t860 VSS 0.10586f
C13292 VDAC_P.n1908 VSS 0.132855f
C13293 VDAC_P.t1154 VSS 0.10586f
C13294 VDAC_P.n1909 VSS 0.132855f
C13295 VDAC_P.t2041 VSS 0.10586f
C13296 VDAC_P.n1910 VSS 0.132855f
C13297 VDAC_P.t712 VSS 0.10586f
C13298 VDAC_P.n1911 VSS 0.132855f
C13299 VDAC_P.t1862 VSS 0.10586f
C13300 VDAC_P.n1912 VSS 0.132855f
C13301 VDAC_P.t964 VSS 0.10586f
C13302 VDAC_P.n1913 VSS 0.132855f
C13303 VDAC_P.t1430 VSS 0.10586f
C13304 VDAC_P.n1914 VSS 0.132855f
C13305 VDAC_P.t1195 VSS 0.10586f
C13306 VDAC_P.n1915 VSS 0.132855f
C13307 VDAC_P.t1206 VSS 0.10586f
C13308 VDAC_P.n1916 VSS 0.132855f
C13309 VDAC_P.t29 VSS 0.10586f
C13310 VDAC_P.n1917 VSS 0.132855f
C13311 VDAC_P.t776 VSS 0.10586f
C13312 VDAC_P.n1918 VSS 0.132855f
C13313 VDAC_P.t502 VSS 0.10586f
C13314 VDAC_P.n1919 VSS 0.132855f
C13315 VDAC_P.t1433 VSS 0.10586f
C13316 VDAC_P.n1920 VSS 0.132855f
C13317 VDAC_P.t434 VSS 0.10586f
C13318 VDAC_P.n1921 VSS 0.132855f
C13319 VDAC_P.t717 VSS 0.10586f
C13320 VDAC_P.n1922 VSS 0.132855f
C13321 VDAC_P.t1863 VSS 0.10586f
C13322 VDAC_P.n1923 VSS 0.132855f
C13323 VDAC_P.t1203 VSS 0.10586f
C13324 VDAC_P.n1924 VSS 0.132855f
C13325 VDAC_P.t1661 VSS 0.10586f
C13326 VDAC_P.n1925 VSS 0.132855f
C13327 VDAC_P.t1916 VSS 0.10586f
C13328 VDAC_P.n1926 VSS 0.132855f
C13329 VDAC_P.t791 VSS 0.10586f
C13330 VDAC_P.n1927 VSS 0.132855f
C13331 VDAC_P.t1019 VSS 0.10586f
C13332 VDAC_P.n1928 VSS 0.132855f
C13333 VDAC_P.t381 VSS 0.10586f
C13334 VDAC_P.n1929 VSS 0.132855f
C13335 VDAC_P.t495 VSS 0.10586f
C13336 VDAC_P.n1930 VSS 0.132855f
C13337 VDAC_P.t228 VSS 0.10586f
C13338 VDAC_P.n1931 VSS 0.132855f
C13339 VDAC_P.t469 VSS 0.10586f
C13340 VDAC_P.n1932 VSS 0.132855f
C13341 VDAC_P.t204 VSS 0.10586f
C13342 VDAC_P.n1933 VSS 0.132855f
C13343 VDAC_P.t1146 VSS 0.10586f
C13344 VDAC_P.n1934 VSS 0.132855f
C13345 VDAC_P.t531 VSS 0.10586f
C13346 VDAC_P.n1935 VSS 0.132855f
C13347 VDAC_P.t1824 VSS 0.10586f
C13348 VDAC_P.n1936 VSS 0.132855f
C13349 VDAC_P.t1925 VSS 0.10586f
C13350 VDAC_P.n1937 VSS 0.132855f
C13351 VDAC_P.t1876 VSS 0.10586f
C13352 VDAC_P.n1938 VSS 0.132855f
C13353 VDAC_P.t1630 VSS 0.10586f
C13354 VDAC_P.n1939 VSS 0.132855f
C13355 VDAC_P.t1900 VSS 0.10586f
C13356 VDAC_P.n1940 VSS 0.132855f
C13357 VDAC_P.t1202 VSS 0.10586f
C13358 VDAC_P.n1941 VSS 0.132855f
C13359 VDAC_P.t1189 VSS 0.10586f
C13360 VDAC_P.n1942 VSS 0.132855f
C13361 VDAC_P.t1928 VSS 0.10586f
C13362 VDAC_P.n1943 VSS 0.12686f
C13363 VDAC_P.t1918 VSS 0.10586f
C13364 VDAC_P.n1944 VSS 0.142819f
C13365 VDAC_P.t41 VSS 0.10586f
C13366 VDAC_P.n1945 VSS 0.142819f
C13367 VDAC_P.t765 VSS 0.10586f
C13368 VDAC_P.n1946 VSS 0.142819f
C13369 VDAC_P.t671 VSS 0.10586f
C13370 VDAC_P.n1947 VSS 0.142819f
C13371 VDAC_P.t153 VSS 0.10586f
C13372 VDAC_P.n1948 VSS 0.142819f
C13373 VDAC_P.t479 VSS 0.10586f
C13374 VDAC_P.n1949 VSS 0.142819f
C13375 VDAC_P.t1632 VSS 0.10586f
C13376 VDAC_P.n1950 VSS 0.142819f
C13377 VDAC_P.t1652 VSS 0.10586f
C13378 VDAC_P.n1951 VSS 0.142819f
C13379 VDAC_P.t16 VSS 0.10586f
C13380 VDAC_P.n1952 VSS 0.142819f
C13381 VDAC_P.t770 VSS 0.10586f
C13382 VDAC_P.n1953 VSS 0.142819f
C13383 VDAC_P.t570 VSS 0.10586f
C13384 VDAC_P.n1954 VSS 0.142819f
C13385 VDAC_P.t663 VSS 0.10586f
C13386 VDAC_P.n1955 VSS 0.142819f
C13387 VDAC_P.t567 VSS 0.10586f
C13388 VDAC_P.n1956 VSS 0.142819f
C13389 VDAC_P.t1794 VSS 0.10586f
C13390 VDAC_P.n1957 VSS 0.142819f
C13391 VDAC_P.t831 VSS 0.10586f
C13392 VDAC_P.n1958 VSS 0.142819f
C13393 VDAC_P.t1439 VSS 0.10586f
C13394 VDAC_P.n1959 VSS 0.142819f
C13395 VDAC_P.t1669 VSS 0.10586f
C13396 VDAC_P.n1960 VSS 0.142819f
C13397 VDAC_P.t753 VSS 0.10586f
C13398 VDAC_P.n1961 VSS 0.142819f
C13399 VDAC_P.t1287 VSS 0.10586f
C13400 VDAC_P.n1962 VSS 0.142819f
C13401 VDAC_P.t1990 VSS 0.10586f
C13402 VDAC_P.n1963 VSS 0.142819f
C13403 VDAC_P.t1207 VSS 0.10586f
C13404 VDAC_P.n1964 VSS 0.142819f
C13405 VDAC_P.t1976 VSS 0.10586f
C13406 VDAC_P.n1965 VSS 0.142819f
C13407 VDAC_P.t1382 VSS 0.10586f
C13408 VDAC_P.n1966 VSS 0.142819f
C13409 VDAC_P.t1770 VSS 0.10586f
C13410 VDAC_P.n1967 VSS 0.142819f
C13411 VDAC_P.t100 VSS 0.10586f
C13412 VDAC_P.n1968 VSS 0.142819f
C13413 VDAC_P.t112 VSS 0.10586f
C13414 VDAC_P.n1969 VSS 0.142819f
C13415 VDAC_P.t1779 VSS 0.10586f
C13416 VDAC_P.n1970 VSS 0.142819f
C13417 VDAC_P.t999 VSS 0.10586f
C13418 VDAC_P.n1971 VSS 0.142819f
C13419 VDAC_P.t924 VSS 0.10586f
C13420 VDAC_P.n1972 VSS 0.137296f
C13421 VDAC_P.t737 VSS 0.10586f
C13422 VDAC_P.n1973 VSS 0.126469f
C13423 VDAC_P.t1938 VSS 0.10586f
C13424 VDAC_P.n1974 VSS 0.132855f
C13425 VDAC_P.t79 VSS 0.10586f
C13426 VDAC_P.n1975 VSS 0.132855f
C13427 VDAC_P.t1091 VSS 0.10586f
C13428 VDAC_P.n1976 VSS 0.132855f
C13429 VDAC_P.t1226 VSS 0.10586f
C13430 VDAC_P.n1977 VSS 0.132855f
C13431 VDAC_P.t1311 VSS 0.10586f
C13432 VDAC_P.n1978 VSS 0.132855f
C13433 VDAC_P.t382 VSS 0.10586f
C13434 VDAC_P.n1979 VSS 0.132855f
C13435 VDAC_P.t996 VSS 0.10586f
C13436 VDAC_P.n1980 VSS 0.132855f
C13437 VDAC_P.t954 VSS 0.10586f
C13438 VDAC_P.n1981 VSS 0.132855f
C13439 VDAC_P.t1424 VSS 0.10586f
C13440 VDAC_P.n1982 VSS 0.132855f
C13441 VDAC_P.t2090 VSS 0.10586f
C13442 VDAC_P.n1983 VSS 0.132855f
C13443 VDAC_P.t1166 VSS 0.10586f
C13444 VDAC_P.n1984 VSS 0.132855f
C13445 VDAC_P.t812 VSS 0.10586f
C13446 VDAC_P.n1985 VSS 0.132855f
C13447 VDAC_P.t702 VSS 0.10586f
C13448 VDAC_P.n1986 VSS 0.132855f
C13449 VDAC_P.t452 VSS 0.10586f
C13450 VDAC_P.n1987 VSS 0.132855f
C13451 VDAC_P.t1909 VSS 0.10586f
C13452 VDAC_P.n1988 VSS 0.132855f
C13453 VDAC_P.t664 VSS 0.10586f
C13454 VDAC_P.n1989 VSS 0.132855f
C13455 VDAC_P.t1023 VSS 0.10586f
C13456 VDAC_P.n1990 VSS 0.132855f
C13457 VDAC_P.t1102 VSS 0.10586f
C13458 VDAC_P.n1991 VSS 0.132855f
C13459 VDAC_P.t1075 VSS 0.10586f
C13460 VDAC_P.n1992 VSS 0.132855f
C13461 VDAC_P.t439 VSS 0.10586f
C13462 VDAC_P.n1993 VSS 0.132855f
C13463 VDAC_P.t1460 VSS 0.10586f
C13464 VDAC_P.n1994 VSS 0.132855f
C13465 VDAC_P.t1875 VSS 0.10586f
C13466 VDAC_P.n1995 VSS 0.132855f
C13467 VDAC_P.t675 VSS 0.10586f
C13468 VDAC_P.n1996 VSS 0.132855f
C13469 VDAC_P.t1903 VSS 0.10586f
C13470 VDAC_P.n1997 VSS 0.132855f
C13471 VDAC_P.t1449 VSS 0.10586f
C13472 VDAC_P.n1998 VSS 0.132855f
C13473 VDAC_P.t454 VSS 0.10586f
C13474 VDAC_P.n1999 VSS 0.132855f
C13475 VDAC_P.t795 VSS 0.10586f
C13476 VDAC_P.n2000 VSS 0.132855f
C13477 VDAC_P.t561 VSS 0.10586f
C13478 VDAC_P.n2001 VSS 0.132855f
C13479 VDAC_P.t847 VSS 0.10586f
C13480 VDAC_P.n2002 VSS 0.132855f
C13481 VDAC_P.t619 VSS 0.10586f
C13482 VDAC_P.n2003 VSS 0.132855f
C13483 VDAC_P.t386 VSS 0.10586f
C13484 VDAC_P.n2004 VSS 0.132855f
C13485 VDAC_P.t1413 VSS 0.10586f
C13486 VDAC_P.n2005 VSS 0.132855f
C13487 VDAC_P.t846 VSS 0.10586f
C13488 VDAC_P.n2006 VSS 0.132855f
C13489 VDAC_P.t1456 VSS 0.10586f
C13490 VDAC_P.n2007 VSS 0.132855f
C13491 VDAC_P.t2098 VSS 0.10586f
C13492 VDAC_P.n2008 VSS 0.132855f
C13493 VDAC_P.t1896 VSS 0.10586f
C13494 VDAC_P.n2009 VSS 0.132855f
C13495 VDAC_P.t37 VSS 0.10586f
C13496 VDAC_P.n2010 VSS 0.132855f
C13497 VDAC_P.t1386 VSS 0.10586f
C13498 VDAC_P.n2011 VSS 0.132855f
C13499 VDAC_P.t876 VSS 0.10586f
C13500 VDAC_P.n2012 VSS 0.132855f
C13501 VDAC_P.t1614 VSS 0.10586f
C13502 VDAC_P.n2013 VSS 0.132855f
C13503 VDAC_P.t1320 VSS 0.10586f
C13504 VDAC_P.n2014 VSS 0.132855f
C13505 VDAC_P.t2027 VSS 0.10586f
C13506 VDAC_P.n2015 VSS 0.132855f
C13507 VDAC_P.t1784 VSS 0.10586f
C13508 VDAC_P.n2016 VSS 0.132855f
C13509 VDAC_P.t2133 VSS 0.10586f
C13510 VDAC_P.n2017 VSS 0.132855f
C13511 VDAC_P.t1330 VSS 0.10586f
C13512 VDAC_P.n2018 VSS 0.132855f
C13513 VDAC_P.t332 VSS 0.10586f
C13514 VDAC_P.n2019 VSS 0.132855f
C13515 VDAC_P.t1781 VSS 0.10586f
C13516 VDAC_P.n2020 VSS 0.132855f
C13517 VDAC_P.t1192 VSS 0.10586f
C13518 VDAC_P.n2021 VSS 0.132855f
C13519 VDAC_P.t1885 VSS 0.10586f
C13520 VDAC_P.n2022 VSS 0.132855f
C13521 VDAC_P.t203 VSS 0.10586f
C13522 VDAC_P.n2023 VSS 0.132855f
C13523 VDAC_P.t787 VSS 0.10586f
C13524 VDAC_P.n2024 VSS 0.132855f
C13525 VDAC_P.t27 VSS 0.10586f
C13526 VDAC_P.n2025 VSS 0.132855f
C13527 VDAC_P.t1944 VSS 0.10586f
C13528 VDAC_P.n2026 VSS 0.132855f
C13529 VDAC_P.t611 VSS 0.10586f
C13530 VDAC_P.n2027 VSS 0.132855f
C13531 VDAC_P.t378 VSS 0.10586f
C13532 VDAC_P.n2028 VSS 0.132855f
C13533 VDAC_P.t665 VSS 0.10586f
C13534 VDAC_P.n2029 VSS 0.132855f
C13535 VDAC_P.t1642 VSS 0.10586f
C13536 VDAC_P.n2030 VSS 0.132855f
C13537 VDAC_P.t1392 VSS 0.10586f
C13538 VDAC_P.n2031 VSS 0.132855f
C13539 VDAC_P.t1866 VSS 0.10586f
C13540 VDAC_P.n2032 VSS 0.132855f
C13541 VDAC_P.t256 VSS 0.10586f
C13542 VDAC_P.n2033 VSS 0.132855f
C13543 VDAC_P.t1756 VSS 0.10586f
C13544 VDAC_P.n2034 VSS 0.132855f
C13545 VDAC_P.t194 VSS 0.10586f
C13546 VDAC_P.n2035 VSS 0.132855f
C13547 VDAC_P.t396 VSS 0.10586f
C13548 VDAC_P.n2036 VSS 0.132855f
C13549 VDAC_P.t806 VSS 0.10586f
C13550 VDAC_P.n2037 VSS 0.132855f
C13551 VDAC_P.t1264 VSS 0.10586f
C13552 VDAC_P.n2038 VSS 0.128057f
C13553 VDAC_P.t1465 VSS 0.10586f
C13554 VDAC_P.n2039 VSS 0.138884f
C13555 VDAC_P.t1342 VSS 0.10586f
C13556 VDAC_P.n2040 VSS 0.144407f
C13557 VDAC_P.t2039 VSS 0.10586f
C13558 VDAC_P.n2041 VSS 0.144407f
C13559 VDAC_P.t1030 VSS 0.10586f
C13560 VDAC_P.n2042 VSS 0.144407f
C13561 VDAC_P.t1796 VSS 0.10586f
C13562 VDAC_P.n2043 VSS 0.144407f
C13563 VDAC_P.t1369 VSS 0.10586f
C13564 VDAC_P.n2044 VSS 0.144407f
C13565 VDAC_P.t1150 VSS 0.10586f
C13566 VDAC_P.n2045 VSS 0.144407f
C13567 VDAC_P.t1939 VSS 0.10586f
C13568 VDAC_P.n2046 VSS 0.144407f
C13569 VDAC_P.t579 VSS 0.10586f
C13570 VDAC_P.n2047 VSS 0.144407f
C13571 VDAC_P.t656 VSS 0.10586f
C13572 VDAC_P.n2048 VSS 0.144407f
C13573 VDAC_P.t208 VSS 0.10586f
C13574 VDAC_P.n2049 VSS 0.144407f
C13575 VDAC_P.t1173 VSS 0.10586f
C13576 VDAC_P.n2050 VSS 0.144407f
C13577 VDAC_P.t979 VSS 0.10586f
C13578 VDAC_P.n2051 VSS 0.144407f
C13579 VDAC_P.t1954 VSS 0.10586f
C13580 VDAC_P.n2052 VSS 0.144407f
C13581 VDAC_P.t893 VSS 0.10586f
C13582 VDAC_P.n2053 VSS 0.144407f
C13583 VDAC_P.t1266 VSS 0.10586f
C13584 VDAC_P.n2054 VSS 0.144407f
C13585 VDAC_P.t1421 VSS 0.10586f
C13586 VDAC_P.n2055 VSS 0.144407f
C13587 VDAC_P.t1148 VSS 0.10586f
C13588 VDAC_P.n2056 VSS 0.144407f
C13589 VDAC_P.t61 VSS 0.10586f
C13590 VDAC_P.n2057 VSS 0.144407f
C13591 VDAC_P.t1851 VSS 0.10586f
C13592 VDAC_P.n2058 VSS 0.144407f
C13593 VDAC_P.t1470 VSS 0.10586f
C13594 VDAC_P.n2059 VSS 0.144407f
C13595 VDAC_P.t775 VSS 0.10586f
C13596 VDAC_P.n2060 VSS 0.144407f
C13597 VDAC_P.t1004 VSS 0.10586f
C13598 VDAC_P.n2061 VSS 0.144407f
C13599 VDAC_P.t1185 VSS 0.10586f
C13600 VDAC_P.n2062 VSS 0.144407f
C13601 VDAC_P.t989 VSS 0.10586f
C13602 VDAC_P.n2063 VSS 0.144407f
C13603 VDAC_P.t1646 VSS 0.10586f
C13604 VDAC_P.n2064 VSS 0.144407f
C13605 VDAC_P.t425 VSS 0.10586f
C13606 VDAC_P.n2065 VSS 0.144407f
C13607 VDAC_P.t1844 VSS 0.10586f
C13608 VDAC_P.n2066 VSS 0.144407f
C13609 VDAC_P.t653 VSS 0.10586f
C13610 VDAC_P.n2067 VSS 0.144407f
C13611 VDAC_P.t2043 VSS 0.10586f
C13612 VDAC_P.n2068 VSS 0.138884f
C13613 VDAC_P.t1842 VSS 0.10586f
C13614 VDAC_P.n2069 VSS 0.128057f
C13615 VDAC_P.t709 VSS 0.10586f
C13616 VDAC_P.n2070 VSS 0.132855f
C13617 VDAC_P.t714 VSS 0.10586f
C13618 VDAC_P.n2071 VSS 0.132855f
C13619 VDAC_P.t343 VSS 0.10586f
C13620 VDAC_P.n2072 VSS 0.132855f
C13621 VDAC_P.t318 VSS 0.10586f
C13622 VDAC_P.n2073 VSS 0.132855f
C13623 VDAC_P.t2110 VSS 0.10586f
C13624 VDAC_P.n2074 VSS 0.132855f
C13625 VDAC_P.t781 VSS 0.10586f
C13626 VDAC_P.n2075 VSS 0.132855f
C13627 VDAC_P.t966 VSS 0.10586f
C13628 VDAC_P.n2076 VSS 0.132855f
C13629 VDAC_P.t725 VSS 0.10586f
C13630 VDAC_P.n2077 VSS 0.132855f
C13631 VDAC_P.t1877 VSS 0.10586f
C13632 VDAC_P.n2078 VSS 0.132855f
C13633 VDAC_P.t109 VSS 0.10586f
C13634 VDAC_P.n2079 VSS 0.132855f
C13635 VDAC_P.t1771 VSS 0.10586f
C13636 VDAC_P.n2080 VSS 0.132855f
C13637 VDAC_P.t1105 VSS 0.10586f
C13638 VDAC_P.n2081 VSS 0.132855f
C13639 VDAC_P.t851 VSS 0.10586f
C13640 VDAC_P.n2082 VSS 0.132855f
C13641 VDAC_P.t2125 VSS 0.10586f
C13642 VDAC_P.n2083 VSS 0.132855f
C13643 VDAC_P.t832 VSS 0.10586f
C13644 VDAC_P.n2084 VSS 0.132855f
C13645 VDAC_P.t890 VSS 0.10586f
C13646 VDAC_P.n2085 VSS 0.132855f
C13647 VDAC_P.t1461 VSS 0.10586f
C13648 VDAC_P.n2086 VSS 0.132855f
C13649 VDAC_P.t1546 VSS 0.10586f
C13650 VDAC_P.n2087 VSS 0.132855f
C13651 VDAC_P.t1249 VSS 0.10586f
C13652 VDAC_P.n2088 VSS 0.132855f
C13653 VDAC_P.t917 VSS 0.10586f
C13654 VDAC_P.n2089 VSS 0.132855f
C13655 VDAC_P.t1143 VSS 0.10586f
C13656 VDAC_P.n2090 VSS 0.132855f
C13657 VDAC_P.t1597 VSS 0.10586f
C13658 VDAC_P.n2091 VSS 0.132855f
C13659 VDAC_P.t2030 VSS 0.10586f
C13660 VDAC_P.n2092 VSS 0.132855f
C13661 VDAC_P.t1491 VSS 0.10586f
C13662 VDAC_P.n2093 VSS 0.132855f
C13663 VDAC_P.t1945 VSS 0.10586f
C13664 VDAC_P.n2094 VSS 0.132855f
C13665 VDAC_P.t651 VSS 0.10586f
C13666 VDAC_P.n2095 VSS 0.132855f
C13667 VDAC_P.t1835 VSS 0.10586f
C13668 VDAC_P.n2096 VSS 0.132855f
C13669 VDAC_P.t1092 VSS 0.10586f
C13670 VDAC_P.n2097 VSS 0.132855f
C13671 VDAC_P.t1625 VSS 0.10586f
C13672 VDAC_P.n2098 VSS 0.132855f
C13673 VDAC_P.t1052 VSS 0.10586f
C13674 VDAC_P.n2099 VSS 0.132855f
C13675 VDAC_P.t1519 VSS 0.10586f
C13676 VDAC_P.n2100 VSS 0.132855f
C13677 VDAC_P.t515 VSS 0.10586f
C13678 VDAC_P.n2101 VSS 0.132855f
C13679 VDAC_P.t800 VSS 0.10586f
C13680 VDAC_P.n2102 VSS 0.132855f
C13681 VDAC_P.t257 VSS 0.10586f
C13682 VDAC_P.n2103 VSS 0.132855f
C13683 VDAC_P.t1364 VSS 0.10586f
C13684 VDAC_P.n2104 VSS 0.132855f
C13685 VDAC_P.t662 VSS 0.10586f
C13686 VDAC_P.n2105 VSS 0.132855f
C13687 VDAC_P.t1788 VSS 0.10586f
C13688 VDAC_P.n2106 VSS 0.132855f
C13689 VDAC_P.t2128 VSS 0.10586f
C13690 VDAC_P.n2107 VSS 0.132855f
C13691 VDAC_P.t275 VSS 0.10586f
C13692 VDAC_P.n2108 VSS 0.132855f
C13693 VDAC_P.t1712 VSS 0.10586f
C13694 VDAC_P.n2109 VSS 0.132855f
C13695 VDAC_P.t1782 VSS 0.10586f
C13696 VDAC_P.n2110 VSS 0.132855f
C13697 VDAC_P.t1144 VSS 0.10586f
C13698 VDAC_P.n2111 VSS 0.132855f
C13699 VDAC_P.t1742 VSS 0.10586f
C13700 VDAC_P.n2112 VSS 0.132855f
C13701 VDAC_P.t1349 VSS 0.10586f
C13702 VDAC_P.n2113 VSS 0.132855f
C13703 VDAC_P.t666 VSS 0.10586f
C13704 VDAC_P.n2114 VSS 0.132855f
C13705 VDAC_P.t167 VSS 0.10586f
C13706 VDAC_P.n2115 VSS 0.132855f
C13707 VDAC_P.t863 VSS 0.10586f
C13708 VDAC_P.n2116 VSS 0.132855f
C13709 VDAC_P.t2014 VSS 0.10586f
C13710 VDAC_P.n2117 VSS 0.132855f
C13711 VDAC_P.t1487 VSS 0.10586f
C13712 VDAC_P.n2118 VSS 0.132855f
C13713 VDAC_P.t470 VSS 0.10586f
C13714 VDAC_P.n2119 VSS 0.132855f
C13715 VDAC_P.t701 VSS 0.10586f
C13716 VDAC_P.n2120 VSS 0.132855f
C13717 VDAC_P.t929 VSS 0.10586f
C13718 VDAC_P.n2121 VSS 0.132855f
C13719 VDAC_P.t647 VSS 0.10586f
C13720 VDAC_P.n2122 VSS 0.132855f
C13721 VDAC_P.t81 VSS 0.10586f
C13722 VDAC_P.n2123 VSS 0.132855f
C13723 VDAC_P.t1564 VSS 0.10586f
C13724 VDAC_P.n2124 VSS 0.132855f
C13725 VDAC_P.t1517 VSS 0.10586f
C13726 VDAC_P.n2125 VSS 0.132855f
C13727 VDAC_P.t2073 VSS 0.10586f
C13728 VDAC_P.n2126 VSS 0.132855f
C13729 VDAC_P.t371 VSS 0.10586f
C13730 VDAC_P.n2127 VSS 0.132855f
C13731 VDAC_P.t943 VSS 0.10586f
C13732 VDAC_P.n2128 VSS 0.132855f
C13733 VDAC_P.t1104 VSS 0.10586f
C13734 VDAC_P.n2129 VSS 0.132855f
C13735 VDAC_P.t1753 VSS 0.10586f
C13736 VDAC_P.n2130 VSS 0.132855f
C13737 VDAC_P.t892 VSS 0.10586f
C13738 VDAC_P.n2131 VSS 0.132855f
C13739 VDAC_P.t342 VSS 0.10586f
C13740 VDAC_P.n2132 VSS 0.132855f
C13741 VDAC_P.t2101 VSS 0.10586f
C13742 VDAC_P.n2133 VSS 0.132855f
C13743 VDAC_P.t1696 VSS 0.10586f
C13744 VDAC_P.n2134 VSS 0.135114f
C13745 C6_N_btm.t1 VSS 1.04079f
C13746 C6_N_btm.n0 VSS 0.153224f
C13747 C6_N_btm.n2 VSS 0.837748f
C13748 C6_N_btm.n3 VSS 1.30605f
C13749 C6_N_btm.n4 VSS 1.89772f
C13750 C6_N_btm.n5 VSS 0.115577f
C13751 C6_N_btm.t55 VSS 0.512522f
C13752 C6_N_btm.t68 VSS 0.532791f
C13753 C6_N_btm.n6 VSS 0.115577f
C13754 C6_N_btm.n7 VSS 0.115577f
C13755 C6_N_btm.t17 VSS 0.512522f
C13756 C6_N_btm.n8 VSS 0.119988f
C13757 C6_N_btm.t12 VSS 0.512522f
C13758 C6_N_btm.n20 VSS 0.159599f
C13759 C6_N_btm.t31 VSS 0.512522f
C13760 C6_N_btm.n21 VSS 0.159599f
C13761 C6_N_btm.n28 VSS 0.115577f
C13762 C6_N_btm.n34 VSS 0.115577f
C13763 C6_N_btm.n35 VSS 0.115577f
C13764 C6_N_btm.t61 VSS 0.512522f
C13765 C6_N_btm.t67 VSS 0.532791f
C13766 C6_N_btm.n36 VSS 0.193911f
C13767 C6_N_btm.t66 VSS 0.532791f
C13768 C6_N_btm.t50 VSS 0.512522f
C13769 C6_N_btm.t8 VSS 0.512522f
C13770 C6_N_btm.n39 VSS 0.193911f
C13771 C6_N_btm.n40 VSS 0.115577f
C13772 C6_N_btm.t57 VSS 0.512522f
C13773 C6_N_btm.t5 VSS 0.512522f
C13774 C6_N_btm.n43 VSS 0.115577f
C13775 C6_N_btm.t29 VSS 0.512522f
C13776 C6_N_btm.t26 VSS 0.512522f
C13777 C6_N_btm.n46 VSS 0.115577f
C13778 C6_N_btm.n47 VSS 0.115577f
C13779 C6_N_btm.t37 VSS 0.512522f
C13780 C6_N_btm.n50 VSS 0.115577f
C13781 C6_N_btm.t53 VSS 0.512522f
C13782 C6_N_btm.t65 VSS 0.512522f
C13783 C6_N_btm.n53 VSS 0.115577f
C13784 C6_N_btm.n54 VSS 0.115577f
C13785 C6_N_btm.t48 VSS 0.512522f
C13786 C6_N_btm.t22 VSS 0.512522f
C13787 C6_N_btm.n57 VSS 0.115577f
C13788 C6_N_btm.t54 VSS 0.512522f
C13789 C6_N_btm.t46 VSS 0.462125f
C13790 C6_N_btm.t32 VSS 0.462125f
C13791 C6_N_btm.t24 VSS 0.462125f
C13792 C6_N_btm.t36 VSS 0.512522f
C13793 C6_N_btm.n69 VSS 0.109928f
C13794 C6_N_btm.t15 VSS 0.462125f
C13795 C6_N_btm.t62 VSS 0.462125f
C13796 C6_N_btm.t4 VSS 0.462125f
C13797 C6_N_btm.t49 VSS 0.462125f
C13798 C6_N_btm.t42 VSS 0.462125f
C13799 C6_N_btm.t11 VSS 0.462125f
C13800 C6_N_btm.t40 VSS 0.462125f
C13801 C6_N_btm.t3 VSS 0.462125f
C13802 C6_N_btm.t30 VSS 0.512522f
C13803 C6_N_btm.n100 VSS 0.119988f
C13804 C6_N_btm.t9 VSS 0.512522f
C13805 C6_N_btm.n101 VSS 0.156187f
C13806 C6_N_btm.t27 VSS 0.462125f
C13807 C6_N_btm.t14 VSS 0.462125f
C13808 C6_N_btm.t33 VSS 0.462125f
C13809 C6_N_btm.t18 VSS 0.462125f
C13810 C6_N_btm.t52 VSS 0.462125f
C13811 C6_N_btm.t25 VSS 0.462125f
C13812 C6_N_btm.t6 VSS 0.462125f
C13813 C6_N_btm.t28 VSS 0.462125f
C13814 C6_N_btm.t13 VSS 0.462125f
C13815 C6_N_btm.t45 VSS 0.462125f
C13816 C6_N_btm.t16 VSS 0.462125f
C13817 C6_N_btm.t2 VSS 0.512522f
C13818 C6_N_btm.n136 VSS 0.156187f
C13819 C6_N_btm.t43 VSS 0.462125f
C13820 C6_N_btm.t7 VSS 0.512522f
C13821 C6_N_btm.t56 VSS 0.462125f
C13822 C6_N_btm.t41 VSS 0.462125f
C13823 C6_N_btm.t19 VSS 0.462125f
C13824 C6_N_btm.t39 VSS 0.462125f
C13825 C6_N_btm.t64 VSS 0.512522f
C13826 C6_N_btm.n154 VSS 0.109928f
C13827 C6_N_btm.t51 VSS 0.462125f
C13828 C6_N_btm.t34 VSS 0.462125f
C13829 C6_N_btm.t20 VSS 0.462125f
C13830 C6_N_btm.t60 VSS 0.512522f
C13831 C6_N_btm.n165 VSS 0.115577f
C13832 C6_N_btm.t44 VSS 0.512522f
C13833 C6_N_btm.t23 VSS 0.512522f
C13834 C6_N_btm.n168 VSS 0.115577f
C13835 C6_N_btm.n169 VSS 0.115577f
C13836 C6_N_btm.t38 VSS 0.512522f
C13837 C6_N_btm.n172 VSS 0.115577f
C13838 C6_N_btm.t10 VSS 0.512522f
C13839 C6_N_btm.t63 VSS 0.512522f
C13840 C6_N_btm.n175 VSS 0.115577f
C13841 C6_N_btm.n176 VSS 0.115577f
C13842 C6_N_btm.t59 VSS 0.512522f
C13843 C6_N_btm.t35 VSS 0.512522f
C13844 C6_N_btm.n179 VSS 0.115577f
C13845 C6_N_btm.t47 VSS 0.512522f
C13846 C6_N_btm.t58 VSS 0.512522f
C13847 C6_N_btm.n182 VSS 0.115577f
C13848 C6_N_btm.n183 VSS 0.193911f
C13849 C6_N_btm.t21 VSS 0.512522f
C13850 C6_N_btm.n186 VSS 0.115577f
C13851 C6_N_btm.t69 VSS 0.513385f
C13852 C6_N_btm.n187 VSS 0.295219f
C13853 VDAC_N.t1522 VSS 0.102761f
C13854 VDAC_N.t1438 VSS 0.102718f
C13855 VDAC_N.n0 VSS 0.114855f
C13856 VDAC_N.t702 VSS 0.102718f
C13857 VDAC_N.t1772 VSS 0.102718f
C13858 VDAC_N.t138 VSS 0.102761f
C13859 VDAC_N.t184 VSS 0.102718f
C13860 VDAC_N.n3 VSS 0.114855f
C13861 VDAC_N.t584 VSS 0.102718f
C13862 VDAC_N.t955 VSS 0.102718f
C13863 VDAC_N.n5 VSS 0.119671f
C13864 VDAC_N.t363 VSS 0.102718f
C13865 VDAC_N.n6 VSS 0.11953f
C13866 VDAC_N.t1397 VSS 0.102718f
C13867 VDAC_N.t1423 VSS 0.102718f
C13868 VDAC_N.t284 VSS 0.102718f
C13869 VDAC_N.t1756 VSS 0.102761f
C13870 VDAC_N.t925 VSS 0.102718f
C13871 VDAC_N.n10 VSS 0.114855f
C13872 VDAC_N.t1791 VSS 0.102718f
C13873 VDAC_N.t627 VSS 0.102718f
C13874 VDAC_N.n15 VSS 0.267352f
C13875 VDAC_N.n16 VSS 0.261101f
C13876 VDAC_N.n17 VSS 0.36829f
C13877 VDAC_N.n18 VSS 0.267352f
C13878 VDAC_N.n19 VSS 0.261101f
C13879 VDAC_N.n20 VSS 0.367761f
C13880 VDAC_N.n21 VSS 0.364104f
C13881 VDAC_N.n22 VSS 2.37284f
C13882 VDAC_N.t1380 VSS 0.105768f
C13883 VDAC_N.n23 VSS 0.137176f
C13884 VDAC_N.t1691 VSS 0.105768f
C13885 VDAC_N.n24 VSS 0.12675f
C13886 VDAC_N.t1588 VSS 0.105768f
C13887 VDAC_N.n25 VSS 0.132739f
C13888 VDAC_N.t469 VSS 0.105768f
C13889 VDAC_N.n26 VSS 0.132739f
C13890 VDAC_N.t1335 VSS 0.105768f
C13891 VDAC_N.n27 VSS 0.132739f
C13892 VDAC_N.t2001 VSS 0.105768f
C13893 VDAC_N.n28 VSS 0.132739f
C13894 VDAC_N.t1441 VSS 0.105768f
C13895 VDAC_N.n29 VSS 0.132739f
C13896 VDAC_N.t1938 VSS 0.105768f
C13897 VDAC_N.n30 VSS 0.132739f
C13898 VDAC_N.t843 VSS 0.105768f
C13899 VDAC_N.n31 VSS 0.132739f
C13900 VDAC_N.t17 VSS 0.105768f
C13901 VDAC_N.n32 VSS 0.132739f
C13902 VDAC_N.t1761 VSS 0.105768f
C13903 VDAC_N.n33 VSS 0.132739f
C13904 VDAC_N.t1303 VSS 0.105768f
C13905 VDAC_N.n34 VSS 0.132739f
C13906 VDAC_N.t1642 VSS 0.105768f
C13907 VDAC_N.n35 VSS 0.132739f
C13908 VDAC_N.t1413 VSS 0.105768f
C13909 VDAC_N.n36 VSS 0.132739f
C13910 VDAC_N.t1862 VSS 0.105768f
C13911 VDAC_N.n37 VSS 0.132739f
C13912 VDAC_N.t1848 VSS 0.105768f
C13913 VDAC_N.n38 VSS 0.132739f
C13914 VDAC_N.t2082 VSS 0.105768f
C13915 VDAC_N.n39 VSS 0.132739f
C13916 VDAC_N.t98 VSS 0.105768f
C13917 VDAC_N.n40 VSS 0.132739f
C13918 VDAC_N.t649 VSS 0.105768f
C13919 VDAC_N.n41 VSS 0.132739f
C13920 VDAC_N.t1354 VSS 0.105768f
C13921 VDAC_N.n42 VSS 0.132739f
C13922 VDAC_N.t1684 VSS 0.105768f
C13923 VDAC_N.n43 VSS 0.132739f
C13924 VDAC_N.t1810 VSS 0.105768f
C13925 VDAC_N.n44 VSS 0.132739f
C13926 VDAC_N.t880 VSS 0.105768f
C13927 VDAC_N.n45 VSS 0.132739f
C13928 VDAC_N.t59 VSS 0.105768f
C13929 VDAC_N.n46 VSS 0.132739f
C13930 VDAC_N.t1840 VSS 0.105768f
C13931 VDAC_N.n47 VSS 0.132739f
C13932 VDAC_N.t2122 VSS 0.105768f
C13933 VDAC_N.n48 VSS 0.132739f
C13934 VDAC_N.t805 VSS 0.105768f
C13935 VDAC_N.n49 VSS 0.132739f
C13936 VDAC_N.t780 VSS 0.105768f
C13937 VDAC_N.n50 VSS 0.132739f
C13938 VDAC_N.t1797 VSS 0.105768f
C13939 VDAC_N.n51 VSS 0.132739f
C13940 VDAC_N.t836 VSS 0.105768f
C13941 VDAC_N.n52 VSS 0.132739f
C13942 VDAC_N.t497 VSS 0.105768f
C13943 VDAC_N.n53 VSS 0.132739f
C13944 VDAC_N.t737 VSS 0.105768f
C13945 VDAC_N.n54 VSS 0.132739f
C13946 VDAC_N.t551 VSS 0.105768f
C13947 VDAC_N.n55 VSS 0.132739f
C13948 VDAC_N.t1553 VSS 0.105768f
C13949 VDAC_N.n56 VSS 0.132739f
C13950 VDAC_N.t555 VSS 0.105768f
C13951 VDAC_N.n57 VSS 0.132739f
C13952 VDAC_N.t1765 VSS 0.105768f
C13953 VDAC_N.n58 VSS 0.132739f
C13954 VDAC_N.t1199 VSS 0.105768f
C13955 VDAC_N.n59 VSS 0.132739f
C13956 VDAC_N.t1881 VSS 0.105768f
C13957 VDAC_N.n60 VSS 0.132739f
C13958 VDAC_N.t375 VSS 0.105768f
C13959 VDAC_N.n61 VSS 0.132739f
C13960 VDAC_N.t842 VSS 0.105768f
C13961 VDAC_N.n62 VSS 0.132739f
C13962 VDAC_N.t1523 VSS 0.105768f
C13963 VDAC_N.n63 VSS 0.132739f
C13964 VDAC_N.t1058 VSS 0.105768f
C13965 VDAC_N.n64 VSS 0.132739f
C13966 VDAC_N.t1158 VSS 0.105768f
C13967 VDAC_N.n65 VSS 0.132739f
C13968 VDAC_N.t1169 VSS 0.105768f
C13969 VDAC_N.n66 VSS 0.132739f
C13970 VDAC_N.t362 VSS 0.105768f
C13971 VDAC_N.n67 VSS 0.132739f
C13972 VDAC_N.t1387 VSS 0.105768f
C13973 VDAC_N.n68 VSS 0.132739f
C13974 VDAC_N.t818 VSS 0.105768f
C13975 VDAC_N.n69 VSS 0.132739f
C13976 VDAC_N.t1304 VSS 0.105768f
C13977 VDAC_N.n70 VSS 0.132739f
C13978 VDAC_N.t2034 VSS 0.105768f
C13979 VDAC_N.n71 VSS 0.132739f
C13980 VDAC_N.t1752 VSS 0.105768f
C13981 VDAC_N.n72 VSS 0.132739f
C13982 VDAC_N.t1079 VSS 0.105768f
C13983 VDAC_N.n73 VSS 0.132739f
C13984 VDAC_N.t868 VSS 0.105768f
C13985 VDAC_N.n74 VSS 0.132739f
C13986 VDAC_N.t1907 VSS 0.105768f
C13987 VDAC_N.n75 VSS 0.132739f
C13988 VDAC_N.t193 VSS 0.105768f
C13989 VDAC_N.n76 VSS 0.132739f
C13990 VDAC_N.t1021 VSS 0.105768f
C13991 VDAC_N.n77 VSS 0.132739f
C13992 VDAC_N.t1557 VSS 0.105768f
C13993 VDAC_N.n78 VSS 0.132739f
C13994 VDAC_N.t1077 VSS 0.105768f
C13995 VDAC_N.n79 VSS 0.132739f
C13996 VDAC_N.t847 VSS 0.105768f
C13997 VDAC_N.n80 VSS 0.132739f
C13998 VDAC_N.t175 VSS 0.105768f
C13999 VDAC_N.n81 VSS 0.132739f
C14000 VDAC_N.t137 VSS 0.105768f
C14001 VDAC_N.n82 VSS 0.132739f
C14002 VDAC_N.t1315 VSS 0.105768f
C14003 VDAC_N.n83 VSS 0.132739f
C14004 VDAC_N.t846 VSS 0.105768f
C14005 VDAC_N.n84 VSS 0.132739f
C14006 VDAC_N.t403 VSS 0.105768f
C14007 VDAC_N.n85 VSS 0.132739f
C14008 VDAC_N.t494 VSS 0.105768f
C14009 VDAC_N.n86 VSS 0.132739f
C14010 VDAC_N.t431 VSS 0.105768f
C14011 VDAC_N.n87 VSS 0.12675f
C14012 VDAC_N.t1028 VSS 0.105768f
C14013 VDAC_N.n88 VSS 0.12675f
C14014 VDAC_N.t187 VSS 0.105768f
C14015 VDAC_N.n89 VSS 0.12675f
C14016 VDAC_N.t1049 VSS 0.105768f
C14017 VDAC_N.n90 VSS 0.12675f
C14018 VDAC_N.t1394 VSS 0.105768f
C14019 VDAC_N.n91 VSS 0.12675f
C14020 VDAC_N.t1733 VSS 0.105768f
C14021 VDAC_N.n92 VSS 0.12675f
C14022 VDAC_N.t712 VSS 0.105768f
C14023 VDAC_N.n93 VSS 0.12675f
C14024 VDAC_N.t713 VSS 0.105768f
C14025 VDAC_N.n94 VSS 0.12675f
C14026 VDAC_N.t1820 VSS 0.105768f
C14027 VDAC_N.n95 VSS 0.12675f
C14028 VDAC_N.t814 VSS 0.105768f
C14029 VDAC_N.n96 VSS 0.12675f
C14030 VDAC_N.t253 VSS 0.105768f
C14031 VDAC_N.n97 VSS 0.12675f
C14032 VDAC_N.t472 VSS 0.105768f
C14033 VDAC_N.n98 VSS 0.12675f
C14034 VDAC_N.t1487 VSS 0.105768f
C14035 VDAC_N.n99 VSS 0.12675f
C14036 VDAC_N.t76 VSS 0.105768f
C14037 VDAC_N.n100 VSS 0.12675f
C14038 VDAC_N.t1786 VSS 0.105768f
C14039 VDAC_N.n101 VSS 0.12675f
C14040 VDAC_N.t1921 VSS 0.105768f
C14041 VDAC_N.n102 VSS 0.12675f
C14042 VDAC_N.t562 VSS 0.105768f
C14043 VDAC_N.n103 VSS 0.12675f
C14044 VDAC_N.t1585 VSS 0.105768f
C14045 VDAC_N.n104 VSS 0.12675f
C14046 VDAC_N.t804 VSS 0.105768f
C14047 VDAC_N.n105 VSS 0.12675f
C14048 VDAC_N.t1006 VSS 0.105768f
C14049 VDAC_N.n106 VSS 0.12675f
C14050 VDAC_N.t297 VSS 0.105768f
C14051 VDAC_N.n107 VSS 0.12675f
C14052 VDAC_N.t57 VSS 0.105768f
C14053 VDAC_N.n108 VSS 0.12675f
C14054 VDAC_N.t1506 VSS 0.105768f
C14055 VDAC_N.n109 VSS 0.12675f
C14056 VDAC_N.t407 VSS 0.105768f
C14057 VDAC_N.n110 VSS 0.12675f
C14058 VDAC_N.t180 VSS 0.105768f
C14059 VDAC_N.n111 VSS 0.12675f
C14060 VDAC_N.t615 VSS 0.105768f
C14061 VDAC_N.n112 VSS 0.12675f
C14062 VDAC_N.t1975 VSS 0.105768f
C14063 VDAC_N.n113 VSS 0.12675f
C14064 VDAC_N.t1694 VSS 0.105768f
C14065 VDAC_N.n114 VSS 0.12675f
C14066 VDAC_N.t835 VSS 0.105768f
C14067 VDAC_N.n115 VSS 0.12675f
C14068 VDAC_N.t2036 VSS 0.105768f
C14069 VDAC_N.n116 VSS 0.12675f
C14070 VDAC_N.t1739 VSS 0.105768f
C14071 VDAC_N.n117 VSS 0.132739f
C14072 VDAC_N.t164 VSS 0.105768f
C14073 VDAC_N.n118 VSS 0.132739f
C14074 VDAC_N.t829 VSS 0.105768f
C14075 VDAC_N.n119 VSS 0.132739f
C14076 VDAC_N.t2091 VSS 0.105768f
C14077 VDAC_N.n120 VSS 0.132739f
C14078 VDAC_N.t808 VSS 0.105768f
C14079 VDAC_N.n121 VSS 0.132739f
C14080 VDAC_N.t1979 VSS 0.105768f
C14081 VDAC_N.n122 VSS 0.132739f
C14082 VDAC_N.t1152 VSS 0.105768f
C14083 VDAC_N.n123 VSS 0.132739f
C14084 VDAC_N.t402 VSS 0.105768f
C14085 VDAC_N.n124 VSS 0.132739f
C14086 VDAC_N.t1396 VSS 0.105768f
C14087 VDAC_N.n125 VSS 0.132739f
C14088 VDAC_N.t1290 VSS 0.105768f
C14089 VDAC_N.n126 VSS 0.132739f
C14090 VDAC_N.t2121 VSS 0.105768f
C14091 VDAC_N.n127 VSS 0.132739f
C14092 VDAC_N.t552 VSS 0.105768f
C14093 VDAC_N.n128 VSS 0.132739f
C14094 VDAC_N.t1022 VSS 0.105768f
C14095 VDAC_N.n129 VSS 0.132739f
C14096 VDAC_N.t638 VSS 0.105768f
C14097 VDAC_N.n130 VSS 0.132739f
C14098 VDAC_N.t295 VSS 0.105768f
C14099 VDAC_N.n131 VSS 0.132739f
C14100 VDAC_N.t1675 VSS 0.105768f
C14101 VDAC_N.n132 VSS 0.132739f
C14102 VDAC_N.t1970 VSS 0.105768f
C14103 VDAC_N.n133 VSS 0.132739f
C14104 VDAC_N.t1457 VSS 0.105768f
C14105 VDAC_N.n134 VSS 0.132739f
C14106 VDAC_N.t1025 VSS 0.105768f
C14107 VDAC_N.n135 VSS 0.132739f
C14108 VDAC_N.t111 VSS 0.105768f
C14109 VDAC_N.n136 VSS 0.132739f
C14110 VDAC_N.t1809 VSS 0.105768f
C14111 VDAC_N.n137 VSS 0.132739f
C14112 VDAC_N.t633 VSS 0.105768f
C14113 VDAC_N.n138 VSS 0.132739f
C14114 VDAC_N.t1705 VSS 0.105768f
C14115 VDAC_N.n139 VSS 0.132739f
C14116 VDAC_N.t1692 VSS 0.105768f
C14117 VDAC_N.n140 VSS 0.132739f
C14118 VDAC_N.t119 VSS 0.105768f
C14119 VDAC_N.n141 VSS 0.132739f
C14120 VDAC_N.t2053 VSS 0.105768f
C14121 VDAC_N.n142 VSS 0.132739f
C14122 VDAC_N.t1432 VSS 0.105768f
C14123 VDAC_N.n143 VSS 0.132739f
C14124 VDAC_N.t1841 VSS 0.105768f
C14125 VDAC_N.n144 VSS 0.132739f
C14126 VDAC_N.t1012 VSS 0.105768f
C14127 VDAC_N.n145 VSS 0.132739f
C14128 VDAC_N.t241 VSS 0.105768f
C14129 VDAC_N.n146 VSS 0.132739f
C14130 VDAC_N.t2012 VSS 0.105768f
C14131 VDAC_N.n147 VSS 0.132739f
C14132 VDAC_N.t626 VSS 0.105768f
C14133 VDAC_N.n148 VSS 0.132739f
C14134 VDAC_N.t285 VSS 0.105768f
C14135 VDAC_N.n149 VSS 0.132739f
C14136 VDAC_N.t1552 VSS 0.105768f
C14137 VDAC_N.n150 VSS 0.132739f
C14138 VDAC_N.t134 VSS 0.105768f
C14139 VDAC_N.n151 VSS 0.132739f
C14140 VDAC_N.t96 VSS 0.105768f
C14141 VDAC_N.n152 VSS 0.132739f
C14142 VDAC_N.t766 VSS 0.105768f
C14143 VDAC_N.n153 VSS 0.132739f
C14144 VDAC_N.t1020 VSS 0.105768f
C14145 VDAC_N.n154 VSS 0.132739f
C14146 VDAC_N.t654 VSS 0.105768f
C14147 VDAC_N.n155 VSS 0.132739f
C14148 VDAC_N.t573 VSS 0.105768f
C14149 VDAC_N.n156 VSS 0.132739f
C14150 VDAC_N.t1024 VSS 0.105768f
C14151 VDAC_N.n157 VSS 0.132739f
C14152 VDAC_N.t293 VSS 0.105768f
C14153 VDAC_N.n158 VSS 0.132739f
C14154 VDAC_N.t793 VSS 0.105768f
C14155 VDAC_N.n159 VSS 0.132739f
C14156 VDAC_N.t454 VSS 0.105768f
C14157 VDAC_N.n160 VSS 0.132739f
C14158 VDAC_N.t1349 VSS 0.105768f
C14159 VDAC_N.n161 VSS 0.132739f
C14160 VDAC_N.t263 VSS 0.105768f
C14161 VDAC_N.n162 VSS 0.132739f
C14162 VDAC_N.t329 VSS 0.105768f
C14163 VDAC_N.n163 VSS 0.132739f
C14164 VDAC_N.t1701 VSS 0.105768f
C14165 VDAC_N.n164 VSS 0.132739f
C14166 VDAC_N.t1125 VSS 0.105768f
C14167 VDAC_N.n165 VSS 0.132739f
C14168 VDAC_N.t809 VSS 0.105768f
C14169 VDAC_N.n166 VSS 0.132739f
C14170 VDAC_N.t2047 VSS 0.105768f
C14171 VDAC_N.n167 VSS 0.132739f
C14172 VDAC_N.t753 VSS 0.105768f
C14173 VDAC_N.n168 VSS 0.132739f
C14174 VDAC_N.t1937 VSS 0.105768f
C14175 VDAC_N.n169 VSS 0.132739f
C14176 VDAC_N.t1940 VSS 0.105768f
C14177 VDAC_N.n170 VSS 0.132739f
C14178 VDAC_N.t877 VSS 0.105768f
C14179 VDAC_N.n171 VSS 0.132739f
C14180 VDAC_N.t2060 VSS 0.105768f
C14181 VDAC_N.n172 VSS 0.132739f
C14182 VDAC_N.t823 VSS 0.105768f
C14183 VDAC_N.n173 VSS 0.132739f
C14184 VDAC_N.t2079 VSS 0.105768f
C14185 VDAC_N.n174 VSS 0.132739f
C14186 VDAC_N.t1976 VSS 0.105768f
C14187 VDAC_N.n175 VSS 0.132739f
C14188 VDAC_N.t997 VSS 0.105768f
C14189 VDAC_N.n176 VSS 0.132739f
C14190 VDAC_N.t1112 VSS 0.105768f
C14191 VDAC_N.n177 VSS 0.132739f
C14192 VDAC_N.t1714 VSS 0.105768f
C14193 VDAC_N.n178 VSS 0.132739f
C14194 VDAC_N.t1316 VSS 0.105768f
C14195 VDAC_N.n179 VSS 0.12675f
C14196 VDAC_N.t262 VSS 0.105768f
C14197 VDAC_N.n180 VSS 0.132739f
C14198 VDAC_N.t779 VSS 0.105768f
C14199 VDAC_N.n181 VSS 0.132739f
C14200 VDAC_N.t1670 VSS 0.105768f
C14201 VDAC_N.n182 VSS 0.132739f
C14202 VDAC_N.t351 VSS 0.105768f
C14203 VDAC_N.n183 VSS 0.132739f
C14204 VDAC_N.t1775 VSS 0.105768f
C14205 VDAC_N.n184 VSS 0.132739f
C14206 VDAC_N.t323 VSS 0.105768f
C14207 VDAC_N.n185 VSS 0.132739f
C14208 VDAC_N.t1671 VSS 0.105768f
C14209 VDAC_N.n186 VSS 0.132739f
C14210 VDAC_N.t2129 VSS 0.105768f
C14211 VDAC_N.n187 VSS 0.132739f
C14212 VDAC_N.t795 VSS 0.105768f
C14213 VDAC_N.n188 VSS 0.132739f
C14214 VDAC_N.t1023 VSS 0.105768f
C14215 VDAC_N.n189 VSS 0.132739f
C14216 VDAC_N.t359 VSS 0.105768f
C14217 VDAC_N.n190 VSS 0.132739f
C14218 VDAC_N.t1911 VSS 0.105768f
C14219 VDAC_N.n191 VSS 0.132739f
C14220 VDAC_N.t1732 VSS 0.105768f
C14221 VDAC_N.n192 VSS 0.132739f
C14222 VDAC_N.t1720 VSS 0.105768f
C14223 VDAC_N.n193 VSS 0.132739f
C14224 VDAC_N.t470 VSS 0.105768f
C14225 VDAC_N.n194 VSS 0.132739f
C14226 VDAC_N.t1479 VSS 0.105768f
C14227 VDAC_N.n195 VSS 0.132739f
C14228 VDAC_N.t418 VSS 0.105768f
C14229 VDAC_N.n196 VSS 0.132739f
C14230 VDAC_N.t337 VSS 0.105768f
C14231 VDAC_N.n197 VSS 0.132739f
C14232 VDAC_N.t1835 VSS 0.105768f
C14233 VDAC_N.n198 VSS 0.132739f
C14234 VDAC_N.t1159 VSS 0.105768f
C14235 VDAC_N.n199 VSS 0.132739f
C14236 VDAC_N.t227 VSS 0.105768f
C14237 VDAC_N.n200 VSS 0.132739f
C14238 VDAC_N.t2066 VSS 0.105768f
C14239 VDAC_N.n201 VSS 0.132739f
C14240 VDAC_N.t399 VSS 0.105768f
C14241 VDAC_N.n202 VSS 0.132739f
C14242 VDAC_N.t1967 VSS 0.105768f
C14243 VDAC_N.n203 VSS 0.132739f
C14244 VDAC_N.t1295 VSS 0.105768f
C14245 VDAC_N.n204 VSS 0.132739f
C14246 VDAC_N.t1867 VSS 0.105768f
C14247 VDAC_N.n205 VSS 0.132739f
C14248 VDAC_N.t676 VSS 0.105768f
C14249 VDAC_N.n206 VSS 0.132739f
C14250 VDAC_N.t231 VSS 0.105768f
C14251 VDAC_N.n207 VSS 0.132739f
C14252 VDAC_N.t252 VSS 0.105768f
C14253 VDAC_N.n208 VSS 0.132739f
C14254 VDAC_N.t785 VSS 0.105768f
C14255 VDAC_N.n209 VSS 0.132739f
C14256 VDAC_N.t151 VSS 0.105768f
C14257 VDAC_N.n210 VSS 0.132739f
C14258 VDAC_N.t848 VSS 0.105768f
C14259 VDAC_N.n211 VSS 0.132739f
C14260 VDAC_N.t961 VSS 0.105768f
C14261 VDAC_N.n212 VSS 0.132739f
C14262 VDAC_N.t788 VSS 0.105768f
C14263 VDAC_N.n213 VSS 0.132739f
C14264 VDAC_N.t1330 VSS 0.105768f
C14265 VDAC_N.n214 VSS 0.132739f
C14266 VDAC_N.t1324 VSS 0.105768f
C14267 VDAC_N.n215 VSS 0.132739f
C14268 VDAC_N.t574 VSS 0.105768f
C14269 VDAC_N.n216 VSS 0.132739f
C14270 VDAC_N.t2029 VSS 0.105768f
C14271 VDAC_N.n217 VSS 0.132739f
C14272 VDAC_N.t248 VSS 0.105768f
C14273 VDAC_N.n218 VSS 0.132739f
C14274 VDAC_N.t1830 VSS 0.105768f
C14275 VDAC_N.n219 VSS 0.132739f
C14276 VDAC_N.t640 VSS 0.105768f
C14277 VDAC_N.n220 VSS 0.132739f
C14278 VDAC_N.t1778 VSS 0.105768f
C14279 VDAC_N.n221 VSS 0.132739f
C14280 VDAC_N.t1375 VSS 0.105768f
C14281 VDAC_N.n222 VSS 0.132739f
C14282 VDAC_N.t1334 VSS 0.105768f
C14283 VDAC_N.n223 VSS 0.132739f
C14284 VDAC_N.t591 VSS 0.105768f
C14285 VDAC_N.n224 VSS 0.132739f
C14286 VDAC_N.t1719 VSS 0.105768f
C14287 VDAC_N.n225 VSS 0.132739f
C14288 VDAC_N.t1042 VSS 0.105768f
C14289 VDAC_N.n226 VSS 0.132739f
C14290 VDAC_N.t1507 VSS 0.105768f
C14291 VDAC_N.n227 VSS 0.132739f
C14292 VDAC_N.t934 VSS 0.105768f
C14293 VDAC_N.n228 VSS 0.132739f
C14294 VDAC_N.t715 VSS 0.105768f
C14295 VDAC_N.n229 VSS 0.132739f
C14296 VDAC_N.t945 VSS 0.105768f
C14297 VDAC_N.n230 VSS 0.132739f
C14298 VDAC_N.t1287 VSS 0.105768f
C14299 VDAC_N.n231 VSS 0.132739f
C14300 VDAC_N.t891 VSS 0.105768f
C14301 VDAC_N.n232 VSS 0.132739f
C14302 VDAC_N.t1660 VSS 0.105768f
C14303 VDAC_N.n233 VSS 0.132739f
C14304 VDAC_N.t405 VSS 0.105768f
C14305 VDAC_N.n234 VSS 0.132739f
C14306 VDAC_N.t2101 VSS 0.105768f
C14307 VDAC_N.n235 VSS 0.132739f
C14308 VDAC_N.t1425 VSS 0.105768f
C14309 VDAC_N.n236 VSS 0.132739f
C14310 VDAC_N.t1889 VSS 0.105768f
C14311 VDAC_N.n237 VSS 0.132739f
C14312 VDAC_N.t1208 VSS 0.105768f
C14313 VDAC_N.n238 VSS 0.132739f
C14314 VDAC_N.t1779 VSS 0.105768f
C14315 VDAC_N.n239 VSS 0.132739f
C14316 VDAC_N.t652 VSS 0.105768f
C14317 VDAC_N.n240 VSS 0.132739f
C14318 VDAC_N.t350 VSS 0.105768f
C14319 VDAC_N.n241 VSS 0.132739f
C14320 VDAC_N.t291 VSS 0.105768f
C14321 VDAC_N.n242 VSS 0.12675f
C14322 VDAC_N.t1236 VSS 0.105768f
C14323 VDAC_N.n243 VSS 0.132739f
C14324 VDAC_N.t1470 VSS 0.105768f
C14325 VDAC_N.n244 VSS 0.132739f
C14326 VDAC_N.t1404 VSS 0.105768f
C14327 VDAC_N.n245 VSS 0.132739f
C14328 VDAC_N.t2056 VSS 0.105768f
C14329 VDAC_N.n246 VSS 0.132739f
C14330 VDAC_N.t150 VSS 0.105768f
C14331 VDAC_N.n247 VSS 0.132739f
C14332 VDAC_N.t1632 VSS 0.105768f
C14333 VDAC_N.n248 VSS 0.132739f
C14334 VDAC_N.t1746 VSS 0.105768f
C14335 VDAC_N.n249 VSS 0.132739f
C14336 VDAC_N.t361 VSS 0.105768f
C14337 VDAC_N.n250 VSS 0.132739f
C14338 VDAC_N.t406 VSS 0.105768f
C14339 VDAC_N.n251 VSS 0.132739f
C14340 VDAC_N.t1245 VSS 0.105768f
C14341 VDAC_N.n252 VSS 0.132739f
C14342 VDAC_N.t162 VSS 0.105768f
C14343 VDAC_N.n253 VSS 0.132739f
C14344 VDAC_N.t1133 VSS 0.105768f
C14345 VDAC_N.n254 VSS 0.132739f
C14346 VDAC_N.t421 VSS 0.105768f
C14347 VDAC_N.n255 VSS 0.132739f
C14348 VDAC_N.t484 VSS 0.105768f
C14349 VDAC_N.n256 VSS 0.132739f
C14350 VDAC_N.t714 VSS 0.105768f
C14351 VDAC_N.n257 VSS 0.132739f
C14352 VDAC_N.t343 VSS 0.105768f
C14353 VDAC_N.n258 VSS 0.132739f
C14354 VDAC_N.t1190 VSS 0.105768f
C14355 VDAC_N.n259 VSS 0.132739f
C14356 VDAC_N.t2110 VSS 0.105768f
C14357 VDAC_N.n260 VSS 0.132739f
C14358 VDAC_N.t1647 VSS 0.105768f
C14359 VDAC_N.n261 VSS 0.132739f
C14360 VDAC_N.t146 VSS 0.105768f
C14361 VDAC_N.n262 VSS 0.132739f
C14362 VDAC_N.t203 VSS 0.105768f
C14363 VDAC_N.n263 VSS 0.132739f
C14364 VDAC_N.t1682 VSS 0.105768f
C14365 VDAC_N.n264 VSS 0.132739f
C14366 VDAC_N.t109 VSS 0.105768f
C14367 VDAC_N.n265 VSS 0.132739f
C14368 VDAC_N.t247 VSS 0.105768f
C14369 VDAC_N.n266 VSS 0.132739f
C14370 VDAC_N.t1097 VSS 0.105768f
C14371 VDAC_N.n267 VSS 0.132739f
C14372 VDAC_N.t131 VSS 0.105768f
C14373 VDAC_N.n268 VSS 0.132739f
C14374 VDAC_N.t2133 VSS 0.105768f
C14375 VDAC_N.n269 VSS 0.132739f
C14376 VDAC_N.t1459 VSS 0.105768f
C14377 VDAC_N.n270 VSS 0.132739f
C14378 VDAC_N.t2023 VSS 0.105768f
C14379 VDAC_N.n271 VSS 0.132739f
C14380 VDAC_N.t1357 VSS 0.105768f
C14381 VDAC_N.n272 VSS 0.132739f
C14382 VDAC_N.t919 VSS 0.105768f
C14383 VDAC_N.n273 VSS 0.132739f
C14384 VDAC_N.t244 VSS 0.105768f
C14385 VDAC_N.n274 VSS 0.132739f
C14386 VDAC_N.t867 VSS 0.105768f
C14387 VDAC_N.n275 VSS 0.132739f
C14388 VDAC_N.t412 VSS 0.105768f
C14389 VDAC_N.n276 VSS 0.132739f
C14390 VDAC_N.t144 VSS 0.105768f
C14391 VDAC_N.n277 VSS 0.132739f
C14392 VDAC_N.t1041 VSS 0.105768f
C14393 VDAC_N.n278 VSS 0.132739f
C14394 VDAC_N.t72 VSS 0.105768f
C14395 VDAC_N.n279 VSS 0.132739f
C14396 VDAC_N.t935 VSS 0.105768f
C14397 VDAC_N.n280 VSS 0.132739f
C14398 VDAC_N.t2004 VSS 0.105768f
C14399 VDAC_N.n281 VSS 0.132739f
C14400 VDAC_N.t730 VSS 0.105768f
C14401 VDAC_N.n282 VSS 0.132739f
C14402 VDAC_N.t908 VSS 0.105768f
C14403 VDAC_N.n283 VSS 0.132739f
C14404 VDAC_N.t1390 VSS 0.105768f
C14405 VDAC_N.n284 VSS 0.132739f
C14406 VDAC_N.t601 VSS 0.105768f
C14407 VDAC_N.n285 VSS 0.132739f
C14408 VDAC_N.t960 VSS 0.105768f
C14409 VDAC_N.n286 VSS 0.132739f
C14410 VDAC_N.t962 VSS 0.105768f
C14411 VDAC_N.n287 VSS 0.132739f
C14412 VDAC_N.t1529 VSS 0.105768f
C14413 VDAC_N.n288 VSS 0.132739f
C14414 VDAC_N.t1666 VSS 0.105768f
C14415 VDAC_N.n289 VSS 0.132739f
C14416 VDAC_N.t1317 VSS 0.105768f
C14417 VDAC_N.n290 VSS 0.132739f
C14418 VDAC_N.t382 VSS 0.105768f
C14419 VDAC_N.n291 VSS 0.132739f
C14420 VDAC_N.t1205 VSS 0.105768f
C14421 VDAC_N.n292 VSS 0.132739f
C14422 VDAC_N.t233 VSS 0.105768f
C14423 VDAC_N.n293 VSS 0.132739f
C14424 VDAC_N.t1089 VSS 0.105768f
C14425 VDAC_N.n294 VSS 0.132739f
C14426 VDAC_N.t1559 VSS 0.105768f
C14427 VDAC_N.n295 VSS 0.132739f
C14428 VDAC_N.t2015 VSS 0.105768f
C14429 VDAC_N.n296 VSS 0.132739f
C14430 VDAC_N.t689 VSS 0.105768f
C14431 VDAC_N.n297 VSS 0.132739f
C14432 VDAC_N.t1909 VSS 0.105768f
C14433 VDAC_N.n298 VSS 0.132739f
C14434 VDAC_N.t1233 VSS 0.105768f
C14435 VDAC_N.n299 VSS 0.132739f
C14436 VDAC_N.t1703 VSS 0.105768f
C14437 VDAC_N.n300 VSS 0.132739f
C14438 VDAC_N.t812 VSS 0.105768f
C14439 VDAC_N.n301 VSS 0.132739f
C14440 VDAC_N.t1591 VSS 0.105768f
C14441 VDAC_N.n302 VSS 0.132739f
C14442 VDAC_N.t533 VSS 0.105768f
C14443 VDAC_N.n303 VSS 0.132739f
C14444 VDAC_N.t1856 VSS 0.105768f
C14445 VDAC_N.n304 VSS 0.132739f
C14446 VDAC_N.t983 VSS 0.105768f
C14447 VDAC_N.n305 VSS 0.12675f
C14448 VDAC_N.t1305 VSS 0.105768f
C14449 VDAC_N.n306 VSS 0.132739f
C14450 VDAC_N.t489 VSS 0.105768f
C14451 VDAC_N.n307 VSS 0.132739f
C14452 VDAC_N.t319 VSS 0.105768f
C14453 VDAC_N.n308 VSS 0.132739f
C14454 VDAC_N.t1659 VSS 0.105768f
C14455 VDAC_N.n309 VSS 0.132739f
C14456 VDAC_N.t2115 VSS 0.105768f
C14457 VDAC_N.n310 VSS 0.132739f
C14458 VDAC_N.t787 VSS 0.105768f
C14459 VDAC_N.n311 VSS 0.132739f
C14460 VDAC_N.t1015 VSS 0.105768f
C14461 VDAC_N.n312 VSS 0.132739f
C14462 VDAC_N.t1264 VSS 0.105768f
C14463 VDAC_N.n313 VSS 0.132739f
C14464 VDAC_N.t1899 VSS 0.105768f
C14465 VDAC_N.n314 VSS 0.132739f
C14466 VDAC_N.t420 VSS 0.105768f
C14467 VDAC_N.n315 VSS 0.132739f
C14468 VDAC_N.t1693 VSS 0.105768f
C14469 VDAC_N.n316 VSS 0.132739f
C14470 VDAC_N.t1420 VSS 0.105768f
C14471 VDAC_N.n317 VSS 0.132739f
C14472 VDAC_N.t1134 VSS 0.105768f
C14473 VDAC_N.n318 VSS 0.132739f
C14474 VDAC_N.t986 VSS 0.105768f
C14475 VDAC_N.n319 VSS 0.132739f
C14476 VDAC_N.t735 VSS 0.105768f
C14477 VDAC_N.n320 VSS 0.132739f
C14478 VDAC_N.t275 VSS 0.105768f
C14479 VDAC_N.n321 VSS 0.132739f
C14480 VDAC_N.t683 VSS 0.105768f
C14481 VDAC_N.n322 VSS 0.132739f
C14482 VDAC_N.t911 VSS 0.105768f
C14483 VDAC_N.n323 VSS 0.132739f
C14484 VDAC_N.t1620 VSS 0.105768f
C14485 VDAC_N.n324 VSS 0.132739f
C14486 VDAC_N.t861 VSS 0.105768f
C14487 VDAC_N.n325 VSS 0.132739f
C14488 VDAC_N.t2118 VSS 0.105768f
C14489 VDAC_N.n326 VSS 0.132739f
C14490 VDAC_N.t1577 VSS 0.105768f
C14491 VDAC_N.n327 VSS 0.132739f
C14492 VDAC_N.t2039 VSS 0.105768f
C14493 VDAC_N.n328 VSS 0.132739f
C14494 VDAC_N.t1368 VSS 0.105768f
C14495 VDAC_N.n329 VSS 0.132739f
C14496 VDAC_N.t1823 VSS 0.105768f
C14497 VDAC_N.n330 VSS 0.132739f
C14498 VDAC_N.t948 VSS 0.105768f
C14499 VDAC_N.n331 VSS 0.132739f
C14500 VDAC_N.t718 VSS 0.105768f
C14501 VDAC_N.n332 VSS 0.132739f
C14502 VDAC_N.t290 VSS 0.105768f
C14503 VDAC_N.n333 VSS 0.132739f
C14504 VDAC_N.t1194 VSS 0.105768f
C14505 VDAC_N.n334 VSS 0.132739f
C14506 VDAC_N.t283 VSS 0.105768f
C14507 VDAC_N.n335 VSS 0.132739f
C14508 VDAC_N.t752 VSS 0.105768f
C14509 VDAC_N.n336 VSS 0.132739f
C14510 VDAC_N.t974 VSS 0.105768f
C14511 VDAC_N.n337 VSS 0.132739f
C14512 VDAC_N.t548 VSS 0.105768f
C14513 VDAC_N.n338 VSS 0.132739f
C14514 VDAC_N.t746 VSS 0.105768f
C14515 VDAC_N.n339 VSS 0.132739f
C14516 VDAC_N.t1217 VSS 0.105768f
C14517 VDAC_N.n340 VSS 0.132739f
C14518 VDAC_N.t1250 VSS 0.105768f
C14519 VDAC_N.n341 VSS 0.132739f
C14520 VDAC_N.t565 VSS 0.105768f
C14521 VDAC_N.n342 VSS 0.132739f
C14522 VDAC_N.t824 VSS 0.105768f
C14523 VDAC_N.n343 VSS 0.132739f
C14524 VDAC_N.t1974 VSS 0.105768f
C14525 VDAC_N.n344 VSS 0.132739f
C14526 VDAC_N.t1461 VSS 0.105768f
C14527 VDAC_N.n345 VSS 0.132739f
C14528 VDAC_N.t1698 VSS 0.105768f
C14529 VDAC_N.n346 VSS 0.132739f
C14530 VDAC_N.t39 VSS 0.105768f
C14531 VDAC_N.n347 VSS 0.132739f
C14532 VDAC_N.t1897 VSS 0.105768f
C14533 VDAC_N.n348 VSS 0.132739f
C14534 VDAC_N.t177 VSS 0.105768f
C14535 VDAC_N.n349 VSS 0.132739f
C14536 VDAC_N.t1685 VSS 0.105768f
C14537 VDAC_N.n350 VSS 0.132739f
C14538 VDAC_N.t364 VSS 0.105768f
C14539 VDAC_N.n351 VSS 0.132739f
C14540 VDAC_N.t799 VSS 0.105768f
C14541 VDAC_N.n352 VSS 0.132739f
C14542 VDAC_N.t2033 VSS 0.105768f
C14543 VDAC_N.n353 VSS 0.132739f
C14544 VDAC_N.t1465 VSS 0.105768f
C14545 VDAC_N.n354 VSS 0.132739f
C14546 VDAC_N.t1923 VSS 0.105768f
C14547 VDAC_N.n355 VSS 0.132739f
C14548 VDAC_N.t84 VSS 0.105768f
C14549 VDAC_N.n356 VSS 0.132739f
C14550 VDAC_N.t1815 VSS 0.105768f
C14551 VDAC_N.n357 VSS 0.132739f
C14552 VDAC_N.t1836 VSS 0.105768f
C14553 VDAC_N.n358 VSS 0.132739f
C14554 VDAC_N.t1182 VSS 0.105768f
C14555 VDAC_N.n359 VSS 0.132739f
C14556 VDAC_N.t2061 VSS 0.105768f
C14557 VDAC_N.n360 VSS 0.132739f
C14558 VDAC_N.t968 VSS 0.105768f
C14559 VDAC_N.n361 VSS 0.132739f
C14560 VDAC_N.t987 VSS 0.105768f
C14561 VDAC_N.n362 VSS 0.132739f
C14562 VDAC_N.t36 VSS 0.105768f
C14563 VDAC_N.n363 VSS 0.132739f
C14564 VDAC_N.t234 VSS 0.105768f
C14565 VDAC_N.n364 VSS 0.132739f
C14566 VDAC_N.t596 VSS 0.105768f
C14567 VDAC_N.n365 VSS 0.132739f
C14568 VDAC_N.t1246 VSS 0.105768f
C14569 VDAC_N.n366 VSS 0.132739f
C14570 VDAC_N.t619 VSS 0.105768f
C14571 VDAC_N.n367 VSS 0.132739f
C14572 VDAC_N.t1032 VSS 0.105768f
C14573 VDAC_N.n368 VSS 0.12675f
C14574 VDAC_N.t2008 VSS 0.105768f
C14575 VDAC_N.n369 VSS 0.132739f
C14576 VDAC_N.t557 VSS 0.105768f
C14577 VDAC_N.n370 VSS 0.132739f
C14578 VDAC_N.t40 VSS 0.105768f
C14579 VDAC_N.n371 VSS 0.132739f
C14580 VDAC_N.t878 VSS 0.105768f
C14581 VDAC_N.n372 VSS 0.132739f
C14582 VDAC_N.t687 VSS 0.105768f
C14583 VDAC_N.n373 VSS 0.132739f
C14584 VDAC_N.t770 VSS 0.105768f
C14585 VDAC_N.n374 VSS 0.132739f
C14586 VDAC_N.t629 VSS 0.105768f
C14587 VDAC_N.n375 VSS 0.132739f
C14588 VDAC_N.t1699 VSS 0.105768f
C14589 VDAC_N.n376 VSS 0.132739f
C14590 VDAC_N.t575 VSS 0.105768f
C14591 VDAC_N.n377 VSS 0.132739f
C14592 VDAC_N.t807 VSS 0.105768f
C14593 VDAC_N.n378 VSS 0.132739f
C14594 VDAC_N.t910 VSS 0.105768f
C14595 VDAC_N.n379 VSS 0.132739f
C14596 VDAC_N.t751 VSS 0.105768f
C14597 VDAC_N.n380 VSS 0.132739f
C14598 VDAC_N.t1933 VSS 0.105768f
C14599 VDAC_N.n381 VSS 0.132739f
C14600 VDAC_N.t790 VSS 0.105768f
C14601 VDAC_N.n382 VSS 0.132739f
C14602 VDAC_N.t1249 VSS 0.105768f
C14603 VDAC_N.n383 VSS 0.132739f
C14604 VDAC_N.t1817 VSS 0.105768f
C14605 VDAC_N.n384 VSS 0.132739f
C14606 VDAC_N.t167 VSS 0.105768f
C14607 VDAC_N.n385 VSS 0.132739f
C14608 VDAC_N.t1605 VSS 0.105768f
C14609 VDAC_N.n386 VSS 0.132739f
C14610 VDAC_N.t18 VSS 0.105768f
C14611 VDAC_N.n387 VSS 0.132739f
C14612 VDAC_N.t1495 VSS 0.105768f
C14613 VDAC_N.n388 VSS 0.132739f
C14614 VDAC_N.t1949 VSS 0.105768f
C14615 VDAC_N.n389 VSS 0.132739f
C14616 VDAC_N.t1389 VSS 0.105768f
C14617 VDAC_N.n390 VSS 0.132739f
C14618 VDAC_N.t1853 VSS 0.105768f
C14619 VDAC_N.n391 VSS 0.132739f
C14620 VDAC_N.t1172 VSS 0.105768f
C14621 VDAC_N.n392 VSS 0.132739f
C14622 VDAC_N.t831 VSS 0.105768f
C14623 VDAC_N.n393 VSS 0.132739f
C14624 VDAC_N.t1212 VSS 0.105768f
C14625 VDAC_N.n394 VSS 0.132739f
C14626 VDAC_N.t2040 VSS 0.105768f
C14627 VDAC_N.n395 VSS 0.132739f
C14628 VDAC_N.t1005 VSS 0.105768f
C14629 VDAC_N.n396 VSS 0.132739f
C14630 VDAC_N.t1600 VSS 0.105768f
C14631 VDAC_N.n397 VSS 0.132739f
C14632 VDAC_N.t1883 VSS 0.105768f
C14633 VDAC_N.n398 VSS 0.132739f
C14634 VDAC_N.t1428 VSS 0.105768f
C14635 VDAC_N.n399 VSS 0.132739f
C14636 VDAC_N.t778 VSS 0.105768f
C14637 VDAC_N.n400 VSS 0.132739f
C14638 VDAC_N.t588 VSS 0.105768f
C14639 VDAC_N.n401 VSS 0.132739f
C14640 VDAC_N.t1090 VSS 0.105768f
C14641 VDAC_N.n402 VSS 0.132739f
C14642 VDAC_N.t1026 VSS 0.105768f
C14643 VDAC_N.n403 VSS 0.132739f
C14644 VDAC_N.t1728 VSS 0.105768f
C14645 VDAC_N.n404 VSS 0.132739f
C14646 VDAC_N.t1806 VSS 0.105768f
C14647 VDAC_N.n405 VSS 0.132739f
C14648 VDAC_N.t436 VSS 0.105768f
C14649 VDAC_N.n406 VSS 0.132739f
C14650 VDAC_N.t810 VSS 0.105768f
C14651 VDAC_N.n407 VSS 0.132739f
C14652 VDAC_N.t183 VSS 0.105768f
C14653 VDAC_N.n408 VSS 0.132739f
C14654 VDAC_N.t666 VSS 0.105768f
C14655 VDAC_N.n409 VSS 0.132739f
C14656 VDAC_N.t1243 VSS 0.105768f
C14657 VDAC_N.n410 VSS 0.132739f
C14658 VDAC_N.t1707 VSS 0.105768f
C14659 VDAC_N.n411 VSS 0.132739f
C14660 VDAC_N.t278 VSS 0.105768f
C14661 VDAC_N.n412 VSS 0.132739f
C14662 VDAC_N.t1489 VSS 0.105768f
C14663 VDAC_N.n413 VSS 0.132739f
C14664 VDAC_N.t535 VSS 0.105768f
C14665 VDAC_N.n414 VSS 0.132739f
C14666 VDAC_N.t1383 VSS 0.105768f
C14667 VDAC_N.n415 VSS 0.132739f
C14668 VDAC_N.t937 VSS 0.105768f
C14669 VDAC_N.n416 VSS 0.132739f
C14670 VDAC_N.t339 VSS 0.105768f
C14671 VDAC_N.n417 VSS 0.132739f
C14672 VDAC_N.t1735 VSS 0.105768f
C14673 VDAC_N.n418 VSS 0.132739f
C14674 VDAC_N.t92 VSS 0.105768f
C14675 VDAC_N.n419 VSS 0.132739f
C14676 VDAC_N.t1627 VSS 0.105768f
C14677 VDAC_N.n420 VSS 0.132739f
C14678 VDAC_N.t543 VSS 0.105768f
C14679 VDAC_N.n421 VSS 0.132739f
C14680 VDAC_N.t800 VSS 0.105768f
C14681 VDAC_N.n422 VSS 0.132739f
C14682 VDAC_N.t259 VSS 0.105768f
C14683 VDAC_N.n423 VSS 0.132739f
C14684 VDAC_N.t1136 VSS 0.105768f
C14685 VDAC_N.n424 VSS 0.132739f
C14686 VDAC_N.t895 VSS 0.105768f
C14687 VDAC_N.n425 VSS 0.132739f
C14688 VDAC_N.t1100 VSS 0.105768f
C14689 VDAC_N.n426 VSS 0.132739f
C14690 VDAC_N.t1286 VSS 0.105768f
C14691 VDAC_N.n427 VSS 0.132739f
C14692 VDAC_N.t2117 VSS 0.105768f
C14693 VDAC_N.n428 VSS 0.132739f
C14694 VDAC_N.t1712 VSS 0.105768f
C14695 VDAC_N.n429 VSS 0.132739f
C14696 VDAC_N.t2010 VSS 0.105768f
C14697 VDAC_N.n430 VSS 0.132739f
C14698 VDAC_N.t1272 VSS 0.105768f
C14699 VDAC_N.n431 VSS 0.12675f
C14700 VDAC_N.t837 VSS 0.105768f
C14701 VDAC_N.n432 VSS 0.132739f
C14702 VDAC_N.t1468 VSS 0.105768f
C14703 VDAC_N.n433 VSS 0.132739f
C14704 VDAC_N.t781 VSS 0.105768f
C14705 VDAC_N.n434 VSS 0.132739f
C14706 VDAC_N.t1991 VSS 0.105768f
C14707 VDAC_N.n435 VSS 0.132739f
C14708 VDAC_N.t176 VSS 0.105768f
C14709 VDAC_N.n436 VSS 0.132739f
C14710 VDAC_N.t493 VSS 0.105768f
C14711 VDAC_N.n437 VSS 0.132739f
C14712 VDAC_N.t1476 VSS 0.105768f
C14713 VDAC_N.n438 VSS 0.132739f
C14714 VDAC_N.t1318 VSS 0.105768f
C14715 VDAC_N.n439 VSS 0.132739f
C14716 VDAC_N.t1228 VSS 0.105768f
C14717 VDAC_N.n440 VSS 0.132739f
C14718 VDAC_N.t566 VSS 0.105768f
C14719 VDAC_N.n441 VSS 0.132739f
C14720 VDAC_N.t527 VSS 0.105768f
C14721 VDAC_N.n442 VSS 0.132739f
C14722 VDAC_N.t888 VSS 0.105768f
C14723 VDAC_N.n443 VSS 0.132739f
C14724 VDAC_N.t922 VSS 0.105768f
C14725 VDAC_N.n444 VSS 0.132739f
C14726 VDAC_N.t1511 VSS 0.105768f
C14727 VDAC_N.n445 VSS 0.132739f
C14728 VDAC_N.t1963 VSS 0.105768f
C14729 VDAC_N.n446 VSS 0.132739f
C14730 VDAC_N.t400 VSS 0.105768f
C14731 VDAC_N.n447 VSS 0.132739f
C14732 VDAC_N.t1865 VSS 0.105768f
C14733 VDAC_N.n448 VSS 0.132739f
C14734 VDAC_N.t660 VSS 0.105768f
C14735 VDAC_N.n449 VSS 0.132739f
C14736 VDAC_N.t1482 VSS 0.105768f
C14737 VDAC_N.n450 VSS 0.132739f
C14738 VDAC_N.t892 VSS 0.105768f
C14739 VDAC_N.n451 VSS 0.132739f
C14740 VDAC_N.t2080 VSS 0.105768f
C14741 VDAC_N.n452 VSS 0.132739f
C14742 VDAC_N.t2103 VSS 0.105768f
C14743 VDAC_N.n453 VSS 0.132739f
C14744 VDAC_N.t232 VSS 0.105768f
C14745 VDAC_N.n454 VSS 0.132739f
C14746 VDAC_N.t462 VSS 0.105768f
C14747 VDAC_N.n455 VSS 0.132739f
C14748 VDAC_N.t404 VSS 0.105768f
C14749 VDAC_N.n456 VSS 0.132739f
C14750 VDAC_N.t410 VSS 0.105768f
C14751 VDAC_N.n457 VSS 0.132739f
C14752 VDAC_N.t1253 VSS 0.105768f
C14753 VDAC_N.n458 VSS 0.132739f
C14754 VDAC_N.t1114 VSS 0.105768f
C14755 VDAC_N.n459 VSS 0.132739f
C14756 VDAC_N.t585 VSS 0.105768f
C14757 VDAC_N.n460 VSS 0.132739f
C14758 VDAC_N.t1784 VSS 0.105768f
C14759 VDAC_N.n461 VSS 0.132739f
C14760 VDAC_N.t1826 VSS 0.105768f
C14761 VDAC_N.n462 VSS 0.132739f
C14762 VDAC_N.t1497 VSS 0.105768f
C14763 VDAC_N.n463 VSS 0.132739f
C14764 VDAC_N.t822 VSS 0.105768f
C14765 VDAC_N.n464 VSS 0.132739f
C14766 VDAC_N.t1281 VSS 0.105768f
C14767 VDAC_N.n465 VSS 0.132739f
C14768 VDAC_N.t1747 VSS 0.105768f
C14769 VDAC_N.n466 VSS 0.132739f
C14770 VDAC_N.t1171 VSS 0.105768f
C14771 VDAC_N.n467 VSS 0.132739f
C14772 VDAC_N.t1639 VSS 0.105768f
C14773 VDAC_N.n468 VSS 0.132739f
C14774 VDAC_N.t1890 VSS 0.105768f
C14775 VDAC_N.n469 VSS 0.132739f
C14776 VDAC_N.t777 VSS 0.105768f
C14777 VDAC_N.n470 VSS 0.132739f
C14778 VDAC_N.t1007 VSS 0.105768f
C14779 VDAC_N.n471 VSS 0.132739f
C14780 VDAC_N.t371 VSS 0.105768f
C14781 VDAC_N.n472 VSS 0.132739f
C14782 VDAC_N.t1953 VSS 0.105768f
C14783 VDAC_N.n473 VSS 0.132739f
C14784 VDAC_N.t1076 VSS 0.105768f
C14785 VDAC_N.n474 VSS 0.132739f
C14786 VDAC_N.t1751 VSS 0.105768f
C14787 VDAC_N.n475 VSS 0.132739f
C14788 VDAC_N.t1532 VSS 0.105768f
C14789 VDAC_N.n476 VSS 0.132739f
C14790 VDAC_N.t642 VSS 0.105768f
C14791 VDAC_N.n477 VSS 0.132739f
C14792 VDAC_N.t545 VSS 0.105768f
C14793 VDAC_N.n478 VSS 0.132739f
C14794 VDAC_N.t432 VSS 0.105768f
C14795 VDAC_N.n479 VSS 0.132739f
C14796 VDAC_N.t1989 VSS 0.105768f
C14797 VDAC_N.n480 VSS 0.132739f
C14798 VDAC_N.t320 VSS 0.105768f
C14799 VDAC_N.n481 VSS 0.132739f
C14800 VDAC_N.t1546 VSS 0.105768f
C14801 VDAC_N.n482 VSS 0.132739f
C14802 VDAC_N.t1460 VSS 0.105768f
C14803 VDAC_N.n483 VSS 0.132739f
C14804 VDAC_N.t1310 VSS 0.105768f
C14805 VDAC_N.n484 VSS 0.132739f
C14806 VDAC_N.t1137 VSS 0.105768f
C14807 VDAC_N.n485 VSS 0.132739f
C14808 VDAC_N.t1760 VSS 0.105768f
C14809 VDAC_N.n486 VSS 0.132739f
C14810 VDAC_N.t530 VSS 0.105768f
C14811 VDAC_N.n487 VSS 0.132739f
C14812 VDAC_N.t48 VSS 0.105768f
C14813 VDAC_N.n488 VSS 0.132739f
C14814 VDAC_N.t1610 VSS 0.105768f
C14815 VDAC_N.n489 VSS 0.132739f
C14816 VDAC_N.t113 VSS 0.105768f
C14817 VDAC_N.n490 VSS 0.132739f
C14818 VDAC_N.t1366 VSS 0.105768f
C14819 VDAC_N.n491 VSS 0.132739f
C14820 VDAC_N.t599 VSS 0.105768f
C14821 VDAC_N.n492 VSS 0.132739f
C14822 VDAC_N.t883 VSS 0.105768f
C14823 VDAC_N.n493 VSS 0.132739f
C14824 VDAC_N.t2090 VSS 0.105768f
C14825 VDAC_N.n494 VSS 0.12675f
C14826 VDAC_N.t446 VSS 0.105768f
C14827 VDAC_N.n495 VSS 0.132739f
C14828 VDAC_N.t1435 VSS 0.105768f
C14829 VDAC_N.n496 VSS 0.132739f
C14830 VDAC_N.t1474 VSS 0.105768f
C14831 VDAC_N.n497 VSS 0.132739f
C14832 VDAC_N.t1221 VSS 0.105768f
C14833 VDAC_N.n498 VSS 0.132739f
C14834 VDAC_N.t857 VSS 0.105768f
C14835 VDAC_N.n499 VSS 0.132739f
C14836 VDAC_N.t1107 VSS 0.105768f
C14837 VDAC_N.n500 VSS 0.132739f
C14838 VDAC_N.t1569 VSS 0.105768f
C14839 VDAC_N.n501 VSS 0.132739f
C14840 VDAC_N.t2035 VSS 0.105768f
C14841 VDAC_N.n502 VSS 0.132739f
C14842 VDAC_N.t387 VSS 0.105768f
C14843 VDAC_N.n503 VSS 0.132739f
C14844 VDAC_N.t975 VSS 0.105768f
C14845 VDAC_N.n504 VSS 0.132739f
C14846 VDAC_N.t333 VSS 0.105768f
C14847 VDAC_N.n505 VSS 0.132739f
C14848 VDAC_N.t475 VSS 0.105768f
C14849 VDAC_N.n506 VSS 0.132739f
C14850 VDAC_N.t140 VSS 0.105768f
C14851 VDAC_N.n507 VSS 0.132739f
C14852 VDAC_N.t1323 VSS 0.105768f
C14853 VDAC_N.n508 VSS 0.132739f
C14854 VDAC_N.t903 VSS 0.105768f
C14855 VDAC_N.n509 VSS 0.132739f
C14856 VDAC_N.t388 VSS 0.105768f
C14857 VDAC_N.n510 VSS 0.132739f
C14858 VDAC_N.t851 VSS 0.105768f
C14859 VDAC_N.n511 VSS 0.132739f
C14860 VDAC_N.t2131 VSS 0.105768f
C14861 VDAC_N.n512 VSS 0.132739f
C14862 VDAC_N.t1098 VSS 0.105768f
C14863 VDAC_N.n513 VSS 0.132739f
C14864 VDAC_N.t2021 VSS 0.105768f
C14865 VDAC_N.n514 VSS 0.132739f
C14866 VDAC_N.t672 VSS 0.105768f
C14867 VDAC_N.n515 VSS 0.132739f
C14868 VDAC_N.t1913 VSS 0.105768f
C14869 VDAC_N.n516 VSS 0.132739f
C14870 VDAC_N.t1748 VSS 0.105768f
C14871 VDAC_N.n517 VSS 0.132739f
C14872 VDAC_N.t1370 VSS 0.105768f
C14873 VDAC_N.n518 VSS 0.132739f
C14874 VDAC_N.t924 VSS 0.105768f
C14875 VDAC_N.n519 VSS 0.132739f
C14876 VDAC_N.t594 VSS 0.105768f
C14877 VDAC_N.n520 VSS 0.132739f
C14878 VDAC_N.t286 VSS 0.105768f
C14879 VDAC_N.n521 VSS 0.132739f
C14880 VDAC_N.t1424 VSS 0.105768f
C14881 VDAC_N.n522 VSS 0.132739f
C14882 VDAC_N.t1874 VSS 0.105768f
C14883 VDAC_N.n523 VSS 0.132739f
C14884 VDAC_N.t1988 VSS 0.105768f
C14885 VDAC_N.n524 VSS 0.132739f
C14886 VDAC_N.t378 VSS 0.105768f
C14887 VDAC_N.n525 VSS 0.132739f
C14888 VDAC_N.t1309 VSS 0.105768f
C14889 VDAC_N.n526 VSS 0.132739f
C14890 VDAC_N.t1222 VSS 0.105768f
C14891 VDAC_N.n527 VSS 0.132739f
C14892 VDAC_N.t1083 VSS 0.105768f
C14893 VDAC_N.n528 VSS 0.132739f
C14894 VDAC_N.t791 VSS 0.105768f
C14895 VDAC_N.n529 VSS 0.132739f
C14896 VDAC_N.t58 VSS 0.105768f
C14897 VDAC_N.n530 VSS 0.132739f
C14898 VDAC_N.t1447 VSS 0.105768f
C14899 VDAC_N.n531 VSS 0.132739f
C14900 VDAC_N.t74 VSS 0.105768f
C14901 VDAC_N.n532 VSS 0.132739f
C14902 VDAC_N.t1341 VSS 0.105768f
C14903 VDAC_N.n533 VSS 0.132739f
C14904 VDAC_N.t913 VSS 0.105768f
C14905 VDAC_N.n534 VSS 0.132739f
C14906 VDAC_N.t1203 VSS 0.105768f
C14907 VDAC_N.n535 VSS 0.132739f
C14908 VDAC_N.t899 VSS 0.105768f
C14909 VDAC_N.n536 VSS 0.132739f
C14910 VDAC_N.t172 VSS 0.105768f
C14911 VDAC_N.n537 VSS 0.132739f
C14912 VDAC_N.t219 VSS 0.105768f
C14913 VDAC_N.n538 VSS 0.132739f
C14914 VDAC_N.t2013 VSS 0.105768f
C14915 VDAC_N.n539 VSS 0.132739f
C14916 VDAC_N.t1736 VSS 0.105768f
C14917 VDAC_N.n540 VSS 0.132739f
C14918 VDAC_N.t1905 VSS 0.105768f
C14919 VDAC_N.n541 VSS 0.132739f
C14920 VDAC_N.t132 VSS 0.105768f
C14921 VDAC_N.n542 VSS 0.132739f
C14922 VDAC_N.t915 VSS 0.105768f
C14923 VDAC_N.n543 VSS 0.132739f
C14924 VDAC_N.t1580 VSS 0.105768f
C14925 VDAC_N.n544 VSS 0.132739f
C14926 VDAC_N.t1150 VSS 0.105768f
C14927 VDAC_N.n545 VSS 0.132739f
C14928 VDAC_N.t220 VSS 0.105768f
C14929 VDAC_N.n546 VSS 0.132739f
C14930 VDAC_N.t256 VSS 0.105768f
C14931 VDAC_N.n547 VSS 0.132739f
C14932 VDAC_N.t946 VSS 0.105768f
C14933 VDAC_N.n548 VSS 0.132739f
C14934 VDAC_N.t980 VSS 0.105768f
C14935 VDAC_N.n549 VSS 0.132739f
C14936 VDAC_N.t230 VSS 0.105768f
C14937 VDAC_N.n550 VSS 0.132739f
C14938 VDAC_N.t1996 VSS 0.105768f
C14939 VDAC_N.n551 VSS 0.132739f
C14940 VDAC_N.t1214 VSS 0.105768f
C14941 VDAC_N.n552 VSS 0.132739f
C14942 VDAC_N.t1191 VSS 0.105768f
C14943 VDAC_N.n553 VSS 0.132739f
C14944 VDAC_N.t512 VSS 0.105768f
C14945 VDAC_N.n554 VSS 0.132739f
C14946 VDAC_N.t506 VSS 0.105768f
C14947 VDAC_N.n555 VSS 0.132739f
C14948 VDAC_N.t1545 VSS 0.105768f
C14949 VDAC_N.n556 VSS 0.132739f
C14950 VDAC_N.t1710 VSS 0.105768f
C14951 VDAC_N.n557 VSS 0.12675f
C14952 VDAC_N.t2044 VSS 0.105768f
C14953 VDAC_N.n558 VSS 0.132739f
C14954 VDAC_N.t1282 VSS 0.105768f
C14955 VDAC_N.n559 VSS 0.132739f
C14956 VDAC_N.t549 VSS 0.105768f
C14957 VDAC_N.n560 VSS 0.132739f
C14958 VDAC_N.t80 VSS 0.105768f
C14959 VDAC_N.n561 VSS 0.132739f
C14960 VDAC_N.t466 VSS 0.105768f
C14961 VDAC_N.n562 VSS 0.132739f
C14962 VDAC_N.t1248 VSS 0.105768f
C14963 VDAC_N.n563 VSS 0.132739f
C14964 VDAC_N.t1570 VSS 0.105768f
C14965 VDAC_N.n564 VSS 0.132739f
C14966 VDAC_N.t1259 VSS 0.105768f
C14967 VDAC_N.n565 VSS 0.132739f
C14968 VDAC_N.t354 VSS 0.105768f
C14969 VDAC_N.n566 VSS 0.132739f
C14970 VDAC_N.t589 VSS 0.105768f
C14971 VDAC_N.n567 VSS 0.132739f
C14972 VDAC_N.t1808 VSS 0.105768f
C14973 VDAC_N.n568 VSS 0.132739f
C14974 VDAC_N.t2050 VSS 0.105768f
C14975 VDAC_N.n569 VSS 0.132739f
C14976 VDAC_N.t1503 VSS 0.105768f
C14977 VDAC_N.n570 VSS 0.132739f
C14978 VDAC_N.t165 VSS 0.105768f
C14979 VDAC_N.n571 VSS 0.132739f
C14980 VDAC_N.t1589 VSS 0.105768f
C14981 VDAC_N.n572 VSS 0.132739f
C14982 VDAC_N.t1500 VSS 0.105768f
C14983 VDAC_N.n573 VSS 0.132739f
C14984 VDAC_N.t1477 VSS 0.105768f
C14985 VDAC_N.n574 VSS 0.132739f
C14986 VDAC_N.t505 VSS 0.105768f
C14987 VDAC_N.n575 VSS 0.132739f
C14988 VDAC_N.t1400 VSS 0.105768f
C14989 VDAC_N.n576 VSS 0.132739f
C14990 VDAC_N.t931 VSS 0.105768f
C14991 VDAC_N.n577 VSS 0.132739f
C14992 VDAC_N.t1036 VSS 0.105768f
C14993 VDAC_N.n578 VSS 0.132739f
C14994 VDAC_N.t1723 VSS 0.105768f
C14995 VDAC_N.n579 VSS 0.132739f
C14996 VDAC_N.t26 VSS 0.105768f
C14997 VDAC_N.n580 VSS 0.132739f
C14998 VDAC_N.t1968 VSS 0.105768f
C14999 VDAC_N.n581 VSS 0.132739f
C15000 VDAC_N.t149 VSS 0.105768f
C15001 VDAC_N.n582 VSS 0.132739f
C15002 VDAC_N.t1520 VSS 0.105768f
C15003 VDAC_N.n583 VSS 0.132739f
C15004 VDAC_N.t870 VSS 0.105768f
C15005 VDAC_N.n584 VSS 0.132739f
C15006 VDAC_N.t1300 VSS 0.105768f
C15007 VDAC_N.n585 VSS 0.132739f
C15008 VDAC_N.t210 VSS 0.105768f
C15009 VDAC_N.n586 VSS 0.132739f
C15010 VDAC_N.t1788 VSS 0.105768f
C15011 VDAC_N.n587 VSS 0.132739f
C15012 VDAC_N.t2088 VSS 0.105768f
C15013 VDAC_N.n588 VSS 0.132739f
C15014 VDAC_N.t569 VSS 0.105768f
C15015 VDAC_N.n589 VSS 0.132739f
C15016 VDAC_N.t1664 VSS 0.105768f
C15017 VDAC_N.n590 VSS 0.132739f
C15018 VDAC_N.t1766 VSS 0.105768f
C15019 VDAC_N.n591 VSS 0.132739f
C15020 VDAC_N.t1369 VSS 0.105768f
C15021 VDAC_N.n592 VSS 0.132739f
C15022 VDAC_N.t1558 VSS 0.105768f
C15023 VDAC_N.n593 VSS 0.132739f
C15024 VDAC_N.t641 VSS 0.105768f
C15025 VDAC_N.n594 VSS 0.132739f
C15026 VDAC_N.t62 VSS 0.105768f
C15027 VDAC_N.n595 VSS 0.132739f
C15028 VDAC_N.t1143 VSS 0.105768f
C15029 VDAC_N.n596 VSS 0.132739f
C15030 VDAC_N.t423 VSS 0.105768f
C15031 VDAC_N.n597 VSS 0.132739f
C15032 VDAC_N.t2006 VSS 0.105768f
C15033 VDAC_N.n598 VSS 0.132739f
C15034 VDAC_N.t417 VSS 0.105768f
C15035 VDAC_N.n599 VSS 0.132739f
C15036 VDAC_N.t1035 VSS 0.105768f
C15037 VDAC_N.n600 VSS 0.132739f
C15038 VDAC_N.t701 VSS 0.105768f
C15039 VDAC_N.n601 VSS 0.132739f
C15040 VDAC_N.t1829 VSS 0.105768f
C15041 VDAC_N.n602 VSS 0.132739f
C15042 VDAC_N.t260 VSS 0.105768f
C15043 VDAC_N.n603 VSS 0.132739f
C15044 VDAC_N.t1717 VSS 0.105768f
C15045 VDAC_N.n604 VSS 0.132739f
C15046 VDAC_N.t24 VSS 0.105768f
C15047 VDAC_N.n605 VSS 0.132739f
C15048 VDAC_N.t127 VSS 0.105768f
C15049 VDAC_N.n606 VSS 0.132739f
C15050 VDAC_N.t2071 VSS 0.105768f
C15051 VDAC_N.n607 VSS 0.132739f
C15052 VDAC_N.t1496 VSS 0.105768f
C15053 VDAC_N.n608 VSS 0.132739f
C15054 VDAC_N.t1955 VSS 0.105768f
C15055 VDAC_N.n609 VSS 0.132739f
C15056 VDAC_N.t2132 VSS 0.105768f
C15057 VDAC_N.n610 VSS 0.132739f
C15058 VDAC_N.t750 VSS 0.105768f
C15059 VDAC_N.n611 VSS 0.132739f
C15060 VDAC_N.t1596 VSS 0.105768f
C15061 VDAC_N.n612 VSS 0.132739f
C15062 VDAC_N.t1258 VSS 0.105768f
C15063 VDAC_N.n613 VSS 0.132739f
C15064 VDAC_N.t287 VSS 0.105768f
C15065 VDAC_N.n614 VSS 0.132739f
C15066 VDAC_N.t840 VSS 0.105768f
C15067 VDAC_N.n615 VSS 0.132739f
C15068 VDAC_N.t1978 VSS 0.105768f
C15069 VDAC_N.n616 VSS 0.132739f
C15070 VDAC_N.t616 VSS 0.105768f
C15071 VDAC_N.n617 VSS 0.132739f
C15072 VDAC_N.t1550 VSS 0.105768f
C15073 VDAC_N.n618 VSS 0.132739f
C15074 VDAC_N.t1361 VSS 0.105768f
C15075 VDAC_N.n619 VSS 0.132739f
C15076 VDAC_N.t1314 VSS 0.105768f
C15077 VDAC_N.n620 VSS 0.12675f
C15078 VDAC_N.t1207 VSS 0.105768f
C15079 VDAC_N.n621 VSS 0.132739f
C15080 VDAC_N.t1771 VSS 0.105768f
C15081 VDAC_N.n622 VSS 0.132739f
C15082 VDAC_N.t559 VSS 0.105768f
C15083 VDAC_N.n623 VSS 0.132739f
C15084 VDAC_N.t1561 VSS 0.105768f
C15085 VDAC_N.n624 VSS 0.132739f
C15086 VDAC_N.t2017 VSS 0.105768f
C15087 VDAC_N.n625 VSS 0.132739f
C15088 VDAC_N.t117 VSS 0.105768f
C15089 VDAC_N.n626 VSS 0.132739f
C15090 VDAC_N.t969 VSS 0.105768f
C15091 VDAC_N.n627 VSS 0.132739f
C15092 VDAC_N.t452 VSS 0.105768f
C15093 VDAC_N.n628 VSS 0.132739f
C15094 VDAC_N.t1803 VSS 0.105768f
C15095 VDAC_N.n629 VSS 0.132739f
C15096 VDAC_N.t1612 VSS 0.105768f
C15097 VDAC_N.n630 VSS 0.132739f
C15098 VDAC_N.t419 VSS 0.105768f
C15099 VDAC_N.n631 VSS 0.132739f
C15100 VDAC_N.t732 VSS 0.105768f
C15101 VDAC_N.n632 VSS 0.132739f
C15102 VDAC_N.t944 VSS 0.105768f
C15103 VDAC_N.n633 VSS 0.132739f
C15104 VDAC_N.t85 VSS 0.105768f
C15105 VDAC_N.n634 VSS 0.132739f
C15106 VDAC_N.t308 VSS 0.105768f
C15107 VDAC_N.n635 VSS 0.132739f
C15108 VDAC_N.t1446 VSS 0.105768f
C15109 VDAC_N.n636 VSS 0.132739f
C15110 VDAC_N.t1148 VSS 0.105768f
C15111 VDAC_N.n637 VSS 0.132739f
C15112 VDAC_N.t528 VSS 0.105768f
C15113 VDAC_N.n638 VSS 0.132739f
C15114 VDAC_N.t161 VSS 0.105768f
C15115 VDAC_N.n639 VSS 0.132739f
C15116 VDAC_N.t1592 VSS 0.105768f
C15117 VDAC_N.n640 VSS 0.132739f
C15118 VDAC_N.t1738 VSS 0.105768f
C15119 VDAC_N.n641 VSS 0.132739f
C15120 VDAC_N.t592 VSS 0.105768f
C15121 VDAC_N.n642 VSS 0.132739f
C15122 VDAC_N.t1526 VSS 0.105768f
C15123 VDAC_N.n643 VSS 0.132739f
C15124 VDAC_N.t1235 VSS 0.105768f
C15125 VDAC_N.n644 VSS 0.132739f
C15126 VDAC_N.t1082 VSS 0.105768f
C15127 VDAC_N.n645 VSS 0.132739f
C15128 VDAC_N.t577 VSS 0.105768f
C15129 VDAC_N.n646 VSS 0.132739f
C15130 VDAC_N.t1593 VSS 0.105768f
C15131 VDAC_N.n647 VSS 0.132739f
C15132 VDAC_N.t914 VSS 0.105768f
C15133 VDAC_N.n648 VSS 0.132739f
C15134 VDAC_N.t391 VSS 0.105768f
C15135 VDAC_N.n649 VSS 0.132739f
C15136 VDAC_N.t1590 VSS 0.105768f
C15137 VDAC_N.n650 VSS 0.132739f
C15138 VDAC_N.t1265 VSS 0.105768f
C15139 VDAC_N.n651 VSS 0.132739f
C15140 VDAC_N.t1837 VSS 0.105768f
C15141 VDAC_N.n652 VSS 0.132739f
C15142 VDAC_N.t311 VSS 0.105768f
C15143 VDAC_N.n653 VSS 0.132739f
C15144 VDAC_N.t825 VSS 0.105768f
C15145 VDAC_N.n654 VSS 0.132739f
C15146 VDAC_N.t1055 VSS 0.105768f
C15147 VDAC_N.n655 VSS 0.132739f
C15148 VDAC_N.t1513 VSS 0.105768f
C15149 VDAC_N.n656 VSS 0.132739f
C15150 VDAC_N.t1969 VSS 0.105768f
C15151 VDAC_N.n657 VSS 0.132739f
C15152 VDAC_N.t663 VSS 0.105768f
C15153 VDAC_N.n658 VSS 0.132739f
C15154 VDAC_N.t143 VSS 0.105768f
C15155 VDAC_N.n659 VSS 0.132739f
C15156 VDAC_N.t1332 VSS 0.105768f
C15157 VDAC_N.n660 VSS 0.132739f
C15158 VDAC_N.t881 VSS 0.105768f
C15159 VDAC_N.n661 VSS 0.132739f
C15160 VDAC_N.t1092 VSS 0.105768f
C15161 VDAC_N.n662 VSS 0.132739f
C15162 VDAC_N.t1230 VSS 0.105768f
C15163 VDAC_N.n663 VSS 0.132739f
C15164 VDAC_N.t1057 VSS 0.105768f
C15165 VDAC_N.n664 VSS 0.132739f
C15166 VDAC_N.t1560 VSS 0.105768f
C15167 VDAC_N.n665 VSS 0.132739f
C15168 VDAC_N.t990 VSS 0.105768f
C15169 VDAC_N.n666 VSS 0.132739f
C15170 VDAC_N.t576 VSS 0.105768f
C15171 VDAC_N.n667 VSS 0.132739f
C15172 VDAC_N.t398 VSS 0.105768f
C15173 VDAC_N.n668 VSS 0.132739f
C15174 VDAC_N.t1364 VSS 0.105768f
C15175 VDAC_N.n669 VSS 0.132739f
C15176 VDAC_N.t342 VSS 0.105768f
C15177 VDAC_N.n670 VSS 0.132739f
C15178 VDAC_N.t301 VSS 0.105768f
C15179 VDAC_N.n671 VSS 0.132739f
C15180 VDAC_N.t1064 VSS 0.105768f
C15181 VDAC_N.n672 VSS 0.132739f
C15182 VDAC_N.t1018 VSS 0.105768f
C15183 VDAC_N.n673 VSS 0.132739f
C15184 VDAC_N.t1473 VSS 0.105768f
C15185 VDAC_N.n674 VSS 0.132739f
C15186 VDAC_N.t1578 VSS 0.105768f
C15187 VDAC_N.n675 VSS 0.132739f
C15188 VDAC_N.t365 VSS 0.105768f
C15189 VDAC_N.n676 VSS 0.132739f
C15190 VDAC_N.t682 VSS 0.105768f
C15191 VDAC_N.n677 VSS 0.132739f
C15192 VDAC_N.t1155 VSS 0.105768f
C15193 VDAC_N.n678 VSS 0.132739f
C15194 VDAC_N.t451 VSS 0.105768f
C15195 VDAC_N.n679 VSS 0.132739f
C15196 VDAC_N.t2058 VSS 0.105768f
C15197 VDAC_N.n680 VSS 0.132739f
C15198 VDAC_N.t1509 VSS 0.105768f
C15199 VDAC_N.n681 VSS 0.132739f
C15200 VDAC_N.t2073 VSS 0.105768f
C15201 VDAC_N.n682 VSS 0.132739f
C15202 VDAC_N.t1403 VSS 0.105768f
C15203 VDAC_N.n683 VSS 0.12675f
C15204 VDAC_N.t128 VSS 0.105768f
C15205 VDAC_N.n684 VSS 0.132739f
C15206 VDAC_N.t1002 VSS 0.105768f
C15207 VDAC_N.n685 VSS 0.132739f
C15208 VDAC_N.t608 VSS 0.105768f
C15209 VDAC_N.n686 VSS 0.132739f
C15210 VDAC_N.t1538 VSS 0.105768f
C15211 VDAC_N.n687 VSS 0.132739f
C15212 VDAC_N.t47 VSS 0.105768f
C15213 VDAC_N.n688 VSS 0.132739f
C15214 VDAC_N.t1306 VSS 0.105768f
C15215 VDAC_N.n689 VSS 0.132739f
C15216 VDAC_N.t97 VSS 0.105768f
C15217 VDAC_N.n690 VSS 0.132739f
C15218 VDAC_N.t1599 VSS 0.105768f
C15219 VDAC_N.n691 VSS 0.132739f
C15220 VDAC_N.t2030 VSS 0.105768f
C15221 VDAC_N.n692 VSS 0.132739f
C15222 VDAC_N.t759 VSS 0.105768f
C15223 VDAC_N.n693 VSS 0.132739f
C15224 VDAC_N.t422 VSS 0.105768f
C15225 VDAC_N.n694 VSS 0.132739f
C15226 VDAC_N.t1385 VSS 0.105768f
C15227 VDAC_N.n695 VSS 0.132739f
C15228 VDAC_N.t483 VSS 0.105768f
C15229 VDAC_N.n696 VSS 0.132739f
C15230 VDAC_N.t79 VSS 0.105768f
C15231 VDAC_N.n697 VSS 0.132739f
C15232 VDAC_N.t289 VSS 0.105768f
C15233 VDAC_N.n698 VSS 0.132739f
C15234 VDAC_N.t2104 VSS 0.105768f
C15235 VDAC_N.n699 VSS 0.132739f
C15236 VDAC_N.t2003 VSS 0.105768f
C15237 VDAC_N.n700 VSS 0.132739f
C15238 VDAC_N.t648 VSS 0.105768f
C15239 VDAC_N.n701 VSS 0.132739f
C15240 VDAC_N.t906 VSS 0.105768f
C15241 VDAC_N.n702 VSS 0.132739f
C15242 VDAC_N.t1604 VSS 0.105768f
C15243 VDAC_N.n703 VSS 0.132739f
C15244 VDAC_N.t1342 VSS 0.105768f
C15245 VDAC_N.n704 VSS 0.132739f
C15246 VDAC_N.t716 VSS 0.105768f
C15247 VDAC_N.n705 VSS 0.132739f
C15248 VDAC_N.t166 VSS 0.105768f
C15249 VDAC_N.n706 VSS 0.132739f
C15250 VDAC_N.t282 VSS 0.105768f
C15251 VDAC_N.n707 VSS 0.132739f
C15252 VDAC_N.t1360 VSS 0.105768f
C15253 VDAC_N.n708 VSS 0.132739f
C15254 VDAC_N.t1842 VSS 0.105768f
C15255 VDAC_N.n709 VSS 0.132739f
C15256 VDAC_N.t71 VSS 0.105768f
C15257 VDAC_N.n710 VSS 0.132739f
C15258 VDAC_N.t114 VSS 0.105768f
C15259 VDAC_N.n711 VSS 0.132739f
C15260 VDAC_N.t659 VSS 0.105768f
C15261 VDAC_N.n712 VSS 0.132739f
C15262 VDAC_N.t610 VSS 0.105768f
C15263 VDAC_N.n713 VSS 0.132739f
C15264 VDAC_N.t10 VSS 0.105768f
C15265 VDAC_N.n714 VSS 0.132739f
C15266 VDAC_N.t433 VSS 0.105768f
C15267 VDAC_N.n715 VSS 0.132739f
C15268 VDAC_N.t1918 VSS 0.105768f
C15269 VDAC_N.n716 VSS 0.132739f
C15270 VDAC_N.t729 VSS 0.105768f
C15271 VDAC_N.n717 VSS 0.132739f
C15272 VDAC_N.t1893 VSS 0.105768f
C15273 VDAC_N.n718 VSS 0.132739f
C15274 VDAC_N.t677 VSS 0.105768f
C15275 VDAC_N.n719 VSS 0.132739f
C15276 VDAC_N.t1783 VSS 0.105768f
C15277 VDAC_N.n720 VSS 0.132739f
C15278 VDAC_N.t95 VSS 0.105768f
C15279 VDAC_N.n721 VSS 0.132739f
C15280 VDAC_N.t1677 VSS 0.105768f
C15281 VDAC_N.n722 VSS 0.132739f
C15282 VDAC_N.t2106 VSS 0.105768f
C15283 VDAC_N.n723 VSS 0.132739f
C15284 VDAC_N.t1543 VSS 0.105768f
C15285 VDAC_N.n724 VSS 0.132739f
C15286 VDAC_N.t1069 VSS 0.105768f
C15287 VDAC_N.n725 VSS 0.132739f
C15288 VDAC_N.t1680 VSS 0.105768f
C15289 VDAC_N.n726 VSS 0.132739f
C15290 VDAC_N.t495 VSS 0.105768f
C15291 VDAC_N.n727 VSS 0.132739f
C15292 VDAC_N.t52 VSS 0.105768f
C15293 VDAC_N.n728 VSS 0.132739f
C15294 VDAC_N.t34 VSS 0.105768f
C15295 VDAC_N.n729 VSS 0.132739f
C15296 VDAC_N.t684 VSS 0.105768f
C15297 VDAC_N.n730 VSS 0.132739f
C15298 VDAC_N.t302 VSS 0.105768f
C15299 VDAC_N.n731 VSS 0.132739f
C15300 VDAC_N.t693 VSS 0.105768f
C15301 VDAC_N.n732 VSS 0.132739f
C15302 VDAC_N.t912 VSS 0.105768f
C15303 VDAC_N.n733 VSS 0.132739f
C15304 VDAC_N.t1834 VSS 0.105768f
C15305 VDAC_N.n734 VSS 0.132739f
C15306 VDAC_N.t1336 VSS 0.105768f
C15307 VDAC_N.n735 VSS 0.132739f
C15308 VDAC_N.t1622 VSS 0.105768f
C15309 VDAC_N.n736 VSS 0.132739f
C15310 VDAC_N.t185 VSS 0.105768f
C15311 VDAC_N.n737 VSS 0.132739f
C15312 VDAC_N.t1178 VSS 0.105768f
C15313 VDAC_N.n738 VSS 0.132739f
C15314 VDAC_N.t1177 VSS 0.105768f
C15315 VDAC_N.n739 VSS 0.132739f
C15316 VDAC_N.t1896 VSS 0.105768f
C15317 VDAC_N.n740 VSS 0.132739f
C15318 VDAC_N.t1902 VSS 0.105768f
C15319 VDAC_N.n741 VSS 0.132739f
C15320 VDAC_N.t75 VSS 0.105768f
C15321 VDAC_N.n742 VSS 0.132739f
C15322 VDAC_N.t850 VSS 0.105768f
C15323 VDAC_N.n743 VSS 0.132739f
C15324 VDAC_N.t1321 VSS 0.105768f
C15325 VDAC_N.n744 VSS 0.132739f
C15326 VDAC_N.t957 VSS 0.105768f
C15327 VDAC_N.n745 VSS 0.132739f
C15328 VDAC_N.t1209 VSS 0.105768f
C15329 VDAC_N.n746 VSS 0.12675f
C15330 VDAC_N.t1216 VSS 0.105768f
C15331 VDAC_N.n747 VSS 0.132739f
C15332 VDAC_N.t1750 VSS 0.105768f
C15333 VDAC_N.n748 VSS 0.132739f
C15334 VDAC_N.t756 VSS 0.105768f
C15335 VDAC_N.n749 VSS 0.132739f
C15336 VDAC_N.t674 VSS 0.105768f
C15337 VDAC_N.n750 VSS 0.132739f
C15338 VDAC_N.t1141 VSS 0.105768f
C15339 VDAC_N.n751 VSS 0.132739f
C15340 VDAC_N.t1106 VSS 0.105768f
C15341 VDAC_N.n752 VSS 0.132739f
C15342 VDAC_N.t2038 VSS 0.105768f
C15343 VDAC_N.n753 VSS 0.132739f
C15344 VDAC_N.t395 VSS 0.105768f
C15345 VDAC_N.n754 VSS 0.132739f
C15346 VDAC_N.t1818 VSS 0.105768f
C15347 VDAC_N.n755 VSS 0.132739f
C15348 VDAC_N.t709 VSS 0.105768f
C15349 VDAC_N.n756 VSS 0.132739f
C15350 VDAC_N.t1374 VSS 0.105768f
C15351 VDAC_N.n757 VSS 0.132739f
C15352 VDAC_N.t1275 VSS 0.105768f
C15353 VDAC_N.n758 VSS 0.132739f
C15354 VDAC_N.t1741 VSS 0.105768f
C15355 VDAC_N.n759 VSS 0.132739f
C15356 VDAC_N.t1515 VSS 0.105768f
C15357 VDAC_N.n760 VSS 0.132739f
C15358 VDAC_N.t1971 VSS 0.105768f
C15359 VDAC_N.n761 VSS 0.132739f
C15360 VDAC_N.t784 VSS 0.105768f
C15361 VDAC_N.n762 VSS 0.132739f
C15362 VDAC_N.t949 VSS 0.105768f
C15363 VDAC_N.n763 VSS 0.132739f
C15364 VDAC_N.t356 VSS 0.105768f
C15365 VDAC_N.n764 VSS 0.132739f
C15366 VDAC_N.t762 VSS 0.105768f
C15367 VDAC_N.n765 VSS 0.132739f
C15368 VDAC_N.t508 VSS 0.105768f
C15369 VDAC_N.n766 VSS 0.132739f
C15370 VDAC_N.t544 VSS 0.105768f
C15371 VDAC_N.n767 VSS 0.132739f
C15372 VDAC_N.t2111 VSS 0.105768f
C15373 VDAC_N.n768 VSS 0.132739f
C15374 VDAC_N.t856 VSS 0.105768f
C15375 VDAC_N.n769 VSS 0.132739f
C15376 VDAC_N.t246 VSS 0.105768f
C15377 VDAC_N.n770 VSS 0.132739f
C15378 VDAC_N.t1572 VSS 0.105768f
C15379 VDAC_N.n771 VSS 0.132739f
C15380 VDAC_N.t1566 VSS 0.105768f
C15381 VDAC_N.n772 VSS 0.132739f
C15382 VDAC_N.t1257 VSS 0.105768f
C15383 VDAC_N.n773 VSS 0.132739f
C15384 VDAC_N.t578 VSS 0.105768f
C15385 VDAC_N.n774 VSS 0.132739f
C15386 VDAC_N.t63 VSS 0.105768f
C15387 VDAC_N.n775 VSS 0.132739f
C15388 VDAC_N.t1800 VSS 0.105768f
C15389 VDAC_N.n776 VSS 0.132739f
C15390 VDAC_N.t1838 VSS 0.105768f
C15391 VDAC_N.n777 VSS 0.132739f
C15392 VDAC_N.t765 VSS 0.105768f
C15393 VDAC_N.n778 VSS 0.132739f
C15394 VDAC_N.t826 VSS 0.105768f
C15395 VDAC_N.n779 VSS 0.132739f
C15396 VDAC_N.t1285 VSS 0.105768f
C15397 VDAC_N.n780 VSS 0.132739f
C15398 VDAC_N.t1749 VSS 0.105768f
C15399 VDAC_N.n781 VSS 0.132739f
C15400 VDAC_N.t603 VSS 0.105768f
C15401 VDAC_N.n782 VSS 0.132739f
C15402 VDAC_N.t129 VSS 0.105768f
C15403 VDAC_N.n783 VSS 0.132739f
C15404 VDAC_N.t1906 VSS 0.105768f
C15405 VDAC_N.n784 VSS 0.132739f
C15406 VDAC_N.t1533 VSS 0.105768f
C15407 VDAC_N.n785 VSS 0.132739f
C15408 VDAC_N.t273 VSS 0.105768f
C15409 VDAC_N.n786 VSS 0.132739f
C15410 VDAC_N.t717 VSS 0.105768f
C15411 VDAC_N.n787 VSS 0.132739f
C15412 VDAC_N.t511 VSS 0.105768f
C15413 VDAC_N.n788 VSS 0.132739f
C15414 VDAC_N.t1096 VSS 0.105768f
C15415 VDAC_N.n789 VSS 0.132739f
C15416 VDAC_N.t55 VSS 0.105768f
C15417 VDAC_N.n790 VSS 0.132739f
C15418 VDAC_N.t1852 VSS 0.105768f
C15419 VDAC_N.n791 VSS 0.132739f
C15420 VDAC_N.t1266 VSS 0.105768f
C15421 VDAC_N.n792 VSS 0.132739f
C15422 VDAC_N.t547 VSS 0.105768f
C15423 VDAC_N.n793 VSS 0.132739f
C15424 VDAC_N.t1672 VSS 0.105768f
C15425 VDAC_N.n794 VSS 0.132739f
C15426 VDAC_N.t1995 VSS 0.105768f
C15427 VDAC_N.n795 VSS 0.132739f
C15428 VDAC_N.t328 VSS 0.105768f
C15429 VDAC_N.n796 VSS 0.132739f
C15430 VDAC_N.t794 VSS 0.105768f
C15431 VDAC_N.n797 VSS 0.132739f
C15432 VDAC_N.t772 VSS 0.105768f
C15433 VDAC_N.n798 VSS 0.132739f
C15434 VDAC_N.t190 VSS 0.105768f
C15435 VDAC_N.n799 VSS 0.132739f
C15436 VDAC_N.t1145 VSS 0.105768f
C15437 VDAC_N.n800 VSS 0.132739f
C15438 VDAC_N.t1792 VSS 0.105768f
C15439 VDAC_N.n801 VSS 0.132739f
C15440 VDAC_N.t154 VSS 0.105768f
C15441 VDAC_N.n802 VSS 0.132739f
C15442 VDAC_N.t352 VSS 0.105768f
C15443 VDAC_N.n803 VSS 0.132739f
C15444 VDAC_N.t1618 VSS 0.105768f
C15445 VDAC_N.n804 VSS 0.132739f
C15446 VDAC_N.t711 VSS 0.105768f
C15447 VDAC_N.n805 VSS 0.132739f
C15448 VDAC_N.t1382 VSS 0.105768f
C15449 VDAC_N.n806 VSS 0.132739f
C15450 VDAC_N.t171 VSS 0.105768f
C15451 VDAC_N.n807 VSS 0.132739f
C15452 VDAC_N.t887 VSS 0.105768f
C15453 VDAC_N.n808 VSS 0.132739f
C15454 VDAC_N.t2098 VSS 0.105768f
C15455 VDAC_N.n809 VSS 0.12675f
C15456 VDAC_N.t1689 VSS 0.105768f
C15457 VDAC_N.n810 VSS 0.132739f
C15458 VDAC_N.t1388 VSS 0.105768f
C15459 VDAC_N.n811 VSS 0.132739f
C15460 VDAC_N.t801 VSS 0.105768f
C15461 VDAC_N.n812 VSS 0.132739f
C15462 VDAC_N.t1033 VSS 0.105768f
C15463 VDAC_N.n813 VSS 0.132739f
C15464 VDAC_N.t1352 VSS 0.105768f
C15465 VDAC_N.n814 VSS 0.132739f
C15466 VDAC_N.t1925 VSS 0.105768f
C15467 VDAC_N.n815 VSS 0.132739f
C15468 VDAC_N.t1844 VSS 0.105768f
C15469 VDAC_N.n816 VSS 0.132739f
C15470 VDAC_N.t1398 VSS 0.105768f
C15471 VDAC_N.n817 VSS 0.132739f
C15472 VDAC_N.t1868 VSS 0.105768f
C15473 VDAC_N.n818 VSS 0.132739f
C15474 VDAC_N.t318 VSS 0.105768f
C15475 VDAC_N.n819 VSS 0.132739f
C15476 VDAC_N.t537 VSS 0.105768f
C15477 VDAC_N.n820 VSS 0.132739f
C15478 VDAC_N.t264 VSS 0.105768f
C15479 VDAC_N.n821 VSS 0.132739f
C15480 VDAC_N.t1914 VSS 0.105768f
C15481 VDAC_N.n822 VSS 0.132739f
C15482 VDAC_N.t353 VSS 0.105768f
C15483 VDAC_N.n823 VSS 0.132739f
C15484 VDAC_N.t1785 VSS 0.105768f
C15485 VDAC_N.n824 VSS 0.132739f
C15486 VDAC_N.t1524 VSS 0.105768f
C15487 VDAC_N.n825 VSS 0.132739f
C15488 VDAC_N.t441 VSS 0.105768f
C15489 VDAC_N.n826 VSS 0.132739f
C15490 VDAC_N.t93 VSS 0.105768f
C15491 VDAC_N.n827 VSS 0.132739f
C15492 VDAC_N.t570 VSS 0.105768f
C15493 VDAC_N.n828 VSS 0.132739f
C15494 VDAC_N.t153 VSS 0.105768f
C15495 VDAC_N.n829 VSS 0.132739f
C15496 VDAC_N.t1328 VSS 0.105768f
C15497 VDAC_N.n830 VSS 0.132739f
C15498 VDAC_N.t501 VSS 0.105768f
C15499 VDAC_N.n831 VSS 0.132739f
C15500 VDAC_N.t468 VSS 0.105768f
C15501 VDAC_N.n832 VSS 0.132739f
C15502 VDAC_N.t706 VSS 0.105768f
C15503 VDAC_N.n833 VSS 0.132739f
C15504 VDAC_N.t1180 VSS 0.105768f
C15505 VDAC_N.n834 VSS 0.132739f
C15506 VDAC_N.t598 VSS 0.105768f
C15507 VDAC_N.n835 VSS 0.132739f
C15508 VDAC_N.t546 VSS 0.105768f
C15509 VDAC_N.n836 VSS 0.132739f
C15510 VDAC_N.t384 VSS 0.105768f
C15511 VDAC_N.n837 VSS 0.132739f
C15512 VDAC_N.t958 VSS 0.105768f
C15513 VDAC_N.n838 VSS 0.132739f
C15514 VDAC_N.t2020 VSS 0.105768f
C15515 VDAC_N.n839 VSS 0.132739f
C15516 VDAC_N.t1442 VSS 0.105768f
C15517 VDAC_N.n840 VSS 0.132739f
C15518 VDAC_N.t671 VSS 0.105768f
C15519 VDAC_N.n841 VSS 0.132739f
C15520 VDAC_N.t630 VSS 0.105768f
C15521 VDAC_N.n842 VSS 0.132739f
C15522 VDAC_N.t1087 VSS 0.105768f
C15523 VDAC_N.n843 VSS 0.132739f
C15524 VDAC_N.t1555 VSS 0.105768f
C15525 VDAC_N.n844 VSS 0.132739f
C15526 VDAC_N.t1954 VSS 0.105768f
C15527 VDAC_N.n845 VSS 0.132739f
C15528 VDAC_N.t1451 VSS 0.105768f
C15529 VDAC_N.n846 VSS 0.132739f
C15530 VDAC_N.t214 VSS 0.105768f
C15531 VDAC_N.n847 VSS 0.132739f
C15532 VDAC_N.t1345 VSS 0.105768f
C15533 VDAC_N.n848 VSS 0.132739f
C15534 VDAC_N.t471 VSS 0.105768f
C15535 VDAC_N.n849 VSS 0.132739f
C15536 VDAC_N.t1213 VSS 0.105768f
C15537 VDAC_N.n850 VSS 0.132739f
C15538 VDAC_N.t465 VSS 0.105768f
C15539 VDAC_N.n851 VSS 0.132739f
C15540 VDAC_N.t332 VSS 0.105768f
C15541 VDAC_N.n852 VSS 0.132739f
C15542 VDAC_N.t1563 VSS 0.105768f
C15543 VDAC_N.n853 VSS 0.132739f
C15544 VDAC_N.t2025 VSS 0.105768f
C15545 VDAC_N.n854 VSS 0.132739f
C15546 VDAC_N.t136 VSS 0.105768f
C15547 VDAC_N.n855 VSS 0.132739f
C15548 VDAC_N.t971 VSS 0.105768f
C15549 VDAC_N.n856 VSS 0.132739f
C15550 VDAC_N.t1764 VSS 0.105768f
C15551 VDAC_N.n857 VSS 0.132739f
C15552 VDAC_N.t1807 VSS 0.105768f
C15553 VDAC_N.n858 VSS 0.132739f
C15554 VDAC_N.t1676 VSS 0.105768f
C15555 VDAC_N.n859 VSS 0.132739f
C15556 VDAC_N.t1162 VSS 0.105768f
C15557 VDAC_N.n860 VSS 0.132739f
C15558 VDAC_N.t1116 VSS 0.105768f
C15559 VDAC_N.n861 VSS 0.132739f
C15560 VDAC_N.t952 VSS 0.105768f
C15561 VDAC_N.n862 VSS 0.132739f
C15562 VDAC_N.t954 VSS 0.105768f
C15563 VDAC_N.n863 VSS 0.132739f
C15564 VDAC_N.t276 VSS 0.105768f
C15565 VDAC_N.n864 VSS 0.132739f
C15566 VDAC_N.t1654 VSS 0.105768f
C15567 VDAC_N.n865 VSS 0.132739f
C15568 VDAC_N.t44 VSS 0.105768f
C15569 VDAC_N.n866 VSS 0.132739f
C15570 VDAC_N.t1226 VSS 0.105768f
C15571 VDAC_N.n867 VSS 0.132739f
C15572 VDAC_N.t613 VSS 0.105768f
C15573 VDAC_N.n868 VSS 0.132739f
C15574 VDAC_N.t1992 VSS 0.105768f
C15575 VDAC_N.n869 VSS 0.132739f
C15576 VDAC_N.t1950 VSS 0.105768f
C15577 VDAC_N.n870 VSS 0.132739f
C15578 VDAC_N.t409 VSS 0.105768f
C15579 VDAC_N.n871 VSS 0.132739f
C15580 VDAC_N.t1718 VSS 0.105768f
C15581 VDAC_N.n872 VSS 0.12675f
C15582 VDAC_N.t1782 VSS 0.105768f
C15583 VDAC_N.n873 VSS 0.132739f
C15584 VDAC_N.t389 VSS 0.105768f
C15585 VDAC_N.n874 VSS 0.132739f
C15586 VDAC_N.t414 VSS 0.105768f
C15587 VDAC_N.n875 VSS 0.132739f
C15588 VDAC_N.t105 VSS 0.105768f
C15589 VDAC_N.n876 VSS 0.132739f
C15590 VDAC_N.t1721 VSS 0.105768f
C15591 VDAC_N.n877 VSS 0.132739f
C15592 VDAC_N.t1153 VSS 0.105768f
C15593 VDAC_N.n878 VSS 0.132739f
C15594 VDAC_N.t1613 VSS 0.105768f
C15595 VDAC_N.n879 VSS 0.132739f
C15596 VDAC_N.t539 VSS 0.105768f
C15597 VDAC_N.n880 VSS 0.132739f
C15598 VDAC_N.t767 VSS 0.105768f
C15599 VDAC_N.n881 VSS 0.132739f
C15600 VDAC_N.t993 VSS 0.105768f
C15601 VDAC_N.n882 VSS 0.132739f
C15602 VDAC_N.t1289 VSS 0.105768f
C15603 VDAC_N.n883 VSS 0.132739f
C15604 VDAC_N.t257 VSS 0.105768f
C15605 VDAC_N.n884 VSS 0.132739f
C15606 VDAC_N.t1268 VSS 0.105768f
C15607 VDAC_N.n885 VSS 0.132739f
C15608 VDAC_N.t1129 VSS 0.105768f
C15609 VDAC_N.n886 VSS 0.132739f
C15610 VDAC_N.t1595 VSS 0.105768f
C15611 VDAC_N.n887 VSS 0.132739f
C15612 VDAC_N.t156 VSS 0.105768f
C15613 VDAC_N.n888 VSS 0.132739f
C15614 VDAC_N.t1483 VSS 0.105768f
C15615 VDAC_N.n889 VSS 0.132739f
C15616 VDAC_N.t1939 VSS 0.105768f
C15617 VDAC_N.n890 VSS 0.132739f
C15618 VDAC_N.t376 VSS 0.105768f
C15619 VDAC_N.n891 VSS 0.132739f
C15620 VDAC_N.t481 VSS 0.105768f
C15621 VDAC_N.n892 VSS 0.132739f
C15622 VDAC_N.t2092 VSS 0.105768f
C15623 VDAC_N.n893 VSS 0.132739f
C15624 VDAC_N.t1731 VSS 0.105768f
C15625 VDAC_N.n894 VSS 0.132739f
C15626 VDAC_N.t28 VSS 0.105768f
C15627 VDAC_N.n895 VSS 0.132739f
C15628 VDAC_N.t520 VSS 0.105768f
C15629 VDAC_N.n896 VSS 0.132739f
C15630 VDAC_N.t271 VSS 0.105768f
C15631 VDAC_N.n897 VSS 0.132739f
C15632 VDAC_N.t1544 VSS 0.105768f
C15633 VDAC_N.n898 VSS 0.132739f
C15634 VDAC_N.t874 VSS 0.105768f
C15635 VDAC_N.n899 VSS 0.132739f
C15636 VDAC_N.t1348 VSS 0.105768f
C15637 VDAC_N.n900 VSS 0.132739f
C15638 VDAC_N.t1498 VSS 0.105768f
C15639 VDAC_N.n901 VSS 0.132739f
C15640 VDAC_N.t1980 VSS 0.105768f
C15641 VDAC_N.n902 VSS 0.132739f
C15642 VDAC_N.t2096 VSS 0.105768f
C15643 VDAC_N.n903 VSS 0.132739f
C15644 VDAC_N.t45 VSS 0.105768f
C15645 VDAC_N.n904 VSS 0.132739f
C15646 VDAC_N.t1688 VSS 0.105768f
C15647 VDAC_N.n905 VSS 0.132739f
C15648 VDAC_N.t1774 VSS 0.105768f
C15649 VDAC_N.n906 VSS 0.132739f
C15650 VDAC_N.t49 VSS 0.105768f
C15651 VDAC_N.n907 VSS 0.132739f
C15652 VDAC_N.t798 VSS 0.105768f
C15653 VDAC_N.n908 VSS 0.132739f
C15654 VDAC_N.t643 VSS 0.105768f
C15655 VDAC_N.n909 VSS 0.132739f
C15656 VDAC_N.t1130 VSS 0.105768f
C15657 VDAC_N.n910 VSS 0.132739f
C15658 VDAC_N.t1149 VSS 0.105768f
C15659 VDAC_N.n911 VSS 0.132739f
C15660 VDAC_N.t819 VSS 0.105768f
C15661 VDAC_N.n912 VSS 0.132739f
C15662 VDAC_N.t2014 VSS 0.105768f
C15663 VDAC_N.n913 VSS 0.132739f
C15664 VDAC_N.t223 VSS 0.105768f
C15665 VDAC_N.n914 VSS 0.132739f
C15666 VDAC_N.t2045 VSS 0.105768f
C15667 VDAC_N.n915 VSS 0.132739f
C15668 VDAC_N.t1377 VSS 0.105768f
C15669 VDAC_N.n916 VSS 0.132739f
C15670 VDAC_N.t141 VSS 0.105768f
C15671 VDAC_N.n917 VSS 0.132739f
C15672 VDAC_N.t500 VSS 0.105768f
C15673 VDAC_N.n918 VSS 0.132739f
C15674 VDAC_N.t81 VSS 0.105768f
C15675 VDAC_N.n919 VSS 0.132739f
C15676 VDAC_N.t988 VSS 0.105768f
C15677 VDAC_N.n920 VSS 0.132739f
C15678 VDAC_N.t425 VSS 0.105768f
C15679 VDAC_N.n921 VSS 0.132739f
C15680 VDAC_N.t2077 VSS 0.105768f
C15681 VDAC_N.n922 VSS 0.132739f
C15682 VDAC_N.t776 VSS 0.105768f
C15683 VDAC_N.n923 VSS 0.132739f
C15684 VDAC_N.t995 VSS 0.105768f
C15685 VDAC_N.n924 VSS 0.132739f
C15686 VDAC_N.t296 VSS 0.105768f
C15687 VDAC_N.n925 VSS 0.132739f
C15688 VDAC_N.t758 VSS 0.105768f
C15689 VDAC_N.n926 VSS 0.132739f
C15690 VDAC_N.t956 VSS 0.105768f
C15691 VDAC_N.n927 VSS 0.132739f
C15692 VDAC_N.t1270 VSS 0.105768f
C15693 VDAC_N.n928 VSS 0.132739f
C15694 VDAC_N.t2105 VSS 0.105768f
C15695 VDAC_N.n929 VSS 0.132739f
C15696 VDAC_N.t440 VSS 0.105768f
C15697 VDAC_N.n930 VSS 0.132739f
C15698 VDAC_N.t1998 VSS 0.105768f
C15699 VDAC_N.n931 VSS 0.132739f
C15700 VDAC_N.t1232 VSS 0.105768f
C15701 VDAC_N.n932 VSS 0.132739f
C15702 VDAC_N.t1562 VSS 0.105768f
C15703 VDAC_N.n933 VSS 0.132739f
C15704 VDAC_N.t1367 VSS 0.105768f
C15705 VDAC_N.n934 VSS 0.132739f
C15706 VDAC_N.t1326 VSS 0.105768f
C15707 VDAC_N.n935 VSS 0.12675f
C15708 VDAC_N.t2019 VSS 0.105768f
C15709 VDAC_N.n936 VSS 0.132739f
C15710 VDAC_N.t456 VSS 0.105768f
C15711 VDAC_N.n937 VSS 0.132739f
C15712 VDAC_N.t499 VSS 0.105768f
C15713 VDAC_N.n938 VSS 0.132739f
C15714 VDAC_N.t884 VSS 0.105768f
C15715 VDAC_N.n939 VSS 0.132739f
C15716 VDAC_N.t1362 VSS 0.105768f
C15717 VDAC_N.n940 VSS 0.132739f
C15718 VDAC_N.t1644 VSS 0.105768f
C15719 VDAC_N.n941 VSS 0.132739f
C15720 VDAC_N.t310 VSS 0.105768f
C15721 VDAC_N.n942 VSS 0.132739f
C15722 VDAC_N.t2086 VSS 0.105768f
C15723 VDAC_N.n943 VSS 0.132739f
C15724 VDAC_N.t488 VSS 0.105768f
C15725 VDAC_N.n944 VSS 0.132739f
C15726 VDAC_N.t950 VSS 0.105768f
C15727 VDAC_N.n945 VSS 0.132739f
C15728 VDAC_N.t516 VSS 0.105768f
C15729 VDAC_N.n946 VSS 0.132739f
C15730 VDAC_N.t838 VSS 0.105768f
C15731 VDAC_N.n947 VSS 0.132739f
C15732 VDAC_N.t33 VSS 0.105768f
C15733 VDAC_N.n948 VSS 0.132739f
C15734 VDAC_N.t1855 VSS 0.105768f
C15735 VDAC_N.n949 VSS 0.132739f
C15736 VDAC_N.t1204 VSS 0.105768f
C15737 VDAC_N.n950 VSS 0.132739f
C15738 VDAC_N.t386 VSS 0.105768f
C15739 VDAC_N.n951 VSS 0.132739f
C15740 VDAC_N.t188 VSS 0.105768f
C15741 VDAC_N.n952 VSS 0.132739f
C15742 VDAC_N.t280 VSS 0.105768f
C15743 VDAC_N.n953 VSS 0.132739f
C15744 VDAC_N.t1099 VSS 0.105768f
C15745 VDAC_N.n954 VSS 0.132739f
C15746 VDAC_N.t1616 VSS 0.105768f
C15747 VDAC_N.n955 VSS 0.132739f
C15748 VDAC_N.t1742 VSS 0.105768f
C15749 VDAC_N.n956 VSS 0.132739f
C15750 VDAC_N.t1184 VSS 0.105768f
C15751 VDAC_N.n957 VSS 0.132739f
C15752 VDAC_N.t1534 VSS 0.105768f
C15753 VDAC_N.n958 VSS 0.132739f
C15754 VDAC_N.t331 VSS 0.105768f
C15755 VDAC_N.n959 VSS 0.132739f
C15756 VDAC_N.t294 VSS 0.105768f
C15757 VDAC_N.n960 VSS 0.132739f
C15758 VDAC_N.t579 VSS 0.105768f
C15759 VDAC_N.n961 VSS 0.132739f
C15760 VDAC_N.t1597 VSS 0.105768f
C15761 VDAC_N.n962 VSS 0.132739f
C15762 VDAC_N.t474 VSS 0.105768f
C15763 VDAC_N.n963 VSS 0.132739f
C15764 VDAC_N.t757 VSS 0.105768f
C15765 VDAC_N.n964 VSS 0.132739f
C15766 VDAC_N.t126 VSS 0.105768f
C15767 VDAC_N.n965 VSS 0.132739f
C15768 VDAC_N.t1271 VSS 0.105768f
C15769 VDAC_N.n966 VSS 0.132739f
C15770 VDAC_N.t255 VSS 0.105768f
C15771 VDAC_N.n967 VSS 0.132739f
C15772 VDAC_N.t1163 VSS 0.105768f
C15773 VDAC_N.n968 VSS 0.132739f
C15774 VDAC_N.t1625 VSS 0.105768f
C15775 VDAC_N.n969 VSS 0.132739f
C15776 VDAC_N.t2085 VSS 0.105768f
C15777 VDAC_N.n970 VSS 0.132739f
C15778 VDAC_N.t121 VSS 0.105768f
C15779 VDAC_N.n971 VSS 0.132739f
C15780 VDAC_N.t1001 VSS 0.105768f
C15781 VDAC_N.n972 VSS 0.132739f
C15782 VDAC_N.t347 VSS 0.105768f
C15783 VDAC_N.n973 VSS 0.132739f
C15784 VDAC_N.t1871 VSS 0.105768f
C15785 VDAC_N.n974 VSS 0.132739f
C15786 VDAC_N.t692 VSS 0.105768f
C15787 VDAC_N.n975 VSS 0.132739f
C15788 VDAC_N.t135 VSS 0.105768f
C15789 VDAC_N.n976 VSS 0.132739f
C15790 VDAC_N.t1140 VSS 0.105768f
C15791 VDAC_N.n977 VSS 0.132739f
C15792 VDAC_N.t1238 VSS 0.105768f
C15793 VDAC_N.n978 VSS 0.132739f
C15794 VDAC_N.t157 VSS 0.105768f
C15795 VDAC_N.n979 VSS 0.132739f
C15796 VDAC_N.t816 VSS 0.105768f
C15797 VDAC_N.n980 VSS 0.132739f
C15798 VDAC_N.t994 VSS 0.105768f
C15799 VDAC_N.n981 VSS 0.132739f
C15800 VDAC_N.t1160 VSS 0.105768f
C15801 VDAC_N.n982 VSS 0.132739f
C15802 VDAC_N.t1530 VSS 0.105768f
C15803 VDAC_N.n983 VSS 0.132739f
C15804 VDAC_N.t1412 VSS 0.105768f
C15805 VDAC_N.n984 VSS 0.132739f
C15806 VDAC_N.t186 VSS 0.105768f
C15807 VDAC_N.n985 VSS 0.132739f
C15808 VDAC_N.t1127 VSS 0.105768f
C15809 VDAC_N.n986 VSS 0.132739f
C15810 VDAC_N.t2128 VSS 0.105768f
C15811 VDAC_N.n987 VSS 0.132739f
C15812 VDAC_N.t2018 VSS 0.105768f
C15813 VDAC_N.n988 VSS 0.132739f
C15814 VDAC_N.t755 VSS 0.105768f
C15815 VDAC_N.n989 VSS 0.132739f
C15816 VDAC_N.t1594 VSS 0.105768f
C15817 VDAC_N.n990 VSS 0.132739f
C15818 VDAC_N.t1379 VSS 0.105768f
C15819 VDAC_N.n991 VSS 0.132739f
C15820 VDAC_N.t686 VSS 0.105768f
C15821 VDAC_N.n992 VSS 0.132739f
C15822 VDAC_N.t1161 VSS 0.105768f
C15823 VDAC_N.n993 VSS 0.132739f
C15824 VDAC_N.t453 VSS 0.105768f
C15825 VDAC_N.n994 VSS 0.132739f
C15826 VDAC_N.t2070 VSS 0.105768f
C15827 VDAC_N.n995 VSS 0.132739f
C15828 VDAC_N.t771 VSS 0.105768f
C15829 VDAC_N.n996 VSS 0.132739f
C15830 VDAC_N.t2081 VSS 0.105768f
C15831 VDAC_N.n997 VSS 0.132739f
C15832 VDAC_N.t373 VSS 0.105768f
C15833 VDAC_N.n998 VSS 0.12675f
C15834 VDAC_N.t637 VSS 0.105768f
C15835 VDAC_N.n999 VSS 0.132739f
C15836 VDAC_N.t921 VSS 0.105768f
C15837 VDAC_N.n1000 VSS 0.132739f
C15838 VDAC_N.t1135 VSS 0.105768f
C15839 VDAC_N.n1001 VSS 0.132739f
C15840 VDAC_N.t1601 VSS 0.105768f
C15841 VDAC_N.n1002 VSS 0.132739f
C15842 VDAC_N.t1043 VSS 0.105768f
C15843 VDAC_N.n1003 VSS 0.132739f
C15844 VDAC_N.t211 VSS 0.105768f
C15845 VDAC_N.n1004 VSS 0.132739f
C15846 VDAC_N.t1943 VSS 0.105768f
C15847 VDAC_N.n1005 VSS 0.132739f
C15848 VDAC_N.t532 VSS 0.105768f
C15849 VDAC_N.n1006 VSS 0.132739f
C15850 VDAC_N.t939 VSS 0.105768f
C15851 VDAC_N.n1007 VSS 0.132739f
C15852 VDAC_N.t580 VSS 0.105768f
C15853 VDAC_N.n1008 VSS 0.132739f
C15854 VDAC_N.t429 VSS 0.105768f
C15855 VDAC_N.n1009 VSS 0.132739f
C15856 VDAC_N.t1084 VSS 0.105768f
C15857 VDAC_N.n1010 VSS 0.132739f
C15858 VDAC_N.t2024 VSS 0.105768f
C15859 VDAC_N.n1011 VSS 0.132739f
C15860 VDAC_N.t1663 VSS 0.105768f
C15861 VDAC_N.n1012 VSS 0.132739f
C15862 VDAC_N.t1075 VSS 0.105768f
C15863 VDAC_N.n1013 VSS 0.132739f
C15864 VDAC_N.t1080 VSS 0.105768f
C15865 VDAC_N.n1014 VSS 0.132739f
C15866 VDAC_N.t523 VSS 0.105768f
C15867 VDAC_N.n1015 VSS 0.132739f
C15868 VDAC_N.t1280 VSS 0.105768f
C15869 VDAC_N.n1016 VSS 0.132739f
C15870 VDAC_N.t1798 VSS 0.105768f
C15871 VDAC_N.n1017 VSS 0.132739f
C15872 VDAC_N.t1652 VSS 0.105768f
C15873 VDAC_N.n1018 VSS 0.132739f
C15874 VDAC_N.t1346 VSS 0.105768f
C15875 VDAC_N.n1019 VSS 0.132739f
C15876 VDAC_N.t1548 VSS 0.105768f
C15877 VDAC_N.n1020 VSS 0.132739f
C15878 VDAC_N.t586 VSS 0.105768f
C15879 VDAC_N.n1021 VSS 0.132739f
C15880 VDAC_N.t1050 VSS 0.105768f
C15881 VDAC_N.n1022 VSS 0.132739f
C15882 VDAC_N.t704 VSS 0.105768f
C15883 VDAC_N.n1023 VSS 0.132739f
C15884 VDAC_N.t1854 VSS 0.105768f
C15885 VDAC_N.n1024 VSS 0.132739f
C15886 VDAC_N.t1409 VSS 0.105768f
C15887 VDAC_N.n1025 VSS 0.132739f
C15888 VDAC_N.t374 VSS 0.105768f
C15889 VDAC_N.n1026 VSS 0.132739f
C15890 VDAC_N.t1297 VSS 0.105768f
C15891 VDAC_N.n1027 VSS 0.132739f
C15892 VDAC_N.t614 VSS 0.105768f
C15893 VDAC_N.n1028 VSS 0.132739f
C15894 VDAC_N.t13 VSS 0.105768f
C15895 VDAC_N.n1029 VSS 0.132739f
C15896 VDAC_N.t841 VSS 0.105768f
C15897 VDAC_N.n1030 VSS 0.132739f
C15898 VDAC_N.t1926 VSS 0.105768f
C15899 VDAC_N.n1031 VSS 0.132739f
C15900 VDAC_N.t1433 VSS 0.105768f
C15901 VDAC_N.n1032 VSS 0.132739f
C15902 VDAC_N.t1895 VSS 0.105768f
C15903 VDAC_N.n1033 VSS 0.132739f
C15904 VDAC_N.t1329 VSS 0.105768f
C15905 VDAC_N.n1034 VSS 0.132739f
C15906 VDAC_N.t1787 VSS 0.105768f
C15907 VDAC_N.n1035 VSS 0.132739f
C15908 VDAC_N.t567 VSS 0.105768f
C15909 VDAC_N.n1036 VSS 0.132739f
C15910 VDAC_N.t855 VSS 0.105768f
C15911 VDAC_N.n1037 VSS 0.132739f
C15912 VDAC_N.t1371 VSS 0.105768f
C15913 VDAC_N.n1038 VSS 0.132739f
C15914 VDAC_N.t1547 VSS 0.105768f
C15915 VDAC_N.n1039 VSS 0.132739f
C15916 VDAC_N.t1071 VSS 0.105768f
C15917 VDAC_N.n1040 VSS 0.132739f
C15918 VDAC_N.t864 VSS 0.105768f
C15919 VDAC_N.n1041 VSS 0.132739f
C15920 VDAC_N.t145 VSS 0.105768f
C15921 VDAC_N.n1042 VSS 0.132739f
C15922 VDAC_N.t228 VSS 0.105768f
C15923 VDAC_N.n1043 VSS 0.132739f
C15924 VDAC_N.t802 VSS 0.105768f
C15925 VDAC_N.n1044 VSS 0.132739f
C15926 VDAC_N.t1452 VSS 0.105768f
C15927 VDAC_N.n1045 VSS 0.132739f
C15928 VDAC_N.t1138 VSS 0.105768f
C15929 VDAC_N.n1046 VSS 0.132739f
C15930 VDAC_N.t9 VSS 0.105768f
C15931 VDAC_N.n1047 VSS 0.132739f
C15932 VDAC_N.t56 VSS 0.105768f
C15933 VDAC_N.n1048 VSS 0.132739f
C15934 VDAC_N.t1846 VSS 0.105768f
C15935 VDAC_N.n1049 VSS 0.132739f
C15936 VDAC_N.t360 VSS 0.105768f
C15937 VDAC_N.n1050 VSS 0.132739f
C15938 VDAC_N.t1630 VSS 0.105768f
C15939 VDAC_N.n1051 VSS 0.132739f
C15940 VDAC_N.t1293 VSS 0.105768f
C15941 VDAC_N.n1052 VSS 0.132739f
C15942 VDAC_N.t1198 VSS 0.105768f
C15943 VDAC_N.n1053 VSS 0.132739f
C15944 VDAC_N.t605 VSS 0.105768f
C15945 VDAC_N.n1054 VSS 0.132739f
C15946 VDAC_N.t1920 VSS 0.105768f
C15947 VDAC_N.n1055 VSS 0.132739f
C15948 VDAC_N.t1922 VSS 0.105768f
C15949 VDAC_N.n1056 VSS 0.132739f
C15950 VDAC_N.t1539 VSS 0.105768f
C15951 VDAC_N.n1057 VSS 0.132739f
C15952 VDAC_N.t1686 VSS 0.105768f
C15953 VDAC_N.n1058 VSS 0.132739f
C15954 VDAC_N.t1327 VSS 0.105768f
C15955 VDAC_N.n1059 VSS 0.132739f
C15956 VDAC_N.t261 VSS 0.105768f
C15957 VDAC_N.n1060 VSS 0.132739f
C15958 VDAC_N.t1215 VSS 0.105768f
C15959 VDAC_N.n1061 VSS 0.12675f
C15960 VDAC_N.t820 VSS 0.105768f
C15961 VDAC_N.n1062 VSS 0.132739f
C15962 VDAC_N.t1574 VSS 0.105768f
C15963 VDAC_N.n1063 VSS 0.132739f
C15964 VDAC_N.t204 VSS 0.105768f
C15965 VDAC_N.n1064 VSS 0.132739f
C15966 VDAC_N.t582 VSS 0.105768f
C15967 VDAC_N.n1065 VSS 0.132739f
C15968 VDAC_N.t1046 VSS 0.105768f
C15969 VDAC_N.n1066 VSS 0.132739f
C15970 VDAC_N.t1816 VSS 0.105768f
C15971 VDAC_N.n1067 VSS 0.132739f
C15972 VDAC_N.t482 VSS 0.105768f
C15973 VDAC_N.n1068 VSS 0.132739f
C15974 VDAC_N.t1405 VSS 0.105768f
C15975 VDAC_N.n1069 VSS 0.132739f
C15976 VDAC_N.t78 VSS 0.105768f
C15977 VDAC_N.n1070 VSS 0.132739f
C15978 VDAC_N.t107 VSS 0.105768f
C15979 VDAC_N.n1071 VSS 0.132739f
C15980 VDAC_N.t174 VSS 0.105768f
C15981 VDAC_N.n1072 VSS 0.132739f
C15982 VDAC_N.t37 VSS 0.105768f
C15983 VDAC_N.n1073 VSS 0.132739f
C15984 VDAC_N.t839 VSS 0.105768f
C15985 VDAC_N.n1074 VSS 0.132739f
C15986 VDAC_N.t1780 VSS 0.105768f
C15987 VDAC_N.n1075 VSS 0.132739f
C15988 VDAC_N.t1378 VSS 0.105768f
C15989 VDAC_N.n1076 VSS 0.132739f
C15990 VDAC_N.t653 VSS 0.105768f
C15991 VDAC_N.n1077 VSS 0.132739f
C15992 VDAC_N.t1166 VSS 0.105768f
C15993 VDAC_N.n1078 VSS 0.132739f
C15994 VDAC_N.t2094 VSS 0.105768f
C15995 VDAC_N.n1079 VSS 0.132739f
C15996 VDAC_N.t229 VSS 0.105768f
C15997 VDAC_N.n1080 VSS 0.132739f
C15998 VDAC_N.t86 VSS 0.105768f
C15999 VDAC_N.n1081 VSS 0.132739f
C16000 VDAC_N.t723 VSS 0.105768f
C16001 VDAC_N.n1082 VSS 0.132739f
C16002 VDAC_N.t1662 VSS 0.105768f
C16003 VDAC_N.n1083 VSS 0.132739f
C16004 VDAC_N.t349 VSS 0.105768f
C16005 VDAC_N.n1084 VSS 0.132739f
C16006 VDAC_N.t1767 VSS 0.105768f
C16007 VDAC_N.n1085 VSS 0.132739f
C16008 VDAC_N.t1085 VSS 0.105768f
C16009 VDAC_N.n1086 VSS 0.132739f
C16010 VDAC_N.t437 VSS 0.105768f
C16011 VDAC_N.n1087 VSS 0.132739f
C16012 VDAC_N.t159 VSS 0.105768f
C16013 VDAC_N.n1088 VSS 0.132739f
C16014 VDAC_N.t1449 VSS 0.105768f
C16015 VDAC_N.n1089 VSS 0.132739f
C16016 VDAC_N.t1019 VSS 0.105768f
C16017 VDAC_N.n1090 VSS 0.132739f
C16018 VDAC_N.t357 VSS 0.105768f
C16019 VDAC_N.n1091 VSS 0.132739f
C16020 VDAC_N.t1799 VSS 0.105768f
C16021 VDAC_N.n1092 VSS 0.132739f
C16022 VDAC_N.t852 VSS 0.105768f
C16023 VDAC_N.n1093 VSS 0.132739f
C16024 VDAC_N.t863 VSS 0.105768f
C16025 VDAC_N.n1094 VSS 0.132739f
C16026 VDAC_N.t860 VSS 0.105768f
C16027 VDAC_N.n1095 VSS 0.132739f
C16028 VDAC_N.t936 VSS 0.105768f
C16029 VDAC_N.n1096 VSS 0.132739f
C16030 VDAC_N.t2043 VSS 0.105768f
C16031 VDAC_N.n1097 VSS 0.132739f
C16032 VDAC_N.t368 VSS 0.105768f
C16033 VDAC_N.n1098 VSS 0.132739f
C16034 VDAC_N.t929 VSS 0.105768f
C16035 VDAC_N.n1099 VSS 0.132739f
C16036 VDAC_N.t1892 VSS 0.105768f
C16037 VDAC_N.n1100 VSS 0.132739f
C16038 VDAC_N.t1414 VSS 0.105768f
C16039 VDAC_N.n1101 VSS 0.132739f
C16040 VDAC_N.t844 VSS 0.105768f
C16041 VDAC_N.n1102 VSS 0.132739f
C16042 VDAC_N.t1358 VSS 0.105768f
C16043 VDAC_N.n1103 VSS 0.132739f
C16044 VDAC_N.t597 VSS 0.105768f
C16045 VDAC_N.n1104 VSS 0.132739f
C16046 VDAC_N.t1872 VSS 0.105768f
C16047 VDAC_N.n1105 VSS 0.132739f
C16048 VDAC_N.t490 VSS 0.105768f
C16049 VDAC_N.n1106 VSS 0.132739f
C16050 VDAC_N.t401 VSS 0.105768f
C16051 VDAC_N.n1107 VSS 0.132739f
C16052 VDAC_N.t1650 VSS 0.105768f
C16053 VDAC_N.n1108 VSS 0.132739f
C16054 VDAC_N.t669 VSS 0.105768f
C16055 VDAC_N.n1109 VSS 0.132739f
C16056 VDAC_N.t726 VSS 0.105768f
C16057 VDAC_N.n1110 VSS 0.132739f
C16058 VDAC_N.t101 VSS 0.105768f
C16059 VDAC_N.n1111 VSS 0.132739f
C16060 VDAC_N.t1661 VSS 0.105768f
C16061 VDAC_N.n1112 VSS 0.132739f
C16062 VDAC_N.t25 VSS 0.105768f
C16063 VDAC_N.n1113 VSS 0.132739f
C16064 VDAC_N.t789 VSS 0.105768f
C16065 VDAC_N.n1114 VSS 0.132739f
C16066 VDAC_N.t1017 VSS 0.105768f
C16067 VDAC_N.n1115 VSS 0.132739f
C16068 VDAC_N.t685 VSS 0.105768f
C16069 VDAC_N.n1116 VSS 0.132739f
C16070 VDAC_N.t1903 VSS 0.105768f
C16071 VDAC_N.n1117 VSS 0.132739f
C16072 VDAC_N.t1227 VSS 0.105768f
C16073 VDAC_N.n1118 VSS 0.132739f
C16074 VDAC_N.t445 VSS 0.105768f
C16075 VDAC_N.n1119 VSS 0.132739f
C16076 VDAC_N.t1516 VSS 0.105768f
C16077 VDAC_N.n1120 VSS 0.132739f
C16078 VDAC_N.t125 VSS 0.105768f
C16079 VDAC_N.n1121 VSS 0.132739f
C16080 VDAC_N.t2041 VSS 0.105768f
C16081 VDAC_N.n1122 VSS 0.132739f
C16082 VDAC_N.t480 VSS 0.105768f
C16083 VDAC_N.n1123 VSS 0.132739f
C16084 VDAC_N.t1929 VSS 0.105768f
C16085 VDAC_N.n1124 VSS 0.12675f
C16086 VDAC_N.t1587 VSS 0.105768f
C16087 VDAC_N.n1125 VSS 0.132739f
C16088 VDAC_N.t1628 VSS 0.105768f
C16089 VDAC_N.n1126 VSS 0.132739f
C16090 VDAC_N.t209 VSS 0.105768f
C16091 VDAC_N.n1127 VSS 0.132739f
C16092 VDAC_N.t981 VSS 0.105768f
C16093 VDAC_N.n1128 VSS 0.132739f
C16094 VDAC_N.t1908 VSS 0.105768f
C16095 VDAC_N.n1129 VSS 0.132739f
C16096 VDAC_N.t1833 VSS 0.105768f
C16097 VDAC_N.n1130 VSS 0.132739f
C16098 VDAC_N.t1004 VSS 0.105768f
C16099 VDAC_N.n1131 VSS 0.132739f
C16100 VDAC_N.t102 VSS 0.105768f
C16101 VDAC_N.n1132 VSS 0.132739f
C16102 VDAC_N.t1078 VSS 0.105768f
C16103 VDAC_N.n1133 VSS 0.132739f
C16104 VDAC_N.t1960 VSS 0.105768f
C16105 VDAC_N.n1134 VSS 0.132739f
C16106 VDAC_N.t1961 VSS 0.105768f
C16107 VDAC_N.n1135 VSS 0.132739f
C16108 VDAC_N.t1512 VSS 0.105768f
C16109 VDAC_N.n1136 VSS 0.132739f
C16110 VDAC_N.t238 VSS 0.105768f
C16111 VDAC_N.n1137 VSS 0.132739f
C16112 VDAC_N.t2130 VSS 0.105768f
C16113 VDAC_N.n1138 VSS 0.132739f
C16114 VDAC_N.t1008 VSS 0.105768f
C16115 VDAC_N.n1139 VSS 0.132739f
C16116 VDAC_N.t27 VSS 0.105768f
C16117 VDAC_N.n1140 VSS 0.132739f
C16118 VDAC_N.t1536 VSS 0.105768f
C16119 VDAC_N.n1141 VSS 0.132739f
C16120 VDAC_N.t450 VSS 0.105768f
C16121 VDAC_N.n1142 VSS 0.132739f
C16122 VDAC_N.t1445 VSS 0.105768f
C16123 VDAC_N.n1143 VSS 0.132739f
C16124 VDAC_N.t1494 VSS 0.105768f
C16125 VDAC_N.n1144 VSS 0.132739f
C16126 VDAC_N.t103 VSS 0.105768f
C16127 VDAC_N.n1145 VSS 0.132739f
C16128 VDAC_N.t1278 VSS 0.105768f
C16129 VDAC_N.n1146 VSS 0.132739f
C16130 VDAC_N.t1115 VSS 0.105768f
C16131 VDAC_N.n1147 VSS 0.132739f
C16132 VDAC_N.t1581 VSS 0.105768f
C16133 VDAC_N.n1148 VSS 0.132739f
C16134 VDAC_N.t1770 VSS 0.105768f
C16135 VDAC_N.n1149 VSS 0.132739f
C16136 VDAC_N.t1469 VSS 0.105768f
C16137 VDAC_N.n1150 VSS 0.132739f
C16138 VDAC_N.t979 VSS 0.105768f
C16139 VDAC_N.n1151 VSS 0.132739f
C16140 VDAC_N.t335 VSS 0.105768f
C16141 VDAC_N.n1152 VSS 0.132739f
C16142 VDAC_N.t1827 VSS 0.105768f
C16143 VDAC_N.n1153 VSS 0.132739f
C16144 VDAC_N.t1147 VSS 0.105768f
C16145 VDAC_N.n1154 VSS 0.132739f
C16146 VDAC_N.t1609 VSS 0.105768f
C16147 VDAC_N.n1155 VSS 0.132739f
C16148 VDAC_N.t2126 VSS 0.105768f
C16149 VDAC_N.n1156 VSS 0.132739f
C16150 VDAC_N.t1501 VSS 0.105768f
C16151 VDAC_N.n1157 VSS 0.132739f
C16152 VDAC_N.t509 VSS 0.105768f
C16153 VDAC_N.n1158 VSS 0.132739f
C16154 VDAC_N.t2116 VSS 0.105768f
C16155 VDAC_N.n1159 VSS 0.132739f
C16156 VDAC_N.t485 VSS 0.105768f
C16157 VDAC_N.n1160 VSS 0.132739f
C16158 VDAC_N.t628 VSS 0.105768f
C16159 VDAC_N.n1161 VSS 0.132739f
C16160 VDAC_N.t1643 VSS 0.105768f
C16161 VDAC_N.n1162 VSS 0.132739f
C16162 VDAC_N.t700 VSS 0.105768f
C16163 VDAC_N.n1163 VSS 0.132739f
C16164 VDAC_N.t1040 VSS 0.105768f
C16165 VDAC_N.n1164 VSS 0.132739f
C16166 VDAC_N.t2135 VSS 0.105768f
C16167 VDAC_N.n1165 VSS 0.132739f
C16168 VDAC_N.t1952 VSS 0.105768f
C16169 VDAC_N.n1166 VSS 0.132739f
C16170 VDAC_N.t982 VSS 0.105768f
C16171 VDAC_N.n1167 VSS 0.132739f
C16172 VDAC_N.t560 VSS 0.105768f
C16173 VDAC_N.n1168 VSS 0.132739f
C16174 VDAC_N.t1486 VSS 0.105768f
C16175 VDAC_N.n1169 VSS 0.132739f
C16176 VDAC_N.t681 VSS 0.105768f
C16177 VDAC_N.n1170 VSS 0.132739f
C16178 VDAC_N.t646 VSS 0.105768f
C16179 VDAC_N.n1171 VSS 0.132739f
C16180 VDAC_N.t1111 VSS 0.105768f
C16181 VDAC_N.n1172 VSS 0.132739f
C16182 VDAC_N.t2072 VSS 0.105768f
C16183 VDAC_N.n1173 VSS 0.132739f
C16184 VDAC_N.t1994 VSS 0.105768f
C16185 VDAC_N.n1174 VSS 0.132739f
C16186 VDAC_N.t747 VSS 0.105768f
C16187 VDAC_N.n1175 VSS 0.132739f
C16188 VDAC_N.t82 VSS 0.105768f
C16189 VDAC_N.n1176 VSS 0.132739f
C16190 VDAC_N.t1365 VSS 0.105768f
C16191 VDAC_N.n1177 VSS 0.132739f
C16192 VDAC_N.t1821 VSS 0.105768f
C16193 VDAC_N.n1178 VSS 0.132739f
C16194 VDAC_N.t307 VSS 0.105768f
C16195 VDAC_N.n1179 VSS 0.132739f
C16196 VDAC_N.t1711 VSS 0.105768f
C16197 VDAC_N.n1180 VSS 0.132739f
C16198 VDAC_N.t1034 VSS 0.105768f
C16199 VDAC_N.n1181 VSS 0.132739f
C16200 VDAC_N.t763 VSS 0.105768f
C16201 VDAC_N.n1182 VSS 0.132739f
C16202 VDAC_N.t1047 VSS 0.105768f
C16203 VDAC_N.n1183 VSS 0.132739f
C16204 VDAC_N.t369 VSS 0.105768f
C16205 VDAC_N.n1184 VSS 0.132739f
C16206 VDAC_N.t941 VSS 0.105768f
C16207 VDAC_N.n1185 VSS 0.132739f
C16208 VDAC_N.t2100 VSS 0.105768f
C16209 VDAC_N.n1186 VSS 0.132739f
C16210 VDAC_N.t1743 VSS 0.105768f
C16211 VDAC_N.n1187 VSS 0.12675f
C16212 VDAC_N.t1598 VSS 0.105768f
C16213 VDAC_N.n1188 VSS 0.132739f
C16214 VDAC_N.t705 VSS 0.105768f
C16215 VDAC_N.n1189 VSS 0.132739f
C16216 VDAC_N.t690 VSS 0.105768f
C16217 VDAC_N.n1190 VSS 0.132739f
C16218 VDAC_N.t99 VSS 0.105768f
C16219 VDAC_N.n1191 VSS 0.132739f
C16220 VDAC_N.t827 VSS 0.105768f
C16221 VDAC_N.n1192 VSS 0.132739f
C16222 VDAC_N.t542 VSS 0.105768f
C16223 VDAC_N.n1193 VSS 0.132739f
C16224 VDAC_N.t773 VSS 0.105768f
C16225 VDAC_N.n1194 VSS 0.132739f
C16226 VDAC_N.t515 VSS 0.105768f
C16227 VDAC_N.n1195 VSS 0.132739f
C16228 VDAC_N.t721 VSS 0.105768f
C16229 VDAC_N.n1196 VSS 0.132739f
C16230 VDAC_N.t951 VSS 0.105768f
C16231 VDAC_N.n1197 VSS 0.132739f
C16232 VDAC_N.t1193 VSS 0.105768f
C16233 VDAC_N.n1198 VSS 0.132739f
C16234 VDAC_N.t461 VSS 0.105768f
C16235 VDAC_N.n1199 VSS 0.132739f
C16236 VDAC_N.t2108 VSS 0.105768f
C16237 VDAC_N.n1200 VSS 0.132739f
C16238 VDAC_N.t1011 VSS 0.105768f
C16239 VDAC_N.n1201 VSS 0.132739f
C16240 VDAC_N.t1224 VSS 0.105768f
C16241 VDAC_N.n1202 VSS 0.132739f
C16242 VDAC_N.t894 VSS 0.105768f
C16243 VDAC_N.n1203 VSS 0.132739f
C16244 VDAC_N.t1508 VSS 0.105768f
C16245 VDAC_N.n1204 VSS 0.132739f
C16246 VDAC_N.t1322 VSS 0.105768f
C16247 VDAC_N.n1205 VSS 0.132739f
C16248 VDAC_N.t1251 VSS 0.105768f
C16249 VDAC_N.n1206 VSS 0.132739f
C16250 VDAC_N.t1110 VSS 0.105768f
C16251 VDAC_N.n1207 VSS 0.132739f
C16252 VDAC_N.t2042 VSS 0.105768f
C16253 VDAC_N.n1208 VSS 0.132739f
C16254 VDAC_N.t904 VSS 0.105768f
C16255 VDAC_N.n1209 VSS 0.132739f
C16256 VDAC_N.t926 VSS 0.105768f
C16257 VDAC_N.n1210 VSS 0.132739f
C16258 VDAC_N.t1393 VSS 0.105768f
C16259 VDAC_N.n1211 VSS 0.132739f
C16260 VDAC_N.t366 VSS 0.105768f
C16261 VDAC_N.n1212 VSS 0.132739f
C16262 VDAC_N.t1279 VSS 0.105768f
C16263 VDAC_N.n1213 VSS 0.132739f
C16264 VDAC_N.t457 VSS 0.105768f
C16265 VDAC_N.n1214 VSS 0.132739f
C16266 VDAC_N.t1062 VSS 0.105768f
C16267 VDAC_N.n1215 VSS 0.132739f
C16268 VDAC_N.t1637 VSS 0.105768f
C16269 VDAC_N.n1216 VSS 0.132739f
C16270 VDAC_N.t1886 VSS 0.105768f
C16271 VDAC_N.n1217 VSS 0.132739f
C16272 VDAC_N.t1419 VSS 0.105768f
C16273 VDAC_N.n1218 VSS 0.132739f
C16274 VDAC_N.t517 VSS 0.105768f
C16275 VDAC_N.n1219 VSS 0.132739f
C16276 VDAC_N.t1313 VSS 0.105768f
C16277 VDAC_N.n1220 VSS 0.132739f
C16278 VDAC_N.t463 VSS 0.105768f
C16279 VDAC_N.n1221 VSS 0.132739f
C16280 VDAC_N.t1164 VSS 0.105768f
C16281 VDAC_N.n1222 VSS 0.132739f
C16282 VDAC_N.t1665 VSS 0.105768f
C16283 VDAC_N.n1223 VSS 0.132739f
C16284 VDAC_N.t2125 VSS 0.105768f
C16285 VDAC_N.n1224 VSS 0.132739f
C16286 VDAC_N.t739 VSS 0.105768f
C16287 VDAC_N.n1225 VSS 0.132739f
C16288 VDAC_N.t2011 VSS 0.105768f
C16289 VDAC_N.n1226 VSS 0.132739f
C16290 VDAC_N.t1288 VSS 0.105768f
C16291 VDAC_N.n1227 VSS 0.132739f
C16292 VDAC_N.t1887 VSS 0.105768f
C16293 VDAC_N.n1228 VSS 0.132739f
C16294 VDAC_N.t1192 VSS 0.105768f
C16295 VDAC_N.n1229 VSS 0.132739f
C16296 VDAC_N.t1542 VSS 0.105768f
C16297 VDAC_N.n1230 VSS 0.132739f
C16298 VDAC_N.t620 VSS 0.105768f
C16299 VDAC_N.n1231 VSS 0.132739f
C16300 VDAC_N.t1102 VSS 0.105768f
C16301 VDAC_N.n1232 VSS 0.132739f
C16302 VDAC_N.t581 VSS 0.105768f
C16303 VDAC_N.n1233 VSS 0.132739f
C16304 VDAC_N.t1744 VSS 0.105768f
C16305 VDAC_N.n1234 VSS 0.132739f
C16306 VDAC_N.t1814 VSS 0.105768f
C16307 VDAC_N.n1235 VSS 0.132739f
C16308 VDAC_N.t664 VSS 0.105768f
C16309 VDAC_N.n1236 VSS 0.132739f
C16310 VDAC_N.t1606 VSS 0.105768f
C16311 VDAC_N.n1237 VSS 0.132739f
C16312 VDAC_N.t1273 VSS 0.105768f
C16313 VDAC_N.n1238 VSS 0.132739f
C16314 VDAC_N.t694 VSS 0.105768f
C16315 VDAC_N.n1239 VSS 0.132739f
C16316 VDAC_N.t1167 VSS 0.105768f
C16317 VDAC_N.n1240 VSS 0.132739f
C16318 VDAC_N.t1631 VSS 0.105768f
C16319 VDAC_N.n1241 VSS 0.132739f
C16320 VDAC_N.t1878 VSS 0.105768f
C16321 VDAC_N.n1242 VSS 0.132739f
C16322 VDAC_N.t1521 VSS 0.105768f
C16323 VDAC_N.n1243 VSS 0.132739f
C16324 VDAC_N.t434 VSS 0.105768f
C16325 VDAC_N.n1244 VSS 0.132739f
C16326 VDAC_N.t1311 VSS 0.105768f
C16327 VDAC_N.n1245 VSS 0.132739f
C16328 VDAC_N.t1879 VSS 0.105768f
C16329 VDAC_N.n1246 VSS 0.132739f
C16330 VDAC_N.t1197 VSS 0.105768f
C16331 VDAC_N.n1247 VSS 0.132739f
C16332 VDAC_N.t845 VSS 0.105768f
C16333 VDAC_N.n1248 VSS 0.132739f
C16334 VDAC_N.t1132 VSS 0.105768f
C16335 VDAC_N.n1249 VSS 0.132739f
C16336 VDAC_N.t1551 VSS 0.105768f
C16337 VDAC_N.n1250 VSS 0.12675f
C16338 VDAC_N.t265 VSS 0.105768f
C16339 VDAC_N.n1251 VSS 0.132739f
C16340 VDAC_N.t192 VSS 0.105768f
C16341 VDAC_N.n1252 VSS 0.132739f
C16342 VDAC_N.t923 VSS 0.105768f
C16343 VDAC_N.n1253 VSS 0.132739f
C16344 VDAC_N.t940 VSS 0.105768f
C16345 VDAC_N.n1254 VSS 0.132739f
C16346 VDAC_N.t1186 VSS 0.105768f
C16347 VDAC_N.n1255 VSS 0.132739f
C16348 VDAC_N.t16 VSS 0.105768f
C16349 VDAC_N.n1256 VSS 0.132739f
C16350 VDAC_N.t1912 VSS 0.105768f
C16351 VDAC_N.n1257 VSS 0.132739f
C16352 VDAC_N.t498 VSS 0.105768f
C16353 VDAC_N.n1258 VSS 0.132739f
C16354 VDAC_N.t744 VSS 0.105768f
C16355 VDAC_N.n1259 VSS 0.132739f
C16356 VDAC_N.t854 VSS 0.105768f
C16357 VDAC_N.n1260 VSS 0.132739f
C16358 VDAC_N.t1188 VSS 0.105768f
C16359 VDAC_N.n1261 VSS 0.132739f
C16360 VDAC_N.t1450 VSS 0.105768f
C16361 VDAC_N.n1262 VSS 0.132739f
C16362 VDAC_N.t65 VSS 0.105768f
C16363 VDAC_N.n1263 VSS 0.132739f
C16364 VDAC_N.t1142 VSS 0.105768f
C16365 VDAC_N.n1264 VSS 0.132739f
C16366 VDAC_N.t538 VSS 0.105768f
C16367 VDAC_N.n1265 VSS 0.132739f
C16368 VDAC_N.t1619 VSS 0.105768f
C16369 VDAC_N.n1266 VSS 0.132739f
C16370 VDAC_N.t142 VSS 0.105768f
C16371 VDAC_N.n1267 VSS 0.132739f
C16372 VDAC_N.t1407 VSS 0.105768f
C16373 VDAC_N.n1268 VSS 0.132739f
C16374 VDAC_N.t513 VSS 0.105768f
C16375 VDAC_N.n1269 VSS 0.132739f
C16376 VDAC_N.t345 VSS 0.105768f
C16377 VDAC_N.n1270 VSS 0.132739f
C16378 VDAC_N.t1757 VSS 0.105768f
C16379 VDAC_N.n1271 VSS 0.132739f
C16380 VDAC_N.t1185 VSS 0.105768f
C16381 VDAC_N.n1272 VSS 0.132739f
C16382 VDAC_N.t1653 VSS 0.105768f
C16383 VDAC_N.n1273 VSS 0.132739f
C16384 VDAC_N.t2107 VSS 0.105768f
C16385 VDAC_N.n1274 VSS 0.132739f
C16386 VDAC_N.t379 VSS 0.105768f
C16387 VDAC_N.n1275 VSS 0.132739f
C16388 VDAC_N.t1997 VSS 0.105768f
C16389 VDAC_N.n1276 VSS 0.132739f
C16390 VDAC_N.t1240 VSS 0.105768f
C16391 VDAC_N.n1277 VSS 0.132739f
C16392 VDAC_N.t907 VSS 0.105768f
C16393 VDAC_N.n1278 VSS 0.132739f
C16394 VDAC_N.t1556 VSS 0.105768f
C16395 VDAC_N.n1279 VSS 0.132739f
C16396 VDAC_N.t1681 VSS 0.105768f
C16397 VDAC_N.n1280 VSS 0.132739f
C16398 VDAC_N.t1417 VSS 0.105768f
C16399 VDAC_N.n1281 VSS 0.132739f
C16400 VDAC_N.t1122 VSS 0.105768f
C16401 VDAC_N.n1282 VSS 0.132739f
C16402 VDAC_N.t1029 VSS 0.105768f
C16403 VDAC_N.n1283 VSS 0.132739f
C16404 VDAC_N.t680 VSS 0.105768f
C16405 VDAC_N.n1284 VSS 0.132739f
C16406 VDAC_N.t426 VSS 0.105768f
C16407 VDAC_N.n1285 VSS 0.132739f
C16408 VDAC_N.t1796 VSS 0.105768f
C16409 VDAC_N.n1286 VSS 0.132739f
C16410 VDAC_N.t198 VSS 0.105768f
C16411 VDAC_N.n1287 VSS 0.132739f
C16412 VDAC_N.t796 VSS 0.105768f
C16413 VDAC_N.n1288 VSS 0.132739f
C16414 VDAC_N.t1170 VSS 0.105768f
C16415 VDAC_N.n1289 VSS 0.132739f
C16416 VDAC_N.t2102 VSS 0.105768f
C16417 VDAC_N.n1290 VSS 0.132739f
C16418 VDAC_N.t920 VSS 0.105768f
C16419 VDAC_N.n1291 VSS 0.132739f
C16420 VDAC_N.t2054 VSS 0.105768f
C16421 VDAC_N.n1292 VSS 0.132739f
C16422 VDAC_N.t213 VSS 0.105768f
C16423 VDAC_N.n1293 VSS 0.132739f
C16424 VDAC_N.t1626 VSS 0.105768f
C16425 VDAC_N.n1294 VSS 0.132739f
C16426 VDAC_N.t1291 VSS 0.105768f
C16427 VDAC_N.n1295 VSS 0.132739f
C16428 VDAC_N.t1861 VSS 0.105768f
C16429 VDAC_N.n1296 VSS 0.132739f
C16430 VDAC_N.t1179 VSS 0.105768f
C16431 VDAC_N.n1297 VSS 0.132739f
C16432 VDAC_N.t1649 VSS 0.105768f
C16433 VDAC_N.n1298 VSS 0.132739f
C16434 VDAC_N.t158 VSS 0.105768f
C16435 VDAC_N.n1299 VSS 0.132739f
C16436 VDAC_N.t1537 VSS 0.105768f
C16437 VDAC_N.n1300 VSS 0.132739f
C16438 VDAC_N.t519 VSS 0.105768f
C16439 VDAC_N.n1301 VSS 0.132739f
C16440 VDAC_N.t727 VSS 0.105768f
C16441 VDAC_N.n1302 VSS 0.132739f
C16442 VDAC_N.t959 VSS 0.105768f
C16443 VDAC_N.n1303 VSS 0.132739f
C16444 VDAC_N.t212 VSS 0.105768f
C16445 VDAC_N.n1304 VSS 0.132739f
C16446 VDAC_N.t853 VSS 0.105768f
C16447 VDAC_N.n1305 VSS 0.132739f
C16448 VDAC_N.t1292 VSS 0.105768f
C16449 VDAC_N.n1306 VSS 0.132739f
C16450 VDAC_N.t31 VSS 0.105768f
C16451 VDAC_N.n1307 VSS 0.132739f
C16452 VDAC_N.t1027 VSS 0.105768f
C16453 VDAC_N.n1308 VSS 0.132739f
C16454 VDAC_N.t464 VSS 0.105768f
C16455 VDAC_N.n1309 VSS 0.132739f
C16456 VDAC_N.t87 VSS 0.105768f
C16457 VDAC_N.n1310 VSS 0.132739f
C16458 VDAC_N.t900 VSS 0.105768f
C16459 VDAC_N.n1311 VSS 0.132739f
C16460 VDAC_N.t1614 VSS 0.105768f
C16461 VDAC_N.n1312 VSS 0.132739f
C16462 VDAC_N.t1708 VSS 0.105768f
C16463 VDAC_N.n1313 VSS 0.12675f
C16464 VDAC_N.t1151 VSS 0.105768f
C16465 VDAC_N.n1314 VSS 0.132739f
C16466 VDAC_N.t239 VSS 0.105768f
C16467 VDAC_N.n1315 VSS 0.132739f
C16468 VDAC_N.t534 VSS 0.105768f
C16469 VDAC_N.n1316 VSS 0.132739f
C16470 VDAC_N.t397 VSS 0.105768f
C16471 VDAC_N.n1317 VSS 0.132739f
C16472 VDAC_N.t269 VSS 0.105768f
C16473 VDAC_N.n1318 VSS 0.132739f
C16474 VDAC_N.t1401 VSS 0.105768f
C16475 VDAC_N.n1319 VSS 0.132739f
C16476 VDAC_N.t943 VSS 0.105768f
C16477 VDAC_N.n1320 VSS 0.132739f
C16478 VDAC_N.t1252 VSS 0.105768f
C16479 VDAC_N.n1321 VSS 0.132739f
C16480 VDAC_N.t459 VSS 0.105768f
C16481 VDAC_N.n1322 VSS 0.132739f
C16482 VDAC_N.t124 VSS 0.105768f
C16483 VDAC_N.n1323 VSS 0.132739f
C16484 VDAC_N.t1535 VSS 0.105768f
C16485 VDAC_N.n1324 VSS 0.132739f
C16486 VDAC_N.t1063 VSS 0.105768f
C16487 VDAC_N.n1325 VSS 0.132739f
C16488 VDAC_N.t1648 VSS 0.105768f
C16489 VDAC_N.n1326 VSS 0.132739f
C16490 VDAC_N.t1472 VSS 0.105768f
C16491 VDAC_N.n1327 VSS 0.132739f
C16492 VDAC_N.t442 VSS 0.105768f
C16493 VDAC_N.n1328 VSS 0.132739f
C16494 VDAC_N.t1427 VSS 0.105768f
C16495 VDAC_N.n1329 VSS 0.132739f
C16496 VDAC_N.t1458 VSS 0.105768f
C16497 VDAC_N.n1330 VSS 0.132739f
C16498 VDAC_N.t621 VSS 0.105768f
C16499 VDAC_N.n1331 VSS 0.132739f
C16500 VDAC_N.t1781 VSS 0.105768f
C16501 VDAC_N.n1332 VSS 0.132739f
C16502 VDAC_N.t563 VSS 0.105768f
C16503 VDAC_N.n1333 VSS 0.132739f
C16504 VDAC_N.t1565 VSS 0.105768f
C16505 VDAC_N.n1334 VSS 0.132739f
C16506 VDAC_N.t514 VSS 0.105768f
C16507 VDAC_N.n1335 VSS 0.132739f
C16508 VDAC_N.t743 VSS 0.105768f
C16509 VDAC_N.n1336 VSS 0.132739f
C16510 VDAC_N.t1917 VSS 0.105768f
C16511 VDAC_N.n1337 VSS 0.132739f
C16512 VDAC_N.t1239 VSS 0.105768f
C16513 VDAC_N.n1338 VSS 0.132739f
C16514 VDAC_N.t1811 VSS 0.105768f
C16515 VDAC_N.n1339 VSS 0.132739f
C16516 VDAC_N.t876 VSS 0.105768f
C16517 VDAC_N.n1340 VSS 0.132739f
C16518 VDAC_N.t77 VSS 0.105768f
C16519 VDAC_N.n1341 VSS 0.132739f
C16520 VDAC_N.t1436 VSS 0.105768f
C16521 VDAC_N.n1342 VSS 0.132739f
C16522 VDAC_N.t1485 VSS 0.105768f
C16523 VDAC_N.n1343 VSS 0.132739f
C16524 VDAC_N.t267 VSS 0.105768f
C16525 VDAC_N.n1344 VSS 0.132739f
C16526 VDAC_N.t1440 VSS 0.105768f
C16527 VDAC_N.n1345 VSS 0.132739f
C16528 VDAC_N.t1843 VSS 0.105768f
C16529 VDAC_N.n1346 VSS 0.132739f
C16530 VDAC_N.t2124 VSS 0.105768f
C16531 VDAC_N.n1347 VSS 0.132739f
C16532 VDAC_N.t178 VSS 0.105768f
C16533 VDAC_N.n1348 VSS 0.132739f
C16534 VDAC_N.t1052 VSS 0.105768f
C16535 VDAC_N.n1349 VSS 0.132739f
C16536 VDAC_N.t1016 VSS 0.105768f
C16537 VDAC_N.n1350 VSS 0.132739f
C16538 VDAC_N.t1973 VSS 0.105768f
C16539 VDAC_N.n1351 VSS 0.132739f
C16540 VDAC_N.t792 VSS 0.105768f
C16541 VDAC_N.n1352 VSS 0.132739f
C16542 VDAC_N.t1726 VSS 0.105768f
C16543 VDAC_N.n1353 VSS 0.132739f
C16544 VDAC_N.t2052 VSS 0.105768f
C16545 VDAC_N.n1354 VSS 0.132739f
C16546 VDAC_N.t438 VSS 0.105768f
C16547 VDAC_N.n1355 VSS 0.132739f
C16548 VDAC_N.t673 VSS 0.105768f
C16549 VDAC_N.n1356 VSS 0.132739f
C16550 VDAC_N.t1234 VSS 0.105768f
C16551 VDAC_N.n1357 VSS 0.132739f
C16552 VDAC_N.t1093 VSS 0.105768f
C16553 VDAC_N.n1358 VSS 0.132739f
C16554 VDAC_N.t1669 VSS 0.105768f
C16555 VDAC_N.n1359 VSS 0.132739f
C16556 VDAC_N.t510 VSS 0.105768f
C16557 VDAC_N.n1360 VSS 0.132739f
C16558 VDAC_N.t1453 VSS 0.105768f
C16559 VDAC_N.n1361 VSS 0.132739f
C16560 VDAC_N.t1734 VSS 0.105768f
C16561 VDAC_N.n1362 VSS 0.132739f
C16562 VDAC_N.t1351 VSS 0.105768f
C16563 VDAC_N.n1363 VSS 0.132739f
C16564 VDAC_N.t139 VSS 0.105768f
C16565 VDAC_N.n1364 VSS 0.132739f
C16566 VDAC_N.t631 VSS 0.105768f
C16567 VDAC_N.n1365 VSS 0.132739f
C16568 VDAC_N.t865 VSS 0.105768f
C16569 VDAC_N.n1366 VSS 0.132739f
C16570 VDAC_N.t1244 VSS 0.105768f
C16571 VDAC_N.n1367 VSS 0.132739f
C16572 VDAC_N.t1481 VSS 0.105768f
C16573 VDAC_N.n1368 VSS 0.132739f
C16574 VDAC_N.t2049 VSS 0.105768f
C16575 VDAC_N.n1369 VSS 0.132739f
C16576 VDAC_N.t703 VSS 0.105768f
C16577 VDAC_N.n1370 VSS 0.132739f
C16578 VDAC_N.t933 VSS 0.105768f
C16579 VDAC_N.n1371 VSS 0.132739f
C16580 VDAC_N.t1956 VSS 0.105768f
C16581 VDAC_N.n1372 VSS 0.132739f
C16582 VDAC_N.t1727 VSS 0.105768f
C16583 VDAC_N.n1373 VSS 0.132739f
C16584 VDAC_N.t1564 VSS 0.105768f
C16585 VDAC_N.n1374 VSS 0.132739f
C16586 VDAC_N.t1218 VSS 0.105768f
C16587 VDAC_N.n1375 VSS 0.132739f
C16588 VDAC_N.t541 VSS 0.105768f
C16589 VDAC_N.n1376 VSS 0.12675f
C16590 VDAC_N.t428 VSS 0.105768f
C16591 VDAC_N.n1377 VSS 0.132739f
C16592 VDAC_N.t194 VSS 0.105768f
C16593 VDAC_N.n1378 VSS 0.132739f
C16594 VDAC_N.t348 VSS 0.105768f
C16595 VDAC_N.n1379 VSS 0.132739f
C16596 VDAC_N.t1864 VSS 0.105768f
C16597 VDAC_N.n1380 VSS 0.132739f
C16598 VDAC_N.t258 VSS 0.105768f
C16599 VDAC_N.n1381 VSS 0.132739f
C16600 VDAC_N.t1408 VSS 0.105768f
C16601 VDAC_N.n1382 VSS 0.132739f
C16602 VDAC_N.t1646 VSS 0.105768f
C16603 VDAC_N.n1383 VSS 0.132739f
C16604 VDAC_N.t667 VSS 0.105768f
C16605 VDAC_N.n1384 VSS 0.132739f
C16606 VDAC_N.t1418 VSS 0.105768f
C16607 VDAC_N.n1385 VSS 0.132739f
C16608 VDAC_N.t611 VSS 0.105768f
C16609 VDAC_N.n1386 VSS 0.132739f
C16610 VDAC_N.t1984 VSS 0.105768f
C16611 VDAC_N.n1387 VSS 0.132739f
C16612 VDAC_N.t21 VSS 0.105768f
C16613 VDAC_N.n1388 VSS 0.132739f
C16614 VDAC_N.t123 VSS 0.105768f
C16615 VDAC_N.n1389 VSS 0.132739f
C16616 VDAC_N.t1113 VSS 0.105768f
C16617 VDAC_N.n1390 VSS 0.132739f
C16618 VDAC_N.t803 VSS 0.105768f
C16619 VDAC_N.n1391 VSS 0.132739f
C16620 VDAC_N.t550 VSS 0.105768f
C16621 VDAC_N.n1392 VSS 0.132739f
C16622 VDAC_N.t73 VSS 0.105768f
C16623 VDAC_N.n1393 VSS 0.132739f
C16624 VDAC_N.t1927 VSS 0.105768f
C16625 VDAC_N.n1394 VSS 0.132739f
C16626 VDAC_N.t112 VSS 0.105768f
C16627 VDAC_N.n1395 VSS 0.132739f
C16628 VDAC_N.t477 VSS 0.105768f
C16629 VDAC_N.n1396 VSS 0.132739f
C16630 VDAC_N.t1900 VSS 0.105768f
C16631 VDAC_N.n1397 VSS 0.132739f
C16632 VDAC_N.t871 VSS 0.105768f
C16633 VDAC_N.n1398 VSS 0.132739f
C16634 VDAC_N.t22 VSS 0.105768f
C16635 VDAC_N.n1399 VSS 0.132739f
C16636 VDAC_N.t1928 VSS 0.105768f
C16637 VDAC_N.n1400 VSS 0.132739f
C16638 VDAC_N.t1951 VSS 0.105768f
C16639 VDAC_N.n1401 VSS 0.132739f
C16640 VDAC_N.t1480 VSS 0.105768f
C16641 VDAC_N.n1402 VSS 0.132739f
C16642 VDAC_N.t1690 VSS 0.105768f
C16643 VDAC_N.n1403 VSS 0.132739f
C16644 VDAC_N.t324 VSS 0.105768f
C16645 VDAC_N.n1404 VSS 0.132739f
C16646 VDAC_N.t1466 VSS 0.105768f
C16647 VDAC_N.n1405 VSS 0.132739f
C16648 VDAC_N.t1340 VSS 0.105768f
C16649 VDAC_N.n1406 VSS 0.132739f
C16650 VDAC_N.t2048 VSS 0.105768f
C16651 VDAC_N.n1407 VSS 0.132739f
C16652 VDAC_N.t1103 VSS 0.105768f
C16653 VDAC_N.n1408 VSS 0.132739f
C16654 VDAC_N.t1624 VSS 0.105768f
C16655 VDAC_N.n1409 VSS 0.132739f
C16656 VDAC_N.t886 VSS 0.105768f
C16657 VDAC_N.n1410 VSS 0.132739f
C16658 VDAC_N.t1359 VSS 0.105768f
C16659 VDAC_N.n1411 VSS 0.132739f
C16660 VDAC_N.t782 VSS 0.105768f
C16661 VDAC_N.n1412 VSS 0.132739f
C16662 VDAC_N.t635 VSS 0.105768f
C16663 VDAC_N.n1413 VSS 0.132739f
C16664 VDAC_N.t1094 VSS 0.105768f
C16665 VDAC_N.n1414 VSS 0.132739f
C16666 VDAC_N.t1131 VSS 0.105768f
C16667 VDAC_N.n1415 VSS 0.132739f
C16668 VDAC_N.t813 VSS 0.105768f
C16669 VDAC_N.n1416 VSS 0.132739f
C16670 VDAC_N.t518 VSS 0.105768f
C16671 VDAC_N.n1417 VSS 0.132739f
C16672 VDAC_N.t1571 VSS 0.105768f
C16673 VDAC_N.n1418 VSS 0.132739f
C16674 VDAC_N.t1031 VSS 0.105768f
C16675 VDAC_N.n1419 VSS 0.132739f
C16676 VDAC_N.t1363 VSS 0.105768f
C16677 VDAC_N.n1420 VSS 0.132739f
C16678 VDAC_N.t1819 VSS 0.105768f
C16679 VDAC_N.n1421 VSS 0.132739f
C16680 VDAC_N.t1828 VSS 0.105768f
C16681 VDAC_N.n1422 VSS 0.132739f
C16682 VDAC_N.t1709 VSS 0.105768f
C16683 VDAC_N.n1423 VSS 0.132739f
C16684 VDAC_N.t14 VSS 0.105768f
C16685 VDAC_N.n1424 VSS 0.132739f
C16686 VDAC_N.t225 VSS 0.105768f
C16687 VDAC_N.n1425 VSS 0.132739f
C16688 VDAC_N.t1045 VSS 0.105768f
C16689 VDAC_N.n1426 VSS 0.132739f
C16690 VDAC_N.t1464 VSS 0.105768f
C16691 VDAC_N.n1427 VSS 0.132739f
C16692 VDAC_N.t1947 VSS 0.105768f
C16693 VDAC_N.n1428 VSS 0.132739f
C16694 VDAC_N.t2084 VSS 0.105768f
C16695 VDAC_N.n1429 VSS 0.132739f
C16696 VDAC_N.t1454 VSS 0.105768f
C16697 VDAC_N.n1430 VSS 0.132739f
C16698 VDAC_N.t636 VSS 0.105768f
C16699 VDAC_N.n1431 VSS 0.132739f
C16700 VDAC_N.t66 VSS 0.105768f
C16701 VDAC_N.n1432 VSS 0.132739f
C16702 VDAC_N.t2093 VSS 0.105768f
C16703 VDAC_N.n1433 VSS 0.132739f
C16704 VDAC_N.t1608 VSS 0.105768f
C16705 VDAC_N.n1434 VSS 0.132739f
C16706 VDAC_N.t998 VSS 0.105768f
C16707 VDAC_N.n1435 VSS 0.132739f
C16708 VDAC_N.t600 VSS 0.105768f
C16709 VDAC_N.n1436 VSS 0.132739f
C16710 VDAC_N.t122 VSS 0.105768f
C16711 VDAC_N.n1437 VSS 0.132739f
C16712 VDAC_N.t1355 VSS 0.105768f
C16713 VDAC_N.n1438 VSS 0.132739f
C16714 VDAC_N.t1298 VSS 0.105768f
C16715 VDAC_N.n1439 VSS 0.12675f
C16716 VDAC_N.t1491 VSS 0.105768f
C16717 VDAC_N.n1440 VSS 0.132739f
C16718 VDAC_N.t2057 VSS 0.105768f
C16719 VDAC_N.n1441 VSS 0.132739f
C16720 VDAC_N.t707 VSS 0.105768f
C16721 VDAC_N.n1442 VSS 0.132739f
C16722 VDAC_N.t1849 VSS 0.105768f
C16723 VDAC_N.n1443 VSS 0.132739f
C16724 VDAC_N.t1124 VSS 0.105768f
C16725 VDAC_N.n1444 VSS 0.132739f
C16726 VDAC_N.t1737 VSS 0.105768f
C16727 VDAC_N.n1445 VSS 0.132739f
C16728 VDAC_N.t2076 VSS 0.105768f
C16729 VDAC_N.n1446 VSS 0.132739f
C16730 VDAC_N.t2016 VSS 0.105768f
C16731 VDAC_N.n1447 VSS 0.132739f
C16732 VDAC_N.t1059 VSS 0.105768f
C16733 VDAC_N.n1448 VSS 0.132739f
C16734 VDAC_N.t416 VSS 0.105768f
C16735 VDAC_N.n1449 VSS 0.132739f
C16736 VDAC_N.t953 VSS 0.105768f
C16737 VDAC_N.n1450 VSS 0.132739f
C16738 VDAC_N.t168 VSS 0.105768f
C16739 VDAC_N.n1451 VSS 0.132739f
C16740 VDAC_N.t774 VSS 0.105768f
C16741 VDAC_N.n1452 VSS 0.132739f
C16742 VDAC_N.t1822 VSS 0.105768f
C16743 VDAC_N.n1453 VSS 0.132739f
C16744 VDAC_N.t1391 VSS 0.105768f
C16745 VDAC_N.n1454 VSS 0.132739f
C16746 VDAC_N.t43 VSS 0.105768f
C16747 VDAC_N.n1455 VSS 0.132739f
C16748 VDAC_N.t1277 VSS 0.105768f
C16749 VDAC_N.n1456 VSS 0.132739f
C16750 VDAC_N.t885 VSS 0.105768f
C16751 VDAC_N.n1457 VSS 0.132739f
C16752 VDAC_N.t100 VSS 0.105768f
C16753 VDAC_N.n1458 VSS 0.132739f
C16754 VDAC_N.t1635 VSS 0.105768f
C16755 VDAC_N.n1459 VSS 0.132739f
C16756 VDAC_N.t1061 VSS 0.105768f
C16757 VDAC_N.n1460 VSS 0.132739f
C16758 VDAC_N.t1525 VSS 0.105768f
C16759 VDAC_N.n1461 VSS 0.132739f
C16760 VDAC_N.t1983 VSS 0.105768f
C16761 VDAC_N.n1462 VSS 0.132739f
C16762 VDAC_N.t1176 VSS 0.105768f
C16763 VDAC_N.n1463 VSS 0.132739f
C16764 VDAC_N.t897 VSS 0.105768f
C16765 VDAC_N.n1464 VSS 0.132739f
C16766 VDAC_N.t116 VSS 0.105768f
C16767 VDAC_N.n1465 VSS 0.132739f
C16768 VDAC_N.t346 VSS 0.105768f
C16769 VDAC_N.n1466 VSS 0.132739f
C16770 VDAC_N.t2123 VSS 0.105768f
C16771 VDAC_N.n1467 VSS 0.132739f
C16772 VDAC_N.t558 VSS 0.105768f
C16773 VDAC_N.n1468 VSS 0.132739f
C16774 VDAC_N.t2009 VSS 0.105768f
C16775 VDAC_N.n1469 VSS 0.132739f
C16776 VDAC_N.t656 VSS 0.105768f
C16777 VDAC_N.n1470 VSS 0.132739f
C16778 VDAC_N.t918 VSS 0.105768f
C16779 VDAC_N.n1471 VSS 0.132739f
C16780 VDAC_N.t1668 VSS 0.105768f
C16781 VDAC_N.n1472 VSS 0.132739f
C16782 VDAC_N.t1350 VSS 0.105768f
C16783 VDAC_N.n1473 VSS 0.132739f
C16784 VDAC_N.t595 VSS 0.105768f
C16785 VDAC_N.n1474 VSS 0.132739f
C16786 VDAC_N.t1146 VSS 0.105768f
C16787 VDAC_N.n1475 VSS 0.132739f
C16788 VDAC_N.t2078 VSS 0.105768f
C16789 VDAC_N.n1476 VSS 0.132739f
C16790 VDAC_N.t1384 VSS 0.105768f
C16791 VDAC_N.n1477 VSS 0.132739f
C16792 VDAC_N.t1858 VSS 0.105768f
C16793 VDAC_N.n1478 VSS 0.132739f
C16794 VDAC_N.t1411 VSS 0.105768f
C16795 VDAC_N.n1479 VSS 0.132739f
C16796 VDAC_N.t1602 VSS 0.105768f
C16797 VDAC_N.n1480 VSS 0.132739f
C16798 VDAC_N.t367 VSS 0.105768f
C16799 VDAC_N.n1481 VSS 0.132739f
C16800 VDAC_N.t1847 VSS 0.105768f
C16801 VDAC_N.n1482 VSS 0.132739f
C16802 VDAC_N.t1165 VSS 0.105768f
C16803 VDAC_N.n1483 VSS 0.132739f
C16804 VDAC_N.t1629 VSS 0.105768f
C16805 VDAC_N.n1484 VSS 0.132739f
C16806 VDAC_N.t2134 VSS 0.105768f
C16807 VDAC_N.n1485 VSS 0.132739f
C16808 VDAC_N.t1519 VSS 0.105768f
C16809 VDAC_N.n1486 VSS 0.132739f
C16810 VDAC_N.t1003 VSS 0.105768f
C16811 VDAC_N.n1487 VSS 0.132739f
C16812 VDAC_N.t1415 VSS 0.105768f
C16813 VDAC_N.n1488 VSS 0.132739f
C16814 VDAC_N.t1877 VSS 0.105768f
C16815 VDAC_N.n1489 VSS 0.132739f
C16816 VDAC_N.t708 VSS 0.105768f
C16817 VDAC_N.n1490 VSS 0.132739f
C16818 VDAC_N.t1763 VSS 0.105768f
C16819 VDAC_N.n1491 VSS 0.132739f
C16820 VDAC_N.t300 VSS 0.105768f
C16821 VDAC_N.n1492 VSS 0.132739f
C16822 VDAC_N.t2120 VSS 0.105768f
C16823 VDAC_N.n1493 VSS 0.132739f
C16824 VDAC_N.t2005 VSS 0.105768f
C16825 VDAC_N.n1494 VSS 0.132739f
C16826 VDAC_N.t872 VSS 0.105768f
C16827 VDAC_N.n1495 VSS 0.132739f
C16828 VDAC_N.t1901 VSS 0.105768f
C16829 VDAC_N.n1496 VSS 0.132739f
C16830 VDAC_N.t1636 VSS 0.105768f
C16831 VDAC_N.n1497 VSS 0.132739f
C16832 VDAC_N.t1586 VSS 0.105768f
C16833 VDAC_N.n1498 VSS 0.132739f
C16834 VDAC_N.t1484 VSS 0.105768f
C16835 VDAC_N.n1499 VSS 0.132739f
C16836 VDAC_N.t306 VSS 0.105768f
C16837 VDAC_N.n1500 VSS 0.132739f
C16838 VDAC_N.t593 VSS 0.105768f
C16839 VDAC_N.n1501 VSS 0.132739f
C16840 VDAC_N.t928 VSS 0.105768f
C16841 VDAC_N.n1502 VSS 0.12675f
C16842 VDAC_N.t710 VSS 0.105768f
C16843 VDAC_N.n1503 VSS 0.132739f
C16844 VDAC_N.t1283 VSS 0.105768f
C16845 VDAC_N.n1504 VSS 0.132739f
C16846 VDAC_N.t314 VSS 0.105768f
C16847 VDAC_N.n1505 VSS 0.132739f
C16848 VDAC_N.t1066 VSS 0.105768f
C16849 VDAC_N.n1506 VSS 0.132739f
C16850 VDAC_N.t1531 VSS 0.105768f
C16851 VDAC_N.n1507 VSS 0.132739f
C16852 VDAC_N.t1894 VSS 0.105768f
C16853 VDAC_N.n1508 VSS 0.132739f
C16854 VDAC_N.t1421 VSS 0.105768f
C16855 VDAC_N.n1509 VSS 0.132739f
C16856 VDAC_N.t1885 VSS 0.105768f
C16857 VDAC_N.n1510 VSS 0.132739f
C16858 VDAC_N.t189 VSS 0.105768f
C16859 VDAC_N.n1511 VSS 0.132739f
C16860 VDAC_N.t1773 VSS 0.105768f
C16861 VDAC_N.n1512 VSS 0.132739f
C16862 VDAC_N.t1091 VSS 0.105768f
C16863 VDAC_N.n1513 VSS 0.132739f
C16864 VDAC_N.t1667 VSS 0.105768f
C16865 VDAC_N.n1514 VSS 0.132739f
C16866 VDAC_N.t2127 VSS 0.105768f
C16867 VDAC_N.n1515 VSS 0.132739f
C16868 VDAC_N.t1422 VSS 0.105768f
C16869 VDAC_N.n1516 VSS 0.132739f
C16870 VDAC_N.t1195 VSS 0.105768f
C16871 VDAC_N.n1517 VSS 0.132739f
C16872 VDAC_N.t245 VSS 0.105768f
C16873 VDAC_N.n1518 VSS 0.132739f
C16874 VDAC_N.t23 VSS 0.105768f
C16875 VDAC_N.n1519 VSS 0.132739f
C16876 VDAC_N.t1549 VSS 0.105768f
C16877 VDAC_N.n1520 VSS 0.132739f
C16878 VDAC_N.t1073 VSS 0.105768f
C16879 VDAC_N.n1521 VSS 0.132739f
C16880 VDAC_N.t1443 VSS 0.105768f
C16881 VDAC_N.n1522 VSS 0.132739f
C16882 VDAC_N.t965 VSS 0.105768f
C16883 VDAC_N.n1523 VSS 0.132739f
C16884 VDAC_N.t1339 VSS 0.105768f
C16885 VDAC_N.n1524 VSS 0.132739f
C16886 VDAC_N.t1795 VSS 0.105768f
C16887 VDAC_N.n1525 VSS 0.132739f
C16888 VDAC_N.t396 VSS 0.105768f
C16889 VDAC_N.n1526 VSS 0.132739f
C16890 VDAC_N.t1579 VSS 0.105768f
C16891 VDAC_N.n1527 VSS 0.132739f
C16892 VDAC_N.t1074 VSS 0.105768f
C16893 VDAC_N.n1528 VSS 0.132739f
C16894 VDAC_N.t1832 VSS 0.105768f
C16895 VDAC_N.n1529 VSS 0.132739f
C16896 VDAC_N.t503 VSS 0.105768f
C16897 VDAC_N.n1530 VSS 0.132739f
C16898 VDAC_N.t1376 VSS 0.105768f
C16899 VDAC_N.n1531 VSS 0.132739f
C16900 VDAC_N.t1825 VSS 0.105768f
C16901 VDAC_N.n1532 VSS 0.132739f
C16902 VDAC_N.t972 VSS 0.105768f
C16903 VDAC_N.n1533 VSS 0.132739f
C16904 VDAC_N.t1410 VSS 0.105768f
C16905 VDAC_N.n1534 VSS 0.132739f
C16906 VDAC_N.t476 VSS 0.105768f
C16907 VDAC_N.n1535 VSS 0.132739f
C16908 VDAC_N.t504 VSS 0.105768f
C16909 VDAC_N.n1536 VSS 0.132739f
C16910 VDAC_N.t502 VSS 0.105768f
C16911 VDAC_N.n1537 VSS 0.132739f
C16912 VDAC_N.t392 VSS 0.105768f
C16913 VDAC_N.n1538 VSS 0.132739f
C16914 VDAC_N.t54 VSS 0.105768f
C16915 VDAC_N.n1539 VSS 0.132739f
C16916 VDAC_N.t1220 VSS 0.105768f
C16917 VDAC_N.n1540 VSS 0.132739f
C16918 VDAC_N.t118 VSS 0.105768f
C16919 VDAC_N.n1541 VSS 0.132739f
C16920 VDAC_N.t623 VSS 0.105768f
C16921 VDAC_N.n1542 VSS 0.132739f
C16922 VDAC_N.t618 VSS 0.105768f
C16923 VDAC_N.n1543 VSS 0.132739f
C16924 VDAC_N.t1189 VSS 0.105768f
C16925 VDAC_N.n1544 VSS 0.132739f
C16926 VDAC_N.t435 VSS 0.105768f
C16927 VDAC_N.n1545 VSS 0.132739f
C16928 VDAC_N.t266 VSS 0.105768f
C16929 VDAC_N.n1546 VSS 0.132739f
C16930 VDAC_N.t1439 VSS 0.105768f
C16931 VDAC_N.n1547 VSS 0.132739f
C16932 VDAC_N.t1999 VSS 0.105768f
C16933 VDAC_N.n1548 VSS 0.132739f
C16934 VDAC_N.t191 VSS 0.105768f
C16935 VDAC_N.n1549 VSS 0.132739f
C16936 VDAC_N.t909 VSS 0.105768f
C16937 VDAC_N.n1550 VSS 0.132739f
C16938 VDAC_N.t1223 VSS 0.105768f
C16939 VDAC_N.n1551 VSS 0.132739f
C16940 VDAC_N.t443 VSS 0.105768f
C16941 VDAC_N.n1552 VSS 0.132739f
C16942 VDAC_N.t970 VSS 0.105768f
C16943 VDAC_N.n1553 VSS 0.132739f
C16944 VDAC_N.t1573 VSS 0.105768f
C16945 VDAC_N.n1554 VSS 0.132739f
C16946 VDAC_N.t2037 VSS 0.105768f
C16947 VDAC_N.n1555 VSS 0.132739f
C16948 VDAC_N.t688 VSS 0.105768f
C16949 VDAC_N.n1556 VSS 0.132739f
C16950 VDAC_N.t35 VSS 0.105768f
C16951 VDAC_N.n1557 VSS 0.132739f
C16952 VDAC_N.t932 VSS 0.105768f
C16953 VDAC_N.n1558 VSS 0.132739f
C16954 VDAC_N.t869 VSS 0.105768f
C16955 VDAC_N.n1559 VSS 0.132739f
C16956 VDAC_N.t12 VSS 0.105768f
C16957 VDAC_N.n1560 VSS 0.132739f
C16958 VDAC_N.t606 VSS 0.105768f
C16959 VDAC_N.n1561 VSS 0.132739f
C16960 VDAC_N.t2063 VSS 0.105768f
C16961 VDAC_N.n1562 VSS 0.132739f
C16962 VDAC_N.t208 VSS 0.105768f
C16963 VDAC_N.n1563 VSS 0.132739f
C16964 VDAC_N.t1910 VSS 0.105768f
C16965 VDAC_N.n1564 VSS 0.132739f
C16966 VDAC_N.t1060 VSS 0.105768f
C16967 VDAC_N.n1565 VSS 0.12675f
C16968 VDAC_N.t1831 VSS 0.105768f
C16969 VDAC_N.n1566 VSS 0.132739f
C16970 VDAC_N.t964 VSS 0.105768f
C16971 VDAC_N.n1567 VSS 0.132739f
C16972 VDAC_N.t875 VSS 0.105768f
C16973 VDAC_N.n1568 VSS 0.132739f
C16974 VDAC_N.t540 VSS 0.105768f
C16975 VDAC_N.n1569 VSS 0.132739f
C16976 VDAC_N.t992 VSS 0.105768f
C16977 VDAC_N.n1570 VSS 0.132739f
C16978 VDAC_N.t2075 VSS 0.105768f
C16979 VDAC_N.n1571 VSS 0.132739f
C16980 VDAC_N.t768 VSS 0.105768f
C16981 VDAC_N.n1572 VSS 0.132739f
C16982 VDAC_N.t1706 VSS 0.105768f
C16983 VDAC_N.n1573 VSS 0.132739f
C16984 VDAC_N.t1088 VSS 0.105768f
C16985 VDAC_N.n1574 VSS 0.132739f
C16986 VDAC_N.t754 VSS 0.105768f
C16987 VDAC_N.n1575 VSS 0.132739f
C16988 VDAC_N.t1724 VSS 0.105768f
C16989 VDAC_N.n1576 VSS 0.132739f
C16990 VDAC_N.t1262 VSS 0.105768f
C16991 VDAC_N.n1577 VSS 0.132739f
C16992 VDAC_N.t1109 VSS 0.105768f
C16993 VDAC_N.n1578 VSS 0.132739f
C16994 VDAC_N.t385 VSS 0.105768f
C16995 VDAC_N.n1579 VSS 0.132739f
C16996 VDAC_N.t1915 VSS 0.105768f
C16997 VDAC_N.n1580 VSS 0.132739f
C16998 VDAC_N.t1312 VSS 0.105768f
C16999 VDAC_N.n1581 VSS 0.132739f
C17000 VDAC_N.t473 VSS 0.105768f
C17001 VDAC_N.n1582 VSS 0.132739f
C17002 VDAC_N.t236 VSS 0.105768f
C17003 VDAC_N.n1583 VSS 0.132739f
C17004 VDAC_N.t698 VSS 0.105768f
C17005 VDAC_N.n1584 VSS 0.132739f
C17006 VDAC_N.t1948 VSS 0.105768f
C17007 VDAC_N.n1585 VSS 0.132739f
C17008 VDAC_N.t1880 VSS 0.105768f
C17009 VDAC_N.n1586 VSS 0.132739f
C17010 VDAC_N.t281 VSS 0.105768f
C17011 VDAC_N.n1587 VSS 0.132739f
C17012 VDAC_N.t728 VSS 0.105768f
C17013 VDAC_N.n1588 VSS 0.132739f
C17014 VDAC_N.t1658 VSS 0.105768f
C17015 VDAC_N.n1589 VSS 0.132739f
C17016 VDAC_N.t1068 VSS 0.105768f
C17017 VDAC_N.n1590 VSS 0.132739f
C17018 VDAC_N.t1430 VSS 0.105768f
C17019 VDAC_N.n1591 VSS 0.132739f
C17020 VDAC_N.t321 VSS 0.105768f
C17021 VDAC_N.n1592 VSS 0.132739f
C17022 VDAC_N.t2000 VSS 0.105768f
C17023 VDAC_N.n1593 VSS 0.132739f
C17024 VDAC_N.t61 VSS 0.105768f
C17025 VDAC_N.n1594 VSS 0.132739f
C17026 VDAC_N.t408 VSS 0.105768f
C17027 VDAC_N.n1595 VSS 0.132739f
C17028 VDAC_N.t1722 VSS 0.105768f
C17029 VDAC_N.n1596 VSS 0.132739f
C17030 VDAC_N.t383 VSS 0.105768f
C17031 VDAC_N.n1597 VSS 0.132739f
C17032 VDAC_N.t1502 VSS 0.105768f
C17033 VDAC_N.n1598 VSS 0.132739f
C17034 VDAC_N.t1229 VSS 0.105768f
C17035 VDAC_N.n1599 VSS 0.132739f
C17036 VDAC_N.t1697 VSS 0.105768f
C17037 VDAC_N.n1600 VSS 0.132739f
C17038 VDAC_N.t1117 VSS 0.105768f
C17039 VDAC_N.n1601 VSS 0.132739f
C17040 VDAC_N.t1583 VSS 0.105768f
C17041 VDAC_N.n1602 VSS 0.132739f
C17042 VDAC_N.t902 VSS 0.105768f
C17043 VDAC_N.n1603 VSS 0.132739f
C17044 VDAC_N.t1471 VSS 0.105768f
C17045 VDAC_N.n1604 VSS 0.132739f
C17046 VDAC_N.t1931 VSS 0.105768f
C17047 VDAC_N.n1605 VSS 0.132739f
C17048 VDAC_N.t1347 VSS 0.105768f
C17049 VDAC_N.n1606 VSS 0.132739f
C17050 VDAC_N.t967 VSS 0.105768f
C17051 VDAC_N.n1607 VSS 0.132739f
C17052 VDAC_N.t1700 VSS 0.105768f
C17053 VDAC_N.n1608 VSS 0.132739f
C17054 VDAC_N.t237 VSS 0.105768f
C17055 VDAC_N.n1609 VSS 0.132739f
C17056 VDAC_N.t1372 VSS 0.105768f
C17057 VDAC_N.n1610 VSS 0.132739f
C17058 VDAC_N.t590 VSS 0.105768f
C17059 VDAC_N.n1611 VSS 0.132739f
C17060 VDAC_N.t1037 VSS 0.105768f
C17061 VDAC_N.n1612 VSS 0.132739f
C17062 VDAC_N.t200 VSS 0.105768f
C17063 VDAC_N.n1613 VSS 0.132739f
C17064 VDAC_N.t1935 VSS 0.105768f
C17065 VDAC_N.n1614 VSS 0.132739f
C17066 VDAC_N.t1924 VSS 0.105768f
C17067 VDAC_N.n1615 VSS 0.132739f
C17068 VDAC_N.t722 VSS 0.105768f
C17069 VDAC_N.n1616 VSS 0.132739f
C17070 VDAC_N.t524 VSS 0.105768f
C17071 VDAC_N.n1617 VSS 0.132739f
C17072 VDAC_N.t622 VSS 0.105768f
C17073 VDAC_N.n1618 VSS 0.132739f
C17074 VDAC_N.t19 VSS 0.105768f
C17075 VDAC_N.n1619 VSS 0.132739f
C17076 VDAC_N.t1528 VSS 0.105768f
C17077 VDAC_N.n1620 VSS 0.132739f
C17078 VDAC_N.t1942 VSS 0.105768f
C17079 VDAC_N.n1621 VSS 0.132739f
C17080 VDAC_N.t1104 VSS 0.105768f
C17081 VDAC_N.n1622 VSS 0.132739f
C17082 VDAC_N.t1490 VSS 0.105768f
C17083 VDAC_N.n1623 VSS 0.132739f
C17084 VDAC_N.t1337 VSS 0.105768f
C17085 VDAC_N.n1624 VSS 0.132739f
C17086 VDAC_N.t650 VSS 0.105768f
C17087 VDAC_N.n1625 VSS 0.132739f
C17088 VDAC_N.t299 VSS 0.105768f
C17089 VDAC_N.n1626 VSS 0.132739f
C17090 VDAC_N.t41 VSS 0.105768f
C17091 VDAC_N.n1627 VSS 0.132739f
C17092 VDAC_N.t1014 VSS 0.105768f
C17093 VDAC_N.n1628 VSS 0.12675f
C17094 VDAC_N.t1054 VSS 0.105768f
C17095 VDAC_N.n1629 VSS 0.132739f
C17096 VDAC_N.t427 VSS 0.105768f
C17097 VDAC_N.n1630 VSS 0.132739f
C17098 VDAC_N.t486 VSS 0.105768f
C17099 VDAC_N.n1631 VSS 0.132739f
C17100 VDAC_N.t201 VSS 0.105768f
C17101 VDAC_N.n1632 VSS 0.132739f
C17102 VDAC_N.t1873 VSS 0.105768f
C17103 VDAC_N.n1633 VSS 0.132739f
C17104 VDAC_N.t665 VSS 0.105768f
C17105 VDAC_N.n1634 VSS 0.132739f
C17106 VDAC_N.t1759 VSS 0.105768f
C17107 VDAC_N.n1635 VSS 0.132739f
C17108 VDAC_N.t60 VSS 0.105768f
C17109 VDAC_N.n1636 VSS 0.132739f
C17110 VDAC_N.t1657 VSS 0.105768f
C17111 VDAC_N.n1637 VSS 0.132739f
C17112 VDAC_N.t2113 VSS 0.105768f
C17113 VDAC_N.n1638 VSS 0.132739f
C17114 VDAC_N.t381 VSS 0.105768f
C17115 VDAC_N.n1639 VSS 0.132739f
C17116 VDAC_N.t521 VSS 0.105768f
C17117 VDAC_N.n1640 VSS 0.132739f
C17118 VDAC_N.t1256 VSS 0.105768f
C17119 VDAC_N.n1641 VSS 0.132739f
C17120 VDAC_N.t1263 VSS 0.105768f
C17121 VDAC_N.n1642 VSS 0.132739f
C17122 VDAC_N.t1725 VSS 0.105768f
C17123 VDAC_N.n1643 VSS 0.132739f
C17124 VDAC_N.t2028 VSS 0.105768f
C17125 VDAC_N.n1644 VSS 0.132739f
C17126 VDAC_N.t1617 VSS 0.105768f
C17127 VDAC_N.n1645 VSS 0.132739f
C17128 VDAC_N.t1053 VSS 0.105768f
C17129 VDAC_N.n1646 VSS 0.132739f
C17130 VDAC_N.t1000 VSS 0.105768f
C17131 VDAC_N.n1647 VSS 0.132739f
C17132 VDAC_N.t1965 VSS 0.105768f
C17133 VDAC_N.n1648 VSS 0.132739f
C17134 VDAC_N.t568 VSS 0.105768f
C17135 VDAC_N.n1649 VSS 0.132739f
C17136 VDAC_N.t947 VSS 0.105768f
C17137 VDAC_N.n1650 VSS 0.132739f
C17138 VDAC_N.t68 VSS 0.105768f
C17139 VDAC_N.n1651 VSS 0.132739f
C17140 VDAC_N.t1274 VSS 0.105768f
C17141 VDAC_N.n1652 VSS 0.132739f
C17142 VDAC_N.t1067 VSS 0.105768f
C17143 VDAC_N.n1653 VSS 0.132739f
C17144 VDAC_N.t1056 VSS 0.105768f
C17145 VDAC_N.n1654 VSS 0.132739f
C17146 VDAC_N.t2002 VSS 0.105768f
C17147 VDAC_N.n1655 VSS 0.132739f
C17148 VDAC_N.t632 VSS 0.105768f
C17149 VDAC_N.n1656 VSS 0.132739f
C17150 VDAC_N.t898 VSS 0.105768f
C17151 VDAC_N.n1657 VSS 0.132739f
C17152 VDAC_N.t1540 VSS 0.105768f
C17153 VDAC_N.n1658 VSS 0.132739f
C17154 VDAC_N.t678 VSS 0.105768f
C17155 VDAC_N.n1659 VSS 0.132739f
C17156 VDAC_N.t1255 VSS 0.105768f
C17157 VDAC_N.n1660 VSS 0.132739f
C17158 VDAC_N.t1118 VSS 0.105768f
C17159 VDAC_N.n1661 VSS 0.132739f
C17160 VDAC_N.t1038 VSS 0.105768f
C17161 VDAC_N.n1662 VSS 0.132739f
C17162 VDAC_N.t1499 VSS 0.105768f
C17163 VDAC_N.n1663 VSS 0.132739f
C17164 VDAC_N.t478 VSS 0.105768f
C17165 VDAC_N.n1664 VSS 0.132739f
C17166 VDAC_N.t199 VSS 0.105768f
C17167 VDAC_N.n1665 VSS 0.132739f
C17168 VDAC_N.t1386 VSS 0.105768f
C17169 VDAC_N.n1666 VSS 0.132739f
C17170 VDAC_N.t655 VSS 0.105768f
C17171 VDAC_N.n1667 VSS 0.132739f
C17172 VDAC_N.t243 VSS 0.105768f
C17173 VDAC_N.n1668 VSS 0.132739f
C17174 VDAC_N.t309 VSS 0.105768f
C17175 VDAC_N.n1669 VSS 0.132739f
C17176 VDAC_N.t873 VSS 0.105768f
C17177 VDAC_N.n1670 VSS 0.132739f
C17178 VDAC_N.t1884 VSS 0.105768f
C17179 VDAC_N.n1671 VSS 0.132739f
C17180 VDAC_N.t1505 VSS 0.105768f
C17181 VDAC_N.n1672 VSS 0.132739f
C17182 VDAC_N.t1957 VSS 0.105768f
C17183 VDAC_N.n1673 VSS 0.132739f
C17184 VDAC_N.t120 VSS 0.105768f
C17185 VDAC_N.n1674 VSS 0.132739f
C17186 VDAC_N.t1859 VSS 0.105768f
C17187 VDAC_N.n1675 VSS 0.132739f
C17188 VDAC_N.t644 VSS 0.105768f
C17189 VDAC_N.n1676 VSS 0.132739f
C17190 VDAC_N.t1753 VSS 0.105768f
C17191 VDAC_N.n1677 VSS 0.132739f
C17192 VDAC_N.t828 VSS 0.105768f
C17193 VDAC_N.n1678 VSS 0.132739f
C17194 VDAC_N.t2064 VSS 0.105768f
C17195 VDAC_N.n1679 VSS 0.132739f
C17196 VDAC_N.t2099 VSS 0.105768f
C17197 VDAC_N.n1680 VSS 0.132739f
C17198 VDAC_N.t1656 VSS 0.105768f
C17199 VDAC_N.n1681 VSS 0.132739f
C17200 VDAC_N.t890 VSS 0.105768f
C17201 VDAC_N.n1682 VSS 0.132739f
C17202 VDAC_N.t1492 VSS 0.105768f
C17203 VDAC_N.n1683 VSS 0.132739f
C17204 VDAC_N.t218 VSS 0.105768f
C17205 VDAC_N.n1684 VSS 0.132739f
C17206 VDAC_N.t1260 VSS 0.105768f
C17207 VDAC_N.n1685 VSS 0.132739f
C17208 VDAC_N.t298 VSS 0.105768f
C17209 VDAC_N.n1686 VSS 0.132739f
C17210 VDAC_N.t1139 VSS 0.105768f
C17211 VDAC_N.n1687 VSS 0.132739f
C17212 VDAC_N.t896 VSS 0.105768f
C17213 VDAC_N.n1688 VSS 0.132739f
C17214 VDAC_N.t42 VSS 0.105768f
C17215 VDAC_N.n1689 VSS 0.132739f
C17216 VDAC_N.t761 VSS 0.105768f
C17217 VDAC_N.n1690 VSS 0.132739f
C17218 VDAC_N.t226 VSS 0.105768f
C17219 VDAC_N.n1691 VSS 0.12675f
C17220 VDAC_N.t20 VSS 0.105768f
C17221 VDAC_N.n1692 VSS 0.132739f
C17222 VDAC_N.t602 VSS 0.105768f
C17223 VDAC_N.n1693 VSS 0.132739f
C17224 VDAC_N.t2059 VSS 0.105768f
C17225 VDAC_N.n1694 VSS 0.132739f
C17226 VDAC_N.t1456 VSS 0.105768f
C17227 VDAC_N.n1695 VSS 0.132739f
C17228 VDAC_N.t1678 VSS 0.105768f
C17229 VDAC_N.n1696 VSS 0.132739f
C17230 VDAC_N.t1044 VSS 0.105768f
C17231 VDAC_N.n1697 VSS 0.132739f
C17232 VDAC_N.t738 VSS 0.105768f
C17233 VDAC_N.n1698 VSS 0.132739f
C17234 VDAC_N.t1211 VSS 0.105768f
C17235 VDAC_N.n1699 VSS 0.132739f
C17236 VDAC_N.t330 VSS 0.105768f
C17237 VDAC_N.n1700 VSS 0.132739f
C17238 VDAC_N.t561 VSS 0.105768f
C17239 VDAC_N.n1701 VSS 0.132739f
C17240 VDAC_N.t224 VSS 0.105768f
C17241 VDAC_N.n1702 VSS 0.132739f
C17242 VDAC_N.t1958 VSS 0.105768f
C17243 VDAC_N.n1703 VSS 0.132739f
C17244 VDAC_N.t741 VSS 0.105768f
C17245 VDAC_N.n1704 VSS 0.132739f
C17246 VDAC_N.t1981 VSS 0.105768f
C17247 VDAC_N.n1705 VSS 0.132739f
C17248 VDAC_N.t312 VSS 0.105768f
C17249 VDAC_N.n1706 VSS 0.132739f
C17250 VDAC_N.t882 VSS 0.105768f
C17251 VDAC_N.n1707 VSS 0.132739f
C17252 VDAC_N.t724 VSS 0.105768f
C17253 VDAC_N.n1708 VSS 0.132739f
C17254 VDAC_N.t1294 VSS 0.105768f
C17255 VDAC_N.n1709 VSS 0.132739f
C17256 VDAC_N.t179 VSS 0.105768f
C17257 VDAC_N.n1710 VSS 0.132739f
C17258 VDAC_N.t94 VSS 0.105768f
C17259 VDAC_N.n1711 VSS 0.132739f
C17260 VDAC_N.t526 VSS 0.105768f
C17261 VDAC_N.n1712 VSS 0.132739f
C17262 VDAC_N.t240 VSS 0.105768f
C17263 VDAC_N.n1713 VSS 0.132739f
C17264 VDAC_N.t1802 VSS 0.105768f
C17265 VDAC_N.n1714 VSS 0.132739f
C17266 VDAC_N.t197 VSS 0.105768f
C17267 VDAC_N.n1715 VSS 0.132739f
C17268 VDAC_N.t358 VSS 0.105768f
C17269 VDAC_N.n1716 VSS 0.132739f
C17270 VDAC_N.t647 VSS 0.105768f
C17271 VDAC_N.n1717 VSS 0.132739f
C17272 VDAC_N.t1729 VSS 0.105768f
C17273 VDAC_N.n1718 VSS 0.132739f
C17274 VDAC_N.t2074 VSS 0.105768f
C17275 VDAC_N.n1719 VSS 0.132739f
C17276 VDAC_N.t1621 VSS 0.105768f
C17277 VDAC_N.n1720 VSS 0.132739f
C17278 VDAC_N.t942 VSS 0.105768f
C17279 VDAC_N.n1721 VSS 0.132739f
C17280 VDAC_N.t719 VSS 0.105768f
C17281 VDAC_N.n1722 VSS 0.132739f
C17282 VDAC_N.t999 VSS 0.105768f
C17283 VDAC_N.n1723 VSS 0.132739f
C17284 VDAC_N.t1299 VSS 0.105768f
C17285 VDAC_N.n1724 VSS 0.132739f
C17286 VDAC_N.t893 VSS 0.105768f
C17287 VDAC_N.n1725 VSS 0.132739f
C17288 VDAC_N.t1916 VSS 0.105768f
C17289 VDAC_N.n1726 VSS 0.132739f
C17290 VDAC_N.t1655 VSS 0.105768f
C17291 VDAC_N.n1727 VSS 0.132739f
C17292 VDAC_N.t2109 VSS 0.105768f
C17293 VDAC_N.n1728 VSS 0.132739f
C17294 VDAC_N.t731 VSS 0.105768f
C17295 VDAC_N.n1729 VSS 0.132739f
C17296 VDAC_N.t1013 VSS 0.105768f
C17297 VDAC_N.n1730 VSS 0.132739f
C17298 VDAC_N.t104 VSS 0.105768f
C17299 VDAC_N.n1731 VSS 0.132739f
C17300 VDAC_N.t1875 VSS 0.105768f
C17301 VDAC_N.n1732 VSS 0.132739f
C17302 VDAC_N.t1128 VSS 0.105768f
C17303 VDAC_N.n1733 VSS 0.132739f
C17304 VDAC_N.t1510 VSS 0.105768f
C17305 VDAC_N.n1734 VSS 0.132739f
C17306 VDAC_N.t556 VSS 0.105768f
C17307 VDAC_N.n1735 VSS 0.132739f
C17308 VDAC_N.t2112 VSS 0.105768f
C17309 VDAC_N.n1736 VSS 0.132739f
C17310 VDAC_N.t1121 VSS 0.105768f
C17311 VDAC_N.n1737 VSS 0.132739f
C17312 VDAC_N.t1704 VSS 0.105768f
C17313 VDAC_N.n1738 VSS 0.132739f
C17314 VDAC_N.t1790 VSS 0.105768f
C17315 VDAC_N.n1739 VSS 0.132739f
C17316 VDAC_N.t336 VSS 0.105768f
C17317 VDAC_N.n1740 VSS 0.132739f
C17318 VDAC_N.t222 VSS 0.105768f
C17319 VDAC_N.n1741 VSS 0.132739f
C17320 VDAC_N.t1261 VSS 0.105768f
C17321 VDAC_N.n1742 VSS 0.132739f
C17322 VDAC_N.t1338 VSS 0.105768f
C17323 VDAC_N.n1743 VSS 0.132739f
C17324 VDAC_N.t169 VSS 0.105768f
C17325 VDAC_N.n1744 VSS 0.132739f
C17326 VDAC_N.t821 VSS 0.105768f
C17327 VDAC_N.n1745 VSS 0.132739f
C17328 VDAC_N.t938 VSS 0.105768f
C17329 VDAC_N.n1746 VSS 0.132739f
C17330 VDAC_N.t769 VSS 0.105768f
C17331 VDAC_N.n1747 VSS 0.132739f
C17332 VDAC_N.t830 VSS 0.105768f
C17333 VDAC_N.n1748 VSS 0.132739f
C17334 VDAC_N.t661 VSS 0.105768f
C17335 VDAC_N.n1749 VSS 0.132739f
C17336 VDAC_N.t1863 VSS 0.105768f
C17337 VDAC_N.n1750 VSS 0.132739f
C17338 VDAC_N.t1183 VSS 0.105768f
C17339 VDAC_N.n1751 VSS 0.132739f
C17340 VDAC_N.t1651 VSS 0.105768f
C17341 VDAC_N.n1752 VSS 0.132739f
C17342 VDAC_N.t444 VSS 0.105768f
C17343 VDAC_N.n1753 VSS 0.132739f
C17344 VDAC_N.t217 VSS 0.105768f
C17345 VDAC_N.n1754 VSS 0.12675f
C17346 VDAC_N.t1399 VSS 0.105768f
C17347 VDAC_N.n1755 VSS 0.132739f
C17348 VDAC_N.t991 VSS 0.105768f
C17349 VDAC_N.n1756 VSS 0.132739f
C17350 VDAC_N.t657 VSS 0.105768f
C17351 VDAC_N.n1757 VSS 0.132739f
C17352 VDAC_N.t889 VSS 0.105768f
C17353 VDAC_N.n1758 VSS 0.132739f
C17354 VDAC_N.t764 VSS 0.105768f
C17355 VDAC_N.n1759 VSS 0.132739f
C17356 VDAC_N.t1645 VSS 0.105768f
C17357 VDAC_N.n1760 VSS 0.132739f
C17358 VDAC_N.t2097 VSS 0.105768f
C17359 VDAC_N.n1761 VSS 0.132739f
C17360 VDAC_N.t1640 VSS 0.105768f
C17361 VDAC_N.n1762 VSS 0.132739f
C17362 VDAC_N.t1009 VSS 0.105768f
C17363 VDAC_N.n1763 VSS 0.132739f
C17364 VDAC_N.t1200 VSS 0.105768f
C17365 VDAC_N.n1764 VSS 0.132739f
C17366 VDAC_N.t1777 VSS 0.105768f
C17367 VDAC_N.n1765 VSS 0.132739f
C17368 VDAC_N.t740 VSS 0.105768f
C17369 VDAC_N.n1766 VSS 0.132739f
C17370 VDAC_N.t670 VSS 0.105768f
C17371 VDAC_N.n1767 VSS 0.132739f
C17372 VDAC_N.t1793 VSS 0.105768f
C17373 VDAC_N.n1768 VSS 0.132739f
C17374 VDAC_N.t748 VSS 0.105768f
C17375 VDAC_N.n1769 VSS 0.132739f
C17376 VDAC_N.t110 VSS 0.105768f
C17377 VDAC_N.n1770 VSS 0.132739f
C17378 VDAC_N.t2114 VSS 0.105768f
C17379 VDAC_N.n1771 VSS 0.132739f
C17380 VDAC_N.t1824 VSS 0.105768f
C17381 VDAC_N.n1772 VSS 0.132739f
C17382 VDAC_N.t2062 VSS 0.105768f
C17383 VDAC_N.n1773 VSS 0.132739f
C17384 VDAC_N.t696 VSS 0.105768f
C17385 VDAC_N.n1774 VSS 0.132739f
C17386 VDAC_N.t1634 VSS 0.105768f
C17387 VDAC_N.n1775 VSS 0.132739f
C17388 VDAC_N.t1860 VSS 0.105768f
C17389 VDAC_N.n1776 VSS 0.132739f
C17390 VDAC_N.t1406 VSS 0.105768f
C17391 VDAC_N.n1777 VSS 0.132739f
C17392 VDAC_N.t317 VSS 0.105768f
C17393 VDAC_N.n1778 VSS 0.132739f
C17394 VDAC_N.t976 VSS 0.105768f
C17395 VDAC_N.n1779 VSS 0.132739f
C17396 VDAC_N.t11 VSS 0.105768f
C17397 VDAC_N.n1780 VSS 0.132739f
C17398 VDAC_N.t1541 VSS 0.105768f
C17399 VDAC_N.n1781 VSS 0.132739f
C17400 VDAC_N.t858 VSS 0.105768f
C17401 VDAC_N.n1782 VSS 0.132739f
C17402 VDAC_N.t1431 VSS 0.105768f
C17403 VDAC_N.n1783 VSS 0.132739f
C17404 VDAC_N.t1462 VSS 0.105768f
C17405 VDAC_N.n1784 VSS 0.132739f
C17406 VDAC_N.t325 VSS 0.105768f
C17407 VDAC_N.n1785 VSS 0.132739f
C17408 VDAC_N.t467 VSS 0.105768f
C17409 VDAC_N.n1786 VSS 0.132739f
C17410 VDAC_N.t1101 VSS 0.105768f
C17411 VDAC_N.n1787 VSS 0.132739f
C17412 VDAC_N.t1567 VSS 0.105768f
C17413 VDAC_N.n1788 VSS 0.132739f
C17414 VDAC_N.t2027 VSS 0.105768f
C17415 VDAC_N.n1789 VSS 0.132739f
C17416 VDAC_N.t207 VSS 0.105768f
C17417 VDAC_N.n1790 VSS 0.132739f
C17418 VDAC_N.t1919 VSS 0.105768f
C17419 VDAC_N.n1791 VSS 0.132739f
C17420 VDAC_N.t1241 VSS 0.105768f
C17421 VDAC_N.n1792 VSS 0.132739f
C17422 VDAC_N.t1813 VSS 0.105768f
C17423 VDAC_N.n1793 VSS 0.132739f
C17424 VDAC_N.t460 VSS 0.105768f
C17425 VDAC_N.n1794 VSS 0.132739f
C17426 VDAC_N.t235 VSS 0.105768f
C17427 VDAC_N.n1795 VSS 0.132739f
C17428 VDAC_N.t1356 VSS 0.105768f
C17429 VDAC_N.n1796 VSS 0.132739f
C17430 VDAC_N.t1126 VSS 0.105768f
C17431 VDAC_N.n1797 VSS 0.132739f
C17432 VDAC_N.t529 VSS 0.105768f
C17433 VDAC_N.n1798 VSS 0.132739f
C17434 VDAC_N.t1344 VSS 0.105768f
C17435 VDAC_N.n1799 VSS 0.132739f
C17436 VDAC_N.t254 VSS 0.105768f
C17437 VDAC_N.n1800 VSS 0.132739f
C17438 VDAC_N.t1812 VSS 0.105768f
C17439 VDAC_N.n1801 VSS 0.132739f
C17440 VDAC_N.t370 VSS 0.105768f
C17441 VDAC_N.n1802 VSS 0.132739f
C17442 VDAC_N.t1804 VSS 0.105768f
C17443 VDAC_N.n1803 VSS 0.132739f
C17444 VDAC_N.t46 VSS 0.105768f
C17445 VDAC_N.n1804 VSS 0.132739f
C17446 VDAC_N.t8 VSS 0.105768f
C17447 VDAC_N.n1805 VSS 0.132739f
C17448 VDAC_N.t496 VSS 0.105768f
C17449 VDAC_N.n1806 VSS 0.132739f
C17450 VDAC_N.t966 VSS 0.105768f
C17451 VDAC_N.n1807 VSS 0.132739f
C17452 VDAC_N.t377 VSS 0.105768f
C17453 VDAC_N.n1808 VSS 0.132739f
C17454 VDAC_N.t206 VSS 0.105768f
C17455 VDAC_N.n1809 VSS 0.132739f
C17456 VDAC_N.t675 VSS 0.105768f
C17457 VDAC_N.n1810 VSS 0.132739f
C17458 VDAC_N.t634 VSS 0.105768f
C17459 VDAC_N.n1811 VSS 0.132739f
C17460 VDAC_N.t1095 VSS 0.105768f
C17461 VDAC_N.n1812 VSS 0.132739f
C17462 VDAC_N.t1673 VSS 0.105768f
C17463 VDAC_N.n1813 VSS 0.132739f
C17464 VDAC_N.t1962 VSS 0.105768f
C17465 VDAC_N.n1814 VSS 0.132739f
C17466 VDAC_N.t1455 VSS 0.105768f
C17467 VDAC_N.n1815 VSS 0.132739f
C17468 VDAC_N.t277 VSS 0.105768f
C17469 VDAC_N.n1816 VSS 0.132739f
C17470 VDAC_N.t1353 VSS 0.105768f
C17471 VDAC_N.n1817 VSS 0.12675f
C17472 VDAC_N.t1202 VSS 0.105768f
C17473 VDAC_N.n1818 VSS 0.132739f
C17474 VDAC_N.t607 VSS 0.105768f
C17475 VDAC_N.n1819 VSS 0.132739f
C17476 VDAC_N.t1936 VSS 0.105768f
C17477 VDAC_N.n1820 VSS 0.132739f
C17478 VDAC_N.t978 VSS 0.105768f
C17479 VDAC_N.n1821 VSS 0.132739f
C17480 VDAC_N.t1437 VSS 0.105768f
C17481 VDAC_N.n1822 VSS 0.132739f
C17482 VDAC_N.t862 VSS 0.105768f
C17483 VDAC_N.n1823 VSS 0.132739f
C17484 VDAC_N.t679 VSS 0.105768f
C17485 VDAC_N.n1824 VSS 0.132739f
C17486 VDAC_N.t83 VSS 0.105768f
C17487 VDAC_N.n1825 VSS 0.132739f
C17488 VDAC_N.t1219 VSS 0.105768f
C17489 VDAC_N.n1826 VSS 0.132739f
C17490 VDAC_N.t1683 VSS 0.105768f
C17491 VDAC_N.n1827 VSS 0.132739f
C17492 VDAC_N.t1982 VSS 0.105768f
C17493 VDAC_N.n1828 VSS 0.132739f
C17494 VDAC_N.t413 VSS 0.105768f
C17495 VDAC_N.n1829 VSS 0.132739f
C17496 VDAC_N.t2031 VSS 0.105768f
C17497 VDAC_N.n1830 VSS 0.132739f
C17498 VDAC_N.t1603 VSS 0.105768f
C17499 VDAC_N.n1831 VSS 0.132739f
C17500 VDAC_N.t155 VSS 0.105768f
C17501 VDAC_N.n1832 VSS 0.132739f
C17502 VDAC_N.t1904 VSS 0.105768f
C17503 VDAC_N.n1833 VSS 0.132739f
C17504 VDAC_N.t1945 VSS 0.105768f
C17505 VDAC_N.n1834 VSS 0.132739f
C17506 VDAC_N.t2068 VSS 0.105768f
C17507 VDAC_N.n1835 VSS 0.132739f
C17508 VDAC_N.t1674 VSS 0.105768f
C17509 VDAC_N.n1836 VSS 0.132739f
C17510 VDAC_N.t1156 VSS 0.105768f
C17511 VDAC_N.n1837 VSS 0.132739f
C17512 VDAC_N.t1242 VSS 0.105768f
C17513 VDAC_N.n1838 VSS 0.132739f
C17514 VDAC_N.t316 VSS 0.105768f
C17515 VDAC_N.n1839 VSS 0.132739f
C17516 VDAC_N.t2032 VSS 0.105768f
C17517 VDAC_N.n1840 VSS 0.132739f
C17518 VDAC_N.t270 VSS 0.105768f
C17519 VDAC_N.n1841 VSS 0.132739f
C17520 VDAC_N.t1168 VSS 0.105768f
C17521 VDAC_N.n1842 VSS 0.132739f
C17522 VDAC_N.t242 VSS 0.105768f
C17523 VDAC_N.n1843 VSS 0.132739f
C17524 VDAC_N.t691 VSS 0.105768f
C17525 VDAC_N.n1844 VSS 0.132739f
C17526 VDAC_N.t662 VSS 0.105768f
C17527 VDAC_N.n1845 VSS 0.132739f
C17528 VDAC_N.t1237 VSS 0.105768f
C17529 VDAC_N.n1846 VSS 0.132739f
C17530 VDAC_N.t1086 VSS 0.105768f
C17531 VDAC_N.n1847 VSS 0.132739f
C17532 VDAC_N.t2022 VSS 0.105768f
C17533 VDAC_N.n1848 VSS 0.132739f
C17534 VDAC_N.t811 VSS 0.105768f
C17535 VDAC_N.n1849 VSS 0.132739f
C17536 VDAC_N.t250 VSS 0.105768f
C17537 VDAC_N.n1850 VSS 0.132739f
C17538 VDAC_N.t1381 VSS 0.105768f
C17539 VDAC_N.n1851 VSS 0.132739f
C17540 VDAC_N.t1839 VSS 0.105768f
C17541 VDAC_N.n1852 VSS 0.132739f
C17542 VDAC_N.t1267 VSS 0.105768f
C17543 VDAC_N.n1853 VSS 0.132739f
C17544 VDAC_N.t879 VSS 0.105768f
C17545 VDAC_N.n1854 VSS 0.132739f
C17546 VDAC_N.t30 VSS 0.105768f
C17547 VDAC_N.n1855 VSS 0.132739f
C17548 VDAC_N.t1623 VSS 0.105768f
C17549 VDAC_N.n1856 VSS 0.132739f
C17550 VDAC_N.t2083 VSS 0.105768f
C17551 VDAC_N.n1857 VSS 0.132739f
C17552 VDAC_N.t393 VSS 0.105768f
C17553 VDAC_N.n1858 VSS 0.132739f
C17554 VDAC_N.t2055 VSS 0.105768f
C17555 VDAC_N.n1859 VSS 0.132739f
C17556 VDAC_N.t1448 VSS 0.105768f
C17557 VDAC_N.n1860 VSS 0.132739f
C17558 VDAC_N.t1845 VSS 0.105768f
C17559 VDAC_N.n1861 VSS 0.132739f
C17560 VDAC_N.t1108 VSS 0.105768f
C17561 VDAC_N.n1862 VSS 0.132739f
C17562 VDAC_N.t734 VSS 0.105768f
C17563 VDAC_N.n1863 VSS 0.132739f
C17564 VDAC_N.t554 VSS 0.105768f
C17565 VDAC_N.n1864 VSS 0.132739f
C17566 VDAC_N.t152 VSS 0.105768f
C17567 VDAC_N.n1865 VSS 0.132739f
C17568 VDAC_N.t2087 VSS 0.105768f
C17569 VDAC_N.n1866 VSS 0.132739f
C17570 VDAC_N.t1568 VSS 0.105768f
C17571 VDAC_N.n1867 VSS 0.132739f
C17572 VDAC_N.t1730 VSS 0.105768f
C17573 VDAC_N.n1868 VSS 0.132739f
C17574 VDAC_N.t304 VSS 0.105768f
C17575 VDAC_N.n1869 VSS 0.132739f
C17576 VDAC_N.t1514 VSS 0.105768f
C17577 VDAC_N.n1870 VSS 0.132739f
C17578 VDAC_N.t1231 VSS 0.105768f
C17579 VDAC_N.n1871 VSS 0.132739f
C17580 VDAC_N.t1072 VSS 0.105768f
C17581 VDAC_N.n1872 VSS 0.132739f
C17582 VDAC_N.t1123 VSS 0.105768f
C17583 VDAC_N.n1873 VSS 0.132739f
C17584 VDAC_N.t448 VSS 0.105768f
C17585 VDAC_N.n1874 VSS 0.132739f
C17586 VDAC_N.t1794 VSS 0.105768f
C17587 VDAC_N.n1875 VSS 0.132739f
C17588 VDAC_N.t1475 VSS 0.105768f
C17589 VDAC_N.n1876 VSS 0.132739f
C17590 VDAC_N.t1582 VSS 0.105768f
C17591 VDAC_N.n1877 VSS 0.132739f
C17592 VDAC_N.t645 VSS 0.105768f
C17593 VDAC_N.n1878 VSS 0.132739f
C17594 VDAC_N.t479 VSS 0.105768f
C17595 VDAC_N.n1879 VSS 0.132739f
C17596 VDAC_N.t1157 VSS 0.105768f
C17597 VDAC_N.n1880 VSS 0.12675f
C17598 VDAC_N.t455 VSS 0.105768f
C17599 VDAC_N.n1881 VSS 0.132739f
C17600 VDAC_N.t564 VSS 0.105768f
C17601 VDAC_N.n1882 VSS 0.132739f
C17602 VDAC_N.t53 VSS 0.105768f
C17603 VDAC_N.n1883 VSS 0.132739f
C17604 VDAC_N.t2089 VSS 0.105768f
C17605 VDAC_N.n1884 VSS 0.132739f
C17606 VDAC_N.t1576 VSS 0.105768f
C17607 VDAC_N.n1885 VSS 0.132739f
C17608 VDAC_N.t1977 VSS 0.105768f
C17609 VDAC_N.n1886 VSS 0.132739f
C17610 VDAC_N.t1144 VSS 0.105768f
C17611 VDAC_N.n1887 VSS 0.132739f
C17612 VDAC_N.t1518 VSS 0.105768f
C17613 VDAC_N.n1888 VSS 0.132739f
C17614 VDAC_N.t196 VSS 0.105768f
C17615 VDAC_N.n1889 VSS 0.132739f
C17616 VDAC_N.t658 VSS 0.105768f
C17617 VDAC_N.n1890 VSS 0.132739f
C17618 VDAC_N.t2119 VSS 0.105768f
C17619 VDAC_N.n1891 VSS 0.132739f
C17620 VDAC_N.t288 VSS 0.105768f
C17621 VDAC_N.n1892 VSS 0.132739f
C17622 VDAC_N.t90 VSS 0.105768f
C17623 VDAC_N.n1893 VSS 0.132739f
C17624 VDAC_N.t1284 VSS 0.105768f
C17625 VDAC_N.n1894 VSS 0.132739f
C17626 VDAC_N.t338 VSS 0.105768f
C17627 VDAC_N.n1895 VSS 0.132739f
C17628 VDAC_N.t1225 VSS 0.105768f
C17629 VDAC_N.n1896 VSS 0.132739f
C17630 VDAC_N.t32 VSS 0.105768f
C17631 VDAC_N.n1897 VSS 0.132739f
C17632 VDAC_N.t274 VSS 0.105768f
C17633 VDAC_N.n1898 VSS 0.132739f
C17634 VDAC_N.t415 VSS 0.105768f
C17635 VDAC_N.n1899 VSS 0.132739f
C17636 VDAC_N.t1762 VSS 0.105768f
C17637 VDAC_N.n1900 VSS 0.132739f
C17638 VDAC_N.t697 VSS 0.105768f
C17639 VDAC_N.n1901 VSS 0.132739f
C17640 VDAC_N.t1554 VSS 0.105768f
C17641 VDAC_N.n1902 VSS 0.132739f
C17642 VDAC_N.t181 VSS 0.105768f
C17643 VDAC_N.n1903 VSS 0.132739f
C17644 VDAC_N.t1713 VSS 0.105768f
C17645 VDAC_N.n1904 VSS 0.132739f
C17646 VDAC_N.t2046 VSS 0.105768f
C17647 VDAC_N.n1905 VSS 0.132739f
C17648 VDAC_N.t1607 VSS 0.105768f
C17649 VDAC_N.n1906 VSS 0.132739f
C17650 VDAC_N.t2067 VSS 0.105768f
C17651 VDAC_N.n1907 VSS 0.132739f
C17652 VDAC_N.t1395 VSS 0.105768f
C17653 VDAC_N.n1908 VSS 0.132739f
C17654 VDAC_N.t989 VSS 0.105768f
C17655 VDAC_N.n1909 VSS 0.132739f
C17656 VDAC_N.t341 VSS 0.105768f
C17657 VDAC_N.n1910 VSS 0.132739f
C17658 VDAC_N.t1745 VSS 0.105768f
C17659 VDAC_N.n1911 VSS 0.132739f
C17660 VDAC_N.t612 VSS 0.105768f
C17661 VDAC_N.n1912 VSS 0.132739f
C17662 VDAC_N.t833 VSS 0.105768f
C17663 VDAC_N.n1913 VSS 0.132739f
C17664 VDAC_N.t2095 VSS 0.105768f
C17665 VDAC_N.n1914 VSS 0.132739f
C17666 VDAC_N.t424 VSS 0.105768f
C17667 VDAC_N.n1915 VSS 0.132739f
C17668 VDAC_N.t1985 VSS 0.105768f
C17669 VDAC_N.n1916 VSS 0.132739f
C17670 VDAC_N.t64 VSS 0.105768f
C17671 VDAC_N.n1917 VSS 0.132739f
C17672 VDAC_N.t1769 VSS 0.105768f
C17673 VDAC_N.n1918 VSS 0.132739f
C17674 VDAC_N.t1444 VSS 0.105768f
C17675 VDAC_N.n1919 VSS 0.132739f
C17676 VDAC_N.t1302 VSS 0.105768f
C17677 VDAC_N.n1920 VSS 0.132739f
C17678 VDAC_N.t380 VSS 0.105768f
C17679 VDAC_N.n1921 VSS 0.132739f
C17680 VDAC_N.t1254 VSS 0.105768f
C17681 VDAC_N.n1922 VSS 0.132739f
C17682 VDAC_N.t1105 VSS 0.105768f
C17683 VDAC_N.n1923 VSS 0.132739f
C17684 VDAC_N.t832 VSS 0.105768f
C17685 VDAC_N.n1924 VSS 0.132739f
C17686 VDAC_N.t458 VSS 0.105768f
C17687 VDAC_N.n1925 VSS 0.132739f
C17688 VDAC_N.t1463 VSS 0.105768f
C17689 VDAC_N.n1926 VSS 0.132739f
C17690 VDAC_N.t786 VSS 0.105768f
C17691 VDAC_N.n1927 VSS 0.132739f
C17692 VDAC_N.t1247 VSS 0.105768f
C17693 VDAC_N.n1928 VSS 0.132739f
C17694 VDAC_N.t38 VSS 0.105768f
C17695 VDAC_N.n1929 VSS 0.132739f
C17696 VDAC_N.t305 VSS 0.105768f
C17697 VDAC_N.n1930 VSS 0.132739f
C17698 VDAC_N.t815 VSS 0.105768f
C17699 VDAC_N.n1931 VSS 0.132739f
C17700 VDAC_N.t1030 VSS 0.105768f
C17701 VDAC_N.n1932 VSS 0.132739f
C17702 VDAC_N.t1493 VSS 0.105768f
C17703 VDAC_N.n1933 VSS 0.132739f
C17704 VDAC_N.t507 VSS 0.105768f
C17705 VDAC_N.n1934 VSS 0.132739f
C17706 VDAC_N.t651 VSS 0.105768f
C17707 VDAC_N.n1935 VSS 0.132739f
C17708 VDAC_N.t1851 VSS 0.105768f
C17709 VDAC_N.n1936 VSS 0.132739f
C17710 VDAC_N.t313 VSS 0.105768f
C17711 VDAC_N.n1937 VSS 0.132739f
C17712 VDAC_N.t1633 VSS 0.105768f
C17713 VDAC_N.n1938 VSS 0.132739f
C17714 VDAC_N.t572 VSS 0.105768f
C17715 VDAC_N.n1939 VSS 0.132739f
C17716 VDAC_N.t775 VSS 0.105768f
C17717 VDAC_N.n1940 VSS 0.132739f
C17718 VDAC_N.t89 VSS 0.105768f
C17719 VDAC_N.n1941 VSS 0.132739f
C17720 VDAC_N.t1584 VSS 0.105768f
C17721 VDAC_N.n1942 VSS 0.132739f
C17722 VDAC_N.t491 VSS 0.105768f
C17723 VDAC_N.n1943 VSS 0.12675f
C17724 VDAC_N.t372 VSS 0.105768f
C17725 VDAC_N.n1944 VSS 0.142694f
C17726 VDAC_N.t1615 VSS 0.105768f
C17727 VDAC_N.n1945 VSS 0.142694f
C17728 VDAC_N.t917 VSS 0.105768f
C17729 VDAC_N.n1946 VSS 0.142694f
C17730 VDAC_N.t1993 VSS 0.105768f
C17731 VDAC_N.n1947 VSS 0.142694f
C17732 VDAC_N.t67 VSS 0.105768f
C17733 VDAC_N.n1948 VSS 0.142694f
C17734 VDAC_N.t1467 VSS 0.105768f
C17735 VDAC_N.n1949 VSS 0.142694f
C17736 VDAC_N.t742 VSS 0.105768f
C17737 VDAC_N.n1950 VSS 0.142694f
C17738 VDAC_N.t1850 VSS 0.105768f
C17739 VDAC_N.n1951 VSS 0.142694f
C17740 VDAC_N.t303 VSS 0.105768f
C17741 VDAC_N.n1952 VSS 0.142694f
C17742 VDAC_N.t216 VSS 0.105768f
C17743 VDAC_N.n1953 VSS 0.142694f
C17744 VDAC_N.t170 VSS 0.105768f
C17745 VDAC_N.n1954 VSS 0.142694f
C17746 VDAC_N.t2007 VSS 0.105768f
C17747 VDAC_N.n1955 VSS 0.142694f
C17748 VDAC_N.t1276 VSS 0.105768f
C17749 VDAC_N.n1956 VSS 0.142694f
C17750 VDAC_N.t1876 VSS 0.105768f
C17751 VDAC_N.n1957 VSS 0.142694f
C17752 VDAC_N.t1679 VSS 0.105768f
C17753 VDAC_N.n1958 VSS 0.142694f
C17754 VDAC_N.t1869 VSS 0.105768f
C17755 VDAC_N.n1959 VSS 0.142694f
C17756 VDAC_N.t587 VSS 0.105768f
C17757 VDAC_N.n1960 VSS 0.142694f
C17758 VDAC_N.t1343 VSS 0.105768f
C17759 VDAC_N.n1961 VSS 0.142694f
C17760 VDAC_N.t1527 VSS 0.105768f
C17761 VDAC_N.n1962 VSS 0.142694f
C17762 VDAC_N.t439 VSS 0.105768f
C17763 VDAC_N.n1963 VSS 0.142694f
C17764 VDAC_N.t487 VSS 0.105768f
C17765 VDAC_N.n1964 VSS 0.142694f
C17766 VDAC_N.t583 VSS 0.105768f
C17767 VDAC_N.n1965 VSS 0.142694f
C17768 VDAC_N.t355 VSS 0.105768f
C17769 VDAC_N.n1966 VSS 0.142694f
C17770 VDAC_N.t215 VSS 0.105768f
C17771 VDAC_N.n1967 VSS 0.142694f
C17772 VDAC_N.t806 VSS 0.105768f
C17773 VDAC_N.n1968 VSS 0.142694f
C17774 VDAC_N.t1966 VSS 0.105768f
C17775 VDAC_N.n1969 VSS 0.142694f
C17776 VDAC_N.t148 VSS 0.105768f
C17777 VDAC_N.n1970 VSS 0.142694f
C17778 VDAC_N.t1768 VSS 0.105768f
C17779 VDAC_N.n1971 VSS 0.142694f
C17780 VDAC_N.t106 VSS 0.105768f
C17781 VDAC_N.n1972 VSS 0.137176f
C17782 VDAC_N.t2065 VSS 0.105768f
C17783 VDAC_N.n1973 VSS 0.126358f
C17784 VDAC_N.t817 VSS 0.105768f
C17785 VDAC_N.n1974 VSS 0.132739f
C17786 VDAC_N.t492 VSS 0.105768f
C17787 VDAC_N.n1975 VSS 0.132739f
C17788 VDAC_N.t449 VSS 0.105768f
C17789 VDAC_N.n1976 VSS 0.132739f
C17790 VDAC_N.t639 VSS 0.105768f
C17791 VDAC_N.n1977 VSS 0.132739f
C17792 VDAC_N.t977 VSS 0.105768f
C17793 VDAC_N.n1978 VSS 0.132739f
C17794 VDAC_N.t195 VSS 0.105768f
C17795 VDAC_N.n1979 VSS 0.132739f
C17796 VDAC_N.t1758 VSS 0.105768f
C17797 VDAC_N.n1980 VSS 0.132739f
C17798 VDAC_N.t1575 VSS 0.105768f
C17799 VDAC_N.n1981 VSS 0.132739f
C17800 VDAC_N.t1010 VSS 0.105768f
C17801 VDAC_N.n1982 VSS 0.132739f
C17802 VDAC_N.t859 VSS 0.105768f
C17803 VDAC_N.n1983 VSS 0.132739f
C17804 VDAC_N.t327 VSS 0.105768f
C17805 VDAC_N.n1984 VSS 0.132739f
C17806 VDAC_N.t390 VSS 0.105768f
C17807 VDAC_N.n1985 VSS 0.132739f
C17808 VDAC_N.t1333 VSS 0.105768f
C17809 VDAC_N.n1986 VSS 0.132739f
C17810 VDAC_N.t866 VSS 0.105768f
C17811 VDAC_N.n1987 VSS 0.132739f
C17812 VDAC_N.t1504 VSS 0.105768f
C17813 VDAC_N.n1988 VSS 0.132739f
C17814 VDAC_N.t1934 VSS 0.105768f
C17815 VDAC_N.n1989 VSS 0.132739f
C17816 VDAC_N.t88 VSS 0.105768f
C17817 VDAC_N.n1990 VSS 0.132739f
C17818 VDAC_N.t609 VSS 0.105768f
C17819 VDAC_N.n1991 VSS 0.132739f
C17820 VDAC_N.t1210 VSS 0.105768f
C17821 VDAC_N.n1992 VSS 0.132739f
C17822 VDAC_N.t1964 VSS 0.105768f
C17823 VDAC_N.n1993 VSS 0.132739f
C17824 VDAC_N.t834 VSS 0.105768f
C17825 VDAC_N.n1994 VSS 0.132739f
C17826 VDAC_N.t1392 VSS 0.105768f
C17827 VDAC_N.n1995 VSS 0.132739f
C17828 VDAC_N.t147 VSS 0.105768f
C17829 VDAC_N.n1996 VSS 0.132739f
C17830 VDAC_N.t1488 VSS 0.105768f
C17831 VDAC_N.n1997 VSS 0.132739f
C17832 VDAC_N.t2069 VSS 0.105768f
C17833 VDAC_N.n1998 VSS 0.132739f
C17834 VDAC_N.t51 VSS 0.105768f
C17835 VDAC_N.n1999 VSS 0.132739f
C17836 VDAC_N.t1308 VSS 0.105768f
C17837 VDAC_N.n2000 VSS 0.132739f
C17838 VDAC_N.t1715 VSS 0.105768f
C17839 VDAC_N.n2001 VSS 0.132739f
C17840 VDAC_N.t1932 VSS 0.105768f
C17841 VDAC_N.n2002 VSS 0.132739f
C17842 VDAC_N.t927 VSS 0.105768f
C17843 VDAC_N.n2003 VSS 0.132739f
C17844 VDAC_N.t699 VSS 0.105768f
C17845 VDAC_N.n2004 VSS 0.132739f
C17846 VDAC_N.t531 VSS 0.105768f
C17847 VDAC_N.n2005 VSS 0.132739f
C17848 VDAC_N.t749 VSS 0.105768f
C17849 VDAC_N.n2006 VSS 0.132739f
C17850 VDAC_N.t522 VSS 0.105768f
C17851 VDAC_N.n2007 VSS 0.132739f
C17852 VDAC_N.t1695 VSS 0.105768f
C17853 VDAC_N.n2008 VSS 0.132739f
C17854 VDAC_N.t571 VSS 0.105768f
C17855 VDAC_N.n2009 VSS 0.132739f
C17856 VDAC_N.t249 VSS 0.105768f
C17857 VDAC_N.n2010 VSS 0.132739f
C17858 VDAC_N.t69 VSS 0.105768f
C17859 VDAC_N.n2011 VSS 0.132739f
C17860 VDAC_N.t394 VSS 0.105768f
C17861 VDAC_N.n2012 VSS 0.132739f
C17862 VDAC_N.t205 VSS 0.105768f
C17863 VDAC_N.n2013 VSS 0.132739f
C17864 VDAC_N.t1946 VSS 0.105768f
C17865 VDAC_N.n2014 VSS 0.132739f
C17866 VDAC_N.t272 VSS 0.105768f
C17867 VDAC_N.n2015 VSS 0.132739f
C17868 VDAC_N.t29 VSS 0.105768f
C17869 VDAC_N.n2016 VSS 0.132739f
C17870 VDAC_N.t326 VSS 0.105768f
C17871 VDAC_N.n2017 VSS 0.132739f
C17872 VDAC_N.t1307 VSS 0.105768f
C17873 VDAC_N.n2018 VSS 0.132739f
C17874 VDAC_N.t1426 VSS 0.105768f
C17875 VDAC_N.n2019 VSS 0.132739f
C17876 VDAC_N.t1972 VSS 0.105768f
C17877 VDAC_N.n2020 VSS 0.132739f
C17878 VDAC_N.t1870 VSS 0.105768f
C17879 VDAC_N.n2021 VSS 0.132739f
C17880 VDAC_N.t1416 VSS 0.105768f
C17881 VDAC_N.n2022 VSS 0.132739f
C17882 VDAC_N.t2051 VSS 0.105768f
C17883 VDAC_N.n2023 VSS 0.132739f
C17884 VDAC_N.t279 VSS 0.105768f
C17885 VDAC_N.n2024 VSS 0.132739f
C17886 VDAC_N.t221 VSS 0.105768f
C17887 VDAC_N.n2025 VSS 0.132739f
C17888 VDAC_N.t1990 VSS 0.105768f
C17889 VDAC_N.n2026 VSS 0.132739f
C17890 VDAC_N.t1687 VSS 0.105768f
C17891 VDAC_N.n2027 VSS 0.132739f
C17892 VDAC_N.t625 VSS 0.105768f
C17893 VDAC_N.n2028 VSS 0.132739f
C17894 VDAC_N.t1789 VSS 0.105768f
C17895 VDAC_N.n2029 VSS 0.132739f
C17896 VDAC_N.t1331 VSS 0.105768f
C17897 VDAC_N.n2030 VSS 0.132739f
C17898 VDAC_N.t1702 VSS 0.105768f
C17899 VDAC_N.n2031 VSS 0.132739f
C17900 VDAC_N.t733 VSS 0.105768f
C17901 VDAC_N.n2032 VSS 0.132739f
C17902 VDAC_N.t1930 VSS 0.105768f
C17903 VDAC_N.n2033 VSS 0.132739f
C17904 VDAC_N.t1944 VSS 0.105768f
C17905 VDAC_N.n2034 VSS 0.132739f
C17906 VDAC_N.t173 VSS 0.105768f
C17907 VDAC_N.n2035 VSS 0.132739f
C17908 VDAC_N.t1206 VSS 0.105768f
C17909 VDAC_N.n2036 VSS 0.132739f
C17910 VDAC_N.t1301 VSS 0.105768f
C17911 VDAC_N.n2037 VSS 0.132739f
C17912 VDAC_N.t1638 VSS 0.105768f
C17913 VDAC_N.n2038 VSS 0.127945f
C17914 VDAC_N.t985 VSS 0.105768f
C17915 VDAC_N.n2039 VSS 0.138762f
C17916 VDAC_N.t315 VSS 0.105768f
C17917 VDAC_N.n2040 VSS 0.144281f
C17918 VDAC_N.t760 VSS 0.105768f
C17919 VDAC_N.n2041 VSS 0.144281f
C17920 VDAC_N.t1517 VSS 0.105768f
C17921 VDAC_N.n2042 VSS 0.144281f
C17922 VDAC_N.t50 VSS 0.105768f
C17923 VDAC_N.n2043 VSS 0.144281f
C17924 VDAC_N.t1857 VSS 0.105768f
C17925 VDAC_N.n2044 VSS 0.144281f
C17926 VDAC_N.t15 VSS 0.105768f
C17927 VDAC_N.n2045 VSS 0.144281f
C17928 VDAC_N.t1120 VSS 0.105768f
C17929 VDAC_N.n2046 VSS 0.144281f
C17930 VDAC_N.t115 VSS 0.105768f
C17931 VDAC_N.n2047 VSS 0.144281f
C17932 VDAC_N.t334 VSS 0.105768f
C17933 VDAC_N.n2048 VSS 0.144281f
C17934 VDAC_N.t536 VSS 0.105768f
C17935 VDAC_N.n2049 VSS 0.144281f
C17936 VDAC_N.t963 VSS 0.105768f
C17937 VDAC_N.n2050 VSS 0.144281f
C17938 VDAC_N.t1119 VSS 0.105768f
C17939 VDAC_N.n2051 VSS 0.144281f
C17940 VDAC_N.t1196 VSS 0.105768f
C17941 VDAC_N.n2052 VSS 0.144281f
C17942 VDAC_N.t745 VSS 0.105768f
C17943 VDAC_N.n2053 VSS 0.144281f
C17944 VDAC_N.t1696 VSS 0.105768f
C17945 VDAC_N.n2054 VSS 0.144281f
C17946 VDAC_N.t1801 VSS 0.105768f
C17947 VDAC_N.n2055 VSS 0.144281f
C17948 VDAC_N.t2026 VSS 0.105768f
C17949 VDAC_N.n2056 VSS 0.144281f
C17950 VDAC_N.t1187 VSS 0.105768f
C17951 VDAC_N.n2057 VSS 0.144281f
C17952 VDAC_N.t1373 VSS 0.105768f
C17953 VDAC_N.n2058 VSS 0.144281f
C17954 VDAC_N.t344 VSS 0.105768f
C17955 VDAC_N.n2059 VSS 0.144281f
C17956 VDAC_N.t133 VSS 0.105768f
C17957 VDAC_N.n2060 VSS 0.144281f
C17958 VDAC_N.t930 VSS 0.105768f
C17959 VDAC_N.n2061 VSS 0.144281f
C17960 VDAC_N.t91 VSS 0.105768f
C17961 VDAC_N.n2062 VSS 0.144281f
C17962 VDAC_N.t1269 VSS 0.105768f
C17963 VDAC_N.n2063 VSS 0.144281f
C17964 VDAC_N.t916 VSS 0.105768f
C17965 VDAC_N.n2064 VSS 0.144281f
C17966 VDAC_N.t1611 VSS 0.105768f
C17967 VDAC_N.n2065 VSS 0.144281f
C17968 VDAC_N.t430 VSS 0.105768f
C17969 VDAC_N.n2066 VSS 0.144281f
C17970 VDAC_N.t1941 VSS 0.105768f
C17971 VDAC_N.n2067 VSS 0.144281f
C17972 VDAC_N.t1173 VSS 0.105768f
C17973 VDAC_N.n2068 VSS 0.138762f
C17974 VDAC_N.t268 VSS 0.105768f
C17975 VDAC_N.n2069 VSS 0.127945f
C17976 VDAC_N.t322 VSS 0.105768f
C17977 VDAC_N.n2070 VSS 0.132739f
C17978 VDAC_N.t1051 VSS 0.105768f
C17979 VDAC_N.n2071 VSS 0.132739f
C17980 VDAC_N.t984 VSS 0.105768f
C17981 VDAC_N.n2072 VSS 0.132739f
C17982 VDAC_N.t1959 VSS 0.105768f
C17983 VDAC_N.n2073 VSS 0.132739f
C17984 VDAC_N.t160 VSS 0.105768f
C17985 VDAC_N.n2074 VSS 0.132739f
C17986 VDAC_N.t1478 VSS 0.105768f
C17987 VDAC_N.n2075 VSS 0.132739f
C17988 VDAC_N.t340 VSS 0.105768f
C17989 VDAC_N.n2076 VSS 0.132739f
C17990 VDAC_N.t182 VSS 0.105768f
C17991 VDAC_N.n2077 VSS 0.132739f
C17992 VDAC_N.t163 VSS 0.105768f
C17993 VDAC_N.n2078 VSS 0.132739f
C17994 VDAC_N.t1048 VSS 0.105768f
C17995 VDAC_N.n2079 VSS 0.132739f
C17996 VDAC_N.t1986 VSS 0.105768f
C17997 VDAC_N.n2080 VSS 0.132739f
C17998 VDAC_N.t624 VSS 0.105768f
C17999 VDAC_N.n2081 VSS 0.132739f
C18000 VDAC_N.t1754 VSS 0.105768f
C18001 VDAC_N.n2082 VSS 0.132739f
C18002 VDAC_N.t695 VSS 0.105768f
C18003 VDAC_N.n2083 VSS 0.132739f
C18004 VDAC_N.t1402 VSS 0.105768f
C18005 VDAC_N.n2084 VSS 0.132739f
C18006 VDAC_N.t1181 VSS 0.105768f
C18007 VDAC_N.n2085 VSS 0.132739f
C18008 VDAC_N.t1755 VSS 0.105768f
C18009 VDAC_N.n2086 VSS 0.132739f
C18010 VDAC_N.t1070 VSS 0.105768f
C18011 VDAC_N.n2087 VSS 0.132739f
C18012 VDAC_N.t783 VSS 0.105768f
C18013 VDAC_N.n2088 VSS 0.132739f
C18014 VDAC_N.t1065 VSS 0.105768f
C18015 VDAC_N.n2089 VSS 0.132739f
C18016 VDAC_N.t1429 VSS 0.105768f
C18017 VDAC_N.n2090 VSS 0.132739f
C18018 VDAC_N.t1891 VSS 0.105768f
C18019 VDAC_N.n2091 VSS 0.132739f
C18020 VDAC_N.t1325 VSS 0.105768f
C18021 VDAC_N.n2092 VSS 0.132739f
C18022 VDAC_N.t905 VSS 0.105768f
C18023 VDAC_N.n2093 VSS 0.132739f
C18024 VDAC_N.t108 VSS 0.105768f
C18025 VDAC_N.n2094 VSS 0.132739f
C18026 VDAC_N.t797 VSS 0.105768f
C18027 VDAC_N.n2095 VSS 0.132739f
C18028 VDAC_N.t1081 VSS 0.105768f
C18029 VDAC_N.n2096 VSS 0.132739f
C18030 VDAC_N.t1776 VSS 0.105768f
C18031 VDAC_N.n2097 VSS 0.132739f
C18032 VDAC_N.t973 VSS 0.105768f
C18033 VDAC_N.n2098 VSS 0.132739f
C18034 VDAC_N.t1320 VSS 0.105768f
C18035 VDAC_N.n2099 VSS 0.132739f
C18036 VDAC_N.t251 VSS 0.105768f
C18037 VDAC_N.n2100 VSS 0.132739f
C18038 VDAC_N.t1740 VSS 0.105768f
C18039 VDAC_N.n2101 VSS 0.132739f
C18040 VDAC_N.t70 VSS 0.105768f
C18041 VDAC_N.n2102 VSS 0.132739f
C18042 VDAC_N.t668 VSS 0.105768f
C18043 VDAC_N.n2103 VSS 0.132739f
C18044 VDAC_N.t1888 VSS 0.105768f
C18045 VDAC_N.n2104 VSS 0.132739f
C18046 VDAC_N.t1882 VSS 0.105768f
C18047 VDAC_N.n2105 VSS 0.132739f
C18048 VDAC_N.t736 VSS 0.105768f
C18049 VDAC_N.n2106 VSS 0.132739f
C18050 VDAC_N.t130 VSS 0.105768f
C18051 VDAC_N.n2107 VSS 0.132739f
C18052 VDAC_N.t292 VSS 0.105768f
C18053 VDAC_N.n2108 VSS 0.132739f
C18054 VDAC_N.t1434 VSS 0.105768f
C18055 VDAC_N.n2109 VSS 0.132739f
C18056 VDAC_N.t1201 VSS 0.105768f
C18057 VDAC_N.n2110 VSS 0.132739f
C18058 VDAC_N.t1174 VSS 0.105768f
C18059 VDAC_N.n2111 VSS 0.132739f
C18060 VDAC_N.t1175 VSS 0.105768f
C18061 VDAC_N.n2112 VSS 0.132739f
C18062 VDAC_N.t1641 VSS 0.105768f
C18063 VDAC_N.n2113 VSS 0.132739f
C18064 VDAC_N.t1898 VSS 0.105768f
C18065 VDAC_N.n2114 VSS 0.132739f
C18066 VDAC_N.t725 VSS 0.105768f
C18067 VDAC_N.n2115 VSS 0.132739f
C18068 VDAC_N.t1987 VSS 0.105768f
C18069 VDAC_N.n2116 VSS 0.132739f
C18070 VDAC_N.t1319 VSS 0.105768f
C18071 VDAC_N.n2117 VSS 0.132739f
C18072 VDAC_N.t901 VSS 0.105768f
C18073 VDAC_N.n2118 VSS 0.132739f
C18074 VDAC_N.t617 VSS 0.105768f
C18075 VDAC_N.n2119 VSS 0.132739f
C18076 VDAC_N.t849 VSS 0.105768f
C18077 VDAC_N.n2120 VSS 0.132739f
C18078 VDAC_N.t553 VSS 0.105768f
C18079 VDAC_N.n2121 VSS 0.132739f
C18080 VDAC_N.t411 VSS 0.105768f
C18081 VDAC_N.n2122 VSS 0.132739f
C18082 VDAC_N.t525 VSS 0.105768f
C18083 VDAC_N.n2123 VSS 0.132739f
C18084 VDAC_N.t1296 VSS 0.105768f
C18085 VDAC_N.n2124 VSS 0.132739f
C18086 VDAC_N.t1805 VSS 0.105768f
C18087 VDAC_N.n2125 VSS 0.132739f
C18088 VDAC_N.t1716 VSS 0.105768f
C18089 VDAC_N.n2126 VSS 0.132739f
C18090 VDAC_N.t447 VSS 0.105768f
C18091 VDAC_N.n2127 VSS 0.132739f
C18092 VDAC_N.t604 VSS 0.105768f
C18093 VDAC_N.n2128 VSS 0.132739f
C18094 VDAC_N.t1154 VSS 0.105768f
C18095 VDAC_N.n2129 VSS 0.132739f
C18096 VDAC_N.t1039 VSS 0.105768f
C18097 VDAC_N.n2130 VSS 0.132739f
C18098 VDAC_N.t720 VSS 0.105768f
C18099 VDAC_N.n2131 VSS 0.132739f
C18100 VDAC_N.t1866 VSS 0.105768f
C18101 VDAC_N.n2132 VSS 0.132739f
C18102 VDAC_N.t996 VSS 0.105768f
C18103 VDAC_N.n2133 VSS 0.132739f
C18104 VDAC_N.t202 VSS 0.105768f
C18105 VDAC_N.n2134 VSS 0.134996f
C18106 a_n2661_46508.n1 VSS 0.733746f
C18107 a_n2661_46508.n3 VSS 0.407886f
C18108 a_n2661_46508.n4 VSS 11.685401f
C18109 a_n2661_46508.n5 VSS 0.132455f
.ends

