magic
tech sky130A
magscale 1 2
timestamp 1713724235
<< viali >>
rect 240 420 290 470
rect -770 240 -720 290
rect -660 240 -610 290
rect -40 240 10 290
rect 130 230 180 280
rect -220 160 -170 210
<< metal1 >>
rect 228 470 302 476
rect 228 460 240 470
rect -650 430 240 460
rect -790 240 -780 300
rect -720 296 -710 300
rect -650 296 -620 430
rect 228 420 240 430
rect 290 420 302 470
rect 228 414 302 420
rect -720 240 -708 296
rect -782 234 -708 240
rect -672 290 -598 296
rect -52 290 22 296
rect -672 240 -660 290
rect -610 240 -598 290
rect -672 234 -598 240
rect -650 200 -620 234
rect -60 230 -50 290
rect 10 234 22 290
rect 118 280 192 286
rect 10 230 20 234
rect 118 230 130 280
rect 180 230 192 280
rect 118 224 192 230
rect -230 216 -220 220
rect -670 140 -660 200
rect -600 140 -590 200
rect -232 160 -220 216
rect -160 195 -150 220
rect 138 195 168 224
rect -160 165 168 195
rect -160 160 -150 165
rect -232 154 -158 160
<< via1 >>
rect -780 290 -720 300
rect -780 240 -770 290
rect -770 240 -720 290
rect -50 240 -40 290
rect -40 240 10 290
rect -50 230 10 240
rect -660 140 -600 200
rect -220 210 -160 220
rect -220 160 -170 210
rect -170 160 -160 210
<< metal2 >>
rect -890 485 -615 515
rect -890 340 -745 370
rect -775 310 -745 340
rect -780 300 -720 310
rect -645 300 -615 485
rect -645 290 10 300
rect -645 270 -50 290
rect -780 230 -720 240
rect -220 220 -160 230
rect -50 220 10 230
rect -660 200 -600 210
rect -890 170 -660 200
rect -220 150 -160 160
rect -660 130 -600 140
rect -205 45 -175 150
rect -890 15 -175 45
use sky130_fd_sc_hd__and2_4  sky130_fd_sc_hd__and2_4_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 -792 0 1 28
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  sky130_fd_sc_hd__or2_4_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 -56 0 1 28
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 -148 0 1 28
box -38 -48 130 592
<< end >>
