magic
tech sky130A
magscale 1 2
timestamp 1715382157
<< metal1 >>
rect 1255 1785 1625 1795
rect 1255 1725 1259 1785
rect 1311 1725 1569 1785
rect 1621 1725 1625 1785
rect 1255 1525 1625 1725
rect 1255 1465 1259 1525
rect 1311 1465 1569 1525
rect 1621 1465 1625 1525
rect 1255 1455 1625 1465
<< via1 >>
rect 1259 1725 1311 1785
rect 1569 1725 1621 1785
rect 1259 1465 1311 1525
rect 1569 1465 1621 1525
<< metal2 >>
rect 1255 1785 1625 1795
rect 1255 1725 1259 1785
rect 1311 1765 1569 1785
rect 1255 1719 1311 1725
rect 1255 1531 1285 1719
rect 1340 1710 1540 1735
rect 1621 1725 1625 1785
rect 1569 1719 1625 1725
rect 1340 1690 1410 1710
rect 1315 1650 1410 1690
rect 1470 1690 1540 1710
rect 1470 1650 1565 1690
rect 1315 1600 1565 1650
rect 1315 1560 1410 1600
rect 1340 1540 1410 1560
rect 1470 1560 1565 1600
rect 1470 1540 1540 1560
rect 1255 1525 1311 1531
rect 1255 1465 1259 1525
rect 1340 1515 1540 1540
rect 1595 1531 1625 1719
rect 1569 1525 1625 1531
rect 1311 1465 1569 1485
rect 1621 1465 1625 1525
rect 1255 1455 1625 1465
<< via2 >>
rect 1410 1650 1470 1710
rect 1410 1540 1470 1600
<< metal3 >>
rect 1410 1715 1470 1810
rect 1400 1710 1480 1715
rect 1400 1650 1410 1710
rect 1470 1650 1480 1710
rect 1400 1600 1480 1650
rect 1400 1540 1410 1600
rect 1470 1540 1480 1600
rect 1400 1535 1480 1540
rect 1410 1440 1470 1535
<< end >>
