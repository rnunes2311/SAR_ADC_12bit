magic
tech sky130A
magscale 1 2
timestamp 1711974973
<< error_p >>
rect -29 481 29 487
rect -29 447 -17 481
rect -29 441 29 447
rect -29 -447 29 -441
rect -29 -481 -17 -447
rect -29 -487 29 -481
<< nwell >>
rect -211 -619 211 619
<< pmos >>
rect -15 -400 15 400
<< pdiff >>
rect -73 388 -15 400
rect -73 -388 -61 388
rect -27 -388 -15 388
rect -73 -400 -15 -388
rect 15 388 73 400
rect 15 -388 27 388
rect 61 -388 73 388
rect 15 -400 73 -388
<< pdiffc >>
rect -61 -388 -27 388
rect 27 -388 61 388
<< nsubdiff >>
rect -175 549 -79 583
rect 79 549 175 583
rect -175 487 -141 549
rect 141 487 175 549
rect -175 -549 -141 -487
rect 141 -549 175 -487
rect -175 -583 -79 -549
rect 79 -583 175 -549
<< nsubdiffcont >>
rect -79 549 79 583
rect -175 -487 -141 487
rect 141 -487 175 487
rect -79 -583 79 -549
<< poly >>
rect -33 481 33 497
rect -33 447 -17 481
rect 17 447 33 481
rect -33 431 33 447
rect -15 400 15 431
rect -15 -431 15 -400
rect -33 -447 33 -431
rect -33 -481 -17 -447
rect 17 -481 33 -447
rect -33 -497 33 -481
<< polycont >>
rect -17 447 17 481
rect -17 -481 17 -447
<< locali >>
rect -175 549 -79 583
rect 79 549 175 583
rect -175 487 -141 549
rect 141 487 175 549
rect -33 447 -17 481
rect 17 447 33 481
rect -61 388 -27 404
rect -61 -404 -27 -388
rect 27 388 61 404
rect 27 -404 61 -388
rect -33 -481 -17 -447
rect 17 -481 33 -447
rect -175 -549 -141 -487
rect 141 -549 175 -487
rect -175 -583 -79 -549
rect 79 -583 175 -549
<< viali >>
rect -17 447 17 481
rect -61 -388 -27 388
rect 27 -388 61 388
rect -17 -481 17 -447
<< metal1 >>
rect -29 481 29 487
rect -29 447 -17 481
rect 17 447 29 481
rect -29 441 29 447
rect -67 388 -21 400
rect -67 -388 -61 388
rect -27 -388 -21 388
rect -67 -400 -21 -388
rect 21 388 67 400
rect 21 -388 27 388
rect 61 -388 67 388
rect 21 -400 67 -388
rect -29 -447 29 -441
rect -29 -481 -17 -447
rect 17 -481 29 -447
rect -29 -487 29 -481
<< properties >>
string FIXED_BBOX -158 -566 158 566
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
