magic
tech sky130A
magscale 1 2
timestamp 1713893667
<< metal1 >>
rect 1740 10449 1770 11600
rect 1725 10439 1785 10449
rect 1780 10379 1785 10439
rect 1725 10369 1785 10379
rect 1815 10325 1845 11600
rect 1800 10315 1860 10325
rect 1855 10255 1860 10315
rect 1800 10245 1860 10255
rect 1725 10156 1785 10166
rect 1780 10096 1785 10156
rect 1725 10086 1785 10096
rect 1740 6360 1770 10086
rect 1800 10002 1860 10012
rect 1855 9942 1860 10002
rect 1800 9932 1860 9942
rect 1815 6360 1845 9932
rect 1890 9856 1920 11600
rect 1875 9846 1935 9856
rect 1930 9786 1935 9846
rect 1875 9776 1935 9786
rect 1965 9731 1995 11600
rect 1950 9721 2010 9731
rect 2005 9661 2010 9721
rect 1950 9651 2010 9661
rect 1875 9576 1935 9586
rect 1930 9516 1935 9576
rect 1875 9506 1935 9516
rect 1890 6360 1920 9506
rect 1950 9469 2010 9479
rect 2005 9409 2010 9469
rect 1950 9399 2010 9409
rect 1965 6360 1995 9399
rect 2040 9361 2070 11600
rect 2025 9351 2085 9361
rect 2080 9291 2085 9351
rect 2025 9281 2085 9291
rect 2115 9237 2145 11600
rect 2100 9227 2160 9237
rect 2155 9167 2160 9227
rect 2100 9157 2160 9167
rect 2025 9068 2085 9078
rect 2080 9008 2085 9068
rect 2025 8998 2085 9008
rect 2040 6360 2070 8998
rect 2100 8914 2160 8924
rect 2155 8854 2160 8914
rect 2100 8844 2160 8854
rect 2115 6360 2145 8844
rect 2190 8768 2220 11600
rect 2175 8758 2235 8768
rect 2230 8698 2235 8758
rect 2175 8688 2235 8698
rect 2265 8643 2295 11600
rect 2250 8633 2310 8643
rect 2305 8573 2310 8633
rect 2250 8563 2310 8573
rect 2175 8488 2235 8498
rect 2230 8428 2235 8488
rect 2175 8418 2235 8428
rect 2190 6360 2220 8418
rect 2250 8381 2310 8391
rect 2305 8321 2310 8381
rect 2250 8311 2310 8321
rect 2265 6360 2295 8311
rect 2341 8292 2370 11600
rect 2340 8273 2370 8292
rect 2325 8263 2385 8273
rect 2380 8203 2385 8263
rect 2325 8193 2385 8203
rect 2415 8149 2445 11600
rect 2400 8139 2460 8149
rect 2455 8079 2460 8139
rect 2400 8069 2460 8079
rect 2325 7980 2385 7990
rect 2380 7920 2385 7980
rect 2325 7910 2385 7920
rect 2340 6360 2370 7910
rect 2400 7826 2460 7836
rect 2455 7766 2460 7826
rect 2400 7756 2460 7766
rect 2415 6360 2445 7756
rect 2490 7680 2520 11600
rect 2475 7670 2535 7680
rect 2530 7610 2535 7670
rect 2475 7600 2535 7610
rect 2565 7555 2595 11600
rect 6107 11416 6167 11426
rect 5447 10672 5477 11410
rect 5522 11097 5552 11410
rect 5521 11090 5552 11097
rect 5506 11080 5566 11090
rect 5506 11020 5511 11080
rect 5506 11010 5566 11020
rect 5521 11002 5551 11010
rect 5446 10668 5477 10672
rect 5522 10974 5551 11002
rect 5431 10658 5491 10668
rect 5431 10598 5436 10658
rect 5431 10588 5491 10598
rect 5446 10575 5477 10588
rect 3760 10430 3770 10530
rect 3940 10430 3950 10530
rect 4090 9890 4100 9990
rect 4270 9890 4280 9990
rect 3760 9340 3770 9440
rect 3940 9340 3950 9440
rect 4090 8800 4100 8900
rect 4270 8800 4280 8900
rect 3760 8250 3770 8350
rect 3940 8250 3950 8350
rect 4090 7710 4100 7810
rect 4270 7710 4280 7810
rect 5447 7555 5477 10575
rect 5522 7680 5552 10974
rect 5597 10757 5627 11410
rect 5672 11181 5701 11410
rect 5671 11174 5701 11181
rect 5656 11164 5716 11174
rect 5656 11104 5661 11164
rect 5656 11094 5716 11104
rect 5671 11086 5701 11094
rect 5596 10753 5627 10757
rect 5581 10743 5641 10753
rect 5581 10683 5586 10743
rect 5581 10673 5641 10683
rect 5596 10660 5627 10673
rect 5597 8149 5627 10660
rect 5672 8292 5701 11086
rect 5747 10842 5777 11410
rect 5822 11258 5852 11410
rect 5807 11248 5867 11258
rect 5807 11188 5812 11248
rect 5807 11178 5867 11188
rect 5746 10838 5777 10842
rect 5731 10828 5791 10838
rect 5731 10768 5736 10828
rect 5731 10758 5791 10768
rect 5746 10745 5777 10758
rect 5747 8643 5777 10745
rect 5822 8768 5852 11178
rect 5897 10927 5927 11410
rect 5972 11342 6002 11410
rect 5957 11332 6017 11342
rect 5957 11272 5962 11332
rect 5957 11262 6017 11272
rect 5896 10923 5927 10927
rect 5881 10913 5941 10923
rect 5881 10853 5886 10913
rect 5881 10843 5941 10853
rect 5896 10783 5927 10843
rect 5897 9237 5927 10783
rect 5972 9343 6002 11262
rect 6047 11013 6077 11410
rect 6107 11356 6112 11416
rect 6107 11346 6167 11356
rect 6046 11008 6077 11013
rect 6031 10998 6091 11008
rect 6031 10938 6036 10998
rect 6031 10928 6091 10938
rect 6046 10920 6077 10928
rect 6047 9761 6077 10920
rect 6122 9906 6152 11346
rect 6107 9896 6167 9906
rect 6107 9836 6112 9896
rect 6107 9826 6167 9836
rect 6032 9751 6092 9761
rect 6032 9691 6037 9751
rect 6032 9681 6092 9691
rect 6107 9576 6167 9586
rect 6107 9516 6112 9576
rect 6107 9506 6167 9516
rect 6032 9448 6092 9458
rect 6032 9388 6037 9448
rect 6032 9378 6092 9388
rect 5957 9333 6017 9343
rect 5957 9273 5962 9333
rect 5957 9263 6017 9273
rect 5882 9227 5942 9237
rect 5882 9167 5887 9227
rect 5882 9157 5942 9167
rect 5957 9068 6017 9078
rect 5957 9008 5962 9068
rect 5957 8998 6017 9008
rect 5882 8914 5942 8924
rect 5882 8854 5887 8914
rect 5882 8844 5942 8854
rect 5807 8758 5867 8768
rect 5807 8698 5812 8758
rect 5807 8688 5867 8698
rect 5732 8633 5792 8643
rect 5732 8573 5737 8633
rect 5732 8563 5792 8573
rect 5807 8488 5867 8498
rect 5807 8428 5812 8488
rect 5807 8418 5867 8428
rect 5732 8381 5792 8391
rect 5732 8321 5737 8381
rect 5732 8311 5792 8321
rect 5672 8273 5702 8292
rect 5657 8263 5717 8273
rect 5657 8203 5662 8263
rect 5657 8193 5717 8203
rect 5582 8139 5642 8149
rect 5582 8079 5587 8139
rect 5582 8069 5642 8079
rect 5657 7980 5717 7990
rect 5657 7920 5662 7980
rect 5657 7910 5717 7920
rect 5582 7826 5642 7836
rect 5582 7766 5587 7826
rect 5582 7756 5642 7766
rect 5507 7670 5567 7680
rect 5507 7610 5512 7670
rect 5507 7600 5567 7610
rect 2550 7545 2610 7555
rect 2605 7485 2610 7545
rect 2550 7475 2610 7485
rect 5432 7545 5492 7555
rect 5432 7485 5437 7545
rect 5432 7475 5492 7485
rect 2475 7400 2535 7410
rect 2530 7340 2535 7400
rect 2475 7330 2535 7340
rect 5507 7400 5567 7410
rect 5507 7340 5512 7400
rect 5507 7330 5567 7340
rect 2490 6360 2520 7330
rect 2550 7293 2610 7303
rect 2605 7233 2610 7293
rect 5432 7293 5492 7303
rect 2550 7223 2610 7233
rect 2565 6360 2595 7223
rect 3760 7170 3770 7270
rect 3940 7170 3950 7270
rect 5432 7233 5437 7293
rect 5432 7223 5492 7233
rect 5447 7120 5477 7223
rect 2625 7090 5477 7120
rect 2625 6360 2655 7090
rect 5522 7060 5552 7330
rect 2685 7030 5552 7060
rect 2685 6360 2715 7030
rect 5597 7000 5627 7756
rect 2745 6975 5627 7000
rect 2745 6970 5626 6975
rect 2745 6360 2775 6970
rect 5672 6940 5702 7910
rect 2805 6910 5702 6940
rect 2805 6360 2835 6910
rect 5747 6880 5777 8311
rect 2865 6850 5777 6880
rect 2865 6360 2895 6850
rect 5822 6820 5852 8418
rect 2925 6790 5853 6820
rect 2925 6360 2955 6790
rect 5897 6760 5927 8844
rect 2985 6730 5927 6760
rect 2985 6360 3015 6730
rect 5972 6700 6002 8998
rect 3045 6670 6002 6700
rect 3045 6360 3075 6670
rect 6047 6640 6077 9378
rect 3105 6610 6077 6640
rect 3105 6360 3135 6610
rect 6122 6580 6152 9506
rect 3165 6550 6152 6580
rect 3165 6360 3195 6550
<< via1 >>
rect 1725 10379 1780 10439
rect 1800 10255 1855 10315
rect 1725 10096 1780 10156
rect 1800 9942 1855 10002
rect 1875 9786 1930 9846
rect 1950 9661 2005 9721
rect 1875 9516 1930 9576
rect 1950 9409 2005 9469
rect 2025 9291 2080 9351
rect 2100 9167 2155 9227
rect 2025 9008 2080 9068
rect 2100 8854 2155 8914
rect 2175 8698 2230 8758
rect 2250 8573 2305 8633
rect 2175 8428 2230 8488
rect 2250 8321 2305 8381
rect 2325 8203 2380 8263
rect 2400 8079 2455 8139
rect 2325 7920 2380 7980
rect 2400 7766 2455 7826
rect 2475 7610 2530 7670
rect 5511 11020 5566 11080
rect 5436 10598 5491 10658
rect 3770 10430 3940 10530
rect 4100 9890 4270 9990
rect 3770 9340 3940 9440
rect 4100 8800 4270 8900
rect 3770 8250 3940 8350
rect 4100 7710 4270 7810
rect 5661 11104 5716 11164
rect 5586 10683 5641 10743
rect 5812 11188 5867 11248
rect 5736 10768 5791 10828
rect 5962 11272 6017 11332
rect 5886 10853 5941 10913
rect 6112 11356 6167 11416
rect 6036 10938 6091 10998
rect 6112 9836 6167 9896
rect 6037 9691 6092 9751
rect 6112 9516 6167 9576
rect 6037 9388 6092 9448
rect 5962 9273 6017 9333
rect 5887 9167 5942 9227
rect 5962 9008 6017 9068
rect 5887 8854 5942 8914
rect 5812 8698 5867 8758
rect 5737 8573 5792 8633
rect 5812 8428 5867 8488
rect 5737 8321 5792 8381
rect 5662 8203 5717 8263
rect 5587 8079 5642 8139
rect 5662 7920 5717 7980
rect 5587 7766 5642 7826
rect 5512 7610 5567 7670
rect 2550 7485 2605 7545
rect 5437 7485 5492 7545
rect 2475 7340 2530 7400
rect 5512 7340 5567 7400
rect 2550 7233 2605 7293
rect 3770 7170 3940 7270
rect 5437 7233 5492 7293
<< metal2 >>
rect 1920 10642 1950 11600
rect 1980 10727 2010 11600
rect 2040 10812 2070 11600
rect 2100 10897 2130 11600
rect 2160 10982 2190 11600
rect 2220 11064 2250 11600
rect 2280 11146 2310 11600
rect 2340 11232 2370 11600
rect 2400 11316 2430 11600
rect 2460 11400 2490 11600
rect 6107 11416 6167 11426
rect 6107 11400 6112 11416
rect 2460 11370 6112 11400
rect 6107 11356 6112 11370
rect 6107 11346 6167 11356
rect 5957 11332 6017 11342
rect 5957 11316 5962 11332
rect 2400 11286 5962 11316
rect 5957 11272 5962 11286
rect 5957 11262 6017 11272
rect 5807 11248 5867 11258
rect 5807 11232 5812 11248
rect 2340 11202 5812 11232
rect 5807 11188 5812 11202
rect 5807 11178 5867 11188
rect 5656 11164 5716 11174
rect 5656 11148 5661 11164
rect 5633 11146 5661 11148
rect 2280 11118 5661 11146
rect 5656 11104 5661 11118
rect 5656 11094 5716 11104
rect 5506 11080 5566 11090
rect 5506 11064 5511 11080
rect 2220 11033 5511 11064
rect 5506 11020 5511 11033
rect 5506 11010 5566 11020
rect 6031 10998 6091 11008
rect 6031 10982 6036 10998
rect 2160 10951 6036 10982
rect 6031 10938 6036 10951
rect 6031 10928 6091 10938
rect 5881 10913 5941 10923
rect 5881 10897 5886 10913
rect 2100 10866 5886 10897
rect 5881 10853 5886 10866
rect 5881 10843 5941 10853
rect 5731 10828 5791 10838
rect 5731 10812 5736 10828
rect 2040 10781 5736 10812
rect 5731 10768 5736 10781
rect 5731 10758 5791 10768
rect 5581 10743 5641 10753
rect 5581 10727 5586 10743
rect 1980 10696 5586 10727
rect 5581 10683 5586 10696
rect 5581 10673 5641 10683
rect 5431 10658 5491 10668
rect 5431 10642 5436 10658
rect 1920 10611 5436 10642
rect 5431 10598 5436 10611
rect 5431 10588 5491 10598
rect 3770 10530 3940 10540
rect 1725 10439 1785 10449
rect 1780 10421 1785 10439
rect 1780 10391 2640 10421
rect 1780 10379 1785 10391
rect 1725 10369 1785 10379
rect 1800 10315 1860 10325
rect 1855 10297 1860 10315
rect 1855 10267 2640 10297
rect 1855 10255 1860 10267
rect 1800 10245 1860 10255
rect 1725 10156 1785 10166
rect 1780 10143 1785 10156
rect 1780 10113 2640 10143
rect 1780 10096 1785 10113
rect 1725 10086 1785 10096
rect 1800 10002 1860 10012
rect 1855 9990 1860 10002
rect 1855 9960 2640 9990
rect 1855 9942 1860 9960
rect 1800 9932 1860 9942
rect 1875 9846 1935 9856
rect 1930 9828 1935 9846
rect 1930 9798 2640 9828
rect 1930 9786 1935 9798
rect 1875 9776 1935 9786
rect 1950 9721 2010 9731
rect 2005 9703 2010 9721
rect 2005 9673 2640 9703
rect 2005 9661 2010 9673
rect 1950 9651 2010 9661
rect 1875 9576 1935 9586
rect 1930 9563 1935 9576
rect 1930 9533 2640 9563
rect 1930 9516 1935 9533
rect 1875 9506 1935 9516
rect 1950 9469 2010 9479
rect 2005 9463 2010 9469
rect 2005 9433 2640 9463
rect 3770 9440 3940 10430
rect 2005 9409 2010 9433
rect 1950 9399 2010 9409
rect 2025 9351 2085 9361
rect 2080 9333 2085 9351
rect 2080 9303 2640 9333
rect 2080 9291 2085 9303
rect 2025 9281 2085 9291
rect 2100 9227 2160 9237
rect 2155 9209 2160 9227
rect 2155 9179 2640 9209
rect 2155 9167 2160 9179
rect 2100 9157 2160 9167
rect 2025 9068 2085 9078
rect 2080 9055 2085 9068
rect 2080 9025 2640 9055
rect 2080 9008 2085 9025
rect 2025 8998 2085 9008
rect 2100 8914 2160 8924
rect 2155 8902 2160 8914
rect 2155 8872 2640 8902
rect 2155 8854 2160 8872
rect 2100 8844 2160 8854
rect 2175 8758 2235 8768
rect 2230 8740 2235 8758
rect 2230 8710 2640 8740
rect 2230 8698 2235 8710
rect 2175 8688 2235 8698
rect 2250 8633 2310 8643
rect 2305 8615 2310 8633
rect 2305 8585 2640 8615
rect 2305 8573 2310 8585
rect 2250 8563 2310 8573
rect 2175 8488 2235 8498
rect 2230 8475 2235 8488
rect 2230 8445 2640 8475
rect 2230 8428 2235 8445
rect 2175 8418 2235 8428
rect 2250 8381 2310 8391
rect 2305 8375 2310 8381
rect 2305 8345 2640 8375
rect 3770 8350 3940 9340
rect 2305 8321 2310 8345
rect 2250 8311 2310 8321
rect 2325 8263 2385 8273
rect 2380 8245 2385 8263
rect 2380 8215 2640 8245
rect 2380 8203 2385 8215
rect 2325 8193 2385 8203
rect 2400 8139 2460 8149
rect 2455 8121 2460 8139
rect 2455 8091 2640 8121
rect 2455 8079 2460 8091
rect 2400 8069 2460 8079
rect 2325 7980 2385 7990
rect 2380 7967 2385 7980
rect 2380 7937 2640 7967
rect 2380 7920 2385 7937
rect 2325 7910 2385 7920
rect 2400 7826 2460 7836
rect 2455 7814 2460 7826
rect 2455 7784 2640 7814
rect 2455 7766 2460 7784
rect 2400 7756 2460 7766
rect 2475 7670 2535 7680
rect 2530 7652 2535 7670
rect 2530 7622 2640 7652
rect 2530 7610 2535 7622
rect 2475 7600 2535 7610
rect 2550 7545 2610 7555
rect 2605 7527 2610 7545
rect 2605 7497 2640 7527
rect 2605 7485 2610 7497
rect 2550 7475 2610 7485
rect 2475 7400 2535 7410
rect 2530 7387 2535 7400
rect 2530 7357 2640 7387
rect 2530 7340 2535 7357
rect 2475 7330 2535 7340
rect 2550 7293 2610 7303
rect 2605 7287 2610 7293
rect 2605 7257 2640 7287
rect 3770 7270 3940 8250
rect 4100 9990 4270 10000
rect 4100 8900 4270 9890
rect 6107 9896 6167 9906
rect 6107 9878 6112 9896
rect 5400 9848 6112 9878
rect 6107 9836 6112 9848
rect 6107 9826 6167 9836
rect 6032 9751 6092 9761
rect 6032 9733 6037 9751
rect 5400 9703 6037 9733
rect 6032 9691 6037 9703
rect 6032 9681 6092 9691
rect 6107 9576 6167 9586
rect 6107 9563 6112 9576
rect 5400 9533 6112 9563
rect 6107 9516 6112 9533
rect 6107 9506 6167 9516
rect 6032 9448 6092 9458
rect 6032 9408 6037 9448
rect 5400 9388 6037 9408
rect 5400 9378 6092 9388
rect 5957 9333 6017 9343
rect 5400 9303 5962 9333
rect 5957 9273 5962 9303
rect 5957 9263 6017 9273
rect 5882 9227 5942 9237
rect 5882 9209 5887 9227
rect 5400 9179 5887 9209
rect 5882 9167 5887 9179
rect 5882 9157 5942 9167
rect 5957 9068 6017 9078
rect 5957 9055 5962 9068
rect 5400 9025 5962 9055
rect 5957 9008 5962 9025
rect 5957 8998 6017 9008
rect 5882 8914 5942 8924
rect 5882 8902 5887 8914
rect 5400 8872 5887 8902
rect 5882 8854 5887 8872
rect 5882 8844 5942 8854
rect 4100 7810 4270 8800
rect 5807 8758 5867 8768
rect 5807 8740 5812 8758
rect 5400 8710 5812 8740
rect 5807 8698 5812 8710
rect 5807 8688 5867 8698
rect 5732 8633 5792 8643
rect 5732 8615 5737 8633
rect 5400 8585 5737 8615
rect 5732 8573 5737 8585
rect 5732 8563 5792 8573
rect 5807 8488 5867 8498
rect 5807 8475 5812 8488
rect 5400 8445 5812 8475
rect 5807 8428 5812 8445
rect 5807 8418 5867 8428
rect 5732 8381 5792 8391
rect 5732 8375 5737 8381
rect 5400 8345 5737 8375
rect 5732 8321 5737 8345
rect 5732 8311 5792 8321
rect 5657 8263 5717 8273
rect 5657 8245 5662 8263
rect 5400 8215 5662 8245
rect 5657 8203 5662 8215
rect 5657 8193 5717 8203
rect 5582 8139 5642 8149
rect 5582 8121 5587 8139
rect 5400 8091 5587 8121
rect 5582 8079 5587 8091
rect 5582 8069 5642 8079
rect 5657 7980 5717 7990
rect 5657 7967 5662 7980
rect 5400 7937 5662 7967
rect 5657 7920 5662 7937
rect 5657 7910 5717 7920
rect 5582 7826 5642 7836
rect 5582 7814 5587 7826
rect 5400 7784 5587 7814
rect 5582 7766 5587 7784
rect 5582 7756 5642 7766
rect 4100 7700 4270 7710
rect 5507 7670 5567 7680
rect 5507 7652 5512 7670
rect 5400 7622 5512 7652
rect 5507 7610 5512 7622
rect 5507 7600 5567 7610
rect 5432 7545 5492 7555
rect 5432 7527 5437 7545
rect 5400 7497 5437 7527
rect 5432 7485 5437 7497
rect 5432 7475 5492 7485
rect 5507 7400 5567 7410
rect 5507 7387 5512 7400
rect 5400 7357 5512 7387
rect 5507 7340 5512 7357
rect 5507 7330 5567 7340
rect 5432 7293 5492 7303
rect 5432 7287 5437 7293
rect 2605 7233 2610 7257
rect 2550 7223 2610 7233
rect 5400 7257 5437 7287
rect 5432 7233 5437 7257
rect 5432 7223 5492 7233
rect 3770 7160 3940 7170
use bbm_unit  bbm_unit_0
timestamp 1713724235
transform -1 0 4607 0 1 9363
box -890 -20 626 620
use bbm_unit_x2  bbm_unit_x2_0
array 0 0 1516 0 2 1088
timestamp 1713891259
transform 1 0 3431 0 1 7187
box -890 -20 626 1164
use bbm_unit_x2  bbm_unit_x2_3
array 0 0 1516 0 1 1088
timestamp 1713891259
transform -1 0 4607 0 1 7187
box -890 -20 626 1164
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 5123 0 -1 10479
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1710522493
transform 1 0 4019 0 -1 10479
box -38 -48 1142 592
<< end >>
