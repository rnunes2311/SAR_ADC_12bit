magic
tech sky130A
timestamp 1712086620
<< metal1 >>
rect 755 270 760 300
rect 790 270 795 300
rect 755 260 795 270
rect 755 240 920 260
rect 755 230 795 240
rect 755 200 760 230
rect 790 200 795 230
<< via1 >>
rect 760 270 790 300
rect 760 200 790 230
<< metal2 >>
rect 755 300 795 305
rect 755 270 760 300
rect 790 270 795 300
rect 755 230 795 270
rect 755 200 760 230
rect 790 200 795 230
rect 755 195 795 200
<< via2 >>
rect 760 270 790 300
rect 760 200 790 230
<< metal3 >>
rect 750 300 920 320
rect 750 270 760 300
rect 790 270 920 300
rect 750 230 920 270
rect 750 200 760 230
rect 790 200 920 230
rect 750 180 920 200
<< mimcap >>
rect 800 290 900 300
rect 800 210 810 290
rect 890 210 900 290
rect 800 200 900 210
<< mimcapcontact >>
rect 810 210 890 290
<< metal4 >>
rect 835 300 865 345
rect 800 290 900 300
rect 800 210 810 290
rect 890 210 900 290
rect 800 200 900 210
rect 835 160 865 200
<< end >>
